GEN|1|1|in principio creavit Deus caelum et terram
GEN|1|2|terra autem erat inanis et vacua et tenebrae super faciem abyssi et spiritus Dei ferebatur super aquas
GEN|1|3|dixitque Deus fiat lux et facta est lux
GEN|1|4|et vidit Deus lucem quod esset bona et divisit lucem ac tenebras
GEN|1|5|appellavitque lucem diem et tenebras noctem factumque est vespere et mane dies unus
GEN|1|6|dixit quoque Deus fiat firmamentum in medio aquarum et dividat aquas ab aquis
GEN|1|7|et fecit Deus firmamentum divisitque aquas quae erant sub firmamento ab his quae erant super firmamentum et factum est ita
GEN|1|8|vocavitque Deus firmamentum caelum et factum est vespere et mane dies secundus
GEN|1|9|dixit vero Deus congregentur aquae quae sub caelo sunt in locum unum et appareat arida factumque est ita
GEN|1|10|et vocavit Deus aridam terram congregationesque aquarum appellavit maria et vidit Deus quod esset bonum
GEN|1|11|et ait germinet terra herbam virentem et facientem semen et lignum pomiferum faciens fructum iuxta genus suum cuius semen in semet ipso sit super terram et factum est ita
GEN|1|12|et protulit terra herbam virentem et adferentem semen iuxta genus suum lignumque faciens fructum et habens unumquodque sementem secundum speciem suam et vidit Deus quod esset bonum
GEN|1|13|factumque est vespere et mane dies tertius
GEN|1|14|dixit autem Deus fiant luminaria in firmamento caeli ut dividant diem ac noctem et sint in signa et tempora et dies et annos
GEN|1|15|ut luceant in firmamento caeli et inluminent terram et factum est ita
GEN|1|16|fecitque Deus duo magna luminaria luminare maius ut praeesset diei et luminare minus ut praeesset nocti et stellas
GEN|1|17|et posuit eas in firmamento caeli ut lucerent super terram
GEN|1|18|et praeessent diei ac nocti et dividerent lucem ac tenebras et vidit Deus quod esset bonum
GEN|1|19|et factum est vespere et mane dies quartus
GEN|1|20|dixit etiam Deus producant aquae reptile animae viventis et volatile super terram sub firmamento caeli
GEN|1|21|creavitque Deus cete grandia et omnem animam viventem atque motabilem quam produxerant aquae in species suas et omne volatile secundum genus suum et vidit Deus quod esset bonum
GEN|1|22|benedixitque eis dicens crescite et multiplicamini et replete aquas maris avesque multiplicentur super terram
GEN|1|23|et factum est vespere et mane dies quintus
GEN|1|24|dixit quoque Deus producat terra animam viventem in genere suo iumenta et reptilia et bestias terrae secundum species suas factumque est ita
GEN|1|25|et fecit Deus bestias terrae iuxta species suas et iumenta et omne reptile terrae in genere suo et vidit Deus quod esset bonum
GEN|1|26|et ait faciamus hominem ad imaginem et similitudinem nostram et praesit piscibus maris et volatilibus caeli et bestiis universaeque terrae omnique reptili quod movetur in terra
GEN|1|27|et creavit Deus hominem ad imaginem suam ad imaginem Dei creavit illum masculum et feminam creavit eos
GEN|1|28|benedixitque illis Deus et ait crescite et multiplicamini et replete terram et subicite eam et dominamini piscibus maris et volatilibus caeli et universis animantibus quae moventur super terram
GEN|1|29|dixitque Deus ecce dedi vobis omnem herbam adferentem semen super terram et universa ligna quae habent in semet ipsis sementem generis sui ut sint vobis in escam
GEN|1|30|et cunctis animantibus terrae omnique volucri caeli et universis quae moventur in terra et in quibus est anima vivens ut habeant ad vescendum et factum est ita
GEN|1|31|viditque Deus cuncta quae fecit et erant valde bona et factum est vespere et mane dies sextus
GEN|2|1|igitur perfecti sunt caeli et terra et omnis ornatus eorum
GEN|2|2|conplevitque Deus die septimo opus suum quod fecerat et requievit die septimo ab universo opere quod patrarat
GEN|2|3|et benedixit diei septimo et sanctificavit illum quia in ipso cessaverat ab omni opere suo quod creavit Deus ut faceret
GEN|2|4|istae generationes caeli et terrae quando creatae sunt in die quo fecit Dominus Deus caelum et terram
GEN|2|5|et omne virgultum agri antequam oreretur in terra omnemque herbam regionis priusquam germinaret non enim pluerat Dominus Deus super terram et homo non erat qui operaretur terram
GEN|2|6|sed fons ascendebat e terra inrigans universam superficiem terrae
GEN|2|7|formavit igitur Dominus Deus hominem de limo terrae et inspiravit in faciem eius spiraculum vitae et factus est homo in animam viventem
GEN|2|8|plantaverat autem Dominus Deus paradisum voluptatis a principio in quo posuit hominem quem formaverat
GEN|2|9|produxitque Dominus Deus de humo omne lignum pulchrum visu et ad vescendum suave lignum etiam vitae in medio paradisi lignumque scientiae boni et mali
GEN|2|10|et fluvius egrediebatur de loco voluptatis ad inrigandum paradisum qui inde dividitur in quattuor capita
GEN|2|11|nomen uni Phison ipse est qui circuit omnem terram Evilat ubi nascitur aurum
GEN|2|12|et aurum terrae illius optimum est ibique invenitur bdellium et lapis onychinus
GEN|2|13|et nomen fluvio secundo Geon ipse est qui circuit omnem terram Aethiopiae
GEN|2|14|nomen vero fluminis tertii Tigris ipse vadit contra Assyrios fluvius autem quartus ipse est Eufrates
GEN|2|15|tulit ergo Dominus Deus hominem et posuit eum in paradiso voluptatis ut operaretur et custodiret illum
GEN|2|16|praecepitque ei dicens ex omni ligno paradisi comede
GEN|2|17|de ligno autem scientiae boni et mali ne comedas in quocumque enim die comederis ex eo morte morieris
GEN|2|18|dixit quoque Dominus Deus non est bonum esse hominem solum faciamus ei adiutorium similem sui
GEN|2|19|formatis igitur Dominus Deus de humo cunctis animantibus terrae et universis volatilibus caeli adduxit ea ad Adam ut videret quid vocaret ea omne enim quod vocavit Adam animae viventis ipsum est nomen eius
GEN|2|20|appellavitque Adam nominibus suis cuncta animantia et universa volatilia caeli et omnes bestias terrae Adam vero non inveniebatur adiutor similis eius
GEN|2|21|inmisit ergo Dominus Deus soporem in Adam cumque obdormisset tulit unam de costis eius et replevit carnem pro ea
GEN|2|22|et aedificavit Dominus Deus costam quam tulerat de Adam in mulierem et adduxit eam ad Adam
GEN|2|23|dixitque Adam hoc nunc os ex ossibus meis et caro de carne mea haec vocabitur virago quoniam de viro sumpta est
GEN|2|24|quam ob rem relinquet homo patrem suum et matrem et adherebit uxori suae et erunt duo in carne una
GEN|2|25|erant autem uterque nudi Adam scilicet et uxor eius et non erubescebant
GEN|3|1|sed et serpens erat callidior cunctis animantibus terrae quae fecerat Dominus Deus qui dixit ad mulierem cur praecepit vobis Deus ut non comederetis de omni ligno paradisi
GEN|3|2|cui respondit mulier de fructu lignorum quae sunt in paradiso vescemur
GEN|3|3|de fructu vero ligni quod est in medio paradisi praecepit nobis Deus ne comederemus et ne tangeremus illud ne forte moriamur
GEN|3|4|dixit autem serpens ad mulierem nequaquam morte moriemini
GEN|3|5|scit enim Deus quod in quocumque die comederitis ex eo aperientur oculi vestri et eritis sicut dii scientes bonum et malum
GEN|3|6|vidit igitur mulier quod bonum esset lignum ad vescendum et pulchrum oculis aspectuque delectabile et tulit de fructu illius et comedit deditque viro suo qui comedit
GEN|3|7|et aperti sunt oculi amborum cumque cognovissent esse se nudos consuerunt folia ficus et fecerunt sibi perizomata
GEN|3|8|et cum audissent vocem Domini Dei deambulantis in paradiso ad auram post meridiem abscondit se Adam et uxor eius a facie Domini Dei in medio ligni paradisi
GEN|3|9|vocavitque Dominus Deus Adam et dixit ei ubi es
GEN|3|10|qui ait vocem tuam audivi in paradiso et timui eo quod nudus essem et abscondi me
GEN|3|11|cui dixit quis enim indicavit tibi quod nudus esses nisi quod ex ligno de quo tibi praeceperam ne comederes comedisti
GEN|3|12|dixitque Adam mulier quam dedisti sociam mihi dedit mihi de ligno et comedi
GEN|3|13|et dixit Dominus Deus ad mulierem quare hoc fecisti quae respondit serpens decepit me et comedi
GEN|3|14|et ait Dominus Deus ad serpentem quia fecisti hoc maledictus es inter omnia animantia et bestias terrae super pectus tuum gradieris et terram comedes cunctis diebus vitae tuae
GEN|3|15|inimicitias ponam inter te et mulierem et semen tuum et semen illius ipsa conteret caput tuum et tu insidiaberis calcaneo eius
GEN|3|16|mulieri quoque dixit multiplicabo aerumnas tuas et conceptus tuos in dolore paries filios et sub viri potestate eris et ipse dominabitur tui
GEN|3|17|ad Adam vero dixit quia audisti vocem uxoris tuae et comedisti de ligno ex quo praeceperam tibi ne comederes maledicta terra in opere tuo in laboribus comedes eam cunctis diebus vitae tuae
GEN|3|18|spinas et tribulos germinabit tibi et comedes herbas terrae
GEN|3|19|in sudore vultus tui vesceris pane donec revertaris in terram de qua sumptus es quia pulvis es et in pulverem reverteris
GEN|3|20|et vocavit Adam nomen uxoris suae Hava eo quod mater esset cunctorum viventium
GEN|3|21|fecit quoque Dominus Deus Adam et uxori eius tunicas pellicias et induit eos
GEN|3|22|et ait ecce Adam factus est quasi unus ex nobis sciens bonum et malum nunc ergo ne forte mittat manum suam et sumat etiam de ligno vitae et comedat et vivat in aeternum
GEN|3|23|emisit eum Dominus Deus de paradiso voluptatis ut operaretur terram de qua sumptus est
GEN|3|24|eiecitque Adam et conlocavit ante paradisum voluptatis cherubin et flammeum gladium atque versatilem ad custodiendam viam ligni vitae
GEN|4|1|Adam vero cognovit Havam uxorem suam quae concepit et peperit Cain dicens possedi hominem per Dominum
GEN|4|2|rursusque peperit fratrem eius Abel fuit autem Abel pastor ovium et Cain agricola
GEN|4|3|factum est autem post multos dies ut offerret Cain de fructibus terrae munera Domino
GEN|4|4|Abel quoque obtulit de primogenitis gregis sui et de adipibus eorum et respexit Dominus ad Abel et ad munera eius
GEN|4|5|ad Cain vero et ad munera illius non respexit iratusque est Cain vehementer et concidit vultus eius
GEN|4|6|dixitque Dominus ad eum quare maestus es et cur concidit facies tua
GEN|4|7|nonne si bene egeris recipies sin autem male statim in foribus peccatum aderit sed sub te erit appetitus eius et tu dominaberis illius
GEN|4|8|dixitque Cain ad Abel fratrem suum egrediamur foras cumque essent in agro consurrexit Cain adversus Abel fratrem suum et interfecit eum
GEN|4|9|et ait Dominus ad Cain ubi est Abel frater tuus qui respondit nescio num custos fratris mei sum
GEN|4|10|dixitque ad eum quid fecisti vox sanguinis fratris tui clamat ad me de terra
GEN|4|11|nunc igitur maledictus eris super terram quae aperuit os suum et suscepit sanguinem fratris tui de manu tua
GEN|4|12|cum operatus fueris eam non dabit tibi fructus suos vagus et profugus eris super terram
GEN|4|13|dixitque Cain ad Dominum maior est iniquitas mea quam ut veniam merear
GEN|4|14|ecce eicis me hodie a facie terrae et a facie tua abscondar et ero vagus et profugus in terra omnis igitur qui invenerit me occidet me
GEN|4|15|dixitque ei Dominus nequaquam ita fiet sed omnis qui occiderit Cain septuplum punietur posuitque Dominus Cain signum ut non eum interficeret omnis qui invenisset eum
GEN|4|16|egressusque Cain a facie Domini habitavit in terra profugus ad orientalem plagam Eden
GEN|4|17|cognovit autem Cain uxorem suam quae concepit et peperit Enoch et aedificavit civitatem vocavitque nomen eius ex nomine filii sui Enoch
GEN|4|18|porro Enoch genuit Irad et Irad genuit Maviahel et Maviahel genuit Matusahel et Matusahel genuit Lamech
GEN|4|19|qui accepit uxores duas nomen uni Ada et nomen alteri Sella
GEN|4|20|genuitque Ada Iabel qui fuit pater habitantium in tentoriis atque pastorum
GEN|4|21|et nomen fratris eius Iubal ipse fuit pater canentium cithara et organo
GEN|4|22|Sella quoque genuit Thubalcain qui fuit malleator et faber in cuncta opera aeris et ferri soror vero Thubalcain Noemma
GEN|4|23|dixitque Lamech uxoribus suis Adae et Sellae audite vocem meam uxores Lamech auscultate sermonem meum quoniam occidi virum in vulnus meum et adulescentulum in livorem meum
GEN|4|24|septuplum ultio dabitur de Cain de Lamech vero septuagies septies
GEN|4|25|cognovit quoque adhuc Adam uxorem suam et peperit filium vocavitque nomen eius Seth dicens posuit mihi Deus semen aliud pro Abel quem occidit Cain
GEN|4|26|sed et Seth natus est filius quem vocavit Enos iste coepit invocare nomen Domini
GEN|5|1|hic est liber generationis Adam in die qua creavit Deus hominem ad similitudinem Dei fecit illum
GEN|5|2|masculum et feminam creavit eos et benedixit illis et vocavit nomen eorum Adam in die qua creati sunt
GEN|5|3|vixit autem Adam centum triginta annis et genuit ad similitudinem et imaginem suam vocavitque nomen eius Seth
GEN|5|4|et facti sunt dies Adam postquam genuit Seth octingenti anni genuitque filios et filias
GEN|5|5|et factum est omne tempus quod vixit Adam anni nongenti triginta et mortuus est
GEN|5|6|vixit quoque Seth centum quinque annos et genuit Enos
GEN|5|7|vixitque Seth postquam genuit Enos octingentis septem annis genuitque filios et filias
GEN|5|8|et facti sunt omnes dies Seth nongentorum duodecim annorum et mortuus est
GEN|5|9|vixit vero Enos nonaginta annis et genuit Cainan
GEN|5|10|post cuius ortum vixit octingentis quindecim annis et genuit filios et filias
GEN|5|11|factique sunt omnes dies Enos nongentorum quinque annorum et mortuus est
GEN|5|12|vixit quoque Cainan septuaginta annis et genuit Malalehel
GEN|5|13|et vixit Cainan postquam genuit Malalehel octingentos quadraginta annos genuitque filios et filias
GEN|5|14|et facti sunt omnes dies Cainan nongenti decem anni et mortuus est
GEN|5|15|vixit autem Malalehel sexaginta quinque annos et genuit Iared
GEN|5|16|et vixit Malalehel postquam genuit Iared octingentis triginta annis et genuit filios et filias
GEN|5|17|et facti sunt omnes dies Malalehel octingenti nonaginta quinque anni et mortuus est
GEN|5|18|vixitque Iared centum sexaginta duobus annis et genuit Enoch
GEN|5|19|et vixit Iared postquam genuit Enoch octingentos annos et genuit filios et filias
GEN|5|20|et facti sunt omnes dies Iared nongenti sexaginta duo anni et mortuus est
GEN|5|21|porro Enoch vixit sexaginta quinque annis et genuit Mathusalam
GEN|5|22|et ambulavit Enoch cum Deo postquam genuit Mathusalam trecentis annis et genuit filios et filias
GEN|5|23|et facti sunt omnes dies Enoch trecenti sexaginta quinque anni
GEN|5|24|ambulavitque cum Deo et non apparuit quia tulit eum Deus
GEN|5|25|vixit quoque Mathusalam centum octoginta septem annos et genuit Lamech
GEN|5|26|et vixit Mathusalam postquam genuit Lamech septingentos octoginta duos annos et genuit filios et filias
GEN|5|27|et facti sunt omnes dies Mathusalae nongenti sexaginta novem anni et mortuus est
GEN|5|28|vixit autem Lamech centum octoginta duobus annis et genuit filium
GEN|5|29|vocavitque nomen eius Noe dicens iste consolabitur nos ab operibus et laboribus manuum nostrarum in terra cui maledixit Dominus
GEN|5|30|vixitque Lamech postquam genuit Noe quingentos nonaginta quinque annos et genuit filios et filias
GEN|5|31|et facti sunt omnes dies Lamech septingenti septuaginta septem anni et mortuus est
GEN|5|32|Noe vero cum quingentorum esset annorum genuit Sem et Ham et Iafeth
GEN|6|1|cumque coepissent homines multiplicari super terram et filias procreassent
GEN|6|2|videntes filii Dei filias eorum quod essent pulchrae acceperunt uxores sibi ex omnibus quas elegerant
GEN|6|3|dixitque Deus non permanebit spiritus meus in homine in aeternum quia caro est eruntque dies illius centum viginti annorum
GEN|6|4|gigantes autem erant super terram in diebus illis postquam enim ingressi sunt filii Dei ad filias hominum illaeque genuerunt isti sunt potentes a saeculo viri famosi
GEN|6|5|videns autem Deus quod multa malitia hominum esset in terra et cuncta cogitatio cordis intenta esset ad malum omni tempore
GEN|6|6|paenituit eum quod hominem fecisset in terra et tactus dolore cordis intrinsecus
GEN|6|7|delebo inquit hominem quem creavi a facie terrae ab homine usque ad animantia a reptili usque ad volucres caeli paenitet enim me fecisse eos
GEN|6|8|Noe vero invenit gratiam coram Domino
GEN|6|9|hae generationes Noe Noe vir iustus atque perfectus fuit in generationibus suis cum Deo ambulavit
GEN|6|10|et genuit tres filios Sem Ham et Iafeth
GEN|6|11|corrupta est autem terra coram Deo et repleta est iniquitate
GEN|6|12|cumque vidisset Deus terram esse corruptam omnis quippe caro corruperat viam suam super terram
GEN|6|13|dixit ad Noe finis universae carnis venit coram me repleta est terra iniquitate a facie eorum et ego disperdam eos cum terra
GEN|6|14|fac tibi arcam de lignis levigatis mansiunculas in arca facies et bitumine linies intrinsecus et extrinsecus
GEN|6|15|et sic facies eam trecentorum cubitorum erit longitudo arcae quinquaginta cubitorum latitudo et triginta cubitorum altitudo illius
GEN|6|16|fenestram in arca facies et in cubito consummabis summitatem ostium autem arcae pones ex latere deorsum cenacula et tristega facies in ea
GEN|6|17|ecce ego adducam diluvii aquas super terram ut interficiam omnem carnem in qua spiritus vitae est subter caelum universa quae in terra sunt consumentur
GEN|6|18|ponamque foedus meum tecum et ingredieris arcam tu et filii tui uxor tua et uxores filiorum tuorum tecum
GEN|6|19|et ex cunctis animantibus universae carnis bina induces in arcam ut vivant tecum masculini sexus et feminini
GEN|6|20|de volucribus iuxta genus suum et de iumentis in genere suo et ex omni reptili terrae secundum genus suum bina de omnibus ingredientur tecum ut possint vivere
GEN|6|21|tolles igitur tecum ex omnibus escis quae mandi possunt et conportabis apud te et erunt tam tibi quam illis in cibum
GEN|6|22|fecit ergo Noe omnia quae praeceperat illi Deus
GEN|7|1|dixitque Dominus ad eum ingredere tu et omnis domus tua arcam te enim vidi iustum coram me in generatione hac
GEN|7|2|ex omnibus animantibus mundis tolle septena septena masculum et feminam de animantibus vero non mundis duo duo masculum et feminam
GEN|7|3|sed et de volatilibus caeli septena septena masculum et feminam ut salvetur semen super faciem universae terrae
GEN|7|4|adhuc enim et post dies septem ego pluam super terram quadraginta diebus et quadraginta noctibus et delebo omnem substantiam quam feci de superficie terrae
GEN|7|5|fecit ergo Noe omnia quae mandaverat ei Dominus
GEN|7|6|eratque sescentorum annorum quando diluvii aquae inundaverunt super terram
GEN|7|7|et ingressus est Noe et filii eius uxor eius et uxores filiorum eius cum eo in arcam propter aquas diluvii
GEN|7|8|de animantibus quoque mundis et inmundis et de volucribus et ex omni quod movetur super terram
GEN|7|9|duo et duo ingressa sunt ad Noe in arcam masculus et femina sicut praeceperat Deus Noe
GEN|7|10|cumque transissent septem dies aquae diluvii inundaverunt super terram
GEN|7|11|anno sescentesimo vitae Noe mense secundo septimodecimo die mensis rupti sunt omnes fontes abyssi magnae et cataractae caeli apertae sunt
GEN|7|12|et facta est pluvia super terram quadraginta diebus et quadraginta noctibus
GEN|7|13|in articulo diei illius ingressus est Noe et Sem et Ham et Iafeth filii eius uxor illius et tres uxores filiorum eius cum eis in arcam
GEN|7|14|ipsi et omne animal secundum genus suum universaque iumenta in genus suum et omne quod movetur super terram in genere suo cunctumque volatile secundum genus suum universae aves omnesque volucres
GEN|7|15|ingressae sunt ad Noe in arcam bina et bina ex omni carne in qua erat spiritus vitae
GEN|7|16|et quae ingressa sunt masculus et femina ex omni carne introierunt sicut praeceperat ei Deus et inclusit eum Dominus de foris
GEN|7|17|factumque est diluvium quadraginta diebus super terram et multiplicatae sunt aquae et elevaverunt arcam in sublime a terra
GEN|7|18|vehementer inundaverunt et omnia repleverunt in superficie terrae porro arca ferebatur super aquas
GEN|7|19|et aquae praevaluerunt nimis super terram opertique sunt omnes montes excelsi sub universo caelo
GEN|7|20|quindecim cubitis altior fuit aqua super montes quos operuerat
GEN|7|21|consumptaque est omnis caro quae movebatur super terram volucrum animantium bestiarum omniumque reptilium quae reptant super terram universi homines
GEN|7|22|et cuncta in quibus spiraculum vitae est in terra mortua sunt
GEN|7|23|et delevit omnem substantiam quae erat super terram ab homine usque ad pecus tam reptile quam volucres caeli et deleta sunt de terra remansit autem solus Noe et qui cum eo erant in arca
GEN|7|24|obtinueruntque aquae terras centum quinquaginta diebus
GEN|8|1|recordatus autem Deus Noe cunctarumque animantium et omnium iumentorum quae erant cum eo in arca adduxit spiritum super terram et inminutae sunt aquae
GEN|8|2|et clausi sunt fontes abyssi et cataractae caeli et prohibitae sunt pluviae de caelo
GEN|8|3|reversaeque aquae de terra euntes et redeuntes et coeperunt minui post centum quinquaginta dies
GEN|8|4|requievitque arca mense septimo vicesima septima die mensis super montes Armeniae
GEN|8|5|at vero aquae ibant et decrescebant usque ad decimum mensem decimo enim mense prima die mensis apparuerunt cacumina montium
GEN|8|6|cumque transissent quadraginta dies aperiens Noe fenestram arcae quam fecerat dimisit corvum
GEN|8|7|qui egrediebatur et revertebatur donec siccarentur aquae super terram
GEN|8|8|emisit quoque columbam post eum ut videret si iam cessassent aquae super faciem terrae
GEN|8|9|quae cum non invenisset ubi requiesceret pes eius reversa est ad eum in arcam aquae enim erant super universam terram extenditque manum et adprehensam intulit in arcam
GEN|8|10|expectatis autem ultra septem diebus aliis rursum dimisit columbam ex arca
GEN|8|11|at illa venit ad eum ad vesperam portans ramum olivae virentibus foliis in ore suo intellexit ergo Noe quod cessassent aquae super terram
GEN|8|12|expectavitque nihilominus septem alios dies et emisit columbam quae non est reversa ultra ad eum
GEN|8|13|igitur sescentesimo primo anno primo mense prima die mensis inminutae sunt aquae super terram et aperiens Noe tectum arcae aspexit viditque quod exsiccata esset superficies terrae
GEN|8|14|mense secundo septima et vicesima die mensis arefacta est terra
GEN|8|15|locutus est autem Deus ad Noe dicens
GEN|8|16|egredere de arca tu et uxor tua filii tui et uxores filiorum tuorum tecum
GEN|8|17|cuncta animantia quae sunt apud te ex omni carne tam in volatilibus quam in bestiis et in universis reptilibus quae reptant super terram educ tecum et ingredimini super terram crescite et multiplicamini super eam
GEN|8|18|egressus est ergo Noe et filii eius uxor illius et uxores filiorum eius cum eo
GEN|8|19|sed et omnia animantia iumenta et reptilia quae repunt super terram secundum genus suum arcam egressa sunt
GEN|8|20|aedificavit autem Noe altare Domino et tollens de cunctis pecoribus et volucribus mundis obtulit holocausta super altare
GEN|8|21|odoratusque est Dominus odorem suavitatis et ait ad eum nequaquam ultra maledicam terrae propter homines sensus enim et cogitatio humani cordis in malum prona sunt ab adulescentia sua non igitur ultra percutiam omnem animantem sicut feci
GEN|8|22|cunctis diebus terrae sementis et messis frigus et aestus aestas et hiemps nox et dies non requiescent
GEN|9|1|benedixitque Deus Noe et filiis eius et dixit ad eos crescite et multiplicamini et implete terram
GEN|9|2|et terror vester ac tremor sit super cuncta animalia terrae et super omnes volucres caeli cum universis quae moventur in terra omnes pisces maris manui vestrae traditi sunt
GEN|9|3|et omne quod movetur et vivit erit vobis in cibum quasi holera virentia tradidi vobis omnia
GEN|9|4|excepto quod carnem cum sanguine non comedetis
GEN|9|5|sanguinem enim animarum vestrarum requiram de manu cunctarum bestiarum et de manu hominis de manu viri et fratris eius requiram animam hominis
GEN|9|6|quicumque effuderit humanum sanguinem fundetur sanguis illius ad imaginem quippe Dei factus est homo
GEN|9|7|vos autem crescite et multiplicamini et ingredimini super terram et implete eam
GEN|9|8|haec quoque dixit Deus ad Noe et ad filios eius cum eo
GEN|9|9|ecce ego statuam pactum meum vobiscum et cum semine vestro post vos
GEN|9|10|et ad omnem animam viventem quae est vobiscum tam in volucribus quam in iumentis et pecudibus terrae cunctis quae egressa sunt de arca et universis bestiis terrae
GEN|9|11|statuam pactum meum vobiscum et nequaquam ultra interficietur omnis caro aquis diluvii neque erit deinceps diluvium dissipans terram
GEN|9|12|dixitque Deus hoc signum foederis quod do inter me et vos et ad omnem animam viventem quae est vobiscum in generationes sempiternas
GEN|9|13|arcum meum ponam in nubibus et erit signum foederis inter me et inter terram
GEN|9|14|cumque obduxero nubibus caelum apparebit arcus meus in nubibus
GEN|9|15|et recordabor foederis mei vobiscum et cum omni anima vivente quae carnem vegetat et non erunt ultra aquae diluvii ad delendam universam carnem
GEN|9|16|eritque arcus in nubibus et videbo illum et recordabor foederis sempiterni quod pactum est inter Deum et inter omnem animam viventem universae carnis quae est super terram
GEN|9|17|dixitque Deus Noe hoc erit signum foederis quod constitui inter me et inter omnem carnem super terram
GEN|9|18|erant igitur filii Noe qui egressi sunt de arca Sem Ham et Iafeth porro Ham ipse est pater Chanaan
GEN|9|19|tres isti sunt filii Noe et ab his disseminatum est omne hominum genus super universam terram
GEN|9|20|coepitque Noe vir agricola exercere terram et plantavit vineam
GEN|9|21|bibensque vinum inebriatus est et nudatus in tabernaculo suo
GEN|9|22|quod cum vidisset Ham pater Chanaan verenda scilicet patris sui esse nuda nuntiavit duobus fratribus suis foras
GEN|9|23|at vero Sem et Iafeth pallium inposuerunt umeris suis et incedentes retrorsum operuerunt verecunda patris sui faciesque eorum aversae erant et patris virilia non viderunt
GEN|9|24|evigilans autem Noe ex vino cum didicisset quae fecerat ei filius suus minor
GEN|9|25|ait maledictus Chanaan servus servorum erit fratribus suis
GEN|9|26|dixitque benedictus Dominus Deus Sem sit Chanaan servus eius
GEN|9|27|dilatet Deus Iafeth et habitet in tabernaculis Sem sitque Chanaan servus eius
GEN|9|28|vixit autem Noe post diluvium trecentis quinquaginta annis
GEN|9|29|et impleti sunt omnes dies eius nongentorum quinquaginta annorum et mortuus est
GEN|10|1|hae generationes filiorum Noe Sem Ham Iafeth natique sunt eis filii post diluvium
GEN|10|2|filii Iafeth Gomer Magog et Madai Iavan et Thubal et Mosoch et Thiras
GEN|10|3|porro filii Gomer Aschenez et Rifath et Thogorma
GEN|10|4|filii autem Iavan Elisa et Tharsis Cetthim et Dodanim
GEN|10|5|ab his divisae sunt insulae gentium in regionibus suis unusquisque secundum linguam et familias in nationibus suis
GEN|10|6|filii autem Ham Chus et Mesraim et Fut et Chanaan
GEN|10|7|filii Chus Saba et Hevila et Sabatha et Regma et Sabathaca filii Regma Saba et Dadan
GEN|10|8|porro Chus genuit Nemrod ipse coepit esse potens in terra
GEN|10|9|et erat robustus venator coram Domino ab hoc exivit proverbium quasi Nemrod robustus venator coram Domino
GEN|10|10|fuit autem principium regni eius Babylon et Arach et Archad et Chalanne in terra Sennaar
GEN|10|11|de terra illa egressus est Assur et aedificavit Nineven et plateas civitatis et Chale
GEN|10|12|Resen quoque inter Nineven et Chale haec est civitas magna
GEN|10|13|at vero Mesraim genuit Ludim et Anamim et Laabim Nepthuim
GEN|10|14|et Phetrusim et Cesluim de quibus egressi sunt Philisthim et Capthurim
GEN|10|15|Chanaan autem genuit Sidonem primogenitum suum Ettheum
GEN|10|16|et Iebuseum et Amorreum Gergeseum
GEN|10|17|Eveum et Araceum Sineum
GEN|10|18|et Aradium Samariten et Amatheum et post haec disseminati sunt populi Chananeorum
GEN|10|19|factique sunt termini Chanaan venientibus a Sidone Geraram usque Gazam donec ingrediaris Sodomam et Gomorram et Adama et Seboim usque Lesa
GEN|10|20|hii filii Ham in cognationibus et linguis et generationibus terrisque et gentibus suis
GEN|10|21|de Sem quoque nati sunt patre omnium filiorum Eber fratre Iafeth maiore
GEN|10|22|filii Sem Aelam et Assur et Arfaxad et Lud et Aram
GEN|10|23|filii Aram Us et Hul et Gether et Mes
GEN|10|24|at vero Arfaxad genuit Sala de quo ortus est Eber
GEN|10|25|natique sunt Eber filii duo nomen uni Faleg eo quod in diebus eius divisa sit terra et nomen fratris eius Iectan
GEN|10|26|qui Iectan genuit Helmodad et Saleph et Asarmoth Iare
GEN|10|27|et Aduram et Uzal Decla
GEN|10|28|et Ebal et Abimahel Saba
GEN|10|29|et Ophir et Evila et Iobab omnes isti filii Iectan
GEN|10|30|et facta est habitatio eorum de Messa pergentibus usque Sephar montem orientalem
GEN|10|31|isti filii Sem secundum cognationes et linguas et regiones in gentibus suis
GEN|10|32|hae familiae Noe iuxta populos et nationes suas ab his divisae sunt gentes in terra post diluvium
GEN|11|1|erat autem terra labii unius et sermonum eorundem
GEN|11|2|cumque proficiscerentur de oriente invenerunt campum in terra Sennaar et habitaverunt in eo
GEN|11|3|dixitque alter ad proximum suum venite faciamus lateres et coquamus eos igni habueruntque lateres pro saxis et bitumen pro cemento
GEN|11|4|et dixerunt venite faciamus nobis civitatem et turrem cuius culmen pertingat ad caelum et celebremus nomen nostrum antequam dividamur in universas terras
GEN|11|5|descendit autem Dominus ut videret civitatem et turrem quam aedificabant filii Adam
GEN|11|6|et dixit ecce unus est populus et unum labium omnibus coeperuntque hoc facere nec desistent a cogitationibus suis donec eas opere conpleant
GEN|11|7|venite igitur descendamus et confundamus ibi linguam eorum ut non audiat unusquisque vocem proximi sui
GEN|11|8|atque ita divisit eos Dominus ex illo loco in universas terras et cessaverunt aedificare civitatem
GEN|11|9|et idcirco vocatum est nomen eius Babel quia ibi confusum est labium universae terrae et inde dispersit eos Dominus super faciem cunctarum regionum
GEN|11|10|hae generationes Sem Sem centum erat annorum quando genuit Arfaxad biennio post diluvium
GEN|11|11|vixitque Sem postquam genuit Arfaxad quingentos annos et genuit filios et filias
GEN|11|12|porro Arfaxad vixit triginta quinque annos et genuit Sale
GEN|11|13|vixitque Arfaxad postquam genuit Sale trecentis tribus annis et genuit filios et filias
GEN|11|14|Sale quoque vixit triginta annis et genuit Eber
GEN|11|15|vixitque Sale postquam genuit Eber quadringentis tribus annis et genuit filios et filias
GEN|11|16|vixit autem Eber triginta quattuor annis et genuit Faleg
GEN|11|17|et vixit Eber postquam genuit Faleg quadringentis triginta annis et genuit filios et filias
GEN|11|18|vixit quoque Faleg triginta annis et genuit Reu
GEN|11|19|vixitque Faleg postquam genuit Reu ducentis novem annis et genuit filios et filias
GEN|11|20|vixit autem Reu triginta duobus annis et genuit Sarug
GEN|11|21|vixitque Reu postquam genuit Sarug ducentis septem annis et genuit filios et filias
GEN|11|22|vixit vero Sarug triginta annis et genuit Nahor
GEN|11|23|vixitque Sarug postquam genuit Nahor ducentos annos et genuit filios et filias
GEN|11|24|vixit autem Nahor viginti novem annis et genuit Thare
GEN|11|25|vixitque Nahor postquam genuit Thare centum decem et novem annos et genuit filios et filias
GEN|11|26|vixitque Thare septuaginta annis et genuit Abram et Nahor et Aran
GEN|11|27|hae sunt autem generationes Thare Thare genuit Abram et Nahor et Aran porro Aran genuit Loth
GEN|11|28|mortuusque est Aran ante Thare patrem suum in terra nativitatis suae in Ur Chaldeorum
GEN|11|29|duxerunt autem Abram et Nahor uxores nomen autem uxoris Abram Sarai et nomen uxoris Nahor Melcha filia Aran patris Melchae et patris Ieschae
GEN|11|30|erat autem Sarai sterilis nec habebat liberos
GEN|11|31|tulit itaque Thare Abram filium suum et Loth filium Aran filium filii sui et Sarai nurum suam uxorem Abram filii sui et eduxit eos de Ur Chaldeorum ut irent in terram Chanaan veneruntque usque Haran et habitaverunt ibi
GEN|11|32|et facti sunt dies Thare ducentorum quinque annorum et mortuus est in Haran
GEN|12|1|dixit autem Dominus ad Abram egredere de terra tua et de cognatione tua et de domo patris tui in terram quam monstrabo tibi
GEN|12|2|faciamque te in gentem magnam et benedicam tibi et magnificabo nomen tuum erisque benedictus
GEN|12|3|benedicam benedicentibus tibi et maledicam maledicentibus tibi atque in te benedicentur universae cognationes terrae
GEN|12|4|egressus est itaque Abram sicut praeceperat ei Dominus et ivit cum eo Loth septuaginta quinque annorum erat Abram cum egrederetur de Haran
GEN|12|5|tulitque Sarai uxorem suam et Loth filium fratris sui universamque substantiam quam possederant et animas quas fecerant in Haran et egressi sunt ut irent in terram Chanaan cumque venissent in eam
GEN|12|6|pertransivit Abram terram usque ad locum Sychem usque ad convallem Inlustrem Chananeus autem tunc erat in terra
GEN|12|7|apparuitque Dominus Abram et dixit ei semini tuo dabo terram hanc qui aedificavit ibi altare Domino qui apparuerat ei
GEN|12|8|et inde transgrediens ad montem qui erat contra orientem Bethel tetendit ibi tabernaculum suum ab occidente habens Bethel et ab oriente Ai aedificavit quoque ibi altare Domino et invocavit nomen eius
GEN|12|9|perrexitque Abram vadens et ultra progrediens ad meridiem
GEN|12|10|facta est autem fames in terra descenditque Abram in Aegyptum ut peregrinaretur ibi praevaluerat enim fames in terra
GEN|12|11|cumque prope esset ut ingrederetur Aegyptum dixit Sarai uxori suae novi quod pulchra sis mulier
GEN|12|12|et quod cum viderint te Aegyptii dicturi sunt uxor ipsius est et interficient me et te reservabunt
GEN|12|13|dic ergo obsecro te quod soror mea sis ut bene sit mihi propter te et vivat anima mea ob gratiam tui
GEN|12|14|cum itaque ingressus esset Abram Aegyptum viderunt Aegyptii mulierem quod esset pulchra nimis
GEN|12|15|et nuntiaverunt principes Pharaoni et laudaverunt eam apud illum et sublata est mulier in domum Pharaonis
GEN|12|16|Abram vero bene usi sunt propter illam fueruntque ei oves et boves et asini et servi et famulae et asinae et cameli
GEN|12|17|flagellavit autem Dominus Pharaonem plagis maximis et domum eius propter Sarai uxorem Abram
GEN|12|18|vocavitque Pharao Abram et dixit ei quidnam est quod fecisti mihi quare non indicasti quod uxor tua esset
GEN|12|19|quam ob causam dixisti esse sororem tuam ut tollerem eam mihi in uxorem nunc igitur ecce coniux tua accipe eam et vade
GEN|12|20|praecepitque Pharao super Abram viris et deduxerunt eum et uxorem illius et omnia quae habebat
GEN|13|1|ascendit ergo Abram de Aegypto ipse et uxor eius et omnia quae habebat et Loth cum eo ad australem plagam
GEN|13|2|erat autem dives valde in possessione argenti et auri
GEN|13|3|reversusque est per iter quo venerat a meridie in Bethel usque ad locum ubi prius fixerat tabernaculum inter Bethel et Ai
GEN|13|4|in loco altaris quod fecerat prius et invocavit ibi nomen Domini
GEN|13|5|sed et Loth qui erat cum Abram fuerunt greges ovium et armenta et tabernacula
GEN|13|6|nec poterat eos capere terra ut habitarent simul erat quippe substantia eorum multa et non quibant habitare communiter
GEN|13|7|unde et facta est rixa inter pastores gregum Abram et Loth eo autem tempore Chananeus et Ferezeus habitabant in illa terra
GEN|13|8|dixit ergo Abram ad Loth ne quaeso sit iurgium inter me et te et inter pastores meos et pastores tuos fratres enim sumus
GEN|13|9|ecce universa terra coram te est recede a me obsecro si ad sinistram ieris ego ad dexteram tenebo si tu dexteram elegeris ego ad sinistram pergam
GEN|13|10|elevatis itaque Loth oculis vidit omnem circa regionem Iordanis quae universa inrigabatur antequam subverteret Dominus Sodomam et Gomorram sicut paradisus Domini et sicut Aegyptus venientibus in Segor
GEN|13|11|elegitque sibi Loth regionem circa Iordanem et recessit ab oriente divisique sunt alterutrum a fratre suo
GEN|13|12|Abram habitavit in terra Chanaan Loth moratus est in oppidis quae erant circa Iordanem et habitavit in Sodomis
GEN|13|13|homines autem Sodomitae pessimi erant et peccatores coram Domino nimis
GEN|13|14|dixitque Dominus ad Abram postquam divisus est Loth ab eo leva oculos tuos et vide a loco in quo nunc es ad aquilonem et ad meridiem ad orientem et ad occidentem
GEN|13|15|omnem terram quam conspicis tibi dabo et semini tuo usque in sempiternum
GEN|13|16|faciamque semen tuum sicut pulverem terrae si quis potest hominum numerare pulverem semen quoque tuum numerare poterit
GEN|13|17|surge et perambula terram in longitudine et in latitudine sua quia tibi daturus sum eam
GEN|13|18|movens igitur Abram tabernaculum suum venit et habitavit iuxta convallem Mambre quod est in Hebron aedificavitque ibi altare Domino
GEN|14|1|factum est autem in illo tempore ut Amrafel rex Sennaar et Arioch rex Ponti et Chodorlahomor rex Aelamitarum et Thadal rex Gentium
GEN|14|2|inirent bellum contra Bara regem Sodomorum et contra Bersa regem Gomorrae et contra Sennaab regem Adamae et contra Semeber regem Seboim contraque regem Balae ipsa est Segor
GEN|14|3|omnes hii convenerunt in vallem Silvestrem quae nunc est mare Salis
GEN|14|4|duodecim enim annis servierant Chodorlahomor et tertiodecimo anno recesserunt ab eo
GEN|14|5|igitur anno quartodecimo venit Chodorlahomor et reges qui erant cum eo percusseruntque Rafaim in Astharothcarnaim et Zuzim cum eis et Emim in Savecariathaim
GEN|14|6|et Chorreos in montibus Seir usque ad campestria Pharan quae est in solitudine
GEN|14|7|reversique sunt et venerunt ad fontem Mesfat ipsa est Cades et percusserunt omnem regionem Amalechitarum et Amorreum qui habitabat in Asasonthamar
GEN|14|8|et egressi sunt rex Sodomorum et rex Gomorrae rexque Adamae et rex Seboim necnon et rex Balae quae est Segor et direxerunt contra eos aciem in valle Silvestri
GEN|14|9|scilicet adversum Chodorlahomor regem Aelamitarum et Thadal regem Gentium et Amrafel regem Sennaar et Arioch regem Ponti quattuor reges adversus quinque
GEN|14|10|vallis autem Silvestris habebat puteos multos bituminis itaque rex Sodomorum et Gomorrae terga verterunt cecideruntque ibi et qui remanserant fugerunt ad montem
GEN|14|11|tulerunt autem omnem substantiam Sodomorum et Gomorrae et universa quae ad cibum pertinent et abierunt
GEN|14|12|necnon et Loth et substantiam eius filium fratris Abram qui habitabat in Sodomis
GEN|14|13|et ecce unus qui evaserat nuntiavit Abram Hebraeo qui habitabat in convalle Mambre Amorrei fratris Eschol et fratris Aner hii enim pepigerant foedus cum Abram
GEN|14|14|quod cum audisset Abram captum videlicet Loth fratrem suum numeravit expeditos vernaculos suos trecentos decem et octo et persecutus est eos usque Dan
GEN|14|15|et divisis sociis inruit super eos nocte percussitque eos et persecutus est usque Hoba quae est ad levam Damasci
GEN|14|16|reduxitque omnem substantiam et Loth fratrem suum cum substantia illius mulieres quoque et populum
GEN|14|17|egressus est autem rex Sodomorum in occursum eius postquam reversus est a caede Chodorlahomor et regum qui cum eo erant in valle Save quae est vallis Regis
GEN|14|18|at vero Melchisedech rex Salem proferens panem et vinum erat enim sacerdos Dei altissimi
GEN|14|19|benedixit ei et ait benedictus Abram Deo excelso qui creavit caelum et terram
GEN|14|20|et benedictus Deus excelsus quo protegente hostes in manibus tuis sunt et dedit ei decimas ex omnibus
GEN|14|21|dixit autem rex Sodomorum ad Abram da mihi animas cetera tolle tibi
GEN|14|22|qui respondit ei levo manum meam ad Dominum Deum excelsum possessorem caeli et terrae
GEN|14|23|quod a filo subteminis usque ad corrigiam caligae non accipiam ex omnibus quae tua sunt ne dicas ego ditavi Abram
GEN|14|24|exceptis his quae comederunt iuvenes et partibus virorum qui venerunt mecum Aner Eschol et Mambre isti accipient partes suas
GEN|15|1|his itaque transactis factus est sermo Domini ad Abram per visionem dicens noli timere Abram ego protector tuus sum et merces tua magna nimis
GEN|15|2|dixitque Abram Domine Deus quid dabis mihi ego vadam absque liberis et filius procuratoris domus meae iste Damascus Eliezer
GEN|15|3|addiditque Abram mihi autem non dedisti semen et ecce vernaculus meus heres meus erit
GEN|15|4|statimque sermo Domini factus est ad eum dicens non erit hic heres tuus sed qui egredietur de utero tuo ipsum habebis heredem
GEN|15|5|eduxitque eum foras et ait illi suspice caelum et numera stellas si potes et dixit ei sic erit semen tuum
GEN|15|6|credidit Domino et reputatum est ei ad iustitiam
GEN|15|7|dixitque ad eum ego Dominus qui eduxi te de Ur Chaldeorum ut darem tibi terram istam et possideres eam
GEN|15|8|at ille ait Domine Deus unde scire possum quod possessurus sim eam
GEN|15|9|respondens Dominus sume inquit mihi vaccam triennem et capram trimam et arietem annorum trium turturem quoque et columbam
GEN|15|10|qui tollens universa haec divisit per medium et utrasque partes contra se altrinsecus posuit aves autem non divisit
GEN|15|11|descenderuntque volucres super cadavera et abigebat eas Abram
GEN|15|12|cumque sol occumberet sopor inruit super Abram et horror magnus et tenebrosus invasit eum
GEN|15|13|dictumque est ad eum scito praenoscens quod peregrinum futurum sit semen tuum in terra non sua et subicient eos servituti et adfligent quadringentis annis
GEN|15|14|verumtamen gentem cui servituri sunt ego iudicabo et post haec egredientur cum magna substantia
GEN|15|15|tu autem ibis ad patres tuos in pace sepultus in senectute bona
GEN|15|16|generatione autem quarta revertentur huc necdum enim conpletae sunt iniquitates Amorreorum usque ad praesens tempus
GEN|15|17|cum ergo occubuisset sol facta est caligo tenebrosa et apparuit clibanus fumans et lampas ignis transiens inter divisiones illas
GEN|15|18|in die illo pepigit Dominus cum Abram foedus dicens semini tuo dabo terram hanc a fluvio Aegypti usque ad fluvium magnum flumen Eufraten
GEN|15|19|Cineos et Cenezeos et Cedmoneos
GEN|15|20|et Hettheos et Ferezeos Rafaim quoque
GEN|15|21|et Amorreos et Chananeos et Gergeseos et Iebuseos
GEN|16|1|igitur Sarai uxor Abram non genuerat liberos sed habens ancillam aegyptiam nomine Agar
GEN|16|2|dixit marito suo ecce conclusit me Dominus ne parerem ingredere ad ancillam meam si forte saltem ex illa suscipiam filios cumque ille adquiesceret deprecanti
GEN|16|3|tulit Agar Aegyptiam ancillam suam post annos decem quam habitare coeperant in terra Chanaan et dedit eam viro suo uxorem
GEN|16|4|qui ingressus est ad eam at illa concepisse se videns despexit dominam suam
GEN|16|5|dixitque Sarai ad Abram inique agis contra me ego dedi ancillam meam in sinum tuum quae videns quod conceperit despectui me habet iudicet Dominus inter me et te
GEN|16|6|cui respondens Abram ecce ait ancilla tua in manu tua est utere ea ut libet adfligente igitur eam Sarai fugam iniit
GEN|16|7|cumque invenisset illam angelus Domini iuxta fontem aquae in solitudine qui est in via Sur
GEN|16|8|dixit ad eam Agar ancilla Sarai unde venis et quo vadis quae respondit a facie Sarai dominae meae ego fugio
GEN|16|9|dixitque ei angelus Domini revertere ad dominam tuam et humiliare sub manibus ipsius
GEN|16|10|et rursum multiplicans inquit multiplicabo semen tuum et non numerabitur prae multitudine
GEN|16|11|ac deinceps ecce ait concepisti et paries filium vocabisque nomen eius Ismahel eo quod audierit Dominus adflictionem tuam
GEN|16|12|hic erit ferus homo manus eius contra omnes et manus omnium contra eum et e regione universorum fratrum suorum figet tabernacula
GEN|16|13|vocavit autem nomen Domini qui loquebatur ad eam Tu Deus qui vidisti me dixit enim profecto hic vidi posteriora videntis me
GEN|16|14|propterea appellavit puteum illum puteum Viventis et videntis me ipse est inter Cades et Barad
GEN|16|15|peperitque Abrae filium qui vocavit nomen eius Ismahel
GEN|16|16|octoginta et sex annorum erat quando peperit ei Agar Ismahelem
GEN|17|1|postquam vero nonaginta et novem annorum esse coeperat apparuit ei Dominus dixitque ad eum ego Deus omnipotens ambula coram me et esto perfectus
GEN|17|2|ponamque foedus meum inter me et te et multiplicabo te vehementer nimis
GEN|17|3|cecidit Abram pronus in faciem
GEN|17|4|dixitque ei Deus ego sum et pactum meum tecum erisque pater multarum gentium
GEN|17|5|nec ultra vocabitur nomen tuum Abram sed appellaberis Abraham quia patrem multarum gentium constitui te
GEN|17|6|faciamque te crescere vehementissime et ponam in gentibus regesque ex te egredientur
GEN|17|7|et statuam pactum meum inter me et te et inter semen tuum post te in generationibus suis foedere sempiterno ut sim Deus tuus et seminis tui post te
GEN|17|8|daboque tibi et semini tuo terram peregrinationis tuae omnem terram Chanaan in possessionem aeternam eroque Deus eorum
GEN|17|9|dixit iterum Deus ad Abraham et tu ergo custodies pactum meum et semen tuum post te in generationibus suis
GEN|17|10|hoc est pactum quod observabitis inter me et vos et semen tuum post te circumcidetur ex vobis omne masculinum
GEN|17|11|et circumcidetis carnem praeputii vestri ut sit in signum foederis inter me et vos
GEN|17|12|infans octo dierum circumcidetur in vobis omne masculinum in generationibus vestris tam vernaculus quam empticius circumcidetur et quicumque non fuerit de stirpe vestra
GEN|17|13|eritque pactum meum in carne vestra in foedus aeternum
GEN|17|14|masculus cuius praeputii caro circumcisa non fuerit delebitur anima illa de populo suo quia pactum meum irritum fecit
GEN|17|15|dixit quoque Deus ad Abraham Sarai uxorem tuam non vocabis Sarai sed Sarram
GEN|17|16|et benedicam ei et ex illa dabo tibi filium cui benedicturus sum eritque in nationes et reges populorum orientur ex eo
GEN|17|17|cecidit Abraham in faciem et risit dicens in corde suo putasne centenario nascetur filius et Sarra nonagenaria pariet
GEN|17|18|dixitque ad Deum utinam Ismahel vivat coram te
GEN|17|19|et ait Deus ad Abraham Sarra uxor tua pariet tibi filium vocabisque nomen eius Isaac et constituam pactum meum illi in foedus sempiternum et semini eius post eum
GEN|17|20|super Ismahel quoque exaudivi te ecce benedicam ei et augebo et multiplicabo eum valde duodecim duces generabit et faciam illum in gentem magnam
GEN|17|21|pactum vero meum statuam ad Isaac quem pariet tibi Sarra tempore isto in anno altero
GEN|17|22|cumque finitus esset sermo loquentis cum eo ascendit Deus ab Abraham
GEN|17|23|tulit autem Abraham Ismahelem filium suum et omnes vernaculos domus suae universosque quos emerat cunctos mares ex omnibus viris domus suae et circumcidit carnem praeputii eorum statim in ipsa die sicut praeceperat ei Deus
GEN|17|24|nonaginta novem erat annorum quando circumcidit carnem praeputii sui
GEN|17|25|et Ismahel filius eius tredecim annos impleverat tempore circumcisionis suae
GEN|17|26|eadem die circumcisus est Abraham et Ismahel filius eius
GEN|17|27|et omnes viri domus illius tam vernaculi quam empticii et alienigenae pariter circumcisi sunt
GEN|18|1|apparuit autem ei Dominus in convalle Mambre sedenti in ostio tabernaculi sui in ipso fervore diei
GEN|18|2|cumque elevasset oculos apparuerunt ei tres viri stantes propter eum quos cum vidisset cucurrit in occursum eorum de ostio tabernaculi et adoravit in terra
GEN|18|3|et dixit Domine si inveni gratiam in oculis tuis ne transeas servum tuum
GEN|18|4|sed adferam pauxillum aquae et lavate pedes vestros et requiescite sub arbore
GEN|18|5|ponam buccellam panis et confortate cor vestrum postea transibitis idcirco enim declinastis ad servum vestrum qui dixerunt fac ut locutus es
GEN|18|6|festinavit Abraham in tabernaculum ad Sarram dixitque ei adcelera tria sata similae commisce et fac subcinericios panes
GEN|18|7|ipse vero ad armentum cucurrit et tulit inde vitulum tenerrimum et optimum deditque puero qui festinavit et coxit illum
GEN|18|8|tulit quoque butyrum et lac et vitulum quem coxerat et posuit coram eis ipse vero stabat iuxta eos sub arbore
GEN|18|9|cumque comedissent dixerunt ad eum ubi est Sarra uxor tua ille respondit ecce in tabernaculo est
GEN|18|10|cui dixit revertens veniam ad te tempore isto vita comite et habebit filium Sarra uxor tua quo audito Sarra risit post ostium tabernaculi
GEN|18|11|erant autem ambo senes provectaeque aetatis et desierant Sarrae fieri muliebria
GEN|18|12|quae risit occulte dicens postquam consenui et dominus meus vetulus est voluptati operam dabo
GEN|18|13|dixit autem Dominus ad Abraham quare risit Sarra dicens num vere paritura sum anus
GEN|18|14|numquid Deo est quicquam difficile iuxta condictum revertar ad te hoc eodem tempore vita comite et habebit Sarra filium
GEN|18|15|negavit Sarra dicens non risi timore perterrita Dominus autem non est inquit ita sed risisti
GEN|18|16|cum ergo surrexissent inde viri direxerunt oculos suos contra Sodomam et Abraham simul gradiebatur deducens eos
GEN|18|17|dixitque Dominus num celare potero Abraham quae gesturus sum
GEN|18|18|cum futurus sit in gentem magnam ac robustissimam et benedicendae sint in illo omnes nationes terrae
GEN|18|19|scio enim quod praecepturus sit filiis suis et domui suae post se ut custodiant viam Domini et faciant iustitiam et iudicium ut adducat Dominus propter Abraham omnia quae locutus est ad eum
GEN|18|20|dixit itaque Dominus clamor Sodomorum et Gomorrae multiplicatus est et peccatum earum adgravatum est nimis
GEN|18|21|descendam et videbo utrum clamorem qui venit ad me opere conpleverint an non est ita ut sciam
GEN|18|22|converteruntque se inde et abierunt Sodomam Abraham vero adhuc stabat coram Domino
GEN|18|23|et adpropinquans ait numquid perdes iustum cum impio
GEN|18|24|si fuerint quinquaginta iusti in civitate peribunt simul et non parces loco illi propter quinquaginta iustos si fuerint in eo
GEN|18|25|absit a te ut rem hanc facias et occidas iustum cum impio fiatque iustus sicut impius non est hoc tuum qui iudicas omnem terram nequaquam facies iudicium
GEN|18|26|dixitque Dominus ad eum si invenero Sodomis quinquaginta iustos in medio civitatis dimittam omni loco propter eos
GEN|18|27|respondens Abraham ait quia semel coepi loquar ad Dominum meum cum sim pulvis et cinis
GEN|18|28|quid si minus quinquaginta iustis quinque fuerint delebis propter quinque universam urbem et ait non delebo si invenero ibi quadraginta quinque
GEN|18|29|rursumque locutus est ad eum sin autem quadraginta inventi fuerint quid facies ait non percutiam propter quadraginta
GEN|18|30|ne quaeso inquit indigneris Domine si loquar quid si inventi fuerint ibi triginta respondit non faciam si invenero ibi triginta
GEN|18|31|quia semel ait coepi loquar ad Dominum meum quid si inventi fuerint ibi viginti dixit non interficiam propter viginti
GEN|18|32|obsecro inquit ne irascaris Domine si loquar adhuc semel quid si inventi fuerint ibi decem dixit non delebo propter decem
GEN|18|33|abiit Dominus postquam cessavit loqui ad Abraham et ille reversus est in locum suum
GEN|19|1|veneruntque duo angeli Sodomam vespere sedente Loth in foribus civitatis qui cum vidisset surrexit et ivit obviam eis adoravitque pronus in terra
GEN|19|2|et dixit obsecro domini declinate in domum pueri vestri et manete ibi lavate pedes vestros et mane proficiscimini in viam vestram qui dixerunt minime sed in platea manebimus
GEN|19|3|conpulit illos oppido ut deverterent ad eum ingressisque domum illius fecit convivium coxit azyma et comederunt
GEN|19|4|prius autem quam irent cubitum viri civitatis vallaverunt domum a puero usque ad senem omnis populus simul
GEN|19|5|vocaveruntque Loth et dixerunt ei ubi sunt viri qui introierunt ad te nocte educ illos huc ut cognoscamus eos
GEN|19|6|egressus ad eos Loth post tergum adcludens ostium ait
GEN|19|7|nolite quaeso fratres mei nolite malum hoc facere
GEN|19|8|habeo duas filias quae necdum cognoverunt virum educam eas ad vos et abutimini eis sicut placuerit vobis dummodo viris istis nihil faciatis mali quia ingressi sunt sub umbraculum tegminis mei
GEN|19|9|at illi dixerunt recede illuc et rursus ingressus es inquiunt ut advena numquid ut iudices te ergo ipsum magis quam hos adfligemus vimque faciebant Loth vehementissime iam prope erat ut refringerent fores
GEN|19|10|et ecce miserunt manum viri et introduxerunt ad se Loth cluseruntque ostium
GEN|19|11|et eos qui erant foris percusserunt caecitate a minimo usque ad maximum ita ut ostium invenire non possent
GEN|19|12|dixerunt autem ad Loth habes hic tuorum quempiam generum aut filios aut filias omnes qui tui sunt educ de urbe hac
GEN|19|13|delebimus enim locum istum eo quod increverit clamor eorum coram Domino qui misit nos ut perdamus illos
GEN|19|14|egressus itaque Loth locutus est ad generos suos qui accepturi erant filias eius et dixit surgite egredimini de loco isto quia delebit Dominus civitatem hanc et visus est eis quasi ludens loqui
GEN|19|15|cumque esset mane cogebant eum angeli dicentes surge et tolle uxorem tuam et duas filias quas habes ne et tu pariter pereas in scelere civitatis
GEN|19|16|dissimulante illo adprehenderunt manum eius et manum uxoris ac duarum filiarum eius eo quod parceret Dominus illi
GEN|19|17|et eduxerunt eum posueruntque extra civitatem ibi locutus est ad eum salva animam tuam noli respicere post tergum nec stes in omni circa regione sed in monte salvum te fac ne et tu simul pereas
GEN|19|18|dixitque Loth ad eos quaeso Domine mi
GEN|19|19|quia invenit servus tuus gratiam coram te et magnificasti misericordiam tuam quam fecisti mecum ut salvares animam meam nec possum in monte salvari ne forte adprehendat me malum et moriar
GEN|19|20|est civitas haec iuxta ad quam possum fugere parva et salvabor in ea numquid non modica est et vivet anima mea
GEN|19|21|dixitque ad eum ecce etiam in hoc suscepi preces tuas ut non subvertam urbem pro qua locutus es
GEN|19|22|festina et salvare ibi quia non potero facere quicquam donec ingrediaris illuc idcirco vocatum est nomen urbis illius Segor
GEN|19|23|sol egressus est super terram et Loth ingressus est in Segor
GEN|19|24|igitur Dominus pluit super Sodomam et Gomorram sulphur et ignem a Domino de caelo
GEN|19|25|et subvertit civitates has et omnem circa regionem universos habitatores urbium et cuncta terrae virentia
GEN|19|26|respiciensque uxor eius post se versa est in statuam salis
GEN|19|27|Abraham autem consurgens mane ubi steterat prius cum Domino
GEN|19|28|intuitus est Sodomam et Gomorram et universam terram regionis illius viditque ascendentem favillam de terra quasi fornacis fumum
GEN|19|29|cum enim subverteret Deus civitates regionis illius recordatus est Abrahae et liberavit Loth de subversione urbium in quibus habitaverat
GEN|19|30|ascenditque Loth de Segor et mansit in monte duae quoque filiae eius cum eo timuerat enim manere in Segor et mansit in spelunca ipse et duae filiae eius
GEN|19|31|dixitque maior ad minorem pater noster senex est et nullus virorum remansit in terra qui possit ingredi ad nos iuxta morem universae terrae
GEN|19|32|veni inebriemus eum vino dormiamusque cum eo ut servare possimus ex patre nostro semen
GEN|19|33|dederunt itaque patri suo bibere vinum nocte illa et ingressa est maior dormivitque cum patre at ille non sensit nec quando accubuit filia nec quando surrexit
GEN|19|34|altera quoque die dixit maior ad minorem ecce dormivi heri cum patre meo demus ei bibere vinum etiam hac nocte et dormies cum eo ut salvemus semen de patre nostro
GEN|19|35|dederunt et illa nocte patri vinum ingressaque minor filia dormivit cum eo et nec tunc quidem sensit quando concubuerit vel quando illa surrexerit
GEN|19|36|conceperunt ergo duae filiae Loth de patre suo
GEN|19|37|peperitque maior filium et vocavit nomen eius Moab ipse est pater Moabitarum usque in praesentem diem
GEN|19|38|minor quoque peperit filium et vocavit nomen eius Ammon id est filius populi mei ipse est pater Ammanitarum usque hodie
GEN|20|1|profectus inde Abraham in terram australem habitavit inter Cades et Sur et peregrinatus est in Geraris
GEN|20|2|dixitque de Sarra uxore sua soror mea est misit ergo Abimelech rex Gerarae et tulit eam
GEN|20|3|venit autem Deus ad Abimelech per somnium noctis et ait ei en morieris propter mulierem quam tulisti habet enim virum
GEN|20|4|Abimelech vero non tetigerat eam et ait Domine num gentem ignorantem et iustam interficies
GEN|20|5|nonne ipse dixit mihi soror mea est et ipsa ait frater meus est in simplicitate cordis mei et munditia manuum mearum feci hoc
GEN|20|6|dixitque ad eum Deus et ego scio quod simplici corde feceris et ideo custodivi te ne peccares in me et non dimisi ut tangeres eam
GEN|20|7|nunc igitur redde uxorem viro suo quia propheta est et orabit pro te et vives si autem nolueris reddere scito quod morte morieris tu et omnia quae tua sunt
GEN|20|8|statimque de nocte consurgens Abimelech vocavit omnes servos suos et locutus est universa verba haec in auribus eorum timueruntque omnes viri valde
GEN|20|9|vocavit autem Abimelech etiam Abraham et dixit ei quid fecisti nobis quid peccavimus in te quia induxisti super me et super regnum meum peccatum grande quae non debuisti facere fecisti nobis
GEN|20|10|rursusque expostulans ait quid vidisti ut hoc faceres
GEN|20|11|respondit Abraham cogitavi mecum dicens forsitan non est timor Dei in loco isto et interficient me propter uxorem meam
GEN|20|12|alias autem et vere soror mea est filia patris mei et non filia matris meae et duxi eam uxorem
GEN|20|13|postquam autem eduxit me Deus de domo patris mei dixi ad eam hanc misericordiam facies mecum in omni loco ad quem ingrediemur dices quod frater tuus sim
GEN|20|14|tulit igitur Abimelech oves et boves et servos et ancillas et dedit Abraham reddiditque illi Sarram uxorem suam
GEN|20|15|et ait terra coram vobis est ubicumque tibi placuerit habita
GEN|20|16|Sarrae autem dixit ecce mille argenteos dedi fratri tuo hoc erit tibi in velamen oculorum ad omnes qui tecum sunt et quocumque perrexeris mementoque te deprehensam
GEN|20|17|orante autem Abraham sanavit Deus Abimelech et uxorem ancillasque eius et pepererunt
GEN|20|18|concluserat enim Deus omnem vulvam domus Abimelech propter Sarram uxorem Abraham
GEN|21|1|visitavit autem Dominus Sarram sicut promiserat et implevit quae locutus est
GEN|21|2|concepitque et peperit filium in senectute sua tempore quo praedixerat ei Deus
GEN|21|3|vocavitque Abraham nomen filii sui quem genuit ei Sarra Isaac
GEN|21|4|et circumcidit eum octavo die sicut praeceperat ei Deus
GEN|21|5|cum centum esset annorum hac quippe aetate patris natus est Isaac
GEN|21|6|dixitque Sarra risum fecit mihi Deus quicumque audierit conridebit mihi
GEN|21|7|rursumque ait quis auditurum crederet Abraham quod Sarra lactaret filium quem peperit ei iam seni
GEN|21|8|crevit igitur puer et ablactatus est fecitque Abraham grande convivium in die ablactationis eius
GEN|21|9|cumque vidisset Sarra filium Agar Aegyptiae ludentem dixit ad Abraham
GEN|21|10|eice ancillam hanc et filium eius non enim erit heres filius ancillae cum filio meo Isaac
GEN|21|11|dure accepit hoc Abraham pro filio suo
GEN|21|12|cui dixit Deus non tibi videatur asperum super puero et super ancilla tua omnia quae dixerit tibi Sarra audi vocem eius quia in Isaac vocabitur tibi semen
GEN|21|13|sed et filium ancillae faciam in gentem magnam quia semen tuum est
GEN|21|14|surrexit itaque Abraham mane et tollens panem et utrem aquae inposuit scapulae eius tradiditque puerum et dimisit eam quae cum abisset errabat in solitudine Bersabee
GEN|21|15|cumque consumpta esset aqua in utre abiecit puerum subter unam arborum quae ibi erant
GEN|21|16|et abiit seditque e regione procul quantum potest arcus iacere dixit enim non videbo morientem puerum et sedens contra levavit vocem suam et flevit
GEN|21|17|exaudivit autem Deus vocem pueri vocavitque angelus Domini Agar de caelo dicens quid agis Agar noli timere exaudivit enim Deus vocem pueri de loco in quo est
GEN|21|18|surge tolle puerum et tene manum illius quia in gentem magnam faciam eum
GEN|21|19|aperuitque oculos eius Deus quae videns puteum aquae abiit et implevit utrem deditque puero bibere
GEN|21|20|et fuit cum eo qui crevit et moratus est in solitudine et factus est iuvenis sagittarius
GEN|21|21|habitavitque in deserto Pharan et accepit illi mater sua uxorem de terra Aegypti
GEN|21|22|eodem tempore dixit Abimelech et Fichol princeps exercitus eius ad Abraham Deus tecum est in universis quae agis
GEN|21|23|iura ergo per Dominum ne noceas mihi et posteris meis stirpique meae sed iuxta misericordiam quam feci tibi facies mihi et terrae in qua versatus es advena
GEN|21|24|dixitque Abraham ego iurabo
GEN|21|25|et increpavit Abimelech propter puteum aquae quem vi abstulerant servi illius
GEN|21|26|respondit Abimelech nescivi quis fecerit hanc rem sed et tu non indicasti mihi et ego non audivi praeter hodie
GEN|21|27|tulit itaque Abraham oves et boves et dedit Abimelech percusseruntque ambo foedus
GEN|21|28|et statuit Abraham septem agnas gregis seorsum
GEN|21|29|cui dixit Abimelech quid sibi volunt septem agnae istae quas stare fecisti seorsum
GEN|21|30|at ille septem inquit agnas accipies de manu mea ut sint in testimonium mihi quoniam ego fodi puteum istum
GEN|21|31|idcirco vocatus est locus ille Bersabee quia ibi uterque iuraverunt
GEN|21|32|et inierunt foedus pro puteo Iuramenti
GEN|21|33|surrexit autem Abimelech et Fichol princeps militiae eius reversique sunt in terram Palestinorum Abraham vero plantavit nemus in Bersabee et invocavit ibi nomen Domini Dei aeterni
GEN|21|34|et fuit colonus terrae Philisthinorum diebus multis
GEN|22|1|quae postquam gesta sunt temptavit Deus Abraham et dixit ad eum Abraham ille respondit adsum
GEN|22|2|ait ei tolle filium tuum unigenitum quem diligis Isaac et vade in terram Visionis atque offer eum ibi holocaustum super unum montium quem monstravero tibi
GEN|22|3|igitur Abraham de nocte consurgens stravit asinum suum ducens secum duos iuvenes et Isaac filium suum cumque concidisset ligna in holocaustum abiit ad locum quem praeceperat ei Deus
GEN|22|4|die autem tertio elevatis oculis vidit locum procul
GEN|22|5|dixitque ad pueros suos expectate hic cum asino ego et puer illuc usque properantes postquam adoraverimus revertemur ad vos
GEN|22|6|tulit quoque ligna holocausti et inposuit super Isaac filium suum ipse vero portabat in manibus ignem et gladium cumque duo pergerent simul
GEN|22|7|dixit Isaac patri suo pater mi at ille respondit quid vis fili ecce inquit ignis et ligna ubi est victima holocausti
GEN|22|8|dixit Abraham Deus providebit sibi victimam holocausti fili mi pergebant ergo pariter
GEN|22|9|veneruntque ad locum quem ostenderat ei Deus in quo aedificavit altare et desuper ligna conposuit cumque conligasset Isaac filium suum posuit eum in altari super struem lignorum
GEN|22|10|extenditque manum et arripuit gladium ut immolaret filium
GEN|22|11|et ecce angelus Domini de caelo clamavit dicens Abraham Abraham qui respondit adsum
GEN|22|12|dixitque ei non extendas manum tuam super puerum neque facias illi quicquam nunc cognovi quod timeas Dominum et non peperceris filio tuo unigenito propter me
GEN|22|13|levavit Abraham oculos viditque post tergum arietem inter vepres herentem cornibus quem adsumens obtulit holocaustum pro filio
GEN|22|14|appellavitque nomen loci illius Dominus videt unde usque hodie dicitur in monte Dominus videbit
GEN|22|15|vocavit autem angelus Domini Abraham secundo de caelo dicens
GEN|22|16|per memet ipsum iuravi dicit Dominus quia fecisti rem hanc et non pepercisti filio tuo unigenito
GEN|22|17|benedicam tibi et multiplicabo semen tuum sicut stellas caeli et velut harenam quae est in litore maris possidebit semen tuum portas inimicorum suorum
GEN|22|18|et benedicentur in semine tuo omnes gentes terrae quia oboedisti voci meae
GEN|22|19|reversus est Abraham ad pueros suos abieruntque Bersabee simul et habitavit ibi
GEN|22|20|his itaque gestis nuntiatum est Abraham quod Melcha quoque genuisset filios Nahor fratri suo
GEN|22|21|Hus primogenitum et Buz fratrem eius Camuhel patrem Syrorum
GEN|22|22|et Chased et Azau Pheldas quoque et Iedlaph
GEN|22|23|ac Bathuel de quo nata est Rebecca octo istos genuit Melcha Nahor fratri Abraham
GEN|22|24|concubina vero illius nomine Roma peperit Tabee et Gaom et Thaas et Maacha
GEN|23|1|vixit autem Sarra centum viginti septem annis
GEN|23|2|et mortua est in civitate Arbee quae est Hebron in terra Chanaan venitque Abraham ut plangeret et fleret eam
GEN|23|3|cumque surrexisset ab officio funeris locutus est ad filios Heth dicens
GEN|23|4|advena sum et peregrinus apud vos date mihi ius sepulchri vobiscum ut sepeliam mortuum meum
GEN|23|5|responderuntque filii Heth
GEN|23|6|audi nos domine princeps Dei es apud nos in electis sepulchris nostris sepeli mortuum tuum nullusque prohibere te poterit quin in monumento eius sepelias mortuum tuum
GEN|23|7|surrexit Abraham et adoravit populum terrae filios videlicet Heth
GEN|23|8|dixitque ad eos si placet animae vestrae ut sepeliam mortuum meum audite me et intercedite apud Ephron filium Soor
GEN|23|9|ut det mihi speluncam duplicem quam habet in extrema parte agri sui pecunia digna tradat mihi eam coram vobis in possessionem sepulchri
GEN|23|10|habitabat autem Ephron in medio filiorum Heth responditque ad Abraham cunctis audientibus qui ingrediebantur portam civitatis illius dicens
GEN|23|11|nequaquam ita fiat domine mi sed magis ausculta quod loquor agrum trado tibi et speluncam quae in eo est praesentibus filiis populi mei sepeli mortuum tuum
GEN|23|12|adoravit Abraham coram populo terrae
GEN|23|13|et locutus est ad Ephron circumstante plebe quaeso ut audias me dabo pecuniam pro agro suscipe eam et sic sepeliam mortuum meum in eo
GEN|23|14|respondit Ephron
GEN|23|15|domine mi audi terram quam postulas quadringentis argenti siclis valet istud est pretium inter me et te sed quantum est hoc sepeli mortuum tuum
GEN|23|16|quod cum audisset Abraham adpendit pecuniam quam Ephron postulaverat audientibus filiis Heth quadringentos siclos argenti et probati monetae publicae
GEN|23|17|confirmatusque est ager quondam Ephronis in quo erat spelunca duplex respiciens Mambre tam ipse quam spelunca et omnes arbores eius in cunctis terminis per circuitum
GEN|23|18|Abrahae in possessionem videntibus filiis Heth et cunctis qui intrabant portam civitatis illius
GEN|23|19|atque ita sepelivit Abraham Sarram uxorem suam in spelunca agri duplici qui respiciebat Mambre haec est Hebron in terra Chanaan
GEN|23|20|et confirmatus est ager et antrum quod erat in eo Abrahae in possessionem monumenti a filiis Heth
GEN|24|1|erat autem Abraham senex dierumque multorum et Dominus in cunctis benedixerat ei
GEN|24|2|dixitque ad servum seniorem domus suae qui praeerat omnibus quae habebat pone manum tuam subter femur meum
GEN|24|3|ut adiurem te per Dominum Deum caeli et terrae ut non accipias uxorem filio meo de filiabus Chananeorum inter quos habito
GEN|24|4|sed ad terram et ad cognationem meam proficiscaris et inde accipias uxorem filio meo Isaac
GEN|24|5|respondit servus si noluerit mulier venire mecum in terram hanc num reducere debeo filium tuum ad locum de quo egressus es
GEN|24|6|dixit Abraham cave nequando reducas illuc filium meum
GEN|24|7|Dominus Deus caeli qui tulit me de domo patris mei et de terra nativitatis meae qui locutus est mihi et iuravit dicens semini tuo dabo terram hanc ipse mittet angelum suum coram te et accipies inde uxorem filio meo
GEN|24|8|sin autem noluerit mulier sequi te non teneberis iuramento filium tantum meum ne reducas illuc
GEN|24|9|posuit ergo servus manum sub femore Abraham domini sui et iuravit illi super sermone hoc
GEN|24|10|tulitque decem camelos de grege domini sui et abiit ex omnibus bonis eius portans secum profectusque perrexit Mesopotamiam ad urbem Nahor
GEN|24|11|cumque camelos fecisset accumbere extra oppidum iuxta puteum aquae vespere eo tempore quo solent mulieres egredi ad hauriendam aquam dixit
GEN|24|12|Domine Deus domini mei Abraham occurre obsecro hodie mihi et fac misericordiam cum domino meo Abraham
GEN|24|13|ecce ego sto propter fontem aquae et filiae habitatorum huius civitatis egredientur ad hauriendam aquam
GEN|24|14|igitur puella cui ego dixero inclina hydriam tuam ut bibam et illa responderit bibe quin et camelis tuis dabo potum ipsa est quam praeparasti servo tuo Isaac et per hoc intellegam quod feceris misericordiam cum domino meo
GEN|24|15|necdum intra se verba conpleverat et ecce Rebecca egrediebatur filia Bathuel filii Melchae uxoris Nahor fratris Abraham habens hydriam in scapula
GEN|24|16|puella decora nimis virgoque pulcherrima et incognita viro descenderat autem ad fontem et impleverat hydriam ac revertebatur
GEN|24|17|occurritque ei servus et ait pauxillum mihi ad sorbendum praebe aquae de hydria tua
GEN|24|18|quae respondit bibe domine mi celeriterque deposuit hydriam super ulnam suam et dedit ei potum
GEN|24|19|cumque ille bibisset adiecit quin et camelis tuis hauriam aquam donec cuncti bibant
GEN|24|20|effundensque hydriam in canalibus recurrit ad puteum ut hauriret aquam et haustam omnibus camelis dedit
GEN|24|21|ille autem contemplabatur eam tacitus scire volens utrum prosperum fecisset iter suum Dominus an non
GEN|24|22|postquam ergo biberunt cameli protulit vir inaures aureas adpendentes siclos duos et armillas totidem pondo siclorum decem
GEN|24|23|dixitque ad eam cuius es filia indica mihi est in domo patris tui locus ad manendum
GEN|24|24|quae respondit filia Bathuelis sum filii Melchae quem peperit Nahor
GEN|24|25|et addidit dicens palearum quoque et faeni plurimum est apud nos et locus spatiosus ad manendum
GEN|24|26|inclinavit se homo et adoravit Dominum
GEN|24|27|dicens benedictus Dominus Deus domini mei Abraham qui non abstulit misericordiam et veritatem suam a domino meo et recto me itinere perduxit in domum fratris domini mei
GEN|24|28|cucurrit itaque puella et nuntiavit in domum matris suae omnia quae audierat
GEN|24|29|habebat autem Rebecca fratrem nomine Laban qui festinus egressus est ad hominem ubi erat fons
GEN|24|30|cumque vidisset inaures et armillas in manibus sororis suae et audisset cuncta verba referentis haec locutus est mihi homo venit ad virum qui stabat iuxta camelos et propter fontem aquae
GEN|24|31|dixitque ad eum ingredere benedicte Domini cur foris stas praeparavi domum et locum camelis
GEN|24|32|et introduxit eum hospitium ac destravit camelos deditque paleas et faenum et aquam ad lavandos pedes camelorum et virorum qui venerant cum eo
GEN|24|33|et adpositus est in conspectu eius panis qui ait non comedam donec loquar sermones meos respondit ei loquere
GEN|24|34|at ille servus inquit Abraham sum
GEN|24|35|et Dominus benedixit domino meo valde magnificatusque est et dedit ei oves et boves argentum et aurum servos et ancillas camelos et asinos
GEN|24|36|et peperit Sarra uxor domini mei filium domino meo in senectute sua deditque illi omnia quae habuerat
GEN|24|37|et adiuravit me dominus meus dicens non accipies uxorem filio meo de filiabus Chananeorum in quorum terra habito
GEN|24|38|sed ad domum patris mei perges et de cognatione mea accipies uxorem filio meo
GEN|24|39|ego vero respondi domino meo quid si noluerit venire mecum mulier
GEN|24|40|Dominus ait in cuius conspectu ambulo mittet angelum suum tecum et diriget viam tuam accipiesque uxorem filio meo de cognatione mea et de domo patris mei
GEN|24|41|innocens eris a maledictione mea cum veneris ad propinquos meos et non dederint tibi
GEN|24|42|veni ergo hodie ad fontem et dixi Domine Deus domini mei Abraham si direxisti viam meam in qua nunc ambulo
GEN|24|43|ecce sto iuxta fontem aquae et virgo quae egredietur ad hauriendam aquam audierit a me da mihi pauxillum aquae ad bibendum ex hydria tua
GEN|24|44|et dixerit mihi et tu bibe et camelis tuis hauriam ipsa est mulier quam praeparavit Dominus filio domini mei
GEN|24|45|dum haec mecum tacitus volverem apparuit Rebecca veniens cum hydria quam portabat in scapula descenditque ad fontem et hausit aquam et aio ad eam da mihi paululum bibere
GEN|24|46|quae festina deposuit hydriam de umero et dixit mihi et tu bibe et camelis tuis potum tribuam bibi et adaquavit camelos
GEN|24|47|interrogavique eam et dixi cuius es filia quae respondit filia Bathuelis sum filii Nahor quem peperit illi Melcha suspendi itaque inaures ad ornandam faciem eius et armillas posui in manibus
GEN|24|48|pronusque adoravi Dominum benedicens Domino Deo domini mei Abraham qui perduxisset me recto itinere ut sumerem filiam fratris domini mei filio eius
GEN|24|49|quam ob rem si facitis misericordiam et veritatem cum domino meo indicate mihi sin autem aliud placet et hoc dicite ut vadam ad dextram sive ad sinistram
GEN|24|50|responderunt Laban et Bathuel a Domino egressus est sermo non possumus extra placitum eius quicquam aliud tecum loqui
GEN|24|51|en Rebecca coram te est tolle eam et proficiscere et sit uxor filii domini tui sicut locutus est Dominus
GEN|24|52|quod cum audisset puer Abraham adoravit in terra Dominum
GEN|24|53|prolatisque vasis argenteis et aureis ac vestibus dedit ea Rebeccae pro munere fratribus quoque eius et matri dona obtulit
GEN|24|54|initoque convivio vescentes pariter et bibentes manserunt ibi surgens autem mane locutus est puer dimittite me ut vadam ad dominum meum
GEN|24|55|responderunt fratres eius et mater maneat puella saltem decem dies apud nos et postea proficiscetur
GEN|24|56|nolite ait me retinere quia Dominus direxit viam meam dimittite me ut pergam ad dominum meum
GEN|24|57|dixerunt vocemus puellam et quaeramus ipsius voluntatem
GEN|24|58|cumque vocata venisset sciscitati sunt vis ire cum homine isto quae ait vadam
GEN|24|59|dimiserunt ergo eam et nutricem illius servumque Abraham et comites eius
GEN|24|60|inprecantes prospera sorori suae atque dicentes soror nostra es crescas in mille milia et possideat semen tuum portas inimicorum suorum
GEN|24|61|igitur Rebecca et puellae illius ascensis camelis secutae sunt virum qui festinus revertebatur ad dominum suum
GEN|24|62|eo tempore Isaac deambulabat per viam quae ducit ad puteum cuius nomen est Viventis et videntis habitabat enim in terra australi
GEN|24|63|et egressus fuerat ad meditandum in agro inclinata iam die cumque levasset oculos vidit camelos venientes procul
GEN|24|64|Rebecca quoque conspecto Isaac descendit de camelo
GEN|24|65|et ait ad puerum quis est ille homo qui venit per agrum in occursum nobis dixit ei ipse est dominus meus at illa tollens cito pallium operuit se
GEN|24|66|servus autem cuncta quae gesserat narravit Isaac
GEN|24|67|qui introduxit eam in tabernaculum Sarrae matris suae et accepit uxorem et in tantum dilexit ut dolorem qui ex morte matris acciderat temperaret
GEN|25|1|Abraham vero aliam duxit uxorem nomine Cetthuram
GEN|25|2|quae peperit ei Zamram et Iexan et Madan et Madian et Iesboch et Sue
GEN|25|3|Iexan quoque genuit Saba et Dadan filii Dadan fuerunt Assurim et Lathusim et Loommim
GEN|25|4|at vero ex Madian ortus est Epha et Opher et Enoch et Abida et Eldaa omnes hii filii Cetthurae
GEN|25|5|deditque Abraham cuncta quae possederat Isaac
GEN|25|6|filiis autem concubinarum largitus est munera et separavit eos ab Isaac filio suo dum adhuc ipse viveret ad plagam orientalem
GEN|25|7|fuerunt autem dies vitae eius centum septuaginta quinque anni
GEN|25|8|et deficiens mortuus est in senectute bona provectaeque aetatis et plenus dierum congregatusque est ad populum suum
GEN|25|9|et sepelierunt eum Isaac et Ismahel filii sui in spelunca duplici quae sita est in agro Ephron filii Soor Hetthei e regione Mambre
GEN|25|10|quem emerat a filiis Heth ibi sepultus est ipse et Sarra uxor eius
GEN|25|11|et post obitum illius benedixit Deus Isaac filio eius qui habitabat iuxta puteum nomine Viventis et videntis
GEN|25|12|hae sunt generationes Ismahel filii Abraham quem peperit ei Agar Aegyptia famula Sarrae
GEN|25|13|et haec nomina filiorum eius in vocabulis et generationibus suis primogenitus Ismahelis Nabaioth dein Cedar et Abdeel et Mabsam
GEN|25|14|Masma quoque et Duma et Massa
GEN|25|15|Adad et Thema Itur et Naphis et Cedma
GEN|25|16|isti sunt filii Ismahel et haec nomina per castella et oppida eorum duodecim principes tribuum suarum
GEN|25|17|anni vitae Ismahel centum triginta septem deficiens mortuus est et adpositus ad populum suum
GEN|25|18|habitavit autem ab Evila usque Sur quae respicit Aegyptum introeuntibus Assyrios coram cunctis fratribus suis obiit
GEN|25|19|hae quoque sunt generationes Isaac filii Abraham Abraham genuit Isaac
GEN|25|20|qui cum quadraginta esset annorum duxit uxorem Rebeccam filiam Bathuel Syri de Mesopotamiam sororem Laban
GEN|25|21|deprecatusque est Dominum pro uxore sua eo quod esset sterilis qui exaudivit eum et dedit conceptum Rebeccae
GEN|25|22|sed conlidebantur in utero eius parvuli quae ait si sic mihi futurum erat quid necesse fuit concipere perrexitque ut consuleret Dominum
GEN|25|23|qui respondens ait duae gentes in utero tuo sunt et duo populi ex ventre tuo dividentur populusque populum superabit et maior minori serviet
GEN|25|24|iam tempus pariendi venerat et ecce gemini in utero repperti sunt
GEN|25|25|qui primus egressus est rufus erat et totus in morem pellis hispidus vocatumque est nomen eius Esau protinus alter egrediens plantam fratris tenebat manu et idcirco appellavit eum Iacob
GEN|25|26|sexagenarius erat Isaac quando nati sunt parvuli
GEN|25|27|quibus adultis factus est Esau vir gnarus venandi et homo agricola Iacob autem vir simplex habitabat in tabernaculis
GEN|25|28|Isaac amabat Esau eo quod de venationibus illius vesceretur et Rebecca diligebat Iacob
GEN|25|29|coxit autem Iacob pulmentum ad quem cum venisset Esau de agro lassus
GEN|25|30|ait da mihi de coctione hac rufa quia oppido lassus sum quam ob causam vocatum est nomen eius Edom
GEN|25|31|cui dixit Iacob vende mihi primogenita tua
GEN|25|32|ille respondit en morior quid mihi proderunt primogenita
GEN|25|33|ait Iacob iura ergo mihi iuravit Esau et vendidit primogenita
GEN|25|34|et sic accepto pane et lentis edulio comedit et bibit et abiit parvipendens quod primogenita vendidisset
GEN|26|1|orta autem fame super terram post eam sterilitatem quae acciderat in diebus Abraham abiit Isaac ad Abimelech regem Palestinorum in Gerara
GEN|26|2|apparuitque ei Dominus et ait ne descendas in Aegyptum sed quiesce in terra quam dixero tibi
GEN|26|3|et peregrinare in ea eroque tecum et benedicam tibi tibi enim et semini tuo dabo universas regiones has conplens iuramentum quod spopondi Abraham patri tuo
GEN|26|4|et multiplicabo semen tuum sicut stellas caeli daboque posteris tuis universas regiones has et benedicentur in semine tuo omnes gentes terrae
GEN|26|5|eo quod oboedierit Abraham voci meae et custodierit praecepta et mandata mea et caerimonias legesque servaverit
GEN|26|6|mansit itaque Isaac in Geraris
GEN|26|7|qui cum interrogaretur a viris loci illius super uxore sua respondit soror mea est timuerat enim confiteri quod sibi esset sociata coniugio reputans ne forte interficerent eum propter illius pulchritudinem
GEN|26|8|cumque pertransissent dies plurimi et ibi demoraretur prospiciens Abimelech Palestinorum rex per fenestram vidit eum iocantem cum Rebecca uxore sua
GEN|26|9|et accersito ait perspicuum est quod uxor tua sit cur mentitus es sororem tuam esse respondit timui ne morerer propter eam
GEN|26|10|dixitque Abimelech quare inposuisti nobis potuit coire quispiam de populo cum uxore tua et induxeras super nos grande peccatum praecepitque omni populo dicens
GEN|26|11|qui tetigerit hominis huius uxorem morte morietur
GEN|26|12|seruit autem Isaac in terra illa et invenit in ipso anno centuplum benedixitque ei Dominus
GEN|26|13|et locupletatus est homo et ibat proficiens atque succrescens donec magnus vehementer effectus est
GEN|26|14|habuit quoque possessionem ovium et armentorum et familiae plurimum ob haec invidentes ei Palestini
GEN|26|15|omnes puteos quos foderant servi patris illius Abraham illo tempore obstruxerunt implentes humo
GEN|26|16|in tantum ut ipse Abimelech diceret ad Isaac recede a nobis quoniam potentior nostri factus es valde
GEN|26|17|et ille discedens veniret ad torrentem Gerarae habitaretque ibi
GEN|26|18|rursum fodit alios puteos quos foderant servi patris sui Abraham et quos illo mortuo olim obstruxerant Philisthim appellavitque eos hisdem nominibus quibus ante pater vocaverat
GEN|26|19|foderunt in torrente et reppererunt aquam vivam
GEN|26|20|sed et ibi iurgium fuit pastorum Gerarae adversum pastores Isaac dicentium nostra est aqua quam ob rem nomen putei ex eo quod acciderat vocavit Calumniam
GEN|26|21|foderunt et alium et pro illo quoque rixati sunt appellavitque eum Inimicitias
GEN|26|22|profectus inde fodit alium puteum pro quo non contenderunt itaque vocavit nomen illius Latitudo dicens nunc dilatavit nos Dominus et fecit crescere super terram
GEN|26|23|ascendit autem ex illo loco in Bersabee
GEN|26|24|ubi apparuit ei Dominus in ipsa nocte dicens ego sum Deus Abraham patris tui noli metuere quia tecum sum benedicam tibi et multiplicabo semen tuum propter servum meum Abraham
GEN|26|25|itaque aedificavit ibi altare et invocato nomine Domini extendit tabernaculum praecepitque servis suis ut foderent puteum
GEN|26|26|ad quem locum cum venissent de Geraris Abimelech et Ochozath amicus illius et Fichol dux militum
GEN|26|27|locutus est eis Isaac quid venistis ad me hominem quem odistis et expulistis a vobis
GEN|26|28|qui responderunt vidimus tecum esse Dominum et idcirco nunc diximus sit iuramentum inter nos et ineamus foedus
GEN|26|29|ut non facias nobis quicquam mali sicut et nos nihil tuorum adtigimus nec fecimus quod te laederet sed cum pace dimisimus auctum benedictione Domini
GEN|26|30|fecit ergo eis convivium et post cibum et potum
GEN|26|31|surgentes mane iuraverunt sibi mutuo dimisitque eos Isaac pacifice in locum suum
GEN|26|32|ecce autem venerunt in ipso die servi Isaac adnuntiantes ei de puteo quem foderant atque dicentes invenimus aquam
GEN|26|33|unde appellavit eum Abundantiam et nomen urbi inpositum est Bersabee usque in praesentem diem
GEN|26|34|Esau vero quadragenarius duxit uxores Iudith filiam Beeri Hetthei et Basemath filiam Helon eiusdem loci
GEN|26|35|quae ambae offenderant animum Isaac et Rebeccae
GEN|27|1|senuit autem Isaac et caligaverunt oculi eius et videre non poterat vocavitque Esau filium suum maiorem et dixit ei fili mi qui respondit adsum
GEN|27|2|cui pater vides inquit quod senuerim et ignorem diem mortis meae
GEN|27|3|sume arma tua faretram et arcum et egredere foras cumque venatu aliquid adprehenderis
GEN|27|4|fac mihi inde pulmentum sicut velle me nosti et adfer ut comedam et benedicat tibi anima mea antequam moriar
GEN|27|5|quod cum audisset Rebecca et ille abisset in agrum ut iussionem patris expleret
GEN|27|6|dixit filio suo Iacob audivi patrem tuum loquentem cum Esau fratre tuo et dicentem ei
GEN|27|7|adfer mihi venationem tuam et fac cibos ut comedam et benedicam tibi coram Domino antequam moriar
GEN|27|8|nunc ergo fili mi adquiesce consiliis meis
GEN|27|9|et pergens ad gregem adfer mihi duos hedos optimos ut faciam ex eis escas patri tuo quibus libenter vescitur
GEN|27|10|quas cum intuleris et comederit benedicat tibi priusquam moriatur
GEN|27|11|cui ille respondit nosti quod Esau frater meus homo pilosus sit et ego lenis
GEN|27|12|si adtractaverit me pater meus et senserit timeo ne putet sibi voluisse inludere et inducat super me maledictionem pro benedictione
GEN|27|13|ad quem mater in me sit ait ista maledictio fili mi tantum audi vocem meam et perge adferque quae dixi
GEN|27|14|abiit et adtulit deditque matri paravit illa cibos sicut noverat velle patrem illius
GEN|27|15|et vestibus Esau valde bonis quas apud se habebat domi induit eum
GEN|27|16|pelliculasque hedorum circumdedit manibus et colli nuda protexit
GEN|27|17|dedit pulmentum et panes quos coxerat tradidit
GEN|27|18|quibus inlatis dixit pater mi et ille respondit audio quis tu es fili mi
GEN|27|19|dixitque Iacob ego sum Esau primogenitus tuus feci sicut praecepisti mihi surge sede et comede de venatione mea ut benedicat mihi anima tua
GEN|27|20|rursum Isaac ad filium suum quomodo inquit tam cito invenire potuisti fili mi qui respondit voluntatis Dei fuit ut cito mihi occurreret quod volebam
GEN|27|21|dixitque Isaac accede huc ut tangam te fili mi et probem utrum tu sis filius meus Esau an non
GEN|27|22|accessit ille ad patrem et palpato eo dixit Isaac vox quidem vox Iacob est sed manus manus sunt Esau
GEN|27|23|et non cognovit eum quia pilosae manus similitudinem maioris expresserant benedicens ergo illi
GEN|27|24|ait tu es filius meus Esau respondit ego sum
GEN|27|25|at ille offer inquit mihi cibos de venatione tua fili mi ut benedicat tibi anima mea quos cum oblatos comedisset obtulit ei etiam vinum quo hausto
GEN|27|26|dixit ad eum accede ad me et da mihi osculum fili mi
GEN|27|27|accessit et osculatus est eum statimque ut sensit vestimentorum illius flagrantiam benedicens ait ecce odor filii mei sicut odor agri cui benedixit Dominus
GEN|27|28|det tibi Deus de rore caeli et de pinguedine terrae abundantiam frumenti et vini
GEN|27|29|et serviant tibi populi et adorent te tribus esto dominus fratrum tuorum et incurventur ante te filii matris tuae qui maledixerit tibi sit maledictus et qui benedixerit benedictionibus repleatur
GEN|27|30|vix Isaac sermonem impleverat et egresso Iacob foras venit Esau
GEN|27|31|coctosque de venatione cibos intulit patri dicens surge pater mi et comede de venatione filii tui ut benedicat mihi anima tua
GEN|27|32|dixitque illi Isaac quis enim es tu qui respondit ego sum primogenitus filius tuus Esau
GEN|27|33|expavit Isaac stupore vehementi et ultra quam credi potest admirans ait quis igitur ille est qui dudum captam venationem adtulit mihi et comedi ex omnibus priusquam tu venires benedixique ei et erit benedictus
GEN|27|34|auditis Esau sermonibus patris inrugiit clamore magno et consternatus ait benedic etiam mihi pater mi
GEN|27|35|qui ait venit germanus tuus fraudulenter et accepit benedictionem tuam
GEN|27|36|at ille subiunxit iuste vocatum est nomen eius Iacob subplantavit enim me en altera vice primogenita mea ante tulit et nunc secundo subripuit benedictionem meam rursumque ad patrem numquid non reservasti ait et mihi benedictionem
GEN|27|37|respondit Isaac dominum tuum illum constitui et omnes fratres eius servituti illius subiugavi frumento et vino stabilivi eum tibi post haec fili mi ultra quid faciam
GEN|27|38|cui Esau num unam inquit tantum benedictionem habes pater mihi quoque obsecro ut benedicas cumque heiulatu magno fleret
GEN|27|39|motus Isaac dixit ad eum in pinguedine terrae et in rore caeli desuper
GEN|27|40|erit benedictio tua vives gladio et fratri tuo servies tempusque veniet cum excutias et solvas iugum eius de cervicibus tuis
GEN|27|41|oderat ergo semper Esau Iacob pro benedictione qua benedixerat ei pater dixitque in corde suo veniant dies luctus patris mei ut occidam Iacob fratrem meum
GEN|27|42|nuntiata sunt haec Rebeccae quae mittens et vocans Iacob filium suum dixit ad eum ecce Esau frater tuus minatur ut occidat te
GEN|27|43|nunc ergo fili audi vocem meam et consurgens fuge ad Laban fratrem meum in Haran
GEN|27|44|habitabisque cum eo dies paucos donec requiescat furor fratris tui
GEN|27|45|et cesset indignatio eius obliviscaturque eorum quae fecisti in eum postea mittam et adducam te inde huc cur utroque orbabor filio in una die
GEN|27|46|dixit quoque Rebecca ad Isaac taedet me vitae meae propter filias Heth si acceperit Iacob uxorem de stirpe huius terrae nolo vivere
GEN|28|1|vocavit itaque Isaac Iacob et benedixit praecepitque ei dicens noli accipere coniugem de genere Chanaan
GEN|28|2|sed vade et proficiscere in Mesopotamiam Syriae ad domum Bathuel patrem matris tuae et accipe tibi inde uxorem de filiabus Laban avunculi tui
GEN|28|3|Deus autem omnipotens benedicat tibi et crescere te faciat atque multiplicet ut sis in turbas populorum
GEN|28|4|et det tibi benedictiones Abraham et semini tuo post te ut possideas terram peregrinationis tuae quam pollicitus est avo tuo
GEN|28|5|cumque dimisisset eum Isaac profectus venit in Mesopotamiam Syriae ad Laban filium Bathuel Syri fratrem Rebeccae matris suae
GEN|28|6|videns autem Esau quod benedixisset pater suus Iacob et misisset eum in Mesopotamiam Syriae ut inde uxorem duceret et quod post benedictionem praecepisset ei dicens non accipies coniugem de filiabus Chanaan
GEN|28|7|quodque oboediens Iacob parentibus isset in Syriam
GEN|28|8|probans quoque quod non libenter aspiceret filias Chanaan pater suus
GEN|28|9|ivit ad Ismahelem et duxit uxorem absque his quas prius habebat Maeleth filiam Ismahel filii Abraham sororem Nabaioth
GEN|28|10|igitur egressus Iacob de Bersabee pergebat Haran
GEN|28|11|cumque venisset ad quendam locum et vellet in eo requiescere post solis occubitum tulit de lapidibus qui iacebant et subponens capiti suo dormivit in eodem loco
GEN|28|12|viditque in somnis scalam stantem super terram et cacumen illius tangens caelum angelos quoque Dei ascendentes et descendentes per eam
GEN|28|13|et Dominum innixum scalae dicentem sibi ego sum Dominus Deus Abraham patris tui et Deus Isaac terram in qua dormis tibi dabo et semini tuo
GEN|28|14|eritque germen tuum quasi pulvis terrae dilataberis ad occidentem et orientem septentrionem et meridiem et benedicentur in te et in semine tuo cunctae tribus terrae
GEN|28|15|et ero custos tuus quocumque perrexeris et reducam te in terram hanc nec dimittam nisi conplevero universa quae dixi
GEN|28|16|cumque evigilasset Iacob de somno ait vere Dominus est in loco isto et ego nesciebam
GEN|28|17|pavensque quam terribilis inquit est locus iste non est hic aliud nisi domus Dei et porta caeli
GEN|28|18|surgens ergo mane tulit lapidem quem subposuerat capiti suo et erexit in titulum fundens oleum desuper
GEN|28|19|appellavitque nomen urbis Bethel quae prius Luza vocabatur
GEN|28|20|vovit etiam votum dicens si fuerit Deus mecum et custodierit me in via per quam ambulo et dederit mihi panem ad vescendum et vestem ad induendum
GEN|28|21|reversusque fuero prospere ad domum patris mei erit mihi Dominus in Deum
GEN|28|22|et lapis iste quem erexi in titulum vocabitur Domus Dei cunctorumque quae dederis mihi decimas offeram tibi
GEN|29|1|profectus ergo Iacob venit ad terram orientalem
GEN|29|2|et vidit puteum in agro tresque greges ovium accubantes iuxta eum nam ex illo adaquabantur pecora et os eius grandi lapide claudebatur
GEN|29|3|morisque erat ut cunctis ovibus congregatis devolverent lapidem et refectis gregibus rursum super os putei ponerent
GEN|29|4|dixitque ad pastores fratres unde estis qui responderunt de Haran
GEN|29|5|quos interrogans numquid ait nostis Laban filium Nahor dixerunt novimus
GEN|29|6|sanusne est inquit valet inquiunt et ecce Rahel filia eius venit cum grege suo
GEN|29|7|dixitque Iacob adhuc multum diei superest nec est tempus ut reducantur ad caulas greges date ante potum ovibus et sic ad pastum eas reducite
GEN|29|8|qui responderunt non possumus donec omnia pecora congregentur et amoveamus lapidem de ore putei ut adaquemus greges
GEN|29|9|adhuc loquebantur et ecce Rahel veniebat cum ovibus patris sui nam gregem ipsa pascebat
GEN|29|10|quam cum vidisset Iacob et sciret consobrinam suam ovesque Laban avunculi sui amovit lapidem quo puteus claudebatur
GEN|29|11|et adaquato grege osculatus est eam elevataque voce flevit
GEN|29|12|et indicavit ei quod frater esset patris eius et filius Rebeccae at illa festinans nuntiavit patri suo
GEN|29|13|qui cum audisset venisse Iacob filium sororis suae cucurrit obviam conplexusque eum et in oscula ruens duxit in domum suam auditis autem causis itineris
GEN|29|14|respondit os meum es et caro mea et postquam expleti sunt dies mensis unius
GEN|29|15|dixit ei num quia frater meus es gratis servies mihi dic quid mercedis accipias
GEN|29|16|habebat vero filias duas nomen maioris Lia minor appellabatur Rahel
GEN|29|17|sed Lia lippis erat oculis Rahel decora facie et venusto aspectu
GEN|29|18|quam diligens Iacob ait serviam tibi pro Rahel filia tua minore septem annis
GEN|29|19|respondit Laban melius est ut tibi eam dem quam viro alteri mane apud me
GEN|29|20|servivit igitur Iacob pro Rahel septem annis et videbantur illi pauci dies prae amoris magnitudine
GEN|29|21|dixitque ad Laban da mihi uxorem meam quia iam tempus expletum est ut ingrediar ad eam
GEN|29|22|qui vocatis multis amicorum turbis ad convivium fecit nuptias
GEN|29|23|et vespere filiam suam Liam introduxit ad eum
GEN|29|24|dans ancillam filiae Zelpham nomine ad quam cum ex more Iacob fuisset ingressus facto mane vidit Liam
GEN|29|25|et dixit ad socerum quid est quod facere voluisti nonne pro Rahel servivi tibi quare inposuisti mihi
GEN|29|26|respondit Laban non est in loco nostro consuetudinis ut minores ante tradamus ad nuptias
GEN|29|27|imple ebdomadem dierum huius copulae et hanc quoque dabo tibi pro opere quo serviturus es mihi septem annis aliis
GEN|29|28|adquievit placito et ebdomade transacta Rahel duxit uxorem
GEN|29|29|cui pater servam Balam dederat
GEN|29|30|tandemque potitus optatis nuptiis amorem sequentis priori praetulit serviens apud eum septem annis aliis
GEN|29|31|videns autem Dominus quod despiceret Liam aperuit vulvam eius sorore sterili permanente
GEN|29|32|quae conceptum genuit filium vocavitque nomen eius Ruben dicens vidit Dominus humilitatem meam nunc amabit me vir meus
GEN|29|33|rursumque concepit et peperit filium et ait quoniam audivit Dominus haberi me contemptui dedit etiam istum mihi vocavitque nomen illius Symeon
GEN|29|34|concepit tertio et genuit alium dixitque nunc quoque copulabitur mihi maritus meus eo quod pepererim illi tres filios et idcirco appellavit nomen eius Levi
GEN|29|35|quarto concepit et peperit filium et ait modo confitebor Domino et ob hoc vocavit eum Iudam cessavitque parere
GEN|30|1|cernens autem Rahel quod infecunda esset invidit sorori et ait marito suo da mihi liberos alioquin moriar
GEN|30|2|cui iratus respondit Iacob num pro Deo ego sum qui privavit te fructu ventris tui
GEN|30|3|at illa habeo inquit famulam Balam ingredere ad eam ut pariat super genua mea et habeam ex ea filios
GEN|30|4|deditque illi Balam in coniugium quae
GEN|30|5|ingresso ad se viro concepit et peperit filium
GEN|30|6|dixitque Rahel iudicavit mihi Dominus et exaudivit vocem meam dans mihi filium et idcirco appellavit nomen illius Dan
GEN|30|7|rursumque Bala concipiens peperit alterum
GEN|30|8|pro quo ait Rahel conparavit me Deus cum sorore mea et invalui vocavitque eum Nepthalim
GEN|30|9|sentiens Lia quod parere desisset Zelpham ancillam suam marito tradidit
GEN|30|10|qua post conceptum edente filium
GEN|30|11|dixit feliciter et idcirco vocavit nomen eius Gad
GEN|30|12|peperit quoque Zelpha alterum
GEN|30|13|dixitque Lia hoc pro beatitudine mea beatam quippe me dicent mulieres propterea appellavit eum Aser
GEN|30|14|egressus autem Ruben tempore messis triticeae in agro repperit mandragoras quos matri Liae detulit dixitque Rahel da mihi partem de mandragoris filii tui
GEN|30|15|illa respondit parumne tibi videtur quod praeripueris maritum mihi nisi etiam mandragoras filii mei tuleris ait Rahel dormiat tecum hac nocte pro mandragoris filii tui
GEN|30|16|redeuntique ad vesperam de agro Iacob egressa est in occursum Lia et ad me inquit intrabis quia mercede conduxi te pro mandragoris filii mei dormivit cum ea nocte illa
GEN|30|17|et exaudivit Deus preces eius concepitque et peperit filium quintum
GEN|30|18|et ait dedit Deus mercedem mihi quia dedi ancillam meam viro meo appellavitque nomen illius Isachar
GEN|30|19|rursum Lia concipiens peperit sextum filium
GEN|30|20|et ait ditavit me Deus dote bona etiam hac vice mecum erit maritus meus eo quod genuerim ei sex filios et idcirco appellavit nomen eius Zabulon
GEN|30|21|post quem peperit filiam nomine Dinam
GEN|30|22|recordatus quoque Dominus Rahelis exaudivit eam et aperuit vulvam illius
GEN|30|23|quae concepit et peperit filium dicens abstulit Deus obprobrium meum
GEN|30|24|et vocavit nomen illius Ioseph dicens addat mihi Dominus filium alterum
GEN|30|25|nato autem Ioseph dixit Iacob socero suo dimitte me ut revertar in patriam et ad terram meam
GEN|30|26|da mihi uxores et liberos meos pro quibus servivi tibi ut abeam tu nosti servitutem qua servivi tibi
GEN|30|27|ait ei Laban inveniam gratiam in conspectu tuo experimento didici quod benedixerit mihi Deus propter te
GEN|30|28|constitue mercedem tuam quam dem tibi
GEN|30|29|at ille respondit tu nosti quomodo servierim tibi et quanta in manibus meis fuerit possessio tua
GEN|30|30|modicum habuisti antequam venirem et nunc dives effectus es benedixitque tibi Dominus ad introitum meum iustum est igitur ut aliquando provideam etiam domui meae
GEN|30|31|dixitque Laban quid dabo tibi at ille ait nihil volo sed si feceris quod postulo iterum pascam et custodiam pecora tua
GEN|30|32|gyra omnes greges tuos et separa cunctas oves varias et sparso vellere et quodcumque furvum et maculosum variumque fuerit tam in ovibus quam in capris erit merces mea
GEN|30|33|respondebitque mihi cras iustitia mea quando placiti tempus advenerit coram te et omnia quae non fuerint varia et maculosa et furva tam in ovibus quam in capris furti me arguent
GEN|30|34|dixit Laban gratum habeo quod petis
GEN|30|35|et separavit in die illo capras et oves hircos et arietes varios atque maculosos cunctum autem gregem unicolorem id est albi et nigri velleris tradidit in manu filiorum suorum
GEN|30|36|et posuit spatium itineris inter se et generum dierum trium qui pascebat reliquos greges eius
GEN|30|37|tollens ergo Iacob virgas populeas virides et amigdalinas et ex platanis ex parte decorticavit eas detractisque corticibus in his quae spoliata fuerant candor apparuit illa vero quae integra erant viridia permanserunt atque in hunc modum color effectus est varius
GEN|30|38|posuitque eas in canalibus ubi effundebatur aqua ut cum venissent greges ad bibendum ante oculos haberent virgas et in aspectu earum conciperent
GEN|30|39|factumque est ut in ipso calore coitus oves intuerentur virgas et parerent maculosa et varia et diverso colore respersa
GEN|30|40|divisitque gregem Iacob et posuit virgas ante oculos arietum erant autem alba quaeque et nigra Laban cetera vero Iacob separatis inter se gregibus
GEN|30|41|igitur quando primo tempore ascendebantur oves ponebat Iacob virgas in canalibus aquarum ante oculos arietum et ovium ut in earum contemplatione conciperent
GEN|30|42|quando vero serotina admissura erat et conceptus extremus non ponebat eas factaque sunt ea quae erant serotina Laban et quae primi temporis Iacob
GEN|30|43|ditatusque est homo ultra modum et habuit greges multos ancillas et servos camelos et asinos
GEN|31|1|postquam autem audivit verba filiorum Laban dicentium tulit Iacob omnia quae fuerunt patris nostri et de illius facultate ditatus factus est inclitus
GEN|31|2|animadvertit quoque faciem Laban quod non esset erga se sicut heri et nudius tertius
GEN|31|3|maxime dicente sibi Domino revertere in terram patrum tuorum et ad generationem tuam eroque tecum
GEN|31|4|misit et vocavit Rahel et Liam in agrum ubi pascebat greges
GEN|31|5|dixitque eis video faciem patris vestri quod non sit erga me sicut heri et nudius tertius Deus autem patris mei fuit mecum
GEN|31|6|et ipsae nostis quod totis viribus meis servierim patri vestro
GEN|31|7|sed pater vester circumvenit me et mutavit mercedem meam decem vicibus et tamen non dimisit eum Deus ut noceret mihi
GEN|31|8|si quando dixit variae erunt mercedes tuae pariebant omnes oves varios fetus quando vero e contrario ait alba quaeque accipies pro mercede omnes greges alba pepererunt
GEN|31|9|tulitque Deus substantiam patris vestri et dedit mihi
GEN|31|10|postquam enim conceptus ovium tempus advenerat levavi oculos meos et vidi in somnis ascendentes mares super feminas varios et maculosos et diversorum colorum
GEN|31|11|dixitque angelus Dei ad me in somnis Iacob et ego respondi adsum
GEN|31|12|qui ait leva oculos tuos et vide universos masculos ascendentes super feminas varios respersos atque maculosos vidi enim omnia quae fecit tibi Laban
GEN|31|13|ego sum Deus Bethel ubi unxisti lapidem et votum vovisti mihi nunc ergo surge et egredere de terra hac revertens in terram nativitatis tuae
GEN|31|14|responderunt Rahel et Lia numquid habemus residui quicquam in facultatibus et hereditate domus patris nostri
GEN|31|15|nonne quasi alienas reputavit nos et vendidit comeditque pretium nostrum
GEN|31|16|sed Deus tulit opes patris nostri et nobis eas tradidit ac filiis nostris unde omnia quae praecepit fac
GEN|31|17|surrexit itaque Iacob et inpositis liberis et coniugibus suis super camelos abiit
GEN|31|18|tulitque omnem substantiam et greges et quicquid in Mesopotamiam quaesierat pergens ad Isaac patrem suum in terram Chanaan
GEN|31|19|eo tempore Laban ierat ad tondendas oves et Rahel furata est idola patris sui
GEN|31|20|noluitque Iacob confiteri socero quod fugeret
GEN|31|21|cumque abisset tam ipse quam omnia quae iuris eius erant et amne transmisso pergeret contra montem Galaad
GEN|31|22|nuntiatum est Laban die tertio quod fugeret Iacob
GEN|31|23|qui adsumptis fratribus suis persecutus est eum diebus septem et conprehendit in monte Galaad
GEN|31|24|viditque in somnis dicentem sibi Dominum cave ne quicquam aspere loquaris contra Iacob
GEN|31|25|iamque Iacob extenderat in monte tabernaculum cum ille consecutus eum cum fratribus suis in eodem monte Galaad fixit tentorium
GEN|31|26|et dixit ad Iacob quare ita egisti ut clam me abigeres filias meas quasi captivas gladio
GEN|31|27|cur ignorante me fugere voluisti nec indicare mihi ut prosequerer te cum gaudio et canticis et tympanis et cithara
GEN|31|28|non es passus ut oscularer filios meos ac filias stulte operatus es et nunc
GEN|31|29|valet quidem manus mea reddere tibi malum sed Deus patris vestri heri dixit mihi cave ne loquaris cum Iacob quicquam durius
GEN|31|30|esto ad tuos ire cupiebas et desiderio tibi erat domus patris tui cur furatus es deos meos
GEN|31|31|respondit Iacob quod inscio te profectus sum timui ne violenter auferres filias tuas
GEN|31|32|quod autem furti arguis apud quemcumque inveneris deos tuos necetur coram fratribus nostris scrutare quicquid tuorum apud me inveneris et aufer haec dicens ignorabat quod Rahel furata esset idola
GEN|31|33|ingressus itaque Laban tabernaculum Iacob et Liae et utriusque famulae non invenit cumque intrasset tentorium Rahelis
GEN|31|34|illa festinans abscondit idola subter stramen cameli et sedit desuper scrutantique omne tentorium et nihil invenienti
GEN|31|35|ait ne irascatur dominus meus quod coram te adsurgere nequeo quia iuxta consuetudinem feminarum nunc accidit mihi sic delusa sollicitudo quaerentis est
GEN|31|36|tumensque Iacob cum iurgio ait quam ob culpam meam et ob quod peccatum sic exarsisti post me
GEN|31|37|et scrutatus es omnem supellectilem meam quid invenisti de cuncta substantia domus tuae pone hic coram fratribus meis et fratribus tuis et iudicent inter me et te
GEN|31|38|idcirco viginti annis fui tecum oves tuae et caprae steriles non fuerunt arietes gregis tui non comedi
GEN|31|39|nec captum a bestia ostendi tibi ego damnum omne reddebam quicquid furto perierat a me exigebas
GEN|31|40|die noctuque aestu urebar et gelu fugiebat somnus ab oculis meis
GEN|31|41|sic per viginti annos in domo tua servivi tibi quattuordecim pro filiabus et sex pro gregibus tuis inmutasti quoque mercedem meam decem vicibus
GEN|31|42|nisi Deus patris mei Abraham et Timor Isaac adfuisset mihi forsitan modo nudum me dimisisses adflictionem meam et laborem manuum mearum respexit Deus et arguit te heri
GEN|31|43|respondit ei Laban filiae et filii et greges tui et omnia quae cernis mea sunt quid possum facere filiis et nepotibus meis
GEN|31|44|veni ergo et ineamus foedus ut sit testimonium inter me et te
GEN|31|45|tulit itaque Iacob lapidem et erexit illum in titulum
GEN|31|46|dixitque fratribus suis adferte lapides qui congregantes fecerunt tumulum comederuntque super eum
GEN|31|47|quem vocavit Laban tumulus Testis et Iacob acervum Testimonii uterque iuxta proprietatem linguae suae
GEN|31|48|dixitque Laban tumulus iste testis erit inter me et te hodie et idcirco appellatum est nomen eius Galaad id est tumulus Testis
GEN|31|49|intueatur Dominus et iudicet inter nos quando recesserimus a nobis
GEN|31|50|si adflixeris filias meas et si introduxeris uxores alias super eas nullus sermonis nostri testis est absque Deo qui praesens respicit
GEN|31|51|dixitque rursus ad Iacob en tumulus hic et lapis quem erexi inter me et te
GEN|31|52|testis erit tumulus inquam iste et lapis sint in testimonio si aut ego transiero illum pergens ad te aut tu praeterieris malum mihi cogitans
GEN|31|53|Deus Abraham et Deus Nahor iudicet inter nos Deus patris eorum iuravit Iacob per Timorem patris sui Isaac
GEN|31|54|immolatisque victimis in monte vocavit fratres suos ut ederent panem qui cum comedissent manserunt ibi
GEN|31|55|Laban vero de nocte consurgens osculatus est filios et filias suas et benedixit illis reversus in locum suum
GEN|32|1|Iacob quoque abiit itinere quo coeperat fueruntque ei obviam angeli Dei
GEN|32|2|quos cum vidisset ait castra Dei sunt haec et appellavit nomen loci illius Manaim id est Castra
GEN|32|3|misit autem et nuntios ante se ad Esau fratrem suum in terram Seir regionis Edom
GEN|32|4|praecepitque eis dicens sic loquimini domino meo Esau haec dicit frater tuus Iacob apud Laban peregrinatus sum et fui usque in praesentem diem
GEN|32|5|habeo boves et asinos oves et servos atque ancillas mittoque nunc legationem ad dominum meum ut inveniam gratiam in conspectu tuo
GEN|32|6|reversi sunt nuntii ad Iacob dicentes venimus ad Esau fratrem tuum et ecce properat in occursum tibi cum quadringentis viris
GEN|32|7|timuit Iacob valde et perterritus divisit populum qui secum erat greges quoque et oves et boves et camelos in duas turmas
GEN|32|8|dicens si venerit Esau ad unam turmam et percusserit eam alia turma quae reliqua est salvabitur
GEN|32|9|dixitque Iacob Deus patris mei Abraham et Deus patris mei Isaac Domine qui dixisti mihi revertere in terram tuam et in locum nativitatis tuae et benefaciam tibi
GEN|32|10|minor sum cunctis miserationibus et veritate quam explesti servo tuo in baculo meo transivi Iordanem istum et nunc cum duabus turmis regredior
GEN|32|11|erue me de manu fratris mei de manu Esau quia valde eum timeo ne forte veniens percutiat matrem cum filiis
GEN|32|12|tu locutus es quod bene mihi faceres et dilatares semen meum sicut harenam maris quae prae multitudine numerari non potest
GEN|32|13|cumque dormisset ibi nocte illa separavit de his quae habebat munera Esau fratri suo
GEN|32|14|capras ducentas hircos viginti oves ducentas arietes viginti
GEN|32|15|camelos fetas cum pullis suis triginta vaccas quadraginta et tauros viginti asinas viginti et pullos earum decem
GEN|32|16|et misit per manus servorum suorum singulos seorsum greges dixitque pueris suis antecedite me et sit spatium inter gregem et gregem
GEN|32|17|et praecepit priori dicens si obvium habueris Esau fratrem meum et interrogaverit te cuius es et quo vadis et cuius sunt ista quae sequeris
GEN|32|18|respondebis servi tui Iacob munera misit domino meo Esau ipse quoque post nos venit
GEN|32|19|similiter mandata dedit secundo ac tertio et cunctis qui sequebantur greges dicens hisdem verbis loquimini ad Esau cum inveneritis eum
GEN|32|20|et addetis ipse quoque servus tuus Iacob iter nostrum insequitur dixit enim placabo illum muneribus quae praecedunt et postea videbo forsitan propitiabitur mihi
GEN|32|21|praecesserunt itaque munera ante eum ipse vero mansit nocte illa in Castris
GEN|32|22|cumque mature surrexisset tulit duas uxores suas et totidem famulas cum undecim filiis et transivit vadum Iaboc
GEN|32|23|transductisque omnibus quae ad se pertinebant
GEN|32|24|remansit solus et ecce vir luctabatur cum eo usque mane
GEN|32|25|qui cum videret quod eum superare non posset tetigit nervum femoris eius et statim emarcuit
GEN|32|26|dixitque ad eum dimitte me iam enim ascendit aurora respondit non dimittam te nisi benedixeris mihi
GEN|32|27|ait ergo quod nomen est tibi respondit Iacob
GEN|32|28|at ille nequaquam inquit Iacob appellabitur nomen tuum sed Israhel quoniam si contra Deum fortis fuisti quanto magis contra homines praevalebis
GEN|32|29|interrogavit eum Iacob dic mihi quo appellaris nomine respondit cur quaeris nomen meum et benedixit ei in eodem loco
GEN|32|30|vocavitque Iacob nomen loci illius Phanuhel dicens vidi Deum facie ad faciem et salva facta est anima mea
GEN|32|31|ortusque est ei statim sol postquam transgressus est Phanuhel ipse vero claudicabat pede
GEN|32|32|quam ob causam non comedunt filii Israhel nervum qui emarcuit in femore Iacob usque in praesentem diem eo quod tetigerit nervum femoris eius et obstipuerit
GEN|33|1|levans autem Iacob oculos suos vidit venientem Esau et cum eo quadringentos viros divisitque filios Liae et Rahel ambarumque famularum
GEN|33|2|et posuit utramque ancillam et liberos earum in principio Liam vero et filios eius in secundo loco Rahel autem et Ioseph novissimos
GEN|33|3|et ipse praegrediens adoravit pronus in terram septies donec adpropinquaret frater eius
GEN|33|4|currens itaque Esau obviam fratri suo amplexatus est eum stringensque collum et osculans flevit
GEN|33|5|levatisque oculis vidit mulieres et parvulos earum et ait quid sibi volunt isti et si ad te pertinent respondit parvuli sunt quos donavit mihi Deus servo tuo
GEN|33|6|et adpropinquantes ancillae et filii earum incurvati sunt
GEN|33|7|accessitque Lia cum liberis suis et cum similiter adorassent extremi Ioseph et Rahel adoraverunt
GEN|33|8|quaenam sunt inquit istae turmae quas obvias habui respondit ut invenirem gratiam coram domino meo
GEN|33|9|et ille habeo ait plurima frater mi sint tua tibi
GEN|33|10|dixit Iacob noli ita obsecro sed si inveni gratiam in oculis tuis accipe munusculum de manibus meis sic enim vidi faciem tuam quasi viderim vultum Dei esto mihi propitius
GEN|33|11|et suscipe benedictionem quam adtuli tibi et quam donavit mihi Deus tribuens omnia vix fratre conpellente suscipiens
GEN|33|12|ait gradiamur simul eroque socius itineris tui
GEN|33|13|dixit Iacob nosti domine mi quod parvulos habeam teneros et oves ac boves fetas mecum quas si plus in ambulando fecero laborare morientur una die cuncti greges
GEN|33|14|praecedat dominus meus ante servum suum et ego sequar paulatim vestigia eius sicut videro posse parvulos meos donec veniam ad dominum meum in Seir
GEN|33|15|respondit Esau oro te ut de populo qui mecum est saltem socii remaneant viae tuae non est inquit necesse hoc uno indigeo ut inveniam gratiam in conspectu domini mei
GEN|33|16|reversus est itaque illo die Esau itinere quo venerat in Seir
GEN|33|17|et Iacob venit in Soccoth ubi aedificata domo et fixis tentoriis appellavit nomen loci illius Soccoth id est Tabernacula
GEN|33|18|transivitque in Salem urbem Sycimorum quae est in terra Chanaan postquam regressus est de Mesopotamiam Syriae et habitavit iuxta oppidum
GEN|33|19|emitque partem agri in qua fixerat tabernaculum a filiis Emor patris Sychem centum agnis
GEN|33|20|et erecto ibi altari invocavit super illud Fortissimum Deum Israhel
GEN|34|1|egressa est autem Dina filia Liae ut videret mulieres regionis illius
GEN|34|2|quam cum vidisset Sychem filius Emor Evei princeps terrae illius adamavit et rapuit et dormivit cum illa vi opprimens virginem
GEN|34|3|et conglutinata est anima eius cum ea tristemque blanditiis delinivit
GEN|34|4|et pergens ad Emor patrem suum accipe mihi inquit puellam hanc coniugem
GEN|34|5|quod cum audisset Iacob absentibus filiis et in pastu occupatis pecorum siluit donec redirent
GEN|34|6|egresso autem Emor patre Sychem ut loqueretur ad Iacob
GEN|34|7|ecce filii eius veniebant de agro auditoque quod acciderat irati sunt valde eo quod foedam rem esset operatus in Israhel et violata filia Iacob rem inlicitam perpetrasset
GEN|34|8|locutus est itaque Emor ad eos Sychem filii mei adhesit anima filiae vestrae date eam illi uxorem
GEN|34|9|et iungamus vicissim conubia filias vestras tradite nobis et filias nostras accipite
GEN|34|10|et habitate nobiscum terra in potestate vestra est exercete negotiamini et possidete eam
GEN|34|11|sed et Sychem ad patrem et ad fratres eius ait inveniam gratiam coram vobis et quaecumque statueritis dabo
GEN|34|12|augete dotem munera postulate libens tribuam quod petieritis tantum date mihi puellam hanc uxorem
GEN|34|13|responderunt filii Iacob Sychem et patri eius in dolo saevientes ob stuprum sororis
GEN|34|14|non possumus facere quod petitis nec dare sororem nostram homini incircumciso quod inlicitum et nefarium est apud nos
GEN|34|15|sed in hoc valebimus foederari si esse volueritis nostri similes et circumcidatur in vobis omne masculini sexus
GEN|34|16|tunc dabimus et accipiemus mutuo filias nostras ac vestras et habitabimus vobiscum erimusque unus populus
GEN|34|17|sin autem circumcidi nolueritis tollemus filiam nostram et recedemus
GEN|34|18|placuit oblatio eorum Emor et Sychem filio eius
GEN|34|19|nec distulit adulescens quin statim quod petebatur expleret amabat enim puellam valde et ipse erat inclitus in omni domo patris sui
GEN|34|20|ingressique portam urbis locuti sunt populo
GEN|34|21|viri isti pacifici sunt et volunt habitare nobiscum negotientur in terra et exerceant eam quae spatiosa et lata cultoribus indiget filias eorum accipiemus uxores et nostras illis dabimus
GEN|34|22|unum est quod differtur tantum bonum si circumcidamus masculos nostros ritum gentis imitantes
GEN|34|23|et substantia eorum et pecora et cuncta quae possident nostra erunt tantum in hoc adquiescamus et habitantes simul unum efficiemus populum
GEN|34|24|adsensi sunt omnes circumcisis cunctis maribus
GEN|34|25|et ecce die tertio quando gravissimus vulnerum dolor est arreptis duo Iacob filii Symeon et Levi fratres Dinae gladiis ingressi sunt urbem confidenter interfectisque omnibus masculis
GEN|34|26|Emor et Sychem pariter necaverunt tollentes Dinam de domo Sychem sororem suam
GEN|34|27|quibus egressis inruerunt super occisos ceteri filii Iacob et depopulati sunt urbem in ultionem stupri
GEN|34|28|oves eorum et armenta et asinos cunctaque vastantes quae in domibus et in agris erant
GEN|34|29|parvulos quoque et uxores eorum duxere captivas
GEN|34|30|quibus patratis audacter Iacob dixit ad Symeon et Levi turbastis me et odiosum fecistis Chananeis et Ferezeis habitatoribus terrae huius nos pauci sumus illi congregati percutient me et delebor ego et domus mea
GEN|34|31|responderunt numquid ut scorto abuti debuere sorore nostra
GEN|35|1|interea locutus est Deus ad Iacob surge et ascende Bethel et habita ibi facque altare Deo qui apparuit tibi quando fugiebas Esau fratrem tuum
GEN|35|2|Iacob vero convocata omni domo sua ait abicite deos alienos qui in medio vestri sunt et mundamini ac mutate vestimenta vestra
GEN|35|3|surgite et ascendamus in Bethel ut faciamus ibi altare Deo qui exaudivit me in die tribulationis meae et fuit socius itineris mei
GEN|35|4|dederunt ergo ei omnes deos alienos quos habebant et inaures quae erant in auribus eorum at ille infodit ea subter terebinthum quae est post urbem Sychem
GEN|35|5|cumque profecti essent terror Dei invasit omnes per circuitum civitates et non sunt ausi persequi recedentes
GEN|35|6|venit igitur Iacob Luzam quae est in terra Chanaan cognomento Bethel ipse et omnis populus cum eo
GEN|35|7|aedificavitque ibi altare et appellavit nomen loci Domus Dei ibi enim apparuit ei Deus cum fugeret fratrem suum
GEN|35|8|eodem tempore mortua est Debbora nutrix Rebeccae et sepulta ad radices Bethel subter quercum vocatumque est nomen loci quercus Fletus
GEN|35|9|apparuit autem iterum Deus Iacob postquam reversus est de Mesopotamiam Syriae benedixitque ei
GEN|35|10|dicens non vocaberis ultra Iacob sed Israhel erit nomen tuum et appellavit eum Israhel
GEN|35|11|dixitque ei ego Deus omnipotens cresce et multiplicare gentes et populi nationum erunt ex te reges de lumbis tuis egredientur
GEN|35|12|terramque quam dedi Abraham et Isaac dabo tibi et semini tuo post te
GEN|35|13|et recessit ab eo
GEN|35|14|ille vero erexit titulum lapideum in loco quo locutus ei fuerat Deus libans super eum libamina et effundens oleum
GEN|35|15|vocansque nomen loci Bethel
GEN|35|16|egressus inde venit verno tempore ad terram quae ducit Efratham in qua cum parturiret Rahel
GEN|35|17|ob difficultatem partus periclitari coepit dixitque ei obsetrix noli timere quia et hunc habebis filium
GEN|35|18|egrediente autem anima prae dolore et inminente iam morte vocavit nomen filii sui Benoni id est filius doloris mei pater vero appellavit eum Beniamin id est filius dexterae
GEN|35|19|mortua est ergo Rahel et sepulta in via quae ducit Efratham haec est Bethleem
GEN|35|20|erexitque Iacob titulum super sepulchrum eius hic est titulus monumenti Rahel usque in praesentem diem
GEN|35|21|egressus inde fixit tabernaculum trans turrem Gregis
GEN|35|22|cumque habitaret in illa regione abiit Ruben et dormivit cum Bala concubina patris sui quod illum minime latuit erant autem filii Iacob duodecim
GEN|35|23|filii Liae primogenitus Ruben et Symeon et Levi et Iudas et Isachar et Zabulon
GEN|35|24|filii Rahel Ioseph et Beniamin
GEN|35|25|filii Balae ancillae Rahelis Dan et Nepthalim
GEN|35|26|filii Zelphae ancillae Liae Gad et Aser hii filii Iacob qui nati sunt ei in Mesopotamiam Syriae
GEN|35|27|venit etiam ad Isaac patrem suum in Mambre civitatem Arbee haec est Hebron in qua peregrinatus est Abraham et Isaac
GEN|35|28|et conpleti sunt dies Isaac centum octoginta annorum
GEN|35|29|consumptusque aetate mortuus est et adpositus populo suo senex et plenus dierum et sepelierunt eum Esau et Iacob filii sui
GEN|36|1|hae sunt autem generationes Esau ipse est Edom
GEN|36|2|Esau accepit uxores de filiabus Chanaan Ada filiam Elom Hetthei et Oolibama filiam Anae filiae Sebeon Evei
GEN|36|3|Basemath quoque filiam Ismahel sororem Nabaioth
GEN|36|4|peperit autem Ada Eliphaz Basemath genuit Rauhel
GEN|36|5|Oolibama edidit Hieus et Hielom et Core hii filii Esau qui nati sunt ei in terra Chanaan
GEN|36|6|tulit autem Esau uxores suas et filios et filias et omnem animam domus suae et substantiam et pecora et cuncta quae habere poterat in terra Chanaan et abiit in alteram regionem recessitque a fratre suo Iacob
GEN|36|7|divites enim erant valde et simul habitare non poterant nec sustinebat eos terra peregrinationis eorum prae multitudine gregum
GEN|36|8|habitavitque Esau in monte Seir ipse est Edom
GEN|36|9|hae sunt generationes Esau patris Edom in monte Seir
GEN|36|10|et haec nomina filiorum eius Eliphaz filius Ada uxoris Esau Rauhel quoque filius Basemath uxoris eius
GEN|36|11|fueruntque filii Eliphaz Theman Omar Sephu et Gatham et Cenez
GEN|36|12|erat autem Thamna concubina Eliphaz filii Esau quae peperit ei Amalech hii sunt filii Adae uxoris Esau
GEN|36|13|filii autem Rauhel Naath et Zara Semma et Meza hii filii Basemath uxoris Esau
GEN|36|14|isti quoque erant filii Oolibama filiae Ana filiae Sebeon uxoris Esau quos genuit ei Hieus et Hielom et Core
GEN|36|15|hii duces filiorum Esau filii Eliphaz primogeniti Esau dux Theman dux Omar dux Sephu dux Cenez
GEN|36|16|dux Core dux Gatham dux Amalech hii filii Eliphaz in terra Edom et hii filii Adae
GEN|36|17|hii quoque filii Rauhel filii Esau dux Naath dux Zara dux Semma dux Meza hii duces Rauhel in terra Edom isti filii Basemath uxoris Esau
GEN|36|18|hii autem filii Oolibama uxoris Esau dux Hieus dux Hielom dux Core hii duces Oolibama filiae Ana uxoris Esau
GEN|36|19|isti filii Esau et hii duces eorum ipse est Edom
GEN|36|20|isti filii Seir Horrei habitatores terrae Lotham et Sobal et Sebeon et Anan
GEN|36|21|Dison et Eser et Disan hii duces Horrei filii Seir in terra Edom
GEN|36|22|facti sunt autem filii Lotham Horrei et Heman erat autem soror Lotham Thamna
GEN|36|23|et isti filii Sobal Alvam et Maneeth et Hebal Sephi et Onam
GEN|36|24|et hii filii Sebeon Ahaia et Anam iste est Ana qui invenit aquas calidas in solitudine cum pasceret asinos Sebeon patris sui
GEN|36|25|habuitque filium Disan et filiam Oolibama
GEN|36|26|et isti filii Disan Amdan et Esban et Iethran et Charan
GEN|36|27|hii quoque filii Eser Balaan et Zevan et Acham
GEN|36|28|habuit autem filios Disan Hus et Aran
GEN|36|29|isti duces Horreorum dux Lothan dux Sobal dux Sebeon dux Ana
GEN|36|30|dux Dison dux Eser dux Disan isti duces Horreorum qui imperaverunt in terra Seir
GEN|36|31|reges autem qui regnaverunt in terra Edom antequam haberent regem filii Israhel fuerunt hii
GEN|36|32|Bale filius Beor nomenque urbis eius Denaba
GEN|36|33|mortuus est autem Bale et regnavit pro eo Iobab filius Zare de Bosra
GEN|36|34|cumque mortuus esset Iobab regnavit pro eo Husan de terra Themanorum
GEN|36|35|hoc quoque mortuo regnavit pro eo Adad filius Badadi qui percussit Madian in regione Moab et nomen urbis eius Ahuith
GEN|36|36|cumque mortuus esset Adad regnavit pro eo Semla de Maserecha
GEN|36|37|hoc quoque mortuo regnavit pro eo Saul de fluvio Rooboth
GEN|36|38|cumque et hic obisset successit in regnum Baalanam filius Achobor
GEN|36|39|isto quoque mortuo regnavit pro eo Adad nomenque urbis eius Phau et appellabatur uxor illius Meezabel filia Matred filiae Mizaab
GEN|36|40|haec ergo nomina Esau in cognationibus et locis et vocabulis suis dux Thamna dux Alva dux Ietheth
GEN|36|41|dux Oolibama dux Ela dux Phinon
GEN|36|42|dux Cenez dux Theman dux Mabsar
GEN|36|43|dux Mabdiel dux Iram hii duces Edom habitantes in terra imperii sui ipse est Esau pater Idumeorum
GEN|37|1|habitavit autem Iacob in terra Chanaan in qua peregrinatus est pater suus
GEN|37|2|et hae sunt generationes eius Ioseph cum sedecim esset annorum pascebat gregem cum fratribus suis adhuc puer et erat cum filiis Balae et Zelphae uxorum patris sui accusavitque fratres suos apud patrem crimine pessimo
GEN|37|3|Israhel autem diligebat Ioseph super omnes filios suos eo quod in senectute genuisset eum fecitque ei tunicam polymitam
GEN|37|4|videntes autem fratres eius quod a patre plus cunctis filiis amaretur oderant eum nec poterant ei quicquam pacificum loqui
GEN|37|5|accidit quoque ut visum somnium referret fratribus quae causa maioris odii seminarium fuit
GEN|37|6|dixitque ad eos audite somnium meum quod vidi
GEN|37|7|putabam ligare nos manipulos in agro et quasi consurgere manipulum meum et stare vestrosque manipulos circumstantes adorare manipulum meum
GEN|37|8|responderunt fratres eius numquid rex noster eris aut subiciemur dicioni tuae haec ergo causa somniorum atque sermonum invidiae et odii fomitem ministravit
GEN|37|9|aliud quoque vidit somnium quod narrans fratribus ait vidi per somnium quasi solem et lunam et stellas undecim adorare me
GEN|37|10|quod cum patri suo et fratribus rettulisset increpavit eum pater et dixit quid sibi vult hoc somnium quod vidisti num ego et mater tua et fratres adorabimus te super terram
GEN|37|11|invidebant igitur ei fratres sui pater vero rem tacitus considerabat
GEN|37|12|cumque fratres illius in pascendis gregibus patris morarentur in Sychem
GEN|37|13|dixit ad eum Israhel fratres tui pascunt oves in Sycimis veni mittam te ad eos quo respondente
GEN|37|14|praesto sum ait vade et vide si cuncta prospera sint erga fratres tuos et pecora et renuntia mihi quid agatur missus de valle Hebron venit in Sychem
GEN|37|15|invenitque eum vir errantem in agro et interrogavit quid quaereret
GEN|37|16|at ille respondit fratres meos quaero indica mihi ubi pascant greges
GEN|37|17|dixitque ei vir recesserunt de loco isto audivi autem eos dicentes eamus in Dothain perrexit ergo Ioseph post fratres suos et invenit eos in Dothain
GEN|37|18|qui cum vidissent eum procul antequam accederet ad eos cogitaverunt illum occidere
GEN|37|19|et mutuo loquebantur ecce somniator venit
GEN|37|20|venite occidamus eum et mittamus in cisternam veterem dicemusque fera pessima devoravit eum et tunc apparebit quid illi prosint somnia sua
GEN|37|21|audiens hoc Ruben nitebatur liberare eum de manibus eorum et dicebat
GEN|37|22|non interficiamus animam eius nec effundatis sanguinem sed proicite eum in cisternam hanc quae est in solitudine manusque vestras servate innoxias hoc autem dicebat volens eripere eum de manibus eorum et reddere patri suo
GEN|37|23|confestim igitur ut pervenit ad fratres nudaverunt eum tunica talari et polymita
GEN|37|24|miseruntque in cisternam quae non habebat aquam
GEN|37|25|et sedentes ut comederent panem viderunt viatores Ismahelitas venire de Galaad et camelos eorum portare aromata et resinam et stacten in Aegyptum
GEN|37|26|dixit ergo Iudas fratribus suis quid nobis prodest si occiderimus fratrem nostrum et celaverimus sanguinem ipsius
GEN|37|27|melius est ut vendatur Ismahelitis et manus nostrae non polluantur frater enim et caro nostra est adquieverunt fratres sermonibus eius
GEN|37|28|et praetereuntibus Madianitis negotiatoribus extrahentes eum de cisterna vendiderunt Ismahelitis viginti argenteis qui duxerunt eum in Aegyptum
GEN|37|29|reversusque Ruben ad cisternam non invenit puerum
GEN|37|30|et scissis vestibus pergens ad fratres ait puer non conparet et ego quo ibo
GEN|37|31|tulerunt autem tunicam eius et in sanguinem hedi quem occiderant tinxerunt
GEN|37|32|mittentes qui ferrent ad patrem et dicerent hanc invenimus vide utrum tunica filii tui sit an non
GEN|37|33|quam cum agnovisset pater ait tunica filii mei est fera pessima comedit eum bestia devoravit Ioseph
GEN|37|34|scissisque vestibus indutus est cilicio lugens filium multo tempore
GEN|37|35|congregatis autem cunctis liberis eius ut lenirent dolorem patris noluit consolationem recipere et ait descendam ad filium meum lugens in infernum et illo perseverante in fletu
GEN|37|36|Madianei vendiderunt Ioseph in Aegypto Putiphar eunucho Pharaonis magistro militiae
GEN|38|1|eo tempore descendens Iudas a fratribus suis divertit ad virum odollamitem nomine Hiram
GEN|38|2|viditque ibi filiam hominis chananei vocabulo Suae et uxore accepta ingressus est ad eam
GEN|38|3|quae concepit et peperit filium vocavitque nomen eius Her
GEN|38|4|rursum concepto fetu natum filium nominavit Onam
GEN|38|5|tertium quoque peperit quem appellavit Sela quo nato parere ultra cessavit
GEN|38|6|dedit autem Iudas uxorem primogenito suo Her nomine Thamar
GEN|38|7|fuitque Her primogenitus Iudae nequam in conspectu Domini et ab eo occisus est
GEN|38|8|dixit ergo Iudas ad Onam filium suum ingredere ad uxorem fratris tui et sociare illi ut suscites semen fratri tuo
GEN|38|9|ille sciens non sibi nasci filios introiens ad uxorem fratris sui semen fundebat in terram ne liberi fratris nomine nascerentur
GEN|38|10|et idcirco percussit eum Dominus quod rem detestabilem faceret
GEN|38|11|quam ob rem dixit Iudas Thamar nurui suae esto vidua in domo patris tui donec crescat Sela filius meus timebat enim ne et ipse moreretur sicut fratres eius quae abiit et habitavit in domo patris sui
GEN|38|12|evolutis autem multis diebus mortua est filia Suae uxor Iudae qui post luctum consolatione suscepta ascendebat ad tonsores ovium suarum ipse et Hiras opilio gregis Odollamita in Thamnas
GEN|38|13|nuntiatumque est Thamar quod socer illius ascenderet in Thamnas ad tondendas oves
GEN|38|14|quae depositis viduitatis vestibus adsumpsit theristrum et mutato habitu sedit in bivio itineris quod ducit Thamnam eo quod crevisset Sela et non eum accepisset maritum
GEN|38|15|quam cum vidisset Iudas suspicatus est esse meretricem operuerat enim vultum suum ne cognosceretur
GEN|38|16|ingrediensque ad eam ait dimitte me ut coeam tecum nesciebat enim quod nurus sua esset qua respondente quid mihi dabis ut fruaris concubitu meo
GEN|38|17|dixit mittam tibi hedum de gregibus rursum illa dicente patiar quod vis si dederis mihi arrabonem donec mittas quod polliceris
GEN|38|18|ait Iudas quid vis tibi pro arrabone dari respondit anulum tuum et armillam et baculum quem manu tenes ad unum igitur coitum concepit mulier
GEN|38|19|et surgens abiit depositoque habitu quem adsumpserat induta est viduitatis vestibus
GEN|38|20|misit autem Iudas hedum per pastorem suum Odollamitem ut reciperet pignus quod dederat mulieri qui cum non invenisset eam
GEN|38|21|interrogavit homines loci illius ubi est mulier quae sedebat in bivio respondentibus cunctis non fuit in loco isto meretrix
GEN|38|22|reversus est ad Iudam et dixit ei non inveni eam sed et homines loci illius dixerunt mihi numquam ibi sedisse scortum
GEN|38|23|ait Iudas habeat sibi certe mendacii nos arguere non poterit ego misi hedum quem promiseram et tu non invenisti eam
GEN|38|24|ecce autem post tres menses nuntiaverunt Iudae dicentes fornicata est Thamar nurus tua et videtur uterus illius intumescere dixit Iudas producite eam ut conburatur
GEN|38|25|quae cum educeretur ad poenam misit ad socerum suum dicens de viro cuius haec sunt concepi cognosce cuius sit anulus et armilla et baculus
GEN|38|26|qui agnitis muneribus ait iustior me est quia non tradidi eam Sela filio meo attamen ultra non cognovit illam
GEN|38|27|instante autem partu apparuerunt gemini in utero atque in ipsa effusione infantum unus protulit manum in qua obsetrix ligavit coccinum dicens
GEN|38|28|iste egreditur prior
GEN|38|29|illo vero retrahente manum egressus est alter dixitque mulier quare divisa est propter te maceria et ob hanc causam vocavit nomen eius Phares
GEN|38|30|postea egressus est frater in cuius manu erat coccinum quem appellavit Zara
GEN|39|1|igitur Ioseph ductus est in Aegyptum emitque eum Putiphar eunuchus Pharaonis princeps exercitus vir aegyptius de manu Ismahelitarum a quibus perductus erat
GEN|39|2|fuitque Dominus cum eo et erat vir in cunctis prospere agens habitabatque in domo domini sui
GEN|39|3|qui optime noverat esse Dominum cum eo et omnia quae gereret ab eo dirigi in manu illius
GEN|39|4|invenitque Ioseph gratiam coram domino suo et ministrabat ei a quo praepositus omnibus gubernabat creditam sibi domum et universa quae tradita fuerant
GEN|39|5|benedixitque Dominus domui Aegyptii propter Ioseph et multiplicavit tam in aedibus quam in agris cunctam eius substantiam
GEN|39|6|nec quicquam aliud noverat nisi panem quo vescebatur erat autem Ioseph pulchra facie et decorus aspectu
GEN|39|7|post multos itaque dies iecit domina oculos suos in Ioseph et ait dormi mecum
GEN|39|8|qui nequaquam adquiescens operi nefario dixit ad eam ecce dominus meus omnibus mihi traditis ignorat quid habeat in domo sua
GEN|39|9|nec quicquam est quod non in mea sit potestate vel non tradiderit mihi praeter te quae uxor eius es quomodo ergo possum malum hoc facere et peccare in Deum meum
GEN|39|10|huiuscemodi verbis per singulos dies et mulier molesta erat adulescenti et ille recusabat stuprum
GEN|39|11|accidit autem ut quadam die intraret Ioseph domum et operis quippiam absque arbitris faceret
GEN|39|12|et illa adprehensa lacinia vestimenti eius diceret dormi mecum qui relicto in manu illius pallio fugit et egressus est foras
GEN|39|13|cumque vidisset mulier vestem in manibus suis et se esse contemptam
GEN|39|14|vocavit homines domus suae et ait ad eos en introduxit virum hebraeum ut inluderet nobis ingressus est ad me ut coiret mecum cumque ego succlamassem
GEN|39|15|et audisset vocem meam reliquit pallium quod tenebam et fugit foras
GEN|39|16|in argumentum ergo fidei retentum pallium ostendit marito revertenti domum
GEN|39|17|et ait ingressus est ad me servus hebraeus quem adduxisti ut inluderet mihi
GEN|39|18|cumque vidisset me clamare reliquit pallium et fugit foras
GEN|39|19|his auditis dominus et nimium credulus verbis coniugis iratus est valde
GEN|39|20|tradiditque Ioseph in carcerem ubi vincti regis custodiebantur et erat ibi clausus
GEN|39|21|fuit autem Dominus cum Ioseph et misertus illius dedit ei gratiam in conspectu principis carceris
GEN|39|22|qui tradidit in manu ipsius universos vinctos qui in custodia tenebantur et quicquid fiebat sub ipso erat
GEN|39|23|nec noverat aliquid cunctis ei creditis Dominus enim erat cum illo et omnia eius opera dirigebat
GEN|40|1|his ita gestis accidit ut peccarent duo eunuchi pincerna regis Aegypti et pistor domino suo
GEN|40|2|iratusque Pharao contra eos nam alter pincernis praeerat alter pistoribus
GEN|40|3|misit eos in carcerem principis militum in quo erat vinctus et Ioseph
GEN|40|4|at custos carceris tradidit eos Ioseph qui et ministrabat eis aliquantum temporis fluxerat et illi in custodia tenebantur
GEN|40|5|videruntque ambo somnium nocte una iuxta interpretationem congruam sibi
GEN|40|6|ad quos cum introisset Ioseph mane et vidisset eos tristes
GEN|40|7|sciscitatus est dicens cur tristior est hodie solito facies vestra
GEN|40|8|qui responderunt somnium vidimus et non est qui interpretetur nobis dixitque ad eos Ioseph numquid non Dei est interpretatio referte mihi quid videritis
GEN|40|9|narravit prior praepositus pincernarum somnium videbam coram me vitem
GEN|40|10|in qua erant tres propagines crescere paulatim gemmas et post flores uvas maturescere
GEN|40|11|calicemque Pharaonis in manu mea tuli ergo uvas et expressi in calicem quem tenebam et tradidi poculum Pharaoni
GEN|40|12|respondit Ioseph haec est interpretatio somnii tres propagines tres adhuc dies sunt
GEN|40|13|post quos recordabitur Pharao magisterii tui et restituet te in gradum pristinum dabisque ei calicem iuxta officium tuum sicut facere ante consueveras
GEN|40|14|tantum memento mei cum tibi bene fuerit et facies mecum misericordiam ut suggeras Pharaoni et educat me de isto carcere
GEN|40|15|quia furto sublatus sum de terra Hebraeorum et hic innocens in lacum missus sum
GEN|40|16|videns pistorum magister quod prudenter somnium dissolvisset ait et ego vidi somnium quod haberem tria canistra farinae super caput meum
GEN|40|17|et in uno canistro quod erat excelsius portare me omnes cibos qui fiunt arte pistoria avesque comedere ex eo
GEN|40|18|respondit Ioseph haec est interpretatio somnii tria canistra tres adhuc dies sunt
GEN|40|19|post quos auferet Pharao caput tuum ac suspendet te in cruce et lacerabunt volucres carnes tuas
GEN|40|20|exin dies tertius natalicius Pharaonis erat qui faciens grande convivium pueris suis recordatus est inter epulas magistri pincernarum et pistorum principis
GEN|40|21|restituitque alterum in locum suum ut porrigeret regi poculum
GEN|40|22|alterum suspendit in patibulo ut coniectoris veritas probaretur
GEN|40|23|et tamen succedentibus prosperis praepositus pincernarum oblitus est interpretis sui
GEN|41|1|post duos annos vidit Pharao somnium putabat se stare super fluvium
GEN|41|2|de quo ascendebant septem boves pulchrae et crassae nimis et pascebantur in locis palustribus
GEN|41|3|aliae quoque septem emergebant de flumine foedae confectaeque macie et pascebantur in ipsa amnis ripa in locis virentibus
GEN|41|4|devoraveruntque eas quarum mira species et habitudo corporum erat expergefactus Pharao
GEN|41|5|rursum dormivit et vidit alterum somnium septem spicae pullulabant in culmo uno plenae atque formonsae
GEN|41|6|aliae quoque totidem spicae tenues et percussae uredine oriebantur
GEN|41|7|devorantes omnem priorum pulchritudinem evigilans post quietem
GEN|41|8|et facto mane pavore perterritus misit ad coniectores Aegypti cunctosque sapientes et accersitis narravit somnium nec erat qui interpretaretur
GEN|41|9|tunc demum reminiscens pincernarum magister ait confiteor peccatum meum
GEN|41|10|iratus rex servis suis me et magistrum pistorum retrudi iussit in carcerem principis militum
GEN|41|11|ubi una nocte uterque vidimus somnium praesagum futurorum
GEN|41|12|erat ibi puer hebraeus eiusdem ducis militum famulus cui narrantes somnia
GEN|41|13|audivimus quicquid postea rei probavit eventus ego enim redditus sum officio meo et ille suspensus est in cruce
GEN|41|14|protinus ad regis imperium eductum de carcere Ioseph totonderunt ac veste mutata obtulerunt ei
GEN|41|15|cui ille ait vidi somnia nec est qui edisserat quae audivi te prudentissime conicere
GEN|41|16|respondit Ioseph absque me Deus respondebit prospera Pharaoni
GEN|41|17|narravit ergo ille quod viderat putabam me stare super ripam fluminis
GEN|41|18|et septem boves de amne conscendere pulchras nimis et obesis carnibus quae in pastu paludis virecta carpebant
GEN|41|19|et ecce has sequebantur aliae septem boves in tantum deformes et macilentae ut numquam tales in terra Aegypti viderim
GEN|41|20|quae devoratis et consumptis prioribus
GEN|41|21|nullum saturitatis dedere vestigium sed simili macie et squalore torpebant evigilans rursum sopore depressus
GEN|41|22|vidi somnium septem spicae pullulabant in culmo uno plenae atque pulcherrimae
GEN|41|23|aliae quoque septem tenues et percussae uredine oriebantur stipula
GEN|41|24|quae priorum pulchritudinem devorarunt narravi coniectoribus somnium et nemo est qui edisserat
GEN|41|25|respondit Ioseph somnium regis unum est quae facturus est Deus ostendit Pharaoni
GEN|41|26|septem boves pulchrae et septem spicae plenae septem ubertatis anni sunt eandemque vim somnii conprehendunt
GEN|41|27|septem quoque boves tenues atque macilentae quae ascenderunt post eas et septem spicae tenues et vento urente percussae septem anni sunt venturae famis
GEN|41|28|qui hoc ordine conplebuntur
GEN|41|29|ecce septem anni venient fertilitatis magnae in universa terra Aegypti
GEN|41|30|quos sequentur septem anni alii tantae sterilitatis ut oblivioni tradatur cuncta retro abundantia consumptura est enim fames omnem terram
GEN|41|31|et ubertatis magnitudinem perditura inopiae magnitudo
GEN|41|32|quod autem vidisti secundo ad eandem rem pertinens somnium firmitatis indicium est eo quod fiat sermo Dei et velocius impleatur
GEN|41|33|nunc ergo provideat rex virum sapientem et industrium et praeficiat eum terrae Aegypti
GEN|41|34|qui constituat praepositos per singulas regiones et quintam partem fructuum per septem annos fertilitatis
GEN|41|35|qui iam nunc futuri sunt congreget in horrea et omne frumentum sub Pharaonis potestate condatur serveturque in urbibus
GEN|41|36|et paretur futurae septem annorum fami quae pressura est Aegyptum et non consumetur terra inopia
GEN|41|37|placuit Pharaoni consilium et cunctis ministris eius
GEN|41|38|locutusque est ad eos num invenire poterimus talem virum qui spiritu Dei plenus sit
GEN|41|39|dixit ergo ad Ioseph quia ostendit Deus tibi omnia quae locutus es numquid sapientiorem et similem tui invenire potero
GEN|41|40|tu eris super domum meam et ad tui oris imperium cunctus populus oboediet uno tantum regni solio te praecedam
GEN|41|41|dicens quoque rursum Pharao ad Ioseph ecce constitui te super universam terram Aegypti
GEN|41|42|tulit anulum de manu sua et dedit in manu eius vestivitque eum stola byssina et collo torquem auream circumposuit
GEN|41|43|fecitque ascendere super currum suum secundum clamante praecone ut omnes coram eo genuflecterent et praepositum esse scirent universae terrae Aegypti
GEN|41|44|dixit quoque rex ad Ioseph ego sum Pharao absque tuo imperio non movebit quisquam manum aut pedem in omni terra Aegypti
GEN|41|45|vertitque nomen illius et vocavit eum lingua aegyptiaca Salvatorem mundi dedit quoque illi uxorem Aseneth filiam Putiphare sacerdotis Heliopoleos egressus itaque Ioseph ad terram Aegypti
GEN|41|46|triginta autem erat annorum quando stetit in conspectu regis Pharaonis circuivit omnes regiones Aegypti
GEN|41|47|venitque fertilitas septem annorum et in manipulos redactae segetes congregatae sunt in horrea Aegypti
GEN|41|48|omnis etiam frugum abundantia in singulis urbibus condita est
GEN|41|49|tantaque fuit multitudo tritici ut harenae maris coaequaretur et copia mensuram excederet
GEN|41|50|nati sunt autem Ioseph filii duo antequam veniret fames quos ei peperit Aseneth filia Putiphare sacerdotis Heliopoleos
GEN|41|51|vocavitque nomen primogeniti Manasse dicens oblivisci me fecit Deus omnium laborum meorum et domum patris mei
GEN|41|52|nomen quoque secundi appellavit Ephraim dicens crescere me fecit Deus in terra paupertatis meae
GEN|41|53|igitur transactis septem annis ubertatis qui fuerant in Aegypto
GEN|41|54|coeperunt venire septem anni inopiae quos praedixerat Ioseph et in universo orbe fames praevaluit in cuncta autem terra Aegypti erat panis
GEN|41|55|qua esuriente clamavit populus ad Pharaonem alimenta petens quibus ille respondit ite ad Ioseph et quicquid vobis dixerit facite
GEN|41|56|crescebat autem cotidie fames in omni terra aperuitque Ioseph universa horrea et vendebat Aegyptiis nam et illos oppresserat fames
GEN|41|57|omnesque provinciae veniebant in Aegyptum ut emerent escas et malum inopiae temperarent
GEN|42|1|audiens autem Iacob quod alimenta venderentur in Aegypto dixit filiis suis quare neglegitis
GEN|42|2|audivi quod triticum venundetur in Aegypto descendite et emite nobis necessaria ut possimus vivere et non consumamur inopia
GEN|42|3|descendentes igitur fratres Ioseph decem ut emerent frumenta in Aegypto
GEN|42|4|Beniamin domi retento ab Iacob qui dixerat fratribus eius ne forte in itinere quicquam patiatur mali
GEN|42|5|ingressi sunt terram Aegypti cum aliis qui pergebant ad emendum erat autem fames in terra Chanaan
GEN|42|6|et Ioseph princeps Aegypti atque ad illius nutum frumenta populis vendebantur cumque adorassent eum fratres sui
GEN|42|7|et agnovisset eos quasi ad alienos durius loquebatur interrogans eos unde venistis qui responderunt de terra Chanaan ut emamus victui necessaria
GEN|42|8|et tamen fratres ipse cognoscens non est agnitus ab eis
GEN|42|9|recordatusque somniorum quae aliquando viderat ait exploratores estis ut videatis infirmiora terrae venistis
GEN|42|10|qui dixerunt non est ita domine sed servi tui venerunt ut emerent cibos
GEN|42|11|omnes filii unius viri sumus pacifici venimus nec quicquam famuli tui machinantur mali
GEN|42|12|quibus ille respondit aliter est inmunita terrae huius considerare venistis
GEN|42|13|et illi duodecim inquiunt servi tui fratres sumus filii viri unius in terra Chanaan minimus cum patre nostro est alius non est super
GEN|42|14|hoc est ait quod locutus sum exploratores estis
GEN|42|15|iam nunc experimentum vestri capiam per salutem Pharaonis non egrediemini hinc donec veniat frater vester minimus
GEN|42|16|mittite e vobis unum et adducat eum vos autem eritis in vinculis donec probentur quae dixistis utrum falsa an vera sint alioquin per salutem Pharaonis exploratores estis
GEN|42|17|tradidit ergo eos custodiae tribus diebus
GEN|42|18|die autem tertio eductis de carcere ait facite quod dixi et vivetis Deum enim timeo
GEN|42|19|si pacifici estis frater vester unus ligetur in carcere vos autem abite et ferte frumenta quae emistis in domos vestras
GEN|42|20|et fratrem vestrum minimum ad me adducite ut possim vestros probare sermones et non moriamini fecerunt ut dixerat
GEN|42|21|et locuti sunt invicem merito haec patimur quia peccavimus in fratrem nostrum videntes angustiam animae illius cum deprecaretur nos et non audivimus idcirco venit super nos ista tribulatio
GEN|42|22|e quibus unus Ruben ait numquid non dixi vobis nolite peccare in puerum et non audistis me en sanguis eius exquiritur
GEN|42|23|nesciebant autem quod intellegeret Ioseph eo quod per interpretem loquebatur ad eos
GEN|42|24|avertitque se parumper et flevit et reversus locutus est ad eos
GEN|42|25|tollens Symeon et ligans illis praesentibus iussitque ministris ut implerent saccos eorum tritico et reponerent pecunias singulorum in sacculis suis datis supra cibariis in via qui fecerunt ita
GEN|42|26|at illi portantes frumenta in asinis profecti sunt
GEN|42|27|apertoque unus sacco ut daret iumento pabulum in diversorio contemplatus pecuniam in ore sacculi
GEN|42|28|dixit fratribus suis reddita est mihi pecunia en habetur in sacco et obstupefacti turbatique dixerunt mutuo quidnam est hoc quod fecit nobis Deus
GEN|42|29|veneruntque ad Iacob patrem suum in terra Chanaan et narraverunt ei omnia quae accidissent sibi dicentes
GEN|42|30|locutus est nobis dominus terrae dure et putavit nos exploratores provinciae
GEN|42|31|cui respondimus pacifici sumus nec ullas molimur insidias
GEN|42|32|duodecim fratres uno patre geniti sumus unus non est super minimus cum patre versatur in terra Chanaan
GEN|42|33|qui ait nobis sic probabo quod pacifici sitis fratrem vestrum unum dimittite apud me et cibaria domibus vestris necessaria sumite et abite
GEN|42|34|fratremque vestrum minimum adducite ad me ut sciam quod non sitis exploratores et istum qui tenetur in vinculis recipere possitis ac deinceps emendi quae vultis habeatis licentiam
GEN|42|35|his dictis cum frumenta effunderent singuli reppererunt in ore saccorum ligatas pecunias exterritisque simul omnibus
GEN|42|36|dixit pater Iacob absque liberis me esse fecistis Ioseph non est super Symeon tenetur in vinculis Beniamin auferetis in me haec mala omnia reciderunt
GEN|42|37|cui respondit Ruben duos filios meos interfice si non reduxero illum tibi trade in manu mea et ego eum restituam
GEN|42|38|at ille non descendet inquit filius meus vobiscum frater eius mortuus est ipse solus remansit si quid ei adversi acciderit in terra ad quam pergitis deducetis canos meos cum dolore ad inferos
GEN|43|1|interim fames omnem terram vehementer premebat
GEN|43|2|consumptisque cibis quos ex Aegypto detulerant dixit Iacob ad filios suos revertimini et emite pauxillum escarum
GEN|43|3|respondit Iudas denuntiavit nobis vir ille sub testificatione iurandi dicens non videbitis faciem meam nisi fratrem vestrum minimum adduxeritis vobiscum
GEN|43|4|si ergo vis mittere eum nobiscum pergemus pariter et ememus tibi necessaria
GEN|43|5|si autem non vis non ibimus vir enim ut saepe diximus denuntiavit nobis dicens non videbitis faciem meam absque fratre vestro minimo
GEN|43|6|dixit eis Israhel in meam hoc fecistis miseriam ut indicaretis ei et alium habere vos fratrem
GEN|43|7|at illi responderunt interrogavit nos homo per ordinem nostram progeniem si pater viveret si haberemus fratrem et nos respondimus ei consequenter iuxta id quod fuerat sciscitatus numquid scire poteramus quod dicturus esset adducite vobiscum fratrem vestrum
GEN|43|8|Iudas quoque dixit patri suo mitte puerum mecum ut proficiscamur et possimus vivere ne moriamur nos et parvuli nostri
GEN|43|9|ego suscipio puerum de manu mea require illum nisi reduxero et tradidero eum tibi ero peccati in te reus omni tempore
GEN|43|10|si non intercessisset dilatio iam vice altera venissemus
GEN|43|11|igitur Israhel pater eorum dixit ad eos si sic necesse est facite quod vultis sumite de optimis terrae fructibus in vasis vestris et deferte viro munera modicum resinae et mellis et styracis et stactes et terebinthi et amigdalarum
GEN|43|12|pecuniamque duplicem ferte vobiscum et illam quam invenistis in sacculis reportate ne forte errore factum sit
GEN|43|13|sed et fratrem vestrum tollite et ite ad virum
GEN|43|14|Deus autem meus omnipotens faciat vobis eum placabilem et remittat vobiscum fratrem vestrum quem tenet et hunc Beniamin ego autem quasi orbatus absque liberis ero
GEN|43|15|tulerunt ergo viri munera et pecuniam duplicem et Beniamin descenderuntque in Aegyptum et steterunt coram Ioseph
GEN|43|16|quos cum ille vidisset et Beniamin simul praecepit dispensatori domus suae dicens introduc viros domum et occide victimas et instrue convivium quoniam mecum sunt comesuri meridie
GEN|43|17|fecit ille sicut fuerat imperatum et introduxit viros domum
GEN|43|18|ibique exterriti dixerunt mutuo propter pecuniam quam rettulimus prius in saccis nostris introducti sumus ut devolvat in nos calumniam et violenter subiciat servituti et nos et asinos nostros
GEN|43|19|quam ob rem in ipsis foribus accedentes ad dispensatorem
GEN|43|20|locuti sunt oramus domine ut audias iam ante descendimus ut emeremus escas
GEN|43|21|quibus emptis cum venissemus ad diversorium aperuimus sacculos nostros et invenimus pecuniam in ore saccorum quam nunc eodem pondere reportamus
GEN|43|22|sed et aliud adtulimus argentum ut emamus quae necessaria sunt non est in nostra conscientia quis eam posuerit in marsuppiis nostris
GEN|43|23|at ille respondit pax vobiscum nolite timere Deus vester et Deus patris vestri dedit vobis thesauros in sacculis vestris nam pecuniam quam dedistis mihi probatam ego habeo eduxitque ad eos Symeon
GEN|43|24|et introductis domum adtulit aquam et laverunt pedes suos deditque pabula asinis eorum
GEN|43|25|illi vero parabant munera donec ingrederetur Ioseph meridie audierant enim quod ibi comesuri essent panem
GEN|43|26|igitur ingressus est Ioseph domum suam obtuleruntque ei munera tenentes in manibus et adoraverunt proni in terram
GEN|43|27|at ille clementer resalutatis eis interrogavit dicens salvusne est pater vester senex de quo dixeratis mihi adhuc vivit
GEN|43|28|qui responderunt sospes est servus tuus pater noster adhuc vivit et incurvati adoraverunt eum
GEN|43|29|adtollens autem oculos Ioseph vidit Beniamin fratrem suum uterinum et ait iste est frater vester parvulus de quo dixeratis mihi et rursum Deus inquit misereatur tui fili mi
GEN|43|30|festinavitque quia commota fuerant viscera eius super fratre suo et erumpebant lacrimae et introiens cubiculum flevit
GEN|43|31|rursusque lota facie egressus continuit se et ait ponite panes
GEN|43|32|quibus adpositis seorsum Ioseph et seorsum fratribus Aegyptiis quoque qui vescebantur simul seorsum inlicitum est enim Aegyptiis comedere cum Hebraeis et profanum putant huiuscemodi convivium
GEN|43|33|sederunt coram eo primogenitus iuxta primogenita sua et minimus iuxta aetatem suam et mirabantur nimis
GEN|43|34|sumptis partibus quas ab eo acceperant maiorque pars venit Beniamin ita ut quinque partibus excederet biberuntque et inebriati sunt cum eo
GEN|44|1|praecepit autem Ioseph dispensatori domus suae dicens imple saccos eorum frumento quantum possunt capere et pone pecuniam singulorum in summitate sacci
GEN|44|2|scyphum autem meum argenteum et pretium quod dedit tritici pone in ore sacci iunioris factumque est ita
GEN|44|3|et orto mane dimissi sunt cum asinis suis
GEN|44|4|iamque urbem exierant et processerant paululum tum Ioseph arcessito dispensatore domus surge inquit persequere viros et adprehensis dicito quare reddidistis malum pro bono
GEN|44|5|scyphum quem furati estis ipse est in quo bibit dominus meus et in quo augurari solet pessimam rem fecistis
GEN|44|6|fecit ille ut iusserat et adprehensis per ordinem locutus est
GEN|44|7|qui responderunt quare sic loquitur dominus noster ut servi tui tantum flagitii commiserint
GEN|44|8|pecuniam quam invenimus in summitate saccorum reportavimus ad te de terra Chanaan et quomodo consequens est ut furati simus de domo domini tui aurum vel argentum
GEN|44|9|apud quemcumque fuerit inventum servorum tuorum quod quaeris moriatur et nos servi erimus domini nostri
GEN|44|10|qui dixit fiat iuxta vestram sententiam apud quem fuerit inventum ipse sit servus meus vos autem eritis innoxii
GEN|44|11|itaque festinato deponentes in terram saccos aperuerunt singuli
GEN|44|12|quos scrutatus incipiens a maiore usque ad minimum invenit scyphum in sacco Beniamin
GEN|44|13|at illi scissis vestibus oneratisque rursum asinis reversi sunt in oppidum
GEN|44|14|primusque Iudas cum fratribus ingressus est ad Ioseph necdum enim de loco abierat omnesque ante eum in terra pariter corruerunt
GEN|44|15|quibus ille ait cur sic agere voluistis an ignoratis quod non sit similis mei in augurandi scientia
GEN|44|16|cui Iudas quid respondebimus inquit domino meo vel quid loquemur aut iusti poterimus obtendere Deus invenit iniquitatem servorum tuorum en omnes servi sumus domini mei et nos et apud quem inventus est scyphus
GEN|44|17|respondit Ioseph absit a me ut sic agam qui furatus est scyphum ipse sit servus meus vos autem abite liberi ad patrem vestrum
GEN|44|18|accedens propius Iudas confidenter ait oro domine mi loquatur servus tuus verbum in auribus tuis et ne irascaris famulo tuo tu es enim post Pharaonem
GEN|44|19|dominus meus interrogasti prius servos tuos habetis patrem aut fratrem
GEN|44|20|et nos respondimus tibi domino meo est nobis pater senex et puer parvulus qui in senecta illius natus est cuius uterinus frater est mortuus et ipsum solum habet mater sua pater vero tenere diligit eum
GEN|44|21|dixistique servis tuis adducite eum ad me et ponam oculos meos super illum
GEN|44|22|suggessimus domino meo non potest puer relinquere patrem suum si enim illum dimiserit morietur
GEN|44|23|et dixisti servis tuis nisi venerit frater vester minimus vobiscum non videbitis amplius faciem meam
GEN|44|24|cum ergo ascendissemus ad famulum tuum patrem nostrum narravimus ei omnia quae locutus est dominus meus
GEN|44|25|et dixit pater noster revertimini et emite nobis parum tritici
GEN|44|26|cui diximus ire non possumus si frater noster minimus descendet nobiscum proficiscemur simul alioquin illo absente non audemus videre faciem viri
GEN|44|27|atque ille respondit vos scitis quod duos genuerit mihi uxor mea
GEN|44|28|egressus est unus et dixistis bestia devoravit eum et hucusque non conparet
GEN|44|29|si tuleritis et istum et aliquid ei in via contigerit deducetis canos meos cum maerore ad inferos
GEN|44|30|igitur si intravero ad servum tuum patrem nostrum et puer defuerit cum anima illius ex huius anima pendeat
GEN|44|31|videritque eum non esse nobiscum morietur et deducent famuli tui canos eius cum dolore ad inferos
GEN|44|32|ego proprie servus tuus qui in meam hunc recepi fidem et spopondi dicens nisi reduxero eum peccati reus ero in patrem meum omni tempore
GEN|44|33|manebo itaque servus tuus pro puero in ministerium domini mei et puer ascendat cum fratribus suis
GEN|44|34|non enim possum redire ad patrem absente puero ne calamitatis quae oppressura est patrem meum testis adsistam
GEN|45|1|non se poterat ultra cohibere Ioseph multis coram adstantibus unde praecepit ut egrederentur cuncti foras et nullus interesset alienus agnitioni mutuae
GEN|45|2|elevavitque vocem cum fletu quam audierunt Aegyptii omnisque domus Pharaonis
GEN|45|3|et dixit fratribus suis ego sum Ioseph adhuc pater meus vivit nec poterant respondere fratres nimio timore perterriti
GEN|45|4|ad quos ille clementer accedite inquit ad me et cum accessissent prope ego sum ait Ioseph frater vester quem vendidistis in Aegypto
GEN|45|5|nolite pavere nec vobis durum esse videatur quod vendidistis me in his regionibus pro salute enim vestra misit me Deus ante vos in Aegyptum
GEN|45|6|biennium est quod fames esse coepit in terra et adhuc quinque anni restant quibus nec arari poterit nec meti
GEN|45|7|praemisitque me Deus ut reservemini super terram et escas ad vivendum habere possitis
GEN|45|8|non vestro consilio sed Dei huc voluntate missus sum qui fecit me quasi patrem Pharaonis et dominum universae domus eius ac principem in omni terra Aegypti
GEN|45|9|festinate et ascendite ad patrem meum et dicetis ei haec mandat filius tuus Ioseph Deus me fecit dominum universae terrae Aegypti descende ad me ne moreris
GEN|45|10|et habita in terra Gessen erisque iuxta me tu et filii tui et filii filiorum tuorum oves tuae et armenta tua et universa quae possides
GEN|45|11|ibique te pascam adhuc enim quinque anni residui sunt famis ne et tu pereas et domus tua et omnia quae possides
GEN|45|12|en oculi vestri et oculi fratris mei Beniamin vident quod os meum loquatur ad vos
GEN|45|13|nuntiate patri meo universam gloriam meam et cuncta quae vidistis in Aegypto festinate et adducite eum ad me
GEN|45|14|cumque amplexatus recidisset in collum Beniamin fratris sui flevit illo quoque flente similiter super collum eius
GEN|45|15|osculatusque est Ioseph omnes fratres suos et ploravit super singulos post quae ausi sunt loqui ad eum
GEN|45|16|auditumque est et celebri sermone vulgatum in aula regis venerunt fratres Ioseph et gavisus est Pharao atque omnis familia eius
GEN|45|17|dixitque ad Ioseph ut imperaret fratribus suis dicens onerantes iumenta ite in terram Chanaan
GEN|45|18|et tollite inde patrem vestrum et cognationem et venite ad me et ego dabo vobis omnia bona Aegypti ut comedatis medullam terrae
GEN|45|19|praecipe etiam ut tollant plaustra de terra Aegypti ad subvectionem parvulorum suorum et coniugum ac dicito tollite patrem vestrum et properate quantocius venientes
GEN|45|20|ne dimittatis quicquam de supellectili vestra quia omnes opes Aegypti vestrae erunt
GEN|45|21|fecerunt filii Israhel ut eis mandatum fuerat quibus dedit Ioseph plaustra secundum Pharaonis imperium et cibaria in itinere
GEN|45|22|singulisque proferri iussit binas stolas Beniamin vero dedit trecentos argenteos cum quinque stolis optimis
GEN|45|23|tantundem pecuniae et vestium mittens patri suo addens eis asinos decem qui subveherent ex omnibus divitiis Aegypti et totidem asinas triticum in itinere panesque portantes
GEN|45|24|dimisit ergo fratres suos et proficiscentibus ait ne irascamini in via
GEN|45|25|qui ascendentes ex Aegypto venerunt in terram Chanaan ad patrem suum Iacob
GEN|45|26|et nuntiaverunt ei dicentes Ioseph vivit et ipse dominatur in omni terra Aegypti quo audito quasi de gravi somno evigilans tamen non credebat eis
GEN|45|27|illi contra referebant omnem ordinem rei cumque vidisset plaustra et universa quae miserat revixit spiritus eius
GEN|45|28|et ait sufficit mihi si adhuc Ioseph filius meus vivit vadam et videbo illum antequam moriar
GEN|46|1|profectusque Israhel cum omnibus quae habebat venit ad puteum Iuramenti et mactatis ibi victimis Deo patris sui Isaac
GEN|46|2|audivit eum per visionem nocte vocantem se et dicentem sibi Iacob Iacob cui respondit ecce adsum
GEN|46|3|ait illi Deus ego sum Fortissimus Deus patris tui noli timere et descende in Aegyptum quia in gentem magnam faciam te ibi
GEN|46|4|ego descendam tecum illuc et ego inde adducam te revertentem Ioseph quoque ponet manum suam super oculos tuos
GEN|46|5|surrexit Iacob a puteo Iuramenti tuleruntque eum filii cum parvulis et uxoribus suis in plaustris quae miserat Pharao ad portandum senem
GEN|46|6|et omnia quae possederat in terra Chanaan venitque in Aegyptum cum omni semine suo
GEN|46|7|filii eius et nepotes filiae et cuncta simul progenies
GEN|46|8|haec sunt autem nomina filiorum Israhel qui ingressi sunt in Aegyptum ipse cum liberis suis primogenitus Ruben
GEN|46|9|filii Ruben Enoch et Phallu et Esrom et Charmi
GEN|46|10|filii Symeon Iemuhel et Iamin et Ahod et Iachin et Saher et Saul filius Chananitidis
GEN|46|11|filii Levi Gerson Caath et Merari
GEN|46|12|filii Iuda Her et Onan et Sela et Phares et Zara mortui sunt autem Her et Onan in terra Chanaan natique sunt filii Phares Esrom et Amul
GEN|46|13|filii Isachar Thola et Phua et Iob et Semron
GEN|46|14|filii Zabulon Sared et Helon et Iahelel
GEN|46|15|hii filii Liae quos genuit in Mesopotamiam Syriae cum Dina filia sua omnes animae filiorum eius et filiarum triginta tres
GEN|46|16|filii Gad Sephion et Haggi Suni et Esebon Heri et Arodi et Areli
GEN|46|17|filii Aser Iamne et Iesua et Iesui et Beria Sara quoque soror eorum filii Beria Heber et Melchihel
GEN|46|18|hii filii Zelphae quam dedit Laban Liae filiae suae et hos genuit Iacob sedecim animas
GEN|46|19|filii Rahel uxoris Iacob Ioseph et Beniamin
GEN|46|20|natique sunt Ioseph filii in terra Aegypti quos genuit ei Aseneth filia Putiphare sacerdotis Heliopoleos Manasses et Ephraim
GEN|46|21|filii Beniamin Bela et Bechor et Asbel Gera et Naaman et Ehi et Ros Mophim et Opphim et Ared
GEN|46|22|hii filii Rahel quos genuit Iacob omnes animae quattuordecim
GEN|46|23|filii Dan Usim
GEN|46|24|filii Nepthalim Iasihel et Guni et Hieser et Sallem
GEN|46|25|hii filii Balae quam dedit Laban Raheli filiae suae et hos genuit Iacob omnes animae septem
GEN|46|26|cunctae animae quae ingressae sunt cum Iacob in Aegyptum et egressae de femore illius absque uxoribus filiorum sexaginta sex
GEN|46|27|filii autem Ioseph qui nati sunt ei in terra Aegypti animae duae omnis anima domus Iacob quae ingressa est Aegyptum fuere septuaginta
GEN|46|28|misit autem Iudam ante se ad Ioseph ut nuntiaret ei et ille occurreret in Gessen
GEN|46|29|quo cum pervenisset iuncto Ioseph curru suo ascendit obviam patri ad eundem locum vidensque eum inruit super collum eius et inter amplexus flevit
GEN|46|30|dixitque pater ad Ioseph iam laetus moriar quia vidi faciem tuam et superstitem te relinquo
GEN|46|31|et ille locutus est ad fratres et ad omnem domum patris sui ascendam et nuntiabo Pharaoni dicamque ei fratres mei et domus patris mei qui erant in terra Chanaan venerunt ad me
GEN|46|32|et sunt viri pastores ovium curamque habent alendorum gregum pecora sua et armenta et omnia quae habere potuerunt adduxerunt secum
GEN|46|33|cumque vocaverit vos et dixerit quod est opus vestrum
GEN|46|34|respondebitis viri pastores sumus servi tui ab infantia nostra usque in praesens et nos et patres nostri haec autem dicetis ut habitare possitis in terra Gessen quia detestantur Aegyptii omnes pastores ovium
GEN|47|1|ingressus ergo Ioseph nuntiavit Pharaoni dicens pater meus et fratres oves eorum et armenta et cuncta quae possident venerunt de terra Chanaan et ecce consistunt in terra Gessen
GEN|47|2|extremos quoque fratrum suorum quinque viros statuit coram rege
GEN|47|3|quos ille interrogavit quid habetis operis responderunt pastores ovium sumus servi tui et nos et patres nostri
GEN|47|4|ad peregrinandum in terra tua venimus quoniam non est herba gregibus servorum tuorum ingravescente fame in regione Chanaan petimusque ut esse nos iubeas servos tuos in terra Gessen
GEN|47|5|dixit itaque rex ad Ioseph pater tuus et fratres tui venerunt ad te
GEN|47|6|terra Aegypti in conspectu tuo est in optimo loco fac habitare eos et trade eis terram Gessen quod si nosti esse in eis viros industrios constitue illos magistros pecorum meorum
GEN|47|7|post haec introduxit Ioseph patrem suum ad regem et statuit eum coram eo qui benedicens illi
GEN|47|8|et interrogatus ab eo quot sunt dies annorum vitae tuae
GEN|47|9|respondit dies peregrinationis vitae meae centum triginta annorum sunt parvi et mali et non pervenerunt usque ad dies patrum meorum quibus peregrinati sunt
GEN|47|10|et benedicto rege egressus est foras
GEN|47|11|Ioseph vero patri et fratribus suis dedit possessionem in Aegypto in optimo loco terrae solo Ramesses ut praeceperat Pharao
GEN|47|12|et alebat eos omnemque domum patris sui praebens cibaria singulis
GEN|47|13|in toto enim orbe panis deerat et oppresserat fames terram maxime Aegypti et Chanaan
GEN|47|14|e quibus omnem pecuniam congregavit pro venditione frumenti et intulit eam in aerarium regis
GEN|47|15|cumque defecisset emptoris pretium venit cuncta Aegyptus ad Ioseph dicens da nobis panes quare morimur coram te deficiente pecunia
GEN|47|16|quibus ille respondit adducite pecora vestra et dabo vobis pro eis cibos si pretium non habetis
GEN|47|17|quae cum adduxissent dedit eis alimenta pro equis et ovibus et bubus et asinis sustentavitque eos illo anno pro commutatione pecorum
GEN|47|18|veneruntque anno secundo et dixerunt ei non celamus dominum nostrum quod deficiente pecunia pecora simul defecerint nec clam te est quod absque corporibus et terra nihil habeamus
GEN|47|19|cur ergo morimur te vidente et nos et terra nostra tui erimus eme nos in servitutem regiam et praebe semina ne pereunte cultore redigatur terra in solitudinem
GEN|47|20|emit igitur Ioseph omnem terram Aegypti vendentibus singulis possessiones suas prae magnitudine famis subiecitque eam Pharaoni
GEN|47|21|et cunctos populos eius a novissimis terminis Aegypti usque ad extremos fines eius
GEN|47|22|praeter terram sacerdotum quae a rege tradita fuerat eis quibus et statuta cibaria ex horreis publicis praebebantur et idcirco non sunt conpulsi vendere possessiones suas
GEN|47|23|dixit ergo Ioseph ad populos en ut cernitis et vos et terram vestram Pharao possidet accipite semina et serite agros
GEN|47|24|ut fruges habere possitis quintam partem regi dabitis quattuor reliquas permitto vobis in sementem et in cibos famulis et liberis vestris
GEN|47|25|qui responderunt salus nostra in manu tua est respiciat nos tantum dominus noster et laeti serviemus regi
GEN|47|26|ex eo tempore usque in praesentem diem in universa terra Aegypti regibus quinta pars solvitur et factum est quasi in legem absque terra sacerdotali quae libera ab hac condicione fuit
GEN|47|27|habitavit ergo Israhel in Aegypto id est in terra Gessen et possedit eam auctusque est et multiplicatus nimis
GEN|47|28|et vixit in ea decem et septem annis factique sunt omnes dies vitae illius centum quadraginta septem annorum
GEN|47|29|cumque adpropinquare cerneret mortis diem vocavit filium suum Ioseph et dixit ad eum si inveni gratiam in conspectu tuo pone manum sub femore meo et facies mihi misericordiam et veritatem ut non sepelias me in Aegypto
GEN|47|30|sed dormiam cum patribus meis et auferas me de hac terra condasque in sepulchro maiorum cui respondit Ioseph ego faciam quod iussisti
GEN|47|31|et ille iura ergo inquit mihi quo iurante adoravit Israhel Deum conversus ad lectuli caput
GEN|48|1|his ita transactis nuntiatum est Ioseph quod aegrotaret pater eius qui adsumptis duobus filiis Manasse et Ephraim ire perrexit
GEN|48|2|dictumque est seni ecce filius tuus Ioseph venit ad te qui confortatus sedit in lectulo
GEN|48|3|et ingresso ad se ait Deus omnipotens apparuit mihi in Luza quae est in terra Chanaan benedixitque mihi
GEN|48|4|et ait ego te augebo et multiplicabo et faciam in turbas populorum daboque tibi terram hanc et semini tuo post te in possessionem sempiternam
GEN|48|5|duo igitur filii tui qui nati sunt tibi in terra Aegypti antequam huc venirem ad te mei erunt Ephraim et Manasses sicut Ruben et Symeon reputabuntur mihi
GEN|48|6|reliquos autem quos genueris post eos tui erunt et nomine fratrum suorum vocabuntur in possessionibus suis
GEN|48|7|mihi enim quando veniebam de Mesopotamiam mortua est Rahel in terra Chanaan in ipso itinere eratque vernum tempus et ingrediebar Ephratam et sepelivi eam iuxta viam Ephratae quae alio nomine appellatur Bethleem
GEN|48|8|videns autem filios eius dixit ad eum qui sunt isti
GEN|48|9|respondit filii mei sunt quos dedit mihi Deus in hoc loco adduc inquit eos ad me ut benedicam illis
GEN|48|10|oculi enim Israhel caligabant prae nimia senectute et clare videre non poterat adplicitosque ad se deosculatus et circumplexus
GEN|48|11|dixit ad filium non sum fraudatus aspectu tuo insuper ostendit mihi Deus semen tuum
GEN|48|12|cumque tulisset eos Ioseph de gremio patris adoravit pronus in terram
GEN|48|13|et posuit Ephraim ad dexteram suam id est ad sinistram Israhel Manassen vero in sinistra sua ad dexteram scilicet patris adplicuitque ambos ad eum
GEN|48|14|qui extendens manum dextram posuit super caput Ephraim iunioris fratris sinistram autem super caput Manasse qui maior natu erat commutans manus
GEN|48|15|benedixitque Ioseph filio suo et ait Deus in cuius conspectu ambulaverunt patres mei Abraham et Isaac Deus qui pascit me ab adulescentia mea usque in praesentem diem
GEN|48|16|angelus qui eruit me de cunctis malis benedicat pueris et invocetur super eos nomen meum nomina quoque patrum meorum Abraham et Isaac et crescant in multitudinem super terram
GEN|48|17|videns autem Ioseph quod posuisset pater suus dexteram manum super caput Ephraim graviter accepit et adprehensam patris manum levare conatus est de capite Ephraim et transferre super caput Manasse
GEN|48|18|dixitque ad patrem non ita convenit pater quia hic est primogenitus pone dexteram tuam super caput eius
GEN|48|19|qui rennuens ait scio fili mi scio et iste quidem erit in populos et multiplicabitur sed frater eius iunior maior illo erit et semen illius crescet in gentes
GEN|48|20|benedixitque eis in ipso tempore dicens in te benedicetur Israhel atque dicetur faciat tibi Deus sicut Ephraim et sicut Manasse constituitque Ephraim ante Manassen
GEN|48|21|et ait ad Ioseph filium suum en ego morior et erit Deus vobiscum reducetque vos ad terram patrum vestrorum
GEN|48|22|do tibi partem unam extra fratres tuos quam tuli de manu Amorrei in gladio et arcu meo
GEN|49|1|vocavit autem Iacob filios suos et ait eis congregamini ut adnuntiem quae ventura sunt vobis diebus novissimis
GEN|49|2|congregamini et audite filii Iacob audite Israhel patrem vestrum
GEN|49|3|Ruben primogenitus meus tu fortitudo mea et principium doloris mei prior in donis maior imperio
GEN|49|4|effusus es sicut aqua non crescas quia ascendisti cubile patris tui et maculasti stratum eius
GEN|49|5|Symeon et Levi fratres vasa iniquitatis bellantia
GEN|49|6|in consilio eorum ne veniat anima mea et in coetu illorum non sit gloria mea quia in furore suo occiderunt virum et in voluntate sua suffoderunt murum
GEN|49|7|maledictus furor eorum quia pertinax et indignatio illorum quia dura dividam eos in Iacob et dispergam illos in Israhel
GEN|49|8|Iuda te laudabunt fratres tui manus tua in cervicibus inimicorum tuorum adorabunt te filii patris tui
GEN|49|9|catulus leonis Iuda a praeda fili mi ascendisti requiescens accubuisti ut leo et quasi leaena quis suscitabit eum
GEN|49|10|non auferetur sceptrum de Iuda et dux de femoribus eius donec veniat qui mittendus est et ipse erit expectatio gentium
GEN|49|11|ligans ad vineam pullum suum et ad vitem o fili mi asinam suam lavabit vino stolam suam et sanguine uvae pallium suum
GEN|49|12|pulchriores oculi eius vino et dentes lacte candidiores
GEN|49|13|Zabulon in litore maris habitabit et in statione navium pertingens usque ad Sidonem
GEN|49|14|Isachar asinus fortis accubans inter terminos
GEN|49|15|vidit requiem quod esset bona et terram quod optima et subposuit umerum suum ad portandum factusque est tributis serviens
GEN|49|16|Dan iudicabit populum suum sicut et alia tribus Israhel
GEN|49|17|fiat Dan coluber in via cerastes in semita mordens ungulas equi ut cadat ascensor eius retro
GEN|49|18|salutare tuum expectabo Domine
GEN|49|19|Gad accinctus proeliabitur ante eum et ipse accingetur retrorsum
GEN|49|20|Aser pinguis panis eius et praebebit delicias regibus
GEN|49|21|Nepthalim cervus emissus et dans eloquia pulchritudinis
GEN|49|22|filius adcrescens Ioseph filius adcrescens et decorus aspectu filiae discurrerunt super murum
GEN|49|23|sed exasperaverunt eum et iurgati sunt invideruntque illi habentes iacula
GEN|49|24|sedit in forti arcus eius et dissoluta sunt vincula brachiorum et manuum illius per manus potentis Iacob inde pastor egressus est lapis Israhel
GEN|49|25|Deus patris tui erit adiutor tuus et Omnipotens benedicet tibi benedictionibus caeli desuper benedictionibus abyssi iacentis deorsum benedictionibus uberum et vulvae
GEN|49|26|benedictiones patris tui confortatae sunt benedictionibus patrum eius donec veniret desiderium collium aeternorum fiant in capite Ioseph et in vertice nazarei inter fratres suos
GEN|49|27|Beniamin lupus rapax mane comedet praedam et vespere dividet spolia
GEN|49|28|omnes hii in tribubus Israhel duodecim haec locutus est eis pater suus benedixitque singulis benedictionibus propriis
GEN|49|29|et praecepit eis dicens ego congregor ad populum meum sepelite me cum patribus meis in spelunca duplici quae est in agro Ephron Hetthei
GEN|49|30|contra Mambre in terra Chanaan quam emit Abraham cum agro ab Ephron Hettheo in possessionem sepulchri
GEN|49|31|ibi sepelierunt eum et Sarram uxorem eius ibi sepultus est Isaac cum Rebecca coniuge ibi et Lia condita iacet
GEN|49|32|finitisque mandatis quibus filios instruebat collegit pedes suos super lectulum et obiit adpositusque est ad populum suum
GEN|49|33|
GEN|50|1|quod cernens Ioseph ruit super faciem patris flens et deosculans eum
GEN|50|2|praecepitque servis suis medicis ut aromatibus condirent patrem
GEN|50|3|quibus iussa explentibus transierunt quadraginta dies iste quippe mos erat cadaverum conditorum flevitque eum Aegyptus septuaginta diebus
GEN|50|4|et expleto planctus tempore locutus est Ioseph ad familiam Pharaonis si inveni gratiam in conspectu vestro loquimini in auribus Pharaonis
GEN|50|5|eo quod pater meus adiuraverit me dicens en morior in sepulchro meo quod fodi mihi in terra Chanaan sepelies me ascendam igitur et sepeliam patrem meum ac revertar
GEN|50|6|dixitque ei Pharao ascende et sepeli patrem tuum sicut adiuratus es
GEN|50|7|quo ascendente ierunt cum eo omnes senes domus Pharaonis cunctique maiores natu terrae Aegypti
GEN|50|8|domus Ioseph cum fratribus suis absque parvulis et gregibus atque armentis quae dereliquerant in terra Gessen
GEN|50|9|habuit quoque in comitatu currus et equites et facta est turba non modica
GEN|50|10|veneruntque ad aream Atad quae sita est trans Iordanem ubi celebrantes exequias planctu magno atque vehementi impleverunt septem dies
GEN|50|11|quod cum vidissent habitatores terrae Chanaan dixerunt planctus magnus est iste Aegyptiis et idcirco appellaverunt nomen loci illius Planctus Aegypti
GEN|50|12|fecerunt ergo filii Iacob sicut praeceperat eis
GEN|50|13|et portantes eum in terram Chanaan sepelierunt in spelunca duplici quam emerat Abraham cum agro in possessionem sepulchri ab Ephron Hettheo contra faciem Mambre
GEN|50|14|reversusque est Ioseph in Aegyptum cum fratribus suis et omni comitatu sepulto patre
GEN|50|15|quo mortuo timentes fratres eius et mutuo conloquentes ne forte memor sit iniuriae quam passus est et reddat nobis malum omne quod fecimus
GEN|50|16|mandaverunt ei pater tuus praecepit nobis antequam moreretur
GEN|50|17|ut haec tibi verbis illius diceremus obsecro ut obliviscaris sceleris fratrum tuorum et peccati atque malitiae quam exercuerunt in te nos quoque oramus ut servis Dei patris tui dimittas iniquitatem hanc quibus auditis flevit Ioseph
GEN|50|18|veneruntque ad eum fratres sui et proni in terram dixerunt servi tui sumus
GEN|50|19|quibus ille respondit nolite timere num Dei possumus rennuere voluntatem
GEN|50|20|vos cogitastis de me malum et Deus vertit illud in bonum ut exaltaret me sicut inpraesentiarum cernitis et salvos faceret multos populos
GEN|50|21|nolite metuere ego pascam vos et parvulos vestros consolatusque est eos et blande ac leniter est locutus
GEN|50|22|et habitavit in Aegypto cum omni domo patris sui vixitque centum decem annis et vidit Ephraim filios usque ad tertiam generationem filii quoque Machir filii Manasse nati sunt in genibus Ioseph
GEN|50|23|quibus transactis locutus est fratribus suis post mortem meam Deus visitabit vos et ascendere faciet de terra ista ad terram quam iuravit Abraham Isaac et Iacob
GEN|50|24|cumque adiurasset eos atque dixisset Deus visitabit vos asportate vobiscum ossa mea de loco isto
GEN|50|25|mortuus est expletis centum decem vitae suae annis et conditus aromatibus repositus est in loculo in Aegypto
GEN|50|26|
EXOD|1|1|haec sunt nomina filiorum Israhel qui ingressi sunt Aegyptum cum Iacob singuli cum domibus suis introierunt
EXOD|1|2|Ruben Symeon Levi Iuda
EXOD|1|3|Isachar Zabulon et Beniamin
EXOD|1|4|Dan et Nepthalim Gad et Aser
EXOD|1|5|erant igitur omnes animae eorum qui egressi sunt de femore Iacob septuaginta Ioseph autem in Aegypto erat
EXOD|1|6|quo mortuo et universis fratribus eius omnique cognatione illa
EXOD|1|7|filii Israhel creverunt et quasi germinantes multiplicati sunt ac roborati nimis impleverunt terram
EXOD|1|8|surrexit interea rex novus super Aegyptum qui ignorabat Ioseph
EXOD|1|9|et ait ad populum suum ecce populus filiorum Israhel multus et fortior nobis
EXOD|1|10|venite sapienter opprimamus eum ne forte multiplicetur et si ingruerit contra nos bellum addatur inimicis nostris expugnatisque nobis egrediatur e terra
EXOD|1|11|praeposuit itaque eis magistros operum ut adfligerent eos oneribus aedificaveruntque urbes tabernaculorum Pharaoni Phiton et Ramesses
EXOD|1|12|quantoque opprimebant eos tanto magis multiplicabantur et crescebant
EXOD|1|13|oderantque filios Israhel Aegyptii et adfligebant inludentes eis
EXOD|1|14|atque ad amaritudinem perducebant vitam eorum operibus duris luti et lateris omnique famulatu quo in terrae operibus premebantur
EXOD|1|15|dixit autem rex Aegypti obsetricibus Hebraeorum quarum una vocabatur Sephra altera Phua
EXOD|1|16|praecipiens eis quando obsetricabitis Hebraeas et partus tempus advenerit si masculus fuerit interficite illum si femina reservate
EXOD|1|17|timuerunt autem obsetrices Deum et non fecerunt iuxta praeceptum regis Aegypti sed conservabant mares
EXOD|1|18|quibus ad se accersitis rex ait quidnam est hoc quod facere voluistis ut pueros servaretis
EXOD|1|19|quae responderunt non sunt hebraeae sicut aegyptiae mulieres ipsae enim obsetricandi habent scientiam et priusquam veniamus ad eas pariunt
EXOD|1|20|bene ergo fecit Deus obsetricibus et crevit populus confortatusque est nimis
EXOD|1|21|et quia timuerant obsetrices Deum aedificavit illis domos
EXOD|1|22|praecepit autem Pharao omni populo suo dicens quicquid masculini sexus natum fuerit in flumen proicite quicquid feminei reservate
EXOD|2|1|egressus est post haec vir de domo Levi accepta uxore stirpis suae
EXOD|2|2|quae concepit et peperit filium et videns eum elegantem abscondit tribus mensibus
EXOD|2|3|cumque iam celare non posset sumpsit fiscellam scirpeam et linivit eam bitumine ac pice posuitque intus infantulum et exposuit eum in carecto ripae fluminis
EXOD|2|4|stante procul sorore eius et considerante eventum rei
EXOD|2|5|ecce autem descendebat filia Pharaonis ut lavaretur in flumine et puellae eius gradiebantur per crepidinem alvei quae cum vidisset fiscellam in papyrione misit unam e famulis suis et adlatam
EXOD|2|6|aperiens cernensque in ea parvulum vagientem miserta eius ait de infantibus Hebraeorum est
EXOD|2|7|cui soror pueri vis inquit ut vadam et vocem tibi hebraeam mulierem quae nutrire possit infantulum
EXOD|2|8|respondit vade perrexit puella et vocavit matrem eius
EXOD|2|9|ad quam locuta filia Pharaonis accipe ait puerum istum et nutri mihi ego tibi dabo mercedem tuam suscepit mulier et nutrivit puerum adultumque tradidit filiae Pharaonis
EXOD|2|10|quem illa adoptavit in locum filii vocavitque nomen eius Mosi dicens quia de aqua tuli eum
EXOD|2|11|in diebus illis postquam creverat Moses egressus ad fratres suos vidit adflictionem eorum et virum aegyptium percutientem quendam de Hebraeis fratribus suis
EXOD|2|12|cumque circumspexisset huc atque illuc et nullum adesse vidisset percussum Aegyptium abscondit sabulo
EXOD|2|13|et egressus die altero conspexit duos Hebraeos rixantes dixitque ei qui faciebat iniuriam quare percutis proximum tuum
EXOD|2|14|qui respondit quis constituit te principem et iudicem super nos num occidere me tu dicis sicut occidisti Aegyptium timuit Moses et ait quomodo palam factum est verbum istud
EXOD|2|15|audivitque Pharao sermonem hunc et quaerebat occidere Mosen qui fugiens de conspectu eius moratus est in terra Madian et sedit iuxta puteum
EXOD|2|16|erant sacerdoti Madian septem filiae quae venerunt ad hauriendas aquas et impletis canalibus adaquare cupiebant greges patris sui
EXOD|2|17|supervenere pastores et eiecerunt eas surrexitque Moses et defensis puellis adaquavit oves earum
EXOD|2|18|quae cum revertissent ad Raguhel patrem suum dixit ad eas cur velocius venistis solito
EXOD|2|19|responderunt vir aegyptius liberavit nos de manu pastorum insuper et hausit aquam nobiscum potumque dedit ovibus
EXOD|2|20|at ille ubi est inquit quare dimisistis hominem vocate eum ut comedat panem
EXOD|2|21|iuravit ergo Moses quod habitaret cum eo accepitque Sefforam filiam eius
EXOD|2|22|quae peperit filium quem vocavit Gersam dicens advena fui in terra aliena
EXOD|2|23|post multum temporis mortuus est rex Aegypti et ingemescentes filii Israhel propter opera vociferati sunt ascenditque clamor eorum ad Deum ab operibus
EXOD|2|24|et audivit gemitum eorum ac recordatus foederis quod pepigerat cum Abraham et Isaac et Iacob
EXOD|2|25|respexit filios Israhel et cognovit eos
EXOD|3|1|Moses autem pascebat oves Iethro cognati sui sacerdotis Madian cumque minasset gregem ad interiora deserti venit ad montem Dei Horeb
EXOD|3|2|apparuitque ei Dominus in flamma ignis de medio rubi et videbat quod rubus arderet et non conbureretur
EXOD|3|3|dixit ergo Moses vadam et videbo visionem hanc magnam quare non conburatur rubus
EXOD|3|4|cernens autem Dominus quod pergeret ad videndum vocavit eum de medio rubi et ait Moses Moses qui respondit adsum
EXOD|3|5|at ille ne adpropies inquit huc solve calciamentum de pedibus tuis locus enim in quo stas terra sancta est
EXOD|3|6|et ait ego sum Deus patris tui Deus Abraham Deus Isaac Deus Iacob abscondit Moses faciem suam non enim audebat aspicere contra Deum
EXOD|3|7|cui ait Dominus vidi adflictionem populi mei in Aegypto et clamorem eius audivi propter duritiam eorum qui praesunt operibus
EXOD|3|8|et sciens dolorem eius descendi ut liberarem eum de manibus Aegyptiorum et educerem de terra illa in terram bonam et spatiosam in terram quae fluit lacte et melle ad loca Chananei et Hetthei et Amorrei Ferezei et Evei et Iebusei
EXOD|3|9|clamor ergo filiorum Israhel venit ad me vidique adflictionem eorum qua ab Aegyptiis opprimuntur
EXOD|3|10|sed veni mittam te ad Pharaonem ut educas populum meum filios Israhel de Aegypto
EXOD|3|11|dixit Moses ad Deum quis ego sum ut vadam ad Pharaonem et educam filios Israhel de Aegypto
EXOD|3|12|qui dixit ei ero tecum et hoc habebis signum quod miserim te cum eduxeris populum de Aegypto immolabis Deo super montem istum
EXOD|3|13|ait Moses ad Deum ecce ego vadam ad filios Israhel et dicam eis Deus patrum vestrorum misit me ad vos si dixerint mihi quod est nomen eius quid dicam eis
EXOD|3|14|dixit Deus ad Mosen ego sum qui sum ait sic dices filiis Israhel qui est misit me ad vos
EXOD|3|15|dixitque iterum Deus ad Mosen haec dices filiis Israhel Dominus Deus patrum vestrorum Deus Abraham Deus Isaac et Deus Iacob misit me ad vos hoc nomen mihi est in aeternum et hoc memoriale meum in generationem et generatione
EXOD|3|16|vade congrega seniores Israhel et dices ad eos Dominus Deus patrum vestrorum apparuit mihi Deus Abraham et Deus Isaac et Deus Iacob dicens visitans visitavi vos et omnia quae acciderunt vobis in Aegypto
EXOD|3|17|et dixi ut educam vos de adflictione Aegypti in terram Chananei et Hetthei et Amorrei Ferezei et Evei et Iebusei ad terram fluentem lacte et melle
EXOD|3|18|et audient vocem tuam ingredierisque tu et seniores Israhel ad regem Aegypti et dices ad eum Dominus Deus Hebraeorum vocavit nos ibimus viam trium dierum per solitudinem ut immolemus Domino Deo nostro
EXOD|3|19|sed ego scio quod non dimittet vos rex Aegypti ut eatis nisi per manum validam
EXOD|3|20|extendam enim manum meam et percutiam Aegyptum in cunctis mirabilibus meis quae facturus sum in medio eorum post haec dimittet vos
EXOD|3|21|daboque gratiam populo huic coram Aegyptiis et cum egrediemini non exibitis vacui
EXOD|3|22|sed postulabit mulier a vicina sua et ab hospita vasa argentea et aurea ac vestes ponetisque eas super filios et filias vestras et spoliabitis Aegyptum
EXOD|4|1|respondens Moses ait non credent mihi neque audient vocem meam sed dicent non apparuit tibi Dominus
EXOD|4|2|dixit ergo ad eum quid est hoc quod tenes in manu tua respondit virga
EXOD|4|3|ait proice eam in terram proiecit et versa est in colubrum ita ut fugeret Moses
EXOD|4|4|dixitque Dominus extende manum tuam et adprehende caudam eius extendit et tenuit versaque est in virgam
EXOD|4|5|ut credant inquit quod apparuerit tibi Dominus Deus patrum tuorum Deus Abraham Deus Isaac Deus Iacob
EXOD|4|6|dixitque Dominus rursum mitte manum in sinum tuum quam cum misisset in sinum protulit leprosam instar nivis
EXOD|4|7|retrahe ait manum in sinum tuum retraxit et protulit iterum et erat similis carni reliquae
EXOD|4|8|si non crediderint inquit tibi neque audierint sermonem signi prioris credent verbo signi sequentis
EXOD|4|9|quod si nec duobus quidem his signis crediderint neque audierint vocem tuam sume aquam fluminis et effunde eam super aridam et quicquid hauseris de fluvio vertetur in sanguinem
EXOD|4|10|ait Moses obsecro Domine non sum eloquens ab heri et nudius tertius et ex quo locutus es ad servum tuum inpeditioris et tardioris linguae sum
EXOD|4|11|dixit Dominus ad eum quis fecit os hominis aut quis fabricatus est mutum et surdum videntem et caecum nonne ego
EXOD|4|12|perge igitur et ego ero in ore tuo doceboque te quid loquaris
EXOD|4|13|at ille obsecro inquit Domine mitte quem missurus es
EXOD|4|14|iratus Dominus in Mosen ait Aaron frater tuus Levites scio quod eloquens sit ecce ipse egreditur in occursum tuum vidensque te laetabitur corde
EXOD|4|15|loquere ad eum et pone verba mea in ore eius ego ero in ore tuo et in ore illius et ostendam vobis quid agere debeatis
EXOD|4|16|ipse loquetur pro te ad populum et erit os tuum tu autem eris ei in his quae ad Deum pertinent
EXOD|4|17|virgam quoque hanc sume in manu tua in qua facturus es signa
EXOD|4|18|abiit Moses et reversus est ad Iethro cognatum suum dixitque ei vadam et revertar ad fratres meos in Aegyptum ut videam si adhuc vivunt cui ait Iethro vade in pace
EXOD|4|19|dixit ergo Dominus ad Mosen in Madian vade revertere in Aegyptum mortui sunt omnes qui quaerebant animam tuam
EXOD|4|20|tulit Moses uxorem et filios suos et inposuit eos super asinum reversusque est in Aegyptum portans virgam Dei in manu sua
EXOD|4|21|dixitque ei Dominus revertenti in Aegyptum vide ut omnia ostenta quae posui in manu tua facias coram Pharaone ego indurabo cor eius et non dimittet populum
EXOD|4|22|dicesque ad eum haec dicit Dominus filius meus primogenitus meus Israhel
EXOD|4|23|dixi tibi dimitte filium meum ut serviat mihi et noluisti dimittere eum ecce ego interficiam filium tuum primogenitum
EXOD|4|24|cumque esset in itinere in diversorio occurrit ei Dominus et volebat occidere eum
EXOD|4|25|tulit ilico Seffora acutissimam petram et circumcidit praeputium filii sui tetigitque pedes eius et ait sponsus sanguinum tu mihi es
EXOD|4|26|et dimisit eum postquam dixerat sponsus sanguinum ob circumcisionem
EXOD|4|27|dixit autem Dominus ad Aaron vade in occursum Mosi in deserto qui perrexit ei obviam in montem Dei et osculatus est eum
EXOD|4|28|narravitque Moses Aaron omnia verba Domini quibus miserat eum et signa quae mandaverat
EXOD|4|29|veneruntque simul et congregaverunt cunctos seniores filiorum Israhel
EXOD|4|30|locutusque est Aaron omnia verba quae dixerat Dominus ad Mosen et fecit signa coram populo
EXOD|4|31|et credidit populus audieruntque quod visitasset Dominus filios Israhel et quod respexisset adflictionem eorum et proni adoraverunt
EXOD|5|1|post haec ingressi sunt Moses et Aaron et dixerunt Pharaoni haec dicit Dominus Deus Israhel dimitte populum meum ut sacrificet mihi in deserto
EXOD|5|2|at ille respondit quis est Dominus ut audiam vocem eius et dimittam Israhel nescio Dominum et Israhel non dimittam
EXOD|5|3|dixerunt Deus Hebraeorum vocavit nos ut eamus viam trium dierum in solitudinem et sacrificemus Domino Deo nostro ne forte accidat nobis pestis aut gladius
EXOD|5|4|ait ad eos rex Aegypti quare Moses et Aaron sollicitatis populum ab operibus suis ite ad onera vestra
EXOD|5|5|dixitque Pharao multus est populus terrae videtis quod turba succreverit quanto magis si dederitis eis requiem ab operibus
EXOD|5|6|praecepit ergo in die illo praefectis operum et exactoribus populi dicens
EXOD|5|7|nequaquam ultra dabitis paleas populo ad conficiendos lateres sicut prius sed ipsi vadant et colligant stipulam
EXOD|5|8|et mensuram laterum quos prius faciebant inponetis super eos nec minuetis quicquam vacant enim et idcirco vociferantur dicentes eamus et sacrificemus Deo nostro
EXOD|5|9|opprimantur operibus et expleant ea ut non adquiescant verbis mendacibus
EXOD|5|10|igitur egressi praefecti operum et exactores ad populum dixerunt sic dicit Pharao non do vobis paleas
EXOD|5|11|ite et colligite sicubi invenire potueritis nec minuetur quicquam de opere vestro
EXOD|5|12|dispersusque est populus per omnem terram Aegypti ad colligendas paleas
EXOD|5|13|praefecti quoque operum instabant dicentes conplete opus vestrum cotidie ut prius facere solebatis quando dabantur vobis paleae
EXOD|5|14|flagellatique sunt qui praeerant operibus filiorum Israhel ab exactoribus Pharaonis dicentibus quare non impletis mensuram laterum sicut prius nec heri nec hodie
EXOD|5|15|veneruntque praepositi filiorum Israhel et vociferati sunt ad Pharaonem dicentes cur ita agis contra servos tuos
EXOD|5|16|paleae non dantur nobis et lateres similiter imperantur en famuli tui flagellis caedimur et iniuste agitur contra populum tuum
EXOD|5|17|qui ait vacatis otio et idcirco dicitis eamus et sacrificemus Domino
EXOD|5|18|ite ergo et operamini paleae non dabuntur vobis et reddetis consuetum numerum laterum
EXOD|5|19|videbantque se praepositi filiorum Israhel in malo eo quod diceretur eis non minuetur quicquam de lateribus per singulos dies
EXOD|5|20|occurreruntque Mosi et Aaron qui stabant ex adverso egredientes a Pharaone
EXOD|5|21|et dixerunt ad eos videat Dominus et iudicet quoniam fetere fecistis odorem nostrum coram Pharao et servis eius et praebuistis ei gladium ut occideret nos
EXOD|5|22|reversusque Moses ad Dominum ait Domine cur adflixisti populum istum quare misisti me
EXOD|5|23|ex eo enim quo ingressus sum ad Pharaonem ut loquerer nomine tuo adflixit populum tuum et non liberasti eos
EXOD|6|1|dixit Dominus ad Mosen nunc videbis quae facturus sum Pharaoni per manum enim fortem dimittet eos et in manu robusta eiciet illos de terra sua
EXOD|6|2|locutusque est Dominus ad Mosen dicens ego Dominus
EXOD|6|3|qui apparui Abraham Isaac et Iacob in Deo omnipotente et nomen meum Adonai non indicavi eis
EXOD|6|4|pepigique cum eis foedus ut darem illis terram Chanaan terram peregrinationis eorum in qua fuerunt advenae
EXOD|6|5|ego audivi gemitum filiorum Israhel quo Aegyptii oppresserunt eos et recordatus sum pacti mei
EXOD|6|6|ideo dic filiis Israhel ego Dominus qui educam vos de ergastulo Aegyptiorum et eruam de servitute ac redimam in brachio excelso et iudiciis magnis
EXOD|6|7|et adsumam vos mihi in populum et ero vester Deus scietisque quod ego sim Dominus Deus vester qui eduxerim vos de ergastulo Aegyptiorum
EXOD|6|8|et induxerim in terram super quam levavi manum meam ut darem eam Abraham Isaac et Iacob daboque illam vobis possidendam ego Dominus
EXOD|6|9|narravit ergo Moses omnia filiis Israhel qui non adquieverunt ei propter angustiam spiritus et opus durissimum
EXOD|6|10|locutusque est Dominus ad Mosen dicens
EXOD|6|11|ingredere et loquere ad Pharao regem Aegypti ut dimittat filios Israhel de terra sua
EXOD|6|12|respondit Moses coram Domino ecce filii Israhel non me audiunt et quomodo audiet me Pharao praesertim cum sim incircumcisus labiis
EXOD|6|13|locutus est Dominus ad Mosen et Aaron et dedit mandatum ad filios Israhel et ad Pharao regem Aegypti ut educerent filios Israhel de terra Aegypti
EXOD|6|14|isti sunt principes domorum per familias suas filii Ruben primogeniti Israhelis Enoch et Phallu Aesrom et Charmi
EXOD|6|15|hae cognationes Ruben filii Symeon Iamuhel et Iamin et Aod Iachin et Soer et Saul filius Chananitidis hae progenies Symeon
EXOD|6|16|et haec nomina filiorum Levi per cognationes suas Gerson et Caath et Merari anni autem vitae Levi fuerunt centum triginta septem
EXOD|6|17|filii Gerson Lobeni et Semei per cognationes suas
EXOD|6|18|filii Caath Amram et Isuar et Hebron et Ozihel annique vitae Caath centum triginta tres
EXOD|6|19|filii Merari Mooli et Musi hae cognationes Levi per familias suas
EXOD|6|20|accepit autem Amram uxorem Iocabed patruelem suam quae peperit ei Aaron et Mosen fueruntque anni vitae Amram centum triginta septem
EXOD|6|21|filii quoque Isuar Core et Napheg et Zechri
EXOD|6|22|filii quoque Ozihel Misahel et Elsaphan et Sethri
EXOD|6|23|accepit autem Aaron uxorem Elisabe filiam Aminadab sororem Naasson quae peperit ei Nadab et Abiu et Eleazar et Ithamar
EXOD|6|24|filii quoque Core Asir et Helcana et Abiasab hae sunt cognationes Coritarum
EXOD|6|25|at vero Eleazar filius Aaron accepit uxorem de filiabus Phutihel quae peperit ei Finees hii sunt principes familiarum leviticarum per cognationes suas
EXOD|6|26|iste est Aaron et Moses quibus praecepit Dominus ut educerent filios Israhel de terra Aegypti per turmas suas
EXOD|6|27|hii sunt qui loquuntur ad Pharao regem Aegypti ut educant filios Israhel de Aegypto iste Moses et Aaron
EXOD|6|28|in die qua locutus est Dominus ad Mosen in terra Aegypti
EXOD|6|29|et locutus est Dominus ad Mosen dicens ego Dominus loquere ad Pharao regem Aegypti omnia quae ego loquor tibi
EXOD|6|30|et ait Moses coram Domino en incircumcisus labiis sum quomodo audiet me Pharao
EXOD|7|1|dixitque Dominus ad Mosen ecce constitui te Deum Pharaonis Aaron frater tuus erit propheta tuus
EXOD|7|2|tu loqueris omnia quae mando tibi ille loquetur ad Pharaonem ut dimittat filios Israhel de terra sua
EXOD|7|3|sed ego indurabo cor eius et multiplicabo signa et ostenta mea in terra Aegypti
EXOD|7|4|et non audiet vos inmittamque manum meam super Aegyptum et educam exercitum et populum meum filios Israhel de terra Aegypti per iudicia maxima
EXOD|7|5|et scient Aegyptii quod ego sim Dominus qui extenderim manum meam super Aegyptum et eduxerim filios Israhel de medio eorum
EXOD|7|6|fecit itaque Moses et Aaron sicut praeceperat Dominus ita egerunt
EXOD|7|7|erat autem Moses octoginta annorum et Aaron octoginta trium quando locuti sunt ad Pharaonem
EXOD|7|8|dixitque Dominus ad Mosen et Aaron
EXOD|7|9|cum dixerit vobis Pharao ostendite signa dices ad Aaron tolle virgam tuam et proice eam coram Pharao ac vertatur in colubrum
EXOD|7|10|ingressi itaque Moses et Aaron ad Pharaonem fecerunt sicut praeceperat Dominus tulitque Aaron virgam coram Pharao et servis eius quae versa est in colubrum
EXOD|7|11|vocavit autem Pharao sapientes et maleficos et fecerunt etiam ipsi per incantationes aegyptias et arcana quaedam similiter
EXOD|7|12|proieceruntque singuli virgas suas quae versae sunt in dracones sed devoravit virga Aaron virgas eorum
EXOD|7|13|induratumque est cor Pharaonis et non audivit eos sicut praeceperat Dominus
EXOD|7|14|dixit autem Dominus ad Mosen ingravatum est cor Pharaonis non vult dimittere populum
EXOD|7|15|vade ad eum mane ecce egredietur ad aquas et stabis in occursum eius super ripam fluminis et virgam quae conversa est in draconem tolles in manu tua
EXOD|7|16|dicesque ad eum Dominus Deus Hebraeorum misit me ad te dicens dimitte populum meum ut mihi sacrificet in deserto et usque ad praesens audire noluisti
EXOD|7|17|haec igitur dicit Dominus in hoc scies quod Dominus sim ecce percutiam virga quae in manu mea est aquam fluminis et vertetur in sanguinem
EXOD|7|18|pisces quoque qui sunt in fluvio morientur et conputrescent aquae et adfligentur Aegyptii bibentes aquam fluminis
EXOD|7|19|dixit quoque Dominus ad Mosen dic ad Aaron tolle virgam tuam et extende manum tuam super aquas Aegypti et super fluvios eorum et rivos ac paludes et omnes lacus aquarum ut vertantur in sanguinem et sit cruor in omni terra Aegypti tam in ligneis vasis quam in saxeis
EXOD|7|20|feceruntque ita Moses et Aaron sicut praeceperat Dominus et elevans virgam percussit aquam fluminis coram Pharao et servis eius quae versa est in sanguinem
EXOD|7|21|et pisces qui erant in flumine mortui sunt conputruitque fluvius et non poterant Aegyptii bibere aquam fluminis et fuit sanguis in tota terra Aegypti
EXOD|7|22|feceruntque similiter malefici Aegyptiorum incantationibus suis et induratum est cor Pharaonis nec audivit eos sicut praeceperat Dominus
EXOD|7|23|avertitque se et ingressus est domum suam nec adposuit cor etiam hac vice
EXOD|7|24|foderunt autem omnes Aegyptii per circuitum fluminis aquam ut biberent non enim poterant bibere de aqua fluminis
EXOD|7|25|impletique sunt septem dies postquam percussit Dominus fluvium
EXOD|8|1|dixitque Dominus ad Mosen ingredere ad Pharao et dices ad eum haec dicit Dominus dimitte populum meum ut sacrificet mihi
EXOD|8|2|sin autem nolueris dimittere ecce ego percutiam omnes terminos tuos ranis
EXOD|8|3|et ebulliet fluvius ranas quae ascendent et ingredientur domum tuam et cubiculum lectuli tui et super stratum tuum et in domos servorum tuorum et in populum tuum et in furnos tuos et in reliquias ciborum tuorum
EXOD|8|4|et ad te et ad populum tuum et ad omnes servos tuos intrabunt ranae
EXOD|8|5|dixitque Dominus ad Mosen dic Aaron extende manum tuam super fluvios et super rivos ac paludes et educ ranas super terram Aegypti
EXOD|8|6|extendit Aaron manum super aquas Aegypti et ascenderunt ranae operueruntque terram Aegypti
EXOD|8|7|fecerunt autem et malefici per incantationes suas similiter eduxeruntque ranas super terram Aegypti
EXOD|8|8|vocavit autem Pharao Mosen et Aaron et dixit orate Dominum ut auferat ranas a me et a populo meo et dimittam populum ut sacrificet Domino
EXOD|8|9|dixitque Moses Pharaoni constitue mihi quando deprecer pro te et pro servis tuis et pro populo tuo ut abigantur ranae a te et a domo tua et tantum in flumine remaneant
EXOD|8|10|qui respondit cras at ille iuxta verbum inquit tuum ut scias quoniam non est sicut Dominus Deus noster
EXOD|8|11|et recedent ranae a te et a domo tua et a servis tuis et a populo tuo tantum in flumine remanebunt
EXOD|8|12|egressique sunt Moses et Aaron a Pharaone et clamavit Moses ad Dominum pro sponsione ranarum quam condixerat Pharaoni
EXOD|8|13|fecitque Dominus iuxta verbum Mosi et mortuae sunt ranae de domibus et de villis et de agris
EXOD|8|14|congregaveruntque eas in inmensos aggeres et conputruit terra
EXOD|8|15|videns autem Pharao quod data esset requies ingravavit cor suum et non audivit eos sicut praeceperat Dominus
EXOD|8|16|dixitque Dominus ad Mosen loquere ad Aaron extende virgam tuam et percute pulverem terrae et sint scinifes in universa terra Aegypti
EXOD|8|17|feceruntque ita et extendit Aaron manu virgam tenens percussitque pulverem terrae et facti sunt scinifes in hominibus et in iumentis omnis pulvis terrae versus est in scinifes per totam terram Aegypti
EXOD|8|18|feceruntque similiter malefici incantationibus suis ut educerent scinifes et non potuerunt erantque scinifes tam in hominibus quam in iumentis
EXOD|8|19|et dixerunt malefici ad Pharao digitus Dei est induratumque est cor Pharaonis et non audivit eos sicut praeceperat Dominus
EXOD|8|20|dixit quoque Dominus ad Mosen consurge diluculo et sta coram Pharaone egreditur enim ad aquas et dices ad eum haec dicit Dominus dimitte populum meum ut sacrificet mihi
EXOD|8|21|quod si non dimiseris eum ecce ego inmittam in te et in servos tuos et in populum tuum et in domos tuas omne genus muscarum et implebuntur domus Aegyptiorum muscis diversi generis et in universa terra in qua fuerint
EXOD|8|22|faciamque mirabilem in die illa terram Gessen in qua populus meus est ut non sint ibi muscae et scias quoniam ego Dominus in medio terrae
EXOD|8|23|ponamque divisionem inter populum meum et populum tuum cras erit signum istud
EXOD|8|24|fecitque Dominus ita et venit musca gravissima in domos Pharaonis et servorum eius et in omnem terram Aegypti corruptaque est terra ab huiuscemodi muscis
EXOD|8|25|vocavit Pharao Mosen et Aaron et ait eis ite sacrificate Deo vestro in terra
EXOD|8|26|et ait Moses non potest ita fieri abominationes enim Aegyptiorum immolabimus Domino Deo nostro quod si mactaverimus ea quae colunt Aegyptii coram eis lapidibus nos obruent
EXOD|8|27|via trium dierum pergemus in solitudine et sacrificabimus Domino Deo nostro sicut praeceperit nobis
EXOD|8|28|dixitque Pharao ego dimittam vos ut sacrificetis Domino Deo vestro in deserto verumtamen longius ne abeatis rogate pro me
EXOD|8|29|et ait Moses egressus a te orabo Dominum et recedet musca a Pharaone et a servis et a populo eius cras verumtamen noli ultra fallere ut non dimittas populum sacrificare Domino
EXOD|8|30|egressusque Moses a Pharao oravit Dominum
EXOD|8|31|qui fecit iuxta verbum illius et abstulit muscas a Pharao et a servis et a populo eius non superfuit ne una quidem
EXOD|8|32|et ingravatum est cor Pharaonis ita ut ne hac quidem vice dimitteret populum
EXOD|9|1|dixit autem Dominus ad Mosen ingredere ad Pharaonem et loquere ad eum haec dicit Dominus Deus Hebraeorum dimitte populum meum ut sacrificet mihi
EXOD|9|2|quod si adhuc rennuis et retines eos
EXOD|9|3|ecce manus mea erit super agros tuos et super equos et asinos et camelos et boves et oves pestis valde gravis
EXOD|9|4|et faciet Dominus mirabile inter possessiones Israhel et possessiones Aegyptiorum ut nihil omnino intereat ex his quae pertinent ad filios Israhel
EXOD|9|5|constituitque Dominus tempus dicens cras faciet Dominus verbum istud in terra
EXOD|9|6|fecit ergo Dominus verbum hoc altero die mortuaque sunt omnia animantia Aegyptiorum de animalibus vero filiorum Israhel nihil omnino periit
EXOD|9|7|et misit Pharao ad videndum nec erat quicquam mortuum de his quae possidebat Israhel ingravatumque est cor Pharaonis et non dimisit populum
EXOD|9|8|et dixit Dominus ad Mosen et Aaron tollite plenas manus cineris de camino et spargat illud Moses in caelum coram Pharao
EXOD|9|9|sitque pulvis super omnem terram Aegypti erunt enim in hominibus et in iumentis vulnera et vesicae turgentes in universa terra Aegypti
EXOD|9|10|tuleruntque cinerem de camino et steterunt contra Pharao et sparsit illud Moses in caelum factaque sunt vulnera vesicarum turgentium in hominibus et in iumentis
EXOD|9|11|nec poterant malefici stare coram Mosen propter vulnera quae in illis erant et in omni terra Aegypti
EXOD|9|12|induravitque Dominus cor Pharaonis et non audivit eos sicut locutus est Dominus ad Mosen
EXOD|9|13|dixit quoque Dominus ad Mosen mane consurge et sta coram Pharao et dices ad eum haec dicit Dominus Deus Hebraeorum dimitte populum meum ut sacrificet mihi
EXOD|9|14|quia in hac vice mittam omnes plagas meas super cor tuum super servos tuos et super populum tuum ut scias quod non sit similis mei in omni terra
EXOD|9|15|nunc enim extendens manum percutiam te et populum tuum peste peribisque de terra
EXOD|9|16|idcirco autem posui te ut ostendam in te fortitudinem meam et narretur nomen meum in omni terra
EXOD|9|17|adhuc retines populum meum et non vis eum dimittere
EXOD|9|18|en pluam hac ipsa hora cras grandinem multam nimis qualis non fuit in Aegypto a die qua fundata est usque in praesens tempus
EXOD|9|19|mitte ergo iam nunc et congrega iumenta tua et omnia quae habes in agro homines enim et iumenta et universa quae inventa fuerint foris nec congregata de agris cecideritque super ea grando morientur
EXOD|9|20|qui timuit verbum Domini de servis Pharao fecit confugere servos suos et iumenta in domos
EXOD|9|21|qui autem neglexit sermonem Domini dimisit servos suos et iumenta in agris
EXOD|9|22|et dixit Dominus ad Mosen extende manum tuam in caelum ut fiat grando in universa terra Aegypti super homines et super iumenta et super omnem herbam agri in terra Aegypti
EXOD|9|23|extenditque Moses virgam in caelum et Dominus dedit tonitrua et grandinem ac discurrentia fulgura super terram pluitque Dominus grandinem super terram Aegypti
EXOD|9|24|et grando et ignis inmixta pariter ferebantur tantaeque fuit magnitudinis quanta ante numquam apparuit in universa terra Aegypti ex quo gens illa condita est
EXOD|9|25|et percussit grando in omni terra Aegypti cuncta quae fuerunt in agris ab homine usque ad iumentum cunctam herbam agri percussit grando et omne lignum regionis confregit
EXOD|9|26|tantum in terra Gessen ubi erant filii Israhel grando non cecidit
EXOD|9|27|misitque Pharao et vocavit Mosen et Aaron dicens ad eos peccavi etiam nunc Dominus iustus ego et populus meus impii
EXOD|9|28|orate Dominum et desinant tonitrua Dei et grando ut dimittam vos et nequaquam hic ultra maneatis
EXOD|9|29|ait Moses cum egressus fuero de urbe extendam palmas meas ad Dominum et cessabunt tonitrua et grando non erit ut scias quia Domini est terra
EXOD|9|30|novi autem quod et tu et servi tui necdum timeatis Dominum Deum
EXOD|9|31|linum ergo et hordeum laesum est eo quod hordeum esset virens et linum iam folliculos germinaret
EXOD|9|32|triticum autem et far non sunt laesa quia serotina erant
EXOD|9|33|egressusque Moses a Pharaone et ex urbe tetendit manus ad Dominum et cessaverunt tonitrua et grando nec ultra stillavit pluvia super terram
EXOD|9|34|videns autem Pharao quod cessasset pluvia et grando et tonitrua auxit peccatum
EXOD|9|35|et ingravatum est cor eius et servorum illius et induratum nimis nec dimisit filios Israhel sicut praeceperat Dominus per manum Mosi
EXOD|10|1|et dixit Dominus ad Mosen ingredere ad Pharao ego enim induravi cor eius et servorum illius ut faciam signa mea haec in eo
EXOD|10|2|et narres in auribus filii tui et nepotum tuorum quotiens contriverim Aegyptios et signa mea fecerim in eis et sciatis quia ego Dominus
EXOD|10|3|introierunt ergo Moses et Aaron ad Pharaonem et dixerunt ad eum haec dicit Dominus Deus Hebraeorum usquequo non vis subici mihi dimitte populum meum ut sacrificet mihi
EXOD|10|4|sin autem resistis et non vis dimittere eum ecce ego inducam cras lucustam in fines tuos
EXOD|10|5|quae operiat superficiem terrae nec quicquam eius appareat sed comedatur quod residuum fuit grandini conrodet enim omnia ligna quae germinant in agris
EXOD|10|6|et implebunt domos tuas et servorum tuorum et omnium Aegyptiorum quantam non viderunt patres tui et avi ex quo orti sunt super terram usque in praesentem diem avertitque se et egressus est a Pharaone
EXOD|10|7|dixerunt autem servi Pharaonis ad eum usquequo patiemur hoc scandalum dimitte homines ut sacrificent Domino Deo suo nonne vides quod perierit Aegyptus
EXOD|10|8|revocaveruntque Mosen et Aaron ad Pharaonem qui dixit eis ite sacrificate Domino Deo vestro quinam sunt qui ituri sunt
EXOD|10|9|ait Moses cum parvulis nostris et senibus pergemus cum filiis et filiabus cum ovibus et armentis est enim sollemnitas Domini nostri
EXOD|10|10|et respondit sic Dominus sit vobiscum quomodo ego dimittam vos et parvulos vestros cui dubium est quod pessime cogitetis
EXOD|10|11|non fiet ita sed ite tantum viri et sacrificate Domino hoc enim et ipsi petistis statimque eiecti sunt de conspectu Pharaonis
EXOD|10|12|dixit autem Dominus ad Mosen extende manum tuam super terram Aegypti ad lucustam ut ascendat super eam et devoret omnem herbam quae residua fuit grandini
EXOD|10|13|extendit Moses virgam super terram Aegypti et Dominus induxit ventum urentem tota illa die ac nocte et mane facto ventus urens levavit lucustas
EXOD|10|14|quae ascenderunt super universam terram Aegypti et sederunt in cunctis finibus Aegyptiorum innumerabiles quales ante illud tempus non fuerant nec postea futurae sunt
EXOD|10|15|operueruntque universam superficiem terrae vastantes omnia devorata est igitur herba terrae et quicquid pomorum in arboribus fuit quae grando dimiserat nihilque omnino virens relictum est in lignis et in herbis terrae in cuncta Aegypto
EXOD|10|16|quam ob rem festinus Pharao vocavit Mosen et Aaron et dixit eis peccavi in Dominum Deum vestrum et in vos
EXOD|10|17|sed nunc dimittite peccatum mihi etiam hac vice et rogate Dominum Deum vestrum ut auferat a me mortem istam
EXOD|10|18|egressusque est de conspectu Pharaonis et oravit Dominum
EXOD|10|19|qui flare fecit ventum ab occidente vehementissimum et arreptam lucustam proiecit in mare Rubrum non remansit ne una quidem in cunctis finibus Aegypti
EXOD|10|20|et induravit Dominus cor Pharaonis nec dimisit filios Israhel
EXOD|10|21|dixit autem Dominus ad Mosen extende manum tuam in caelum et sint tenebrae super terram Aegypti tam densae ut palpari queant
EXOD|10|22|extendit Moses manum in caelum et factae sunt tenebrae horribiles in universa terra Aegypti tribus diebus
EXOD|10|23|nemo vidit fratrem suum nec movit se de loco in quo erat ubicumque autem habitabant filii Israhel lux erat
EXOD|10|24|vocavitque Pharao Mosen et Aaron et dixit eis ite sacrificate Domino oves tantum vestrae et armenta remaneant parvuli vestri eant vobiscum
EXOD|10|25|ait Moses hostias quoque et holocausta dabis nobis quae offeramus Domino Deo nostro
EXOD|10|26|cuncti greges pergent nobiscum non remanebit ex eis ungula quae necessaria sunt in cultum Domini Dei nostri praesertim cum ignoremus quid debeat immolari donec ad ipsum locum perveniamus
EXOD|10|27|induravit autem Dominus cor Pharaonis et noluit dimittere eos
EXOD|10|28|dixitque Pharao ad eum recede a me cave ne ultra videas faciem meam quocumque die apparueris mihi morieris
EXOD|10|29|respondit Moses ita fiat ut locutus es non videbo ultra faciem tuam
EXOD|11|1|et dixit Dominus ad Mosen adhuc una plaga tangam Pharaonem et Aegyptum et post haec dimittet vos et exire conpellet
EXOD|11|2|dices ergo omni plebi ut postulet vir ab amico suo et mulier a vicina sua vasa argentea et aurea
EXOD|11|3|dabit autem Dominus gratiam populo coram Aegyptiis fuitque Moses vir magnus valde in terra Aegypti coram servis Pharao et omni populo
EXOD|11|4|et ait haec dicit Dominus media nocte egrediar in Aegyptum
EXOD|11|5|et morietur omne primogenitum in terra Aegyptiorum a primogenito Pharaonis qui sedet in solio eius usque ad primogenitum ancillae quae est ad molam et omnia primogenita iumentorum
EXOD|11|6|eritque clamor magnus in universa terra Aegypti qualis nec ante fuit nec postea futurus est
EXOD|11|7|apud omnes autem filios Israhel non muttiet canis ab homine usque ad pecus ut sciatis quanto miraculo dividat Dominus Aegyptios et Israhel
EXOD|11|8|descendentque omnes servi tui isti ad me et adorabunt me dicentes egredere tu et omnis populus qui subiectus est tibi post haec egrediemur
EXOD|11|9|et exivit a Pharaone iratus nimis dixit autem Dominus ad Mosen non audiet vos Pharao ut multa signa fiant in terra Aegypti
EXOD|11|10|Moses autem et Aaron fecerunt omnia ostenta quae scripta sunt coram Pharaone et induravit Dominus cor Pharaonis nec dimisit filios Israhel de terra sua
EXOD|12|1|dixit quoque Dominus ad Mosen et Aaron in terra Aegypti
EXOD|12|2|mensis iste vobis principium mensuum primus erit in mensibus anni
EXOD|12|3|loquimini ad universum coetum filiorum Israhel et dicite eis decima die mensis huius tollat unusquisque agnum per familias et domos suas
EXOD|12|4|sin autem minor est numerus ut sufficere possit ad vescendum agnum adsumet vicinum suum qui iunctus est domui eius iuxta numerum animarum quae sufficere possunt ad esum agni
EXOD|12|5|erit autem agnus absque macula masculus anniculus iuxta quem ritum tolletis et hedum
EXOD|12|6|et servabitis eum usque ad quartamdecimam diem mensis huius immolabitque eum universa multitudo filiorum Israhel ad vesperam
EXOD|12|7|et sument de sanguine ac ponent super utrumque postem et in superliminaribus domorum in quibus comedent illum
EXOD|12|8|et edent carnes nocte illa assas igni et azymos panes cum lactucis agrestibus
EXOD|12|9|non comedetis ex eo crudum quid nec coctum aqua sed assum tantum igni caput cum pedibus eius et intestinis vorabitis
EXOD|12|10|nec remanebit ex eo quicquam usque mane si quid residui fuerit igne conburetis
EXOD|12|11|sic autem comedetis illum renes vestros accingetis calciamenta habebitis in pedibus tenentes baculos in manibus et comedetis festinantes est enim phase id est transitus Domini
EXOD|12|12|et transibo per terram Aegypti nocte illa percutiamque omne primogenitum in terra Aegypti ab homine usque ad pecus et in cunctis diis Aegypti faciam iudicia ego Dominus
EXOD|12|13|erit autem sanguis vobis in signum in aedibus in quibus eritis et videbo sanguinem ac transibo vos nec erit in vobis plaga disperdens quando percussero terram Aegypti
EXOD|12|14|habebitis autem hanc diem in monumentum et celebrabitis eam sollemnem Domino in generationibus vestris cultu sempiterno
EXOD|12|15|septem diebus azyma comedetis in die primo non erit fermentum in domibus vestris quicumque comederit fermentatum peribit anima illa de Israhel a primo die usque ad diem septimum
EXOD|12|16|dies prima erit sancta atque sollemnis et dies septima eadem festivitate venerabilis nihil operis facietis in eis exceptis his quae ad vescendum pertinent
EXOD|12|17|et observabitis azyma in eadem enim ipsa die educam exercitum vestrum de terra Aegypti et custodietis diem istum in generationes vestras ritu perpetuo
EXOD|12|18|primo mense quartadecima die mensis ad vesperam comedetis azyma usque ad diem vicesimam primam eiusdem mensis ad vesperam
EXOD|12|19|septem diebus fermentum non invenietur in domibus vestris qui comederit fermentatum peribit anima eius de coetu Israhel tam de advenis quam de indigenis terrae
EXOD|12|20|omne fermentatum non comedetis in cunctis habitaculis vestris edetis azyma
EXOD|12|21|vocavit autem Moses omnes seniores filiorum Israhel et dixit ad eos ite tollentes animal per familias vestras immolate phase
EXOD|12|22|fasciculumque hysopi tinguite sanguine qui est in limine et aspergite ex eo superliminare et utrumque postem nullus vestrum egrediatur ostium domus suae usque mane
EXOD|12|23|transibit enim Dominus percutiens Aegyptios cumque viderit sanguinem in superliminari et in utroque poste transcendet ostium et non sinet percussorem ingredi domos vestras et laedere
EXOD|12|24|custodi verbum istud legitimum tibi et filiis tuis usque in aeternum
EXOD|12|25|cumque introieritis terram quam Dominus daturus est vobis ut pollicitus est observabitis caerimonias istas
EXOD|12|26|et cum dixerint vobis filii vestri quae est ista religio
EXOD|12|27|dicetis eis victima transitus Domini est quando transivit super domos filiorum Israhel in Aegypto percutiens Aegyptios et domos nostras liberans incurvatusque populus adoravit
EXOD|12|28|et egressi filii Israhel fecerunt sicut praeceperat Dominus Mosi et Aaron
EXOD|12|29|factum est autem in noctis medio percussit Dominus omne primogenitum in terra Aegypti a primogenito Pharaonis qui sedebat in solio eius usque ad primogenitum captivae quae erat in carcere et omne primogenitum iumentorum
EXOD|12|30|surrexitque Pharao nocte et omnes servi eius cunctaque Aegyptus et ortus est clamor magnus in Aegypto neque enim erat domus in qua non iaceret mortuus
EXOD|12|31|vocatisque Mosen et Aaron nocte ait surgite egredimini a populo meo et vos et filii Israhel ite immolate Domino sicut dicitis
EXOD|12|32|oves vestras et armenta adsumite ut petieratis et abeuntes benedicite mihi
EXOD|12|33|urguebantque Aegyptii populum de terra exire velociter dicentes omnes moriemur
EXOD|12|34|tulit igitur populus conspersam farinam antequam fermentaretur et ligans in palliis posuit super umeros suos
EXOD|12|35|feceruntque filii Israhel sicut praeceperat Moses et petierunt ab Aegyptiis vasa argentea et aurea vestemque plurimam
EXOD|12|36|dedit autem Dominus gratiam populo coram Aegyptiis ut commodarent eis et spoliaverunt Aegyptios
EXOD|12|37|profectique sunt filii Israhel de Ramesse in Soccoth sescenta ferme milia peditum virorum absque parvulis
EXOD|12|38|sed et vulgus promiscuum innumerabile ascendit cum eis oves et armenta et animantia diversi generis multa nimis
EXOD|12|39|coxeruntque farinam quam dudum conspersam de Aegypto tulerant et fecerunt subcinericios panes azymos neque enim poterant fermentari cogentibus exire Aegyptiis et nullam facere sinentibus moram nec pulmenti quicquam occurrerant praeparare
EXOD|12|40|habitatio autem filiorum Israhel qua manserant in Aegypto fuit quadringentorum triginta annorum
EXOD|12|41|quibus expletis eadem die egressus est omnis exercitus Domini de terra Aegypti
EXOD|12|42|nox est ista observabilis Domini quando eduxit eos de terra Aegypti hanc observare debent omnes filii Israhel in generationibus suis
EXOD|12|43|dixitque Dominus ad Mosen et Aaron haec est religio phase omnis alienigena non comedet ex eo
EXOD|12|44|omnis autem servus empticius circumcidetur et sic comedet
EXOD|12|45|advena et mercennarius non edent ex eo
EXOD|12|46|in una domo comedetur nec efferetis de carnibus eius foras nec os illius confringetis
EXOD|12|47|omnis coetus filiorum Israhel faciet illud
EXOD|12|48|quod si quis peregrinorum in vestram voluerit transire coloniam et facere phase Domini circumcidetur prius omne masculinum eius et tunc rite celebrabit eritque sicut indigena terrae si quis autem circumcisus non fuerit non vescetur ex eo
EXOD|12|49|eadem lex erit indigenae et colono qui peregrinatur apud vos
EXOD|12|50|fecerunt omnes filii Israhel sicut praeceperat Dominus Mosi et Aaron
EXOD|12|51|et in eadem die eduxit Dominus filios Israhel de terra Aegypti per turmas suas
EXOD|13|1|locutusque est Dominus ad Mosen dicens
EXOD|13|2|sanctifica mihi omne primogenitum quod aperit vulvam in filiis Israhel tam de hominibus quam de iumentis mea sunt enim omnia
EXOD|13|3|et ait Moses ad populum mementote diei huius in qua egressi estis de Aegypto et de domo servitutis quoniam in manu forti eduxit vos Dominus de loco isto ut non comedatis fermentatum panem
EXOD|13|4|hodie egredimini mense novarum frugum
EXOD|13|5|cumque te introduxerit Dominus in terram Chananei et Hetthei et Amorrei et Evei et Iebusei quam iuravit patribus tuis ut daret tibi terram fluentem lacte et melle celebrabis hunc morem sacrorum mense isto
EXOD|13|6|septem diebus vesceris azymis et in die septimo erit sollemnitas Domini
EXOD|13|7|azyma comedetis septem diebus non apparebit apud te aliquid fermentatum nec in cunctis finibus tuis
EXOD|13|8|narrabisque filio tuo in die illo dicens hoc est quod fecit Dominus mihi quando egressus sum de Aegypto
EXOD|13|9|et erit quasi signum in manu tua et quasi monumentum ante oculos tuos et ut lex Domini semper in ore tuo in manu enim forti eduxit te Dominus de Aegypto
EXOD|13|10|custodies huiuscemodi cultum statuto tempore a diebus in dies
EXOD|13|11|cumque introduxerit te in terram Chananei sicut iuravit tibi et patribus tuis et dederit eam tibi
EXOD|13|12|separabis omne quod aperit vulvam Domino et quod primitivum est in pecoribus tuis quicquid habueris masculini sexus consecrabis Domino
EXOD|13|13|primogenitum asini mutabis ove quod si non redemeris interficies omne autem primogenitum hominis de filiis tuis pretio redimes
EXOD|13|14|cumque interrogaverit te filius tuus cras dicens quid est hoc respondebis ei in manu forti eduxit nos Dominus de Aegypto de domo servitutis
EXOD|13|15|nam cum induratus esset Pharao et nollet nos dimittere occidit Dominus omne primogenitum in terra Aegypti a primogenito hominis usque ad primogenitum iumentorum idcirco immolo Domino omne quod aperit vulvam masculini sexus et omnia primogenita filiorum meorum redimo
EXOD|13|16|erit igitur quasi signum in manu tua et quasi adpensum quid ob recordationem inter oculos tuos eo quod in manu forti eduxerit nos Dominus de Aegypto
EXOD|13|17|igitur cum emisisset Pharao populum non eos duxit Dominus per viam terrae Philisthim quae vicina est reputans ne forte paeniteret eum si vidisset adversum se bella consurgere et reverteretur in Aegyptum
EXOD|13|18|sed circumduxit per viam deserti quae est iuxta mare Rubrum et armati ascenderunt filii Israhel de terra Aegypti
EXOD|13|19|tulit quoque Moses ossa Ioseph secum eo quod adiurasset filios Israhel dicens visitabit vos Deus efferte ossa mea hinc vobiscum
EXOD|13|20|profectique de Soccoth castrametati sunt in Etham in extremis finibus solitudinis
EXOD|13|21|Dominus autem praecedebat eos ad ostendendam viam per diem in columna nubis et per noctem in columna ignis ut dux esset itineris utroque tempore
EXOD|13|22|numquam defuit columna nubis per diem nec columna ignis per noctem coram populo
EXOD|14|1|locutus est autem Dominus ad Mosen dicens
EXOD|14|2|loquere filiis Israhel reversi castrametentur e regione Phiahiroth quae est inter Magdolum et mare contra Beelsephon in conspectu eius castra ponetis super mare
EXOD|14|3|dicturusque est Pharao super filiis Israhel coartati sunt in terra conclusit eos desertum
EXOD|14|4|et indurabo cor eius ac persequetur vos et glorificabor in Pharao et in omni exercitu eius scientque Aegyptii quia ego sum Dominus feceruntque ita
EXOD|14|5|et nuntiatum est regi Aegyptiorum quod fugisset populus inmutatumque est cor Pharaonis et servorum eius super populo et dixerunt quid voluimus facere ut dimitteremus Israhel ne serviret nobis
EXOD|14|6|iunxit ergo currum et omnem populum suum adsumpsit secum
EXOD|14|7|tulitque sescentos currus electos quicquid in Aegypto curruum fuit et duces totius exercitus
EXOD|14|8|induravitque Dominus cor Pharaonis regis Aegypti et persecutus est filios Israhel at illi egressi erant in manu excelsa
EXOD|14|9|cumque persequerentur Aegyptii vestigia praecedentium reppererunt eos in castris super mare omnis equitatus et currus Pharaonis et universus exercitus erant in Ahiroth contra Beelsephon
EXOD|14|10|cumque adpropinquasset Pharao levantes filii Israhel oculos viderunt Aegyptios post se et timuerunt valde clamaveruntque ad Dominum
EXOD|14|11|et dixerunt ad Mosen forsitan non erant sepulchra in Aegypto ideo tulisti nos ut moreremur in solitudine quid hoc facere voluisti ut educeres nos ex Aegypto
EXOD|14|12|nonne iste est sermo quem loquebamur ad te in Aegypto dicentes recede a nobis ut serviamus Aegyptiis multo enim melius est servire eis quam mori in solitudine
EXOD|14|13|et ait Moses ad populum nolite timere state et videte magnalia Domini quae facturus est hodie Aegyptios enim quos nunc videtis nequaquam ultra videbitis usque in sempiternum
EXOD|14|14|Dominus pugnabit pro vobis et vos tacebitis
EXOD|14|15|dixitque Dominus ad Mosen quid clamas ad me loquere filiis Israhel ut proficiscantur
EXOD|14|16|tu autem eleva virgam tuam et extende manum super mare et divide illud ut gradiantur filii Israhel in medio mari per siccum
EXOD|14|17|ego autem indurabo cor Aegyptiorum ut persequantur vos et glorificabor in Pharaone et in omni exercitu eius in curribus et in equitibus illius
EXOD|14|18|et scient Aegyptii quia ego sum Dominus cum glorificatus fuero in Pharaone et in curribus atque in equitibus eius
EXOD|14|19|tollensque se angelus Dei qui praecedebat castra Israhel abiit post eos et cum eo pariter columna nubis priora dimittens post tergum
EXOD|14|20|stetit inter castra Aegyptiorum et castra Israhel et erat nubes tenebrosa et inluminans noctem ut ad se invicem toto noctis tempore accedere non valerent
EXOD|14|21|cumque extendisset Moses manum super mare abstulit illud Dominus flante vento vehementi et urente tota nocte et vertit in siccum divisaque est aqua
EXOD|14|22|et ingressi sunt filii Israhel per medium maris sicci erat enim aqua quasi murus a dextra eorum et leva
EXOD|14|23|persequentesque Aegyptii ingressi sunt post eos omnis equitatus Pharaonis currus eius et equites per medium maris
EXOD|14|24|iamque advenerat vigilia matutina et ecce respiciens Dominus super castra Aegyptiorum per columnam ignis et nubis interfecit exercitum eorum
EXOD|14|25|et subvertit rotas curruum ferebanturque in profundum dixerunt ergo Aegyptii fugiamus Israhelem Dominus enim pugnat pro eis contra nos
EXOD|14|26|et ait Dominus ad Mosen extende manum tuam super mare ut revertantur aquae ad Aegyptios super currus et equites eorum
EXOD|14|27|cumque extendisset Moses manum contra mare reversum est primo diluculo ad priorem locum fugientibusque Aegyptiis occurrerunt aquae et involvit eos Dominus in mediis fluctibus
EXOD|14|28|reversaeque sunt aquae et operuerunt currus et equites cuncti exercitus Pharaonis qui sequentes ingressi fuerant mare ne unus quidem superfuit ex eis
EXOD|14|29|filii autem Israhel perrexerunt per medium sicci maris et aquae eis erant quasi pro muro a dextris et a sinistris
EXOD|14|30|liberavitque Dominus in die illo Israhel de manu Aegyptiorum
EXOD|14|31|et viderunt Aegyptios mortuos super litus maris et manum magnam quam exercuerat Dominus contra eos timuitque populus Dominum et crediderunt Domino et Mosi servo eius
EXOD|15|1|tunc cecinit Moses et filii Israhel carmen hoc Domino et dixerunt cantemus Domino gloriose enim magnificatus est equum et ascensorem deiecit in mare
EXOD|15|2|fortitudo mea et laus mea Dominus et factus est mihi in salutem iste Deus meus et glorificabo eum Deus patris mei et exaltabo eum
EXOD|15|3|Dominus quasi vir pugnator Omnipotens nomen eius
EXOD|15|4|currus Pharaonis et exercitum eius proiecit in mare electi principes eius submersi sunt in mari Rubro
EXOD|15|5|abyssi operuerunt eos descenderunt in profundum quasi lapis
EXOD|15|6|dextera tua Domine magnifice in fortitudine dextera tua Domine percussit inimicum
EXOD|15|7|et in multitudine gloriae tuae deposuisti adversarios meos misisti iram tuam quae devoravit eos ut stipulam
EXOD|15|8|et in spiritu furoris tui congregatae sunt aquae stetit unda fluens congregatae sunt abyssi in medio mari
EXOD|15|9|dixit inimicus persequar et conprehendam dividam spolia implebitur anima mea evaginabo gladium meum interficiet eos manus mea
EXOD|15|10|flavit spiritus tuus et operuit eos mare submersi sunt quasi plumbum in aquis vehementibus
EXOD|15|11|quis similis tui in fortibus Domine quis similis tui magnificus in sanctitate terribilis atque laudabilis et faciens mirabilia
EXOD|15|12|extendisti manum tuam et devoravit eos terra
EXOD|15|13|dux fuisti in misericordia tua populo quem redemisti et portasti eum in fortitudine tua ad habitaculum sanctum tuum
EXOD|15|14|adtenderunt populi et irati sunt dolores obtinuerunt habitatores Philisthim
EXOD|15|15|tunc conturbati sunt principes Edom robustos Moab obtinuit tremor obriguerunt omnes habitatores Chanaan
EXOD|15|16|inruat super eos formido et pavor in magnitudine brachii tui fiant inmobiles quasi lapis donec pertranseat populus tuus Domine donec pertranseat populus tuus iste quem possedisti
EXOD|15|17|introduces eos et plantabis in monte hereditatis tuae firmissimo habitaculo tuo quod operatus es Domine sanctuarium Domine quod firmaverunt manus tuae
EXOD|15|18|Dominus regnabit in aeternum et ultra
EXOD|15|19|ingressus est enim equus Pharao cum curribus et equitibus eius in mare et reduxit super eos Dominus aquas maris filii autem Israhel ambulaverunt per siccum in medio eius
EXOD|15|20|sumpsit ergo Maria prophetis soror Aaron tympanum in manu egressaeque sunt omnes mulieres post eam cum tympanis et choris
EXOD|15|21|quibus praecinebat dicens cantemus Domino gloriose enim magnificatus est equum et ascensorem eius deiecit in mare
EXOD|15|22|tulit autem Moses Israhel de mari Rubro et egressi sunt in desertum Sur ambulaveruntque tribus diebus per solitudinem et non inveniebant aquam
EXOD|15|23|et venerunt in Marath nec poterant bibere aquas de Mara eo quod essent amarae unde et congruum loco nomen inposuit vocans illud Mara id est amaritudinem
EXOD|15|24|et murmuravit populus contra Mosen dicens quid bibemus
EXOD|15|25|at ille clamavit ad Dominum qui ostendit ei lignum quod cum misisset in aquas in dulcedinem versae sunt ibi constituit ei praecepta atque iudicia et ibi temptavit eum
EXOD|15|26|dicens si audieris vocem Domini Dei tui et quod rectum est coram eo feceris et oboedieris mandatis eius custodierisque omnia praecepta illius cunctum languorem quem posui in Aegypto non inducam super te ego enim Dominus sanator tuus
EXOD|15|27|venerunt autem in Helim ubi erant duodecim fontes aquarum et septuaginta palmae et castrametati sunt iuxta aquas
EXOD|16|1|profectique sunt de Helim et venit omnis multitudo filiorum Israhel in desertum Sin quod est inter Helim et Sinai quintodecimo die mensis secundi postquam egressi sunt de terra Aegypti
EXOD|16|2|et murmuravit omnis congregatio filiorum Israhel contra Mosen et contra Aaron in solitudine
EXOD|16|3|dixeruntque ad eos filii Israhel utinam mortui essemus per manum Domini in terra Aegypti quando sedebamus super ollas carnium et comedebamus panes in saturitate cur eduxistis nos in desertum istud ut occideretis omnem multitudinem fame
EXOD|16|4|dixit autem Dominus ad Mosen ecce ego pluam vobis panes de caelo egrediatur populus et colligat quae sufficiunt per singulos dies ut temptem eum utrum ambulet in lege mea an non
EXOD|16|5|die autem sexta parent quod inferant et sit duplum quam colligere solebant per singulos dies
EXOD|16|6|dixeruntque Moses et Aaron ad omnes filios Israhel vespere scietis quod Dominus eduxerit vos de terra Aegypti
EXOD|16|7|et mane videbitis gloriam Domini audivit enim murmur vestrum contra Dominum nos vero quid sumus quia mussitatis contra nos
EXOD|16|8|et ait Moses dabit Dominus vobis vespere carnes edere et mane panes in saturitate eo quod audierit murmurationes vestras quibus murmurati estis contra eum nos enim quid sumus nec contra nos est murmur vestrum sed contra Dominum
EXOD|16|9|dixitque Moses ad Aaron dic universae congregationi filiorum Israhel accedite coram Domino audivit enim murmur vestrum
EXOD|16|10|cumque loqueretur Aaron ad omnem coetum filiorum Israhel respexerunt ad solitudinem et ecce gloria Domini apparuit in nube
EXOD|16|11|locutus est autem Dominus ad Mosen dicens
EXOD|16|12|audivi murmurationes filiorum Israhel loquere ad eos vespere comedetis carnes et mane saturabimini panibus scietisque quod sim Dominus Deus vester
EXOD|16|13|factum est ergo vespere et ascendens coturnix operuit castra mane quoque ros iacuit per circuitum castrorum
EXOD|16|14|cumque operuisset superficiem terrae apparuit in solitudine minutum et quasi pilo tunsum in similitudinem pruinae super terram
EXOD|16|15|quod cum vidissent filii Israhel dixerunt ad invicem man hu quod significat quid est hoc ignorabant enim quid esset quibus ait Moses iste est panis quem dedit Dominus vobis ad vescendum
EXOD|16|16|hic est sermo quem praecepit Dominus colligat ex eo unusquisque quantum sufficiat ad vescendum gomor per singula capita iuxta numerum animarum vestrarum quae habitant in tabernaculo sic tolletis
EXOD|16|17|feceruntque ita filii Israhel et collegerunt alius plus alius minus
EXOD|16|18|et mensi sunt ad mensuram gomor nec qui plus collegerat habuit amplius nec qui minus paraverat repperit minus sed singuli iuxta id quod edere poterant congregarunt
EXOD|16|19|dixitque Moses ad eos nullus relinquat ex eo in mane
EXOD|16|20|qui non audierunt eum sed dimiserunt quidam ex eis usque mane et scatere coepit vermibus atque conputruit et iratus est contra eos Moses
EXOD|16|21|colligebant autem mane singuli quantum sufficere poterat ad vescendum cumque incaluisset sol liquefiebat
EXOD|16|22|in die vero sexta collegerunt cibos duplices id est duo gomor per singulos homines venerunt autem omnes principes multitudinis et narraverunt Mosi
EXOD|16|23|qui ait eis hoc est quod locutus est Dominus requies sabbati sanctificata erit Domino cras quodcumque operandum est facite et quae coquenda sunt coquite quicquid autem reliquum fuerit reponite usque in mane
EXOD|16|24|feceruntque ita ut praeceperat Moses et non conputruit neque vermis inventus est in eo
EXOD|16|25|dixitque Moses comedite illud hodie quia sabbatum est Domino non invenietur hodie in agro
EXOD|16|26|sex diebus colligite in die autem septimo sabbatum est Domino idcirco non invenietur
EXOD|16|27|venit septima dies et egressi de populo ut colligerent non invenerunt
EXOD|16|28|dixit autem Dominus ad Mosen usquequo non vultis custodire mandata mea et legem meam
EXOD|16|29|videte quod Dominus dederit vobis sabbatum et propter hoc tribuerit vobis die sexto cibos duplices maneat unusquisque apud semet ipsum nullus egrediatur de loco suo die septimo
EXOD|16|30|et sabbatizavit populus die septimo
EXOD|16|31|appellavitque domus Israhel nomen eius man quod erat quasi semen coriandri album gustusque eius quasi similae cum melle
EXOD|16|32|dixit autem Moses iste est sermo quem praecepit Dominus imple gomor ex eo et custodiatur in futuras retro generationes ut noverint panem quo alui vos in solitudine quando educti estis de terra Aegypti
EXOD|16|33|dixitque Moses ad Aaron sume vas unum et mitte ibi man quantum potest capere gomor et repone coram Domino ad servandum in generationes vestras
EXOD|16|34|sicut praecepit Dominus Mosi posuitque illud Aaron in tabernaculo reservandum
EXOD|16|35|filii autem Israhel comederunt man quadraginta annis donec venirent in terram habitabilem hoc cibo aliti sunt usquequo tangerent fines terrae Chanaan
EXOD|16|36|gomor autem decima pars est oephi
EXOD|17|1|igitur profecta omnis multitudo filiorum Israhel de deserto Sin per mansiones suas iuxta sermonem Domini castrametata est in Raphidim ubi non erat aqua ad bibendum populo
EXOD|17|2|qui iurgatus contra Mosen ait da nobis aquam ut bibamus quibus respondit Moses quid iurgamini contra me cur temptatis Dominum
EXOD|17|3|sitivit ergo populus ibi pro aquae penuria et murmuravit contra Mosen dicens cur nos exire fecisti de Aegypto ut occideres et nos et liberos nostros ac iumenta siti
EXOD|17|4|clamavit autem Moses ad Dominum dicens quid faciam populo huic adhuc pauxillum et lapidabunt me
EXOD|17|5|ait Dominus ad Mosen antecede populum et sume tecum de senibus Israhel et virgam qua percussisti fluvium tolle in manu tua et vade
EXOD|17|6|en ego stabo coram te ibi super petram Horeb percutiesque petram et exibit ex ea aqua ut bibat populus fecit Moses ita coram senibus Israhel
EXOD|17|7|et vocavit nomen loci illius Temptatio propter iurgium filiorum Israhel et quia temptaverunt Dominum dicentes estne Dominus in nobis an non
EXOD|17|8|venit autem Amalech et pugnabat contra Israhel in Raphidim
EXOD|17|9|dixitque Moses ad Iosue elige viros et egressus pugna contra Amalech cras ego stabo in vertice collis habens virgam Dei in manu mea
EXOD|17|10|fecit Iosue ut locutus ei erat Moses et pugnavit contra Amalech Moses autem et Aaron et Hur ascenderunt super verticem collis
EXOD|17|11|cumque levaret Moses manus vincebat Israhel sin autem paululum remisisset superabat Amalech
EXOD|17|12|manus autem Mosi erant graves sumentes igitur lapidem posuerunt subter eum in quo sedit Aaron autem et Hur sustentabant manus eius ex utraque parte et factum est ut manus ipsius non lassarentur usque ad occasum solis
EXOD|17|13|fugavitque Iosue Amalech et populum eius in ore gladii
EXOD|17|14|dixit autem Dominus ad Mosen scribe hoc ob monumentum in libro et trade auribus Iosue delebo enim memoriam Amalech sub caelo
EXOD|17|15|aedificavitque Moses altare et vocavit nomen eius Dominus exaltatio mea dicens
EXOD|17|16|quia manus solii Domini et bellum Dei erit contra Amalech a generatione in generationem
EXOD|18|1|cumque audisset Iethro sacerdos Madian cognatus Mosi omnia quae fecerat Deus Mosi et Israhel populo suo eo quod eduxisset Dominus Israhel de Aegypto
EXOD|18|2|tulit Sefforam uxorem Mosi quam remiserat
EXOD|18|3|et duos filios eius quorum unus vocabatur Gersan dicente patre advena fui in terra aliena
EXOD|18|4|alter vero Eliezer Deus enim ait patris mei adiutor meus et eruit me de gladio Pharaonis
EXOD|18|5|venit ergo Iethro cognatus Mosi et filii eius et uxor ad Mosen in desertum ubi erat castrametatus iuxta montem Dei
EXOD|18|6|et mandavit Mosi dicens ego cognatus tuus Iethro venio ad te et uxor tua et duo filii tui cum ea
EXOD|18|7|qui egressus in occursum cognati sui adoravit et osculatus est eum salutaveruntque se mutuo verbis pacificis cumque intrasset tabernaculum
EXOD|18|8|narravit Moses cognato suo cuncta quae fecerat Deus Pharaoni et Aegyptiis propter Israhel universum laborem qui accidisset eis in itinere quo liberarat eos Dominus
EXOD|18|9|laetatusque est Iethro super omnibus bonis quae fecerat Dominus Israheli eo quod eruisset eum de manu Aegyptiorum
EXOD|18|10|et ait benedictus Dominus qui liberavit vos de manu Aegyptiorum et de manu Pharaonis qui eruit populum suum de manu Aegypti
EXOD|18|11|nunc cognovi quia magnus Dominus super omnes deos eo quod superbe egerint contra illos
EXOD|18|12|obtulit ergo Iethro cognatus Mosi holocausta et hostias Deo veneruntque Aaron et omnes senes Israhel ut comederent panem cum eo coram Domino
EXOD|18|13|altero autem die sedit Moses ut iudicaret populum qui adsistebat Mosi de mane usque ad vesperam
EXOD|18|14|quod cum vidisset cognatus eius omnia scilicet quae agebat in populo ait quid est hoc quod facis in plebe cur solus sedes et omnis populus praestolatur de mane usque ad vesperam
EXOD|18|15|cui respondit Moses venit ad me populus quaerens sententiam Dei
EXOD|18|16|cumque acciderit eis aliqua disceptatio veniunt ad me ut iudicem inter eos et ostendam praecepta Dei et leges eius
EXOD|18|17|at ille non bonam inquit rem facis
EXOD|18|18|stulto labore consumeris et tu et populus iste qui tecum est ultra vires tuas est negotium solus illud non poteris sustinere
EXOD|18|19|sed audi verba mea atque consilia et erit Deus tecum esto tu populo in his quae ad Deum pertinent ut referas quae dicuntur ad eum
EXOD|18|20|ostendasque populo caerimonias et ritum colendi viamque per quam ingredi debeant et opus quod facere
EXOD|18|21|provide autem de omni plebe viros potentes et timentes Deum in quibus sit veritas et qui oderint avaritiam et constitue ex eis tribunos et centuriones et quinquagenarios et decanos
EXOD|18|22|qui iudicent populum omni tempore quicquid autem maius fuerit referant ad te et ipsi minora tantummodo iudicent leviusque tibi sit partito in alios onere
EXOD|18|23|si hoc feceris implebis imperium Dei et praecepta eius poteris sustentare et omnis hic populus revertetur cum pace ad loca sua
EXOD|18|24|quibus auditis Moses fecit omnia quae ille suggesserat
EXOD|18|25|et electis viris strenuis de cuncto Israhel constituit eos principes populi tribunos et centuriones et quinquagenarios et decanos
EXOD|18|26|qui iudicabant plebem omni tempore quicquid autem gravius erat referebant ad eum faciliora tantummodo iudicantes
EXOD|18|27|dimisitque cognatum qui reversus abiit in terram suam
EXOD|19|1|mense tertio egressionis Israhel de terra Aegypti in die hac venerunt in solitudinem Sinai
EXOD|19|2|nam profecti de Raphidim et pervenientes usque in desertum Sinai castrametati sunt in eodem loco ibique Israhel fixit tentoria e regione montis
EXOD|19|3|Moses autem ascendit ad Deum vocavitque eum Dominus de monte et ait haec dices domui Iacob et adnuntiabis filiis Israhel
EXOD|19|4|vos ipsi vidistis quae fecerim Aegyptiis quomodo portaverim vos super alas aquilarum et adsumpserim mihi
EXOD|19|5|si ergo audieritis vocem meam et custodieritis pactum meum eritis mihi in peculium de cunctis populis mea est enim omnis terra
EXOD|19|6|et vos eritis mihi regnum sacerdotale et gens sancta haec sunt verba quae loqueris ad filios Israhel
EXOD|19|7|venit Moses et convocatis maioribus natu populi exposuit omnes sermones quos mandaverat Dominus
EXOD|19|8|responditque universus populus simul cuncta quae locutus est Dominus faciemus cumque rettulisset Moses verba populi ad Dominum
EXOD|19|9|ait ei Dominus iam nunc veniam ad te in caligine nubis ut audiat me populus loquentem ad te et credat tibi in perpetuum nuntiavit ergo Moses verba populi ad Dominum
EXOD|19|10|qui dixit ei vade ad populum et sanctifica illos hodie et cras laventque vestimenta sua
EXOD|19|11|et sint parati in diem tertium die enim tertio descendet Dominus coram omni plebe super montem Sinai
EXOD|19|12|constituesque terminos populo per circuitum et dices cavete ne ascendatis in montem nec tangatis fines illius omnis qui tetigerit montem morte morietur
EXOD|19|13|manus non tanget eum sed lapidibus opprimetur aut confodietur iaculis sive iumentum fuerit sive homo non vivet cum coeperit clangere bucina tunc ascendant in montem
EXOD|19|14|descenditque Moses de monte ad populum et sanctificavit eum cumque lavissent vestimenta sua
EXOD|19|15|ait ad eos estote parati in diem tertium ne adpropinquetis uxoribus vestris
EXOD|19|16|iam advenerat tertius dies et mane inclaruerat et ecce coeperunt audiri tonitrua ac micare fulgura et nubes densissima operire montem clangorque bucinae vehementius perstrepebat timuit populus qui erat in castris
EXOD|19|17|cumque eduxisset eos Moses in occursum Dei de loco castrorum steterunt ad radices montis
EXOD|19|18|totus autem mons Sinai fumabat eo quod descendisset Dominus super eum in igne et ascenderet fumus ex eo quasi de fornace eratque mons omnis terribilis
EXOD|19|19|et sonitus bucinae paulatim crescebat in maius et prolixius tendebatur Moses loquebatur et Dominus respondebat ei
EXOD|19|20|descenditque Dominus super montem Sinai in ipso montis vertice et vocavit Mosen in cacumen eius quo cum ascendisset
EXOD|19|21|dixit ad eum descende et contestare populum ne forte velint transcendere terminos ad videndum Dominum et pereat ex eis plurima multitudo
EXOD|19|22|sacerdotes quoque qui accedunt ad Dominum sanctificentur ne percutiat eos
EXOD|19|23|dixitque Moses ad Dominum non poterit vulgus ascendere in montem Sinai tu enim testificatus es et iussisti dicens pone terminos circa montem et sanctifica illum
EXOD|19|24|cui ait Dominus vade descende ascendesque tu et Aaron tecum sacerdotes autem et populus ne transeant terminos nec ascendant ad Dominum ne forte interficiat illos
EXOD|19|25|descendit Moses ad populum et omnia narravit eis
EXOD|20|1|locutus quoque est Dominus cunctos sermones hos
EXOD|20|2|ego sum Dominus Deus tuus qui eduxi te de terra Aegypti de domo servitutis
EXOD|20|3|non habebis deos alienos coram me
EXOD|20|4|non facies tibi sculptile neque omnem similitudinem quae est in caelo desuper et quae in terra deorsum nec eorum quae sunt in aquis sub terra
EXOD|20|5|non adorabis ea neque coles ego sum Dominus Deus tuus fortis zelotes visitans iniquitatem patrum in filiis in tertiam et quartam generationem eorum qui oderunt me
EXOD|20|6|et faciens misericordiam in milia his qui diligunt me et custodiunt praecepta mea
EXOD|20|7|non adsumes nomen Domini Dei tui in vanum nec enim habebit insontem Dominus eum qui adsumpserit nomen Domini Dei sui frustra
EXOD|20|8|memento ut diem sabbati sanctifices
EXOD|20|9|sex diebus operaberis et facies omnia opera tua
EXOD|20|10|septimo autem die sabbati Domini Dei tui non facies omne opus tu et filius tuus et filia tua servus tuus et ancilla tua iumentum tuum et advena qui est intra portas tuas
EXOD|20|11|sex enim diebus fecit Dominus caelum et terram et mare et omnia quae in eis sunt et requievit in die septimo idcirco benedixit Dominus diei sabbati et sanctificavit eum
EXOD|20|12|honora patrem tuum et matrem tuam ut sis longevus super terram quam Dominus Deus tuus dabit tibi
EXOD|20|13|non occides
EXOD|20|14|non moechaberis
EXOD|20|15|non furtum facies
EXOD|20|16|non loqueris contra proximum tuum falsum testimonium
EXOD|20|17|non concupisces domum proximi tui nec desiderabis uxorem eius non servum non ancillam non bovem non asinum nec omnia quae illius sunt
EXOD|20|18|cunctus autem populus videbat voces et lampadas et sonitum bucinae montemque fumantem et perterriti ac pavore concussi steterunt procul
EXOD|20|19|dicentes Mosi loquere tu nobis et audiemus non loquatur nobis Dominus ne forte moriamur
EXOD|20|20|et ait Moses ad populum nolite timere ut enim probaret vos venit Deus et ut terror illius esset in vobis et non peccaretis
EXOD|20|21|stetitque populus de longe Moses autem accessit ad caliginem in qua erat Deus
EXOD|20|22|dixit praeterea Dominus ad Mosen haec dices filiis Israhel vos vidistis quod de caelo locutus sum vobis
EXOD|20|23|non facietis mecum deos argenteos nec deos aureos facietis vobis
EXOD|20|24|altare de terra facietis mihi et offeretis super eo holocausta et pacifica vestra oves vestras et boves in omni loco in quo memoria fuerit nominis mei veniam ad te et benedicam tibi
EXOD|20|25|quod si altare lapideum feceris mihi non aedificabis illud de sectis lapidibus si enim levaveris cultrum tuum super eo polluetur
EXOD|20|26|non ascendes per gradus ad altare meum ne reveletur turpitudo tua
EXOD|21|1|haec sunt iudicia quae propones eis
EXOD|21|2|si emeris servum hebraeum sex annis serviet tibi in septimo egredietur liber gratis
EXOD|21|3|cum quali veste intraverit cum tali exeat si habens uxorem et uxor egredietur simul
EXOD|21|4|sin autem dominus dederit illi uxorem et peperit filios et filias mulier et liberi eius erunt domini sui ipse vero exibit cum vestitu suo
EXOD|21|5|quod si dixerit servus diligo dominum meum et uxorem ac liberos non egrediar liber
EXOD|21|6|offeret eum dominus diis et adplicabitur ad ostium et postes perforabitque aurem eius subula et erit ei servus in saeculum
EXOD|21|7|si quis vendiderit filiam suam in famulam non egredietur sicut ancillae exire consuerunt
EXOD|21|8|si displicuerit oculis domini sui cui tradita fuerit dimittet eam populo autem alieno vendendi non habet potestatem si spreverit eam
EXOD|21|9|sin autem filio suo desponderit eam iuxta morem filiarum faciet illi
EXOD|21|10|quod si alteram ei acceperit providebit puellae nuptias et vestimenta et pretium pudicitiae non negabit
EXOD|21|11|si tria ista non fecerit egredietur gratis absque pecunia
EXOD|21|12|qui percusserit hominem volens occidere morte moriatur
EXOD|21|13|qui autem non est insidiatus sed Deus illum tradidit in manu eius constituam tibi locum quo fugere debeat
EXOD|21|14|si quis de industria occiderit proximum suum et per insidias ab altari meo evelles eum ut moriatur
EXOD|21|15|qui percusserit patrem suum et matrem morte moriatur
EXOD|21|16|qui furatus fuerit hominem et vendiderit eum convictus noxae morte moriatur
EXOD|21|17|qui maledixerit patri suo et matri morte moriatur
EXOD|21|18|si rixati fuerint viri et percusserit alter proximum suum lapide vel pugno et ille mortuus non fuerit sed iacuerit in lectulo
EXOD|21|19|si surrexerit et ambulaverit foris super baculum suum innocens erit qui percussit ita tamen ut operas eius et inpensas in medicos restituat
EXOD|21|20|qui percusserit servum suum vel ancillam virga et mortui fuerint in manibus eius criminis reus erit
EXOD|21|21|sin autem uno die supervixerit vel duobus non subiacebit poenae quia pecunia illius est
EXOD|21|22|si rixati fuerint viri et percusserit quis mulierem praegnantem et abortivum quidem fecerit sed ipsa vixerit subiacebit damno quantum expetierit maritus mulieris et arbitri iudicarint
EXOD|21|23|sin autem mors eius fuerit subsecuta reddet animam pro anima
EXOD|21|24|oculum pro oculo dentem pro dente manum pro manu pedem pro pede
EXOD|21|25|adustionem pro adustione vulnus pro vulnere livorem pro livore
EXOD|21|26|si percusserit quispiam oculum servi sui aut ancillae et luscos eos fecerit dimittet liberos pro oculo quem eruit
EXOD|21|27|dentem quoque si excusserit servo vel ancillae suae similiter dimittet eos liberos
EXOD|21|28|si bos cornu petierit virum aut mulierem et mortui fuerint lapidibus obruetur et non comedentur carnes eius dominusque bovis innocens erit
EXOD|21|29|quod si bos cornipeta fuerit ab heri et nudius tertius et contestati sunt dominum eius nec reclusit eum occideritque virum aut mulierem et bos lapidibus obruetur et dominum illius occident
EXOD|21|30|quod si pretium ei fuerit inpositum dabit pro anima sua quicquid fuerit postulatus
EXOD|21|31|filium quoque et filiam si cornu percusserit simili sententiae subiacebit
EXOD|21|32|si servum ancillamque invaserit triginta siclos argenti dabit domino bos vero lapidibus opprimetur
EXOD|21|33|si quis aperuerit cisternam et foderit et non operuerit eam cecideritque bos vel asinus in eam
EXOD|21|34|dominus cisternae reddet pretium iumentorum quod autem mortuum est ipsius erit
EXOD|21|35|si bos alienus bovem alterius vulnerarit et ille mortuus fuerit vendent bovem vivum et divident pretium cadaver autem mortui inter se dispertient
EXOD|21|36|sin autem sciebat quod bos cornipeta esset ab heri et nudius tertius et non custodivit eum dominus suus reddet bovem pro bove et cadaver integrum accipiet
EXOD|22|1|si quis furatus fuerit bovem aut ovem et occiderit vel vendiderit quinque boves pro uno bove restituet et quattuor oves pro una ove
EXOD|22|2|si effringens fur domum sive suffodiens fuerit inventus et accepto vulnere mortuus fuerit percussor non erit reus sanguinis
EXOD|22|3|quod si orto sole hoc fecerit homicidium perpetravit et ipse morietur si non habuerit quod pro furto reddat venundabitur
EXOD|22|4|si inventum fuerit apud eum quod furatus est vivens sive bos sive asinus sive ovis duplum restituet
EXOD|22|5|si laeserit quispiam agrum vel vineam et dimiserit iumentum suum ut depascatur aliena quicquid optimum habuerit in agro suo vel in vinea pro damni aestimatione restituet
EXOD|22|6|si egressus ignis invenerit spinas et conprehenderit acervos frugum sive stantes segetes in agris reddet damnum qui ignem succenderit
EXOD|22|7|si quis commendaverit amico pecuniam aut vas in custodiam et ab eo qui susceperat furto ablata fuerint si invenitur fur duplum reddet
EXOD|22|8|si latet dominus domus adplicabitur ad deos et iurabit quod non extenderit manum in rem proximi sui
EXOD|22|9|ad perpetrandam fraudem tam in bove quam in asino et ove ac vestimento et quicquid damnum inferre potest ad deos utriusque causa perveniet et si illi iudicaverint duplum restituet proximo suo
EXOD|22|10|si quis commendaverit proximo suo asinum bovem ovem et omne iumentum ad custodiam et mortuum fuerit aut debilitatum vel captum ab hostibus nullusque hoc viderit
EXOD|22|11|iusiurandum erit in medio quod non extenderit manum ad rem proximi sui suscipietque dominus iuramentum et ille reddere non cogetur
EXOD|22|12|quod si furto ablatum fuerit restituet damnum domino
EXOD|22|13|si comestum a bestia deferet ad eum quod occisum est et non restituet
EXOD|22|14|qui a proximo suo quicquam horum mutuo postularit et debilitatum aut mortuum fuerit domino non praesente reddere conpelletur
EXOD|22|15|quod si inpraesentiarum fuit dominus non restituet maxime si conductum venerat pro mercede operis sui
EXOD|22|16|si seduxerit quis virginem necdum desponsatam et dormierit cum ea dotabit eam et habebit uxorem
EXOD|22|17|si pater virginis dare noluerit reddet pecuniam iuxta modum dotis quam virgines accipere consuerunt
EXOD|22|18|maleficos non patieris vivere
EXOD|22|19|qui coierit cum iumento morte moriatur
EXOD|22|20|qui immolat diis occidetur praeter Domino soli
EXOD|22|21|advenam non contristabis neque adfliges eum advenae enim et ipsi fuistis in terra Aegypti
EXOD|22|22|viduae et pupillo non nocebitis
EXOD|22|23|si laeseritis eos vociferabuntur ad me et ego audiam clamorem eorum
EXOD|22|24|et indignabitur furor meus percutiamque vos gladio et erunt uxores vestrae viduae et filii vestri pupilli
EXOD|22|25|si pecuniam mutuam dederis populo meo pauperi qui habitat tecum non urgues eum quasi exactor nec usuris opprimes
EXOD|22|26|si pignus a proximo tuo acceperis vestimentum ante solis occasum redde ei
EXOD|22|27|ipsum enim est solum quo operitur indumentum carnis eius nec habet aliud in quo dormiat si clamaverit ad me exaudiam eum quia misericors sum
EXOD|22|28|diis non detrahes et principi populi tui non maledices
EXOD|22|29|decimas tuas et primitias non tardabis offerre primogenitum filiorum tuorum dabis mihi
EXOD|22|30|de bubus quoque et ovibus similiter facies septem diebus sit cum matre sua die octavo reddes illum mihi
EXOD|22|31|viri sancti eritis mihi carnem quae a bestiis fuerit praegustata non comedetis sed proicietis canibus
EXOD|23|1|non suscipies vocem mendacii nec iunges manum tuam ut pro impio dicas falsum testimonium
EXOD|23|2|non sequeris turbam ad faciendum malum nec in iudicio plurimorum adquiesces sententiae ut a vero devies
EXOD|23|3|pauperis quoque non misereberis in negotio
EXOD|23|4|si occurreris bovi inimici tui aut asino erranti reduc ad eum
EXOD|23|5|si videris asinum odientis te iacere sub onere non pertransibis sed sublevabis cum eo
EXOD|23|6|non declinabis in iudicio pauperis
EXOD|23|7|mendacium fugies insontem et iustum non occides quia aversor impium
EXOD|23|8|nec accipias munera quae excaecant etiam prudentes et subvertunt verba iustorum
EXOD|23|9|peregrino molestus non eris scitis enim advenarum animas quia et ipsi peregrini fuistis in terra Aegypti
EXOD|23|10|sex annis seminabis terram tuam et congregabis fruges eius
EXOD|23|11|anno autem septimo dimittes eam et requiescere facies ut comedant pauperes populi tui et quicquid reliqui fuerit edant bestiae agri ita facies in vinea et in oliveto tuo
EXOD|23|12|sex diebus operaberis septima die cessabis ut requiescat bos et asinus tuus et refrigeretur filius ancillae tuae et advena
EXOD|23|13|omnia quae dixi vobis custodite et per nomen externorum deorum non iurabitis neque audietur ex ore vestro
EXOD|23|14|tribus vicibus per singulos annos mihi festa celebrabitis
EXOD|23|15|sollemnitatem azymorum custodies septem diebus comedes azyma sicut praecepi tibi tempore mensis novorum quando egressus es de Aegypto non apparebis in conspectu meo vacuus
EXOD|23|16|et sollemnitatem messis primitivorum operis tui quaecumque serueris in agro sollemnitatem quoque in exitu anni quando congregaveris omnes fruges tuas de agro
EXOD|23|17|ter in anno apparebit omne masculinum tuum coram Domino Deo
EXOD|23|18|non immolabis super fermento sanguinem victimae meae nec remanebit adeps sollemnitatis meae usque mane
EXOD|23|19|primitias frugum terrae tuae deferes in domum Domini Dei tui nec coques hedum in lacte matris suae
EXOD|23|20|ecce ego mittam angelum meum qui praecedat te et custodiat in via et introducat ad locum quem paravi
EXOD|23|21|observa eum et audi vocem eius nec contemnendum putes quia non dimittet cum peccaveritis et est nomen meum in illo
EXOD|23|22|quod si audieris vocem eius et feceris omnia quae loquor inimicus ero inimicis tuis et adfligam adfligentes te
EXOD|23|23|praecedetque te angelus meus et introducet te ad Amorreum et Hettheum et Ferezeum Chananeumque et Eveum et Iebuseum quos ego contribo
EXOD|23|24|non adorabis deos eorum nec coles eos non facies opera eorum sed destrues eos et confringes statuas eorum
EXOD|23|25|servietisque Domino Deo vestro ut benedicam panibus tuis et aquis et auferam infirmitatem de medio tui
EXOD|23|26|non erit infecunda nec sterilis in terra tua numerum dierum tuorum implebo
EXOD|23|27|terrorem meum mittam in praecursum tuum et occidam omnem populum ad quem ingredieris cunctorumque inimicorum tuorum coram te terga vertam
EXOD|23|28|emittens crabrones prius qui fugabunt Eveum et Chananeum et Hettheum antequam introeas
EXOD|23|29|non eiciam eos a facie tua anno uno ne terra in solitudinem redigatur et crescant contra te bestiae
EXOD|23|30|paulatim expellam eos de conspectu tuo donec augearis et possideas terram
EXOD|23|31|ponam autem terminos tuos a mari Rubro usque ad mare Palestinorum et a deserto usque ad Fluvium tradam manibus vestris habitatores terrae et eiciam eos de conspectu vestro
EXOD|23|32|non inibis cum eis foedus nec cum diis eorum
EXOD|23|33|non habitent in terra tua ne forte peccare te faciant in me si servieris diis eorum quod tibi certo erit in scandalum
EXOD|24|1|Mosi quoque dixit ascende ad Dominum tu et Aaron Nadab et Abiu et septuaginta senes ex Israhel et adorabitis procul
EXOD|24|2|solusque Moses ascendet ad Dominum et illi non adpropinquabunt nec populus ascendet cum eo
EXOD|24|3|venit ergo Moses et narravit plebi omnia verba Domini atque iudicia responditque cunctus populus una voce omnia verba Domini quae locutus est faciemus
EXOD|24|4|scripsit autem Moses universos sermones Domini et mane consurgens aedificavit altare ad radices montis et duodecim titulos per duodecim tribus Israhel
EXOD|24|5|misitque iuvenes de filiis Israhel et obtulerunt holocausta immolaveruntque victimas pacificas Domino vitulos
EXOD|24|6|tulit itaque Moses dimidiam partem sanguinis et misit in crateras partem autem residuam fudit super altare
EXOD|24|7|adsumensque volumen foederis legit audiente populo qui dixerunt omnia quae locutus est Dominus faciemus et erimus oboedientes
EXOD|24|8|ille vero sumptum sanguinem respersit in populum et ait hic est sanguis foederis quod pepigit Dominus vobiscum super cunctis sermonibus his
EXOD|24|9|ascenderuntque Moses et Aaron Nadab et Abiu et septuaginta de senioribus Israhel
EXOD|24|10|et viderunt Deum Israhel sub pedibus eius quasi opus lapidis sapphirini et quasi caelum cum serenum est
EXOD|24|11|nec super eos qui procul recesserant de filiis Israhel misit manum suam videruntque Deum et comederunt ac biberunt
EXOD|24|12|dixit autem Dominus ad Mosen ascende ad me in montem et esto ibi daboque tibi tabulas lapideas et legem ac mandata quae scripsi ut doceas eos
EXOD|24|13|surrexerunt Moses et Iosue minister eius ascendensque Moses in montem Dei
EXOD|24|14|senioribus ait expectate hic donec revertamur ad vos habetis Aaron et Hur vobiscum si quid natum fuerit quaestionis referetis ad eos
EXOD|24|15|cumque ascendisset Moses operuit nubes montem
EXOD|24|16|et habitavit gloria Domini super Sinai tegens illum nube sex diebus septimo autem die vocavit eum de medio caliginis
EXOD|24|17|erat autem species gloriae Domini quasi ignis ardens super verticem montis in conspectu filiorum Israhel
EXOD|24|18|ingressusque Moses medium nebulae ascendit in montem et fuit ibi quadraginta diebus et quadraginta noctibus
EXOD|25|1|locutusque est Dominus ad Mosen dicens
EXOD|25|2|loquere filiis Israhel ut tollant mihi primitias ab omni homine qui offert ultroneus accipietis eas
EXOD|25|3|haec sunt autem quae accipere debetis aurum et argentum et aes
EXOD|25|4|hyacinthum et purpuram coccumque bis tinctum et byssum pilos caprarum
EXOD|25|5|et pelles arietum rubricatas pelles ianthinas et ligna setthim
EXOD|25|6|oleum ad luminaria concinnanda aromata in unguentum et thymiama boni odoris
EXOD|25|7|lapides onychinos et gemmas ad ornandum ephod ac rationale
EXOD|25|8|facientque mihi sanctuarium et habitabo in medio eorum
EXOD|25|9|iuxta omnem similitudinem tabernaculi quod ostendam tibi et omnium vasorum in cultum eius sicque facietis illud
EXOD|25|10|arcam de lignis setthim conpingite cuius longitudo habeat duos semis cubitos latitudo cubitum et dimidium altitudo cubitum similiter ac semissem
EXOD|25|11|et deaurabis eam auro mundissimo intus et foris faciesque supra coronam auream per circuitum
EXOD|25|12|et quattuor circulos aureos quos pones per quattuor arcae angulos duo circuli sint in latere uno et duo in altero
EXOD|25|13|facies quoque vectes de lignis setthim et operies eos auro
EXOD|25|14|inducesque per circulos qui sunt in arcae lateribus ut portetur in eis
EXOD|25|15|qui semper erunt in circulis nec umquam extrahentur ab eis
EXOD|25|16|ponesque in arcam testificationem quam dabo tibi
EXOD|25|17|facies et propitiatorium de auro mundissimo duos cubitos et dimidium tenebit longitudo eius cubitum ac semissem latitudo
EXOD|25|18|duos quoque cherubin aureos et productiles facies ex utraque parte oraculi
EXOD|25|19|cherub unus sit in latere uno et alter in altero
EXOD|25|20|utrumque latus propitiatorii tegant expandentes alas et operientes oraculum respiciantque se mutuo versis vultibus in propitiatorium quo operienda est arca
EXOD|25|21|in qua pones testimonium quod dabo tibi
EXOD|25|22|inde praecipiam et loquar ad te supra propitiatorio scilicet ac medio duorum cherubin qui erunt super arcam testimonii cuncta quae mandabo per te filiis Israhel
EXOD|25|23|facies et mensam de lignis setthim habentem duos cubitos longitudinis et in latitudine cubitum et in altitudine cubitum ac semissem
EXOD|25|24|et inaurabis eam auro purissimo faciesque illi labium aureum per circuitum
EXOD|25|25|et ipsi labio coronam interrasilem altam quattuor digitis et super illam alteram coronam aureolam
EXOD|25|26|quattuor quoque circulos aureos praeparabis et pones eos in quattuor angulis eiusdem mensae per singulos pedes
EXOD|25|27|subter coronam erunt circuli aurei ut mittantur vectes per eos et possit mensa portari
EXOD|25|28|ipsosque vectes facies de lignis setthim et circumdabis auro ad subvehendam mensam
EXOD|25|29|parabis et acetabula ac fialas turibula et cyatos in quibus offerenda sunt libamina ex auro purissimo
EXOD|25|30|et pones super mensam panes propositionis in conspectu meo semper
EXOD|25|31|facies et candelabrum ductile de auro mundissimo hastile eius et calamos scyphos et spherulas ac lilia ex ipso procedentia
EXOD|25|32|sex calami egredientur de lateribus tres ex uno latere et tres ex altero
EXOD|25|33|tres scyphi quasi in nucis modum per calamos singulos spherulaque simul et lilium et tres similiter scyphi instar nucis in calamo altero spherulaque et lilium hoc erit opus sex calamorum qui producendi sunt de hastili
EXOD|25|34|in ipso autem candelabro erunt quattuor scyphi in nucis modum spherulaeque per singulos et lilia
EXOD|25|35|spherula sub duobus calamis per tria loca qui simul sex fiunt procedentes de hastili uno
EXOD|25|36|et spherae igitur et calami ex ipso erunt universa ductilia de auro purissimo
EXOD|25|37|facies et lucernas septem et pones eas super candelabrum ut luceant ex adverso
EXOD|25|38|emunctoria quoque et ubi quae emuncta sunt extinguantur fient de auro purissimo
EXOD|25|39|omne pondus candelabri cum universis vasis suis habebit talentum auri mundissimi
EXOD|25|40|inspice et fac secundum exemplar quod tibi in monte monstratum est
EXOD|26|1|tabernaculum vero ita fiet decem cortinas de bysso retorta et hyacintho ac purpura coccoque bis tincto variatas opere plumario facies
EXOD|26|2|longitudo cortinae unius habebit viginti octo cubitos latitudo quattuor cubitorum erit unius mensurae fient universa tentoria
EXOD|26|3|quinque cortinae sibi iungentur mutuo et aliae quinque nexu simili coherebunt
EXOD|26|4|ansulas hyacinthinas in lateribus ac summitatibus facies cortinarum ut possint invicem copulari
EXOD|26|5|quinquagenas ansulas cortina habebit in utraque parte ita insertas ut ansa contra ansam veniat et altera alteri possit aptari
EXOD|26|6|facies et quinquaginta circulos aureos quibus cortinarum vela iungenda sunt ut unum tabernaculum fiat
EXOD|26|7|facies et saga cilicina undecim ad operiendum tectum tabernaculi
EXOD|26|8|longitudo sagi unius habebit triginta cubitos et latitudo quattuor aequa erit mensura sagorum omnium
EXOD|26|9|e quibus quinque iunges seorsum et sex sibi mutuo copulabis ita ut sextum sagum in fronte tecti duplices
EXOD|26|10|facies et quinquaginta ansas in ora sagi unius ut coniungi cum altero queat et quinquaginta ansas in ora sagi alterius ut cum altero copuletur
EXOD|26|11|quinquaginta fibulas aeneas quibus iungantur ansae et unum ex omnibus operimentum fiat
EXOD|26|12|quod autem superfuerit in sagis quae parantur tecto id est unum sagum quod amplius est ex medietate eius operies posteriora tabernaculi
EXOD|26|13|et cubitus ex una parte pendebit et alter ex altera qui plus est in sagorum longitudine utrumque latus tabernaculi protegens
EXOD|26|14|facies et operimentum aliud tecto de pellibus arietum rubricatis et super hoc rursum aliud operimentum de ianthinis pellibus
EXOD|26|15|facies et tabulas stantes tabernaculi de lignis setthim
EXOD|26|16|quae singulae denos cubitos in longitudine habeant et in latitudine singulos ac semissem
EXOD|26|17|in lateribus tabulae duae incastraturae fient quibus tabula alteri tabulae conectatur atque in hunc modum cunctae tabulae parabuntur
EXOD|26|18|quarum viginti erunt in latere meridiano quod vergit ad austrum
EXOD|26|19|quibus quadraginta bases argenteas fundes ut binae bases singulis tabulis per duos angulos subiciantur
EXOD|26|20|in latere quoque secundo tabernaculi quod vergit ad aquilonem viginti tabulae erunt
EXOD|26|21|quadraginta habentes bases argenteas binae bases singulis tabulis subponentur
EXOD|26|22|ad occidentalem vero plagam tabernaculi facies sex tabulas
EXOD|26|23|et rursum alias duas quae in angulis erigantur post tergum tabernaculi
EXOD|26|24|eruntque coniunctae a deorsum usque sursum et una omnes conpago retinebit duabus quoque tabulis quae in angulis ponendae sunt similis iunctura servabitur
EXOD|26|25|et erunt simul tabulae octo bases earum argenteae sedecim duabus basibus per unam tabulam supputatis
EXOD|26|26|facies et vectes de lignis setthim quinque ad continendas tabulas in uno latere tabernaculi
EXOD|26|27|et quinque alios in altero et eiusdem numeri ad occidentalem plagam
EXOD|26|28|qui mittentur per medias tabulas a summo usque ad summum
EXOD|26|29|ipsasque tabulas deaurabis et fundes eis anulos aureos per quos vectes tabulata contineant quos operies lamminis aureis
EXOD|26|30|et eriges tabernaculum iuxta exemplum quod tibi in monte monstratum est
EXOD|26|31|facies et velum de hyacintho et purpura coccoque bis tincto et bysso retorta opere plumario et pulchra varietate contextum
EXOD|26|32|quod adpendes ante quattuor columnas de lignis setthim quae ipsae quidem deauratae erunt et habebunt capita aurea sed bases argenteas
EXOD|26|33|inseretur autem velum per circulos intra quod pones arcam testimonii et quo sanctuarium et sanctuarii sanctuaria dividentur
EXOD|26|34|pones et propitiatorium super arcam testimonii in sancta sanctorum
EXOD|26|35|mensamque extra velum et contra mensam candelabrum in latere tabernaculi meridiano mensa enim stabit in parte aquilonis
EXOD|26|36|facies et tentorium in introitu tabernaculi de hyacintho et purpura coccoque bis tincto et bysso retorta opere plumarii
EXOD|26|37|et quinque columnas deaurabis lignorum setthim ante quas ducetur tentorium quarum erunt capita aurea et bases aeneae
EXOD|27|1|facies et altare de lignis setthim quod habebit quinque cubitos in longitudine et totidem in latitudine id est quadrum et tres cubitos in altitudine
EXOD|27|2|cornua autem per quattuor angulos ex ipso erunt et operies illud aere
EXOD|27|3|faciesque in usus eius lebetas ad suscipiendos cineres et forcipes atque fuscinulas et ignium receptacula omnia vasa ex aere fabricabis
EXOD|27|4|craticulamque in modum retis aeneam per cuius quattuor angulos erunt quattuor anuli aenei
EXOD|27|5|quos pones subter arulam altaris eritque craticula usque ad altaris medium
EXOD|27|6|facies et vectes altaris de lignis setthim duos quos operies lamminis aeneis
EXOD|27|7|et induces per circulos eruntque ex utroque latere altaris ad portandum
EXOD|27|8|non solidum sed inane et cavum intrinsecus facies illud sicut tibi in monte monstratum est
EXOD|27|9|facies et atrium tabernaculi in cuius plaga australi contra meridiem erunt tentoria de bysso retorta centum cubitos unum latus tenebit in longitudine
EXOD|27|10|et columnas viginti cum basibus totidem aeneis quae capita cum celaturis suis habebunt argentea
EXOD|27|11|similiter in latere aquilonis per longum erunt tentoria centum cubitorum columnae viginti et bases aeneae eiusdem numeri et capita earum cum celaturis suis argentea
EXOD|27|12|in latitudine vero atrii quod respicit ad occidentem erunt tentoria per quinquaginta cubitos et columnae decem basesque totidem
EXOD|27|13|in ea quoque atrii latitudine quae respicit ad orientem quinquaginta cubiti erunt
EXOD|27|14|in quibus quindecim cubitorum tentoria lateri uno deputabuntur columnaeque tres et bases totidem
EXOD|27|15|et in latere altero erunt tentoria cubitos obtinentia quindecim columnas tres et bases totidem
EXOD|27|16|in introitu vero atrii fiet tentorium cubitorum viginti ex hyacintho et purpura coccoque bis tincto et bysso retorta opere plumarii columnas habebit quattuor cum basibus totidem
EXOD|27|17|omnes columnae atrii per circuitum vestitae erunt argenti lamminis capitibus argenteis et basibus aeneis
EXOD|27|18|in longitudine occupabit atrium cubitos centum in latitudine quinquaginta altitudo quinque cubitorum erit fietque de bysso retorta et habebit bases aeneas
EXOD|27|19|cuncta vasa tabernaculi in omnes usus et caerimonias tam paxillos eius quam atrii ex aere facies
EXOD|27|20|praecipe filiis Israhel ut adferant tibi oleum de arboribus olivarum purissimum piloque contusum ut ardeat lucerna semper
EXOD|27|21|in tabernaculo testimonii extra velum quod oppansum est testimonio et conlocabunt eam Aaron et filii eius ut usque mane luceat coram Domino perpetuus erit cultus per successiones eorum a filiis Israhel
EXOD|28|1|adplica quoque ad te Aaron fratrem tuum cum filiis suis de medio filiorum Israhel ut sacerdotio fungantur mihi Aaron Nadab et Abiu Eleazar et Ithamar
EXOD|28|2|faciesque vestem sanctam fratri tuo in gloriam et decorem
EXOD|28|3|et loqueris cunctis sapientibus corde quos replevi spiritu prudentiae ut faciant vestes Aaron in quibus sanctificatus ministret mihi
EXOD|28|4|haec autem erunt vestimenta quae facient rationale et superumerale tunicam et lineam strictam cidarim et balteum facient vestimenta sancta Aaron fratri tuo et filiis eius ut sacerdotio fungantur mihi
EXOD|28|5|accipientque aurum et hyacinthum et purpuram coccumque bis tinctum et byssum
EXOD|28|6|facient autem superumerale de auro et hyacintho ac purpura coccoque bis tincto et bysso retorta opere polymito
EXOD|28|7|duas oras iunctas habebit in utroque latere summitatum ut in unum redeant
EXOD|28|8|ipsaque textura et cuncta operis varietas erit ex auro et hyacintho et purpura coccoque bis tincto et bysso retorta
EXOD|28|9|sumesque duos lapides onychinos et sculpes in eis nomina filiorum Israhel
EXOD|28|10|sex nomina in lapide uno et sex reliqua in altero iuxta ordinem nativitatis eorum
EXOD|28|11|opere sculptoris et celatura gemmarii sculpes eos nominibus filiorum Israhel inclusos auro atque circumdatos
EXOD|28|12|et pones in utroque latere superumeralis memoriale filiis Israhel portabitque Aaron nomina eorum coram Domino super utrumque umerum ob recordationem
EXOD|28|13|facies et uncinos ex auro
EXOD|28|14|et duas catenulas auri purissimi sibi invicem coherentes quas inseres uncinis
EXOD|28|15|rationale quoque iudicii facies opere polymito iuxta texturam superumeralis ex auro hyacintho et purpura coccoque bis tincto et bysso retorta
EXOD|28|16|quadrangulum erit et duplex mensuram palmi habebit tam in longitudine quam in latitudine
EXOD|28|17|ponesque in eo quattuor ordines lapidum in primo versu erit lapis sardius et topazius et zmaragdus
EXOD|28|18|in secundo carbunculus sapphyrus et iaspis
EXOD|28|19|in tertio ligyrius achates et amethistus
EXOD|28|20|in quarto chrysolitus onychinus et berillus inclusi auro erunt per ordines suos
EXOD|28|21|habebuntque nomina filiorum Israhel duodecim nominibus celabuntur singuli lapides nominibus singulorum per duodecim tribus
EXOD|28|22|facies in rationali catenas sibi invicem coherentes ex auro purissimo
EXOD|28|23|et duos anulos aureos quos pones in utraque rationalis summitate
EXOD|28|24|catenasque aureas iunges anulis qui sunt in marginibus eius
EXOD|28|25|et ipsarum catenarum extrema duobus copulabis uncinis in utroque latere superumeralis quod rationale respicit
EXOD|28|26|facies et duos anulos aureos quos pones in summitatibus rationalis et in oris quae e regione sunt superumeralis et posteriora eius aspiciunt
EXOD|28|27|nec non et alios duos anulos aureos qui ponendi sunt in utroque latere superumeralis deorsum quod respicit contra faciem iuncturae inferioris ut aptari possit cum superumerali
EXOD|28|28|et stringatur rationale anulis suis cum anulis superumeralis vitta hyacinthina ut maneat iunctura fabrefacta et a se invicem rationale et superumerale nequeant separari
EXOD|28|29|portabitque Aaron nomina filiorum Israhel in rationali iudicii super pectus suum quando ingreditur sanctuarium memoriale coram Domino in aeternum
EXOD|28|30|pones autem in rationali iudicii doctrinam et veritatem quae erunt in pectore Aaron quando ingreditur coram Domino et gestabit iudicium filiorum Israhel in pectore suo in conspectu Domini semper
EXOD|28|31|facies et tunicam superumeralis totam hyacinthinam
EXOD|28|32|in cuius medio supra erit capitium et ora per gyrum eius textilis sicut fieri solet in extremis vestium partibus ne facile rumpatur
EXOD|28|33|deorsum vero ad pedes eiusdem tunicae per circuitum quasi mala punica facies ex hyacintho et purpura et cocco bis tincto mixtis in medio tintinabulis
EXOD|28|34|ita ut tintinabulum sit aureum et malum rursumque tintinabulum aliud aureum et malum punicum
EXOD|28|35|et vestietur ea Aaron in officio ministerii ut audiatur sonitus quando ingreditur et egreditur sanctuarium in conspectu Domini et non moriatur
EXOD|28|36|facies et lamminam de auro purissimo in qua sculpes opere celatoris Sanctum Domino
EXOD|28|37|ligabisque eam vitta hyacinthina et erit super tiaram
EXOD|28|38|inminens fronti pontificis portabitque Aaron iniquitates eorum quae obtulerint et sanctificaverint filii Israhel in cunctis muneribus et donariis suis erit autem lammina semper in fronte eius ut placatus eis sit Dominus
EXOD|28|39|stringesque tunicam bysso et tiaram byssinam facies et balteum opere plumarii
EXOD|28|40|porro filiis Aaron tunicas lineas parabis et balteos ac tiaras in gloriam et decorem
EXOD|28|41|vestiesque his omnibus Aaron fratrem tuum et filios eius cum eo et cunctorum consecrabis manus sanctificabisque illos ut sacerdotio fungantur mihi
EXOD|28|42|facies et feminalia linea ut operiant carnem turpitudinis suae a renibus usque ad femina
EXOD|28|43|et utentur eis Aaron et filii eius quando ingredientur tabernaculum testimonii vel quando adpropinquant ad altare ut ministrent in sanctuario ne iniquitatis rei moriantur legitimum sempiternum erit Aaron et semini eius post eum
EXOD|29|1|sed et hoc facies ut mihi in sacerdotio consecrentur tolle vitulum de armento et arietes duos inmaculatos
EXOD|29|2|panesque azymos et crustula absque fermento quae conspersa sint oleo lagana quoque azyma oleo lita de simila triticea cuncta facies
EXOD|29|3|et posita in canistro offeres vitulum autem et duos arietes
EXOD|29|4|et Aaron ac filios eius adplicabis ad ostium tabernaculi testimonii cumque laveris patrem cum filiis aqua
EXOD|29|5|indues Aaron vestimentis suis id est linea et tunica et superumerali et rationali quod constringes balteo
EXOD|29|6|et pones tiaram in capite eius et lamminam sanctam super tiaram
EXOD|29|7|et oleum unctionis fundes super caput eius atque hoc ritu consecrabitur
EXOD|29|8|filios quoque illius adplicabis et indues tunicis lineis cingesque balteo
EXOD|29|9|Aaron scilicet et liberos eius et inpones eis mitras eruntque sacerdotes mei in religione perpetua postquam initiaveris manus eorum
EXOD|29|10|adplicabis et vitulum coram tabernaculo testimonii inponentque Aaron et filii eius manus super caput illius
EXOD|29|11|et mactabis eum in conspectu Domini iuxta ostium tabernaculi testimonii
EXOD|29|12|sumptumque de sanguine vituli pones super cornua altaris digito tuo reliquum autem sanguinem fundes iuxta basim eius
EXOD|29|13|sumes et adipem totum qui operit intestina et reticulum iecoris ac duos renes et adipem qui super eos est et offeres incensum super altare
EXOD|29|14|carnes vero vituli et corium et fimum conbures foris extra castra eo quod pro peccato sit
EXOD|29|15|unum quoque arietum sumes super cuius caput ponent Aaron et filii eius manus
EXOD|29|16|quem cum mactaveris tolles de sanguine eius et fundes circa altare
EXOD|29|17|ipsum autem arietem secabis in frusta lotaque intestina eius ac pedes pones super concisas carnes et super caput illius
EXOD|29|18|et offeres totum arietem in incensum super altare oblatio est Domini odor suavissimus victimae Dei
EXOD|29|19|tolles quoque arietem alterum super cuius caput Aaron et filii eius ponent manus
EXOD|29|20|quem cum immolaveris sumes de sanguine ipsius et pones super extremum dextrae auriculae Aaron et filiorum eius et super pollices manus eorum et pedis dextri fundesque sanguinem super altare per circuitum
EXOD|29|21|cumque tuleris de sanguine qui est super altare et de oleo unctionis asperges Aaron et vestes eius filios et vestimenta eorum consecratisque et ipsis et vestibus
EXOD|29|22|tolles adipem de ariete et caudam et arvinam quae operit vitalia ac reticulum iecoris et duos renes atque adipem qui super eos est armumque dextrum eo quod sit aries consecrationum
EXOD|29|23|tortam panis unius crustulum conspersum oleo laganum de canistro azymorum quod positum est in conspectu Domini
EXOD|29|24|ponesque omnia super manus Aaron et filiorum eius et sanctificabis eos elevans coram Domino
EXOD|29|25|suscipiesque universa de manibus eorum et incendes super altare in holocaustum odorem suavissimum in conspectu Domini quia oblatio eius est
EXOD|29|26|sumes quoque pectusculum de ariete quo initiatus est Aaron sanctificabisque illud elatum coram Domino et cedet in partem tuam
EXOD|29|27|sanctificabis et pectusculum consecratum et armum quem de ariete separasti
EXOD|29|28|quo initiatus est Aaron et filii eius cedentque in partem Aaron et filiorum eius iure perpetuo a filiis Israhel quia primitiva sunt et initia de victimis eorum pacificis quae offerunt Domino
EXOD|29|29|vestem autem sanctam qua utitur Aaron habebunt filii eius post eum ut unguantur in ea et consecrentur manus eorum
EXOD|29|30|septem diebus utetur illa qui pontifex pro eo fuerit constitutus de filiis eius et qui ingredietur tabernaculum testimonii ut ministret in sanctuario
EXOD|29|31|arietem autem consecrationum tolles et coques carnes eius in loco sancto
EXOD|29|32|quibus vescetur Aaron et filii eius panes quoque qui sunt in canistro in vestibulo tabernaculi testimonii comedent
EXOD|29|33|ut sit placabile sacrificium et sanctificentur offerentium manus alienigena non vescetur ex eis quia sancti sunt
EXOD|29|34|quod si remanserit de carnibus consecratis sive de panibus usque mane conbures reliquias igni non comedentur quia sanctificata sunt
EXOD|29|35|omnia quae praecepi tibi facies super Aaron et filiis eius septem diebus consecrabis manus eorum
EXOD|29|36|et vitulum pro peccato offeres per singulos dies ad expiandum mundabisque altare cum immolaris expiationis hostiam et ungues illud in sanctificationem
EXOD|29|37|septem diebus expiabis altare et sanctificabis et erit sanctum sanctorum omnis qui tetigerit illud sanctificabitur
EXOD|29|38|hoc est quod facies in altari agnos anniculos duos per singulos dies iugiter
EXOD|29|39|unum agnum mane et alterum vespere
EXOD|29|40|decimam partem similae conspersae oleo tunso quod habeat mensuram quartam partem hin et vinum ad libandum eiusdem mensurae in agno uno
EXOD|29|41|alterum vero agnum offeres ad vesperam iuxta ritum matutinae oblationis et iuxta ea quae diximus in odorem suavitatis
EXOD|29|42|sacrificium Domino oblatione perpetua in generationes vestras ad ostium tabernaculi testimonii coram Domino ubi constituam ut loquar ad te
EXOD|29|43|ibique praecipiam filiis Israhel et sanctificabitur altare in gloria mea
EXOD|29|44|sanctificabo et tabernaculum testimonii cum altari et Aaron cum filiis eius ut sacerdotio fungantur mihi
EXOD|29|45|et habitabo in medio filiorum Israhel eroque eis Deus
EXOD|29|46|et scient quia ego Dominus Deus eorum qui eduxi eos de terra Aegypti ut manerem inter illos ego Dominus Deus ipsorum
EXOD|30|1|facies quoque altare in adolendum thymiama de lignis setthim
EXOD|30|2|habens cubitum longitudinis et alterum latitudinis id est quadrangulum et duos cubitos in altitudine cornua ex ipso procedent
EXOD|30|3|vestiesque illud auro purissimo tam craticulam eius quam parietes per circuitum et cornua faciesque ei coronam aureolam per gyrum
EXOD|30|4|et duos anulos aureos sub corona per singula latera ut mittantur in eos vectes et altare portetur
EXOD|30|5|ipsos quoque vectes facies de lignis setthim et inaurabis
EXOD|30|6|ponesque altare contra velum quod ante arcam pendet testimonii coram propitiatorio quo tegitur testimonium ubi loquar tibi
EXOD|30|7|et adolebit incensum super eo Aaron suave fraglans mane quando conponet lucernas incendet illud
EXOD|30|8|et quando conlocat eas ad vesperum uret thymiama sempiternum coram Domino in generationes vestras
EXOD|30|9|non offeretis super eo thymiama conpositionis alterius nec oblationem et victimam nec liba libabitis
EXOD|30|10|et deprecabitur Aaron super cornua eius semel per annum in sanguine quod oblatum est pro peccato et placabit super eo in generationibus vestris sanctum sanctorum erit Domino
EXOD|30|11|locutusque est Dominus ad Mosen dicens
EXOD|30|12|quando tuleris summam filiorum Israhel iuxta numerum dabunt singuli pretium pro animabus suis Domino et non erit plaga in eis cum fuerint recensiti
EXOD|30|13|hoc autem dabit omnis qui transit ad nomen dimidium sicli iuxta mensuram templi siclus viginti obolos habet media pars sicli offeretur Domino
EXOD|30|14|qui habetur in numero a viginti annis et supra dabit pretium
EXOD|30|15|dives non addet ad medium sicli et pauper nihil minuet
EXOD|30|16|susceptamque pecuniam quae conlata est a filiis Israhel trades in usus tabernaculi testimonii ut sit monumentum eorum coram Domino et propitietur animabus illorum
EXOD|30|17|locutusque est Dominus ad Mosen dicens
EXOD|30|18|facies et labium aeneum cum basi sua ad lavandum ponesque illud inter tabernaculum testimonii et altare et missa aqua
EXOD|30|19|lavabunt in eo Aaron et filii eius manus suas ac pedes
EXOD|30|20|quando ingressuri sunt tabernaculum testimonii et quando accessuri ad altare ut offerant in eo thymiama Domino
EXOD|30|21|ne forte moriantur legitimum sempiternum erit ipsi et semini eius per successiones
EXOD|30|22|locutusque est Dominus ad Mosen
EXOD|30|23|dicens sume tibi aromata prima et zmyrnae electae quingentos siclos et cinnamomi medium id est ducentos quinquaginta calami similiter ducentos quinquaginta
EXOD|30|24|cassiae autem quingentos siclos in pondere sanctuarii olei de olivetis mensuram hin
EXOD|30|25|faciesque unctionis oleum sanctum unguentum conpositum opere unguentarii
EXOD|30|26|et ungues ex eo tabernaculum testimonii et arcam testamenti
EXOD|30|27|mensamque cum vasis suis candelabrum et utensilia eius altaria thymiamatis
EXOD|30|28|et holocausti et universam supellectilem quae ad cultum eorum pertinent
EXOD|30|29|sanctificabisque omnia et erunt sancta sanctorum qui tetigerit ea sanctificabitur
EXOD|30|30|Aaron et filios eius ungues sanctificabisque eos ut sacerdotio fungantur mihi
EXOD|30|31|filiis quoque Israhel dices hoc oleum unctionis sanctum erit mihi in generationes vestras
EXOD|30|32|caro hominis non unguetur ex eo et iuxta conpositionem eius non facietis aliud quia sanctificatum est et sanctum erit vobis
EXOD|30|33|homo quicumque tale conposuerit et dederit ex eo alieno exterminabitur de populo suo
EXOD|30|34|dixitque Dominus ad Mosen sume tibi aromata stacten et onycha galbanen boni odoris et tus lucidissimum aequalis ponderis erunt omnia
EXOD|30|35|faciesque thymiama conpositum opere unguentarii mixtum diligenter et purum et sanctificatione dignissimum
EXOD|30|36|cumque in tenuissimum pulverem universa contuderis pones ex eo coram testimonio tabernaculi in quo loco apparebo tibi sanctum sanctorum erit vobis thymiama
EXOD|30|37|talem conpositionem non facietis in usus vestros quia sanctum est Domino
EXOD|30|38|homo quicumque fecerit simile ut odore illius perfruatur peribit de populis suis
EXOD|31|1|locutusque est Dominus ad Mosen dicens
EXOD|31|2|ecce vocavi ex nomine Beselehel filium Uri filii Hur de tribu Iuda
EXOD|31|3|et implevi eum spiritu Dei sapientia intellegentia et scientia in omni opere
EXOD|31|4|ad excogitandum fabre quicquid fieri potest ex auro et argento et aere
EXOD|31|5|marmore et gemmis et diversitate lignorum
EXOD|31|6|dedique ei socium Hooliab filium Achisamech de tribu Dan et in corde omnis eruditi posui sapientiam ut faciant cuncta quae praecepi tibi
EXOD|31|7|tabernaculum foederis et arcam testimonii et propitiatorium quod super eam est et cuncta vasa tabernaculi
EXOD|31|8|mensamque et vasa eius candelabrum purissimum cum vasis suis et altaria thymiamatis
EXOD|31|9|et holocausti et omnia vasa eorum labium cum basi sua
EXOD|31|10|vestes sanctas in ministerio Aaron sacerdoti et filiis eius ut fungantur officio suo in sacris
EXOD|31|11|oleum unctionis et thymiama aromatum in sanctuario omnia quae praecepi tibi facient
EXOD|31|12|et locutus est Dominus ad Mosen dicens
EXOD|31|13|loquere filiis Israhel et dices ad eos videte ut sabbatum meum custodiatis quia signum est inter me et vos in generationibus vestris ut sciatis quia ego Dominus qui sanctifico vos
EXOD|31|14|custodite sabbatum sanctum est enim vobis qui polluerit illud morte morietur qui fecerit in eo opus peribit anima illius de medio populi sui
EXOD|31|15|sex diebus facietis opus in die septimo sabbatum est requies sancta Domino omnis qui fecerit opus in hac die morietur
EXOD|31|16|custodiant filii Israhel sabbatum et celebrent illud in generationibus suis pactum est sempiternum
EXOD|31|17|inter me et filios Israhel signumque perpetuum sex enim diebus fecit Dominus caelum et terram et in septimo ab opere cessavit
EXOD|31|18|dedit quoque Mosi conpletis huiuscemodi sermonibus in monte Sinai duas tabulas testimonii lapideas scriptas digito Dei
EXOD|32|1|videns autem populus quod moram faceret descendendi de monte Moses congregatus adversus Aaron ait surge fac nobis deos qui nos praecedant Mosi enim huic viro qui nos eduxit de terra Aegypti ignoramus quid acciderit
EXOD|32|2|dixitque ad eos Aaron tollite inaures aureas de uxorum filiorumque et filiarum vestrarum auribus et adferte ad me
EXOD|32|3|fecit populus quae iusserat deferens inaures ad Aaron
EXOD|32|4|quas cum ille accepisset formavit opere fusorio et fecit ex eis vitulum conflatilem dixeruntque hii sunt dii tui Israhel qui te eduxerunt de terra Aegypti
EXOD|32|5|quod cum vidisset Aaron aedificavit altare coram eo et praeconis voce clamavit dicens cras sollemnitas Domini est
EXOD|32|6|surgentesque mane obtulerunt holocausta et hostias pacificas et sedit populus comedere ac bibere et surrexerunt ludere
EXOD|32|7|locutus est autem Dominus ad Mosen vade descende peccavit populus tuus quem eduxisti de terra Aegypti
EXOD|32|8|recesserunt cito de via quam ostendisti eis feceruntque sibi vitulum conflatilem et adoraverunt atque immolantes ei hostias dixerunt isti sunt dii tui Israhel qui te eduxerunt de terra Aegypti
EXOD|32|9|rursumque ait Dominus ad Mosen cerno quod populus iste durae cervicis sit
EXOD|32|10|dimitte me ut irascatur furor meus contra eos et deleam eos faciamque te in gentem magnam
EXOD|32|11|Moses autem orabat Dominum Deum suum dicens cur Domine irascitur furor tuus contra populum tuum quem eduxisti de terra Aegypti in fortitudine magna et in manu robusta
EXOD|32|12|ne quaeso dicant Aegyptii callide eduxit eos ut interficeret in montibus et deleret e terra quiescat ira tua et esto placabilis super nequitia populi tui
EXOD|32|13|recordare Abraham Isaac et Israhel servorum tuorum quibus iurasti per temet ipsum dicens multiplicabo semen vestrum sicut stellas caeli et universam terram hanc de qua locutus sum dabo semini vestro et possidebitis eam semper
EXOD|32|14|placatusque est Dominus ne faceret malum quod locutus fuerat adversus populum suum
EXOD|32|15|et reversus est Moses de monte portans duas tabulas testimonii manu scriptas ex utraque parte
EXOD|32|16|et factas opere Dei scriptura quoque Dei erat sculpta in tabulis
EXOD|32|17|audiens autem Iosue tumultum populi vociferantis dixit ad Mosen ululatus pugnae auditur in castris
EXOD|32|18|qui respondit non est clamor adhortantium ad pugnam neque vociferatio conpellentium ad fugam sed vocem cantantium ego audio
EXOD|32|19|cumque adpropinquasset ad castra vidit vitulum et choros iratusque valde proiecit de manu tabulas et confregit eas ad radices montis
EXOD|32|20|arripiensque vitulum quem fecerant conbusit et contrivit usque ad pulverem quem sparsit in aqua et dedit ex eo potum filiis Israhel
EXOD|32|21|dixitque ad Aaron quid tibi fecit hic populus ut induceres super eum peccatum maximum
EXOD|32|22|cui ille respondit ne indignetur dominus meus tu enim nosti populum istum quod pronus sit ad malum
EXOD|32|23|dixerunt mihi fac nobis deos qui praecedant nos huic enim Mosi qui nos eduxit de terra Aegypti nescimus quid acciderit
EXOD|32|24|quibus ego dixi quis vestrum habet aurum tulerunt et dederunt mihi et proieci illud in ignem egressusque est hic vitulus
EXOD|32|25|videns ergo Moses populum quod esset nudatus spoliaverat enim eum Aaron propter ignominiam sordis et inter hostes nudum constituerat
EXOD|32|26|et stans in porta castrorum ait si quis est Domini iungatur mihi congregatique sunt ad eum omnes filii Levi
EXOD|32|27|quibus ait haec dicit Dominus Deus Israhel ponat vir gladium super femur suum ite et redite de porta usque ad portam per medium castrorum et occidat unusquisque fratrem et amicum et proximum suum
EXOD|32|28|fecerunt filii Levi iuxta sermonem Mosi cecideruntque in die illo quasi tria milia hominum
EXOD|32|29|et ait Moses consecrastis manus vestras hodie Domino unusquisque in filio et fratre suo ut detur vobis benedictio
EXOD|32|30|facto autem die altero locutus est Moses ad populum peccastis peccatum maximum ascendam ad Dominum si quo modo eum quivero deprecari pro scelere vestro
EXOD|32|31|reversusque ad Dominum ait obsecro peccavit populus iste peccatum magnum feceruntque sibi deos aureos aut dimitte eis hanc noxam
EXOD|32|32|aut si non facis dele me de libro tuo quem scripsisti
EXOD|32|33|cui respondit Dominus qui peccaverit mihi delebo eum de libro meo
EXOD|32|34|tu autem vade et duc populum istum quo locutus sum tibi angelus meus praecedet te ego autem in die ultionis visitabo et hoc peccatum eorum
EXOD|32|35|percussit ergo Dominus populum pro reatu vituli quem fecit Aaron
EXOD|33|1|locutusque est Dominus ad Mosen vade ascende de loco isto tu et populus tuus quem eduxisti de terra Aegypti in terram quam iuravi Abraham Isaac et Iacob dicens semini tuo dabo eam
EXOD|33|2|et mittam praecursorem tui angelum ut eiciam Chananeum et Amorreum et Hettheum et Ferezeum et Eveum et Iebuseum
EXOD|33|3|et intres in terram fluentem lacte et melle non enim ascendam tecum quia populus durae cervicis est ne forte disperdam te in via
EXOD|33|4|audiens populus sermonem hunc pessimum luxit et nullus ex more indutus est cultu suo
EXOD|33|5|dixitque Dominus ad Mosen loquere filiis Israhel populus durae cervicis es semel ascendam in medio tui et delebo te iam nunc depone ornatum tuum ut sciam quid faciam tibi
EXOD|33|6|deposuerunt ergo filii Israhel ornatum suum a monte Horeb
EXOD|33|7|Moses quoque tollens tabernaculum tetendit extra castra procul vocavitque nomen eius tabernaculum foederis et omnis populus qui habebat aliquam quaestionem egrediebatur ad tabernaculum foederis extra castra
EXOD|33|8|cumque egrederetur Moses ad tabernaculum surgebat universa plebs et stabat unusquisque in ostio papilionis sui aspiciebantque tergum Mosi donec ingrederetur tentorium
EXOD|33|9|ingresso autem illo tabernaculum foederis descendebat columna nubis et stabat ad ostium loquebaturque cum Mosi
EXOD|33|10|cernentibus universis quod columna nubis staret ad ostium tabernaculi stabantque ipsi et adorabant per fores tabernaculorum suorum
EXOD|33|11|loquebatur autem Dominus ad Mosen facie ad faciem sicut loqui solet homo ad amicum suum cumque ille reverteretur in castra minister eius Iosue filius Nun puer non recedebat de tabernaculo
EXOD|33|12|dixit autem Moses ad Dominum praecipis ut educam populum istum et non indicas mihi quem missurus es mecum praesertim cum dixeris novi te ex nomine et invenisti gratiam coram me
EXOD|33|13|si ergo inveni gratiam in conspectu tuo ostende mihi viam tuam ut sciam te et inveniam gratiam ante oculos tuos respice populum tuum gentem hanc
EXOD|33|14|dixitque Dominus facies mea praecedet te et requiem dabo tibi
EXOD|33|15|et ait Moses si non tu ipse praecedes ne educas nos de loco isto
EXOD|33|16|in quo enim scire poterimus ego et populus tuus invenisse nos gratiam in conspectu tuo nisi ambulaveris nobiscum ut glorificemur ab omnibus populis qui habitant super terram
EXOD|33|17|dixit autem Dominus ad Mosen et verbum istud quod locutus es faciam invenisti enim gratiam coram me et te ipsum novi ex nomine
EXOD|33|18|qui ait ostende mihi gloriam tuam
EXOD|33|19|respondit ego ostendam omne bonum tibi et vocabo in nomine Domini coram te et miserebor cui voluero et clemens ero in quem mihi placuerit
EXOD|33|20|rursumque ait non poteris videre faciem meam non enim videbit me homo et vivet
EXOD|33|21|et iterum ecce inquit est locus apud me stabis super petram
EXOD|33|22|cumque transibit gloria mea ponam te in foramine petrae et protegam dextera mea donec transeam
EXOD|33|23|tollamque manum meam et videbis posteriora mea faciem autem meam videre non poteris
EXOD|34|1|ac deinceps praecide ait tibi duas tabulas lapideas instar priorum et scribam super eas verba quae habuerunt tabulae quas fregisti
EXOD|34|2|esto paratus mane ut ascendas statim in montem Sinai stabisque mecum super verticem montis
EXOD|34|3|nullus ascendat tecum nec videatur quispiam per totum montem boves quoque et oves non pascantur e contra
EXOD|34|4|excidit ergo duas tabulas lapideas quales ante fuerant et de nocte consurgens ascendit in montem Sinai sicut ei praeceperat Dominus portans secum tabulas
EXOD|34|5|cumque descendisset Dominus per nubem stetit Moses cum eo invocans nomen Domini
EXOD|34|6|quo transeunte coram eo ait Dominator Domine Deus misericors et clemens patiens et multae miserationis ac verus
EXOD|34|7|qui custodis misericordiam in milia qui aufers iniquitatem et scelera atque peccata nullusque apud te per se innocens est qui reddis iniquitatem patrum in filiis ac nepotibus in tertiam et quartam progeniem
EXOD|34|8|festinusque Moses curvatus est pronus in terram et adorans
EXOD|34|9|ait si inveni gratiam in conspectu tuo Domine obsecro ut gradiaris nobiscum populus enim durae cervicis est et auferas iniquitates nostras atque peccata nosque possideas
EXOD|34|10|respondit Dominus ego inibo pactum videntibus cunctis signa faciam quae numquam sunt visa super terram nec in ullis gentibus ut cernat populus in cuius es medio opus Domini terribile quod facturus sum
EXOD|34|11|observa cuncta quae hodie mando tibi ego ipse eiciam ante faciem tuam Amorreum et Chananeum et Hettheum Ferezeum quoque et Eveum et Iebuseum
EXOD|34|12|cave ne umquam cum habitatoribus terrae illius iungas amicitias quae tibi sint in ruinam
EXOD|34|13|sed aras eorum destrue confringe statuas lucosque succide
EXOD|34|14|noli adorare deum alienum Dominus Zelotes nomen eius Deus est aemulator
EXOD|34|15|ne ineas pactum cum hominibus illarum regionum ne cum fornicati fuerint cum diis suis et adoraverint simulacra eorum vocet te quispiam ut comedas de immolatis
EXOD|34|16|nec uxorem de filiabus eorum accipies filiis tuis ne postquam ipsae fuerint fornicatae fornicari faciant et filios tuos in deos suos
EXOD|34|17|deos conflatiles non facies tibi
EXOD|34|18|sollemnitatem azymorum custodies septem diebus vesceris azymis sicut praecepi tibi in tempore mensis novorum mense enim verni temporis egressus es de Aegypto
EXOD|34|19|omne quod aperit vulvam generis masculini meum erit de cunctis animantibus tam de bubus quam de ovibus meum erit
EXOD|34|20|primogenitum asini redimes ove sin autem nec pretium pro eo dederis occidetur primogenitum filiorum tuorum redimes nec apparebis in conspectu meo vacuus
EXOD|34|21|sex diebus operaberis die septimo cessabis arare et metere
EXOD|34|22|sollemnitatem ebdomadarum facies tibi in primitiis frugum messis tuae triticeae et sollemnitatem quando redeunte anni tempore cuncta conduntur
EXOD|34|23|tribus temporibus anni apparebit omne masculinum tuum in conspectu omnipotentis Domini Dei Israhel
EXOD|34|24|cum enim tulero gentes a facie tua et dilatavero terminos tuos nullus insidiabitur terrae tuae ascendente te et apparente in conspectu Domini Dei tui ter in anno
EXOD|34|25|non immolabis super fermento sanguinem hostiae meae neque residebit mane de victima sollemnitatis phase
EXOD|34|26|primitias frugum terrae tuae offeres in domum Domini Dei tui non coques hedum in lacte matris suae
EXOD|34|27|dixitque Dominus ad Mosen scribe tibi verba haec quibus et tecum et cum Israhel pepigi foedus
EXOD|34|28|fecit ergo ibi cum Domino quadraginta dies et quadraginta noctes panem non comedit et aquam non bibit et scripsit in tabulis verba foederis decem
EXOD|34|29|cumque descenderet Moses de monte Sinai tenebat duas tabulas testimonii et ignorabat quod cornuta esset facies sua ex consortio sermonis Dei
EXOD|34|30|videntes autem Aaron et filii Israhel cornutam Mosi faciem timuerunt prope accedere
EXOD|34|31|vocatique ab eo reversi sunt tam Aaron quam principes synagogae et postquam locutus est
EXOD|34|32|venerunt ad eum etiam omnes filii Israhel quibus praecepit cuncta quae audierat a Domino in monte Sinai
EXOD|34|33|impletisque sermonibus posuit velamen super faciem suam
EXOD|34|34|quod ingressus ad Dominum et loquens cum eo auferebat donec exiret et tunc loquebatur ad filios Israhel omnia quae sibi fuerant imperata
EXOD|34|35|qui videbant faciem egredientis Mosi esse cornutam sed operiebat rursus ille faciem suam si quando loquebatur ad eos
EXOD|35|1|igitur congregata omni turba filiorum Israhel dixit ad eos haec sunt quae iussit Dominus fieri
EXOD|35|2|sex diebus facietis opus septimus dies erit vobis sanctus sabbatum et requies Domini qui fecerit opus in eo occidetur
EXOD|35|3|non succendetis ignem in omnibus habitaculis vestris per diem sabbati
EXOD|35|4|et ait Moses ad omnem catervam filiorum Israhel iste est sermo quem praecepit Dominus dicens
EXOD|35|5|separate apud vos primitias Domino omnis voluntarius et proni animi offerat eas Domino aurum et argentum et aes
EXOD|35|6|hyacinthum purpuram coccumque bis tinctum et byssum pilos caprarum
EXOD|35|7|et pelles arietum rubricatas et ianthinas
EXOD|35|8|ligna setthim
EXOD|35|9|et oleum ad luminaria concinnanda et ut conficiatur unguentum et thymiama suavissimum
EXOD|35|10|lapides onychinos et gemmas ad ornatum superumeralis et rationalis
EXOD|35|11|quisquis vestrum est sapiens veniat et faciat quod Dominus imperavit
EXOD|35|12|tabernaculum scilicet et tectum eius atque operimentum anulos et tabulata cum vectibus paxillos et bases
EXOD|35|13|arcam et vectes propitiatorium et velum quod ante illud oppanditur
EXOD|35|14|mensam cum vectibus et vasis et propositionis panibus
EXOD|35|15|candelabrum ad luminaria sustentanda vasa illius et lucernas et oleum ad nutrimenta ignium
EXOD|35|16|altare thymiamatis et vectes oleum unctionis et thymiama ex aromatibus tentorium ad ostium tabernaculi
EXOD|35|17|altare holocausti et craticulam eius aeneam cum vectibus et vasis suis labrum et basim eius
EXOD|35|18|cortinas atrii cum columnis et basibus tentorium in foribus vestibuli
EXOD|35|19|paxillos tabernaculi et atrii cum funiculis suis
EXOD|35|20|vestimenta quorum usus est in ministerio sanctuarii vestes Aaron pontificis ac filiorum eius ut sacerdotio fungantur mihi
EXOD|35|21|egressaque omnis multitudo filiorum Israhel de conspectu Mosi
EXOD|35|22|obtulit mente promptissima atque devota primitias Domino ad faciendum opus tabernaculi testimonii quicquid in cultum et ad vestes sanctas necessarium erat
EXOD|35|23|viri cum mulieribus praebuerunt armillas et inaures anulos et dextralia omne vas aureum in donaria Domini separatum est
EXOD|35|24|si quis habuit hyacinthum purpuram coccumque bis tinctum byssum et pilos caprarum pelles arietum rubricatas et ianthinas
EXOD|35|25|argenti et aeris metalla obtulerunt Domino lignaque setthim in varios usus
EXOD|35|26|sed et mulieres doctae dederunt quae neverant hyacinthum purpuram et vermiculum ac byssum
EXOD|35|27|et pilos caprarum sponte propria cuncta tribuentes
EXOD|35|28|principes vero obtulerunt lapides onychinos et gemmas ad superumerale et rationale
EXOD|35|29|aromataque et oleum ad luminaria concinnanda et ad praeparandum unguentum ac thymiama odoris suavissimi conponendum
EXOD|35|30|omnes viri et mulieres mente devota obtulerunt donaria ut fierent opera quae iusserat Dominus per manum Mosi cuncti filii Israhel voluntaria Domino dedicaverunt
EXOD|35|31|dixitque Moses ad filios Israhel ecce vocavit Dominus ex nomine Beselehel filium Uri filii Hur de tribu Iuda
EXOD|35|32|implevitque eum spiritu Dei sapientiae et intellegentiae et scientiae omni doctrina
EXOD|35|33|ad excogitandum et faciendum opus in auro et argento et aere sculpendisque lapidibus et opere carpentario quicquid fabre adinveniri potest
EXOD|35|34|dedit in corde eius Hooliab quoque filium Achisamech de tribu Dan
EXOD|35|35|ambos erudivit sapientia ut faciant opera abietarii polymitarii ac plumarii de hyacintho et purpura coccoque bis tincto et bysso et texant omnia ac nova quaeque repperiant
EXOD|36|1|fecit ergo Beselehel et Hooliab et omnis vir sapiens quibus dedit Dominus sapientiam et intellectum ut scirent fabre operari quae in usus sanctuarii necessaria sunt et quae praecepit Dominus
EXOD|36|2|cumque vocasset eos Moses et omnem eruditum virum cui dederat Deus sapientiam et qui sponte sua obtulerant se ad faciendum opus
EXOD|36|3|tradidit eis universa donaria filiorum Israhel qui cum instarent operi cotidie mane vota populus offerebat
EXOD|36|4|unde artifices venire conpulsi
EXOD|36|5|dixerunt Mosi plus offert populus quam necessarium est
EXOD|36|6|iussit ergo Moses praeconis voce cantari nec vir nec mulier quicquam ultra offerat in opere sanctuarii sicque cessatum est a muneribus offerendis
EXOD|36|7|eo quod oblata sufficerent et superabundarent
EXOD|36|8|feceruntque omnes corde sapientes ad explendum opus tabernaculi cortinas decem de bysso retorta et hyacintho et purpura coccoque bis tincto opere vario et arte polymita
EXOD|36|9|quarum una habebat in longitudine viginti octo cubitos et in latitudine quattuor una mensura erat omnium cortinarum
EXOD|36|10|coniunxitque cortinas quinque alteram alteri et alias quinque sibi invicem copulavit
EXOD|36|11|fecit et ansas hyacinthinas in ora cortinae unius ex utroque latere et in ora cortinae alterius similiter
EXOD|36|12|ut contra se invicem venirent ansae et mutuo iungerentur
EXOD|36|13|unde et quinquaginta fudit circulos aureos qui morderent cortinarum ansas et fieret unum tabernaculum
EXOD|36|14|fecit et saga undecim de pilis caprarum ad operiendum tectum tabernaculi
EXOD|36|15|unum sagum habebat in longitudine cubitos triginta et in latitudine cubitos quattuor unius mensurae erant omnia saga
EXOD|36|16|quorum quinque iunxit seorsum et sex alia separatim
EXOD|36|17|fecitque ansas quinquaginta in ora sagi unius et quinquaginta in ora sagi alterius ut sibi invicem iungerentur
EXOD|36|18|et fibulas aeneas quinquaginta quibus necteretur tectum et unum pallium ex omnibus sagis fieret
EXOD|36|19|fecit et opertorium tabernaculi de pellibus arietum rubricatis aliudque desuper velamentum de pellibus ianthinis
EXOD|36|20|fecit et tabulas tabernaculi de lignis setthim stantes
EXOD|36|21|decem cubitorum erat longitudo tabulae unius et unum ac semis cubitum latitudo retinebat
EXOD|36|22|binae incastraturae erant per singulas tabulas ut altera alteri iungeretur sic fecit in omnibus tabulis tabernaculi
EXOD|36|23|e quibus viginti ad plagam meridianam erant contra austrum
EXOD|36|24|cum quadraginta basibus argenteis duae bases sub una tabula ponebantur ex utraque angulorum parte ubi incastraturae laterum in angulis terminantur
EXOD|36|25|ad plagam quoque tabernaculi quae respicit ad aquilonem fecit viginti tabulas
EXOD|36|26|cum quadraginta argenteis basibus duas bases per singulas tabulas
EXOD|36|27|contra occidentem vero id est ad eam partem tabernaculi quae mare respicit fecit sex tabulas
EXOD|36|28|et duas alias per singulos angulos tabernaculi retro
EXOD|36|29|quae iunctae erant deorsum usque sursum et in unam conpagem pariter ferebantur ita fecit ex utraque parte per angulos
EXOD|36|30|ut octo essent simul tabulae et haberent bases argenteas sedecim binas scilicet bases sub singulis tabulis
EXOD|36|31|fecit et vectes de lignis setthim quinque ad continendas tabulas unius lateris tabernaculi
EXOD|36|32|et quinque alios ad alterius lateris tabulas coaptandas et extra hos quinque alios vectes ad occidentalem plagam tabernaculi contra mare
EXOD|36|33|fecit quoque vectem alium qui per medias tabulas ab angulo usque ad angulum perveniret
EXOD|36|34|ipsa autem tabulata deauravit et circulos eorum fecit aureos per quos vectes induci possint quos et ipsos aureis lamminis operuit
EXOD|36|35|fecit et velum de hyacintho purpura vermiculo ac bysso retorta opere polymitario varium atque distinctum
EXOD|36|36|et quattuor columnas de lignis setthim quas cum capitibus deauravit fusis basibus earum argenteis
EXOD|36|37|fecit et tentorium in introitu tabernaculi ex hyacintho purpura vermiculo byssoque retorta opere plumarii
EXOD|36|38|et columnas quinque cum capitibus suis quas operuit auro basesque earum fudit aeneas
EXOD|37|1|fecit autem Beselehel et arcam de lignis setthim habentem duos semis cubitos in longitudinem et cubitum ac semissem in latitudinem altitudo quoque uno cubito fuit et dimidio vestivitque eam auro purissimo intus ac foris
EXOD|37|2|et fecit illi coronam auream per gyrum
EXOD|37|3|conflans quattuor anulos aureos per quattuor angulos eius duos anulos in latere uno et duos in altero
EXOD|37|4|vectes quoque fecit de lignis setthim quos vestivit auro
EXOD|37|5|et quos misit in anulos qui erant in lateribus arcae ad portandum eam
EXOD|37|6|fecit et propitiatorium id est oraculum de auro mundissimo duorum cubitorum et dimidio in longitudine et cubito ac semisse in latitudine
EXOD|37|7|duos etiam cherubin ex auro ductili quos posuit ex utraque parte propitiatorii
EXOD|37|8|cherub unum in summitate huius partis et cherub alterum in summitate partis alterius duos cherubin in singulis summitatibus propitiatorii
EXOD|37|9|extendentes alas et tegentes propitiatorium seque mutuo et illud respectantes
EXOD|37|10|fecit et mensam de lignis setthim in longitudine duorum cubitorum et in latitudine unius cubiti quae habebat in altitudine cubitum ac semissem
EXOD|37|11|circumdeditque eam auro mundissimo et fecit illi labium aureum per gyrum
EXOD|37|12|ipsique labio coronam interrasilem quattuor digitorum et super eandem alteram coronam auream
EXOD|37|13|fudit et quattuor circulos aureos quos posuit in quattuor angulis per singulos pedes mensae
EXOD|37|14|contra coronam misitque in eos vectes ut possit mensa portari
EXOD|37|15|ipsos quoque vectes fecit de lignis setthim et circumdedit eos auro
EXOD|37|16|et vasa ad diversos usus mensae acetabula fialas cyatos et turibula ex auro puro in quibus offerenda sunt liba
EXOD|37|17|fecit et candelabrum ductile de auro mundissimo de cuius vecte calami scyphi spherulae ac lilia procedebant
EXOD|37|18|sex in utroque latere tres calami ex parte una et tres ex altera
EXOD|37|19|tres scyphi in nucis modum per calamos singulos spherulaeque simul et lilia et tres scyphi instar nucis in calamo altero spherulaeque simul et lilia aequum erat opus sex calamorum qui procedebant de stipite candelabri
EXOD|37|20|in ipso autem vecte erant quattuor scyphi in nucis modum spherulaeque per singulos et lilia
EXOD|37|21|et spherae sub duobus calamis per loca tria qui simul sex fiunt calami procedentes de vecte uno
EXOD|37|22|et spherae igitur et calami ex ipso erant universa ductilia de auro purissimo
EXOD|37|23|fecit et lucernas septem cum emunctoriis suis et vasa ubi quae emuncta sunt extinguuntur de auro mundissimo
EXOD|37|24|talentum auri adpendebat candelabrum cum omnibus vasis suis
EXOD|37|25|fecit et altare thymiamatis de lignis setthim habens per quadrum singulos cubitos et in altitudine duos e cuius angulis procedebant cornua
EXOD|37|26|vestivitque illud auro purissimo cum craticula ac parietibus et cornibus
EXOD|37|27|fecitque ei coronam aureolam per gyrum et duos anulos aureos sub corona per singula latera ut mittantur in eos vectes et possit altare portari
EXOD|37|28|ipsos autem vectes fecit de lignis setthim et operuit lamminis aureis
EXOD|37|29|conposuit et oleum ad sanctificationis unguentum et thymiama de aromatibus mundissimis opere pigmentarii
EXOD|38|1|fecit et altare holocausti de lignis setthim quinque cubitorum per quadrum et trium in altitudine
EXOD|38|2|cuius cornua de angulis procedebant operuitque illud aeneis lamminis
EXOD|38|3|et in usus eius paravit ex aere vasa diversa lebetas forcipes fuscinulas uncinos et ignium receptacula
EXOD|38|4|craticulamque eius in modum retis fecit aeneam et subter eam in altaris medio arulam
EXOD|38|5|fusis quattuor anulis per totidem retiaculi summitates ad inmittendos vectes ad portandum
EXOD|38|6|quos et ipsos fecit de lignis setthim et operuit lamminis aeneis
EXOD|38|7|induxitque in circulos qui in altaris lateribus eminebant ipsum autem altare non erat solidum sed cavum ex tabulis et intus vacuum
EXOD|38|8|fecit et labrum aeneum cum base sua de speculis mulierum quae excubabant in ostio tabernaculi
EXOD|38|9|et atrium in cuius australi plaga erant tentoria de bysso retorta cubitorum centum
EXOD|38|10|columnae aeneae viginti cum basibus suis capita columnarum et tota operis celatura argentea
EXOD|38|11|aeque ad septentrionalis plagam tentoria columnae basesque et capita columnarum eiusdem et mensurae et operis ac metalli erant
EXOD|38|12|in ea vero plaga quae occidentem respicit fuere tentoria cubitorum quinquaginta columnae decem cum basibus suis aeneae et capita columnarum celata argentea
EXOD|38|13|porro contra orientem quinquaginta cubitorum paravit tentoria
EXOD|38|14|e quibus quindecim cubitos columnarum trium cum basibus suis unum tenebat latus
EXOD|38|15|et in parte altera quia utraque introitum tabernaculi facit quindecim aeque cubitorum erant tentoria columnae tres et bases totidem
EXOD|38|16|cuncta atrii tentoria byssus torta texuerat
EXOD|38|17|bases columnarum fuere aeneae capita autem earum cum celaturis suis argentea sed et ipsas columnas atrii vestivit argento
EXOD|38|18|et in introitu eius opere plumario fecit tentorium ex hyacintho purpura vermiculo ac bysso retorta quod habebat viginti cubitos in longitudine altitudo vero quinque cubitorum erat iuxta mensuram quam cuncta atrii habebant tentoria
EXOD|38|19|columnae autem ingressus fuere quattuor cum basibus aeneis capitaque earum et celaturae argenteae
EXOD|38|20|paxillos quoque tabernaculi et atrii per gyrum fecit aeneos
EXOD|38|21|haec sunt instrumenta tabernaculi testimonii quae numerata sunt iuxta praeceptum Mosi in caerimonias Levitarum per manum Ithamar filii Aaron sacerdotis
EXOD|38|22|quas Beselehel filius Uri filii Hur de tribu Iuda Domino per Mosen iubente conpleverat
EXOD|38|23|iuncto sibi socio Hooliab filio Achisamech de tribu Dan qui et ipse artifex lignorum egregius fuit et polymitarius atque plumarius ex hyacintho purpura vermiculo et bysso
EXOD|38|24|omne aurum quod expensum est in opere sanctuarii et quod oblatum in donariis viginti novem talentorum fuit et septingentorum triginta siclorum ad mensuram sanctuarii
EXOD|38|25|oblatum est autem ab his qui transierant ad numerum a viginti annis et supra de sescentis tribus milibus et quingentis quinquaginta armatorum
EXOD|38|26|fuerunt praeterea centum talenta argenti e quibus conflatae sunt bases sanctuarii et introitus ubi velum pendet
EXOD|38|27|centum bases factae sunt de talentis centum singulis talentis per bases singulas supputatis
EXOD|38|28|de mille autem septingentis et septuaginta quinque fecit capita columnarum quas et ipsas vestivit argento
EXOD|38|29|aeris quoque oblata sunt talenta septuaginta duo milia et quadringenti supra sicli
EXOD|38|30|ex quibus fusae sunt bases in introitu tabernaculi testimonii et altare aeneum cum craticula sua omniaque vasa quae ad usum eius pertinent
EXOD|38|31|et bases atrii tam in circuitu quam in ingressu eius et paxilli tabernaculi atque atrii per gyrum
EXOD|39|1|de hyacintho vero et purpura vermiculo ac bysso fecit vestes quibus indueretur Aaron quando ministrabat in sanctis sicut praecepit Dominus Mosi
EXOD|39|2|fecit igitur superumerale de auro hyacintho et purpura coccoque bis tincto et bysso retorta
EXOD|39|3|opere polymitario inciditque bratteas aureas et extenuavit in fila ut possint torqueri cum priorum colorum subtemine
EXOD|39|4|duasque oras sibi invicem copulatas in utroque latere summitatum
EXOD|39|5|et balteum ex hisdem coloribus sicut praeceperat Dominus Mosi
EXOD|39|6|paravit et duos lapides onychinos adstrictos et inclusos auro et sculptos arte gemmaria nominibus filiorum Israhel
EXOD|39|7|posuitque eos in lateribus superumeralis in monumentum filiorum Israhel sicut praeceperat Dominus Mosi
EXOD|39|8|fecit et rationale opere polymito iuxta opus superumeralis ex auro hyacintho purpura coccoque bis tincto et bysso retorta
EXOD|39|9|quadrangulum duplex mensurae palmi
EXOD|39|10|et posuit in eo gemmarum ordines quattuor in primo versu erat sardius topazius zmaragdus
EXOD|39|11|in secundo carbunculus sapphyrus iaspis
EXOD|39|12|in tertio ligyrius achates amethistus
EXOD|39|13|in quarto chrysolitus onychinus berillus circumdati et inclusi auro per ordines suos
EXOD|39|14|ipsique lapides duodecim sculpti erant nominibus duodecim tribuum Israhel singuli per nomina singulorum
EXOD|39|15|fecerunt in rationali et catenulas sibi invicem coherentes de auro purissimo
EXOD|39|16|et duos uncinos totidemque anulos aureos porro anulos posuerunt in utroque latere rationalis
EXOD|39|17|e quibus penderent duae catenae aureae quas inseruerunt uncinis qui in superumeralis angulis eminebant
EXOD|39|18|haec et ante et retro ita conveniebant sibi ut superumerale et rationale mutuo necterentur
EXOD|39|19|stricta ad balteum et anulis fortius copulata quos iungebat vitta hyacinthina ne laxe fluerent et a se invicem moverentur sicut praecepit Dominus Mosi
EXOD|39|20|fecerunt quoque tunicam superumeralis totam hyacinthinam
EXOD|39|21|et capitium in superiori parte contra medium oramque per gyrum capitii textilem
EXOD|39|22|deorsum autem ad pedes mala punica ex hyacintho purpura vermiculo ac bysso retorta
EXOD|39|23|et tintinabula de auro mundissimo quae posuerunt inter mala granata in extrema parte tunicae per gyrum
EXOD|39|24|tintinabulum aureum et malum punicum quibus ornatus incedebat pontifex quando ministerio fungebatur sicut praecepit Dominus Mosi
EXOD|39|25|fecerunt et tunicas byssinas opere textili Aaron et filiis eius
EXOD|39|26|et mitras cum coronulis suis ex bysso
EXOD|39|27|feminalia quoque linea byssina
EXOD|39|28|cingulum vero de bysso retorta hyacintho purpura ac vermiculo distinctum arte plumaria sicut praecepit Dominus Mosi
EXOD|39|29|fecerunt et lamminam sacrae venerationis de auro purissimo scripseruntque in ea opere gemmario Sanctum Domini
EXOD|39|30|et strinxerunt eam cum mitra vitta hyacinthina sicut praecepit Dominus Mosi
EXOD|39|31|perfectum est igitur omne opus tabernaculi et tecti testimonii feceruntque filii Israhel cuncta quae praeceperat Dominus Mosi
EXOD|39|32|et obtulerunt tabernaculum et tectum et universam supellectilem anulos tabulas vectes columnas ac bases
EXOD|39|33|opertorium de pellibus arietum rubricatis et aliud operimentum de ianthinis pellibus
EXOD|39|34|velum arcam vectes propitiatorium
EXOD|39|35|mensam cum vasis et propositionis panibus
EXOD|39|36|candelabrum lucernas et utensilia eorum cum oleo
EXOD|39|37|altare aureum et unguentum thymiama ex aromatibus
EXOD|39|38|et tentorium in introitu tabernaculi
EXOD|39|39|altare aeneum retiaculum vectes et vasa eius omnia labrum cum basi sua tentoria atrii et columnas cum basibus suis
EXOD|39|40|tentorium in introitu atrii funiculosque illius et paxillos nihil ex vasis defuit quae in ministerium tabernaculi et in tectum foederis iussa sunt fieri
EXOD|39|41|vestes quoque quibus sacerdotes utuntur in sanctuario Aaron scilicet et filii eius
EXOD|39|42|obtulerunt filii Israhel sicut praeceperat Dominus
EXOD|39|43|quae postquam Moses cuncta vidit expleta benedixit eis
EXOD|40|1|locutusque est Dominus ad Mosen dicens
EXOD|40|2|mense primo die prima mensis eriges tabernaculum testimonii
EXOD|40|3|et pones in eo arcam dimittesque ante illam velum
EXOD|40|4|et inlata mensa pones super eam quae rite praecepta sunt candelabrum stabit cum lucernis suis
EXOD|40|5|et altare aureum in quo adoletur incensum coram arca testimonii tentorium in introitu tabernaculi pones
EXOD|40|6|et ante illud altare holocausti
EXOD|40|7|labrum inter altare et tabernaculum quod implebis aqua
EXOD|40|8|circumdabisque atrium tentoriis et ingressum eius
EXOD|40|9|et adsumpto unctionis oleo ungues tabernaculum cum vasis suis ut sanctificentur
EXOD|40|10|altare holocausti et omnia vasa eius
EXOD|40|11|labrum cum basi sua omnia unctionis oleo consecrabis ut sint sancta sanctorum
EXOD|40|12|adplicabisque Aaron et filios eius ad fores tabernaculi testimonii et lotos aqua
EXOD|40|13|indues sanctis vestibus ut ministrent mihi et unctio eorum in sacerdotium proficiat sempiternum
EXOD|40|14|fecitque Moses omnia quae praeceperat Dominus
EXOD|40|15|igitur mense primo anni secundi in prima die mensis conlocatum est tabernaculum
EXOD|40|16|erexitque illud Moses et posuit tabulas ac bases et vectes statuitque columnas
EXOD|40|17|et expandit tectum super tabernaculum inposito desuper operimento sicut Dominus imperarat
EXOD|40|18|posuit et testimonium in arca subditis infra vectibus et oraculum desuper
EXOD|40|19|cumque intulisset arcam in tabernaculum adpendit ante eam velum ut expleret Domini iussionem
EXOD|40|20|posuit et mensam in tabernaculo testimonii ad plagam septentrionalem extra velum
EXOD|40|21|ordinatis coram propositionis panibus sicut praeceperat Dominus Mosi
EXOD|40|22|posuit et candelabrum in tabernaculum testimonii e regione mensae in parte australi
EXOD|40|23|locatis per ordinem lucernis iuxta praeceptum Domini
EXOD|40|24|posuit et altare aureum sub tecto testimonii contra velum
EXOD|40|25|et adolevit super eo incensum aromatum sicut iusserat Dominus
EXOD|40|26|posuit et tentorium in introitu tabernaculi
EXOD|40|27|et altare holocausti in vestibulo testimonii offerens in eo holocaustum et sacrificia ut Dominus imperarat
EXOD|40|28|labrum quoque statuit inter tabernaculum testimonii et altare implens illud aqua
EXOD|40|29|laveruntque Moses et Aaron ac filii eius manus suas et pedes
EXOD|40|30|cum ingrederentur tectum foederis et accederent ad altare sicut praeceperat Dominus
EXOD|40|31|erexit et atrium per gyrum tabernaculi et altaris ducto in introitu eius tentorio postquam cuncta perfecta sunt
EXOD|40|32|operuit nubes tabernaculum testimonii et gloria Domini implevit illud
EXOD|40|33|nec poterat Moses ingredi tectum foederis nube operiente omnia et maiestate Domini coruscante quia cuncta nubes operuerat
EXOD|40|34|si quando nubes tabernaculum deserebat proficiscebantur filii Israhel per turmas suas
EXOD|40|35|si pendebat desuper manebant in eodem loco
EXOD|40|36|nubes quippe Domini incubabat per diem tabernaculo et ignis in nocte videntibus populis Israhel per cunctas mansiones suas
LEV|1|1|vocavit autem Mosen et locutus est ei Dominus de tabernaculo testimonii dicens
LEV|1|2|loquere filiis Israhel et dices ad eos homo qui obtulerit ex vobis hostiam Domino de pecoribus id est de bubus et ovibus offerens victimas
LEV|1|3|si holocaustum fuerit eius oblatio ac de armento masculum inmaculatum offeret ad ostium tabernaculi testimonii ad placandum sibi Dominum
LEV|1|4|ponetque manus super caput hostiae et acceptabilis erit atque in expiationem eius proficiens
LEV|1|5|immolabitque vitulum coram Domino et offerent filii Aaron sacerdotes sanguinem eius fundentes super altaris circuitum quod est ante ostium tabernaculi
LEV|1|6|detractaque pelle hostiae artus in frusta concident
LEV|1|7|et subicient in altari ignem strue lignorum ante conposita
LEV|1|8|et membra quae caesa sunt desuper ordinantes caput videlicet et cuncta quae adherent iecori
LEV|1|9|intestinis et pedibus lotis aqua adolebitque ea sacerdos super altare in holocaustum et suavem odorem Domino
LEV|1|10|quod si de pecoribus oblatio est de ovibus sive de capris holocaustum anniculum et absque macula offeret
LEV|1|11|immolabitque ad latus altaris quod respicit ad aquilonem coram Domino sanguinem vero illius fundent super altare filii Aaron per circuitum
LEV|1|12|dividentque membra caput et omnia quae adherent iecori et inponent super ligna quibus subiciendus est ignis
LEV|1|13|intestina vero et pedes lavabunt aqua et oblata omnia adolebit sacerdos super altare in holocaustum et odorem suavissimum Domino
LEV|1|14|sin autem de avibus holocausti oblatio fuerit Domino de turturibus et pullis columbae
LEV|1|15|offeret eam sacerdos ad altare et retorto ad collum capite ac rupto vulneris loco decurrere faciet sanguinem super crepidinem altaris
LEV|1|16|vesiculam vero gutturis et plumas proiciet propter altare ad orientalem plagam in loco in quo cineres effundi solent
LEV|1|17|confringetque ascellas eius et non secabit nec ferro dividet eam et adolebit super altare lignis igne subposito holocaustum est et oblatio suavissimi odoris Domino
LEV|2|1|anima cum obtulerit oblationem sacrificii Domino simila erit eius oblatio fundetque super eam oleum et ponet tus
LEV|2|2|ac deferet ad filios Aaron sacerdotes quorum unus tollet pugillum plenum similae et olei ac totum tus et ponet memoriale super altare in odorem suavissimum Domino
LEV|2|3|quod autem reliquum fuerit de sacrificio erit Aaron et filiorum eius sanctum sanctorum de oblationibus Domini
LEV|2|4|cum autem obtuleris sacrificium coctum in clibano de simila panes scilicet absque fermento conspersos oleo et lagana azyma oleo lita
LEV|2|5|si oblatio tua fuerit de sartagine similae conspersae oleo et absque fermento
LEV|2|6|divides eam minutatim et fundes supra oleum
LEV|2|7|sin autem de craticula sacrificium aeque simila oleo conspergetur
LEV|2|8|quam offeres Domino tradens manibus sacerdotis
LEV|2|9|qui cum obtulerit eam tollet memoriale de sacrificio et adolebit super altare in odorem suavitatis Domino
LEV|2|10|quicquid autem reliquum est erit Aaron et filiorum eius sanctum sanctorum de oblationibus Domini
LEV|2|11|omnis oblatio quae offertur Domino absque fermento fiet nec quicquam fermenti ac mellis adolebitur in sacrificio Domini
LEV|2|12|primitias tantum eorum offeretis et munera super altare vero non ponentur in odorem suavitatis
LEV|2|13|quicquid obtuleris sacrificii sale condies nec auferes sal foederis Dei tui de sacrificio tuo in omni oblatione offeres sal
LEV|2|14|sin autem obtuleris munus primarum frugum tuarum Domino de spicis adhuc virentibus torres eas igni et confringes in morem farris et sic offeres primitias tuas Domino
LEV|2|15|fundens supra oleum et tus inponens quia oblatio Domini est
LEV|2|16|de qua adolebit sacerdos in memoriam muneris partem farris fracti et olei ac totum tus
LEV|3|1|quod si hostia pacificorum fuerit eius oblatio et de bubus voluerit offerre marem sive feminam inmaculata offeret coram Domino
LEV|3|2|ponetque manum super caput victimae suae quae immolabitur in introitu tabernaculi fundentque filii Aaron sacerdotes sanguinem per circuitum altaris
LEV|3|3|et offerent de hostia pacificorum in oblationem Domini adipem qui operit vitalia et quicquid pinguedinis intrinsecus est
LEV|3|4|duos renes cum adipe quo teguntur ilia et reticulum iecoris cum renunculis
LEV|3|5|adolebuntque ea super altare in holocaustum lignis igne subposito in oblationem suavissimi odoris Domino
LEV|3|6|si vero de ovibus fuerit eius oblatio et pacificorum hostia sive masculum sive feminam obtulerit inmaculata erunt
LEV|3|7|si agnum obtulerit coram Domino
LEV|3|8|ponet manum super caput victimae suae quae immolabitur in vestibulo tabernaculi testimonii fundentque filii Aaron sanguinem eius per altaris circuitum
LEV|3|9|et offerent de pacificorum hostia sacrificium Domino adipem et caudam totam
LEV|3|10|cum renibus et pinguedinem quae operit ventrem atque universa vitalia et utrumque renunculum cum adipe qui est iuxta ilia reticulumque iecoris cum renunculis
LEV|3|11|et adolebit ea sacerdos super altare in pabulum ignis et oblationis Domini
LEV|3|12|si capra fuerit eius oblatio et obtulerit eam Domino
LEV|3|13|ponet manum suam super caput eius immolabitque eam in introitu tabernaculi testimonii et fundent filii Aaron sanguinem eius per altaris circuitum
LEV|3|14|tollentque ex ea in pastum ignis dominici adipem qui operit ventrem et qui tegit universa vitalia
LEV|3|15|duos renunculos cum reticulo qui est super eos iuxta ilia et arvinam iecoris cum renunculis
LEV|3|16|adolebitque ea sacerdos super altare in alimoniam ignis et suavissimi odoris omnis adeps Domini erit
LEV|3|17|iure perpetuo in generationibus et cunctis habitaculis vestris nec adipes nec sanguinem omnino comedetis
LEV|4|1|locutusque est Dominus ad Mosen dicens
LEV|4|2|loquere filiis Israhel anima cum peccaverit per ignorantiam et de universis mandatis Domini quae praecepit ut non fierent quippiam fecerit
LEV|4|3|si sacerdos qui est unctus peccaverit delinquere faciens populum offeret pro peccato suo vitulum inmaculatum Domino
LEV|4|4|et adducet illum ad ostium tabernaculi testimonii coram Domino ponetque manum super caput eius et immolabit eum Domino
LEV|4|5|hauriet quoque de sanguine vituli inferens illud in tabernaculum testimonii
LEV|4|6|cumque intinxerit digitum in sanguinem asperget eo septies coram Domino contra velum sanctuarii
LEV|4|7|ponetque de eodem sanguine super cornua altaris thymiamatis gratissimi Domino quod est in tabernaculo testimonii omnem autem reliquum sanguinem fundet in basim altaris holocausti in introitu tabernaculi
LEV|4|8|et adipem vituli auferet pro peccato tam eum qui operit vitalia quam omnia quae intrinsecus sunt
LEV|4|9|duos renunculos et reticulum quod est super eos iuxta ilia et adipem iecoris cum renunculis
LEV|4|10|sicut aufertur de vitulo hostiae pacificorum et adolebit ea super altare holocausti
LEV|4|11|pellem vero et omnes carnes cum capite et pedibus et intestinis et fimo
LEV|4|12|et reliquo corpore efferet extra castra in locum mundum ubi cineres effundi solent incendetque ea super lignorum struem quae in loco effusorum cinerum cremabuntur
LEV|4|13|quod si omnis turba Israhel ignoraverit et per inperitiam fecerit quod contra mandatum Domini est
LEV|4|14|et postea intellexerit peccatum suum offeret vitulum pro peccato adducetque eum ad ostium tabernaculi
LEV|4|15|et ponent seniores populi manus super caput eius coram Domino immolatoque vitulo in conspectu Domini
LEV|4|16|inferet sacerdos qui unctus est de sanguine eius in tabernaculum testimonii
LEV|4|17|tincto digito aspergens septies contra velum
LEV|4|18|ponetque de eodem sanguine in cornibus altaris quod est coram Domino in tabernaculo testimonii reliquum autem sanguinem fundet iuxta basim altaris holocaustorum quod est in ostio tabernaculi testimonii
LEV|4|19|omnemque eius adipem tollet et adolebit super altare
LEV|4|20|sic faciens et de hoc vitulo quomodo fecit et prius et rogante pro eis sacerdote propitius erit Dominus
LEV|4|21|ipsum autem vitulum efferet extra castra atque conburet sicut et priorem vitulum quia pro peccato est multitudinis
LEV|4|22|si peccaverit princeps et fecerit unum e pluribus per ignorantiam quod Domini lege prohibetur
LEV|4|23|et postea intellexerit peccatum suum offeret hostiam Domino hircum de capris inmaculatum
LEV|4|24|ponetque manum suam super caput eius cumque immolaverit eum in loco ubi solet mactari holocaustum coram Domino quia pro peccato est
LEV|4|25|tinguet sacerdos digitum in sanguine hostiae pro peccato tangens cornua altaris holocausti et reliquum fundens ad basim eius
LEV|4|26|adipem vero adolebit supra sicut in victimis pacificorum fieri solet rogabitque pro eo et pro peccato eius ac dimittetur ei
LEV|4|27|quod si peccaverit anima per ignorantiam de populo terrae ut faciat quicquam ex his quae Domini lege prohibentur atque delinquat
LEV|4|28|et cognoverit peccatum suum offeret capram inmaculatam
LEV|4|29|ponetque manum super caput hostiae quae pro peccato est et immolabit eam in loco holocausti
LEV|4|30|tolletque sacerdos de sanguine in digito suo et tangens cornua altaris holocausti reliquum fundet ad basim eius
LEV|4|31|omnem autem auferens adipem sicut auferri solet de victimis pacificorum adolebit super altare in odorem suavitatis Domino rogabitque pro eo et dimittetur ei
LEV|4|32|sin autem de pecoribus obtulerit victimam pro peccato ovem scilicet inmaculatam
LEV|4|33|ponet manum super caput eius et immolabit eam in loco ubi solent holocaustorum caedi hostiae
LEV|4|34|sumetque sacerdos de sanguine eius digito suo et tangens cornua altaris holocausti reliquum fundet ad basim eius
LEV|4|35|omnem quoque auferens adipem sicut auferri solet adeps arietis qui immolatur pro pacificis et cremabit super altare in incensum Domini rogabitque pro eo et pro peccato eius et dimittetur illi
LEV|5|1|si peccaverit anima et audierit vocem iurantis testisque fuerit quod aut ipse vidit aut conscius est nisi indicaverit portabit iniquitatem suam
LEV|5|2|anima quae tetigerit aliquid inmundum sive quod occisum a bestia est aut per se mortuum vel quodlibet aliud reptile et oblita fuerit inmunditiae suae rea est et deliquit
LEV|5|3|et si tetigerit quicquam de inmunditia hominis iuxta omnem inpuritatem qua pollui solet oblitaque cognoverit postea subiacebit delicto
LEV|5|4|anima quae iuraverit et protulerit labiis suis ut vel male quid faceret vel bene et id ipsum iuramento et sermone firmaverit oblitaque postea intellexerit delictum suum
LEV|5|5|agat paenitentiam pro peccato
LEV|5|6|et offerat agnam de gregibus sive capram orabitque pro eo sacerdos et pro peccato eius
LEV|5|7|sin autem non potuerit offerre pecus offerat duos turtures vel duos pullos columbarum Domino unum pro peccato et alterum in holocaustum
LEV|5|8|dabitque eos sacerdoti qui primum offerens pro peccato retorquebit caput eius ad pinnulas ita ut collo hereat et non penitus abrumpatur
LEV|5|9|et asperget de sanguine eius parietem altaris quicquid autem reliquum fuerit faciet destillare ad fundamentum eius quia pro peccato est
LEV|5|10|alterum vero adolebit holocaustum ut fieri solet rogabitque pro eo sacerdos et pro peccato eius et dimittetur ei
LEV|5|11|quod si non quiverit manus eius offerre duos turtures vel duos pullos columbae offeret pro peccato similam partem oephi decimam non mittet in eam oleum nec turis aliquid inponet quia pro peccato est
LEV|5|12|tradetque eam sacerdoti qui plenum ex toto pugillum hauriens cremabit super altare in monumentum eius qui obtulit
LEV|5|13|rogans pro illo et expians reliquam vero partem ipse habebit in munere
LEV|5|14|locutus est Dominus ad Mosen dicens
LEV|5|15|anima si praevaricans caerimonias per errorem in his quae Domino sunt sanctificata peccaverit offeret pro delicto suo arietem inmaculatum de gregibus qui emi potest duobus siclis iuxta pondus sanctuarii
LEV|5|16|ipsumque quod intulit damni restituet et quintam partem ponet supra tradens sacerdoti qui rogabit pro eo offerens arietem et dimittetur ei
LEV|5|17|anima si peccaverit per ignorantiam feceritque unum ex his quae Domini lege prohibentur et peccati rea intellexerit iniquitatem suam
LEV|5|18|offeret arietem inmaculatum de gregibus sacerdoti iuxta mensuram aestimationemque peccati qui orabit pro eo quod nesciens fecerit et dimittetur ei
LEV|5|19|quia per errorem deliquit in Dominum
LEV|6|1|locutus est Dominus ad Mosen dicens
LEV|6|2|anima quae peccaverit et contempto Domino negaverit depositum proximo suo quod fidei eius creditum fuerat vel vi aliquid extorserit aut calumniam fecerit
LEV|6|3|sive rem perditam invenerit et infitians insuper peierarit et quodlibet aliud ex pluribus fecerit in quibus peccare solent homines
LEV|6|4|convicta delicti reddet
LEV|6|5|omnia quae per fraudem voluit obtinere integra et quintam insuper partem domino cui damnum intulerat
LEV|6|6|pro peccato autem suo offeret arietem inmaculatum de grege et dabit eum sacerdoti iuxta aestimationem mensuramque delicti
LEV|6|7|qui rogabit pro eo coram Domino et dimittetur illi pro singulis quae faciendo peccaverit
LEV|6|8|locutus est Dominus ad Mosen dicens
LEV|6|9|praecipe Aaron et filiis eius haec est lex holocausti cremabitur in altari tota nocte usque mane ignis ex eodem altari erit
LEV|6|10|vestietur sacerdos tunica et feminalibus lineis tolletque cineres quos vorans ignis exusit et ponens iuxta altare
LEV|6|11|spoliabitur prioribus vestimentis indutusque aliis efferet eos extra castra et in loco mundissimo usque ad favillam consumi faciet
LEV|6|12|ignis autem in altari semper ardebit quem nutriet sacerdos subiciens ligna mane per singulos dies et inposito holocausto desuper adolebit adipes pacificorum
LEV|6|13|ignis est iste perpetuus qui numquam deficiet in altari
LEV|6|14|haec est lex sacrificii et libamentorum quae offerent filii Aaron coram Domino et coram altari
LEV|6|15|tollet sacerdos pugillum similae quae conspersa est oleo et totum tus quod super similam positum est adolebitque illud in altari in monumentum odoris suavissimi Domino
LEV|6|16|reliquam autem partem similae comedet Aaron cum filiis suis absque fermento et comedet in loco sancto atrii tabernaculi
LEV|6|17|ideo autem non fermentabitur quia pars eius in Domini offertur incensum sanctum sanctorum erit sicut pro peccato atque delicto
LEV|6|18|mares tantum stirpis Aaron comedent illud legitimum ac sempiternum est in generationibus vestris de sacrificiis Domini omnis qui tetigerit illa sanctificabitur
LEV|6|19|et locutus est Dominus ad Mosen dicens
LEV|6|20|haec est oblatio Aaron et filiorum eius quam offerre debent Domino in die unctionis suae decimam partem oephi offerent similae in sacrificio sempiterno medium eius mane et medium vespere
LEV|6|21|quae in sartagine oleo conspersa frigetur offeret autem eam calidam in odorem suavissimum Domino
LEV|6|22|sacerdos qui patri iure successerit et tota cremabitur in altari
LEV|6|23|omne enim sacrificium sacerdotum igne consumetur nec quisquam comedet ex eo
LEV|6|24|locutus est Dominus ad Mosen dicens
LEV|6|25|loquere Aaron et filiis eius ista est lex hostiae pro peccato in loco ubi offertur holocaustum immolabitur coram Domino sanctum sanctorum est
LEV|6|26|sacerdos qui offert comedet eam in loco sancto in atrio tabernaculi
LEV|6|27|quicquid tetigerit carnes eius sanctificabitur si de sanguine illius vestis fuerit aspersa lavabitur in loco sancto
LEV|6|28|vas autem fictile in quo cocta est confringetur quod si vas aeneum fuerit defricabitur et lavabitur aqua
LEV|6|29|omnis masculus de genere sacerdotali vescetur carnibus eius quia sanctum sanctorum est
LEV|6|30|hostia enim quae caeditur pro peccato cuius sanguis infertur in tabernaculum testimonii ad expiandum in sanctuario non comedetur sed conburetur igni
LEV|7|1|haec quoque est lex hostiae pro delicto sancta sanctorum est
LEV|7|2|idcirco ubi immolatur holocaustum mactabitur et victima pro delicto sanguis eius per gyrum fundetur altaris
LEV|7|3|offerent ex ea caudam et adipem qui operit vitalia
LEV|7|4|duos renunculos et pinguedinem quae iuxta ilia est reticulumque iecoris cum renunculis
LEV|7|5|et adolebit ea sacerdos super altare incensum est Domini pro delicto
LEV|7|6|omnis masculus de sacerdotali genere in loco sancto vescetur his carnibus quia sanctum sanctorum est
LEV|7|7|sicut pro peccato offertur hostia ita et pro delicto utriusque hostiae lex una erit ad sacerdotem qui eam obtulerit pertinebit
LEV|7|8|sacerdos qui offert holocausti victimam habebit pellem eius
LEV|7|9|et omne sacrificium similae quod coquitur in clibano et quicquid in craticula vel in sartagine praeparatur eius erit sacerdotis a quo offertur
LEV|7|10|sive oleo conspersa sive arida fuerit cunctis filiis Aaron aequa mensura per singulos dividetur
LEV|7|11|haec est lex hostiae pacificorum quae offertur Domino
LEV|7|12|si pro gratiarum actione fuerit oblatio offerent panes absque fermento conspersos oleo et lagana azyma uncta oleo coctamque similam et collyridas olei admixtione conspersas
LEV|7|13|panes quoque fermentatos cum hostia gratiarum quae immolatur pro pacificis
LEV|7|14|ex quibus unus pro primitiis offeretur Domino et erit sacerdotis qui fundet hostiae sanguinem
LEV|7|15|cuius carnes eadem comedentur die nec remanebit ex eis quicquam usque mane
LEV|7|16|si voto vel sponte quisquam obtulerit hostiam eadem similiter edetur die sed et si quid in crastinum remanserit vesci licitum est
LEV|7|17|quicquid autem tertius invenerit dies ignis absumet
LEV|7|18|si quis de carnibus victimae pacificorum die tertio comederit irrita fiet oblatio nec proderit offerenti quin potius quaecumque anima tali se edulio contaminarit praevaricationis rea erit
LEV|7|19|caro quae aliquid tetigerit inmundum non comedetur sed conburetur igni qui fuerit mundus vescetur ea
LEV|7|20|anima polluta quae ederit de carnibus hostiae pacificorum quae oblata est Domino peribit de populis suis
LEV|7|21|et quae tetigerit inmunditiam hominis vel iumenti sive omnis rei quae polluere potest et comederit de huiuscemodi carnibus interibit de populis suis
LEV|7|22|locutusque est Dominus ad Mosen dicens
LEV|7|23|loquere filiis Israhel adipem bovis et ovis et caprae non comedetis
LEV|7|24|adipem cadaveris morticini et eius animalis quod a bestia captum est habebitis in usus varios
LEV|7|25|si quis adipem qui offerri debet in incensum Domini comederit peribit de populo suo
LEV|7|26|sanguinem quoque omnis animalis non sumetis in cibo tam de avibus quam de pecoribus
LEV|7|27|omnis anima quae ederit sanguinem peribit de populis suis
LEV|7|28|locutus est Dominus ad Mosen dicens
LEV|7|29|loquere filiis Israhel qui offert victimam pacificorum Domino offerat simul et sacrificium id est libamenta eius
LEV|7|30|tenebit manibus adipem hostiae et pectusculum cumque ambo oblata Domino consecrarit tradet sacerdoti
LEV|7|31|qui adolebit adipem super altare pectusculum autem erit Aaron et filiorum eius
LEV|7|32|armus quoque dexter de pacificorum hostiis cedet in primitias sacerdotis
LEV|7|33|qui obtulerit sanguinem et adipem filiorum Aaron ipse habebit et armum dextrum in portione sua
LEV|7|34|pectusculum enim elationis et armum separationis tuli a filiis Israhel de hostiis eorum pacificis et dedi Aaron sacerdoti ac filiis eius lege perpetua ab omni populo Israhel
LEV|7|35|haec est unctio Aaron et filiorum eius in caerimoniis Domini die qua obtulit eos Moses ut sacerdotio fungerentur
LEV|7|36|et quae praecepit dari eis Dominus a filiis Israhel religione perpetua in generationibus suis
LEV|7|37|ista est lex holocausti et sacrificii pro peccato atque delicto et pro consecratione et pacificorum victimis
LEV|7|38|quas constituit Dominus Mosi in monte Sinai quando mandavit filiis Israhel ut offerrent oblationes suas Domino in deserto Sinai
LEV|8|1|locutusque est Dominus ad Mosen dicens
LEV|8|2|tolle Aaron cum filiis suis vestes eorum et unctionis oleum vitulum pro peccato duos arietes canistrum cum azymis
LEV|8|3|et congregabis omnem coetum ad ostium tabernaculi
LEV|8|4|fecit Moses ut Dominus imperarat congregataque omni turba ante fores
LEV|8|5|ait iste est sermo quem iussit Dominus fieri
LEV|8|6|statimque obtulit Aaron et filios eius cumque lavisset eos
LEV|8|7|vestivit pontificem subucula linea accingens eum balteo et induens tunica hyacinthina et desuper umerale inposuit
LEV|8|8|quod adstringens cingulo aptavit rationali in quo erat doctrina et veritas
LEV|8|9|cidarim quoque texit caput et super eam contra frontem posuit lamminam auream consecratam in sanctificationem sicut praeceperat ei Dominus
LEV|8|10|tulit et unctionis oleum quo levit tabernaculum cum omni supellectili sua
LEV|8|11|cumque sanctificans aspersisset altare septem vicibus unxit illud et omnia vasa eius labrumque cum basi sua sanctificavit oleo
LEV|8|12|quod fundens super caput Aaron unxit eum et consecravit
LEV|8|13|filios quoque eius oblatos vestivit tunicis lineis et cinxit balteo inposuitque mitras ut iusserat Dominus
LEV|8|14|obtulit et vitulum pro peccato cumque super caput eius posuissent Aaron et filii eius manus suas
LEV|8|15|immolavit eum hauriens sanguinem et tincto digito tetigit cornua altaris per gyrum quo expiato et sanctificato fudit reliquum sanguinem ad fundamenta eius
LEV|8|16|adipem autem qui erat super vitalia et reticulum iecoris duosque renunculos cum arvinulis suis adolevit super altare
LEV|8|17|vitulum cum pelle carnibus et fimo cremans extra castra sicut praeceperat Dominus
LEV|8|18|obtulit et arietem in holocaustum super cuius caput cum inposuissent Aaron et filii eius manus suas
LEV|8|19|immolavit eum et fudit sanguinem eius per altaris circuitum
LEV|8|20|ipsumque arietem in frusta concidens caput eius et artus et adipem adolevit igni
LEV|8|21|lotis prius intestinis et pedibus totumque simul arietem incendit super altare eo quod esset holocaustum suavissimi odoris Domino sicut praeceperat ei
LEV|8|22|obtulit et arietem secundum in consecrationem sacerdotum posueruntque super caput illius Aaron et filii eius manus suas
LEV|8|23|quem cum immolasset Moses sumens de sanguine tetigit extremum auriculae dextrae Aaron et pollicem manus eius dextrae similiter et pedis
LEV|8|24|obtulit et filios Aaron cumque de sanguine arietis immolati tetigisset extremum auriculae singulorum dextrae et pollices manus ac pedis dextri reliquum fudit super altare per circuitum
LEV|8|25|adipem vero et caudam omnemque pinguedinem quae operit intestina reticulumque iecoris et duos renes cum adipibus suis et armo dextro separavit
LEV|8|26|tollens autem de canistro azymorum quod erat coram Domino panem absque fermento et collyridam conspersam oleo laganumque posuit super adipes et armum dextrum
LEV|8|27|tradens simul omnia Aaron et filiis eius qui postquam levaverunt ea coram Domino
LEV|8|28|rursum suscepta de manibus eorum adolevit super altare holocausti eo quod consecrationis esset oblatio in odorem suavitatis sacrificii Domini
LEV|8|29|tulit et pectusculum elevans illud coram Domino de ariete consecrationis in partem suam sicut praeceperat ei Dominus
LEV|8|30|adsumensque unguentum et sanguinem qui erat in altari aspersit super Aaron et vestimenta eius et super filios illius ac vestes eorum
LEV|8|31|cumque sanctificasset eos in vestitu suo praecepit eis dicens coquite carnes ante fores tabernaculi et ibi comedite eas panes quoque consecrationis edite qui positi sunt in canistro sicut praecepit mihi dicens Aaron et filii eius comedent eos
LEV|8|32|quicquid autem reliquum fuerit de carne et panibus ignis absumet
LEV|8|33|de ostio quoque tabernaculi non exibitis septem diebus usque ad diem quo conplebitur tempus consecrationis vestrae septem enim diebus finitur consecratio
LEV|8|34|sicut et inpraesentiarum factum est ut ritus sacrificii conpleretur
LEV|8|35|die ac nocte manebitis in tabernaculo observantes custodias Domini ne moriamini sic enim mihi praeceptum est
LEV|8|36|feceruntque Aaron et filii eius cuncta quae locutus est Dominus per manum Mosi
LEV|9|1|facto autem octavo die vocavit Moses Aaron et filios eius ac maiores natu Israhel dixitque ad Aaron
LEV|9|2|tolle de armento vitulum pro peccato et arietem in holocaustum utrumque inmaculatos et offer illos coram Domino
LEV|9|3|et ad filios Israhel loqueris tollite hircum pro peccato et vitulum atque agnum anniculos et sine macula in holocaustum
LEV|9|4|bovem et arietem pro pacificis et immolate eos coram Domino in sacrificio singulorum similam oleo conspersam offerentes hodie enim Dominus apparebit vobis
LEV|9|5|tulerunt ergo cuncta quae iusserat Moses ad ostium tabernaculi ubi cum omnis staret multitudo
LEV|9|6|ait Moses iste est sermo quem praecepit Dominus facite et apparebit vobis gloria eius
LEV|9|7|dixit et ad Aaron accede ad altare et immola pro peccato tuo offer holocaustum et deprecare pro te et pro populo cumque mactaveris hostiam populi ora pro eo sicut praecepit Dominus
LEV|9|8|statimque Aaron accedens ad altare immolavit vitulum pro peccato suo
LEV|9|9|cuius sanguinem obtulerunt ei filii sui in quo tinguens digitum tetigit cornua altaris et fudit residuum ad basim eius
LEV|9|10|adipemque et renunculos ac reticulum iecoris quae sunt pro peccato adolevit super altare sicut praeceperat Dominus Mosi
LEV|9|11|carnes vero et pellem eius extra castra conbusit igni
LEV|9|12|immolavit et holocausti victimam obtuleruntque ei filii sui sanguinem eius quem fudit per altaris circuitum
LEV|9|13|ipsam etiam hostiam in frusta concisam cum capite et membris singulis obtulerunt quae omnia super altare cremavit igni
LEV|9|14|lotis prius aqua intestinis et pedibus
LEV|9|15|et pro peccato populi offerens mactavit hircum expiatoque altari
LEV|9|16|fecit holocaustum
LEV|9|17|addens in sacrificio libamenta quae pariter offeruntur et adolens ea super altare absque caerimoniis holocausti matutini
LEV|9|18|immolavit et bovem atque arietem hostias pacificas populi obtuleruntque ei filii sui sanguinem quem fudit super altare in circuitu
LEV|9|19|adipes autem bovis et caudam arietis renunculosque cum adipibus suis et reticulum iecoris
LEV|9|20|posuerunt super pectora cumque cremati essent adipes in altari
LEV|9|21|pectora eorum et armos dextros separavit Aaron elevans coram Domino sicut praeceperat Moses
LEV|9|22|et tendens manum contra populum benedixit eis sicque conpletis hostiis pro peccato et holocaustis et pacificis descendit
LEV|9|23|ingressi autem Moses et Aaron tabernaculum testimonii et deinceps egressi benedixerunt populo apparuitque gloria Domini omni multitudini
LEV|9|24|et ecce egressus ignis a Domino devoravit holocaustum et adipes qui erant super altare quod cum vidissent turbae laudaverunt Dominum ruentes in facies suas
LEV|10|1|arreptisque Nadab et Abiu filii Aaron turibulis posuerunt ignem et incensum desuper offerentes coram Domino ignem alienum quod eis praeceptum non erat
LEV|10|2|egressusque ignis a Domino devoravit eos et mortui sunt coram Domino
LEV|10|3|dixitque Moses ad Aaron hoc est quod locutus est Dominus sanctificabor in his qui adpropinquant mihi et in conspectu omnis populi glorificabor quod audiens tacuit Aaron
LEV|10|4|vocatis autem Moses Misahel et Elsaphan filios Ozihel patrui Aaron ait ad eos ite et colligite fratres vestros de conspectu sanctuarii et asportate extra castra
LEV|10|5|confestimque pergentes tulerunt eos sicut iacebant vestitos lineis tunicis et eiecerunt foras ut sibi fuerat imperatum
LEV|10|6|locutus est Moses ad Aaron et ad Eleazar atque Ithamar filios eius capita vestra nolite nudare et vestimenta nolite scindere ne forte moriamini et super omnem coetum oriatur indignatio fratres vestri et omnis domus Israhel plangant incendium quod Dominus suscitavit
LEV|10|7|vos autem non egredimini fores tabernaculi alioquin peribitis oleum quippe sanctae unctionis est super vos qui fecerunt omnia iuxta praeceptum Mosi
LEV|10|8|dixit quoque Dominus ad Aaron
LEV|10|9|vinum et omne quod inebriare potest non bibetis tu et filii tui quando intratis tabernaculum testimonii ne moriamini quia praeceptum est sempiternum in generationes vestras
LEV|10|10|et ut habeatis scientiam discernendi inter sanctum et profanum inter pollutum et mundum
LEV|10|11|doceatisque filios Israhel omnia legitima mea quae locutus est Dominus ad eos per manum Mosi
LEV|10|12|locutusque est Moses ad Aaron et ad Eleazar atque Ithamar filios eius qui residui erant tollite sacrificium quod remansit de oblatione Domini et comedite illud absque fermento iuxta altare quia sanctum sanctorum est
LEV|10|13|comedetis autem in loco sancto quod datum est tibi et filiis tuis de oblationibus Domini sicut praeceptum est mihi
LEV|10|14|pectusculum quoque quod oblatum est et armum qui separatus est edetis in loco mundissimo tu et filii tui ac filiae tuae tecum tibi enim ac liberis tuis reposita sunt de hostiis salutaribus filiorum Israhel
LEV|10|15|eo quod armum et pectus et adipes qui cremantur in altari elevaverint coram Domino et pertineant ad te et ad filios tuos lege perpetua sicut praecepit Dominus
LEV|10|16|inter haec hircum qui oblatus fuerat pro peccato cum quaereret Moses exustum repperit iratusque contra Eleazar et Ithamar filios Aaron qui remanserant ait
LEV|10|17|cur non comedistis hostiam pro peccato in loco sancto quae sancta sanctorum est et data vobis ut portetis iniquitatem multitudinis et rogetis pro ea in conspectu Domini
LEV|10|18|praesertim cum de sanguine illius non sit inlatum intra sancta et comedere eam debueritis in sanctuario sicut praeceptum est mihi
LEV|10|19|respondit Aaron oblata est hodie victima pro peccato et holocaustum coram Domino mihi autem accidit quod vides quomodo potui comedere eam aut placere Domino in caerimoniis mente lugubri
LEV|10|20|quod cum audisset Moses recepit satisfactionem
LEV|11|1|locutus est Dominus ad Mosen et Aaron dicens
LEV|11|2|dicite filiis Israhel haec sunt animalia quae comedere debetis de cunctis animantibus terrae
LEV|11|3|omne quod habet divisam ungulam et ruminat in pecoribus comedetis
LEV|11|4|quicquid autem ruminat quidem et habet ungulam sed non dividit eam sicut camelus et cetera non comedetis illud et inter inmunda reputabitis
LEV|11|5|chyrogryllius qui ruminat ungulamque non dividit inmundus est
LEV|11|6|lepus quoque nam et ipse ruminat sed ungulam non dividit
LEV|11|7|et sus qui cum ungulam dividat non ruminat
LEV|11|8|horum carnibus non vescemini nec cadavera contingetis quia inmunda sunt vobis
LEV|11|9|haec sunt quae gignuntur in aquis et vesci licitum est omne quod habet pinnulas et squamas tam in mari quam in fluminibus et stagnis comedetis
LEV|11|10|quicquid autem pinnulas et squamas non habet eorum quae in aquis moventur et vivunt abominabile vobis
LEV|11|11|et execrandum erit carnes eorum non comedetis et morticina vitabitis
LEV|11|12|cuncta quae non habent pinnulas et squamas in aquis polluta erunt
LEV|11|13|haec sunt quae de avibus comedere non debetis et vitanda sunt vobis aquilam et grypem et alietum
LEV|11|14|milvum ac vulturem iuxta genus suum
LEV|11|15|et omne corvini generis in similitudinem suam
LEV|11|16|strutionem et noctuam et larum et accipitrem iuxta genus suum
LEV|11|17|bubonem et mergulum et ibin
LEV|11|18|cycnum et onocrotalum et porphirionem
LEV|11|19|erodionem et charadrion iuxta genus suum opupam quoque et vespertilionem
LEV|11|20|omne de volucribus quod graditur super quattuor pedes abominabile erit vobis
LEV|11|21|quicquid autem ambulat quidem super quattuor pedes sed habet longiora retro crura per quae salit super terram
LEV|11|22|comedere debetis ut est brucus in genere suo et attacus atque ophiomachus ac lucusta singula iuxta genus suum
LEV|11|23|quicquid autem ex volucribus quattuor tantum habet pedes execrabile erit vobis
LEV|11|24|et quicumque morticina eorum tetigerit polluetur et erit inmundus usque ad vesperum
LEV|11|25|et si necesse fuerit ut portet quippiam horum mortuum lavabit vestimenta sua et inmundus erit usque ad solis occasum
LEV|11|26|omne animal quod habet quidem ungulam sed non dividit eam nec ruminat inmundum erit et quicquid tetigerit illud contaminabitur
LEV|11|27|quod ambulat super manus ex cunctis animantibus quae incedunt quadrupedia inmundum erit qui tetigerit morticina eorum polluetur usque ad vesperum
LEV|11|28|et qui portaverit huiuscemodi cadavera lavabit vestimenta sua et inmundus erit usque ad vesperum quia omnia haec inmunda sunt vobis
LEV|11|29|hoc quoque inter polluta reputabitur de his quae moventur in terra mustela et mus et corcodillus singula iuxta genus suum
LEV|11|30|migale et cameleon et stelio ac lacerta et talpa
LEV|11|31|omnia haec inmunda sunt qui tetigerit morticina eorum inmundus erit usque ad vesperum
LEV|11|32|et super quod ceciderit quicquam de morticinis eorum polluetur tam vas ligneum et vestimentum quam pelles et cilicia et in quocumque fit opus tinguentur aqua et polluta erunt usque ad vesperum et sic postea mundabuntur
LEV|11|33|vas autem fictile in quo horum quicquam intro ceciderit polluetur et idcirco frangendum est
LEV|11|34|omnis cibus quem comeditis si fusa fuerit super eum aqua inmundus erit et omne liquens quod bibitur de universo vase inmundum erit
LEV|11|35|et quicquid de morticinis istiusmodi ceciderit super illud inmundum erit sive clibani sive cytropodes destruentur et inmundi erunt
LEV|11|36|fontes vero et cisternae et omnis aquarum congregatio munda erit qui morticinum eorum tetigerit polluetur
LEV|11|37|si ceciderint super sementem non polluent eam
LEV|11|38|sin autem quispiam aqua sementem perfuderit et postea morticinis tacta fuerit ilico polluetur
LEV|11|39|si mortuum fuerit animal quod licet vobis comedere qui cadaver eius tetigerit inmundus erit usque ad vesperum
LEV|11|40|et qui comederit ex eo quippiam sive portaverit lavabit vestimenta sua et inmundus erit usque ad vesperum
LEV|11|41|omne quod reptat super terram abominabile erit nec adsumetur in cibum
LEV|11|42|quicquid super pectus quadrupes graditur et multos habet pedes sive per humum trahitur non comedetis quia abominabile est
LEV|11|43|nolite contaminare animas vestras nec tangatis quicquam eorum ne inmundi sitis
LEV|11|44|ego enim sum Dominus Deus vester sancti estote quoniam et ego sanctus sum ne polluatis animas vestras in omni reptili quod movetur super terram
LEV|11|45|ego sum Dominus qui eduxi vos de terra Aegypti ut essem vobis in Deum sancti eritis quia et ego sanctus sum
LEV|11|46|ista est lex animantium et volucrum et omnis animae viventis quae movetur in aqua et reptat in terra
LEV|11|47|ut differentias noveritis mundi et inmundi et sciatis quid comedere et quid respuere debeatis
LEV|12|1|locutus est Dominus ad Mosen dicens
LEV|12|2|loquere filiis Israhel et dices ad eos mulier si suscepto semine pepererit masculum inmunda erit septem diebus iuxta dies separationis menstruae
LEV|12|3|et die octavo circumcidetur infantulus
LEV|12|4|ipsa vero triginta tribus diebus manebit in sanguine purificationis suae omne sanctum non tanget nec ingredietur sanctuarium donec impleantur dies purificationis eius
LEV|12|5|sin autem feminam pepererit inmunda erit duabus ebdomadibus iuxta ritum fluxus menstrui et sexaginta ac sex diebus manebit in sanguine purificationis suae
LEV|12|6|cumque expleti fuerint dies purificationis eius pro filio sive pro filia deferet agnum anniculum in holocaustum et pullum columbae sive turturem pro peccato ad ostium tabernaculi testimonii et tradet sacerdoti
LEV|12|7|qui offeret illa coram Domino et rogabit pro ea et sic mundabitur a profluvio sanguinis sui ista est lex parientis masculum ac feminam
LEV|12|8|quod si non invenerit manus eius nec potuerit offerre agnum sumet duos turtures vel duos pullos columbae unum in holocaustum et alterum pro peccato orabitque pro ea sacerdos et sic mundabitur
LEV|13|1|locutus est Dominus ad Mosen et Aaron dicens
LEV|13|2|homo in cuius carne et cute ortus fuerit diversus color sive pustula aut quasi lucens quippiam id est plaga leprae adducetur ad Aaron sacerdotem vel ad unum quemlibet filiorum eius
LEV|13|3|qui cum viderit lepram in cute et pilos in album mutatos colorem ipsamque speciem leprae humiliorem cute et carne reliqua plaga leprae est et ad arbitrium eius separabitur
LEV|13|4|sin autem lucens candor fuerit in cute nec humilior carne reliqua et pili coloris pristini recludet eum sacerdos septem diebus
LEV|13|5|et considerabit die septimo et siquidem lepra ultra non creverit nec transierit in cute priores terminos rursum includet eum septem diebus aliis
LEV|13|6|et die septimo contemplabitur si obscurior fuerit lepra et non creverit in cute mundabit eum quia scabies est lavabitque homo vestimenta sua et mundus erit
LEV|13|7|quod si postquam a sacerdote visus est et redditus munditiae iterum lepra creverit adducetur ad eum
LEV|13|8|et inmunditiae condemnabitur
LEV|13|9|plaga leprae si fuerit in homine adducetur ad sacerdotem
LEV|13|10|et videbit eum cumque color albus in cute fuerit et capillorum mutarit aspectum ipsa quoque caro viva apparuerit
LEV|13|11|lepra vetustissima iudicabitur atque inolita cuti contaminabit itaque eum sacerdos et non recludet quia perspicue inmunditia est
LEV|13|12|sin autem effloruerit discurrens lepra in cute et operuerit omnem carnem a capite usque ad pedes quicquid sub aspectu oculorum cadit
LEV|13|13|considerabit eum sacerdos et teneri lepra mundissima iudicabit eo quod omnis in candorem versa sit et idcirco homo mundus erit
LEV|13|14|quando vero caro vivens in eo apparuerit
LEV|13|15|tunc sacerdotis iudicio polluetur et inter inmundos reputabitur caro enim viva si lepra aspergatur inmunda est
LEV|13|16|quod si rursum versa fuerit in alborem et totum hominem operuerit
LEV|13|17|considerabit eum sacerdos et mundum esse decernet
LEV|13|18|caro et cutis in qua ulcus natum est et sanatum
LEV|13|19|et in loco ulceris cicatrix apparuerit alba sive subrufa adducetur homo ad sacerdotem
LEV|13|20|qui cum viderit locum leprae humiliorem carne reliqua et pilos versos in candorem contaminabit eum plaga enim leprae orta est in ulcere
LEV|13|21|quod si pilus coloris est pristini et cicatrix subobscura et vicina carne non est humilior recludet eum septem diebus
LEV|13|22|et siquidem creverit adiudicabit eum leprae
LEV|13|23|sin autem steterit in loco suo ulceris est cicatrix et homo mundus erit
LEV|13|24|caro et cutis quam ignis exuserit et sanata albam sive rufam habuerit cicatricem
LEV|13|25|considerabit eam sacerdos et ecce versa est in alborem et locus eius reliqua cute humilior contaminabit eum quia plaga leprae in cicatrice orta est
LEV|13|26|quod si pilorum color non fuerit inmutatus nec humilior plaga carne reliqua et ipsa leprae species fuerit subobscura recludet eum septem diebus
LEV|13|27|et die septimo contemplabitur si creverit in cute lepra contaminabit eum
LEV|13|28|sin autem in loco suo candor steterit non satis clarus plaga conbustionis est et idcirco mundabitur quia cicatrix est conbusturae
LEV|13|29|vir sive mulier in cuius capite vel barba germinarit lepra videbit eos sacerdos
LEV|13|30|et siquidem humilior fuerit locus carne reliqua et capillus flavus solitoque subtilior contaminabit eos quia lepra capitis ac barbae est
LEV|13|31|sin autem viderit et locum maculae aequalem vicinae carni et capillum nigrum recludet eos septem diebus
LEV|13|32|et die septimo intuebitur si non creverit macula et capillus sui coloris est et locus plagae carni reliquae aequalis
LEV|13|33|radetur homo absque loco maculae et includetur septem diebus aliis
LEV|13|34|si die septimo visa fuerit stetisse plaga in loco suo nec humilior carne reliqua mundabit eum lotisque vestibus mundus erit
LEV|13|35|sin autem post emundationem rursus creverit macula in cute
LEV|13|36|non quaeret amplius utrum capillus in flavum colorem sit commutatus quia aperte inmundus est
LEV|13|37|porro si steterit macula et capilli nigri fuerint noverit hominem esse sanatum et confidenter eum pronuntiet mundum
LEV|13|38|vir et mulier in cuius cute candor apparuerit
LEV|13|39|intuebitur eos sacerdos si deprehenderit subobscurum alborem lucere in cute sciat non esse lepram sed maculam coloris candidi et hominem mundum
LEV|13|40|vir de cuius capite capilli fluunt calvus ac mundus est
LEV|13|41|et si a fronte ceciderint pili recalvaster et mundus est
LEV|13|42|sin autem in calvitio sive in recalvatione albus vel rufus color fuerit exortus
LEV|13|43|et hoc sacerdos viderit condemnabit eum haut dubiae leprae quae orta est in calvitio
LEV|13|44|quicumque ergo maculatus fuerit lepra et separatus ad arbitrium sacerdotis
LEV|13|45|habebit vestimenta dissuta caput nudum os veste contectum contaminatum ac sordidum se clamabit
LEV|13|46|omni tempore quo leprosus est et inmundus solus habitabit extra castra
LEV|13|47|vestis lanea sive linea quae lepram habuerit
LEV|13|48|in stamine atque subtemine aut certe pellis vel quicquid ex pelle confectum est
LEV|13|49|si alba aut rufa macula fuerit infecta lepra reputabitur ostendeturque sacerdoti
LEV|13|50|qui consideratam recludet septem diebus
LEV|13|51|et die septimo rursus aspiciens si crevisse deprehenderit lepra perseverans est pollutum iudicabit vestimentum et omne in quo fuerit inventa
LEV|13|52|et idcirco conburetur flammis
LEV|13|53|quod si eam viderit non crevisse
LEV|13|54|praecipiet et lavabunt id in quo lepra est recludetque illud septem diebus aliis
LEV|13|55|et cum viderit faciem quidem pristinam non reversam nec tamen crevisse lepram inmundum iudicabit et igne conburet eo quod infusa sit in superficie vestimenti vel per totum lepra
LEV|13|56|sin autem obscurior fuerit locus leprae postquam vestis est lota abrumpet eum et a solido dividet
LEV|13|57|quod si ultra apparuerit in his locis quae prius inmaculata erant lepra volatilis et vaga debet igne conburi
LEV|13|58|si cessaverit lavabit ea quae pura sunt secundo et munda erunt
LEV|13|59|ista est lex leprae vestimenti lanei et linei staminis atque subteminis omnisque supellectilis pelliciae quomodo mundari debeat vel contaminari
LEV|14|1|locutusque est Dominus ad Mosen dicens
LEV|14|2|hic est ritus leprosi quando mundandus est adducetur ad sacerdotem
LEV|14|3|qui egressus e castris cum invenerit lepram esse mundatam
LEV|14|4|praecipiet ei qui purificatur ut offerat pro se duos passeres vivos quos vesci licitum est et lignum cedrinum vermiculumque et hysopum
LEV|14|5|et unum e passeribus immolari iubebit in vase fictili super aquas viventes
LEV|14|6|alium autem vivum cum ligno cedrino et cocco et hysopo tinguet in sanguine passeris immolati
LEV|14|7|quo asperget illum qui mundandus est septies ut iure purgetur et dimittet passerem vivum ut in agrum avolet
LEV|14|8|cumque laverit homo vestimenta sua radet omnes pilos corporis et lavabitur aqua purificatusque ingredietur castra ita dumtaxat ut maneat extra tabernaculum suum septem diebus
LEV|14|9|et die septimo radat capillos capitis barbamque et supercilia ac totius corporis pilos et lotis rursum vestibus et corpore
LEV|14|10|die octavo adsumet duos agnos inmaculatos et ovem anniculam absque macula et tres decimas similae in sacrificium quae conspersa sit oleo et seorsum olei sextarium
LEV|14|11|cumque sacerdos purificans hominem statuerit eum et haec omnia coram Domino in ostio tabernaculi testimonii
LEV|14|12|tollet agnum et offeret eum pro delicto oleique sextarium et oblatis ante Dominum omnibus
LEV|14|13|immolabit agnum ubi immolari solet hostia pro peccato et holocaustum id est in loco sancto sicut enim pro peccato ita et pro delicto ad sacerdotem pertinet hostia sancta sanctorum est
LEV|14|14|adsumensque sacerdos de sanguine hostiae quae immolata est pro delicto ponet super extremum auriculae dextrae eius qui mundatur et super pollices manus dextrae et pedis
LEV|14|15|et de olei sextario mittet in manum suam sinistram
LEV|14|16|tinguetque digitum dextrum in eo et asperget septies contra Dominum
LEV|14|17|quod autem reliquum est olei in leva manu fundet super extremum auriculae dextrae eius qui mundatur et super pollices manus ac pedis dextri et super sanguinem qui fusus est pro delicto
LEV|14|18|et super caput eius
LEV|14|19|rogabitque pro eo coram Domino et faciet sacrificium pro peccato tunc immolabit holocaustum
LEV|14|20|et ponet illud in altari cum libamentis suis et homo rite mundabitur
LEV|14|21|quod si pauper est et non potest manus eius invenire quae dicta sunt adsumet agnum pro delicto ad oblationem ut roget pro eo sacerdos decimamque partem similae conspersae oleo in sacrificium et olei sextarium
LEV|14|22|duosque turtures sive duos pullos columbae quorum sit unus pro peccato et alter in holocaustum
LEV|14|23|offeretque ea die octavo purificationis suae sacerdoti ad ostium tabernaculi testimonii coram Domino
LEV|14|24|qui suscipiens agnum pro delicto et sextarium olei levabit simul
LEV|14|25|immolatoque agno de sanguine eius ponet super extremum auriculae dextrae illius qui mundatur et super pollices manus eius ac pedis dextri
LEV|14|26|olei vero partem mittet in manum suam sinistram
LEV|14|27|in quo tinguens digitum dextrae manus asperget septies contra Dominum
LEV|14|28|tangetque extremum dextrae auriculae illius qui mundatur et pollices manus ac pedis dextri in loco sanguinis qui effusus est pro delicto
LEV|14|29|reliquam autem partem olei quae est in sinistra manu mittet super caput purificati ut placet pro eo Dominum
LEV|14|30|et turturem sive pullum columbae offeret
LEV|14|31|unum pro delicto et alterum in holocaustum cum libamentis suis
LEV|14|32|hoc est sacrificium leprosi qui habere non potest omnia in emundationem sui
LEV|14|33|locutus est Dominus ad Mosen et Aaron dicens
LEV|14|34|cum ingressi fueritis terram Chanaan quam ego dabo vobis in possessionem si fuerit plaga leprae in aedibus
LEV|14|35|ibit cuius est domus nuntians sacerdoti et dicet quasi plaga leprae videtur mihi esse in domo mea
LEV|14|36|at ille praecipiet ut efferant universa de domo priusquam ingrediatur eam et videat utrum lepra sit ne inmunda fiant omnia quae in domo sunt intrabitque postea ut consideret domus lepram
LEV|14|37|et cum viderit in parietibus illius quasi valliculas pallore sive rubore deformes et humiliores superficie reliqua
LEV|14|38|egredietur ostium domus et statim claudet eam septem diebus
LEV|14|39|reversusque die septimo considerabit eam si invenerit crevisse lepram
LEV|14|40|iubebit erui lapides in quibus lepra est et proici eos extra civitatem in loco inmundo
LEV|14|41|domum autem ipsam radi intrinsecus per circuitum et spargi pulverem rasurae extra urbem in loco inmundo
LEV|14|42|lapidesque alios reponi pro his qui ablati fuerint et luto alio liniri domum
LEV|14|43|sin autem postquam eruti sunt lapides et pulvis elatus et alia terra lita
LEV|14|44|ingressus sacerdos viderit reversam lepram et parietes aspersos maculis lepra est perseverans et inmunda domus
LEV|14|45|quam statim destruent et lapides eius ac ligna atque universum pulverem proicient extra oppidum in loco inmundo
LEV|14|46|qui intraverit domum quando clausa est inmundus erit usque ad vesperum
LEV|14|47|et qui dormierit in ea et comederit quippiam lavabit vestimenta sua
LEV|14|48|quod si introiens sacerdos viderit lepram non crevisse in domo postquam denuo lita est purificabit eam reddita sanitate
LEV|14|49|et in purificationem eius sumet duos passeres lignumque cedrinum et vermiculum atque hysopum
LEV|14|50|et immolato uno passere in vase fictili super aquas vivas
LEV|14|51|tollet lignum cedrinum et hysopum et coccum et passerem vivum et intinguet omnia in sanguine passeris immolati atque in aquis viventibus et asperget domum septies
LEV|14|52|purificabitque eam tam in sanguine passeris quam in aquis viventibus et in passere vivo lignoque cedrino et hysopo atque vermiculo
LEV|14|53|cumque dimiserit passerem avolare in agrum libere orabit pro domo et iure mundabitur
LEV|14|54|ista est lex omnis leprae et percussurae
LEV|14|55|leprae vestium et domorum
LEV|14|56|cicatricis et erumpentium papularum lucentis maculae et in varias species coloribus inmutatis
LEV|14|57|ut possit sciri quo tempore mundum quid vel inmundum sit
LEV|15|1|locutusque est Dominus ad Mosen et Aaron dicens
LEV|15|2|loquimini filiis Israhel et dicite eis vir qui patitur fluxum seminis inmundus erit
LEV|15|3|et tunc iudicabitur huic vitio subiacere cum per momenta singula adheserit carni illius atque concreverit foedus humor
LEV|15|4|omne stratum in quo dormierit inmundum erit et ubicumque sederit
LEV|15|5|si quis hominum tetigerit lectum eius lavabit vestimenta sua et ipse lotus aqua inmundus erit usque ad vesperum
LEV|15|6|si sederit ubi ille sederat et ipse lavabit vestimenta sua et lotus aqua inmundus erit usque ad vesperum
LEV|15|7|qui tetigerit carnem eius lavabit vestimenta sua et ipse lotus aqua inmundus erit usque ad vesperum
LEV|15|8|si salivam huiuscemodi homo iecerit super eum qui mundus est lavabit vestem suam et lotus aqua inmundus erit usque ad vesperum
LEV|15|9|sagma super quo sederit inmundum erit
LEV|15|10|et quicquid sub eo fuerit qui fluxum seminis patitur pollutum erit usque ad vesperum qui portaverit horum aliquid lavabit vestem suam et ipse lotus aqua inmundus erit usque ad vesperum
LEV|15|11|omnis quem tetigerit qui talis est non lotis ante manibus lavabit vestimenta sua et lotus aqua inmundus erit usque ad vesperum
LEV|15|12|vas fictile quod tetigerit confringetur vas autem ligneum lavabitur aqua
LEV|15|13|si sanatus fuerit qui huiuscemodi sustinet passionem numerabit septem dies post emundationem sui et lotis vestibus ac toto corpore in aquis viventibus erit mundus
LEV|15|14|die autem octavo sumet duos turtures aut duos pullos columbae et veniet in conspectu Domini ad ostium tabernaculi testimonii dabitque eos sacerdoti
LEV|15|15|qui faciet unum pro peccato et alterum in holocaustum rogabitque pro eo coram Domino ut emundetur a fluxu seminis sui
LEV|15|16|vir de quo egreditur semen coitus lavabit aqua omne corpus suum et inmundus erit usque ad vesperum
LEV|15|17|vestem et pellem quam habuerit lavabit aqua et inmunda erit usque ad vesperum
LEV|15|18|mulier cum qua coierit lavabitur aqua et inmunda erit usque ad vesperum
LEV|15|19|mulier quae redeunte mense patitur fluxum sanguinis septem diebus separabitur
LEV|15|20|omnis qui tetigerit eam inmundus erit usque ad vesperum
LEV|15|21|et in quo dormierit vel sederit diebus separationis suae polluetur
LEV|15|22|qui tetigerit lectum eius lavabit vestimenta sua et ipse lotus aqua inmundus erit usque ad vesperum
LEV|15|23|omne vas super quo illa sederit quisquis adtigerit lavabit vestimenta sua et lotus aqua pollutus erit usque ad vesperum
LEV|15|24|si coierit cum ea vir tempore sanguinis menstrualis inmundus erit septem diebus et omne stratum in quo dormierit polluetur
LEV|15|25|mulier quae patitur multis diebus fluxum sanguinis non in tempore menstruali vel quae post menstruum sanguinem fluere non cessat quamdiu huic subiacet passioni inmunda erit quasi sit in tempore menstruo
LEV|15|26|omne stratum in quo dormierit et vas in quo sederit pollutum erit
LEV|15|27|quicumque tetigerit eam lavabit vestimenta sua et ipse lotus aqua inmundus erit usque ad vesperum
LEV|15|28|si steterit sanguis et fluere cessarit numerabit septem dies purificationis suae
LEV|15|29|et octavo die offeret pro se sacerdoti duos turtures vel duos pullos columbae ad ostium tabernaculi testimonii
LEV|15|30|qui unum faciet pro peccato et alterum in holocaustum rogabitque pro ea coram Domino et pro fluxu inmunditiae eius
LEV|15|31|docebitis ergo filios Israhel ut caveant inmunditiam et non moriantur in sordibus suis cum polluerint tabernaculum meum quod est inter eos
LEV|15|32|ista est lex eius qui patitur fluxum seminis et qui polluitur coitu
LEV|15|33|et quae menstruis temporibus separatur vel quae iugi fluit sanguine et hominis qui dormierit cum ea
LEV|16|1|locutusque est Dominus ad Mosen post mortem duum filiorum Aaron quando offerentes ignem alienum interfecti sunt
LEV|16|2|et praecepit ei dicens loquere ad Aaron fratrem tuum ne omni tempore ingrediatur sanctuarium quod est intra velum coram propitiatorio quo tegitur arca ut non moriatur quia in nube apparebo super oraculum
LEV|16|3|nisi haec ante fecerit vitulum offeret pro peccato et arietem in holocaustum
LEV|16|4|tunica linea vestietur feminalibus lineis verecunda celabit accingetur zona linea cidarim lineam inponet capiti haec enim vestimenta sunt sancta quibus cunctis cum lotus fuerit induetur
LEV|16|5|suscipietque ab universa multitudine filiorum Israhel duos hircos pro peccato et unum arietem in holocaustum
LEV|16|6|cumque obtulerit vitulum et oraverit pro se et pro domo sua
LEV|16|7|duos hircos stare faciet coram Domino in ostio tabernaculi testimonii
LEV|16|8|mittens super utrumque sortem unam Domino et alteram capro emissario
LEV|16|9|cuius sors exierit Domino offeret illum pro peccato
LEV|16|10|cuius autem in caprum emissarium statuet eum vivum coram Domino ut fundat preces super eo et emittat illum in solitudinem
LEV|16|11|his rite celebratis offeret vitulum et rogans pro se et pro domo sua immolabit eum
LEV|16|12|adsumptoque turibulo quod de prunis altaris impleverit et hauriens manu conpositum thymiama in incensum ultra velum intrabit in sancta
LEV|16|13|ut positis super ignem aromatibus nebula eorum et vapor operiat oraculum quod est super testimonium et non moriatur
LEV|16|14|tollet quoque de sanguine vituli et asperget digito septies contra propitiatorium ad orientem
LEV|16|15|cumque mactaverit hircum pro peccato populi inferet sanguinem eius intra velum sicut praeceptum est de sanguine vituli ut aspergat e regione oraculi
LEV|16|16|et expiet sanctuarium ab inmunditiis filiorum Israhel et a praevaricationibus eorum cunctisque peccatis iuxta hunc ritum faciet tabernaculo testimonii quod fixum est inter eos in medio sordium habitationis eorum
LEV|16|17|nullus hominum sit in tabernaculo quando pontifex ingreditur sanctuarium ut roget pro se et pro domo sua et pro universo coetu Israhel donec egrediatur
LEV|16|18|cum autem exierit ad altare quod coram Domino est oret pro se et sumptum sanguinem vituli atque hirci fundat super cornua eius per gyrum
LEV|16|19|aspergensque digito septies expiet et sanctificet illud ab inmunditiis filiorum Israhel
LEV|16|20|postquam emundarit sanctuarium et tabernaculum et altare tunc offerat hircum viventem
LEV|16|21|et posita utraque manu super caput eius confiteatur omnes iniquitates filiorum Israhel et universa delicta atque peccata eorum quae inprecans capiti eius emittet illum per hominem paratum in desertum
LEV|16|22|cumque portaverit hircus omnes iniquitates eorum in terram solitariam et dimissus fuerit in deserto
LEV|16|23|revertetur Aaron in tabernaculum testimonii et depositis vestibus quibus prius indutus erat cum intraret sanctuarium relictisque ibi
LEV|16|24|lavabit carnem suam in loco sancto indueturque vestimentis suis et postquam egressus obtulerit holocaustum suum ac plebis rogabit tam pro se quam pro populo
LEV|16|25|et adipem qui oblatus est pro peccatis adolebit super altare
LEV|16|26|ille vero qui dimiserit caprum emissarium lavabit vestimenta sua et corpus aqua et sic ingredietur in castra
LEV|16|27|vitulum autem et hircum qui pro peccato fuerant immolati et quorum sanguis inlatus est ut in sanctuario expiatio conpleretur asportabunt foras castra et conburent igni tam pelles quam carnes eorum et fimum
LEV|16|28|et quicumque conbuserit ea lavabit vestimenta sua et carnem aqua et sic ingredietur in castra
LEV|16|29|eritque hoc vobis legitimum sempiternum mense septimo decima die mensis adfligetis animas vestras nullumque facietis opus sive indigena sive advena qui peregrinatur inter vos
LEV|16|30|in hac die expiatio erit vestri atque mundatio ab omnibus peccatis vestris coram Domino mundabimini
LEV|16|31|sabbatum enim requietionis est et adfligetis animas vestras religione perpetua
LEV|16|32|expiabit autem sacerdos qui unctus fuerit et cuius initiatae manus ut sacerdotio fungatur pro patre suo indueturque stola linea et vestibus sanctis
LEV|16|33|et expiabit sanctuarium et tabernaculum testimonii atque altare sacerdotes quoque et universum populum
LEV|16|34|eritque hoc vobis legitimum sempiternum ut oretis pro filiis Israhel et pro cunctis peccatis eorum semel in anno fecit igitur sicut praeceperat Dominus Mosi
LEV|17|1|et locutus est Dominus ad Mosen dicens
LEV|17|2|loquere Aaron et filiis eius et cunctis filiis Israhel et dices ad eos iste est sermo quem mandavit Dominus dicens
LEV|17|3|homo quilibet de domo Israhel si occiderit bovem aut ovem sive capram in castris vel extra castra
LEV|17|4|et non obtulerit ad ostium tabernaculi oblationem Domino sanguinis reus erit quasi sanguinem fuderit sic peribit de medio populi sui
LEV|17|5|ideo offerre debent sacerdoti filii Israhel hostias suas quas occidunt in agro ut sanctificentur Domino ante ostium tabernaculi testimonii et immolent eas hostias pacificas Domino
LEV|17|6|fundetque sacerdos sanguinem super altare Domini ad ostium tabernaculi testimonii et adolebit adipem in odorem suavitatis Domino
LEV|17|7|et nequaquam ultra immolabunt hostias suas daemonibus cum quibus fornicati sunt legitimum sempiternum erit illis et posteris eorum
LEV|17|8|et ad ipsos dices homo de domo Israhel et de advenis qui peregrinantur apud vos qui obtulerit holocaustum sive victimam
LEV|17|9|et ad ostium tabernaculi testimonii non adduxerit eam ut offeratur Domino interibit de populo suo
LEV|17|10|homo quilibet de domo Israhel et de advenis qui peregrinantur inter eos si comederit sanguinem obfirmabo faciem meam contra animam illius et disperdam eam de populo suo
LEV|17|11|quia anima carnis in sanguine est et ego dedi illum vobis ut super altare in eo expietis pro animabus vestris et sanguis pro animae piaculo sit
LEV|17|12|idcirco dixi filiis Israhel omnis anima ex vobis non comedet sanguinem nec ex advenis qui peregrinantur inter vos
LEV|17|13|homo quicumque de filiis Israhel et de advenis qui peregrinantur apud vos si venatione atque aucupio ceperit feram vel avem quibus vesci licitum est fundat sanguinem eius et operiat illum terra
LEV|17|14|anima enim omnis carnis in sanguine est unde dixi filiis Israhel sanguinem universae carnis non comedetis quia anima carnis in sanguine est et quicumque comederit illum interibit
LEV|17|15|anima quae comederit morticinum vel captum a bestia tam de indigenis quam de advenis lavabit vestes suas et semet ipsum aqua et contaminatus erit usque ad vesperum et hoc ordine mundus fiet
LEV|17|16|quod si non laverit vestimenta sua nec corpus portabit iniquitatem suam
LEV|18|1|locutusque est Dominus ad Mosen dicens
LEV|18|2|loquere filiis Israhel et dices ad eos ego Dominus Deus vester
LEV|18|3|iuxta consuetudinem terrae Aegypti in qua habitastis non facietis et iuxta morem regionis Chanaan ad quam ego introducturus sum vos non agetis nec in legitimis eorum ambulabitis
LEV|18|4|facietis iudicia mea et praecepta servabitis et ambulabitis in eis ego Dominus Deus vester
LEV|18|5|custodite leges meas atque iudicia quae faciens homo vivet in eis ego Dominus
LEV|18|6|omnis homo ad proximam sanguinis sui non accedet ut revelet turpitudinem eius ego Dominus
LEV|18|7|turpitudinem patris et turpitudinem matris tuae non discoperies mater tua est non revelabis turpitudinem eius
LEV|18|8|turpitudinem uxoris patris tui non discoperies turpitudo enim patris tui est
LEV|18|9|turpitudinem sororis tuae ex patre sive ex matre quae domi vel foris genita est non revelabis
LEV|18|10|turpitudinem filiae filii tui vel neptis ex filia non revelabis quia turpitudo tua est
LEV|18|11|turpitudinem filiae uxoris patris tui quam peperit patri tuo et est soror tua non revelabis
LEV|18|12|turpitudinem sororis patris tui non discoperies quia caro est patris tui
LEV|18|13|turpitudinem sororis matris tuae non revelabis eo quod caro sit matris tuae
LEV|18|14|turpitudinem patrui tui non revelabis nec accedes ad uxorem eius quae tibi adfinitate coniungitur
LEV|18|15|turpitudinem nurus tuae non revelabis quia uxor filii tui est nec discoperies ignominiam eius
LEV|18|16|turpitudinem uxoris fratris tui non revelabis quia turpitudo fratris tui est
LEV|18|17|turpitudinem uxoris tuae et filiae eius non revelabis filiam filii eius et filiam filiae illius non sumes ut reveles ignominiam eius quia caro illius sunt et talis coitus incestus est
LEV|18|18|sororem uxoris tuae in pelicatum illius non accipies nec revelabis turpitudinem eius adhuc illa vivente
LEV|18|19|ad mulierem quae patitur menstrua non accedes nec revelabis foeditatem eius
LEV|18|20|cum uxore proximi tui non coibis nec seminis commixtione maculaberis
LEV|18|21|de semine tuo non dabis ut consecretur idolo Moloch nec pollues nomen Dei tui ego Dominus
LEV|18|22|cum masculo non commisceberis coitu femineo quia abominatio est
LEV|18|23|cum omni pecore non coibis nec maculaberis cum eo mulier non subcumbet iumento nec miscebitur ei quia scelus est
LEV|18|24|ne polluamini in omnibus his quibus contaminatae sunt universae gentes quas ego eiciam ante conspectum vestrum
LEV|18|25|et quibus polluta est terra cuius ego scelera visitabo ut evomat habitatores suos
LEV|18|26|custodite legitima mea atque iudicia et non faciat ex omnibus abominationibus istis tam indigena quam colonus qui peregrinatur apud vos
LEV|18|27|omnes enim execrationes istas fecerunt accolae terrae qui fuerunt ante vos et polluerunt eam
LEV|18|28|cavete ergo ne et vos similiter evomat cum paria feceritis sicut evomuit gentem quae fuit ante vos
LEV|18|29|omnis anima quae fecerit de abominationibus his quippiam peribit de medio populi sui
LEV|18|30|custodite mandata mea nolite facere quae fecerunt hii qui fuerunt ante vos et ne polluamini in eis ego Dominus Deus vester
LEV|19|1|locutus est Dominus ad Mosen dicens
LEV|19|2|loquere ad omnem coetum filiorum Israhel et dices ad eos sancti estote quia ego sanctus sum Dominus Deus vester
LEV|19|3|unusquisque matrem et patrem suum timeat sabbata mea custodite ego Dominus Deus vester
LEV|19|4|nolite converti ad idola nec deos conflatiles faciatis vobis ego Dominus Deus vester
LEV|19|5|si immolaveritis hostiam pacificorum Domino ut sit placabilis
LEV|19|6|eo die quo fuerit immolata comedetis eam et die altero quicquid autem residuum fuerit in diem tertium igne conburetis
LEV|19|7|si quis post biduum comederit ex ea profanus erit et impietatis reus
LEV|19|8|portabit iniquitatem suam quia sanctum Domini polluit et peribit anima illa de populo suo
LEV|19|9|cum messueris segetes terrae tuae non tondebis usque ad solum superficiem terrae nec remanentes spicas colliges
LEV|19|10|neque in vinea tua racemos et grana decidentia congregabis sed pauperibus et peregrinis carpenda dimittes ego Dominus Deus vester
LEV|19|11|non facietis furtum non mentiemini nec decipiet unusquisque proximum suum
LEV|19|12|non peierabis in nomine meo nec pollues nomen Dei tui ego Dominus
LEV|19|13|non facies calumniam proximo tuo nec vi opprimes eum non morabitur opus mercennarii apud te usque mane
LEV|19|14|non maledices surdo nec coram caeco pones offendiculum sed timebis Deum tuum quia ego sum Dominus
LEV|19|15|non facies quod iniquum est nec iniuste iudicabis nec consideres personam pauperis nec honores vultum potentis iuste iudica proximo tuo
LEV|19|16|non eris criminator et susurro in populis non stabis contra sanguinem proximi tui ego Dominus
LEV|19|17|ne oderis fratrem tuum in corde tuo sed publice argue eum ne habeas super illo peccatum
LEV|19|18|non quaeres ultionem nec memor eris iniuriae civium tuorum diliges amicum tuum sicut temet ipsum ego Dominus
LEV|19|19|leges meas custodite iumenta tua non facies coire cum alterius generis animantibus agrum non seres diverso semine veste quae ex duobus texta est non indueris
LEV|19|20|homo si dormierit cum muliere coitu seminis quae sit ancilla etiam nubilis et tamen pretio non redempta nec libertate donata vapulabunt ambo et non morientur quia non fuit libera
LEV|19|21|pro delicto autem suo offeret Domino ad ostium tabernaculi testimonii arietem
LEV|19|22|orabitque pro eo sacerdos et pro delicto eius coram Domino et repropitiabitur ei dimitteturque peccatum
LEV|19|23|quando ingressi fueritis terram et plantaveritis in ea ligna pomifera auferetis praeputia eorum poma quae germinant inmunda erunt vobis nec edetis ex eis
LEV|19|24|quarto anno omnis fructus eorum sanctificabitur laudabilis Domino
LEV|19|25|quinto autem anno comedetis fructus congregantes poma quae proferunt ego Dominus Deus vester
LEV|19|26|non comedetis cum sanguine non augurabimini nec observabitis somnia
LEV|19|27|neque in rotundum adtondebitis comam nec radatis barbam
LEV|19|28|et super mortuo non incidetis carnem vestram neque figuras aliquas et stigmata facietis vobis ego Dominus
LEV|19|29|ne prostituas filiam tuam et contaminetur terra et impleatur piaculo
LEV|19|30|sabbata mea custodite et sanctuarium meum metuite ego Dominus
LEV|19|31|ne declinetis ad magos nec ab ariolis aliquid sciscitemini ut polluamini per eos ego Dominus Deus vester
LEV|19|32|coram cano capite consurge et honora personam senis et time Deum tuum ego sum Dominus
LEV|19|33|si habitaverit advena in terra vestra et moratus fuerit inter vos ne exprobretis ei
LEV|19|34|sed sit inter vos quasi indigena et diligetis eum quasi vosmet ipsos fuistis enim et vos advenae in terra Aegypti ego Dominus Deus vester
LEV|19|35|nolite facere iniquum aliquid in iudicio in regula in pondere in mensura
LEV|19|36|statera iusta et aequa sint pondera iustus modius aequusque sextarius ego Dominus Deus vester qui eduxi vos de terra Aegypti
LEV|19|37|custodite omnia praecepta mea et universa iudicia et facite ea ego Dominus
LEV|20|1|locutusque est Dominus ad Mosen dicens
LEV|20|2|haec loqueris filiis Israhel homo de filiis Israhel et de advenis qui habitant in Israhel si quis dederit de semine suo idolo Moloch morte moriatur populus terrae lapidabit eum
LEV|20|3|et ego ponam faciem meam contra illum succidamque eum de medio populi sui eo quod dederit de semine suo Moloch et contaminaverit sanctuarium meum ac polluerit nomen sanctum meum
LEV|20|4|quod si neglegens populus terrae et quasi parvipendens imperium meum dimiserit hominem qui dederit de semine suo Moloch nec voluerit eum occidere
LEV|20|5|ponam faciem meam super hominem illum et cognationem eius succidamque et ipsum et omnes qui consenserunt ei ut fornicarentur cum Moloch de medio populi sui
LEV|20|6|anima quae declinaverit ad magos et ariolos et fornicata fuerit cum eis ponam faciem meam contra eam et interficiam illam de medio populi sui
LEV|20|7|sanctificamini et estote sancti quia ego Dominus Deus vester
LEV|20|8|custodite praecepta mea et facite ea ego Dominus qui sanctifico vos
LEV|20|9|qui maledixerit patri suo et matri morte moriatur patri matrique maledixit sanguis eius sit super eum
LEV|20|10|si moechatus quis fuerit cum uxore alterius et adulterium perpetrarit cum coniuge proximi sui morte moriantur et moechus et adultera
LEV|20|11|qui dormierit cum noverca sua et revelaverit ignominiam patris sui morte moriantur ambo sanguis eorum sit super eos
LEV|20|12|si quis dormierit cum nuru sua uterque moriantur quia scelus operati sunt sanguis eorum sit super eos
LEV|20|13|qui dormierit cum masculo coitu femineo uterque operati sunt nefas morte moriantur sit sanguis eorum super eos
LEV|20|14|qui supra uxorem filiam duxerit matrem eius scelus operatus est vivus ardebit cum eis nec permanebit tantum nefas in medio vestri
LEV|20|15|qui cum iumento et pecore coierit morte moriatur pecus quoque occidite
LEV|20|16|mulier quae subcubuerit cuilibet iumento simul interficietur cum eo sanguis eorum sit super eos
LEV|20|17|qui acceperit sororem suam filiam patris sui vel filiam matris suae et viderit turpitudinem eius illaque conspexerit fratris ignominiam nefariam rem operati sunt occidentur in conspectu populi sui eo quod turpitudinem suam mutuo revelarint et portabunt iniquitatem suam
LEV|20|18|qui coierit cum muliere in fluxu menstruo et revelaverit turpitudinem eius ipsaque aperuerit fontem sanguinis sui interficientur ambo de medio populi sui
LEV|20|19|turpitudinem materterae tuae et amitae tuae non discoperies qui hoc fecerit ignominiam carnis suae nudavit portabunt ambo iniquitatem suam
LEV|20|20|qui coierit cum uxore patrui vel avunculi sui et revelaverit ignominiam cognationis suae portabunt ambo peccatum suum absque liberis morientur
LEV|20|21|qui duxerit uxorem fratris sui rem facit inlicitam turpitudinem fratris sui revelavit absque filiis erunt
LEV|20|22|custodite leges meas atque iudicia et facite ea ne et vos evomat terra quam intraturi estis et habitaturi
LEV|20|23|nolite ambulare in legitimis nationum quas ego expulsurus sum ante vos omnia enim haec fecerunt et abominatus sum eos
LEV|20|24|vobis autem loquor possidete terram eorum quam dabo vobis in hereditatem terram fluentem lacte et melle ego Dominus Deus vester qui separavi vos a ceteris populis
LEV|20|25|separate ergo et vos iumentum mundum ab inmundo et avem mundam ab inmunda ne polluatis animas vestras in pecore et in avibus et cunctis quae moventur in terra et quae vobis ostendi esse polluta
LEV|20|26|eritis sancti mihi quia sanctus ego sum Dominus et separavi vos a ceteris populis ut essetis mei
LEV|20|27|vir sive mulier in quibus pythonicus vel divinationis fuerit spiritus morte moriantur lapidibus obruent eos sanguis eorum sit super illos
LEV|21|1|dixit quoque Dominus ad Mosen loquere ad sacerdotes filios Aaron et dices eis ne contaminetur sacerdos in mortibus civium suorum
LEV|21|2|nisi tantum in consanguineis ac propinquis id est super matre et patre et filio ac filia fratre quoque
LEV|21|3|et sorore virgine quae non est nupta viro
LEV|21|4|sed nec in principe populi sui contaminabitur
LEV|21|5|non radent caput nec barbam neque in carnibus suis facient incisuras
LEV|21|6|sancti erunt Deo suo et non polluent nomen eius incensum enim Domini et panes Dei sui offerunt et ideo sancti erunt
LEV|21|7|scortum et vile prostibulum non ducet uxorem nec eam quae repudiata est a marito quia consecratus est Deo suo
LEV|21|8|et panes propositionis offert sit ergo sanctus quia et ego sanctus sum Dominus qui sanctifico vos
LEV|21|9|sacerdotis filia si deprehensa fuerit in stupro et violaverit nomen patris sui flammis exuretur
LEV|21|10|pontifex id est sacerdos maximus inter fratres suos super cuius caput fusum est unctionis oleum et cuius manus in sacerdotio consecratae sunt vestitusque est sanctis vestibus caput suum non discoperiet vestimenta non scindet
LEV|21|11|et ad omnem mortuum non ingredietur omnino super patre quoque suo et matre non contaminabitur
LEV|21|12|nec egredietur de sanctis ne polluat sanctuarium Domini quia oleum sanctae unctionis Dei sui super eum est ego Dominus
LEV|21|13|virginem ducet uxorem
LEV|21|14|viduam et repudiatam et sordidam atque meretricem non accipiet sed puellam de populo suo
LEV|21|15|ne commisceat stirpem generis sui vulgo gentis suae quia ego Dominus qui sanctifico eum
LEV|21|16|locutusque est Dominus ad Mosen dicens
LEV|21|17|loquere ad Aaron homo de semine tuo per familias qui habuerit maculam non offeret panes Deo suo
LEV|21|18|nec accedet ad ministerium eius si caecus fuerit si claudus si vel parvo vel grandi et torto naso
LEV|21|19|si fracto pede si manu
LEV|21|20|si gibbus si lippus si albuginem habens in oculo si iugem scabiem si inpetiginem in corpore vel hirniosus
LEV|21|21|omnis qui habuerit maculam de semine Aaron sacerdotis non accedet offerre hostias Domino nec panes Deo suo
LEV|21|22|vescetur tamen panibus qui offeruntur in sanctuario
LEV|21|23|ita dumtaxat ut intra velum non ingrediatur nec accedat ad altare quia maculam habet et contaminare non debet sanctuarium meum ego Dominus qui sanctifico eos
LEV|21|24|locutus est ergo Moses ad Aaron et filios eius et ad omnem Israhel cuncta quae sibi fuerant imperata
LEV|22|1|locutus quoque est Dominus ad Mosen dicens
LEV|22|2|loquere ad Aaron et ad filios eius ut caveant ab his quae consecrata sunt filiorum Israhel et non contaminent nomen sanctificatorum mihi quae ipsi offerunt ego Dominus
LEV|22|3|dic ad eos et ad posteros eorum omnis homo qui accesserit de stirpe vestra ad ea quae consecrata sunt et quae obtulerunt filii Israhel Domino in quo est inmunditia peribit coram Domino ego sum Dominus
LEV|22|4|homo de semine Aaron qui fuerit leprosus aut patiens fluxum seminis non vescetur de his quae sanctificata sunt mihi donec sanetur qui tetigerit inmundum super mortuo et ex quo egreditur semen quasi coitus
LEV|22|5|et qui tangit reptile et quodlibet inmundum cuius tactus est sordidus
LEV|22|6|inmundus erit usque ad vesperum et non vescetur his quae sanctificata sunt sed cum laverit carnem suam aqua
LEV|22|7|et occubuerit sol tunc mundatus vescetur de sanctificatis quia cibus illius est
LEV|22|8|morticinum et captum a bestia non comedent nec polluentur in eis ego sum Dominus
LEV|22|9|custodient praecepta mea ut non subiaceant peccato et moriantur in sanctuario cum polluerint illud ego Dominus qui sanctifico eos
LEV|22|10|omnis alienigena non comedet de sanctificatis inquilinus sacerdotis et mercennarius non vescentur ex eis
LEV|22|11|quem autem sacerdos emerit et qui vernaculus domus eius fuerit hii comedent ex eis
LEV|22|12|si filia sacerdotis cuilibet ex populo nupta fuerit de his quae sanctificata sunt et de primitiis non vescetur
LEV|22|13|sin autem vidua vel repudiata et absque liberis reversa fuerit ad domum patris sui sicut puella consuerat aletur cibis patris sui omnis alienigena comedendi ex eis non habet potestatem
LEV|22|14|qui comederit de sanctificatis per ignorantiam addet quintam partem cum eo quod comedit et dabit sacerdoti in sanctuarium
LEV|22|15|nec contaminabunt sanctificata filiorum Israhel quae offerunt Domino
LEV|22|16|ne forte sustineant iniquitatem delicti sui cum sanctificata comederint ego Dominus qui sanctifico eos
LEV|22|17|locutus est Dominus ad Mosen dicens
LEV|22|18|loquere ad Aaron et filios eius et ad omnes filios Israhel dicesque ad eos homo de domo Israhel et de advenis qui habitant apud vos qui obtulerit oblationem suam vel vota solvens vel sponte offerens quicquid illud obtulerit in holocaustum Domini
LEV|22|19|ut offeratur per vos masculus inmaculatus erit ex bubus et ex ovibus et ex capris
LEV|22|20|si maculam habuerit non offeretis neque erit acceptabile
LEV|22|21|homo qui obtulerit victimam pacificorum Domino vel vota solvens vel sponte offerens tam de bubus quam de ovibus inmaculatum offeret ut acceptabile sit omnis macula non erit in eo
LEV|22|22|si caecum fuerit si fractum si cicatricem habens si papulas aut scabiem vel inpetiginem non offeretis ea Domino neque adolebitis ex eis super altare Domini
LEV|22|23|bovem et ovem aure et cauda amputatis voluntarie offerre potes votum autem ex his solvi non potest
LEV|22|24|omne animal quod vel contritis vel tunsis vel sectis ablatisque testiculis est non offeretis Domino et in terra vestra hoc omnino ne faciatis
LEV|22|25|de manu alienigenae non offeretis panes Deo vestro et quicquid aliud dare voluerint quia corrupta et maculata sunt omnia non suscipietis ea
LEV|22|26|locutusque est Dominus ad Mosen dicens
LEV|22|27|bos ovis et capra cum genita fuerint septem diebus erunt sub ubere matris suae die autem octavo et deinceps offerri poterunt Domino
LEV|22|28|sive illa bos sive ovis non immolabuntur una die cum fetibus suis
LEV|22|29|si immolaveritis hostiam pro gratiarum actione Domino ut possit esse placabilis
LEV|22|30|eodem die comedetis eam non remanebit quicquam in mane alterius diei ego Dominus
LEV|22|31|custodite mandata mea et facite ea ego Dominus
LEV|22|32|ne polluatis nomen meum sanctum ut sanctificer in medio filiorum Israhel ego Dominus qui sanctifico vos
LEV|22|33|et eduxi de terra Aegypti ut essem vobis in Deum ego Dominus
LEV|23|1|locutus est Dominus ad Mosen dicens
LEV|23|2|loquere filiis Israhel et dices ad eos hae sunt feriae Domini quas vocabitis sanctas
LEV|23|3|sex diebus facietis opus dies septimus quia sabbati requies est vocabitur sanctus omne opus non facietis in eo sabbatum Domini est in cunctis habitationibus vestris
LEV|23|4|hae sunt ergo feriae Domini sanctae quas celebrare debetis temporibus suis
LEV|23|5|mense primo quartadecima die mensis ad vesperum phase Domini est
LEV|23|6|et quintadecima die mensis huius sollemnitas azymorum Domini est septem diebus azyma comedetis
LEV|23|7|dies primus erit vobis celeberrimus sanctusque omne opus servile non facietis in eo
LEV|23|8|sed offeretis sacrificium in igne Domino septem diebus dies autem septimus erit celebrior et sanctior nullumque servile opus fiet in eo
LEV|23|9|locutusque est Dominus ad Mosen dicens
LEV|23|10|loquere filiis Israhel et dices ad eos cum ingressi fueritis terram quam ego dabo vobis et messueritis segetem feretis manipulos spicarum primitias messis vestrae ad sacerdotem
LEV|23|11|qui elevabit fasciculum coram Domino ut acceptabile sit pro vobis altero die sabbati et sanctificabit illum
LEV|23|12|atque in eodem die quo manipulus consecratur caedetur agnus inmaculatus anniculus in holocaustum Domini
LEV|23|13|et libamenta offerentur cum eo duae decimae similae conspersae oleo in incensum Domini odoremque suavissimum liba quoque vini quarta pars hin
LEV|23|14|panem et pulentam et pultes non comedetis ex segete usque ad diem qua offeratis ex ea Deo vestro praeceptum est sempiternum in generationibus cunctisque habitaculis vestris
LEV|23|15|numerabitis ergo ab altero die sabbati in quo obtulistis manipulum primitiarum septem ebdomadas plenas
LEV|23|16|usque ad alteram diem expletionis ebdomadae septimae id est quinquaginta dies et sic offeretis sacrificium novum Domino
LEV|23|17|ex omnibus habitaculis vestris panes primitiarum duos de duabus decimis similae fermentatae quos coquetis in primitias Domini
LEV|23|18|offeretisque cum panibus septem agnos inmaculatos anniculos et vitulum de armento unum et arietes duos et erunt in holocausto cum libamentis suis in odorem suavissimum Domino
LEV|23|19|facietis et hircum pro peccato duosque agnos anniculos hostias pacificorum
LEV|23|20|cumque elevaverit eos sacerdos cum panibus primitiarum coram Domino cedent in usum eius
LEV|23|21|et vocabitis hunc diem celeberrimum atque sanctissimum omne opus servile non facietis in eo legitimum sempiternum erit in cunctis habitaculis et generationibus vestris
LEV|23|22|postquam autem messueritis segetem terrae vestrae non secabitis eam usque ad solum nec remanentes spicas colligetis sed pauperibus et peregrinis dimittetis eas ego Dominus Deus vester
LEV|23|23|locutusque est Dominus ad Mosen dicens
LEV|23|24|loquere filiis Israhel mense septimo prima die mensis erit vobis sabbatum memorabile clangentibus tubis et vocabitur sanctum
LEV|23|25|omne opus servile non facietis in eo et offeretis holocaustum Domino
LEV|23|26|locutusque est Dominus ad Mosen dicens
LEV|23|27|decimo die mensis huius septimi dies expiationum erit celeberrimus et vocabitur sanctus adfligetisque animas vestras in eo et offeretis holocaustum Domino
LEV|23|28|omne opus non facietis in tempore diei huius quia dies propitiationis est ut propitietur vobis Dominus Deus vester
LEV|23|29|omnis anima quae adflicta non fuerit die hoc peribit de populis suis
LEV|23|30|et quae operis quippiam fecerit delebo eam de populo suo
LEV|23|31|nihil ergo operis facietis in eo legitimum sempiternum erit vobis in cunctis generationibus et habitationibus vestris
LEV|23|32|sabbatum requietionis est adfligetis animas vestras die nono mensis a vespero usque ad vesperum celebrabitis sabbata vestra
LEV|23|33|et locutus est Dominus ad Mosen dicens
LEV|23|34|loquere filiis Israhel a quintodecimo die mensis huius septimi erunt feriae tabernaculorum septem diebus Domino
LEV|23|35|dies primus vocabitur celeberrimus atque sanctissimus omne opus servile non facietis
LEV|23|36|et septem diebus offeretis holocausta Domino dies quoque octavus erit celeberrimus atque sanctissimus et offeretis holocaustum Domino est enim coetus atque collectae omne opus servile non facietis in eo
LEV|23|37|hae sunt feriae Domini quas vocabitis celeberrimas et sanctissimas offeretisque in eis oblationes Domino holocausta et libamenta iuxta ritum uniuscuiusque diei
LEV|23|38|exceptis sabbatis Domini donisque vestris et quae offertis ex voto vel quae sponte tribuitis Domino
LEV|23|39|a quintodecimo ergo die mensis septimi quando congregaveritis omnes fructus terrae vestrae celebrabitis ferias Domini septem diebus die primo et die octavo erit sabbatum id est requies
LEV|23|40|sumetisque vobis die primo fructus arboris pulcherrimae spatulasque palmarum et ramos ligni densarum frondium et salices de torrente et laetabimini coram Domino Deo vestro
LEV|23|41|celebrabitisque sollemnitatem eius septem diebus per annum legitimum sempiternum erit in generationibus vestris mense septimo festa celebrabitis
LEV|23|42|et habitabitis in umbraculis septem diebus omnis qui de genere est Israhel manebit in tabernaculis
LEV|23|43|ut discant posteri vestri quod in tabernaculis habitare fecerim filios Israhel cum educerem eos de terra Aegypti ego Dominus Deus vester
LEV|23|44|locutusque est Moses super sollemnitatibus Domini ad filios Israhel
LEV|24|1|et locutus est Dominus ad Mosen dicens
LEV|24|2|praecipe filiis Israhel ut adferant tibi oleum de olivis purissimum ac lucidum ad concinnandas lucernas iugiter
LEV|24|3|extra velum testimonii in tabernaculo foederis ponetque eas Aaron a vespere usque in mane coram Domino cultu rituque perpetuo in generationibus vestris
LEV|24|4|super candelabro mundissimo ponentur semper in conspectu Domini
LEV|24|5|accipies quoque similam et coques ex ea duodecim panes qui singuli habebunt duas decimas
LEV|24|6|quorum senos altrinsecus super mensam purissimam coram Domino statues
LEV|24|7|et pones super eos tus lucidissimum ut sit panis in monumentum oblationis Domini
LEV|24|8|per singula sabbata mutabuntur coram Domino suscepti a filiis Israhel foedere sempiterno
LEV|24|9|eruntque Aaron et filiorum eius ut comedant eos in loco sancto quia sanctum sanctorum est de sacrificiis Domini iure perpetuo
LEV|24|10|ecce autem egressus filius mulieris israhelitis quem pepererat de viro aegyptio inter filios Israhel iurgatus est in castris cum viro israhelite
LEV|24|11|cumque blasphemasset nomen et maledixisset ei adductus est ad Mosen vocabatur autem mater eius Salumith filia Dabri de tribu Dan
LEV|24|12|miseruntque eum in carcerem donec nossent quid iuberet Dominus
LEV|24|13|qui locutus est ad Mosen
LEV|24|14|dicens educ blasphemum extra castra et ponant omnes qui audierunt manus suas super caput eius et lapidet eum populus universus
LEV|24|15|et ad filios Israhel loqueris homo qui maledixerit Deo suo portabit peccatum suum
LEV|24|16|et qui blasphemaverit nomen Domini morte moriatur lapidibus opprimet eum omnis multitudo sive ille civis seu peregrinus fuerit qui blasphemaverit nomen Domini morte moriatur
LEV|24|17|qui percusserit et occiderit hominem morte moriatur
LEV|24|18|qui percusserit animal reddat vicarium id est animam pro anima
LEV|24|19|qui inrogaverit maculam cuilibet civium suorum sicut fecit fiet ei
LEV|24|20|fracturam pro fractura oculum pro oculo dentem pro dente restituet qualem inflixerit maculam talem sustinere cogetur
LEV|24|21|qui percusserit iumentum reddet aliud qui percusserit hominem punietur
LEV|24|22|aequum iudicium sit inter vos sive peregrinus sive civis peccaverit quia ego sum Dominus Deus vester
LEV|24|23|locutusque est Moses ad filios Israhel et eduxerunt eum qui blasphemaverat extra castra ac lapidibus oppresserunt feceruntque filii Israhel sicut praeceperat Dominus Mosi
LEV|25|1|locutusque est Dominus ad Mosen in monte Sinai dicens
LEV|25|2|loquere filiis Israhel et dices ad eos quando ingressi fueritis terram quam ego dabo vobis sabbatizet sabbatum Domini
LEV|25|3|sex annis seres agrum tuum et sex annis putabis vineam tuam colligesque fructus eius
LEV|25|4|septimo autem anno sabbatum erit terrae requietionis Domini agrum non seres et vineam non putabis
LEV|25|5|quae sponte gignit humus non metes et uvas primitiarum tuarum non colliges quasi vindemiam annus enim requietionis terrae est
LEV|25|6|sed erunt vobis in cibum tibi et servo tuo ancillae et mercennario tuo et advenae qui peregrinantur apud te
LEV|25|7|iumentis tuis et pecoribus omnia quae nascuntur praebebunt cibum
LEV|25|8|numerabis quoque tibi septem ebdomades annorum id est septem septies quae simul faciunt annos quadraginta novem
LEV|25|9|et clanges bucina mense septimo decima die mensis propitiationis tempore in universa terra vestra
LEV|25|10|sanctificabisque annum quinquagesimum et vocabis remissionem cunctis habitatoribus terrae tuae ipse est enim iobeleus revertetur homo ad possessionem suam et unusquisque rediet ad familiam pristinam
LEV|25|11|quia iobeleus est et quinquagesimus annus non seretis neque metetis sponte in agro nascentia et primitias vindemiae non colligetis
LEV|25|12|ob sanctificationem iobelei sed statim ablata comedetis
LEV|25|13|anno iobelei redient omnes ad possessiones suas
LEV|25|14|quando vendes quippiam civi tuo vel emes ab eo ne contristes fratrem tuum sed iuxta numerum annorum iobelei emes ab eo
LEV|25|15|et iuxta supputationem frugum vendet tibi
LEV|25|16|quanto plus anni remanserint post iobeleum tanto crescet et pretium et quanto minus temporis numeraveris tanto minoris et emptio constabit tempus enim frugum vendet tibi
LEV|25|17|nolite adfligere contribules vestros sed timeat unusquisque Deum suum quia ego Dominus Deus vester
LEV|25|18|facite praecepta mea et iudicia custodite et implete ea ut habitare possitis in terra absque ullo pavore
LEV|25|19|et gignat vobis humus fructus suos quibus vescamini usque ad saturitatem nullius impetum formidantes
LEV|25|20|quod si dixeritis quid comedemus anno septimo si non seruerimus neque collegerimus fruges nostras
LEV|25|21|dabo benedictionem meam vobis anno sexto et faciet fructus trium annorum
LEV|25|22|seretisque anno octavo et comedetis veteres fruges usque ad nonum annum donec nova nascantur edetis vetera
LEV|25|23|terra quoque non veniet in perpetuum quia mea est et vos advenae et coloni mei estis
LEV|25|24|unde cuncta regio possessionis vestrae sub redemptionis condicione vendetur
LEV|25|25|si adtenuatus frater tuus vendiderit possessiunculam suam et voluerit propinquus eius potest redimere quod ille vendiderat
LEV|25|26|sin autem non habuerit proximum et ipse pretium ad redimendum potuerit invenire
LEV|25|27|conputabuntur fructus ex eo tempore quo vendidit et quod reliquum est reddet emptori sicque recipiet possessionem suam
LEV|25|28|quod si non invenerit manus eius ut reddat pretium habebit emptor quod emerat usque ad annum iobeleum in ipso enim omnis venditio redit ad dominum et ad possessorem pristinum
LEV|25|29|qui vendiderit domum intra urbis muros habebit licentiam redimendi donec unus impleatur annus
LEV|25|30|si non redemerit et anni circulus fuerit evolutus emptor possidebit eam et posteri eius in perpetuum et redimi non poterit etiam in iobeleo
LEV|25|31|sin autem in villa fuerit domus quae muros non habet agrorum iure vendetur si ante redempta non fuerit in iobeleo revertetur ad dominum
LEV|25|32|aedes Levitarum quae in urbibus sunt semper possunt redimi
LEV|25|33|si redemptae non fuerint in iobeleo revertentur ad dominos quia domus urbium leviticarum pro possessionibus sunt inter filios Israhel
LEV|25|34|suburbana autem eorum non venient quia possessio sempiterna est
LEV|25|35|si adtenuatus fuerit frater tuus et infirmus manu et susceperis eum quasi advenam et peregrinum et vixerit tecum
LEV|25|36|ne accipias usuras ab eo nec amplius quam dedisti time Deum tuum ut vivere possit frater tuus apud te
LEV|25|37|pecuniam tuam non dabis ei ad usuram et frugum superabundantiam non exiges
LEV|25|38|ego Dominus Deus vester qui eduxi vos de terra Aegypti ut darem vobis terram Chanaan et essem vester Deus
LEV|25|39|si paupertate conpulsus vendiderit se tibi frater tuus non eum opprimes servitute famulorum
LEV|25|40|sed quasi mercennarius et colonus erit usque ad annum iobeleum operabitur apud te
LEV|25|41|et postea egredietur cum liberis suis et revertetur ad cognationem et ad possessionem patrum suorum
LEV|25|42|mei enim servi sunt et ego eduxi eos de terra Aegypti non venient condicione servorum
LEV|25|43|ne adfligas eum per potentiam sed metuito Deum tuum
LEV|25|44|servus et ancilla sint vobis de nationibus quae in circuitu vestro sunt
LEV|25|45|et de advenis qui peregrinantur apud vos vel qui ex his nati fuerint in terra vestra hos habebitis famulos
LEV|25|46|et hereditario iure transmittetis ad posteros ac possidebitis in aeternum fratres autem vestros filios Israhel ne opprimatis per potentiam
LEV|25|47|si invaluerit apud vos manus advenae atque peregrini et adtenuatus frater tuus vendiderit se ei aut cuiquam de stirpe eius
LEV|25|48|post venditionem potest redimi qui voluerit ex fratribus suis redimet eum
LEV|25|49|et patruus et patruelis et consanguineus et adfinis sin autem et ipse potuerit redimet se
LEV|25|50|supputatis dumtaxat annis a tempore venditionis suae usque ad annum iobeleum et pecunia qua venditus fuerat iuxta annorum numerum et rationem mercennarii supputata
LEV|25|51|si plures fuerint anni qui remanent usque ad iobeleum secundum hos reddet et pretium
LEV|25|52|si pauci ponet rationem cum eo iuxta annorum numerum et reddet emptori quod reliquum est annorum
LEV|25|53|quibus ante servivit mercedibus inputatis non adfliget eum violenter in conspectu tuo
LEV|25|54|quod si per haec redimi non potuerit anno iobeleo egredietur cum liberis suis
LEV|25|55|mei sunt enim servi filii Israhel quos eduxi de terra Aegypti
LEV|26|1|ego Dominus Deus vester non facietis vobis idolum et sculptile nec titulos erigetis nec insignem lapidem ponetis in terra vestra ut adoretis eum ego enim sum Dominus Deus vester
LEV|26|2|custodite sabbata mea et pavete ad sanctuarium meum ego Dominus
LEV|26|3|si in praeceptis meis ambulaveritis et mandata mea custodieritis et feceritis ea dabo vobis pluvias temporibus suis
LEV|26|4|et terra gignet germen suum et pomis arbores replebuntur
LEV|26|5|adprehendet messium tritura vindemiam et vindemia occupabit sementem et comedetis panem vestrum in saturitatem et absque pavore habitabitis in terra vestra
LEV|26|6|dabo pacem in finibus vestris dormietis et non erit qui exterreat auferam malas bestias et gladius non transibit terminos vestros
LEV|26|7|persequemini inimicos vestros et corruent coram vobis
LEV|26|8|persequentur quinque de vestris centum alienos et centum ex vobis decem milia cadent inimici vestri in conspectu vestro gladio
LEV|26|9|respiciam vos et crescere faciam multiplicabimini et firmabo pactum meum vobiscum
LEV|26|10|comedetis vetustissima veterum et vetera novis supervenientibus proicietis
LEV|26|11|ponam tabernaculum meum in medio vestri et non abiciet vos anima mea
LEV|26|12|ambulabo inter vos et ero vester Deus vosque eritis populus meus
LEV|26|13|ego Dominus Deus vester qui eduxi vos de terra Aegyptiorum ne serviretis eis et qui confregi catenas cervicum vestrarum ut incederetis erecti
LEV|26|14|quod si non audieritis me nec feceritis omnia mandata mea
LEV|26|15|si spreveritis leges meas et iudicia mea contempseritis ut non faciatis ea quae a me constituta sunt et ad irritum perducatis pactum meum
LEV|26|16|ego quoque haec faciam vobis visitabo vos velociter in egestate et ardore qui conficiat oculos vestros et consumat animas frustra seretis sementem quae ab hostibus devorabitur
LEV|26|17|ponam faciem meam contra vos et corruetis coram hostibus vestris et subiciemini his qui oderunt vos fugietis nemine persequente
LEV|26|18|sin autem nec sic oboedieritis mihi addam correptiones vestras septuplum propter peccata vestra
LEV|26|19|et conteram superbiam duritiae vestrae daboque caelum vobis desuper sicut ferrum et terram aeneam
LEV|26|20|consumetur in cassum labor vester non proferet terra germen nec arbores poma praebebunt
LEV|26|21|si ambulaveritis ex adverso mihi nec volueritis audire me addam plagas vestras usque in septuplum propter peccata vestra
LEV|26|22|emittamque in vos bestias agri quae consumant et vos et pecora vestra et ad paucitatem cuncta redigant desertaeque fiant viae vestrae
LEV|26|23|quod si nec sic volueritis recipere disciplinam sed ambulaveritis ex adverso mihi
LEV|26|24|ego quoque contra vos adversus incedam et percutiam vos septies propter peccata vestra
LEV|26|25|inducamque super vos gladium ultorem foederis mei cumque confugeritis in urbes mittam pestilentiam in medio vestri et trademini hostium manibus
LEV|26|26|postquam confregero baculum panis vestri ita ut decem mulieres in uno clibano coquant panes et reddant eos ad pondus et comedetis et non saturabimini
LEV|26|27|sin autem nec per haec audieritis me sed ambulaveritis contra me
LEV|26|28|et ego incedam adversum vos in furore contrario et corripiam vos septem plagis propter peccata vestra
LEV|26|29|ita ut comedatis carnes filiorum et filiarum vestrarum
LEV|26|30|destruam excelsa vestra et simulacra confringam cadetis inter ruinas idolorum vestrorum et abominabitur vos anima mea
LEV|26|31|in tantum ut urbes vestras redigam in solitudinem et deserta faciam sanctuaria vestra nec recipiam ultra odorem suavissimum
LEV|26|32|disperdamque terram vestram et stupebunt super ea inimici vestri cum habitatores illius fuerint
LEV|26|33|vos autem dispergam in gentes et evaginabo post vos gladium eritque terra vestra deserta et civitates dirutae
LEV|26|34|tunc placebunt terrae sabbata sua cunctis diebus solitudinis suae quando fueritis
LEV|26|35|in terra hostili sabbatizabit et requiescet in sabbatis solitudinis suae eo quod non requieverit in sabbatis vestris quando habitabatis in ea
LEV|26|36|et qui de vobis remanserint dabo pavorem in cordibus eorum in regionibus hostium terrebit eos sonitus folii volantis et ita fugient quasi gladium cadent nullo sequente
LEV|26|37|et corruent singuli super fratres suos quasi bella fugientes nemo vestrum inimicis audebit resistere
LEV|26|38|peribitis inter gentes et hostilis vos terra consumet
LEV|26|39|quod si et de his aliqui remanserint tabescent in iniquitatibus suis in terra inimicorum suorum et propter peccata patrum suorum et sua adfligentur
LEV|26|40|donec confiteantur iniquitates suas et maiorum suorum quibus praevaricati sunt in me et ambulaverunt ex adverso mihi
LEV|26|41|ambulabo igitur et ego contra eos et inducam illos in terram hostilem donec erubescat incircumcisa mens eorum tunc orabunt pro impietatibus suis
LEV|26|42|et recordabor foederis mei quod pepigi cum Iacob et Isaac et Abraham terrae quoque memor ero
LEV|26|43|quae cum relicta fuerit ab eis conplacebit sibi in sabbatis suis patiens solitudinem propter illos ipsi vero rogabunt pro peccatis suis eo quod abiecerint iudicia mea et leges meas despexerint
LEV|26|44|et tamen etiam cum essent in terra hostili non penitus abieci eos neque sic despexi ut consumerentur et irritum facerem pactum meum cum eis ego enim sum Dominus Deus eorum
LEV|26|45|et recordabor foederis mei pristini quando eduxi eos de terra Aegypti in conspectu gentium ut essem Deus eorum ego Dominus Deus haec sunt praecepta atque iudicia et leges quas dedit Dominus inter se et inter filios Israhel in monte Sinai per manum Mosi
LEV|26|46|
LEV|27|1|locutusque est Dominus ad Mosen dicens
LEV|27|2|loquere filiis Israhel et dices ad eos homo qui votum fecerit et spoponderit Deo animam suam sub aestimatione dabit pretium
LEV|27|3|si fuerit masculus a vicesimo usque ad sexagesimum annum dabit quinquaginta siclos argenti ad mensuram sanctuarii
LEV|27|4|si mulier triginta
LEV|27|5|a quinto autem anno usque ad vicesimum masculus dabit viginti siclos femina decem
LEV|27|6|ab uno mense usque ad annum quintum pro masculo dabuntur quinque sicli pro femina tres
LEV|27|7|sexagenarius et ultra masculus dabit quindecim siclos femina decem
LEV|27|8|si pauper fuerit et aestimationem reddere non valebit stabit coram sacerdote et quantum ille aestimaverit et viderit eum posse reddere tantum dabit
LEV|27|9|animal autem quod immolari potest Domino si quis voverit sanctum erit
LEV|27|10|et mutari non poterit id est nec melius malo nec peius bono quod si mutaverit et ipsum quod mutatum est et illud pro quo mutatum est consecratum erit Domino
LEV|27|11|animal inmundum quod immolari Domino non potest si quis voverit adducetur ante sacerdotem
LEV|27|12|qui diiudicans utrum bonum an malum sit statuet pretium
LEV|27|13|quod si dare voluerit is qui offert addet supra aestimationis quintam partem
LEV|27|14|homo si voverit domum suam et sanctificaverit Domino considerabit eam sacerdos utrum bona an mala sit et iuxta pretium quod ab eo fuerit constitutum venundabitur
LEV|27|15|sin autem ille qui voverat voluerit redimere eam dabit quintam partem aestimationis supra et habebit domum
LEV|27|16|quod si agrum possessionis suae voverit et consecraverit Domino iuxta mensuram sementis aestimabitur pretium si triginta modiis hordei seritur terra quinquaginta siclis veniet argenti
LEV|27|17|si statim ab anno incipientis iobelei voverit agrum quanto valere potest tanto aestimabitur
LEV|27|18|sin autem post aliquantum temporis supputabit sacerdos pecuniam iuxta annorum qui reliqui sunt numerum usque ad iobeleum et detrahetur ex pretio
LEV|27|19|quod si voluerit redimere agrum ille qui voverat addet quintam partem aestimatae pecuniae et possidebit eum
LEV|27|20|sin autem noluerit redimere sed alteri cuilibet fuerit venundatus ultra eum qui voverat redimere non poterit
LEV|27|21|quia cum iobelei venerit dies sanctificatus erit Domino et possessio consecrata ad ius pertinet sacerdotum
LEV|27|22|si ager emptus et non de possessione maiorum sanctificatus fuerit Domino
LEV|27|23|supputabit sacerdos iuxta annorum numerum usque ad iobeleum pretium et dabit ille qui voverat eum Domino
LEV|27|24|in iobeleo autem revertetur ad priorem dominum qui vendiderat eum et habuerat in sortem possessionis suae
LEV|27|25|omnis aestimatio siclo sanctuarii ponderabitur siclus viginti obolos habet
LEV|27|26|primogenita quae ad Dominum pertinent nemo sanctificare poterit et vovere sive bos sive ovis fuerit Domini sunt
LEV|27|27|quod si inmundum est animal redimet qui obtulit iuxta aestimationem tuam et addet quintam partem pretii si redimere noluerit vendetur alteri quantocumque a te fuerit aestimatum
LEV|27|28|omne quod Domino consecratur sive homo fuerit sive animal sive ager non veniet nec redimi poterit quicquid semel fuerit consecratum sanctum sanctorum erit Domino
LEV|27|29|et omnis consecratio quae offertur ab homine non redimetur sed morte morietur
LEV|27|30|omnes decimae terrae sive de frugibus sive de pomis arborum Domini sunt et illi sanctificantur
LEV|27|31|si quis autem voluerit redimere decimas suas addet quintam partem earum
LEV|27|32|omnium decimarum boves et oves et caprae quae sub pastoris virga transeunt quicquid decimum venerit sanctificabitur Domino
LEV|27|33|non eligetur nec bonum nec malum nec altero commutabitur si quis mutaverit et quod mutatum est et pro quo mutatum est sanctificabitur Domino et non redimetur
LEV|27|34|haec sunt praecepta quae mandavit Dominus Mosi ad filios Israhel in monte Sinai
NUM|1|1|locutusque est Dominus ad Mosen in deserto Sinai in tabernaculo foederis prima die mensis secundi anno altero egressionis eorum ex Aegypto dicens
NUM|1|2|tollite summam universae congregationis filiorum Israhel per cognationes et domos suas et nomina singulorum quicquid sexus est masculini
NUM|1|3|a vicesimo anno et supra omnium virorum fortium ex Israhel et numerabitis eos per turmas suas tu et Aaron
NUM|1|4|eruntque vobiscum principes tribuum ac domorum in cognationibus suis
NUM|1|5|quorum ista sunt nomina de Ruben Elisur filius Sedeur
NUM|1|6|de Symeon Salamihel filius Surisaddai
NUM|1|7|de Iuda Naasson filius Aminadab
NUM|1|8|de Isachar Nathanahel filius Suar
NUM|1|9|de Zabulon Heliab filius Helon
NUM|1|10|filiorum autem Ioseph de Ephraim Helisama filius Ammiud de Manasse Gamalihel filius Phadassur
NUM|1|11|de Beniamin Abidan filius Gedeonis
NUM|1|12|de Dan Ahiezer filius Amisaddai
NUM|1|13|de Aser Phegihel filius Ochran
NUM|1|14|de Gad Heliasaph filius Duhel
NUM|1|15|de Nepthali Ahira filius Henan
NUM|1|16|hii nobilissimi principes multitudinis per tribus et cognationes suas et capita exercitus Israhel
NUM|1|17|quos tulerunt Moses et Aaron cum omni vulgi multitudine
NUM|1|18|et congregaverunt primo die mensis secundi recensentes eos per cognationes et domos ac familias et capita et nomina singulorum a vicesimo anno et supra
NUM|1|19|sicut praeceperat Dominus Mosi numeratique sunt in deserto Sinai
NUM|1|20|de Ruben primogenito Israhelis per generationes et familias ac domos suas et nomina capitum singulorum omne quod sexus est masculini a vicesimo anno et supra procedentium ad bellum
NUM|1|21|quadraginta sex milia quingenti
NUM|1|22|de filiis Symeon per generationes et familias ac domos cognationum suarum recensiti sunt per nomina et capita singulorum omne quod sexus est masculini a vicesimo anno et supra procedentium ad bellum
NUM|1|23|quinquaginta novem milia trecenti
NUM|1|24|de filiis Gad per generationes et familias ac domos cognationum suarum recensiti sunt per nomina singulorum a viginti annis et supra omnes qui ad bella procederent
NUM|1|25|quadraginta quinque milia sescenti quinquaginta
NUM|1|26|de filiis Iuda per generationes et familias ac domos cognationum suarum per nomina singulorum a vicesimo anno et supra omnes qui poterant ad bella procedere
NUM|1|27|recensiti sunt septuaginta quattuor milia sescenti
NUM|1|28|de filiis Isachar per generationes et familias ac domos cognationum suarum per nomina singulorum a vicesimo anno et supra omnes qui ad bella procederent
NUM|1|29|recensiti sunt quinquaginta quattuor milia quadringenti
NUM|1|30|de filiis Zabulon per generationes et familias ac domos cognationum suarum recensiti sunt per nomina singulorum a vicesimo anno et supra omnes qui poterant ad bella procedere
NUM|1|31|quinquaginta septem milia quadringenti
NUM|1|32|de filiis Ioseph filiorum Ephraim per generationes et familias ac domos cognationum suarum recensiti sunt per nomina singulorum a vicesimo anno et supra omnes qui poterant ad bella procedere
NUM|1|33|quadraginta milia quingenti
NUM|1|34|porro filiorum Manasse per generationes et familias ac domos cognationum suarum recensiti sunt per nomina singulorum a viginti annis et supra omnes qui poterant ad bella procedere
NUM|1|35|triginta duo milia ducenti
NUM|1|36|de filiis Beniamin per generationes et familias ac domos cognationum suarum recensiti sunt nominibus singulorum a vicesimo anno et supra omnes qui poterant ad bella procedere
NUM|1|37|triginta quinque milia quadringenti
NUM|1|38|de filiis Dan per generationes et familias ac domos cognationum suarum recensiti sunt nominibus singulorum a vicesimo anno et supra omnes qui poterant ad bella procedere
NUM|1|39|sexaginta duo milia septingenti
NUM|1|40|de filiis Aser per generationes et familias ac domos cognationum suarum recensiti sunt per nomina singulorum a vicesimo anno et supra omnes qui poterant ad bella procedere
NUM|1|41|quadraginta milia et mille quingenti
NUM|1|42|de filiis Nepthali per generationes et familias ac domos cognationum suarum recensiti sunt nominibus singulorum a vicesimo anno et supra omnes qui poterant ad bella procedere
NUM|1|43|quinquaginta tria milia quadringenti
NUM|1|44|hii sunt quos numeraverunt Moses et Aaron et duodecim principes Israhel singulos per domos cognationum suarum
NUM|1|45|fueruntque omnes filiorum Israhel per domos et familias suas a vicesimo anno et supra qui poterant ad bella procedere
NUM|1|46|sescenta tria milia virorum quingenti quinquaginta
NUM|1|47|Levitae autem in tribu familiarum suarum non sunt numerati cum eis
NUM|1|48|locutusque est Dominus ad Mosen dicens
NUM|1|49|tribum Levi noli numerare neque ponas summam eorum cum filiis Israhel
NUM|1|50|sed constitue eos super tabernaculum testimonii cuncta vasa eius et quicquid ad caerimonias pertinet ipsi portabunt tabernaculum et omnia utensilia eius et erunt in ministerio ac per gyrum tabernaculi metabuntur
NUM|1|51|cum proficiscendum fuerit deponent Levitae tabernaculum cum castra metanda erigent quisquis externorum accesserit occidetur
NUM|1|52|metabuntur autem castra filii Israhel unusquisque per turmas et cuneos atque exercitum suum
NUM|1|53|porro Levitae per gyrum tabernaculi figent tentoria ne fiat indignatio super multitudinem filiorum Israhel et excubabunt in custodiis tabernaculi testimonii
NUM|1|54|fecerunt ergo filii Israhel iuxta omnia quae praeceperat Dominus Mosi
NUM|2|1|locutusque est Dominus ad Mosen et Aaron dicens
NUM|2|2|singuli per turmas signa atque vexilla et domos cognationum suarum castrametabuntur filiorum Israhel per gyrum tabernaculi foederis
NUM|2|3|ad orientem Iudas figet tentoria per turmas exercitus sui eritque princeps filiorum eius Naasson filius Aminadab
NUM|2|4|et omnis de stirpe eius summa pugnantium septuaginta quattuor milia sescentorum
NUM|2|5|iuxta eum castrametati sunt de tribu Isachar quorum princeps fuit Nathanahel filius Suar
NUM|2|6|et omnis numerus pugnatorum eius quinquaginta quattuor milia quadringenti
NUM|2|7|in tribu Zabulon princeps fuit Heliab filius Helon
NUM|2|8|omnis de stirpe eius exercitus pugnatorum quinquaginta septem milia quadringenti
NUM|2|9|universi qui in castris Iudae adnumerati sunt fuerunt centum octoginta sex milia quadringenti et per turmas suas primi egredientur
NUM|2|10|in castris filiorum Ruben ad meridianam plagam erit princeps Elisur filius Sedeur
NUM|2|11|et cunctus exercitus pugnatorum eius qui numerati sunt quadraginta sex milia quingenti
NUM|2|12|iuxta eum castrametati sunt de tribu Symeon quorum princeps fuit Salamihel filius Surisaddai
NUM|2|13|et cunctus exercitus pugnatorum eius qui numerati sunt quinquaginta novem milia trecenti
NUM|2|14|in tribu Gad princeps fuit Heliasaph filius Duhel
NUM|2|15|et cunctus exercitus pugnatorum eius qui numerati sunt quadraginta quinque milia sescenti quinquaginta
NUM|2|16|omnes qui recensiti sunt in castris Ruben centum quinquaginta milia et mille quadringenti quinquaginta per turmas suas in secundo loco proficiscentur
NUM|2|17|levabitur autem tabernaculum testimonii per officia Levitarum et turmas eorum quomodo erigetur ita et deponetur singuli per loca et ordines suos proficiscentur
NUM|2|18|ad occidentalem plagam erunt castra filiorum Ephraim quorum princeps fuit Helisama filius Ammiud
NUM|2|19|cunctus exercitus pugnatorum eius qui numerati sunt quadraginta milia quingenti
NUM|2|20|et cum eis tribus filiorum Manasse quorum princeps fuit Gamalihel filius Phadassur
NUM|2|21|cunctus exercitus pugnatorum eius qui numerati sunt triginta duo milia ducenti
NUM|2|22|in tribu filiorum Beniamin princeps fuit Abidan filius Gedeonis
NUM|2|23|et cunctus exercitus pugnatorum eius qui recensiti sunt triginta quinque milia quadringenti
NUM|2|24|omnes qui numerati sunt in castris Ephraim centum octo milia centum per turmas suas tertii proficiscentur
NUM|2|25|ad aquilonis partem castrametati sunt filii Dan quorum princeps fuit Ahiezer filius Amisaddai
NUM|2|26|cunctus exercitus pugnatorum eius qui numerati sunt sexaginta duo milia septingenti
NUM|2|27|iuxta eum fixere tentoria de tribu Aser quorum princeps fuit Phegihel filius Ochran
NUM|2|28|cunctus exercitus pugnatorum eius qui numerati sunt quadraginta milia et mille quingenti
NUM|2|29|de tribu filiorum Nepthalim princeps fuit Ahira filius Henan
NUM|2|30|cunctus exercitus pugnatorum eius quinquaginta tria milia quadringenti
NUM|2|31|omnes qui numerati sunt in castris Dan fuerunt centum quinquaginta septem milia sescenti et novissimi proficiscentur
NUM|2|32|hic numerus filiorum Israhel per domos cognationum suarum et turmas divisi exercitus sescenta tria milia quingenti quinquaginta
NUM|2|33|Levitae autem non sunt numerati inter filios Israhel sic enim praecepit Dominus Mosi
NUM|2|34|feceruntque filii Israhel iuxta omnia quae mandaverat Dominus castrametati sunt per turmas suas et profecti per familias ac domos patrum suorum
NUM|3|1|haec sunt generationes Aaron et Mosi in die qua locutus est Dominus ad Mosen in monte Sinai
NUM|3|2|et haec nomina filiorum Aaron primogenitus eius Nadab dein Abiu et Eleazar et Ithamar
NUM|3|3|haec nomina filiorum Aaron sacerdotum qui uncti sunt et quorum repletae et consecratae manus ut sacerdotio fungerentur
NUM|3|4|mortui sunt Nadab et Abiu cum offerrent ignem alienum in conspectu Domini in deserto Sinai absque liberis functique sunt sacerdotio Eleazar et Ithamar coram Aaron patre suo
NUM|3|5|locutus est Dominus ad Mosen dicens
NUM|3|6|adplica tribum Levi et fac stare in conspectu Aaron sacerdotis ut ministrent ei et excubent
NUM|3|7|et observent quicquid ad cultum pertinet multitudinis coram tabernaculo testimonii
NUM|3|8|et custodiant vasa tabernaculi servientes in ministerio eius
NUM|3|9|dabisque dono Levitas
NUM|3|10|Aaron et filiis eius quibus traditi sunt a filiis Israhel Aaron autem et filios eius constitues super cultum sacerdotii externus qui ad ministrandum accesserit morietur
NUM|3|11|locutusque est Dominus ad Mosen dicens
NUM|3|12|ego tuli Levitas a filiis Israhel pro omni primogenito qui aperit vulvam in filiis Israhel eruntque Levitae mei
NUM|3|13|meum est enim omne primogenitum ex quo percussi primogenitos in terra Aegypti sanctificavi mihi quicquid primum nascitur in Israhel ab homine usque ad pecus mei sunt ego Dominus
NUM|3|14|locutus est Dominus ad Mosen in deserto Sinai dicens
NUM|3|15|numera filios Levi per domos patrum suorum et familias omnem masculum ab uno mense et supra
NUM|3|16|numeravit Moses ut praeceperat Dominus
NUM|3|17|et inventi sunt filii Levi per nomina sua Gerson et Caath et Merari
NUM|3|18|filii Gerson Lebni et Semei
NUM|3|19|filii Caath Amram et Iessaar Hebron et Ozihel
NUM|3|20|filii Merari Mooli et Musi
NUM|3|21|de Gerson fuere familiae duae lebnitica et semeitica
NUM|3|22|quarum numeratus est populus sexus masculini ab uno mense et supra septem milia quingentorum
NUM|3|23|hii post tabernaculum metabuntur ad occidentem
NUM|3|24|sub principe Eliasaph filio Lahel
NUM|3|25|et habebunt excubias in tabernaculo foederis
NUM|3|26|ipsum tabernaculum et operimentum eius tentorium quod trahitur ante fores tecti foederis et cortinas atrii tentorium quoque quod adpenditur in introitu atrii tabernaculi et quicquid ad ritum altaris pertinet funes tabernaculi et omnia utensilia eius
NUM|3|27|cognatio Caath habebit populos Amramitas et Iessaaritas et Hebronitas et Ozihelitas hae sunt familiae Caathitarum recensitae per nomina sua
NUM|3|28|omnes generis masculini ab uno mense et supra octo milia sescenti habebunt excubias sanctuarii
NUM|3|29|et castrametabuntur ad meridianam plagam
NUM|3|30|princepsque eorum erit Elisaphan filius Ozihel
NUM|3|31|et custodient arcam mensamque et candelabrum altaria et vasa sanctuarii in quibus ministratur et velum cunctamque huiuscemodi supellectilem
NUM|3|32|princeps autem principum Levitarum Eleazar filius Aaron sacerdotis erit super excubitores custodiae sanctuarii
NUM|3|33|at vero de Merari erunt populi Moolitae et Musitae recensiti per nomina sua
NUM|3|34|omnes generis masculini ab uno mense et supra sex milia ducenti
NUM|3|35|princeps eorum Surihel filius Abiahihel in plaga septentrionali castrametabuntur
NUM|3|36|erunt sub custodia eorum tabulae tabernaculi et vectes et columnae ac bases earum et omnia quae ad cultum huiuscemodi pertinent
NUM|3|37|columnaeque atrii per circuitum cum basibus suis et paxilli cum funibus
NUM|3|38|castrametabuntur ante tabernaculum foederis id est ad orientalem plagam Moses et Aaron cum filiis suis habentes custodiam sanctuarii in medio filiorum Israhel quisquis alienus accesserit morietur
NUM|3|39|omnes Levitae quos numeraverunt Moses et Aaron iuxta praeceptum Domini per familias suas in genere masculino a mense uno et supra fuerunt viginti duo milia
NUM|3|40|et ait Dominus ad Mosen numera primogenitos sexus masculini de filiis Israhel a mense uno et supra et habebis summam eorum
NUM|3|41|tollesque Levitas mihi pro omni primogenito filiorum Israhel ego sum Dominus et pecora eorum pro universis primogenitis pecoris filiorum Israhel
NUM|3|42|recensuit Moses sicut praeceperat Dominus primogenitos filiorum Israhel
NUM|3|43|et fuerunt masculi per nomina sua a mense uno et supra viginti duo milia ducenti septuaginta tres
NUM|3|44|locutusque est Dominus ad Mosen
NUM|3|45|tolle Levitas pro primogenitis filiorum Israhel et pecora Levitarum pro pecoribus eorum eruntque Levitae mei ego sum Dominus
NUM|3|46|in pretio autem ducentorum septuaginta trium qui excedunt numerum Levitarum de primogenitis filiorum Israhel
NUM|3|47|accipies quinque siclos per singula capita ad mensuram sanctuarii siclus habet obolos viginti
NUM|3|48|dabisque pecuniam Aaron et filiis eius pretium eorum qui supra sunt
NUM|3|49|tulit igitur Moses pecuniam eorum qui fuerant amplius et quos redemerant a Levitis
NUM|3|50|pro primogenitis filiorum Israhel mille trecentorum sexaginta quinque siclorum iuxta pondus sanctuarii
NUM|3|51|et dedit eam Aaroni et filiis eius iuxta verbum quod praeceperat sibi Dominus
NUM|4|1|locutusque est Dominus ad Mosen et Aaron dicens
NUM|4|2|tolle summam filiorum Caath de medio Levitarum per domos et familias suas
NUM|4|3|a tricesimo anno et supra usque ad quinquagesimum annum omnium qui ingrediuntur ut stent et ministrent in tabernaculo foederis
NUM|4|4|hic est cultus filiorum Caath tabernaculum foederis et sanctum sanctorum
NUM|4|5|ingredientur Aaron et filii eius quando movenda sunt castra et deponent velum quod pendet ante fores involventque eo arcam testimonii
NUM|4|6|et operient rursum velamine ianthinarum pellium extendentque desuper pallium totum hyacinthinum et inducent vectes
NUM|4|7|mensam quoque propositionis involvent hyacinthino pallio et ponent cum ea turibula et mortariola cyatos et crateras ad liba fundenda panes semper in ea erunt
NUM|4|8|extendentque desuper pallium coccineum quod rursum operient velamento ianthinarum pellium et inducent vectes
NUM|4|9|sument et pallium hyacinthinum quo operient candelabrum cum lucernis et forcipibus suis et emunctoriis et cunctis vasis olei quae ad concinnandas lucernas necessaria sunt
NUM|4|10|et super omnia ponent operimentum ianthinarum pellium et inducent vectes
NUM|4|11|nec non et altare aureum involvent hyacinthino vestimento et extendent desuper operimentum ianthinarum pellium inducentque vectes
NUM|4|12|omnia vasa quibus ministratur in sanctuario involvent hyacinthino pallio et extendent desuper operimentum ianthinarum pellium inducentque vectes
NUM|4|13|sed et altare mundabunt cinere et involvent illud purpureo vestimento
NUM|4|14|ponentque cum eo omnia vasa quibus in ministerio eius utuntur id est ignium receptacula fuscinulas ac tridentes uncinos et vatilla cuncta vasa altaris operient simul velamine ianthinarum pellium et inducent vectes
NUM|4|15|cumque involverint Aaron et filii eius sanctuarium et omnia vasa eius in commotione castrorum tunc intrabunt filii Caath ut portent involuta et non tangant vasa sanctuarii ne moriantur ista sunt onera filiorum Caath in tabernaculo foederis
NUM|4|16|super quos erit Eleazar filius Aaron sacerdotis ad cuius pertinet curam oleum ad concinnandas lucernas et conpositionis incensum et sacrificium quod semper offertur et oleum unctionis et quicquid ad cultum tabernaculi pertinet omniumque vasorum quae in sanctuario sunt
NUM|4|17|locutusque est Dominus ad Mosen et Aaron dicens
NUM|4|18|nolite perdere populum Caath de medio Levitarum
NUM|4|19|sed hoc facite eis ut vivant et non moriantur si tetigerint sancta sanctorum Aaron et filii eius intrabunt ipsique disponent opera singulorum et divident quid portare quis debeat
NUM|4|20|alii nulla curiositate videant quae sunt in sanctuario priusquam involvantur alioquin morientur
NUM|4|21|locutus est Dominus ad Mosen dicens
NUM|4|22|tolle summam etiam filiorum Gerson per domos ac familias et cognationes suas
NUM|4|23|a triginta annis et supra usque ad annos quinquaginta numera omnes qui ingrediuntur et ministrant in tabernaculo foederis
NUM|4|24|hoc est officium familiae Gersonitarum
NUM|4|25|ut portent cortinas tabernaculi et tectum foederis operimentum aliud et super omnia velamen ianthinum tentoriumque quod pendet in introitu foederis tabernaculi
NUM|4|26|cortinas atrii et velum in introitu quod est ante tabernaculum omnia quae ad altare pertinent funiculos et vasa ministerii
NUM|4|27|iubente Aaron et filiis eius portabunt filii Gerson et scient singuli cui debeant oneri mancipari
NUM|4|28|hic est cultus familiae Gersonitarum in tabernaculo foederis eruntque sub manu Ithamar filii Aaron sacerdotis
NUM|4|29|filios quoque Merari per familias et domos patrum suorum recensebis
NUM|4|30|a triginta annis et supra usque ad annos quinquaginta omnes qui ingrediuntur ad officium ministerii sui et cultum foederis testimonii
NUM|4|31|haec sunt onera eorum portabunt tabulas tabernaculi et vectes eius columnas et bases earum
NUM|4|32|columnas quoque atrii per circuitum cum basibus et paxillis et funibus suis omnia vasa et supellectilem ad numerum accipient sicque portabunt
NUM|4|33|hoc est officium familiae Meraritarum et ministerium in tabernaculo foederis eruntque sub manu Ithamar filii Aaron sacerdotis
NUM|4|34|recensuerunt igitur Moses et Aaron et principes synagogae filios Caath per cognationes et domos patrum suorum
NUM|4|35|a triginta annis et supra usque ad annum quinquagesimum omnes qui ingrediuntur ad ministerium tabernaculi foederis
NUM|4|36|et inventi sunt duo milia septingenti quinquaginta
NUM|4|37|hic est numerus populi Caath qui intrat tabernaculum foederis hos numeravit Moses et Aaron iuxta sermonem Domini per manum Mosi
NUM|4|38|numerati sunt et filii Gerson per cognationes et domos patrum suorum
NUM|4|39|a triginta annis et supra usque ad annum quinquagesimum omnes qui ingrediuntur ut ministrent in tabernaculo foederis
NUM|4|40|et inventi sunt duo milia sescenti triginta
NUM|4|41|hic est populus Gersonitarum quos numeraverunt Moses et Aaron iuxta verbum Domini
NUM|4|42|numerati sunt et filii Merari per cognationes et domos patrum suorum
NUM|4|43|a triginta annis et supra usque ad annum quinquagesimum omnes qui ingrediuntur ad explendos ritus tabernaculi foederis
NUM|4|44|et inventi sunt tria milia ducenti
NUM|4|45|hic est numerus filiorum Merari quos recensuerunt Moses et Aaron iuxta imperium Domini per manum Mosi
NUM|4|46|omnes qui recensiti sunt de Levitis et quos fecit ad nomen Moses et Aaron et principes Israhel per cognationes et domos patrum suorum
NUM|4|47|a triginta annis et supra usque ad annum quinquagesimum ingredientes ad ministerium tabernaculi et onera portanda
NUM|4|48|fuerunt simul octo milia quingenti octoginta
NUM|4|49|iuxta verbum Domini recensuit eos Moses unumquemque iuxta officium et onera sua sicut praeceperat ei Dominus
NUM|5|1|locutusque est Dominus ad Mosen dicens
NUM|5|2|praecipe filiis Israhel ut eiciant de castris omnem leprosum et qui semine fluit pollutusque est super mortuo
NUM|5|3|tam masculum quam feminam eicite de castris ne contaminent ea cum habitaverim vobiscum
NUM|5|4|feceruntque ita filii Israhel et eiecerunt eos extra castra sicut locutus erat Dominus Mosi
NUM|5|5|locutus est Dominus ad Mosen dicens
NUM|5|6|loquere ad filios Israhel vir sive mulier cum fecerint ex omnibus peccatis quae solent hominibus accidere et per neglegentiam transgressi fuerint mandatum Domini atque deliquerint
NUM|5|7|confitebuntur peccatum suum et reddent ipsum caput quintamque partem desuper ei in quem peccaverint
NUM|5|8|sin autem non fuerit qui recipiat dabunt Domino et erit sacerdotis excepto ariete qui offertur pro expiatione ut sit placabilis hostia
NUM|5|9|omnes quoque primitiae quas offerunt filii Israhel ad sacerdotem pertinent
NUM|5|10|et quicquid in sanctuarium offertur a singulis et traditur manibus sacerdotis ipsius erit
NUM|5|11|locutus est Dominus ad Mosen dicens
NUM|5|12|loquere ad filios Israhel et dices ad eos vir cuius uxor erraverit maritumque contemnens
NUM|5|13|dormierit cum altero viro et hoc maritus deprehendere non quiverit sed latet adulterium et testibus argui non potest quia non est inventa in stupro
NUM|5|14|si spiritus zelotypiae concitaverit virum contra uxorem suam quae vel polluta est vel falsa suspicione appetitur
NUM|5|15|adducet eam ad sacerdotem et offeret oblationem pro illa decimam partem sati farinae hordiaciae non fundet super eam oleum nec inponet tus quia sacrificium zelotypiae est et oblatio investigans adulterium
NUM|5|16|offeret igitur eam sacerdos et statuet coram Domino
NUM|5|17|adsumetque aquam sanctam in vase fictili et pauxillum terrae de pavimento tabernaculi mittet in eam
NUM|5|18|cumque steterit mulier in conspectu Domini discoperiet caput eius et ponet super manus illius sacrificium recordationis et oblationem zelotypiae ipse autem tenebit aquas amarissimas in quibus cum execratione maledicta congessit
NUM|5|19|adiurabitque eam et dicet si non dormivit vir alienus tecum et si non polluta es deserto mariti toro non te nocebunt aquae istae amarissimae in quas maledicta congessi
NUM|5|20|sin autem declinasti a viro tuo atque polluta es et concubuisti cum altero
NUM|5|21|his maledictionibus subiacebis det te Dominus in maledictionem exemplumque cunctorum in populo suo putrescere faciat femur tuum et tumens uterus disrumpatur
NUM|5|22|ingrediantur aquae maledictae in ventrem tuum et utero tumescente putrescat femur et respondebit mulier amen amen
NUM|5|23|scribetque sacerdos in libello ista maledicta et delebit ea aquis amarissimis in quas maledicta congessit
NUM|5|24|et dabit ei bibere quas cum exhauserit
NUM|5|25|tollet sacerdos de manu eius sacrificium zelotypiae et elevabit illud coram Domino inponetque super altare ita dumtaxat ut prius
NUM|5|26|pugillum sacrificii tollat de eo quod offertur et incendat super altare et sic potum det mulieri aquas amarissimas
NUM|5|27|quas cum biberit si polluta est et contempto viro adulterii rea pertransibunt eam aquae maledictionis et inflato ventre conputrescet femur eritque mulier in maledictionem et in exemplum omni populo
NUM|5|28|quod si polluta non fuerit erit innoxia et faciet liberos
NUM|5|29|ista est lex zelotypiae si declinaverit mulier a viro suo et si polluta fuerit
NUM|5|30|maritusque zelotypiae spiritu concitatus adduxerit eam in conspectu Domini et fecerit ei sacerdos iuxta omnia quae scripta sunt
NUM|5|31|maritus absque culpa erit et illa recipiet iniquitatem suam
NUM|6|1|locutus est Dominus ad Mosen dicens
NUM|6|2|loquere ad filios Israhel et dices ad eos vir sive mulier cum fecerit votum ut sanctificentur et se voluerint Domino consecrare
NUM|6|3|vino et omni quod inebriare potest abstinebunt acetum ex vino et ex qualibet alia potione et quicquid de uva exprimitur non bibent uvas recentes siccasque non comedent
NUM|6|4|cunctis diebus quibus ex voto Domino consecrantur quicquid ex vinea esse potest ab uva passa usque ad acinum non comedent
NUM|6|5|omni tempore separationis suae novacula non transibit super caput eius usque ad conpletum diem quo Domino consecratur sanctus erit crescente caesarie capitis eius
NUM|6|6|omni tempore consecrationis suae super mortuum non ingredietur
NUM|6|7|nec super patris quidem et matris et fratris sororisque funere contaminabitur quia consecratio Dei sui super caput eius est
NUM|6|8|omnes dies separationis suae sanctus erit Domino
NUM|6|9|sin autem mortuus fuerit subito quispiam coram eo polluetur caput consecrationis eius quod radet ilico et in eadem die purgationis suae et rursum septima
NUM|6|10|in octavo autem die offeret duos turtures vel duos pullos columbae sacerdoti in introitu foederis testimonii
NUM|6|11|facietque sacerdos unum pro peccato et alterum in holocaustum et deprecabitur pro eo quia peccavit super mortuo sanctificabitque caput eius in die illo
NUM|6|12|et consecrabit Domino dies separationis illius offerens agnum anniculum pro peccato ita tamen ut dies priores irriti fiant quoniam polluta est sanctificatio eius
NUM|6|13|ista est lex consecrationis cum dies quos ex voto decreverat conplebuntur adducet eum ad ostium tabernaculi foederis
NUM|6|14|et offeret oblationem eius Domino agnum anniculum inmaculatum in holocaustum et ovem anniculam inmaculatam pro peccato et arietem inmaculatum hostiam pacificam
NUM|6|15|canistrum quoque panum azymorum qui conspersi sunt oleo et lagana absque fermento uncta oleo ac libamina singulorum
NUM|6|16|quae offeret sacerdos coram Domino et faciet tam pro peccato quam in holocaustum
NUM|6|17|arietem vero immolabit hostiam pacificam Domino offerens simul canistrum azymorum et libamenta quae ex more debentur
NUM|6|18|tunc radetur nazareus ante ostium tabernaculi foederis caesarie consecrationis suae tolletque capillos eius et ponet super ignem qui est subpositus sacrificio pacificorum
NUM|6|19|et armum coctum arietis tortamque absque fermento unam de canistro et laganum azymum unum et tradet in manibus nazarei postquam rasum fuerit caput eius
NUM|6|20|susceptaque rursum ab eo elevabit in conspectu Domini et sanctificata sacerdotis erunt sicut pectusculum quod separari iussum est et femur post haec potest bibere nazareus vinum
NUM|6|21|ista est lex nazarei cum voverit oblationem suam Domino tempore consecrationis suae exceptis his quae invenerit manus eius iuxta quod mente devoverat ita faciet ad perfectionem sanctificationis suae
NUM|6|22|locutus est Dominus ad Mosen dicens
NUM|6|23|loquere Aaron et filiis eius sic benedicetis filiis Israhel et dicetis eis
NUM|6|24|benedicat tibi Dominus et custodiat te
NUM|6|25|ostendat Dominus faciem suam tibi et misereatur tui
NUM|6|26|convertat Dominus vultum suum ad te et det tibi pacem
NUM|6|27|invocabunt nomen meum super filios Israhel et ego benedicam eis
NUM|7|1|factum est autem in die qua conplevit Moses tabernaculum et erexit illud unxitque et sanctificavit cum omnibus vasis suis altare similiter et vasa eius
NUM|7|2|obtulerunt principes Israhel et capita familiarum qui erant per singulas tribus praefecti eorum qui numerati fuerant
NUM|7|3|munera coram Domino sex plaustra tecta cum duodecim bubus unum plaustrum obtulere duo duces et unum bovem singuli obtuleruntque ea in conspectu tabernaculi
NUM|7|4|ait autem Dominus ad Mosen
NUM|7|5|suscipe ab eis ut serviant in ministerio tabernaculi et tradas ea Levitis iuxta ordinem ministerii sui
NUM|7|6|itaque cum suscepisset Moses plaustra et boves tradidit eos Levitis
NUM|7|7|duo plaustra et quattuor boves dedit filiis Gerson iuxta id quod habebant necessarium
NUM|7|8|quattuor alia plaustra et octo boves dedit filiis Merari secundum officia et cultum suum sub manu Ithamar filii Aaron sacerdotis
NUM|7|9|filiis autem Caath non dedit plaustra et boves quia in sanctuario serviunt et onera propriis portant umeris
NUM|7|10|igitur obtulerunt duces in dedicationem altaris die qua unctum est oblationem suam ante altare
NUM|7|11|dixitque Dominus ad Mosen singuli duces per singulos dies offerant munera in dedicationem altaris
NUM|7|12|primo die obtulit oblationem suam Naasson filius Aminadab de tribu Iuda
NUM|7|13|fueruntque in ea acetabulum argenteum pondo centum triginta siclorum fiala argentea habens septuaginta siclos iuxta pondus sanctuarii utrumque plenum simila conspersa oleo in sacrificium
NUM|7|14|mortariolum ex decem siclis aureis plenum incenso
NUM|7|15|bovem et arietem et agnum anniculum in holocaustum
NUM|7|16|hircumque pro peccato
NUM|7|17|et in sacrificio pacificorum boves duos arietes quinque hircos quinque agnos anniculos quinque haec est oblatio Naasson filii Aminadab
NUM|7|18|secundo die obtulit Nathanahel filius Suar dux de tribu Isachar
NUM|7|19|acetabulum argenteum adpendens centum triginta siclos fialam argenteam habentem septuaginta siclos iuxta pondus sanctuarii utrumque plenum simila conspersa oleo in sacrificium
NUM|7|20|mortariolum aureum habens decem siclos plenum incenso
NUM|7|21|bovem de armento et arietem et agnum anniculum in holocaustum
NUM|7|22|hircumque pro peccato
NUM|7|23|et in sacrificio pacificorum boves duos arietes quinque hircos quinque agnos anniculos quinque haec fuit oblatio Nathanahel filii Suar
NUM|7|24|tertio die princeps filiorum Zabulon Heliab filius Helon
NUM|7|25|obtulit acetabulum argenteum adpendens centum triginta siclos fialam argenteam habentem septuaginta siclos ad pondus sanctuarii utrumque plenum simila conspersa oleo in sacrificium
NUM|7|26|mortariolum aureum adpendens decem siclos plenum incenso
NUM|7|27|bovem de armento et arietem et agnum anniculum in holocaustum
NUM|7|28|hircumque pro peccato
NUM|7|29|et in sacrificio pacificorum boves duos arietes quinque hircos quinque agnos anniculos quinque haec est oblatio Heliab filii Helon
NUM|7|30|die quarto princeps filiorum Ruben Helisur filius Sedeur
NUM|7|31|obtulit acetabulum argenteum adpendens centum triginta siclos fialam argenteam habentem septuaginta siclos ad pondus sanctuarii utrumque plenum simila conspersa oleo in sacrificium
NUM|7|32|mortariolum aureum adpendens decem siclos plenum incenso
NUM|7|33|bovem de armento et arietem et agnum anniculum in holocaustum
NUM|7|34|hircumque pro peccato
NUM|7|35|et in hostias pacificorum boves duos arietes quinque hircos quinque agnos anniculos quinque haec fuit oblatio Helisur filii Sedeur
NUM|7|36|die quinto princeps filiorum Symeon Salamihel filius Surisaddai
NUM|7|37|obtulit acetabulum argenteum adpendens centum triginta siclos fialam argenteam habentem septuaginta siclos ad pondus sanctuarii utrumque plenum simila conspersa oleo in sacrificium
NUM|7|38|mortariolum aureum adpendens decem siclos plenum incenso
NUM|7|39|bovem de armento et arietem et agnum anniculum in holocaustum
NUM|7|40|hircumque pro peccato
NUM|7|41|et in hostias pacificorum boves duos arietes quinque hircos quinque agnos anniculos quinque haec fuit oblatio Salamihel filii Surisaddai
NUM|7|42|die sexto princeps filiorum Gad Heliasaph filius Duhel
NUM|7|43|obtulit acetabulum argenteum adpendens centum triginta siclos fialam argenteam habentem septuaginta siclos ad pondus sanctuarii utrumque plenum simila conspersa oleo in sacrificium
NUM|7|44|mortariolum aureum adpendens siclos decem plenum incenso
NUM|7|45|bovem de armento et arietem et agnum anniculum in holocaustum
NUM|7|46|hircumque pro peccato
NUM|7|47|et in hostias pacificorum boves duos arietes quinque hircos quinque agnos anniculos quinque haec fuit oblatio Heliasaph filii Duhel
NUM|7|48|die septimo princeps filiorum Ephraim Helisama filius Ammiud
NUM|7|49|obtulit acetabulum argenteum adpendens centum triginta siclos fialam argenteam habentem septuaginta siclos ad pondus sanctuarii utrumque plenum simila conspersa oleo in sacrificium
NUM|7|50|mortariolum aureum adpendens decem siclos plenum incenso
NUM|7|51|bovem de armento et arietem et agnum anniculum in holocaustum
NUM|7|52|hircumque pro peccato
NUM|7|53|et in hostias pacificas boves duos arietes quinque hircos quinque agnos anniculos quinque haec fuit oblatio Helisama filii Ammiud
NUM|7|54|die octavo princeps filiorum Manasse Gamalihel filius Phadassur
NUM|7|55|obtulit acetabulum argenteum adpendens centum triginta siclos fialam argenteam habentem septuaginta siclos ad pondus sanctuarii utrumque plenum simila conspersa oleo in sacrificium
NUM|7|56|mortariolum aureum adpendens decem siclos plenum incenso
NUM|7|57|bovem de armento et arietem et agnum anniculum in holocaustum
NUM|7|58|hircumque pro peccato
NUM|7|59|et in hostias pacificorum boves duos arietes quinque hircos quinque agnos anniculos quinque haec fuit oblatio Gamalihel filii Phadassur
NUM|7|60|die nono princeps filiorum Beniamin Abidan filius Gedeonis
NUM|7|61|obtulit acetabulum argenteum adpendens centum triginta siclos fialam argenteam habentem septuaginta siclos ad pondus sanctuarii utrumque plenum simila conspersa oleo in sacrificium
NUM|7|62|mortariolum aureum adpendens decem siclos plenum incenso
NUM|7|63|bovem de armento et arietem et agnum anniculum in holocaustum
NUM|7|64|hircumque pro peccato
NUM|7|65|et in hostias pacificorum boves duos arietes quinque hircos quinque agnos anniculos quinque haec fuit oblatio Abidan filii Gedeonis
NUM|7|66|die decimo princeps filiorum Dan Ahiezer filius Amisaddai
NUM|7|67|obtulit acetabulum argenteum adpendens centum triginta siclos fialam argenteam habentem septuaginta siclos ad pondus sanctuarii utrumque plenum simila conspersa oleo in sacrificium
NUM|7|68|mortariolum aureum adpendens decem siclos plenum incenso
NUM|7|69|bovem de armento et arietem et agnum anniculum in holocaustum
NUM|7|70|hircumque pro peccato
NUM|7|71|et in hostias pacificorum boves duos arietes quinque hircos quinque agnos anniculos quinque haec fuit oblatio Ahiezer filii Amisaddai
NUM|7|72|die undecimo princeps filiorum Aser Phagaihel filius Ochran
NUM|7|73|obtulit acetabulum argenteum adpendens centum triginta siclos fialam argenteam habentem septuaginta siclos ad pondus sanctuarii utrumque plenum simila conspersa oleo in sacrificium
NUM|7|74|mortariolum aureum adpendens decem siclos plenum incenso
NUM|7|75|bovem de armento et arietem et agnum anniculum in holocaustum
NUM|7|76|hircumque pro peccato
NUM|7|77|et in hostias pacificorum boves duos arietes quinque hircos quinque agnos anniculos quinque haec fuit oblatio Phagaihel filii Ochran
NUM|7|78|die duodecimo princeps filiorum Nepthalim Achira filius Henan
NUM|7|79|obtulit acetabulum argenteum adpendens centum triginta siclos fialam argenteam habentem septuaginta siclos ad pondus sanctuarii utrumque plenum simila conspersa oleo in sacrificium
NUM|7|80|mortariolum aureum adpendens decem siclos plenum incenso
NUM|7|81|bovem de armento et arietem et agnum anniculum in holocaustum
NUM|7|82|hircumque pro peccato
NUM|7|83|et in hostias pacificorum boves duos arietes quinque hircos quinque agnos anniculos quinque haec fuit oblatio Achira filii Henan
NUM|7|84|haec in dedicatione altaris oblata sunt a principibus Israhel in die qua consecratum est acetabula argentea duodecim fialae argenteae duodecim mortariola aurea duodecim
NUM|7|85|ita ut centum triginta argenti siclos haberet unum acetabulum et septuaginta siclos una fiala id est in commune vasorum omnium ex argento sicli duo milia quadringenti pondere sanctuarii
NUM|7|86|mortariola aurea duodecim plena incenso denos siclos adpendentia pondere sanctuarii id est simul auri sicli centum viginti
NUM|7|87|boves de armento in holocaustum duodecim arietes duodecim agni anniculi duodecim et libamenta eorum hirci duodecim pro peccato
NUM|7|88|hostiae pacificorum boves viginti quattuor arietes sexaginta hirci sexaginta agni anniculi sexaginta haec oblata sunt in dedicatione altaris quando unctum est
NUM|7|89|cumque ingrederetur Moses tabernaculum foederis ut consuleret oraculum audiebat vocem loquentis ad se de propitiatorio quod erat super arcam testimonii inter duos cherubin unde et loquebatur ei
NUM|8|1|locutus est Dominus ad Mosen dicens
NUM|8|2|loquere Aaroni et dices ad eum cum posueris septem lucernas contra eam partem quam candelabrum respicit lucere debebunt
NUM|8|3|fecitque Aaron et inposuit lucernas super candelabrum ut praeceperat Dominus Mosi
NUM|8|4|haec autem erat factura candelabri ex auro ductili tam medius stipes quam cuncta ex utroque calamorum latera nascebantur iuxta exemplum quod ostendit Dominus Mosi ita operatus est candelabrum
NUM|8|5|et locutus est Dominus ad Mosen dicens
NUM|8|6|tolle Levitas de medio filiorum Israhel et purificabis eos
NUM|8|7|iuxta hunc ritum aspergantur aqua lustrationis et radant omnes pilos carnis suae cumque laverint vestimenta sua et mundati fuerint
NUM|8|8|tollant bovem de armentis et libamentum eius similam oleo conspersam bovem autem alterum de armento tu accipies pro peccato
NUM|8|9|et adplicabis Levitas coram tabernaculo foederis convocata omni multitudine filiorum Israhel
NUM|8|10|cumque Levitae fuerint coram Domino ponent filii Israhel manus suas super eos
NUM|8|11|et offeret Aaron Levitas munus in conspectu Domini a filiis Israhel ut serviant in ministerio eius
NUM|8|12|Levitae quoque ponent manus suas super capita boum e quibus unum facies pro peccato et alterum in holocaustum Domini ut depreceris pro eis
NUM|8|13|statuesque Levitas in conspectu Aaron et filiorum eius et consecrabis oblatos Domino
NUM|8|14|ac separabis de medio filiorum Israhel ut sint mei
NUM|8|15|et postea ingrediantur tabernaculum foederis ut serviant mihi sicque purificabis et consecrabis eos in oblationem Domini quoniam dono donati sunt mihi a filiis Israhel
NUM|8|16|pro primogenitis quae aperiunt omnem vulvam in Israhel accepi eos
NUM|8|17|mea sunt omnia primogenita filiorum Israhel tam ex hominibus quam ex iumentis ex die quo percussi omnem primogenitum in terra Aegypti sanctificavi eos mihi
NUM|8|18|et tuli Levitas pro cunctis primogenitis filiorum Israhel
NUM|8|19|tradidique eos dono Aaroni et filiis eius de medio populi ut serviant mihi pro Israhel in tabernaculo foederis et orent pro eis ne sit in populo plaga si ausi fuerint accedere ad sanctuarium
NUM|8|20|feceruntque Moses et Aaron et omnis multitudo filiorum Israhel super Levitas quae praeceperat Dominus Mosi
NUM|8|21|purificatique sunt et laverunt vestimenta sua elevavitque eos Aaron in conspectu Domini et oravit pro eis
NUM|8|22|ut purificati ingrederentur ad officia sua in tabernaculum foederis coram Aaron et filiis eius sicut praeceperat Dominus Mosi de Levitis ita factum est
NUM|8|23|locutus est Dominus ad Mosen dicens
NUM|8|24|haec est lex Levitarum a viginti quinque annis et supra ingredientur ut ministrent in tabernaculo foederis
NUM|8|25|cumque quinquagesimum annum aetatis impleverint servire cessabunt
NUM|8|26|eruntque ministri fratrum suorum in tabernaculo foederis ut custodiant quae sibi fuerint commendata opera autem ipsa non faciant sic dispones Levitas in custodiis suis
NUM|9|1|locutus est Dominus ad Mosen in deserto Sinai anno secundo postquam egressi sunt de terra Aegypti mense primo dicens
NUM|9|2|faciant filii Israhel phase in tempore suo
NUM|9|3|quartadecima die mensis huius ad vesperam iuxta omnes caerimonias et iustificationes eius
NUM|9|4|praecepitque Moses filiis Israhel ut facerent phase
NUM|9|5|qui fecerunt tempore suo quartadecima die mensis ad vesperam in monte Sinai iuxta omnia quae mandaverat Dominus Mosi fecerunt filii Israhel
NUM|9|6|ecce autem quidam inmundi super animam hominis qui non poterant facere pascha in die illo accedentes ad Mosen et Aaron
NUM|9|7|dixerunt eis inmundi sumus super animam hominis quare fraudamur ut non valeamus offerre oblationem Domino in tempore suo inter filios Israhel
NUM|9|8|quibus respondit Moses state ut consulam quid praecipiat Dominus de vobis
NUM|9|9|locutusque est Dominus ad Mosen dicens
NUM|9|10|loquere filiis Israhel homo qui fuerit inmundus super anima sive in via procul in gente vestra faciat phase Domino
NUM|9|11|mense secundo quartadecima die mensis ad vesperam cum azymis et lactucis agrestibus comedent illud
NUM|9|12|non relinquent ex eo quippiam usque mane et os eius non confringent omnem ritum phase observabunt
NUM|9|13|si quis autem et mundus est et in itinere non fuit et tamen non fecit phase exterminabitur anima illa de populis suis quia sacrificium Domino non obtulit tempore suo peccatum suum ipse portabit
NUM|9|14|peregrinus quoque et advena si fuerit apud vos faciet phase Domini iuxta caerimonias et iustificationes eius praeceptum idem erit apud vos tam advenae quam indigenae
NUM|9|15|igitur die qua erectum est tabernaculum operuit illud nubes a vespere autem super tentorium erat quasi species ignis usque mane
NUM|9|16|sic fiebat iugiter per diem operiebat illud nubes et per noctem quasi species ignis
NUM|9|17|cumque ablata fuisset nubes quae tabernaculum protegebat tunc proficiscebantur filii Israhel et in loco ubi stetisset nubes ibi castrametabantur
NUM|9|18|ad imperium Domini proficiscebantur et ad imperium illius figebant tabernaculum cunctis diebus quibus stabat nubes super tabernaculum manebant in eodem loco
NUM|9|19|et si evenisset ut multo tempore maneret super illud erant filii Israhel in excubiis Domini et non proficiscebantur
NUM|9|20|quotquot diebus fuisset nubes super tabernaculum ad imperium Domini erigebant tentoria et ad imperium illius deponebant
NUM|9|21|si fuisset nubes a vespere usque mane et statim diluculo tabernaculum reliquisset proficiscebantur et si post diem et noctem recessisset dissipabant tentoria
NUM|9|22|si biduo aut uno mense vel longiori tempore fuisset super tabernaculum manebant filii Israhel in eodem loco et non proficiscebantur statim autem ut recessisset movebant castra
NUM|9|23|per verbum Domini figebant tentoria et per verbum illius proficiscebantur erantque in excubiis Domini iuxta imperium eius per manum Mosi
NUM|10|1|locutus est Dominus ad Mosen dicens
NUM|10|2|fac tibi duas tubas argenteas ductiles quibus convocare possis multitudinem quando movenda sunt castra
NUM|10|3|cumque increpueris tubis congregabitur ad te omnis turba ad ostium foederis tabernaculi
NUM|10|4|si semel clangueris venient ad te principes et capita multitudinis Israhel
NUM|10|5|sin autem prolixior atque concisus clangor increpuerit movebunt castra primi qui sunt ad orientalem plagam
NUM|10|6|in secundo autem sonitu et pari ululatu tubae levabunt tentoria qui habitant ad meridiem et iuxta hunc modum reliqui facient ululantibus tubis in profectione
NUM|10|7|quando autem congregandus est populus simplex tubarum clangor erit et non concise ululabunt
NUM|10|8|filii Aaron sacerdotes clangent tubis eritque hoc legitimum sempiternum in generationibus vestris
NUM|10|9|si exieritis ad bellum de terra vestra contra hostes qui dimicant adversum vos clangetis ululantibus tubis et erit recordatio vestri coram Domino Deo vestro ut eruamini de manibus inimicorum vestrorum
NUM|10|10|si quando habebitis epulum et dies festos et kalendas canetis tubis super holocaustis et pacificis victimis ut sint vobis in recordationem Dei vestri ego Dominus Deus vester
NUM|10|11|anno secundo mense secundo vicesima die mensis elevata est nubes de tabernaculo foederis
NUM|10|12|profectique sunt filii Israhel per turmas suas de deserto Sinai et recubuit nubes in solitudine Pharan
NUM|10|13|moveruntque castra primi iuxta imperium Domini in manu Mosi
NUM|10|14|filii Iuda per turmas suas quorum princeps erat Naasson filius Aminadab
NUM|10|15|in tribu filiorum Isachar fuit princeps Nathanahel filius Suar
NUM|10|16|in tribu Zabulon erat princeps Heliab filius Helon
NUM|10|17|depositumque est tabernaculum quod portantes egressi sunt filii Gerson et Merari
NUM|10|18|profectique sunt et filii Ruben per turmas et ordinem suum quorum princeps erat Helisur filius Sedeur
NUM|10|19|in tribu autem filiorum Symeon princeps fuit Salamihel filius Surisaddai
NUM|10|20|porro in tribu Gad erat princeps Heliasaph filius Duhel
NUM|10|21|profectique sunt et Caathitae portantes sanctuarium tamdiu tabernaculum portabatur donec venirent ad erectionis locum
NUM|10|22|moverunt castra et filii Ephraim per turmas suas in quorum exercitu princeps erat Helisama filius Ammiud
NUM|10|23|in tribu autem filiorum Manasse princeps fuit Gamalihel filius Phadassur
NUM|10|24|et in tribu Beniamin dux Abidan filius Gedeonis
NUM|10|25|novissimi castrorum omnium profecti sunt filii Dan per turmas suas in quorum exercitu princeps fuit Ahiezer filius Amisaddai
NUM|10|26|in tribu autem filiorum Aser erat princeps Phagaihel filius Ochran
NUM|10|27|et in tribu filiorum Nepthalim princeps Achira filius Henan
NUM|10|28|haec sunt castra et profectiones filiorum Israhel per turmas suas quando egrediebantur
NUM|10|29|dixitque Moses Hobab filio Rahuhel Madianiti cognato suo proficiscimur ad locum quem Dominus daturus est nobis veni nobiscum ut benefaciamus tibi quia Dominus bona promisit Israheli
NUM|10|30|cui ille respondit non vadam tecum sed revertar in terram meam in qua natus sum
NUM|10|31|et ille noli inquit nos relinquere tu enim nosti in quibus locis per desertum castra ponere debeamus et eris ductor noster
NUM|10|32|cumque nobiscum veneris quicquid optimum fuerit ex opibus quas nobis traditurus est Dominus dabimus tibi
NUM|10|33|profecti sunt ergo de monte Domini via trium dierum arcaque foederis Domini praecedebat eos per dies tres providens castrorum locum
NUM|10|34|nubes quoque Domini super eos erat per diem cum incederent
NUM|10|35|cumque elevaretur arca dicebat Moses surge Domine et dissipentur inimici tui et fugiant qui oderunt te a facie tua
NUM|10|36|cum autem deponeretur aiebat revertere Domine ad multitudinem exercitus Israhel
NUM|11|1|interea ortum est murmur populi quasi dolentium pro labore contra Dominum quod cum audisset iratus est et accensus in eos ignis Domini devoravit extremam castrorum partem
NUM|11|2|cumque clamasset populus ad Mosen oravit Moses Dominum et absortus est ignis
NUM|11|3|vocavitque nomen loci illius Incensio eo quod succensus fuisset contra eos ignis Domini
NUM|11|4|vulgus quippe promiscuum quod ascenderat cum eis flagravit desiderio sedens et flens iunctis sibi pariter filiis Israhel et ait quis dabit nobis ad vescendum carnes
NUM|11|5|recordamur piscium quos comedebamus in Aegypto gratis in mentem nobis veniunt cucumeres et pepones porrique et cepae et alia
NUM|11|6|anima nostra arida est nihil aliud respiciunt oculi nostri nisi man
NUM|11|7|erat autem man quasi semen coriandri coloris bdellii
NUM|11|8|circuibatque populus et colligens illud frangebat mola sive terebat in mortario coquens in olla et faciens ex eo tortulas saporis quasi panis oleati
NUM|11|9|cumque descenderet nocte super castra ros descendebat pariter et man
NUM|11|10|audivit ergo Moses flentem populum per familias singulos per ostia tentorii sui iratusque est furor Domini valde sed et Mosi intoleranda res visa est
NUM|11|11|et ait ad Dominum cur adflixisti servum tuum quare non invenio gratiam coram te et cur inposuisti pondus universi populi huius super me
NUM|11|12|numquid ego concepi omnem hanc multitudinem vel genui eam ut dicas mihi porta eos in sinu tuo sicut portare solet nutrix infantulum et defer in terram pro qua iurasti patribus eorum
NUM|11|13|unde mihi carnes ut dem tantae multitudini flent contra me dicentes da nobis carnes ut comedamus
NUM|11|14|non possum solus sustinere omnem hunc populum quia gravis mihi est
NUM|11|15|sin aliter tibi videtur obsecro ut interficias me et inveniam gratiam in oculis tuis ne tantis adficiar malis
NUM|11|16|et dixit Dominus ad Mosen congrega mihi septuaginta viros de senibus Israhel quos tu nosti quod senes populi sint ac magistri et duces eos ad ostium tabernaculi foederis faciesque ibi stare tecum
NUM|11|17|ut descendam et loquar tibi et auferam de spiritu tuo tradamque eis ut sustentent tecum onus populi et non tu solus graveris
NUM|11|18|populo quoque dices sanctificamini cras comedetis carnes ego enim audivi vos dicere quis dabit nobis escas carnium bene nobis erat in Aegypto ut det vobis Dominus carnes et comedatis
NUM|11|19|non uno die nec duobus vel quinque aut decem nec viginti quidem
NUM|11|20|sed usque ad mensem dierum donec exeat per nares vestras et vertatur in nausiam eo quod reppuleritis Dominum qui in medio vestri est et fleveritis coram eo dicentes quare egressi sumus ex Aegypto
NUM|11|21|et ait Moses sescenta milia peditum huius populi sunt et tu dicis dabo eis esum carnium mense integro
NUM|11|22|numquid ovium et boum multitudo caedetur ut possit sufficere ad cibum vel omnes pisces maris in unum congregabuntur ut eos satient
NUM|11|23|cui respondit Dominus numquid manus Domini invalida est iam nunc videbis utrum meus sermo opere conpleatur
NUM|11|24|venit igitur Moses et narravit populo verba Domini congregans septuaginta viros de senibus Israhel quos stare fecit circa tabernaculum
NUM|11|25|descenditque Dominus per nubem et locutus est ad eum auferens de spiritu qui erat in Mosen et dans septuaginta viris cumque requievisset in eis spiritus prophetaverunt nec ultra cessarunt
NUM|11|26|remanserant autem in castris duo viri quorum unus vocabatur Heldad et alter Medad super quos requievit spiritus nam et ipsi descripti fuerant et non exierant ad tabernaculum
NUM|11|27|cumque prophetarent in castris cucurrit puer et nuntiavit Mosi dicens Heldad et Medad prophetant in castris
NUM|11|28|statim Iosue filius Nun minister Mosi et electus e pluribus ait domine mi Moses prohibe eos
NUM|11|29|at ille quid inquit aemularis pro me quis tribuat ut omnis populus prophetet et det eis Dominus spiritum suum
NUM|11|30|reversusque est Moses et maiores natu Israhel in castra
NUM|11|31|ventus autem egrediens a Domino arreptas trans mare coturnices detulit et dimisit in castra itinere quantum uno die confici potest ex omni parte castrorum per circuitum volabantque in aere duobus cubitis altitudine super terram
NUM|11|32|surgens ergo populus toto die illo et nocte ac die altero congregavit coturnicum qui parum decem choros et siccaverunt eas per gyrum castrorum
NUM|11|33|adhuc carnes erant in dentibus eorum nec defecerat huiuscemodi cibus et ecce furor Domini concitatus in populum percussit eum plaga magna nimis
NUM|11|34|vocatusque est ille locus sepulchra Concupiscentiae ibi enim sepelierunt populum qui desideraverat egressi autem de sepulchris Concupiscentiae venerunt in Aseroth et manserunt ibi
NUM|11|35|
NUM|12|1|locutaque est Maria et Aaron contra Mosen propter uxorem eius aethiopissam
NUM|12|2|et dixerunt num per solum Mosen locutus est Dominus nonne et nobis similiter est locutus quod cum audisset Dominus
NUM|12|3|erat enim Moses vir mitissimus super omnes homines qui morabantur in terra
NUM|12|4|statim locutus est ad eum et ad Aaron et Mariam egredimini vos tantum tres ad tabernaculum foederis cumque fuissent egressi
NUM|12|5|descendit Dominus in columna nubis et stetit in introitu tabernaculi vocans Aaron et Mariam qui cum issent
NUM|12|6|dixit ad eos audite sermones meos si quis fuerit inter vos propheta Domini in visione apparebo ei vel per somnium loquar ad illum
NUM|12|7|at non talis servus meus Moses qui in omni domo mea fidelissimus est
NUM|12|8|ore enim ad os loquor ei et palam non per enigmata et figuras Dominum videt quare igitur non timuistis detrahere servo meo Mosi
NUM|12|9|iratusque contra eos abiit
NUM|12|10|nubes quoque recessit quae erat super tabernaculum et ecce Maria apparuit candens lepra quasi nix cumque respexisset eam Aaron et vidisset perfusam lepra
NUM|12|11|ait ad Mosen obsecro domine mi ne inponas nobis hoc peccatum quod stulte commisimus
NUM|12|12|ne fiat haec quasi mortua et ut abortivum quod proicitur de vulva matris suae ecce iam medium carnis eius devoratum est lepra
NUM|12|13|clamavitque Moses ad Dominum dicens Deus obsecro sana eam
NUM|12|14|cui respondit Dominus si pater eius spuisset in faciem illius nonne debuerat saltem septem dierum rubore suffundi separetur septem diebus extra castra et postea revocabitur
NUM|12|15|exclusa est itaque Maria extra castra septem diebus et populus non est motus de loco illo donec revocata est Maria
NUM|12|16|
NUM|13|1|profectus est de Aseroth fixis tentoriis in deserto Pharan
NUM|13|2|ibi locutus est Dominus ad Mosen dicens
NUM|13|3|mitte viros qui considerent terram Chanaan quam daturus sum filiis Israhel singulos de singulis tribubus ex principibus
NUM|13|4|fecit Moses quod Dominus imperarat de deserto Pharan mittens principes viros quorum ista sunt nomina
NUM|13|5|de tribu Ruben Semmua filium Zecchur
NUM|13|6|de tribu Symeon Saphat filium Huri
NUM|13|7|de tribu Iuda Chaleb filium Iepphonne
NUM|13|8|de tribu Isachar Igal filium Ioseph
NUM|13|9|de tribu Ephraim Osee filium Nun
NUM|13|10|de tribu Beniamin Phalti filium Raphu
NUM|13|11|de tribu Zabulon Geddihel filium Sodi
NUM|13|12|de tribu Ioseph sceptri Manasse Gaddi filium Susi
NUM|13|13|de tribu Dan Ammihel filium Gemalli
NUM|13|14|de tribu Aser Sthur filium Michahel
NUM|13|15|de tribu Nepthali Naabbi filium Vaphsi
NUM|13|16|de tribu Gad Guhel filium Machi
NUM|13|17|haec sunt nomina virorum quos misit Moses ad considerandam terram vocavitque Osee filium Nun Iosue
NUM|13|18|misit ergo eos Moses ad considerandam terram Chanaan et dixit ad eos ascendite per meridianam plagam cumque veneritis ad montes
NUM|13|19|considerate terram qualis sit et populum qui habitator est eius utrum fortis sit an infirmus pauci numero an plures
NUM|13|20|ipsa terra bona an mala urbes quales muratae an absque muris
NUM|13|21|humus pinguis an sterilis nemorosa an absque arboribus confortamini et adferte nobis de fructibus terrae erat autem tempus quando iam praecoquae uvae vesci possunt
NUM|13|22|cumque ascendissent exploraverunt terram a deserto Sin usque Roob intrantibus Emath
NUM|13|23|ascenderuntque ad meridiem et venerunt in Hebron ubi erant Ahiman et Sisai et Tholmai filii Enach nam Hebron septem annis ante Tanim urbem Aegypti condita est
NUM|13|24|pergentesque usque ad torrentem Botri absciderunt palmitem cum uva sua quem portaverunt in vecte duo viri de malis quoque granatis et de ficis loci illius tulerunt
NUM|13|25|qui appellatus est Neelescol id est torrens Botri eo quod botrum inde portassent filii Israhel
NUM|13|26|reversique exploratores terrae post quadraginta dies omni regione circuita
NUM|13|27|venerunt ad Mosen et Aaron et ad omnem coetum filiorum Israhel in desertum Pharan quod est in Cades locutique eis et omni multitudini ostenderunt fructus terrae
NUM|13|28|et narraverunt dicentes venimus in terram ad quam misisti nos quae re vera fluit lacte et melle ut ex his fructibus cognosci potest
NUM|13|29|sed cultores fortissimos habet et urbes grandes atque muratas stirpem Enach vidimus ibi
NUM|13|30|Amalech habitat in meridie Hettheus et Iebuseus et Amorreus in montanis Chananeus vero moratur iuxta mare et circa fluenta Iordanis
NUM|13|31|inter haec Chaleb conpescens murmur populi qui oriebatur contra Mosen ait ascendamus et possideamus terram quoniam poterimus obtinere eam
NUM|13|32|alii vero qui fuerant cum eo dicebant nequaquam ad hunc populum valemus ascendere quia fortior nobis est
NUM|13|33|detraxeruntque terrae quam inspexerant apud filios Israhel dicentes terram quam lustravimus devorat habitatores suos populum quem aspeximus procerae staturae est
NUM|13|34|ibi vidimus monstra quaedam filiorum Enach de genere giganteo quibus conparati quasi lucustae videbamur
NUM|14|1|igitur vociferans omnis turba flevit nocte illa
NUM|14|2|et murmurati sunt contra Mosen et Aaron cuncti filii Israhel dicentes
NUM|14|3|utinam mortui essemus in Aegypto et non in hac vasta solitudine utinam pereamus et non inducat nos Dominus in terram istam ne cadamus gladio et uxores ac liberi nostri ducantur captivi nonne melius est reverti in Aegyptum
NUM|14|4|dixeruntque alter ad alterum constituamus nobis ducem et revertamur in Aegyptum
NUM|14|5|quo audito Moses et Aaron ceciderunt proni in terram coram omni multitudine filiorum Israhel
NUM|14|6|at vero Iosue filius Nun et Chaleb filius Iepphonne qui et ipsi lustraverant terram sciderunt vestimenta sua
NUM|14|7|et ad omnem multitudinem filiorum Israhel locuti sunt terram quam circuivimus valde bona est
NUM|14|8|si propitius fuerit Dominus inducet nos in eam et tradet humum lacte et melle manantem
NUM|14|9|nolite rebelles esse contra Dominum neque timeatis populum terrae huius quia sicut panem ita eos possumus devorare recessit ab illis omne praesidium Dominus nobiscum est nolite metuere
NUM|14|10|cumque clamaret omnis multitudo et lapidibus eos vellet opprimere apparuit gloria Domini super tectum foederis cunctis filiis Israhel
NUM|14|11|et dixit Dominus ad Mosen usquequo detrahet mihi populus iste quousque non credent mihi in omnibus signis quae feci coram eis
NUM|14|12|feriam igitur eos pestilentia atque consumam te autem faciam principem super gentem magnam et fortiorem quam haec est
NUM|14|13|et ait Moses ad Dominum ut audiant Aegyptii de quorum medio eduxisti populum istum
NUM|14|14|et habitatores terrae huius qui audierunt quod tu Domine in populo isto sis et facie videaris ad faciem et nubes tua protegat illos et in columna nubis praecedas eos per diem et in columna ignis per noctem
NUM|14|15|quod occideris tantam multitudinem quasi unum hominem et dicant
NUM|14|16|non poterat introducere populum in terram pro qua iuraverat idcirco occidit eos in solitudine
NUM|14|17|magnificetur ergo fortitudo Domini sicut iurasti dicens
NUM|14|18|Dominus patiens et multae misericordiae auferens iniquitatem et scelera nullumque innoxium derelinquens qui visitas peccata patrum in filios in tertiam et quartam generationem
NUM|14|19|dimitte obsecro peccatum populi tui huius secundum magnitudinem misericordiae tuae sicut propitius fuisti egredientibus de Aegypto usque ad locum istum
NUM|14|20|dixitque Dominus dimisi iuxta verbum tuum
NUM|14|21|vivo ego et implebitur gloria Domini universa terra
NUM|14|22|attamen omnes homines qui viderunt maiestatem meam et signa quae feci in Aegypto et in solitudine et temptaverunt me iam per decem vices nec oboedierunt voci meae
NUM|14|23|non videbunt terram pro qua iuravi patribus eorum nec quisquam ex illis qui detraxit mihi intuebitur eam
NUM|14|24|servum meum Chaleb qui plenus alio spiritu secutus est me inducam in terram hanc quam circuivit et semen eius possidebit eam
NUM|14|25|quoniam Amalechites et Chananeus habitant in vallibus cras movete castra et revertimini in solitudinem per viam maris Rubri
NUM|14|26|locutusque est Dominus ad Mosen et Aaron dicens
NUM|14|27|usquequo multitudo haec pessima murmurat contra me querellas filiorum Israhel audivi
NUM|14|28|dic ergo eis vivo ego ait Dominus sicut locuti estis audiente me sic faciam vobis
NUM|14|29|in solitudine hac iacebunt cadavera vestra omnes qui numerati estis a viginti annis et supra et murmurastis contra me
NUM|14|30|non intrabitis terram super quam levavi manum meam ut habitare vos facerem praeter Chaleb filium Iepphonne et Iosue filium Nun
NUM|14|31|parvulos autem vestros de quibus dixistis quod praedae hostibus forent introducam ut videant terram quae vobis displicuit
NUM|14|32|vestra cadavera iacebunt in solitudine
NUM|14|33|filii vestri erunt vagi in deserto annis quadraginta et portabunt fornicationem vestram donec consumantur cadavera patrum in deserto
NUM|14|34|iuxta numerum quadraginta dierum quibus considerastis terram annus pro die inputabitur et quadraginta annis recipietis iniquitates vestras et scietis ultionem meam
NUM|14|35|quoniam sicut locutus sum ita faciam omni multitudini huic pessimae quae consurrexit adversum me in solitudine hac deficiet et morietur
NUM|14|36|igitur omnes viri quos miserat Moses ad contemplandam terram et qui reversi murmurare fecerant contra eum omnem multitudinem detrahentes terrae quod esset mala
NUM|14|37|mortui sunt atque percussi in conspectu Domini
NUM|14|38|Iosue autem filius Nun et Chaleb filius Iepphonne vixerunt ex omnibus qui perrexerant ad considerandam terram
NUM|14|39|locutusque est Moses universa verba haec ad omnes filios Israhel et luxit populus nimis
NUM|14|40|et ecce mane primo surgentes ascenderunt verticem montis atque dixerunt parati sumus ascendere ad locum de quo Dominus locutus est quia peccavimus
NUM|14|41|quibus Moses cur inquit transgredimini verbum Domini quod vobis non cedet in prosperum
NUM|14|42|nolite ascendere non enim est Dominus vobiscum ne corruatis coram inimicis vestris
NUM|14|43|Amalechites et Chananeus ante vos sunt quorum gladio corruetis eo quod nolueritis adquiescere Domino nec erit Dominus vobiscum
NUM|14|44|at illi contenebrati ascenderunt in verticem montis arca autem testamenti Domini et Moses non recesserunt de castris
NUM|14|45|descenditque Amalechites et Chananeus qui habitabant in monte et percutiens eos atque concidens persecutus est usque Horma
NUM|15|1|locutus est Dominus ad Mosen dicens
NUM|15|2|loquere ad filios Israhel et dices ad eos cum ingressi fueritis terram habitationis vestrae quam ego dabo vobis
NUM|15|3|et feceritis oblationem Domino in holocaustum aut victimam vota solventes vel sponte offerentes munera aut in sollemnitatibus vestris adolentes odorem suavitatis Domino de bubus sive de ovibus
NUM|15|4|offeret quicumque immolaverit victimam sacrificium similae decimam partem oephi conspersae oleo quod mensuram habebit quartam partem hin
NUM|15|5|et vinum ad liba fundenda eiusdem mensurae dabit in holocausto sive in victima per agnos singulos
NUM|15|6|et arietis erit sacrificium similae duarum decimarum quae conspersa sit oleo tertiae partis hin
NUM|15|7|et vinum ad libamentum tertiae partis eiusdem mensurae offeret in odorem suavitatis Domino
NUM|15|8|quando vero de bubus feceris holocaustum aut hostiam ut impleas votum vel pacificas victimas
NUM|15|9|dabis per singulos boves similae tres decimas conspersae oleo quod habeat medium mensurae hin
NUM|15|10|et vinum ad liba fundenda eiusdem mensurae in oblationem suavissimi odoris Domino
NUM|15|11|sic facietis
NUM|15|12|per singulos boves et arietes et agnos et hedos
NUM|15|13|tam indigenae quam peregrini
NUM|15|14|eodem ritu offerent sacrificia
NUM|15|15|unum praeceptum erit atque iudicium tam vobis quam advenis terrae
NUM|15|16|locutus est Dominus ad Mosen dicens
NUM|15|17|loquere filiis Israhel et dices ad eos
NUM|15|18|cum veneritis in terram quam dabo vobis
NUM|15|19|et comederitis de panibus regionis illius separabitis primitias Domino
NUM|15|20|de cibis vestris sicut de areis primitias separatis
NUM|15|21|ita et de pulmentis dabitis primitiva Domino
NUM|15|22|quod si per ignorantiam praeterieritis quicquam horum quae locutus est Dominus ad Mosen
NUM|15|23|et mandavit per eum ad vos a die qua coepit iubere et ultra
NUM|15|24|oblitaque fuerit facere multitudo offeret vitulum de armento holocaustum in odorem suavissimum Domino et sacrificium eius ac liba ut caerimoniae postulant hircumque pro peccato
NUM|15|25|et rogabit sacerdos pro omni multitudine filiorum Israhel et dimittetur eis quoniam non sponte peccaverunt nihilominus offerentes incensum Domino pro se et pro peccato atque errore suo
NUM|15|26|et dimittetur universae plebi filiorum Israhel et advenis qui peregrinantur inter vos quoniam culpa est omnis populi per ignorantiam
NUM|15|27|quod si anima una nesciens peccaverit offeret capram anniculam pro peccato suo
NUM|15|28|et deprecabitur pro ea sacerdos quod inscia peccaverit coram Domino inpetrabitque ei veniam et dimittetur illi
NUM|15|29|tam indigenis quam advenis una lex erit omnium qui peccaverint ignorantes
NUM|15|30|anima vero quae per superbiam aliquid commiserit sive civis sit ille sive peregrinus quoniam adversum Dominum rebellis fuit peribit de populo suo
NUM|15|31|verbum enim Domini contempsit et praeceptum illius fecit irritum idcirco delebitur et portabit iniquitatem suam
NUM|15|32|factum est autem cum essent filii Israhel in solitudine et invenissent hominem colligentem ligna in die sabbati
NUM|15|33|obtulerunt eum Mosi et Aaron et universae multitudini
NUM|15|34|qui recluserunt eum in carcerem nescientes quid super eo facere deberent
NUM|15|35|dixitque Dominus ad Mosen morte moriatur homo iste obruat eum lapidibus omnis turba extra castra
NUM|15|36|cumque eduxissent eum foras obruerunt lapidibus et mortuus est sicut praeceperat Dominus
NUM|15|37|dixit quoque Dominus ad Mosen
NUM|15|38|loquere filiis Israhel et dices ad eos ut faciant sibi fimbrias per angulos palliorum ponentes in eis vittas hyacinthinas
NUM|15|39|quas cum viderint recordentur omnium mandatorum Domini nec sequantur cogitationes suas et oculos per res varias fornicantes
NUM|15|40|sed magis memores praeceptorum Domini faciant ea sintque sancti Deo suo
NUM|15|41|ego Dominus Deus vester qui eduxi vos de terra Aegypti ut essem vester Deus
NUM|16|1|ecce autem Core filius Isaar filii Caath filii Levi et Dathan atque Abiram filii Heliab Hon quoque filius Pheleth de filiis Ruben
NUM|16|2|surrexerunt contra Mosen aliique filiorum Israhel ducenti quinquaginta viri proceres synagogae et qui tempore concilii per nomina vocabantur
NUM|16|3|cumque stetissent adversum Mosen et Aaron dixerunt sufficiat vobis quia omnis multitudo sanctorum est et in ipsis est Dominus cur elevamini super populum Domini
NUM|16|4|quod cum audisset Moses cecidit pronus in faciem
NUM|16|5|locutusque ad Core et ad omnem multitudinem mane inquit notum faciet Dominus qui ad se pertineant et sanctos adplicabit sibi et quos elegerit adpropinquabunt ei
NUM|16|6|hoc igitur facite tollat unusquisque turibula sua tu Core et omne concilium tuum
NUM|16|7|et hausto cras igne ponite desuper thymiama coram Domino et quemcumque elegerit ipse erit sanctus multum erigimini filii Levi
NUM|16|8|dixitque rursum ad Core audite filii Levi
NUM|16|9|num parum vobis est quod separavit vos Deus Israhel ab omni populo et iunxit sibi ut serviretis ei in cultu tabernaculi et staretis coram frequentia populi et ministraretis ei
NUM|16|10|idcirco ad se fecit accedere te et omnes fratres tuos filios Levi ut vobis etiam sacerdotium vindicetis
NUM|16|11|et omnis globus tuus stet contra Dominum quid est enim Aaron ut murmuretis contra eum
NUM|16|12|misit ergo Moses ut vocaret Dathan et Abiram filios Heliab qui responderunt non venimus
NUM|16|13|numquid parum est tibi quod eduxisti nos de terra quae lacte et melle manabat ut occideres in deserto nisi et dominatus fueris nostri
NUM|16|14|re vera induxisti nos in terram quae fluit rivis lactis et mellis et dedisti nobis possessiones agrorum et vinearum an et oculos nostros vis eruere non venimus
NUM|16|15|iratusque Moses valde ait ad Dominum ne respicias sacrificia eorum tu scis quod ne asellum quidem umquam acceperim ab eis nec adflixerim quempiam eorum
NUM|16|16|dixitque ad Core tu et omnis congregatio tua state seorsum coram Domino et Aaron die crastino separatim
NUM|16|17|tollite singuli turibula vestra et ponite super ea incensum offerentes Domino ducenta quinquaginta turibula Aaron quoque teneat turibulum suum
NUM|16|18|quod cum fecissent stantibus Mosen et Aaron
NUM|16|19|et coacervassent adversum eos omnem multitudinem ad ostium tabernaculi apparuit cunctis gloria Domini
NUM|16|20|locutusque Dominus ad Mosen et Aaron ait
NUM|16|21|separamini de medio congregationis huius ut eos repente disperdam
NUM|16|22|qui ceciderunt proni in faciem atque dixerunt fortissime Deus spirituum universae carnis num uno peccante contra omnes tua ira desaeviet
NUM|16|23|et ait Dominus ad Mosen
NUM|16|24|praecipe universo populo ut separetur a tabernaculis Core et Dathan et Abiram
NUM|16|25|surrexitque Moses et abiit ad Dathan et Abiram et sequentibus eum senioribus Israhel
NUM|16|26|dixit ad turbam recedite a tabernaculis hominum impiorum et nolite tangere quae ad eos pertinent ne involvamini in peccatis eorum
NUM|16|27|cumque recessissent a tentoriis eorum per circuitum Dathan et Abiram egressi stabant in introitu papilionum suorum cum uxoribus et liberis omnique frequentia
NUM|16|28|et ait Moses in hoc scietis quod Dominus miserit me ut facerem universa quae cernitis et non ex proprio ea corde protulerim
NUM|16|29|si consueta hominum morte interierint et visitaverit eos plaga qua et ceteri visitari solent non misit me Dominus
NUM|16|30|sin autem novam rem fecerit Dominus ut aperiens terra os suum degluttiat eos et omnia quae ad illos pertinent descenderintque viventes in infernum scietis quod blasphemaverint Dominum
NUM|16|31|confestim igitur ut cessavit loqui disrupta est terra sub pedibus eorum
NUM|16|32|et aperiens os suum devoravit illos cum tabernaculis suis et universa substantia
NUM|16|33|descenderuntque vivi in infernum operti humo et perierunt de medio multitudinis
NUM|16|34|at vero omnis Israhel qui stabat per gyrum fugit ad clamorem pereuntium dicens ne forte et nos terra degluttiat
NUM|16|35|sed et ignis egressus a Domino interfecit ducentos quinquaginta viros qui offerebant incensum
NUM|16|36|locutusque est Dominus ad Mosen dicens
NUM|16|37|praecipe Eleazaro filio Aaron sacerdotis ut tollat turibula quae iacent in incendio et ignem huc illucque dispergat quoniam sanctificata sunt
NUM|16|38|in mortibus peccatorum producatque ea in lamminas et adfigat altari eo quod oblatum sit in eis incensum Domino et sanctificata sint ut cernant ea pro signo et monumento filii Israhel
NUM|16|39|tulit ergo Eleazar sacerdos turibula aenea in quibus obtulerant hii quos incendium devoravit et produxit ea in lamminas adfigens altari
NUM|16|40|ut haberent postea filii Israhel quibus commonerentur ne quis accedat alienigena et qui non est de semine Aaron ad offerendum incensum Domino ne patiatur sicut passus est Core et omnis congregatio eius loquente Domino ad Mosen
NUM|16|41|murmuravit autem omnis multitudo filiorum Israhel sequenti die contra Mosen et Aaron dicens vos interfecistis populum Domini
NUM|16|42|cumque oreretur seditio et tumultus incresceret
NUM|16|43|Moses et Aaron fugerunt ad tabernaculum foederis quod postquam ingressi sunt operuit nubes et apparuit gloria Domini
NUM|16|44|dixitque Dominus ad Mosen
NUM|16|45|recedite de medio huius multitudinis etiam nunc delebo eos cumque iacerent in terra
NUM|16|46|dixit Moses ad Aaron tolle turibulum et hausto igne de altari mitte incensum desuper pergens cito ad populum ut roges pro eis iam enim egressa est ira a Domino et plaga desaevit
NUM|16|47|quod cum fecisset Aaron et cucurrisset ad mediam multitudinem quam iam vastabat incendium obtulit thymiama
NUM|16|48|et stans inter mortuos ac viventes pro populo deprecatus est et plaga cessavit
NUM|16|49|fuerunt autem qui percussi sunt quattuordecim milia hominum et septingenti absque his qui perierant in seditione Core
NUM|16|50|reversusque est Aaron ad Mosen ad ostium tabernaculi foederis postquam quievit interitus
NUM|17|1|et locutus est Dominus ad Mosen dicens
NUM|17|2|loquere ad filios Israhel et accipe ab eis virgas singulas per cognationes suas a cunctis principibus tribuum virgas duodecim et uniuscuiusque nomen superscribes virgae suae
NUM|17|3|nomen autem Aaron erit in tribu Levi et una virga cunctas eorum familias continebit
NUM|17|4|ponesque eas in tabernaculo foederis coram testimonio ubi loquar ad te
NUM|17|5|quem ex his elegero germinabit virga eius et cohibebo a me querimonias filiorum Israhel quibus contra vos murmurant
NUM|17|6|locutusque est Moses ad filios Israhel et dederunt ei omnes principes virgas per singulas tribus fueruntque virgae duodecim absque virga Aaron
NUM|17|7|quas cum posuisset Moses coram Domino in tabernaculo testimonii
NUM|17|8|sequenti die regressus invenit germinasse virgam Aaron in domo Levi et turgentibus gemmis eruperant flores qui foliis dilatatis in amigdalas deformati sunt
NUM|17|9|protulit ergo Moses omnes virgas de conspectu Domini ad cunctos filios Israhel videruntque et receperunt singuli virgas suas
NUM|17|10|dixitque Dominus ad Mosen refer virgam Aaron in tabernaculum testimonii ut servetur ibi in signum rebellium filiorum et quiescant querellae eorum a me ne moriantur
NUM|17|11|fecitque Moses sicut praeceperat Dominus
NUM|17|12|dixerunt autem filii Israhel ad Mosen ecce consumpti sumus omnes perivimus
NUM|17|13|quicumque accedit ad tabernaculum Domini moritur num usque ad internicionem cuncti delendi sumus
NUM|18|1|dixitque Dominus ad Aaron tu et filii tui et domus patris tui tecum portabitis iniquitatem sanctuarii et tu et filii tui simul sustinebitis peccata sacerdotii vestri
NUM|18|2|sed et fratres tuos de tribu Levi et sceptro patris tui sume tecum praestoque sint et ministrent tibi tu autem et filii tui ministrabitis in tabernaculo testimonii
NUM|18|3|excubabuntque Levitae ad praecepta tua et ad cuncta opera tabernaculi ita dumtaxat ut ad vasa sanctuarii et altare non accedant ne et illi moriantur et vos pereatis simul
NUM|18|4|sint autem tecum et excubent in custodiis tabernaculi et in omnibus caerimoniis eius alienigena non miscebitur vobis
NUM|18|5|excubate in custodia sanctuarii et in ministerio altaris ne oriatur indignatio super filios Israhel
NUM|18|6|ego dedi vobis fratres vestros Levitas de medio filiorum Israhel et tradidi donum Domino ut serviant in ministeriis tabernaculi eius
NUM|18|7|tu autem et filii tui custodite sacerdotium vestrum et omnia quae ad cultum altaris pertinent et intra velum sunt per sacerdotes administrabuntur si quis externus accesserit occidetur
NUM|18|8|locutus est Dominus ad Aaron ecce dedi tibi custodiam primitiarum mearum omnia quae sanctificantur a filiis Israhel tibi tradidi et filiis tuis pro officio sacerdotali legitima sempiterna
NUM|18|9|haec ergo accipies de his quae sanctificantur et oblata sunt Domino omnis oblatio et sacrificium et quicquid pro peccato atque delicto redditur mihi et cedet in sancta sanctorum tuum erit et filiorum tuorum
NUM|18|10|in sanctuario comedes illud mares tantum edent ex eo quia consecratum est tibi
NUM|18|11|primitias autem quas voverint et obtulerint filii Israhel tibi dedi et filiis ac filiabus tuis iure perpetuo qui mundus est in domo tua vescetur eis
NUM|18|12|omnem medullam olei et vini ac frumenti quicquid offerunt primitiarum Domino tibi dedi
NUM|18|13|universa frugum initia quas gignit humus et Domino deportantur cedent in usus tuos qui mundus est in domo tua vescetur eis
NUM|18|14|omne quod ex voto reddiderint filii Israhel tuum erit
NUM|18|15|quicquid primum erumpet e vulva cunctae carnis quam offerunt Domino sive ex hominibus sive de pecoribus fuerit tui iuris erit ita dumtaxat ut pro hominis primogenito pretium accipias et omne animal quod inmundum est redimi facias
NUM|18|16|cuius redemptio erit post unum mensem siclis argenti quinque pondere sanctuarii siclus viginti obolos habet
NUM|18|17|primogenitum autem bovis et ovis et caprae non facies redimi quia sanctificata sunt Domino sanguinem tantum eorum fundes super altare et adipes adolebis in suavissimum odorem Domino
NUM|18|18|carnes vero in usum tuum cedent sicut pectusculum consecratum et armus dexter tua erunt
NUM|18|19|omnes primitias sanctuarii quas offerunt filii Israhel Domino tibi dedi et filiis ac filiabus tuis iure perpetuo pactum salis est sempiternum coram Domino tibi ac filiis tuis
NUM|18|20|dixitque Dominus ad Aaron in terra eorum nihil possidebitis nec habebitis partem inter eos ego pars et hereditas tua in medio filiorum Israhel
NUM|18|21|filiis autem Levi dedi omnes decimas Israhelis in possessionem pro ministerio quo serviunt mihi in tabernaculo foederis
NUM|18|22|ut non accedant ultra filii Israhel ad tabernaculum nec committant peccatum mortiferum
NUM|18|23|solis filiis Levi mihi in tabernaculo servientibus et portantibus peccata populi legitimum sempiternum erit in generationibus vestris nihil aliud possidebunt
NUM|18|24|decimarum oblatione contenti quas in usus eorum et necessaria separavi
NUM|18|25|locutusque est Dominus ad Mosen dicens
NUM|18|26|praecipe Levitis atque denuntia cum acceperitis a filiis Israhel decimas quas dedi vobis primitias earum offerte Domino id est decimam partem decimae
NUM|18|27|ut reputetur vobis in oblationem primitivorum tam de areis quam de torcularibus
NUM|18|28|et universis quorum accipitis primitias offerte Domino et date Aaron sacerdoti
NUM|18|29|omnia quae offertis ex decimis et in donaria Domini separatis optima et electa erunt
NUM|18|30|dicesque ad eos si praeclara et meliora quaeque obtuleritis ex decimis reputabitur vobis quasi de area et torculari dederitis primitias
NUM|18|31|et comedetis eas in omnibus locis vestris tam vos quam familiae vestrae quia pretium est pro ministerio quo servitis in tabernaculo testimonii
NUM|18|32|et non peccabitis super hoc egregia vobis et pinguia reservantes ne polluatis oblationes filiorum Israhel et moriamini
NUM|19|1|locutusque est Dominus ad Mosen et Aaron dicens
NUM|19|2|ista est religio victimae quam constituit Dominus praecipe filiis Israhel ut adducant ad te vaccam rufam aetatis integrae in qua nulla sit macula nec portaverit iugum
NUM|19|3|tradetisque eam Eleazaro sacerdoti qui eductam extra castra immolabit in conspectu omnium
NUM|19|4|et tinguens digitum in sanguine eius asperget contra fores tabernaculi septem vicibus
NUM|19|5|conburetque eam cunctis videntibus tam pelle et carnibus eius quam sanguine et fimo flammae traditis
NUM|19|6|lignum quoque cedrinum et hysopum coccumque bis tinctum sacerdos mittet in flammam quae vaccam vorat
NUM|19|7|et tunc demum lotis vestibus et corpore suo ingredietur in castra commaculatusque erit usque ad vesperam
NUM|19|8|sed et ille qui conbuserit eam lavabit vestimenta sua et corpus et inmundus erit usque ad vesperam
NUM|19|9|colliget autem vir mundus cineres vaccae et effundet eos extra castra in loco purissimo ut sint multitudini filiorum Israhel in custodiam et in aquam aspersionis quia pro peccato vacca conbusta est
NUM|19|10|cumque laverit qui vaccae portaverat cineres vestimenta sua inmundus erit usque ad vesperum habebunt hoc filii Israhel et advenae qui habitant inter eos sanctum iure perpetuo
NUM|19|11|qui tetigerit cadaver hominis et propter hoc septem diebus fuerit inmundus
NUM|19|12|aspergetur ex hac aqua die tertio et septimo et sic mundabitur si die tertio aspersus non fuerit septimo non poterit emundari
NUM|19|13|omnis qui tetigerit humanae animae morticinum et aspersus hac commixtione non fuerit polluet tabernaculum Domini et peribit ex Israhel quia aqua expiationis non est aspersus inmundus erit et manebit spurcitia eius super eum
NUM|19|14|ista est lex hominis qui moritur in tabernaculo omnes qui ingrediuntur tentorium illius et universa vasa quae ibi sunt polluta erunt septem diebus
NUM|19|15|vas quod non habuerit operculum nec ligaturam desuper inmundum erit
NUM|19|16|si quis in agro tetigerit cadaver occisi hominis aut per se mortui sive os illius vel sepulchrum inmundus erit septem diebus
NUM|19|17|tollent de cineribus conbustionis atque peccati et mittent aquas vivas super eos in vas
NUM|19|18|in quibus cum homo mundus tinxerit hysopum asperget eo omne tentorium et cunctam supellectilem et homines huiuscemodi contagione pollutos
NUM|19|19|atque hoc modo mundus lustrabit inmundum tertio et septimo die expiatusque die septimo lavabit et se et vestimenta sua et mundus erit ad vesperam
NUM|19|20|si quis hoc ritu non fuerit expiatus peribit anima illius de medio ecclesiae quia sanctuarium Domini polluit et non est aqua lustrationis aspersus
NUM|19|21|erit hoc praeceptum legitimum sempiternum ipse quoque qui aspergit aquas lavabit vestimenta sua omnis qui tetigerit aquas expiationis inmundus erit usque ad vesperam
NUM|19|22|quicquid tetigerit inmundus inmundum faciet et anima quae horum quippiam tetigerit inmunda erit usque ad vesperum
NUM|20|1|veneruntque filii Israhel et omnis multitudo in desertum Sin mense primo et mansit populus in Cades mortuaque est ibi Maria et sepulta in eodem loco
NUM|20|2|cumque indigeret aqua populus coierunt adversum Mosen et Aaron
NUM|20|3|et versi in seditionem dixerunt utinam perissemus inter fratres nostros coram Domino
NUM|20|4|cur eduxistis ecclesiam Domini in solitudinem ut et nos et nostra iumenta moriantur
NUM|20|5|quare nos fecistis ascendere de Aegypto et adduxistis in locum istum pessimum qui seri non potest qui nec ficum gignit nec vineas nec mala granata insuper et aquam non habet ad bibendum
NUM|20|6|ingressusque Moses et Aaron dimissa multitudine tabernaculum foederis corruerunt proni in terram et apparuit gloria Domini super eos
NUM|20|7|locutusque est Dominus ad Mosen dicens
NUM|20|8|tolle virgam et congrega populum tu et Aaron frater tuus et loquimini ad petram coram eis et illa dabit aquas cumque eduxeris aquam de petra bibet omnis multitudo et iumenta eius
NUM|20|9|tulit igitur Moses virgam quae erat in conspectu Domini sicut praeceperat ei
NUM|20|10|congregata multitudine ante petram dixitque eis audite rebelles et increduli num de petra hac vobis aquam poterimus eicere
NUM|20|11|cumque elevasset Moses manum percutiens virga bis silicem egressae sunt aquae largissimae ita ut et populus biberet et iumenta
NUM|20|12|dixitque Dominus ad Mosen et Aaron quia non credidistis mihi ut sanctificaretis me coram filiis Israhel non introducetis hos populos in terram quam dabo eis
NUM|20|13|haec est aqua Contradictionis ubi iurgati sunt filii Israhel contra Dominum et sanctificatus est in eis
NUM|20|14|misit interea nuntios Moses de Cades ad regem Edom qui dicerent haec mandat frater tuus Israhel nosti omnem laborem qui adprehendit nos
NUM|20|15|quomodo descenderint patres nostri in Aegyptum et habitaverimus ibi multo tempore adflixerintque nos Aegyptii et patres nostros
NUM|20|16|et quomodo clamaverimus ad Dominum et exaudierit nos miseritque angelum qui eduxerit nos de Aegypto ecce in urbe Cades quae est in extremis finibus tuis positi
NUM|20|17|obsecramus ut nobis transire liceat per terram tuam non ibimus per agros nec per vineas non bibemus aquas de puteis tuis sed gradiemur via publica nec ad dextram nec ad sinistram declinantes donec transeamus terminos tuos
NUM|20|18|cui respondit Edom non transibis per me alioquin armatus occurram tibi
NUM|20|19|dixeruntque filii Israhel per tritam gradiemur viam et si biberimus aquas tuas nos et pecora nostra dabimus quod iustum est nulla erit in pretio difficultas tantum velociter transeamus
NUM|20|20|at ille respondit non transibis statimque egressus est obvius cum infinita multitudine et manu forti
NUM|20|21|nec voluit adquiescere deprecanti ut concederet transitum per fines suos quam ob rem devertit ab eo Israhel
NUM|20|22|cumque castra movissent de Cades venerunt in montem Or qui est in finibus terrae Edom
NUM|20|23|ubi locutus est Dominus ad Mosen
NUM|20|24|pergat inquit Aaron ad populos suos non enim intrabit terram quam dedi filiis Israhel eo quod incredulus fuerit ori meo ad aquas Contradictionis
NUM|20|25|tolle Aaron et filium eius cum eo et duces eos in montem Or
NUM|20|26|cumque nudaveris patrem veste sua indues ea Eleazarum filium eius et Aaron colligetur et morietur ibi
NUM|20|27|fecit Moses ut praeceperat Dominus et ascenderunt in montem Or coram omni multitudine
NUM|20|28|cumque Aaron spoliasset vestibus suis induit eis Eleazarum filium eius
NUM|20|29|illo mortuo in montis supercilio descendit cum Eleazaro
NUM|20|30|omnis autem multitudo videns occubuisse Aaron flevit super eo triginta diebus per cunctas familias suas
NUM|21|1|quod cum audisset Chananeus rex Arad qui habitabat ad meridiem venisse scilicet Israhel per exploratorum viam pugnavit contra illum et victor existens duxit ex eo praedam
NUM|21|2|at Israhel voto se Domino obligans ait si tradideris populum istum in manu mea delebo urbes eius
NUM|21|3|exaudivitque Dominus preces Israhel et tradidit Chananeum quem ille interfecit subversis urbibus eius et vocavit nomen loci illius Horma id est anathema
NUM|21|4|profecti sunt autem et de monte Or per viam quae ducit ad mare Rubrum ut circumirent terram Edom et taedere coepit populum itineris ac laboris
NUM|21|5|locutusque contra Deum et Mosen ait cur eduxisti nos de Aegypto ut moreremur in solitudine deest panis non sunt aquae anima nostra iam nausiat super cibo isto levissimo
NUM|21|6|quam ob rem misit Dominus in populum ignitos serpentes ad quorum plagas et mortes plurimorum
NUM|21|7|venerunt ad Mosen atque dixerunt peccavimus quia locuti sumus contra Dominum et te ora ut tollat a nobis serpentes oravit Moses pro populo
NUM|21|8|et locutus est Dominus ad eum fac serpentem et pone eum pro signo qui percussus aspexerit eum vivet
NUM|21|9|fecit ergo Moses serpentem aeneum et posuit pro signo quem cum percussi aspicerent sanabantur
NUM|21|10|profectique filii Israhel castrametati sunt in Oboth
NUM|21|11|unde egressi fixere tentoria in Hieabarim in solitudine quae respicit Moab contra orientalem plagam
NUM|21|12|et inde moventes venerunt ad torrentem Zared
NUM|21|13|quem relinquentes castrametati sunt contra Arnon quae est in deserto et prominet in finibus Amorrei siquidem Arnon terminus est Moab dividens Moabitas et Amorreos
NUM|21|14|unde dicitur in libro bellorum Domini sicut fecit in mari Rubro sic faciet in torrentibus Arnon
NUM|21|15|scopuli torrentium inclinati sunt ut requiescerent in Ar et recumberent in finibus Moabitarum
NUM|21|16|ex eo loco apparuit puteus super quo locutus est Dominus ad Mosen congrega populum et dabo ei aquam
NUM|21|17|tunc cecinit Israhel carmen istud ascendat puteus concinebant
NUM|21|18|puteus quem foderunt principes et paraverunt duces multitudinis in datore legis et in baculis suis de solitudine Matthana
NUM|21|19|de Matthana Nahalihel de Nahalihel in Bamoth
NUM|21|20|de Bamoth vallis est in regione Moab in vertice Phasga et quod respicit contra desertum
NUM|21|21|misit autem Israhel nuntios ad Seon regem Amorreorum dicens
NUM|21|22|obsecro ut transire mihi liceat per terram tuam non declinabimus in agros et vineas non bibemus aquas ex puteis via regia gradiemur donec transeamus terminos tuos
NUM|21|23|qui concedere noluit ut transiret Israhel per fines suos quin potius exercitu congregato egressus est obviam in desertum et venit in Iasa pugnavitque contra eum
NUM|21|24|a quo percussus est in ore gladii et possessa est terra eius ab Arnon usque Iebboc et filios Ammon quia forti praesidio tenebantur termini Ammanitarum
NUM|21|25|tulit ergo Israhel omnes civitates eius et habitavit in urbibus Amorrei in Esebon scilicet et viculis eius
NUM|21|26|urbs Esebon fuit regis Seon Amorrei qui pugnavit contra regem Moab et tulit omnem terram quae dicionis illius fuerat usque Arnon
NUM|21|27|idcirco dicitur in proverbio venite in Esebon aedificetur et construatur civitas Seon
NUM|21|28|ignis egressus est de Esebon flamma de oppido Seon et devoravit Ar Moabitarum et habitatores excelsorum Arnon
NUM|21|29|vae tibi Moab peristi popule Chamos dedit filios eius in fugam et filias in captivitatem regi Amorreorum Seon
NUM|21|30|iugum ipsorum disperiit ab Esebon usque Dibon lassi pervenerunt in Nophe et usque Medaba
NUM|21|31|habitavit itaque Israhel in terra Amorrei
NUM|21|32|misitque Moses qui explorarent Iazer cuius ceperunt viculos et possederunt habitatores
NUM|21|33|verteruntque se et ascenderunt per viam Basan et occurrit eis Og rex Basan cum omni populo suo pugnaturus in Edrai
NUM|21|34|dixitque Dominus ad Mosen ne timeas eum quia in manu tua tradidi illum et omnem populum ac terram eius faciesque illi sicut fecisti Seon regi Amorreorum habitatori Esebon
NUM|21|35|percusserunt igitur et hunc cum filiis suis universumque populum eius usque ad internicionem et possederunt terram illius
NUM|22|1|profectique castrametati sunt in campestribus Moab ubi trans Iordanem Hierichus sita est
NUM|22|2|videns autem Balac filius Sepphor omnia quae fecerat Israhel Amorreo
NUM|22|3|et quod pertimuissent eum Moabitae et impetum eius ferre non possent
NUM|22|4|dixit ad maiores natu Madian ita delebit hic populus omnes qui in nostris finibus commorantur quomodo solet bos herbas usque ad radices carpere ipse erat eo tempore rex in Moab
NUM|22|5|misit ergo nuntios ad Balaam filium Beor ariolum qui habitabat super flumen terrae filiorum Ammon ut vocarent eum et dicerent ecce egressus est populus ex Aegypto qui operuit superficiem terrae sedens contra me
NUM|22|6|veni igitur et maledic populo huic quia fortior me est si quo modo possim percutere et eicere eum de terra mea novi enim quod benedictus sit cui benedixeris et maledictus in quem maledicta congesseris
NUM|22|7|perrexerunt seniores Moab et maiores natu Madian habentes divinationis pretium in manibus cumque venissent ad Balaam et narrassent ei omnia verba Balac
NUM|22|8|ille respondit manete hic nocte et respondebo quicquid mihi dixerit Dominus manentibus illis apud Balaam venit Deus et ait ad eum
NUM|22|9|quid sibi volunt homines isti apud te
NUM|22|10|respondit Balac filius Sepphor rex Moabitarum misit ad me
NUM|22|11|dicens ecce populus qui egressus est de Aegypto operuit superficiem terrae veni et maledic ei si quo modo possim pugnans abicere eum
NUM|22|12|dixitque Deus ad Balaam noli ire cum eis neque maledicas populo quia benedictus est
NUM|22|13|qui mane consurgens dixit ad principes ite in terram vestram quia prohibuit me Deus venire vobiscum
NUM|22|14|reversi principes dixerunt ad Balac noluit Balaam venire nobiscum
NUM|22|15|rursum ille multo plures et nobiliores quam ante miserat misit
NUM|22|16|qui cum venissent ad Balaam dixerunt sic dicit Balac filius Sepphor ne cuncteris venire ad me
NUM|22|17|paratum honorare te et quicquid volueris dare veni et maledic populo isti
NUM|22|18|respondit Balaam si dederit mihi Balac plenam domum suam argenti et auri non potero inmutare verbum Domini Dei mei ut vel plus vel minus loquar
NUM|22|19|obsecro ut hic maneatis etiam hac nocte et scire queam quid mihi rursum respondeat Dominus
NUM|22|20|venit ergo Deus ad Balaam nocte et ait ei si vocare te venerunt homines isti surge et vade cum eis ita dumtaxat ut quod tibi praecepero facias
NUM|22|21|surrexit Balaam mane et strata asina profectus est cum eis
NUM|22|22|et iratus est Deus stetitque angelus Domini in via contra Balaam qui sedebat asinae et duos pueros habebat secum
NUM|22|23|cernens asina angelum stantem in via evaginato gladio avertit se de itinere et ibat per agrum quam cum verberaret Balaam et vellet ad semitam reducere
NUM|22|24|stetit angelus in angustiis duarum maceriarum quibus vineae cingebantur
NUM|22|25|quem videns asina iunxit se parieti et adtrivit sedentis pedem at ille iterum verberabat
NUM|22|26|et nihilominus angelus ad locum angustum transiens ubi nec ad dextram nec ad sinistram poterat deviari obvius stetit
NUM|22|27|cumque vidisset asina stantem angelum concidit sub pedibus sedentis qui iratus vehementius caedebat fuste latera
NUM|22|28|aperuitque Dominus os asinae et locuta est quid feci tibi cur percutis me ecce iam tertio
NUM|22|29|respondit Balaam quia commeruisti et inlusisti mihi utinam haberem gladium ut te percuterem
NUM|22|30|dixit asina nonne animal tuum sum cui semper sedere consuesti usque in praesentem diem dic quid simile umquam fecerim tibi at ille ait numquam
NUM|22|31|protinus aperuit Dominus oculos Balaam et vidit angelum stantem in via evaginato gladio adoravitque eum pronus in terram
NUM|22|32|cui angelus cur inquit tertio verberas asinam tuam ego veni ut adversarer tibi quia perversa est via tua mihique contraria
NUM|22|33|et nisi asina declinasset de via dans locum resistenti te occidissem et illa viveret
NUM|22|34|dixit Balaam peccavi nesciens quod tu stares contra me et nunc si displicet tibi ut vadam revertar
NUM|22|35|ait angelus vade cum istis et cave ne aliud quam praecepero tibi loquaris ivit igitur cum principibus
NUM|22|36|quod cum audisset Balac egressus est in occursum eius in oppido Moabitarum quod situm est in extremis finibus Arnon
NUM|22|37|dixitque ad Balaam misi nuntios ut vocarent te cur non statim venisti ad me an quia mercedem adventui tuo reddere nequeo
NUM|22|38|cui ille respondit ecce adsum numquid loqui potero aliud nisi quod Deus posuerit in ore meo
NUM|22|39|perrexerunt ergo simul et venerunt in urbem quae in extremis regni eius finibus erat
NUM|22|40|cumque occidisset Balac boves et oves misit ad Balaam et principes qui cum eo erant munera
NUM|22|41|mane autem facto duxit eum ad excelsa Baal et intuitus est extremam partem populi
NUM|23|1|dixitque Balaam ad Balac aedifica mihi hic septem aras et para totidem vitulos eiusdemque numeri arietes
NUM|23|2|cumque fecisset iuxta sermonem Balaam inposuerunt simul vitulum et arietem super aram
NUM|23|3|dixitque Balaam ad Balac sta paulisper iuxta holocaustum tuum donec vadam si forte occurrat mihi Dominus et quodcumque imperaverit loquar tibi
NUM|23|4|cumque abisset velociter occurrit ei Deus locutusque ad eum Balaam septem inquit aras erexi et inposui vitulum et arietem desuper
NUM|23|5|Dominus autem posuit verbum in ore eius et ait revertere ad Balac et haec loqueris
NUM|23|6|reversus invenit stantem Balac iuxta holocaustum suum et omnes principes Moabitarum
NUM|23|7|adsumptaque parabola sua dixit de Aram adduxit me Balac rex Moabitarum de montibus orientis veni inquit et maledic Iacob propera et detestare Israhel
NUM|23|8|quomodo maledicam cui non maledixit Deus qua ratione detester quem Dominus non detestatur
NUM|23|9|de summis silicibus videbo eum et de collibus considerabo illum populus solus habitabit et inter gentes non reputabitur
NUM|23|10|quis dinumerare possit pulverem Iacob et nosse numerum stirpis Israhel moriatur anima mea morte iustorum et fiant novissima mea horum similia
NUM|23|11|dixitque Balac ad Balaam quid est hoc quod agis ut malediceres inimicis vocavi te et tu e contrario benedicis eis
NUM|23|12|cui ille respondit num aliud possum loqui nisi quod iusserit Dominus
NUM|23|13|dixit ergo Balac veni mecum in alterum locum unde partem Israhelis videas et totum videre non possis inde maledicito ei
NUM|23|14|cumque duxisset eum in locum sublimem super verticem montis Phasga aedificavit Balaam septem aras et inpositis supra vitulo atque ariete
NUM|23|15|dixit ad Balac sta hic iuxta holocaustum tuum donec ego pergam obvius
NUM|23|16|cui cum Dominus occurrisset posuissetque verbum in ore eius ait revertere ad Balac et haec loqueris ei
NUM|23|17|reversus invenit eum stantem iuxta holocaustum suum et principes Moabitarum cum eo ad quem Balac quid inquit locutus est Dominus
NUM|23|18|at ille adsumpta parabola sua ait sta Balac et ausculta audi fili Sepphor
NUM|23|19|non est Deus quasi homo ut mentiatur nec ut filius hominis ut mutetur dixit ergo et non faciet locutus est et non implebit
NUM|23|20|ad benedicendum adductus sum benedictionem prohibere non valeo
NUM|23|21|non est idolum in Iacob nec videtur simulacrum in Israhel Dominus Deus eius cum eo est et clangor victoriae regis in illo
NUM|23|22|Deus eduxit eum de Aegypto cuius fortitudo similis est rinocerotis
NUM|23|23|non est augurium in Iacob nec divinatio in Israhel temporibus suis dicetur Iacob et Israheli quid operatus sit Deus
NUM|23|24|ecce populus ut leaena consurget et quasi leo erigetur non accubabit donec devoret praedam et occisorum sanguinem bibat
NUM|23|25|dixitque Balac ad Balaam nec maledicas ei nec benedicas
NUM|23|26|et ille nonne ait dixi tibi quod quicquid mihi Deus imperaret hoc facerem
NUM|23|27|et ait Balac ad eum veni et ducam te ad alium locum si forte placeat Deo ut inde maledicas eis
NUM|23|28|cumque duxisset eum super verticem montis Phogor qui respicit solitudinem
NUM|23|29|dixit ei Balaam aedifica mihi hic septem aras et para totidem vitulos eiusdemque numeri arietes
NUM|23|30|fecit Balac ut Balaam dixerat inposuitque vitulos et arietes per singulas aras
NUM|24|1|cumque vidisset Balaam quod placeret Domino ut benediceret Israheli nequaquam abiit ut ante perrexerat ut augurium quaereret sed dirigens contra desertum vultum suum
NUM|24|2|et elevans oculos vidit Israhel in tentoriis commorantem per tribus suas et inruente in se spiritu Dei
NUM|24|3|adsumpta parabola ait dixit Balaam filius Beor dixit homo cuius obturatus est oculus
NUM|24|4|dixit auditor sermonum Dei qui visionem Omnipotentis intuitus est qui cadit et sic aperiuntur oculi eius
NUM|24|5|quam pulchra tabernacula tua Iacob et tentoria tua Israhel
NUM|24|6|ut valles nemorosae ut horti iuxta fluvios inrigui ut tabernacula quae fixit Dominus quasi cedri propter aquas
NUM|24|7|fluet aqua de situla eius et semen illius erit in aquas multas tolletur propter Agag rex eius et auferetur regnum illius
NUM|24|8|Deus eduxit illum de Aegypto cuius fortitudo similis est rinocerotis devorabunt gentes hostes illius ossaque eorum confringent et perforabunt sagittis
NUM|24|9|accubans dormivit ut leo et quasi leaena quam suscitare nullus audebit qui benedixerit tibi erit ipse benedictus qui maledixerit in maledictione reputabitur
NUM|24|10|iratusque Balac contra Balaam conplosis manibus ait ad maledicendum inimicis meis vocavi te quibus e contrario tertio benedixisti
NUM|24|11|revertere ad locum tuum decreveram quidem magnifice honorare te sed Dominus privavit te honore disposito
NUM|24|12|respondit Balaam ad Balac nonne nuntiis tuis quos misisti ad me dixi
NUM|24|13|si dederit mihi Balac plenam domum suam argenti et auri non potero praeterire sermonem Domini Dei mei ut vel boni quid vel mali proferam ex corde meo sed quicquid Dominus dixerit hoc loquar
NUM|24|14|verumtamen pergens ad populum meum dabo consilium quid populus tuus huic populo faciat extremo tempore
NUM|24|15|sumpta igitur parabola rursum ait dixit Balaam filius Beor dixit homo cuius obturatus est oculus
NUM|24|16|dixit auditor sermonum Dei qui novit doctrinam Altissimi et visiones Omnipotentis videt qui cadens apertos habet oculos
NUM|24|17|videbo eum sed non modo intuebor illum sed non prope orietur stella ex Iacob et consurget virga de Israhel et percutiet duces Moab vastabitque omnes filios Seth
NUM|24|18|et erit Idumea possessio eius hereditas Seir cedet inimicis suis Israhel vero fortiter aget
NUM|24|19|de Iacob erit qui dominetur et perdat reliquias civitatis
NUM|24|20|cumque vidisset Amalech adsumens parabolam ait principium gentium Amalech cuius extrema perdentur
NUM|24|21|vidit quoque Cineum et adsumpta parabola ait robustum est quidem habitaculum tuum sed si in petra posueris nidum tuum
NUM|24|22|et fueris electus de stirpe Cain quamdiu poteris permanere Assur enim capiet te
NUM|24|23|adsumptaque parabola iterum locutus est heu quis victurus est quando ista faciet Deus
NUM|24|24|venient in trieribus de Italia superabunt Assyrios vastabuntque Hebraeos et ad extremum etiam ipsi peribunt
NUM|24|25|surrexitque Balaam et reversus est in locum suum Balac quoque via qua venerat rediit
NUM|25|1|morabatur autem eo tempore Israhel in Setthim et fornicatus est populus cum filiabus Moab
NUM|25|2|quae vocaverunt eos ad sacrificia sua at illi comederunt et adoraverunt deos earum
NUM|25|3|initiatusque est Israhel Beelphegor et iratus Dominus
NUM|25|4|ait ad Mosen tolle cunctos principes populi et suspende eos contra solem in patibulis ut avertatur furor meus ab Israhel
NUM|25|5|dixitque Moses ad iudices Israhel occidat unusquisque proximos suos qui initiati sunt Beelphegor
NUM|25|6|et ecce unus de filiis Israhel intravit coram fratribus suis ad scortum madianitin vidente Mose et omni turba filiorum Israhel qui flebant ante fores tabernaculi
NUM|25|7|quod cum vidisset Finees filius Eleazari filii Aaron sacerdotis surrexit de medio multitudinis et arrepto pugione
NUM|25|8|ingressus est post virum israhelitem in lupanar et perfodit ambos simul virum scilicet et mulierem in locis genitalibus cessavitque plaga a filiis Israhel
NUM|25|9|et occisi sunt viginti quattuor milia homines
NUM|25|10|dixitque Dominus ad Mosen
NUM|25|11|Finees filius Eleazari filii Aaron sacerdotis avertit iram meam a filiis Israhel quia zelo meo commotus est contra eos ut non ipse delerem filios Israhel in zelo meo
NUM|25|12|idcirco loquere ad eos ecce do ei pacem foederis mei
NUM|25|13|et erit tam ipsi quam semini illius pactum sacerdotii sempiternum quia zelatus est pro Deo suo et expiavit scelus filiorum Israhel
NUM|25|14|erat autem nomen viri israhelitae qui occisus est cum Madianitide Zambri filius Salu dux de cognatione et tribu Symeonis
NUM|25|15|porro mulier madianitis quae pariter interfecta est vocabatur Chozbi filia Sur principis nobilissimi Madianitarum
NUM|25|16|locutusque est Dominus ad Mosen dicens
NUM|25|17|hostes vos sentiant Madianitae et percutite eos
NUM|25|18|quia et ipsi hostiliter egerunt contra vos et decepere insidiis per idolum Phogor et Chozbi filiam ducis Madian sororem suam quae percussa est in die plagae pro sacrilegio Phogor
NUM|26|1|postquam noxiorum sanguis effusus est dixit Dominus ad Mosen et Eleazarum filium Aaron sacerdotem
NUM|26|2|numerate omnem summam filiorum Israhel a viginti annis et supra per domos et cognationes suas cunctos qui possunt ad bella procedere
NUM|26|3|locuti sunt itaque Moses et Eleazar sacerdos in campestribus Moab super Iordanem contra Hierichum ad eos qui erant
NUM|26|4|a viginti annis et supra sicut Dominus imperarat quorum iste est numerus
NUM|26|5|Ruben primogenitus Israhel huius filius Enoch a quo familia Enochitarum et Phallu a quo familia Phalluitarum
NUM|26|6|et Esrom a quo familia Esromitarum et Charmi a quo familia Charmitarum
NUM|26|7|hae sunt familiae de stirpe Ruben quarum numerus inventus est quadraginta tria milia et septingenti triginta
NUM|26|8|filius Phallu Heliab
NUM|26|9|huius filii Namuhel et Dathan et Abiram isti sunt Dathan et Abiram principes populi qui surrexerunt contra Mosen et Aaron in seditione Core quando adversum Dominum rebellaverunt
NUM|26|10|et aperiens terra os suum devoravit Core morientibus plurimis quando conbusit ignis ducentos quinquaginta viros et factum est grande miraculum
NUM|26|11|ut Core pereunte filii illius non perirent
NUM|26|12|filii Symeon per cognationes suas Namuhel ab hoc familia Namuhelitarum Iamin ab hoc familia Iaminitarum Iachin ab hoc familia Iachinitarum
NUM|26|13|Zare ab hoc familia Zareitarum Saul ab hoc familia Saulitarum
NUM|26|14|hae sunt familiae de stirpe Symeon quarum omnis numerus fuit viginti duo milia ducentorum
NUM|26|15|filii Gad per cognationes suas Sephon ab hoc familia Sephonitarum Aggi ab hoc familia Aggitarum Suni ab hoc familia Sunitarum
NUM|26|16|Ozni ab hoc familia Oznitarum Heri ab hoc familia Heritarum
NUM|26|17|Arod ab hoc familia Aroditarum Arihel ab hoc familia Arihelitarum
NUM|26|18|istae sunt familiae Gad quarum omnis numerus fuit quadraginta milia quingentorum
NUM|26|19|filii Iuda Her et Onan qui ambo mortui sunt in terra Chanaan
NUM|26|20|fueruntque filii Iuda per cognationes suas Sela a quo familia Selanitarum Phares a quo familia Pharesitarum Zare a quo familia Zareitarum
NUM|26|21|porro filii Phares Esrom a quo familia Esromitarum et Amul a quo familia Amulitarum
NUM|26|22|istae sunt familiae Iuda quarum omnis numerus fuit septuaginta milia quingentorum
NUM|26|23|filii Isachar per cognationes suas Thola a quo familia Tholaitarum Phua a quo familia Phuaitarum
NUM|26|24|Iasub a quo familia Iasubitarum Semran a quo familia Semranitarum
NUM|26|25|hae sunt cognationes Isachar quarum numerus fuit sexaginta quattuor milia trecentorum
NUM|26|26|filii Zabulon per cognationes suas Sared a quo familia Sareditarum Helon a quo familia Helonitarum Ialel a quo familia Ialelitarum
NUM|26|27|hae sunt cognationes Zabulon quarum numerus fuit sexaginta milia quingentorum
NUM|26|28|filii Ioseph per cognationes suas Manasse et Ephraim
NUM|26|29|de Manasse ortus est Machir a quo familia Machiritarum Machir genuit Galaad a quo familia Galaaditarum
NUM|26|30|Galaad habuit filios Hiezer a quo familia Hiezeritarum et Elec a quo familia Elecarum
NUM|26|31|et Asrihel a quo familia Asrihelitarum et Sechem a quo familia Sechemitarum
NUM|26|32|et Semida a quo familia Semidatarum et Epher a quo familia Epheritarum
NUM|26|33|fuit autem Epher pater Salphaad qui filios non habebat sed tantum filias quarum ista sunt nomina Maala et Noa et Egla et Melcha et Thersa
NUM|26|34|hae sunt familiae Manasse et numerus earum quinquaginta duo milia septingentorum
NUM|26|35|filii autem Ephraim per cognationes suas fuerunt hii Suthala a quo familia Suthalitarum Becher a quo familia Becheritarum Tehen a quo familia Tehenitarum
NUM|26|36|porro filius Suthala fuit Heran a quo familia Heranitarum
NUM|26|37|hae sunt cognationes filiorum Ephraim quarum numerus triginta duo milia quingentorum
NUM|26|38|isti sunt filii Ioseph per familias suas filii Beniamin in cognationibus suis Bale a quo familia Baleitarum Azbel a quo familia Azbelitarum Ahiram a quo familia Ahiramitarum
NUM|26|39|Supham a quo familia Suphamitarum Hupham a quo familia Huphamitarum
NUM|26|40|filii Bale Hered et Noeman de Hered familia Hereditarum de Noeman familia Noemitarum
NUM|26|41|hii sunt filii Beniamin per cognationes suas quorum numerus quadraginta quinque milia sescentorum
NUM|26|42|filii Dan per cognationes suas Suham a quo familia Suhamitarum hae cognationes Dan per familias suas
NUM|26|43|omnes fuere Suhamitae quorum numerus erat sexaginta quattuor milia quadringentorum
NUM|26|44|filii Aser per cognationes suas Iemna a quo familia Iemnaitarum Iessui a quo familia Iessuitarum Brie a quo familia Brieitarum
NUM|26|45|filii Brie Haber a quo familia Haberitarum et Melchihel a quo familia Melchihelitarum
NUM|26|46|nomen autem filiae Aser fuit Sara
NUM|26|47|hae cognationes filiorum Aser et numerus eorum quinquaginta tria milia quadringentorum
NUM|26|48|filii Nepthalim per cognationes suas Iessihel a quo familia Iessihelitarum Guni a quo familia Gunitarum
NUM|26|49|Iesser a quo familia Iesseritarum Sellem a quo familia Sellemitarum
NUM|26|50|hae sunt cognationes filiorum Nepthalim per familias suas quorum numerus quadraginta quinque milia quadringentorum
NUM|26|51|ista est summa filiorum Israhel qui recensiti sunt sescenta milia et mille septingenti triginta
NUM|26|52|locutusque est Dominus ad Mosen dicens
NUM|26|53|istis dividetur terra iuxta numerum vocabulorum in possessiones suas
NUM|26|54|pluribus maiorem partem dabis et paucioribus minorem singulis sicut nunc recensiti sunt tradetur possessio
NUM|26|55|ita dumtaxat ut sors terram tribubus dividat et familiis
NUM|26|56|quicquid sorte contigerit hoc vel plures accipient vel pauciores
NUM|26|57|hic quoque est numerus filiorum Levi per familias suas Gerson a quo familia Gersonitarum Caath a quo familia Caathitarum Merari a quo familia Meraritarum
NUM|26|58|hae sunt familiae Levi familia Lobni familia Hebroni familia Mooli familia Musi familia Cori at vero Caath genuit Amram
NUM|26|59|qui habuit uxorem Iochabed filiam Levi quae nata est ei in Aegypto haec genuit viro suo Amram filios Aaron et Mosen et Mariam sororem eorum
NUM|26|60|de Aaron orti sunt Nadab et Abiu et Eleazar et Ithamar
NUM|26|61|quorum Nadab et Abiu mortui sunt cum obtulissent ignem alienum coram Domino
NUM|26|62|fueruntque omnes qui numerati sunt viginti tria milia generis masculini ab uno mense et supra quia non sunt recensiti inter filios Israhel nec eis cum ceteris data possessio
NUM|26|63|hic est numerus filiorum Israhel qui descripti sunt a Mosen et Eleazaro sacerdote in campestribus Moab supra Iordanem contra Hiericho
NUM|26|64|inter quos nullus fuit eorum qui ante numerati sunt a Mose et Aaron in deserto Sinai
NUM|26|65|praedixerat enim Dominus quod omnes morerentur in solitudine nullusque remansit ex eis nisi Chaleb filius Iepphonne et Iosue filius Nun
NUM|27|1|accesserunt autem filiae Salphaad filii Epher filii Galaad filii Machir filii Manasse qui fuit filius Ioseph quarum sunt nomina Maala et Noa et Egla et Melcha et Thersa
NUM|27|2|steteruntque coram Mosen et Eleazaro sacerdote et cunctis principibus populi ad ostium tabernaculi foederis atque dixerunt
NUM|27|3|pater noster mortuus est in deserto nec fuit in seditione quae concitata est contra Dominum sub Core sed in peccato suo mortuus est hic non habuit mares filios cur tollitur nomen illius de familia sua quia non habet filium date nobis possessionem inter cognatos patris nostri
NUM|27|4|rettulitque Moses causam earum ad iudicium Domini
NUM|27|5|qui dixit ad eum
NUM|27|6|iustam rem postulant filiae Salphaad da eis possessionem inter cognatos patris sui et ei in hereditate succedant
NUM|27|7|ad filios autem Israhel loqueris haec
NUM|27|8|homo cum mortuus fuerit absque filio ad filiam eius transibit hereditas
NUM|27|9|si filiam non habuerit habebit successores fratres suos
NUM|27|10|quod si et fratres non fuerint dabitis hereditatem fratribus patris eius
NUM|27|11|sin autem nec patruos habuerit dabitur hereditas his qui ei proximi sunt eritque hoc filiis Israhel sanctum lege perpetua sicut praecepit Dominus Mosi
NUM|27|12|dixit quoque Dominus ad Mosen ascende in montem istum Abarim et contemplare inde terram quam daturus sum filiis Israhel
NUM|27|13|cumque videris eam ibis et tu ad populum tuum sicut ivit frater tuus Aaron
NUM|27|14|quia offendistis me in deserto Sin in contradictione multitudinis nec sanctificare me voluistis coram ea super aquas hae sunt aquae Contradictionis in Cades deserti Sin
NUM|27|15|cui respondit Moses
NUM|27|16|provideat Dominus Deus spirituum omnis carnis hominem qui sit super multitudinem hanc
NUM|27|17|et possit exire et intrare ante eos et educere illos vel introducere ne sit populus Domini sicut oves absque pastore
NUM|27|18|dixitque Dominus ad eum tolle Iosue filium Nun virum in quo est spiritus et pone manum tuam super eum
NUM|27|19|qui stabit coram Eleazaro sacerdote et omni multitudine
NUM|27|20|et dabis ei praecepta cunctis videntibus et partem gloriae tuae ut audiat eum omnis synagoga filiorum Israhel
NUM|27|21|pro hoc si quid agendum erit Eleazar sacerdos consulet Dominum ad verbum eius egredietur et ingredietur ipse et omnes filii Israhel cum eo et cetera multitudo
NUM|27|22|fecit Moses ut praeceperat Dominus cumque tulisset Iosue statuit eum coram Eleazaro sacerdote et omni frequentia populi
NUM|27|23|et inpositis capiti eius manibus cuncta replicavit quae mandaverat Dominus
NUM|28|1|dixit quoque Dominus ad Mosen
NUM|28|2|praecipe filiis Israhel et dices ad eos oblationem meam et panes et incensum odoris suavissimi offerte per tempora sua
NUM|28|3|haec sunt sacrificia quae offerre debetis agnos anniculos inmaculatos duos cotidie in holocaustum sempiternum
NUM|28|4|unum offeretis mane et alterum ad vesperam
NUM|28|5|decimam partem oephi similae quae conspersa sit oleo purissimo et habeat quartam partem hin
NUM|28|6|holocaustum iuge est quod obtulistis in monte Sinai in odorem suavissimum incensi Domini
NUM|28|7|et libabitis vini quartam partem hin per agnos singulos in sanctuario Domini
NUM|28|8|alterumque agnum similiter offeretis ad vesperam iuxta omnem ritum sacrificii matutini et libamentorum eius oblationem suavissimi odoris Domino
NUM|28|9|die autem sabbati offeretis duos agnos anniculos inmaculatos et duas decimas similae oleo conspersae in sacrificio et liba
NUM|28|10|quae rite funduntur per singula sabbata in holocausto sempiterno
NUM|28|11|in kalendis autem id est in mensuum exordiis offeretis holocaustum Domino vitulos de armento duos arietem unum agnos anniculos septem inmaculatos
NUM|28|12|et tres decimas similae oleo conspersae in sacrificio per singulos vitulos et duas decimas similae oleo conspersae per singulos arietes
NUM|28|13|et decimam decimae similae ex oleo in sacrificio per agnos singulos holocaustum suavissimi odoris atque incensi est Domino
NUM|28|14|libamenta autem vini quae per singulas fundenda sunt victimas ista erunt media pars hin per vitulos singulos tertia per arietem quarta per agnum hoc erit holocaustum per omnes menses qui sibi anno vertente succedunt
NUM|28|15|hircus quoque offeretur Domino pro peccatis in holocaustum sempiternum cum libamentis suis
NUM|28|16|mense autem primo quartadecima die mensis phase Domini erit
NUM|28|17|et quintadecima die sollemnitas septem diebus vescentur azymis
NUM|28|18|quarum dies prima venerabilis et sancta erit omne opus servile non facietis in ea
NUM|28|19|offeretisque incensum holocaustum Domino vitulos de armento duos arietem unum agnos anniculos inmaculatos septem
NUM|28|20|et sacrificia singulorum ex simila quae conspersa sit oleo tres decimas per singulos vitulos et duas decimas per arietem
NUM|28|21|et decimam decimae per agnos singulos id est per septem agnos
NUM|28|22|et hircum pro peccato unum ut expietur pro vobis
NUM|28|23|praeter holocaustum matutinum quod semper offertis
NUM|28|24|ita facietis per singulos dies septem dierum in fomitem ignis et in odorem suavissimum Domino qui surget de holocausto et de libationibus singulorum
NUM|28|25|dies quoque septimus celeberrimus et sanctus erit vobis omne opus servile non facietis in eo
NUM|28|26|dies etiam primitivorum quando offertis novas fruges Domino expletis ebdomadibus venerabilis et sancta erit omne opus servile non facietis in ea
NUM|28|27|offeretisque holocaustum in odorem suavissimum Domino vitulos de armento duos arietem unum et agnos anniculos inmaculatos septem
NUM|28|28|atque in sacrificiis eorum similae oleo conspersae tres decimas per singulos vitulos per arietes duas
NUM|28|29|per agnos decimam decimae qui simul sunt agni septem hircum quoque
NUM|28|30|qui mactatur pro expiatione praeter holocaustum sempiternum et liba eius
NUM|28|31|inmaculata offeretis omnia cum libationibus suis
NUM|29|1|mensis etiam septimi prima dies venerabilis et sancta erit vobis omne opus servile non facietis in ea quia dies clangoris est et tubarum
NUM|29|2|offeretisque holocaustum in odorem suavissimum Domino vitulum de armento unum arietem unum agnos anniculos inmaculatos septem
NUM|29|3|et in sacrificiis eorum similae oleo conspersae tres decimas per singulos vitulos duas decimas per arietem
NUM|29|4|unam decimam per agnum qui simul sunt agni septem
NUM|29|5|et hircum pro peccato qui offertur in expiationem populi
NUM|29|6|praeter holocaustum kalendarum cum sacrificiis suis et holocaustum sempiternum cum libationibus solitis hisdem caerimoniis offeretis in odorem suavissimum incensum Domino
NUM|29|7|decima quoque dies mensis huius septimi erit vobis sancta atque venerabilis et adfligetis animas vestras omne opus servile non facietis in ea
NUM|29|8|offeretisque holocaustum Domino in odorem suavissimum vitulum de armento unum arietem unum agnos anniculos inmaculatos septem
NUM|29|9|et in sacrificiis eorum similae oleo conspersae tres decimas per vitulos singulos duas decimas per arietem
NUM|29|10|decimam decimae per agnos singulos qui sunt simul septem agni
NUM|29|11|et hircum pro peccato absque his quae offerri pro delicto solent in expiationem et holocaustum sempiternum in sacrificio et libaminibus eorum
NUM|29|12|quintadecima vero die mensis septimi quae vobis erit sancta atque venerabilis omne opus servile non facietis in ea sed celebrabitis sollemnitatem Domino septem diebus
NUM|29|13|offeretisque holocaustum in odorem suavissimum Domino vitulos de armento tredecim arietes duos agnos anniculos quattuordecim inmaculatos
NUM|29|14|et in libamentis eorum similae oleo conspersae tres decimas per vitulos singulos qui sunt simul vituli tredecim et duas decimas arieti uno id est simul arietibus duobus
NUM|29|15|et decimam decimae agnis singulis qui sunt simul agni quattuordecim
NUM|29|16|et hircum pro peccato absque holocausto sempiterno et sacrificio et libamine eius
NUM|29|17|in die altero offeres vitulos de armento duodecim arietes duos agnos anniculos inmaculatos quattuordecim
NUM|29|18|sacrificiaque et libamina singulorum per vitulos et arietes et agnos rite celebrabis
NUM|29|19|et hircum pro peccato absque holocausto sempiterno sacrificioque eius et libamine
NUM|29|20|die tertio offeres vitulos undecim arietes duos agnos anniculos inmaculatos quattuordecim
NUM|29|21|sacrificiaque et libamina singulorum per vitulos et arietes et agnos rite celebrabis
NUM|29|22|et hircum pro peccato absque holocausto sempiterno et sacrificio et libamine eius
NUM|29|23|die quarto offeres vitulos decem arietes duos agnos anniculos inmaculatos quattuordecim
NUM|29|24|sacrificiaque eorum et libamina singulorum per vitulos et arietes et agnos rite celebrabis
NUM|29|25|et hircum pro peccato absque holocausto sempiterno sacrificioque eius et libamine
NUM|29|26|die quinto offeres vitulos novem arietes duos agnos anniculos inmaculatos quattuordecim
NUM|29|27|sacrificiaque et libamina singulorum per vitulos et arietes et agnos rite celebrabis
NUM|29|28|et hircum pro peccato absque holocausto sempiterno sacrificioque eius et libamine
NUM|29|29|die sexto offeres vitulos octo arietes duos agnos anniculos inmaculatos quattuordecim
NUM|29|30|sacrificiaque et libamina singulorum per vitulos et arietes et agnos rite celebrabis
NUM|29|31|et hircum pro peccato absque holocausto sempiterno sacrificioque eius et libamine
NUM|29|32|die septimo offeres vitulos septem arietes duos agnos anniculos inmaculatos quattuordecim
NUM|29|33|sacrificiaque et libamina singulorum per vitulos et arietes et agnos rite celebrabis
NUM|29|34|et hircum pro peccato absque holocausto sempiterno sacrificioque eius et libamine
NUM|29|35|die octavo qui est celeberrimus omne opus servile non facietis
NUM|29|36|offerentes holocaustum in odorem suavissimum Domino vitulum unum arietem unum agnos anniculos inmaculatos septem
NUM|29|37|sacrificiaque et libamina singulorum per vitulos et arietes et agnos rite celebrabis
NUM|29|38|et hircum pro peccato absque holocausto sempiterno sacrificioque eius et libamine
NUM|29|39|haec offeretis Domino in sollemnitatibus vestris praeter vota et oblationes spontaneas in holocausto in sacrificio in libamine et in hostiis pacificis
NUM|30|1|narravitque Moses filiis Israhel omnia quae ei Dominus imperarat
NUM|30|2|et locutus est ad principes tribuum filiorum Israhel iste est sermo quem praecepit Dominus
NUM|30|3|si quis virorum votum Domino voverit aut se constrinxerit iuramento non faciet irritum verbum suum sed omne quod promisit implebit
NUM|30|4|mulier si quippiam voverit et se constrinxerit iuramento quae est in domo patris sui et in aetate adhuc puellari si cognoverit pater votum quod pollicita est et iuramentum quo obligavit animam suam et tacuerit voti rea erit
NUM|30|5|quicquid pollicita est et iuravit opere conplebit
NUM|30|6|sin autem statim ut audierit contradixerit pater et vota et iuramenta eius irrita erunt nec obnoxia tenebitur sponsioni eo quod contradixerit pater
NUM|30|7|si maritum habuerit et voverit aliquid et semel verbum de ore eius egrediens animam illius obligaverit iuramento
NUM|30|8|quo die audierit vir et non contradixerit voti rea erit reddet quodcumque promiserat
NUM|30|9|sin autem audiens statim contradixerit et irritas fecerit pollicitationes eius verbaque quibus obstrinxerat animam suam propitius ei erit Dominus
NUM|30|10|vidua et repudiata quicquid voverint reddent
NUM|30|11|uxor in domo viri cum se voto constrinxerit et iuramento
NUM|30|12|si audierit vir et tacuerit nec contradixerit sponsioni reddet quodcumque promiserat
NUM|30|13|sin autem extemplo contradixerit non tenebitur promissionis rea quia maritus contradixit et Dominus ei propitius erit
NUM|30|14|si voverit et iuramento se constrinxerit ut per ieiunium vel ceterarum rerum abstinentiam adfligat animam suam in arbitrio viri erit ut faciat sive non faciat
NUM|30|15|quod si audiens vir tacuerit et in alteram diem distulerit sententiam quicquid voverat atque promiserat reddet quia statim ut audivit tacuit
NUM|30|16|sin autem contradixerit postquam rescivit portabit ipse iniquitatem eius
NUM|30|17|istae sunt leges quas constituit Dominus Mosi inter virum et uxorem inter patrem et filiam quae in puellari adhuc aetate est vel quae manet in parentis domo
NUM|31|1|locutusque est Dominus ad Mosen dicens
NUM|31|2|ulciscere prius filios Israhel de Madianitis et sic colligeris ad populum tuum
NUM|31|3|statimque Moses armate inquit ex vobis viros ad pugnam qui possint ultionem Domini expetere de Madianitis
NUM|31|4|mille viri de singulis tribubus eligantur Israhel qui mittantur ad bellum
NUM|31|5|dederuntque millenos de cunctis tribubus id est duodecim milia expeditorum ad pugnam
NUM|31|6|quos misit Moses cum Finees filio Eleazari sacerdotis vasa quoque sancta et tubas ad clangendum tradidit ei
NUM|31|7|cumque pugnassent contra Madianitas atque vicissent omnes mares occiderunt
NUM|31|8|et reges eorum Evi et Recem et Sur et Ur et Rebe quinque principes gentis Balaam quoque filium Beor interfecerunt gladio
NUM|31|9|ceperuntque mulieres eorum et parvulos omniaque pecora et cunctam supellectilem quicquid habere potuerant depopulati sunt
NUM|31|10|tam urbes quam viculos et castella flamma consumpsit
NUM|31|11|et tulerunt praedam et universa quae ceperant tam ex hominibus quam ex iumentis
NUM|31|12|et adduxerunt ad Mosen et Eleazarum sacerdotem et ad omnem multitudinem filiorum Israhel reliqua etiam utensilia portaverunt ad castra in campestribus Moab iuxta Iordanem contra Hiericho
NUM|31|13|egressi sunt autem Moses et Eleazar sacerdos et omnes principes synagogae in occursum eorum extra castra
NUM|31|14|iratusque Moses principibus exercitus tribunis et centurionibus qui venerant de bello
NUM|31|15|ait cur feminas reservastis
NUM|31|16|nonne istae sunt quae deceperunt filios Israhel ad suggestionem Balaam et praevaricari vos fecerunt in Domino super peccato Phogor unde et percussus est populus
NUM|31|17|ergo cunctos interficite quicquid est generis masculini etiam in parvulis et mulieres quae noverunt viros in coitu iugulate
NUM|31|18|puellas autem et omnes feminas virgines reservate vobis
NUM|31|19|et manete extra castra septem diebus qui occiderit hominem vel occisum tetigerit lustrabitur die tertio et septimo
NUM|31|20|et de omni praeda sive vestimentum fuerit sive vas et aliquid in utensilia praeparatum de caprarum pellibus et pilis et ligno expiabitur
NUM|31|21|Eleazar quoque sacerdos ad viros exercitus qui pugnaverant sic locutus est hoc est praeceptum legis quod mandavit Dominus Mosi
NUM|31|22|aurum et argentum et aes et ferrum et stagnum et plumbum
NUM|31|23|et omne quod potest transire per flammas igne purgabitur quicquid autem ignem non potest sustinere aqua expiationis sanctificabitur
NUM|31|24|et lavabitis vestimenta vestra die septimo et purificati postea castra intrabitis
NUM|31|25|dixitque Dominus ad Mosen
NUM|31|26|tollite summam eorum quae capta sunt ab homine usque ad pecus tu et Eleazar sacerdos et principes vulgi
NUM|31|27|dividesque ex aequo praedam inter eos qui pugnaverunt et egressi sunt ad bellum et inter omnem reliquam multitudinem
NUM|31|28|et separabis partem Domino ab his qui pugnaverunt et fuerunt in bello unam animam de quingentis tam ex hominibus quam ex bubus et asinis et ovibus
NUM|31|29|et dabis eam Eleazaro sacerdoti quia primitiae Domini sunt
NUM|31|30|ex media quoque parte filiorum Israhel accipies quinquagesimum caput hominum et boum et asinorum et ovium cunctarumque animantium et dabis ea Levitis qui excubant in custodiis tabernaculi Domini
NUM|31|31|feceruntque Moses et Eleazar sicut praeceperat Dominus
NUM|31|32|fuit autem praeda quam exercitus ceperat ovium sescenta septuaginta quinque milia
NUM|31|33|boum septuaginta duo milia
NUM|31|34|asinorum sexaginta milia et mille
NUM|31|35|animae hominum sexus feminei quae non cognoverant viros triginta duo milia
NUM|31|36|dataque est media pars his qui in proelio fuerant ovium trecenta triginta septem milia quingenta
NUM|31|37|e quibus in partem Domini supputatae sunt oves sescentae septuaginta quinque
NUM|31|38|et de bubus triginta sex milibus boves septuaginta duo
NUM|31|39|de asinis triginta milibus quingentis asini sexaginta unus
NUM|31|40|de animabus hominum sedecim milibus cesserunt in partem Domini triginta duae animae
NUM|31|41|tradiditque Moses numerum primitiarum Domini Eleazaro sacerdoti sicut ei fuerat imperatum
NUM|31|42|ex media parte filiorum Israhel quam separaverat his qui in proelio fuerant
NUM|31|43|de media vero parte quae contigerat reliquae multitudini id est de ovium trecentis triginta septem milibus quingentis
NUM|31|44|et de bubus triginta sex milibus
NUM|31|45|et de asinis triginta milibus quingentis
NUM|31|46|et de hominibus sedecim milibus
NUM|31|47|tulit Moses quinquagesimum caput et dedit Levitis qui excubant in tabernaculo Domini sicut praeceperat Dominus
NUM|31|48|cumque accessissent principes exercitus ad Mosen et tribuni centurionesque dixerunt
NUM|31|49|nos servi tui recensuimus numerum pugnatorum quos habuimus sub manu nostra et ne unus quidem defuit
NUM|31|50|ob hanc causam offerimus in donariis Domini singuli quod in praeda auri potuimus invenire periscelides et armillas anulos et dextralia ac murenulas ut depreceris pro nobis Dominum
NUM|31|51|susceperuntque Moses et Eleazar sacerdos omne aurum in diversis speciebus
NUM|31|52|pondo sedecim milia septingentos quinquaginta siclos a tribunis et centurionibus
NUM|31|53|unusquisque enim quod in praeda rapuerat suum erat
NUM|31|54|et susceptum intulerunt in tabernaculum testimonii in monumentum filiorum Israhel coram Domino
NUM|32|1|filii autem Ruben et Gad habebant pecora multa et erat illis in iumentis infinita substantia cumque vidissent Iazer et Galaad aptas alendis animalibus
NUM|32|2|venerunt ad Mosen et ad Eleazarum sacerdotem et principes multitudinis atque dixerunt
NUM|32|3|Atharoth et Dibon et Iazer et Nemra Esbon et Eleale et Sabam et Nebo et Beon
NUM|32|4|terram quam percussit Dominus in conspectu filiorum Israhel regionis uberrimae est ad pastum animalium et nos servi tui habemus iumenta plurima
NUM|32|5|precamurque si invenimus gratiam coram te ut des nobis famulis tuis eam in possessionem ne facias nos transire Iordanem
NUM|32|6|quibus respondit Moses numquid fratres vestri ibunt ad pugnam et vos hic sedebitis
NUM|32|7|cur subvertitis mentes filiorum Israhel ne transire audeant in locum quem eis daturus est Dominus
NUM|32|8|nonne ita egerunt patres vestri quando misi de Cadesbarne ad explorandam terram
NUM|32|9|cumque venissent usque ad vallem Botri lustrata omni regione subverterunt cor filiorum Israhel ut non intrarent fines quos eis Dominus dedit
NUM|32|10|qui iratus iuravit dicens
NUM|32|11|si videbunt homines isti qui ascenderunt ex Aegypto a viginti annis et supra terram quam sub iuramento pollicitus sum Abraham Isaac et Iacob et noluerunt sequi me
NUM|32|12|praeter Chaleb filium Iepphonne Cenezeum et Iosue filium Nun isti impleverunt voluntatem meam
NUM|32|13|iratusque Dominus adversum Israhel circumduxit eum per desertum quadraginta annis donec consumeretur universa generatio quae fecerat malum in conspectu eius
NUM|32|14|et ecce inquit vos surrexistis pro patribus vestris incrementa et alumni hominum peccatorum ut augeretis furorem Domini contra Israhel
NUM|32|15|qui si nolueritis sequi eum in solitudine populum derelinquet et vos causa eritis necis omnium
NUM|32|16|at illi prope accedentes dixerunt caulas ovium fabricabimus et stabula iumentorum parvulis quoque nostris urbes munitas
NUM|32|17|nos autem ipsi armati et accincti pergemus ad proelium ante filios Israhel donec introducamus eos ad loca sua parvuli nostri et quicquid habere possumus erunt in urbibus muratis propter habitatorum insidias
NUM|32|18|non revertemur in domos nostras usquequo possideant filii Israhel hereditatem suam
NUM|32|19|nec quicquam quaeremus trans Iordanem quia iam habemus possessionem nostram in orientali eius plaga
NUM|32|20|quibus Moses ait si facitis quod promittitis expediti pergite coram Domino ad pugnam
NUM|32|21|et omnis vir bellator armatus Iordanem transeat donec subvertat Dominus inimicos suos
NUM|32|22|et subiciatur ei omnis terra tunc eritis inculpabiles et apud Dominum et apud Israhel et obtinebitis regiones quas vultis coram Domino
NUM|32|23|sin autem quod dicitis non feceritis nulli dubium quin peccetis in Dominum et scitote quoniam peccatum vestrum adprehendet vos
NUM|32|24|aedificate ergo urbes parvulis vestris et caulas ac stabula ovibus ac iumentis et quod polliciti estis implete
NUM|32|25|dixeruntque filii Gad et Ruben ad Mosen servi tui sumus faciemus quod iubet dominus noster
NUM|32|26|parvulos nostros et mulieres et pecora ac iumenta relinquemus in urbibus Galaad
NUM|32|27|nos autem famuli tui omnes expediti pergemus ad bellum sicut tu domine loqueris
NUM|32|28|praecepit ergo Moses Eleazaro sacerdoti et Iosue filio Nun et principibus familiarum per tribus Israhel et dixit ad eos
NUM|32|29|si transierint filii Gad et filii Ruben vobiscum Iordanem omnes armati ad bellum coram Domino et vobis fuerit terra subiecta date eis Galaad in possessionem
NUM|32|30|sin autem noluerint transire vobiscum in terram Chanaan inter vos habitandi accipiant loca
NUM|32|31|responderuntque filii Gad et filii Ruben sicut locutus est Dominus servis suis ita faciemus
NUM|32|32|ipsi armati pergemus coram Domino in terram Chanaan et possessionem iam suscepisse nos confitemur trans Iordanem
NUM|32|33|dedit itaque Moses filiis Gad et Ruben et dimidiae tribui Manasse filii Ioseph regnum Seon regis Amorrei et regnum Og regis Basan et terram eorum cum urbibus suis per circuitum
NUM|32|34|igitur extruxerunt filii Gad Dibon et Atharoth et Aroer
NUM|32|35|Etrothsophan et Iazer Iecbaa
NUM|32|36|et Bethnemra et Betharan urbes munitas et caulas pecoribus suis
NUM|32|37|filii vero Ruben aedificaverunt Esbon et Eleale et Cariathaim
NUM|32|38|et Nabo et Baalmeon versis nominibus Sabama quoque inponentes vocabula urbibus quas extruxerant
NUM|32|39|porro filii Machir filii Manasse perrexerunt in Galaad et vastaverunt eam interfecto Amorreo habitatore eius
NUM|32|40|dedit ergo Moses terram Galaad Machir filio Manasse qui habitavit in ea
NUM|32|41|Iair autem filius Manasse abiit et occupavit vicos eius quos appellavit Avothiair id est villas Iair
NUM|32|42|Nobe quoque perrexit et adprehendit Canath cum viculis suis vocavitque eam ex nomine suo Nobe
NUM|33|1|hae sunt mansiones filiorum Israhel qui egressi sunt de Aegypto per turmas suas in manu Mosi et Aaron
NUM|33|2|quas descripsit Moses iuxta castrorum loca quae Domini iussione mutabant
NUM|33|3|profecti igitur de Ramesse mense primo quintadecima die mensis primi altera die phase filii Israhel in manu excelsa videntibus cunctis Aegyptiis
NUM|33|4|et sepelientibus primogenitos quos percusserat Dominus nam et in diis eorum exercuerat ultionem
NUM|33|5|castrametati sunt in Soccoth
NUM|33|6|et de Soccoth venerunt in Aetham quae est in extremis finibus solitudinis
NUM|33|7|inde egressi venerunt contra Phiahiroth quae respicit Beelsephon et castrametati sunt ante Magdolum
NUM|33|8|profectique de Phiahiroth transierunt per medium mare in solitudinem et ambulantes tribus diebus per desertum Aetham castrametati sunt in Mara
NUM|33|9|profectique de Mara venerunt in Helim ubi erant duodecim fontes aquarum et palmae septuaginta ibique castrametati sunt
NUM|33|10|sed et inde egressi fixere tentoria super mare Rubrum profectique de mari Rubro
NUM|33|11|castrametati sunt in deserto Sin
NUM|33|12|unde egressi venerunt in Dephca
NUM|33|13|profectique de Dephca castrametati sunt in Alus
NUM|33|14|egressi de Alus Raphidim fixere tentoria ubi aqua populo defuit ad bibendum
NUM|33|15|profectique de Raphidim castrametati sunt in deserto Sinai
NUM|33|16|sed et de solitudine Sinai egressi venerunt ad sepulchra Concupiscentiae
NUM|33|17|profectique de sepulchris Concupiscentiae castrametati sunt in Aseroth
NUM|33|18|et de Aseroth venerunt in Rethma
NUM|33|19|profectique de Rethma castrametati sunt in Remmonphares
NUM|33|20|unde egressi venerunt in Lebna
NUM|33|21|et de Lebna castrametati sunt in Ressa
NUM|33|22|egressi de Ressa venerunt in Ceelatha
NUM|33|23|unde profecti castrametati sunt in monte Sepher
NUM|33|24|egressi de monte Sepher venerunt in Arada
NUM|33|25|inde proficiscentes castrametati sunt in Maceloth
NUM|33|26|profectique de Maceloth venerunt in Thaath
NUM|33|27|de Thaath castrametati sunt in Thare
NUM|33|28|unde egressi fixerunt tentoria in Methca
NUM|33|29|et de Methca castrametati sunt in Esmona
NUM|33|30|profectique de Esmona venerunt in Moseroth
NUM|33|31|et de Moseroth castrametati sunt in Baneiacan
NUM|33|32|egressique de Baneiacan venerunt in montem Gadgad
NUM|33|33|unde profecti castrametati sunt in Hietebatha
NUM|33|34|et de Hietebatha venerunt in Ebrona
NUM|33|35|egressique de Ebrona castrametati sunt in Asiongaber
NUM|33|36|inde profecti venerunt in desertum Sin haec est Cades
NUM|33|37|egressique de Cades castrametati sunt in monte Hor in extremis finibus terrae Edom
NUM|33|38|ascenditque Aaron sacerdos montem Hor iubente Domino et ibi mortuus est anno quadragesimo egressionis filiorum Israhel ex Aegypto mense quinto prima die mensis
NUM|33|39|cum esset annorum centum viginti trium
NUM|33|40|audivitque Chananeus rex Arad qui habitabat ad meridiem in terra Chanaan venisse filios Israhel
NUM|33|41|et profecti de monte Hor castrametati sunt in Salmona
NUM|33|42|unde egressi venerunt in Phinon
NUM|33|43|profectique de Phinon castrametati sunt in Oboth
NUM|33|44|et de Oboth venerunt in Ieabarim quae est in finibus Moabitarum
NUM|33|45|profectique de Ieabarim fixere tentoria in Dibongad
NUM|33|46|unde egressi castrametati sunt in Elmondeblathaim
NUM|33|47|egressi de Elmondeblathaim venerunt ad montes Abarim contra Nabo
NUM|33|48|profectique de montibus Abarim transierunt ad campestria Moab super Iordanem contra Hiericho
NUM|33|49|ibique castrametati sunt de Bethsimon usque ad Belsattim in planioribus locis Moabitarum
NUM|33|50|ubi locutus est Dominus ad Mosen
NUM|33|51|praecipe filiis Israhel et dic ad eos quando transieritis Iordanem intrantes terram Chanaan
NUM|33|52|disperdite cunctos habitatores regionis illius confringite titulos et statuas comminuite atque omnia excelsa vastate
NUM|33|53|mundantes terram et habitantes in ea ego enim dedi vobis illam in possessionem
NUM|33|54|quam dividetis vobis sorte pluribus dabitis latiorem et paucis angustiorem singulis ut sors ceciderit ita tribuetur hereditas per tribus et familias possessio dividetur
NUM|33|55|sin autem nolueritis interficere habitatores terrae qui remanserint erunt vobis quasi clavi in oculis et lanceae in lateribus et adversabuntur vobis in terra habitationis vestrae
NUM|33|56|et quicquid illis facere cogitaram vobis faciam
NUM|34|1|locutus est Dominus ad Mosen
NUM|34|2|praecipe filiis Israhel et dices ad eos cum ingressi fueritis terram Chanaan et in possessionem vobis sorte ceciderit his finibus terminabitur
NUM|34|3|pars meridiana incipiet a solitudine Sin quae est iuxta Edom et habebit terminos contra orientem mare Salsissimum
NUM|34|4|qui circumibunt australem plagam per ascensum Scorpionis ita ut transeant Senna et perveniant in meridiem usque ad Cadesbarne unde egredientur confinia ad villam nomine Addar et tendent usque Asemona
NUM|34|5|ibitque per gyrum terminus ab Asemona usque ad torrentem Aegypti et maris Magni litore finietur
NUM|34|6|plaga autem occidentalis a mari Magno incipiet et ipso fine cludetur
NUM|34|7|porro ad septentrionalem plagam a mari Magno termini incipient pervenientes usque ad montem Altissimum
NUM|34|8|a quo venies in Emath usque ad terminos Sedada
NUM|34|9|ibuntque confinia usque Zephrona et villam Henan hii erunt termini in parte aquilonis
NUM|34|10|inde metabuntur fines contra orientalem plagam de villa Henan usque Sephama
NUM|34|11|et de Sephama descendent termini in Rebla contra fontem inde pervenient contra orientem ad mare Chenereth
NUM|34|12|et tendent usque Iordanem et ad ultimum Salsissimo cludentur mari hanc habebitis terram per fines suos in circuitu
NUM|34|13|praecepitque Moses filiis Israhel dicens haec erit terra quam possidebitis sorte et quam iussit dari Dominus novem tribubus et dimidiae tribui
NUM|34|14|tribus enim filiorum Ruben per familias suas et tribus filiorum Gad iuxta cognationum numerum media quoque tribus Manasse
NUM|34|15|id est duae semis tribus acceperunt partem suam trans Iordanem contra Hiericho ad orientalem plagam
NUM|34|16|et ait Dominus ad Mosen
NUM|34|17|haec sunt nomina virorum qui terram vobis divident Eleazar sacerdos et Iosue filius Nun
NUM|34|18|et singuli principes de tribubus singulis
NUM|34|19|quorum ista sunt vocabula de tribu Iuda Chaleb filius Iepphonne
NUM|34|20|de tribu Symeon Samuhel filius Ammiud
NUM|34|21|de tribu Beniamin Helidad filius Chaselon
NUM|34|22|de tribu filiorum Dan Bocci filius Iogli
NUM|34|23|filiorum Ioseph de tribu Manasse Hannihel filius Ephod
NUM|34|24|de tribu Ephraim Camuhel filius Sephtan
NUM|34|25|de tribu Zabulon Elisaphan filius Pharnach
NUM|34|26|de tribu Isachar dux Faltihel filius Ozan
NUM|34|27|de tribu Aser Ahiud filius Salomi
NUM|34|28|de tribu Nepthali Phedahel filius Ameiud
NUM|34|29|hii sunt quibus praecepit Dominus ut dividerent filiis Israhel terram Chanaan
NUM|35|1|haec quoque locutus est Dominus ad Mosen in campestribus Moab super Iordanem contra Hiericho
NUM|35|2|praecipe filiis Israhel ut dent Levitis de possessionibus suis
NUM|35|3|urbes ad habitandum et suburbana earum per circuitum ut ipsi in oppidis maneant et suburbana sint pecoribus ac iumentis
NUM|35|4|quae a muris civitatum forinsecus per circuitum mille passuum spatio tendentur
NUM|35|5|contra orientem duo milia erunt cubiti et contra meridiem similiter duo milia ad mare quoque quod respicit occidentem eadem mensura erit et septentrionalis plaga aequali termino finietur eruntque urbes in medio et foris suburbana
NUM|35|6|de ipsis autem oppidis quae Levitis dabitis sex erunt in fugitivorum auxilia separata ut fugiat ad ea qui fuderit sanguinem exceptis his alia quadraginta duo oppida
NUM|35|7|id est simul quadraginta octo cum suburbanis suis
NUM|35|8|ipsaeque urbes quae dabuntur de possessionibus filiorum Israhel ab his qui plus habent plures auferentur et qui minus pauciores singuli iuxta mensuram hereditatis suae dabunt oppida Levitis
NUM|35|9|ait Dominus ad Mosen
NUM|35|10|loquere filiis Israhel et dices ad eos quando transgressi fueritis Iordanem in terram Chanaan
NUM|35|11|decernite quae urbes esse debeant in praesidia fugitivorum qui nolentes sanguinem fuderint
NUM|35|12|in quibus cum fuerit profugus cognatus occisi eum non poterit occidere donec stet in conspectu multitudinis et causa illius iudicetur
NUM|35|13|de ipsis autem urbibus quae ad fugitivorum subsidia separantur
NUM|35|14|tres erunt trans Iordanem et tres in terra Chanaan
NUM|35|15|tam filiis Israhel quam advenis atque peregrinis ut confugiat ad eas qui nolens sanguinem fuderit
NUM|35|16|si quis ferro percusserit et mortuus fuerit qui percussus est reus erit homicidii et ipse morietur
NUM|35|17|si lapidem iecerit et ictus occubuerit similiter punietur
NUM|35|18|si ligno percussus interierit percussoris sanguine vindicabitur
NUM|35|19|propinquus occisi homicidam interficiet statim ut adprehenderit eum percutiet
NUM|35|20|si per odium quis hominem inpulerit vel iecerit quippiam in eum per insidias
NUM|35|21|aut cum esset inimicus manu percusserit et ille mortuus fuerit percussor homicidii reus erit cognatus occisi statim ut invenerit eum iugulabit
NUM|35|22|quod si fortuito et absque odio
NUM|35|23|et inimicitiis quicquam horum fecerit
NUM|35|24|et hoc audiente populo fuerit conprobatum atque inter percussorem et propinquum sanguinis quaestio ventilata
NUM|35|25|liberabitur innocens de ultoris manu et reducetur per sententiam in urbem ad quam confugerat manebitque ibi donec sacerdos magnus qui oleo sancto unctus est moriatur
NUM|35|26|si interfector extra fines urbium quae exulibus deputatae sunt
NUM|35|27|fuerit inventus et percussus ab eo qui ultor est sanguinis absque noxa erit qui eum occiderit
NUM|35|28|debuerat enim profugus usque ad mortem pontificis in urbe residere postquam autem ille obierit homicida revertetur in terram suam
NUM|35|29|haec sempiterna erunt et legitima in cunctis habitationibus vestris
NUM|35|30|homicida sub testibus punietur ad unius testimonium nullus condemnabitur
NUM|35|31|non accipietis pretium ab eo qui reus est sanguinis statim et ipse morietur
NUM|35|32|exules et profugi ante mortem pontificis nullo modo in urbes suas reverti poterunt
NUM|35|33|ne polluatis terram habitationis vestrae quae insontium cruore maculatur nec aliter expiari potest nisi per eius sanguinem qui alterius sanguinem fuderit
NUM|35|34|atque ita emundabitur vestra possessio me commorante vobiscum ego enim sum Dominus qui habito inter filios Israhel
NUM|36|1|accesserunt autem et principes familiarum Galaad filii Machir filii Manasse de stirpe filiorum Ioseph locutique sunt Mosi coram principibus Israhel atque dixerunt
NUM|36|2|tibi domino nostro praecepit Dominus ut terram sorte divideres filiis Israhel et ut filiabus Salphaad fratris nostri dares possessionem debitam patri
NUM|36|3|quas si alterius tribus homines uxores acceperint sequetur possessio sua et translata ad aliam tribum de nostra hereditate minuetur
NUM|36|4|atque ita fiet ut cum iobeleus id est quinquagesimus annus remissionis advenerit confundatur sortium distributio et aliorum possessio ad alios transeat
NUM|36|5|respondit Moses filiis Israhel et Domino praecipiente ait recte tribus filiorum Ioseph locuta est
NUM|36|6|et haec lex super filiabus Salphaad a Domino promulgata est nubant quibus volunt tantum ut suae tribus hominibus
NUM|36|7|ne commisceatur possessio filiorum Israhel de tribu in tribum omnes enim viri ducent uxores de tribu et cognatione sua
NUM|36|8|et cunctae feminae maritos de eadem tribu accipient ut hereditas permaneat in familiis
NUM|36|9|nec sibi misceantur tribus sed ta maneant
NUM|36|10|ut a Domino separatae sunt feceruntque filiae Salphaad ut fuerat imperatum
NUM|36|11|et nupserunt Maala et Thersa et Egla et Melcha et Noa filiis patrui sui
NUM|36|12|de familia Manasse qui fuit filius Ioseph et possessio quae illis fuerat adtributa mansit in tribu et familia patris earum
NUM|36|13|haec sunt mandata atque iudicia quae praecepit Dominus per manum Mosi ad filios Israhel in campestribus Moab super Iordanem contra Hiericho
DEUT|1|1|haec sunt verba quae locutus est Moses ad omnem Israhel trans Iordanem in solitudine campestri contra mare Rubrum inter Pharan et Thophel et Laban et Aseroth ubi auri est plurimum
DEUT|1|2|undecim diebus de Horeb per viam montis Seir usque Cadesbarne
DEUT|1|3|quadragesimo anno undecimo mense prima die mensis locutus est Moses ad filios Israhel omnia quae praeceperat illi Dominus ut diceret eis
DEUT|1|4|postquam percussit Seon regem Amorreorum qui habitavit in Esebon et Og regem Basan qui mansit in Aseroth et in Edrai
DEUT|1|5|trans Iordanem in terra Moab coepitque Moses explanare legem et dicere
DEUT|1|6|Dominus Deus noster locutus est ad nos in Horeb dicens sufficit vobis quod in hoc monte mansistis
DEUT|1|7|revertimini et venite ad montem Amorreorum et ad cetera quae ei proxima sunt campestria atque montana et humiliora loca contra meridiem et iuxta litus maris terram Chananeorum et Libani usque ad flumen magnum Eufraten
DEUT|1|8|en inquit tradidi vobis ingredimini et possidete eam super qua iuravit Dominus patribus vestris Abraham et Isaac et Iacob ut daret illam eis et semini eorum post eos
DEUT|1|9|dixique vobis illo in tempore
DEUT|1|10|non possum solus sustinere vos quia Dominus Deus vester multiplicavit vos et estis hodie sicut stellae caeli plurimae
DEUT|1|11|Dominus Deus patrum vestrorum addat ad hunc numerum multa milia et benedicat vobis sicut locutus est
DEUT|1|12|non valeo solus vestra negotia sustinere et pondus ac iurgia
DEUT|1|13|date e vobis viros sapientes et gnaros et quorum conversatio sit probata in tribubus vestris ut ponam eos vobis principes
DEUT|1|14|tunc respondistis mihi bona res est quam vis facere
DEUT|1|15|tulique de tribubus vestris viros sapientes et nobiles et constitui eos principes tribunos et centuriones et quinquagenarios ac decanos qui docerent vos singula
DEUT|1|16|praecepique eis dicens audite illos et quod iustum est iudicate sive civis sit ille sive peregrinus
DEUT|1|17|nulla erit distantia personarum ita parvum audietis ut magnum nec accipietis cuiusquam personam quia Dei iudicium est quod si difficile vobis aliquid visum fuerit referte ad me et ego audiam
DEUT|1|18|praecepique omnia quae facere deberetis
DEUT|1|19|profecti autem de Horeb transivimus per heremum terribilem et maximam quam vidistis per viam montis Amorrei sicut praeceperat Dominus Deus noster nobis cumque venissemus in Cadesbarne
DEUT|1|20|dixi vobis venistis ad montem Amorrei quem Dominus Deus noster daturus est nobis
DEUT|1|21|vide terram quam Dominus Deus tuus dat tibi ascende et posside eam sicut locutus est Dominus Deus patribus tuis noli metuere nec quicquam paveas
DEUT|1|22|et accessistis ad me omnes atque dixistis mittamus viros qui considerent terram et renuntient per quod iter debeamus ascendere et ad quas pergere civitates
DEUT|1|23|cumque mihi sermo placuisset misi e vobis duodecim viros singulos de tribubus suis
DEUT|1|24|qui cum perrexissent et ascendissent in montana venerunt usque ad vallem Botri et considerata terra
DEUT|1|25|sumentes de fructibus eius ut ostenderent ubertatem adtulerunt ad nos atque dixerunt bona est terra quam Dominus Deus noster daturus est nobis
DEUT|1|26|et noluistis ascendere sed increduli ad sermonem Domini Dei nostri
DEUT|1|27|murmurati estis in tabernaculis vestris atque dixistis odit nos Dominus et idcirco eduxit nos de terra Aegypti ut traderet in manu Amorrei atque deleret
DEUT|1|28|quo ascendemus nuntii terruerunt cor nostrum dicentes maxima multitudo est et nobis in statura procerior urbes magnae et ad caelum usque munitae filios Enacim vidimus ibi
DEUT|1|29|et dixi vobis nolite metuere nec timeatis eos
DEUT|1|30|Dominus Deus qui ductor est vester pro vobis ipse pugnabit sicut fecit in Aegypto videntibus cunctis
DEUT|1|31|et in solitudine ipse vidisti portavit te Dominus Deus tuus ut solet homo gestare parvulum filium suum in omni via per quam ambulasti donec veniretis ad locum istum
DEUT|1|32|et nec sic quidem credidistis Domino Deo vestro
DEUT|1|33|qui praecessit vos in via et metatus est locum in quo tentoria figere deberetis nocte ostendens vobis iter per ignem et die per columnam nubis
DEUT|1|34|cumque audisset Dominus vocem sermonum vestrorum iratus iuravit et ait
DEUT|1|35|non videbit quispiam de hominibus generationis huius pessimae terram bonam quam sub iuramento pollicitus sum patribus vestris
DEUT|1|36|praeter Chaleb filium Iepphonne ipse enim videbit eam et ipsi dabo terram quam calcavit et filiis eius quia secutus est Dominum
DEUT|1|37|nec miranda indignatio in populum cum mihi quoque iratus Dominus propter vos dixerit nec tu ingredieris illuc
DEUT|1|38|sed Iosue filius Nun minister tuus ipse intrabit pro te hunc exhortare et robora et ipse terram sorte dividat Israheli
DEUT|1|39|parvuli vestri de quibus dixistis quod captivi ducerentur et filii qui hodie boni ac mali ignorant distantiam ipsi ingredientur et ipsis dabo terram et possidebunt eam
DEUT|1|40|vos autem revertimini et abite in solitudinem per viam maris Rubri
DEUT|1|41|et respondistis mihi peccavimus Domino ascendemus atque pugnabimus sicut praecepit Dominus Deus noster cumque instructi armis pergeretis in montem
DEUT|1|42|ait mihi Dominus dic ad eos nolite ascendere neque pugnetis non enim sum vobiscum ne cadatis coram inimicis vestris
DEUT|1|43|locutus sum et non audistis sed adversantes imperio Domini et tumentes superbia ascendistis in montem
DEUT|1|44|itaque egressus Amorreus qui habitabat in montibus et obviam veniens persecutus est vos sicut solent apes persequi et cecidit de Seir usque Horma
DEUT|1|45|cumque reversi ploraretis coram Domino non audivit vos nec voci vestrae voluit adquiescere
DEUT|1|46|sedistis ergo in Cadesbarne multo tempore
DEUT|2|1|profectique inde venimus in solitudinem quae ducit ad mare Rubrum sicut mihi dixerat Dominus et circumivimus montem Seir longo tempore
DEUT|2|2|dixitque Dominus ad me
DEUT|2|3|sufficit vobis circumire montem istum ite contra aquilonem
DEUT|2|4|et populo praecipe dicens transibitis per terminos fratrum vestrorum filiorum Esau qui habitant in Seir et timebunt vos
DEUT|2|5|videte ergo diligenter ne moveamini contra eos neque enim dabo vobis de terra eorum quantum potest unius pedis calcare vestigium quia in possessionem Esau dedi montem Seir
DEUT|2|6|cibos emetis ab eis pecunia et comedetis aquam emptam haurietis et bibetis
DEUT|2|7|Dominus Deus tuus benedixit tibi in omni opere manuum tuarum novit iter tuum quomodo transieris solitudinem hanc magnam per quadraginta annos habitans tecum Dominus Deus tuus et nihil tibi defuit
DEUT|2|8|cumque transissemus fratres nostros filios Esau qui habitabant in Seir per viam campestrem de Helath et de Asiongaber venimus ad iter quod ducit in desertum Moab
DEUT|2|9|dixitque Dominus ad me non pugnes contra Moabitas nec ineas adversum eos proelium non enim dabo tibi quicquam de terra eorum quia filiis Loth tradidi Ar in possessionem
DEUT|2|10|Emim primi fuerunt habitatores eius populus magnus et validus et tam excelsus ut de Enacim stirpe
DEUT|2|11|quasi gigantes crederentur et essent similes filiorum Enacim denique Moabitae appellant eos Emim
DEUT|2|12|in Seir autem prius habitaverunt Horim quibus expulsis atque deletis habitaverunt filii Esau sicut fecit Israhel in terra possessionis suae quam dedit ei Dominus
DEUT|2|13|surgentes ergo ut transiremus torrentem Zared venimus ad eum
DEUT|2|14|tempus autem quo ambulavimus de Cadesbarne usque ad transitum torrentis Zared triginta octo annorum fuit donec consumeretur omnis generatio hominum bellatorum de castris sicut iuraverat Dominus
DEUT|2|15|cuius manus fuit adversum eos ut interirent de castrorum medio
DEUT|2|16|postquam autem universi ceciderunt pugnatores
DEUT|2|17|locutus est Dominus ad me dicens
DEUT|2|18|tu transibis hodie terminos Moab urbem nomine Ar
DEUT|2|19|et accedens in vicina filiorum Ammon cave ne pugnes contra eos nec movearis ad proelium non enim dabo tibi de terra filiorum Ammon quia filiis Loth dedi eam in possessionem
DEUT|2|20|terra gigantum reputata est et in ipsa olim habitaverunt gigantes quos Ammanitae vocant Zomzommim
DEUT|2|21|populus magnus et multus et procerae longitudinis sicut Enacim quos delevit Dominus a facie eorum et fecit illos habitare pro eis
DEUT|2|22|sicut fecerat filiis Esau qui habitant in Seir delens Horreos et terram eorum illis tradens quam possident usque in praesens
DEUT|2|23|Eveos quoque qui habitabant in Aserim usque Gazam Cappadoces expulerunt qui egressi de Cappadocia deleverunt eos et habitaverunt pro illis
DEUT|2|24|surgite et transite torrentem Arnon ecce tradidi in manu tua Seon regem Esebon Amorreum et terram eius incipe possidere et committe adversum eum proelium
DEUT|2|25|hodie incipiam mittere terrorem atque formidinem tuam in populos qui habitant sub omni caelo ut audito nomine tuo paveant et in morem parturientium contremescant et dolore teneantur
DEUT|2|26|misi ergo nuntios de solitudine Cademoth ad Seon regem Esebon verbis pacificis dicens
DEUT|2|27|transibimus per terram tuam publica gradiemur via non declinabimus neque ad dextram neque ad sinistram
DEUT|2|28|alimenta pretio vende nobis ut vescamur aquam pecunia tribue et sic bibemus tantum est ut nobis concedas transitum
DEUT|2|29|sicut fecerunt filii Esau qui habitant in Seir et Moabitae qui morantur in Ar donec veniamus ad Iordanem et transeamus in terram quam Dominus Deus noster daturus est nobis
DEUT|2|30|noluitque Seon rex Esebon dare nobis transitum quia induraverat Dominus Deus tuus spiritum eius et obfirmaverat cor illius ut traderetur in manus tuas sicut nunc vides
DEUT|2|31|dixitque Dominus ad me ecce coepi tradere tibi Seon et terram eius incipe possidere eam
DEUT|2|32|egressusque est Seon obviam nobis cum omni populo suo ad proelium in Iesa
DEUT|2|33|et tradidit eum Dominus Deus noster nobis percussimusque eum cum filiis et omni populo suo
DEUT|2|34|cunctasque urbes in tempore illo cepimus interfectis habitatoribus earum viris ac mulieribus et parvulis non reliquimus in eis quicquam
DEUT|2|35|absque iumentis quae in partem venere praedantium et spoliis urbium quas cepimus
DEUT|2|36|ab Aroer quae est super ripam torrentis Arnon oppido quod in valle situm est usque Galaad non fuit vicus et civitas quae nostras effugeret manus omnes tradidit Dominus Deus noster nobis
DEUT|2|37|absque terra filiorum Ammon ad quam non accessimus et cunctis quae adiacent torrenti Ieboc et urbibus montanis universisque locis a quibus nos prohibuit Dominus Deus noster
DEUT|3|1|itaque conversi ascendimus per iter Basan egressusque est Og rex Basan in occursum nobis cum populo suo ad bellandum in Edrai
DEUT|3|2|dixitque Dominus ad me ne timeas eum quia in manu tua traditus est cum omni populo ac terra sua faciesque ei sicut fecisti Seon regi Amorreorum qui habitavit in Esebon
DEUT|3|3|tradidit ergo Dominus Deus noster in manibus nostris etiam Og regem Basan et universum populum eius percussimusque eos usque ad internicionem
DEUT|3|4|vastantes cunctas civitates illius uno tempore non fuit oppidum quod nos effugeret sexaginta urbes omnem regionem Argob regni Og in Basan
DEUT|3|5|cunctae urbes erant munitae muris altissimis portisque et vectibus absque oppidis innumeris quae non habebant muros
DEUT|3|6|et delevimus eos sicut feceramus Seon regi Esebon disperdentes omnem civitatem virosque ac mulieres et parvulos
DEUT|3|7|iumenta autem et spolia urbium diripuimus
DEUT|3|8|tulimusque illo in tempore terram de manu duorum regum Amorreorum qui erant trans Iordanem a torrente Arnon usque ad montem Hermon
DEUT|3|9|quem Sidonii Sarion vocant et Amorrei Sanir
DEUT|3|10|omnes civitates quae sitae sunt in planitie et universam terram Galaad et Basan usque Selcha et Edrai civitates regni Og in Basan
DEUT|3|11|solus quippe Og rex Basan restiterat de stirpe gigantum monstratur lectus eius ferreus qui est in Rabbath filiorum Ammon novem cubitos habens longitudinis et quattuor latitudinis ad mensuram cubiti virilis manus
DEUT|3|12|terramque possedimus in tempore illo ab Aroer quae est super ripam torrentis Arnon usque ad mediam partem montis Galaad et civitates illius dedi Ruben et Gad
DEUT|3|13|reliquam autem partem Galaad et omnem Basan regni Og tradidi mediae tribui Manasse omnem regionem Argob cuncta Basan vocatur terra gigantum
DEUT|3|14|Iair filius Manasse possedit omnem regionem Argob usque ad terminos Gesuri et Machathi vocavitque ex nomine suo Basan Avothiair id est villas Iair usque in praesentem diem
DEUT|3|15|Machir quoque dedi Galaad
DEUT|3|16|et tribubus Ruben et Gad dedi terram Galaad usque ad torrentem Arnon medium torrentis et finium usque ad torrentem Ieboc qui est terminus filiorum Ammon
DEUT|3|17|et planitiem solitudinis atque Iordanem et terminos Chenereth usque ad mare Deserti quod est Salsissimum ad radices montis Phasga contra orientem
DEUT|3|18|praecepique vobis in tempore illo dicens Dominus Deus vester dat vobis terram hanc in hereditatem expediti praecedite fratres vestros filios Israhel omnes viri robusti
DEUT|3|19|absque uxoribus et parvulis ac iumentis novi enim quod plura habeatis pecora et in urbibus remanere debebunt quas tradidi vobis
DEUT|3|20|donec requiem tribuat Dominus fratribus vestris sicut vobis tribuit et possideant etiam ipsi terram quam daturus est eis trans Iordanem tunc revertetur unusquisque in possessionem suam quam dedi vobis
DEUT|3|21|Iosue quoque in tempore illo praecepi dicens oculi tui viderunt quae fecit Dominus Deus vester duobus his regibus sic faciet omnibus regnis ad quae transiturus es
DEUT|3|22|ne timeas eos Dominus enim Deus vester pugnabit pro vobis
DEUT|3|23|precatusque sum Dominum in tempore illo dicens
DEUT|3|24|Domine Deus tu coepisti ostendere servo tuo magnitudinem tuam manumque fortissimam neque enim est alius Deus vel in caelo vel in terra qui possit facere opera tua et conparari fortitudini tuae
DEUT|3|25|transibo igitur et videbo terram hanc optimam trans Iordanem et montem istum egregium et Libanum
DEUT|3|26|iratusque est Dominus mihi propter vos nec exaudivit me sed dixit mihi sufficit tibi nequaquam ultra loquaris de hac re ad me
DEUT|3|27|ascende cacumen Phasgae et oculos tuos circumfer ad occidentem et aquilonem austrumque et orientem et aspice nec enim transibis Iordanem istum
DEUT|3|28|praecipe Iosue et corrobora eum atque conforta quia ipse praecedet populum istum et dividet eis terram quam visurus es
DEUT|3|29|mansimusque in valle contra fanum Phogor
DEUT|4|1|et nunc Israhel audi praecepta et iudicia quae ego doceo te ut faciens ea vivas et ingrediens possideas terram quam Dominus Deus patrum vestrorum daturus est vobis
DEUT|4|2|non addetis ad verbum quod vobis loquor neque auferetis ex eo custodite mandata Domini Dei vestri quae ego praecipio vobis
DEUT|4|3|oculi vestri viderunt omnia quae fecit Dominus contra Beelphegor quomodo contriverit omnes cultores eius de medio vestri
DEUT|4|4|vos autem qui adheretis Domino Deo vestro vivitis universi usque in praesentem diem
DEUT|4|5|scitis quod docuerim vos praecepta atque iustitias sicut mandavit mihi Dominus Deus meus sic facietis ea in terra quam possessuri estis
DEUT|4|6|et observabitis et implebitis opere haec est enim vestra sapientia et intellectus coram populis ut audientes universa praecepta haec dicant en populus sapiens et intellegens gens magna
DEUT|4|7|nec est alia natio tam grandis quae habeat deos adpropinquantes sibi sicut Dominus Deus noster adest cunctis obsecrationibus nostris
DEUT|4|8|quae est enim alia gens sic inclita ut habeat caerimonias iustaque iudicia et universam legem quam ego proponam hodie ante oculos vestros
DEUT|4|9|custodi igitur temet ipsum et animam tuam sollicite ne obliviscaris verborum quae viderunt oculi tui et ne excedant de corde tuo cunctis diebus vitae tuae docebis ea filios ac nepotes tuos
DEUT|4|10|diem in quo stetisti coram Domino Deo tuo in Horeb quando Dominus locutus est mihi dicens congrega ad me populum ut audiat sermones meos et discat timere me omni tempore quo vivit in terra doceantque filios suos
DEUT|4|11|et accessistis ad radices montis qui ardebat usque ad caelum erantque in eo tenebrae nubes et caligo
DEUT|4|12|locutusque est Dominus ad vos de medio ignis vocem verborum eius audistis et formam penitus non vidistis
DEUT|4|13|et ostendit vobis pactum suum quod praecepit ut faceretis et decem verba quae scripsit in duabus tabulis lapideis
DEUT|4|14|mihique mandavit in illo tempore ut docerem vos caerimonias et iudicia quae facere deberetis in terra quam possessuri estis
DEUT|4|15|custodite igitur sollicite animas vestras non vidistis aliquam similitudinem in die qua locutus est Dominus vobis in Horeb de medio ignis
DEUT|4|16|ne forte decepti faciatis vobis sculptam similitudinem aut imaginem masculi vel feminae
DEUT|4|17|similitudinem omnium iumentorum quae sunt super terram vel avium sub caelo volantium
DEUT|4|18|atque reptilium quae moventur in terra sive piscium qui sub terra morantur in aquis
DEUT|4|19|ne forte oculis elevatis ad caelum videas solem et lunam et omnia astra caeli et errore deceptus adores ea et colas quae creavit Dominus Deus tuus in ministerium cunctis gentibus quae sub caelo sunt
DEUT|4|20|vos autem tulit Dominus et eduxit de fornace ferrea Aegypti ut haberet populum hereditarium sicut est in praesenti die
DEUT|4|21|iratusque est Dominus contra me propter sermones vestros et iuravit ut non transirem Iordanem nec ingrederer terram optimam quam daturus est vobis
DEUT|4|22|ecce morior in hac humo non transibo Iordanem vos transibitis et possidebitis terram egregiam
DEUT|4|23|cave nequando obliviscaris pacti Domini Dei tui quod pepigit tecum et facias tibi sculptam similitudinem eorum quae fieri Dominus prohibuit
DEUT|4|24|quia Dominus Deus tuus ignis consumens est Deus aemulator
DEUT|4|25|si genueritis filios ac nepotes et morati fueritis in terra deceptique feceritis vobis aliquam similitudinem patrantes malum coram Domino Deo vestro ut eum ad iracundiam provocetis
DEUT|4|26|testes invoco hodie caelum et terram cito perituros vos esse de terra quam transito Iordane possessuri estis non habitabitis in ea longo tempore sed delebit vos Dominus
DEUT|4|27|atque disperget in omnes gentes et remanebitis pauci in nationibus ad quas vos ducturus est Dominus
DEUT|4|28|ibique servietis diis qui hominum manu fabricati sunt ligno et lapidi qui non vident non audiunt non comedunt non odorantur
DEUT|4|29|cumque quaesieris ibi Dominum Deum tuum invenies eum si tamen toto corde quaesieris et tota tribulatione animae tuae
DEUT|4|30|postquam te invenerint omnia quae praedicta sunt novissimo tempore reverteris ad Dominum Deum tuum et audies vocem eius
DEUT|4|31|quia Deus misericors Dominus Deus tuus est non dimittet te nec omnino delebit neque obliviscetur pacti in quo iuravit patribus tuis
DEUT|4|32|interroga de diebus antiquis qui fuerunt ante te ex die quo creavit Deus hominem super terram a summo caeli usque ad summum eius si facta est aliquando huiuscemodi res aut umquam cognitum est
DEUT|4|33|ut audiret populus vocem Dei loquentis de medio ignis sicut tu audisti et vixisti
DEUT|4|34|si fecit Deus ut ingrederetur et tolleret sibi gentem de medio nationum per temptationes signa atque portenta per pugnam et robustam manum extentumque brachium et horribiles visiones iuxta omnia quae fecit pro vobis Dominus Deus vester in Aegypto videntibus oculis tuis
DEUT|4|35|ut scires quoniam Dominus ipse est Deus et non est alius praeter unum
DEUT|4|36|de caelo te fecit audire vocem suam ut doceret te et in terra ostendit tibi ignem suum maximum et audisti verba illius de medio ignis
DEUT|4|37|quia dilexit patres tuos et elegit semen eorum post eos eduxitque te praecedens in virtute sua magna ex Aegypto
DEUT|4|38|ut deleret nationes maximas et fortiores te in introitu tuo et introduceret te daretque tibi terram earum in possessionem sicut cernis in praesenti die
DEUT|4|39|scito ergo hodie et cogitato in corde tuo quod Dominus ipse sit Deus in caelo sursum et in terra deorsum et non sit alius
DEUT|4|40|custodi praecepta eius atque mandata quae ego praecipio tibi ut bene sit tibi et filiis tuis post te et permaneas multo tempore super terram quam Dominus Deus tuus daturus est tibi
DEUT|4|41|tunc separavit Moses tres civitates trans Iordanem ad orientalem plagam
DEUT|4|42|ut confugiat ad eas qui occiderit nolens proximum suum nec fuerit inimicus ante unum et alterum diem et ad harum aliquam urbium possit evadere
DEUT|4|43|Bosor in solitudine quae sita est in terra campestri de tribu Ruben et Ramoth in Galaad quae est in tribu Gad et Golam in Basan quae est in tribu Manasse
DEUT|4|44|ista est lex quam proposuit Moses coram filiis Israhel
DEUT|4|45|et haec testimonia et caerimoniae atque iudicia quae locutus est ad filios Israhel quando egressi sunt de Aegypto
DEUT|4|46|trans Iordanem in valle contra fanum Phogor in terra Seon regis Amorrei qui habitavit in Esebon quem percussit Moses filii quoque Israhel egressi ex Aegypto
DEUT|4|47|possederunt terram eius et terram Og regis Basan duorum regum Amorreorum qui erant trans Iordanem ad solis ortum
DEUT|4|48|ab Aroer quae sita est super ripam torrentis Arnon usque ad montem Sion qui est et Hermon
DEUT|4|49|omnem planitiem trans Iordanem ad orientalem plagam usque ad mare Solitudinis et usque ad radices montis Phasga
DEUT|5|1|vocavitque Moses omnem Israhelem et dixit ad eum audi Israhel caerimonias atque iudicia quae ego loquor in auribus vestris hodie discite ea et opere conplete
DEUT|5|2|Dominus Deus noster pepigit nobiscum foedus in Horeb
DEUT|5|3|non cum patribus nostris iniit pactum sed nobiscum qui inpraesentiarum sumus et vivimus
DEUT|5|4|facie ad faciem locutus est nobis in monte de medio ignis
DEUT|5|5|ego sequester et medius fui inter Dominum et vos in tempore illo ut adnuntiarem vobis verba eius timuistis enim ignem et non ascendistis in montem et ait
DEUT|5|6|ego Dominus Deus tuus qui eduxi te de terra Aegypti de domo servitutis
DEUT|5|7|non habebis deos alienos in conspectu meo
DEUT|5|8|non facies tibi sculptile nec similitudinem omnium quae in caelo sunt desuper et quae in terra deorsum et quae versantur in aquis sub terra
DEUT|5|9|non adorabis ea et non coles ego enim sum Dominus Deus tuus Deus aemulator reddens iniquitatem patrum super filios in tertiam et quartam generationem his qui oderunt me
DEUT|5|10|et faciens misericordiam in multa milia diligentibus me et custodientibus praecepta mea
DEUT|5|11|non usurpabis nomen Domini Dei tui frustra quia non erit inpunitus qui super re vana nomen eius adsumpserit
DEUT|5|12|observa diem sabbati ut sanctifices eum sicut praecepit tibi Dominus Deus tuus
DEUT|5|13|sex diebus operaberis et facies omnia opera tua
DEUT|5|14|septimus dies sabbati est id est requies Domini Dei tui non facies in eo quicquam operis tu et filius tuus et filia servus et ancilla et bos et asinus et omne iumentum tuum et peregrinus qui est intra portas tuas ut requiescat servus et ancilla tua sicut et tu
DEUT|5|15|memento quod et ipse servieris in Aegypto et eduxerit te inde Dominus Deus tuus in manu forti et brachio extento idcirco praecepit tibi ut observares diem sabbati
DEUT|5|16|honora patrem tuum et matrem sicut praecepit tibi Dominus Deus tuus ut longo vivas tempore et bene sit tibi in terra quam Dominus Deus tuus daturus est tibi
DEUT|5|17|non occides
DEUT|5|18|neque moechaberis
DEUT|5|19|furtumque non facies
DEUT|5|20|nec loqueris contra proximum tuum falsum testimonium
DEUT|5|21|non concupisces uxorem proximi tui non domum non agrum non servum non ancillam non bovem non asinum et universa quae illius sunt
DEUT|5|22|haec verba locutus est Dominus ad omnem multitudinem vestram in monte de medio ignis et nubis et caliginis voce magna nihil addens amplius et scripsit ea in duabus tabulis lapideis quas tradidit mihi
DEUT|5|23|vos autem postquam audistis vocem de medio tenebrarum et montem ardere vidistis accessistis ad me omnes principes tribuum et maiores natu atque dixistis
DEUT|5|24|ecce ostendit nobis Dominus Deus noster maiestatem et magnitudinem suam vocem eius audivimus de medio ignis et probavimus hodie quod loquente Deo cum homine vixerit homo
DEUT|5|25|cur ergo morimur et devorabit nos ignis hic maximus si enim audierimus ultra vocem Domini Dei nostri moriemur
DEUT|5|26|quid est omnis caro ut audiat vocem Dei viventis qui de medio ignis loquitur sicut nos audivimus et possit vivere
DEUT|5|27|tu magis accede et audi cuncta quae dixerit Dominus Deus noster tibi loquerisque ad nos et nos audientes faciemus ea
DEUT|5|28|quod cum audisset Dominus ait ad me audivi vocem verborum populi huius quae locuti sunt tibi bene omnia sunt locuti
DEUT|5|29|quis det talem eos habere mentem ut timeant me et custodiant universa mandata mea in omni tempore ut bene sit eis et filiis eorum in sempiternum
DEUT|5|30|vade et dic eis revertimini in tentoria vestra
DEUT|5|31|tu vero hic sta mecum et loquar tibi omnia mandata et caerimonias atque iudicia quae docebis eos ut faciant ea in terra quam dabo illis in possessionem
DEUT|5|32|custodite igitur et facite quae praecepit Dominus Deus vobis non declinabitis neque ad dextram neque ad sinistram
DEUT|5|33|sed per viam quam praecepit Dominus Deus vester ambulabitis ut vivatis et bene sit vobis et protelentur dies in terra possessionis vestrae
DEUT|6|1|haec sunt praecepta et caerimoniae atque iudicia quae mandavit Dominus Deus vester ut docerem vos et faciatis ea in terra ad quam transgredimini possidendam
DEUT|6|2|ut timeas Dominum Deum tuum et custodias omnia mandata et praecepta eius quae ego praecipio tibi et filiis ac nepotibus tuis cunctis diebus vitae tuae ut prolongentur dies tui
DEUT|6|3|audi Israhel et observa ut facias et bene sit tibi et multipliceris amplius sicut pollicitus est Dominus Deus patrum tuorum tibi terram lacte et melle manantem
DEUT|6|4|audi Israhel Dominus Deus noster Dominus unus est
DEUT|6|5|diliges Dominum Deum tuum ex toto corde tuo et ex tota anima tua et ex tota fortitudine tua
DEUT|6|6|eruntque verba haec quae ego praecipio tibi hodie in corde tuo
DEUT|6|7|et narrabis ea filiis tuis et meditaberis sedens in domo tua et ambulans in itinere dormiens atque consurgens
DEUT|6|8|et ligabis ea quasi signum in manu tua eruntque et movebuntur inter oculos tuos
DEUT|6|9|scribesque ea in limine et ostiis domus tuae
DEUT|6|10|cumque introduxerit te Dominus Deus tuus in terram pro qua iuravit patribus tuis Abraham Isaac et Iacob et dederit tibi civitates magnas et optimas quas non aedificasti
DEUT|6|11|domos plenas cunctarum opum quas non extruxisti cisternas quas non fodisti vineta et oliveta quae non plantasti
DEUT|6|12|et comederis et saturatus fueris
DEUT|6|13|cave diligenter ne obliviscaris Domini qui eduxit te de terra Aegypti de domo servitutis Dominum Deum tuum timebis et ipsi servies ac per nomen illius iurabis
DEUT|6|14|non ibitis post deos alienos cunctarum gentium quae in circuitu vestro sunt
DEUT|6|15|quoniam Deus aemulator Dominus Deus tuus in medio tui nequando irascatur furor Domini Dei tui contra te et auferat te de superficie terrae
DEUT|6|16|non temptabis Dominum Deum tuum sicut temptasti in loco temptationis
DEUT|6|17|custodi praecepta Domini Dei tui ac testimonia et caerimonias quas praecepit tibi
DEUT|6|18|et fac quod placitum est et bonum in conspectu Domini ut bene sit tibi et ingressus possideas terram optimam de qua iuravit Dominus patribus tuis
DEUT|6|19|ut deleret omnes inimicos tuos coram te sicut locutus est
DEUT|6|20|cum interrogaverit te filius tuus cras dicens quid sibi volunt testimonia haec et caerimoniae atque iudicia quae praecepit Dominus Deus noster nobis
DEUT|6|21|dices ei servi eramus Pharaonis in Aegypto et eduxit nos Dominus de Aegypto in manu forti
DEUT|6|22|fecitque signa atque prodigia magna et pessima in Aegypto contra Pharaonem et omnem domum illius in conspectu nostro
DEUT|6|23|et eduxit nos inde ut introductis daret terram super qua iuravit patribus nostris
DEUT|6|24|praecepitque nobis Dominus ut faciamus omnia legitima haec et timeamus Dominum Deum nostrum et bene sit nobis cunctis diebus vitae nostrae sicut est hodie
DEUT|6|25|eritque nostri misericors si custodierimus et fecerimus omnia praecepta eius coram Domino Deo nostro sicut mandavit nobis
DEUT|7|1|cum introduxerit te Dominus Deus tuus in terram quam possessurus ingredieris et deleverit gentes multas coram te Hettheum et Gergeseum et Amorreum Chananeum et Ferezeum et Eveum et Iebuseum septem gentes multo maioris numeri quam tu es et robustiores te
DEUT|7|2|tradideritque eas Dominus Deus tuus tibi percuties eas usque ad internicionem non inibis cum eis foedus nec misereberis earum
DEUT|7|3|neque sociabis cum eis coniugia filiam tuam non dabis filio eius nec filiam illius accipies filio tuo
DEUT|7|4|quia seducet filium tuum ne sequatur me et ut magis serviat diis alienis irasceturque furor Domini et delebit te cito
DEUT|7|5|quin potius haec facietis eis aras eorum subvertite confringite statuas lucosque succidite et sculptilia conburite
DEUT|7|6|quia populus sanctus es Domino Deo tuo te elegit Dominus Deus tuus ut sis ei populus peculiaris de cunctis populis qui sunt super terram
DEUT|7|7|non quia cunctas gentes numero vincebatis vobis iunctus est Dominus et elegit vos cum omnibus sitis populis pauciores
DEUT|7|8|sed quia dilexit vos Dominus et custodivit iuramentum quod iuravit patribus vestris eduxitque vos in manu forti et redemit de domo servitutis de manu Pharaonis regis Aegypti
DEUT|7|9|et scies quia Dominus Deus tuus ipse est Deus fortis et fidelis custodiens pactum et misericordiam diligentibus se et his qui custodiunt praecepta eius in mille generationes
DEUT|7|10|et reddens odientibus se statim ita ut disperdat eos et ultra non differat protinus eis restituens quod merentur
DEUT|7|11|custodi ergo praecepta et caerimonias atque iudicia quae ego mando tibi hodie ut facias
DEUT|7|12|si postquam audieris haec iudicia custodieris ea et feceris custodiet et Dominus Deus tuus tibi pactum et misericordiam quam iuravit patribus tuis
DEUT|7|13|et diliget te ac multiplicabit benedicetque fructui ventris tui et fructui terrae tuae frumento tuo atque vindemiae oleo et armentis gregibus ovium tuarum super terram pro qua iuravit patribus tuis ut daret eam tibi
DEUT|7|14|benedictus eris inter omnes populos non erit apud te sterilis utriusque sexus tam in hominibus quam in gregibus tuis
DEUT|7|15|auferet Dominus a te omnem languorem et infirmitates Aegypti pessimas quas novisti non inferet tibi sed cunctis hostibus tuis
DEUT|7|16|devorabis omnes populos quos Dominus Deus tuus daturus est tibi non parcet eis oculus tuus nec servies diis eorum ne sint in ruinam tui
DEUT|7|17|si dixeris in corde tuo plures sunt gentes istae quam ego quomodo potero delere eas
DEUT|7|18|noli metuere sed recordare quae fecerit Dominus Deus tuus Pharaoni et cunctis Aegyptiis
DEUT|7|19|plagas maximas quas viderunt oculi tui et signa atque portenta manumque robustam et extentum brachium ut educeret te Dominus Deus tuus sic faciet cunctis populis quos metuis
DEUT|7|20|insuper et crabrones mittet Dominus Deus tuus in eos donec deleat omnes atque disperdat qui te fugerint et latere potuerint
DEUT|7|21|non timebis eos quia Dominus Deus tuus in medio tui est Deus magnus et terribilis
DEUT|7|22|ipse consumet nationes has in conspectu tuo paulatim atque per partes non poteris delere eas pariter ne forte multiplicentur contra te bestiae terrae
DEUT|7|23|dabitque eos Dominus Deus tuus in conspectu tuo et interficiet illos donec penitus deleantur
DEUT|7|24|tradet reges eorum in manus tuas et disperdes nomina eorum sub caelo nullus poterit resistere tibi donec conteras eos
DEUT|7|25|sculptilia eorum igne conbures non concupisces argentum et aurum de quibus facta sunt neque adsumes ex eis tibi quicquam ne offendas propter ea quia abominatio est Domini Dei tui
DEUT|7|26|nec inferes quippiam ex idolo in domum tuam ne fias anathema sicut et illud est quasi spurcitiam detestaberis et velut inquinamentum ac sordes abominationi habebis quia anathema est
DEUT|8|1|omne mandatum quod ego praecipio tibi hodie cave diligenter ut facias ut possitis vivere et multiplicemini ingressique possideatis terram pro qua iuravit Dominus patribus vestris
DEUT|8|2|et recordaberis cuncti itineris per quod adduxit te Dominus Deus tuus quadraginta annis per desertum ut adfligeret te atque temptaret et nota fierent quae in tuo animo versabantur utrum custodires mandata illius an non
DEUT|8|3|adflixit te penuria et dedit tibi cibum manna quem ignorabas tu et patres tui ut ostenderet tibi quod non in solo pane vivat homo sed in omni verbo quod egreditur ex ore Domini
DEUT|8|4|vestimentum tuum quo operiebaris nequaquam vetustate defecit et pes tuus non est subtritus en quadragesimus annus est
DEUT|8|5|ut recogites in corde tuo quia sicut erudit homo filium suum sic Dominus Deus tuus erudivit te
DEUT|8|6|ut custodias mandata Domini Dei tui et ambules in viis eius et timeas eum
DEUT|8|7|Dominus enim Deus tuus introducet te in terram bonam terram rivorum aquarumque et fontium in cuius campis et montibus erumpunt fluviorum abyssi
DEUT|8|8|terram frumenti hordei vinearum in qua ficus et mala granata et oliveta nascuntur terram olei ac mellis
DEUT|8|9|ubi absque ulla penuria comedes panem tuum et rerum omnium abundantia perfrueris cuius lapides ferrum sunt et de montibus eius aeris metalla fodiuntur
DEUT|8|10|ut cum comederis et satiatus fueris benedicas Domino Deo tuo pro terra optima quam dedit tibi
DEUT|8|11|observa et cave nequando obliviscaris Domini Dei tui et neglegas mandata eius atque iudicia et caerimonias quas ego praecipio tibi hodie
DEUT|8|12|ne postquam comederis et satiatus domos pulchras aedificaveris et habitaveris in eis
DEUT|8|13|habuerisque armenta et ovium greges argenti et auri cunctarumque rerum copiam
DEUT|8|14|elevetur cor tuum et non reminiscaris Domini Dei tui qui eduxit te de terra Aegypti de domo servitutis
DEUT|8|15|et ductor tuus fuit in solitudine magna atque terribili in qua erat serpens flatu adurens et scorpio ac dipsas et nullae omnino aquae qui eduxit rivos de petra durissima
DEUT|8|16|et cibavit te manna in solitudine quod nescierunt patres tui et postquam adflixit ac probavit ad extremum misertus est tui
DEUT|8|17|ne diceres in corde tuo fortitudo mea et robur manus meae haec mihi omnia praestiterunt
DEUT|8|18|sed recorderis Domini Dei tui quod ipse tibi vires praebuerit ut impleret pactum suum super quo iuravit patribus tuis sicut praesens indicat dies
DEUT|8|19|sin autem oblitus Domini Dei tui secutus fueris alienos deos coluerisque illos et adoraveris ecce nunc praedico tibi quod omnino dispereas
DEUT|8|20|sicut gentes quas delevit Dominus in introitu tuo ita et vos peribitis si inoboedientes fueritis voci Domini Dei vestri
DEUT|9|1|audi Israhel tu transgredieris hodie Iordanem ut possideas nationes maximas et fortiores te civitates ingentes et ad caelum usque muratas
DEUT|9|2|populum magnum atque sublimem filios Enacim quos ipse vidisti et audisti quibus nullus potest ex adverso resistere
DEUT|9|3|scies ergo hodie quod Dominus Deus tuus ipse transibit ante te ignis devorans atque consumens qui conterat eos et deleat atque disperdat ante faciem tuam velociter sicut locutus est tibi
DEUT|9|4|ne dicas in corde tuo cum deleverit eos Dominus Deus tuus in conspectu tuo propter iustitiam meam introduxit me Dominus ut terram hanc possiderem cum propter impietates suas istae deletae sint nationes
DEUT|9|5|neque enim propter iustitias tuas et aequitatem cordis tui ingredieris ut possideas terras eorum sed quia illae egerunt impie te introeunte deletae sunt et ut conpleret verbum suum Dominus quod sub iuramento pollicitus est patribus tuis Abraham Isaac et Iacob
DEUT|9|6|scito igitur quod non propter iustitias tuas Dominus Deus tuus dederit tibi terram hanc optimam in possessionem cum durissimae cervicis sis populus
DEUT|9|7|memento et ne obliviscaris quomodo ad iracundiam provocaveris Dominum Deum tuum in solitudine ex eo die quo es egressus ex Aegypto usque ad locum istum semper adversum Dominum contendisti
DEUT|9|8|nam et in Horeb provocasti eum et iratus delere te voluit
DEUT|9|9|quando ascendi in montem ut acciperem tabulas lapideas tabulas pacti quod pepigit vobiscum Dominus et perseveravi in monte quadraginta diebus ac noctibus panem non comedens et aquam non bibens
DEUT|9|10|deditque mihi Dominus duas tabulas lapideas scriptas digito Dei et continentes omnia verba quae vobis in monte locutus est de medio ignis quando contio populi congregata est
DEUT|9|11|cumque transissent quadraginta dies et totidem noctes dedit mihi Dominus duas tabulas lapideas tabulas foederis
DEUT|9|12|dixitque mihi surge et descende hinc cito quia populus tuus quos eduxisti de Aegypto deseruerunt velociter viam quam demonstrasti eis feceruntque sibi conflatile
DEUT|9|13|rursumque ait Dominus ad me cerno quod populus iste durae cervicis sit
DEUT|9|14|dimitte me ut conteram eum et deleam nomen eius sub caelo et constituam te super gentem quae hac maior et fortior sit
DEUT|9|15|cumque de monte ardente descenderem et duas tabulas foederis utraque tenerem manu
DEUT|9|16|vidissemque vos peccasse Domino Deo vestro et fecisse vobis vitulum conflatilem ac deseruisse velociter viam eius quam vobis ostenderat
DEUT|9|17|proieci tabulas de manibus meis confregique eas in conspectu vestro
DEUT|9|18|et procidi ante Dominum sicut prius quadraginta diebus et noctibus panem non comedens et aquam non bibens propter omnia peccata vestra quae gessistis contra Dominum et eum ad iracundiam provocastis
DEUT|9|19|timui enim indignationem et iram illius qua adversum vos concitatus delere vos voluit et exaudivit me Dominus etiam hac vice
DEUT|9|20|adversum Aaron quoque vehementer iratus voluit eum conterere et pro illo similiter deprecatus sum
DEUT|9|21|peccatum autem vestrum quod feceratis id est vitulum arripiens igne conbusi et in frusta comminuens omninoque in pulverem redigens proieci in torrentem qui de monte descendit
DEUT|9|22|in Incendio quoque et in Temptatione et in sepulchris Concupiscentiae provocastis Dominum
DEUT|9|23|et quando misit vos de Cadesbarne dicens ascendite et possidete terram quam dedi vobis et contempsistis imperium Domini Dei vestri et non credidistis ei neque vocem eius audire voluistis
DEUT|9|24|sed semper fuistis rebelles a die qua nosse vos coepi
DEUT|9|25|et iacui coram Domino quadraginta diebus ac noctibus quibus eum suppliciter deprecabar ne deleret vos ut fuerat comminatus
DEUT|9|26|et orans dixi Domine Deus ne disperdas populum tuum et hereditatem tuam quam redemisti in magnitudine tua quos eduxisti de Aegypto in manu forti
DEUT|9|27|recordare servorum tuorum Abraham Isaac et Iacob ne aspicias duritiam populi huius et impietatem atque peccatum
DEUT|9|28|ne forte dicant habitatores terrae de qua eduxisti nos non poterat Dominus introducere eos in terram quam pollicitus est eis et oderat illos idcirco eduxit ut interficeret eos in solitudine
DEUT|9|29|qui sunt populus tuus et hereditas tua quos eduxisti in fortitudine tua magna et in brachio tuo extento
DEUT|10|1|in tempore illo dixit Dominus ad me dola tibi duas tabulas lapideas sicut priores fuerunt et ascende ad me in montem faciesque arcam ligneam
DEUT|10|2|et scribam in tabulis verba quae fuerunt in his quas ante confregisti ponesque eas in arca
DEUT|10|3|feci igitur arcam de lignis setthim cumque dolassem duas tabulas lapideas instar priorum ascendi in montem habens eas in manibus
DEUT|10|4|scripsitque in tabulis iuxta id quod prius scripserat verba decem quae locutus est Dominus ad vos in monte de medio ignis quando populus congregatus est et dedit eas mihi
DEUT|10|5|reversusque de monte descendi et posui tabulas in arcam quam feceram quae hucusque ibi sunt sicut mihi praecepit Dominus
DEUT|10|6|filii autem Israhel castra moverunt ex Beroth filiorum Iacan in Musera ubi Aaron mortuus ac sepultus est pro quo sacerdotio functus est filius eius Eleazar
DEUT|10|7|inde venerunt in Gadgad de quo loco profecti castrametati sunt in Ietabatha in terra aquarum atque torrentium
DEUT|10|8|eo tempore separavit tribum Levi ut portaret arcam foederis Domini et staret coram eo in ministerio ac benediceret in nomine illius usque in praesentem diem
DEUT|10|9|quam ob rem non habuit Levi partem neque possessionem cum fratribus suis quia ipse Dominus possessio eius est sicut promisit ei Dominus Deus tuus
DEUT|10|10|ego autem steti in monte sicut prius quadraginta diebus ac noctibus exaudivitque me Dominus etiam hac vice et te perdere noluit
DEUT|10|11|dixitque mihi vade et praecede populum ut ingrediatur et possideat terram quam iuravi patribus eorum ut traderem eis
DEUT|10|12|et nunc Israhel quid Dominus Deus tuus petit a te nisi ut timeas Dominum Deum tuum et ambules in viis eius et diligas eum ac servias Domino Deo tuo in toto corde tuo et in tota anima tua
DEUT|10|13|custodiasque mandata Domini et caerimonias eius quas ego hodie praecipio ut bene sit tibi
DEUT|10|14|en Domini Dei tui caelum est et caelum caeli terra et omnia quae in ea sunt
DEUT|10|15|et tamen patribus tuis conglutinatus est Dominus et amavit eos elegitque semen eorum post eos id est vos de cunctis gentibus sicut hodie conprobatur
DEUT|10|16|circumcidite igitur praeputium cordis vestri et cervicem vestram ne induretis amplius
DEUT|10|17|quia Dominus Deus vester ipse est Deus deorum et Dominus dominantium Deus magnus et potens et terribilis qui personam non accipit nec munera
DEUT|10|18|facit iudicium pupillo et viduae amat peregrinum et dat ei victum atque vestitum
DEUT|10|19|et vos ergo amate peregrinos quia et ipsi fuistis advenae in terra Aegypti
DEUT|10|20|Dominum Deum tuum timebis et ei servies ipsi adherebis iurabisque in nomine illius
DEUT|10|21|ipse est laus tua et Deus tuus qui fecit tibi haec magnalia et terribilia quae viderunt oculi tui
DEUT|10|22|in septuaginta animabus descenderunt patres tui in Aegyptum et ecce nunc multiplicavit te Dominus Deus tuus sicut astra caeli
DEUT|11|1|ama itaque Dominum Deum tuum et observa praecepta eius et caerimonias iudicia atque mandata omni tempore
DEUT|11|2|cognoscite hodie quae ignorant filii vestri qui non viderunt disciplinam Domini Dei vestri magnalia eius et robustam manum extentumque brachium
DEUT|11|3|signa et opera quae fecit in medio Aegypti Pharaoni regi et universae terrae eius
DEUT|11|4|omnique exercitui Aegyptiorum et equis ac curribus quomodo operuerint eos aquae Rubri maris cum vos persequerentur et deleverit eos Dominus usque in praesentem diem
DEUT|11|5|vobisque quae fecerit in solitudine donec veniretis ad hunc locum
DEUT|11|6|et Dathan atque Abiram filiis Heliab qui fuit filius Ruben quos aperto ore suo terra absorbuit cum domibus et tabernaculis et universa substantia eorum quam habebant in medio Israhelis
DEUT|11|7|oculi vestri viderunt omnia opera Domini magna quae fecit
DEUT|11|8|ut custodiatis universa mandata illius quae ego hodie praecipio vobis et possitis introire et possidere terram ad quam ingredimini
DEUT|11|9|multoque in ea vivatis tempore quam sub iuramento pollicitus est Dominus patribus vestris et semini eorum lacte et melle manantem
DEUT|11|10|terra enim ad quam ingredieris possidendam non est sicut terra Aegypti de qua existi ubi iacto semine in hortorum morem aquae ducuntur inriguae
DEUT|11|11|sed montuosa est et campestris de caelo expectans pluvias
DEUT|11|12|quam Dominus Deus tuus semper invisit et oculi illius in ea sunt a principio anni usque ad finem eius
DEUT|11|13|si ergo oboedieritis mandatis meis quae hodie praecipio vobis ut diligatis Dominum Deum vestrum et serviatis ei in toto corde vestro et in tota anima vestra
DEUT|11|14|dabo pluviam terrae vestrae temporivam et serotinam ut colligatis frumentum et vinum et oleum
DEUT|11|15|faenum ex agris ad pascenda iumenta et ut ipsi comedatis ac saturemini
DEUT|11|16|cavete ne forte decipiatur cor vestrum et recedatis a Domino serviatisque diis alienis et adoretis eos
DEUT|11|17|iratusque Dominus claudat caelum et pluviae non descendant nec terra det germen suum pereatisque velociter de terra optima quam Dominus daturus est vobis
DEUT|11|18|ponite haec verba mea in cordibus et in animis vestris et suspendite ea pro signo in manibus et inter vestros oculos conlocate
DEUT|11|19|docete filios vestros ut illa meditentur quando sederis in domo tua et ambulaveris in via et accubueris atque surrexeris
DEUT|11|20|scribes ea super postes et ianuas domus tuae
DEUT|11|21|ut multiplicentur dies tui et filiorum tuorum in terra quam iuravit Dominus patribus tuis ut daret eis quamdiu caelum inminet terrae
DEUT|11|22|si enim custodieritis mandata quae ego praecipio vobis et feceritis ea ut diligatis Dominum Deum vestrum et ambuletis in omnibus viis eius adherentes ei
DEUT|11|23|disperdet Dominus omnes gentes istas ante faciem vestram et possidebitis eas quae maiores et fortiores vobis sunt
DEUT|11|24|omnis locus quem calcaverit pes vester vester erit a deserto et Libano a flumine magno Eufraten usque ad mare occidentale erunt termini vestri
DEUT|11|25|nullus stabit contra vos terrorem vestrum et formidinem dabit Dominus Deus vester super omnem terram quam calcaturi estis sicut locutus est vobis
DEUT|11|26|en propono in conspectu vestro hodie benedictionem et maledictionem
DEUT|11|27|benedictionem si oboedieritis mandatis Domini Dei vestri quae ego praecipio vobis
DEUT|11|28|maledictionem si non audieritis mandata Domini Dei vestri sed recesseritis de via quam ego nunc ostendo vobis et ambulaveritis post deos alienos quos ignoratis
DEUT|11|29|cum introduxerit te Dominus Deus tuus in terram ad quam pergis habitandam pones benedictionem super montem Garizim maledictionem super montem Hebal
DEUT|11|30|qui sunt trans Iordanem post viam quae vergit ad solis occubitum in terra Chananei qui habitat in campestribus contra Galgalam quae est iuxta vallem tendentem et intrantem procul
DEUT|11|31|vos enim transibitis Iordanem ut possideatis terram quam Dominus Deus vester daturus est vobis et habeatis ac possideatis illam
DEUT|11|32|videte ergo ut impleatis caerimonias atque iudicia quae ego hodie ponam in conspectu vestro
DEUT|12|1|haec sunt praecepta atque iudicia quae facere debetis in terra quam Dominus Deus patrum tuorum daturus est tibi ut possideas eam cunctis diebus quibus super humum gradieris
DEUT|12|2|subvertite omnia loca in quibus coluerunt gentes quas possessuri estis deos suos super montes excelsos et colles et subter omne lignum frondosum
DEUT|12|3|dissipate aras earum et confringite statuas lucos igne conburite et idola comminuite disperdite nomina eorum de locis illis
DEUT|12|4|non facietis ita Domino Deo vestro
DEUT|12|5|sed ad locum quem elegerit Dominus Deus vester de cunctis tribubus vestris ut ponat nomen suum ibi et habitet in eo venietis
DEUT|12|6|et offeretis in illo loco holocausta et victimas vestras decimas et primitias manuum vestrarum et vota atque donaria primogenita boum et ovium
DEUT|12|7|et comedetis ibi in conspectu Domini Dei vestri ac laetabimini in cunctis ad quae miseritis manum vos et domus vestrae in quibus benedixerit vobis Dominus Deus vester
DEUT|12|8|non facietis ibi quae nos hic facimus hodie singuli quod sibi rectum videtur
DEUT|12|9|neque enim usque in praesens tempus venistis ad requiem et possessionem quam Dominus Deus daturus est vobis
DEUT|12|10|transibitis Iordanem et habitabitis in terram quam Dominus Deus vester daturus est vobis ut requiescatis a cunctis hostibus per circuitum et absque ullo timore habitetis
DEUT|12|11|in loco quem elegerit Dominus Deus vester ut sit nomen eius in eo illuc omnia quae praecipio conferetis holocausta et hostias ac decimas et primitias manuum vestrarum et quicquid praecipuum est in muneribus quae vovistis Domino
DEUT|12|12|ibi epulabimini coram Domino Deo vestro vos filii ac filiae vestrae famuli et famulae atque Levites qui in vestris urbibus commorantur neque enim habet aliam partem et possessionem inter vos
DEUT|12|13|cave ne offeras holocausta tua in omni loco quem videris
DEUT|12|14|sed in eo quem elegerit Dominus in una tribuum tuarum offeres hostias et facies quaecumque praecipio tibi
DEUT|12|15|sin autem comedere volueris et te esus carnium delectarit occide et comede iuxta benedictionem Domini Dei tui quam dedit tibi in urbibus tuis sive inmundum fuerit hoc est maculatum et debile sive mundum hoc est integrum et sine macula quod offerri licet sicut capream et cervum comedes
DEUT|12|16|absque esu dumtaxat sanguinis quod super terram quasi aquam effundes
DEUT|12|17|non poteris comedere in oppidis tuis decimam frumenti et vini et olei tui primogenita armentorum et pecorum et omnia quae voveris et sponte offerre volueris et primitias manuum tuarum
DEUT|12|18|sed coram Domino Deo tuo comedes ea in loco quem elegerit Dominus Deus tuus tu et filius tuus ac filia servus et famula atque Levites qui manet in urbibus tuis et laetaberis et reficieris coram Domino Deo tuo in cunctis ad quae extenderis manum tuam
DEUT|12|19|cave ne derelinquas Leviten omni tempore quo versaris in terra
DEUT|12|20|quando dilataverit Dominus Deus tuus terminos tuos sicut locutus est tibi et volueris vesci carnibus quas desiderat anima tua
DEUT|12|21|locus autem quem elegerit Dominus Deus tuus ut sit nomen eius ibi si procul fuerit occides de armentis et pecoribus quae habueris sicut praecepi tibi et comedes in oppidis tuis ut tibi placet
DEUT|12|22|sicut comeditur caprea et cervus ita vesceris eis et mundus et inmundus in commune vescentur
DEUT|12|23|hoc solum cave ne sanguinem comedas sanguis enim eorum pro anima est et idcirco non debes animam comedere cum carnibus
DEUT|12|24|sed super terram fundes quasi aquam
DEUT|12|25|ut sit tibi bene et filiis tuis post te cum feceris quod placet in conspectu Domini
DEUT|12|26|quae autem sanctificaveris et voveris Domino tolles et venies ad locum quem elegerit Dominus
DEUT|12|27|et offeres oblationes tuas carnem et sanguinem super altare Domini Dei tui sanguinem hostiarum fundes in altari carnibus autem ipse vesceris
DEUT|12|28|observa et audi omnia quae ego praecipio tibi ut bene sit tibi et filiis tuis post te in sempiternum cum feceris quod bonum est et placitum in conspectu Domini Dei tui
DEUT|12|29|quando disperderit Dominus Deus tuus ante faciem tuam gentes ad quas ingredieris possidendas et possederis eas atque habitaveris in terra earum
DEUT|12|30|cave ne imiteris eas postquam te fuerint introeunte subversae et requiras caerimonias earum dicens sicut coluerunt gentes istae deos suos ita et ego colam
DEUT|12|31|non facies similiter Domino Deo tuo omnes enim abominationes quas aversatur Dominus fecerunt diis suis offerentes filios et filias et conburentes igne
DEUT|12|32|quod praecipio tibi hoc tantum facito Domino nec addas quicquam nec minuas
DEUT|13|1|si surrexerit in medio tui prophetes aut qui somnium vidisse se dicat et praedixerit signum atque portentum
DEUT|13|2|et evenerit quod locutus est et dixerit tibi eamus et sequamur deos alienos quos ignoras et serviamus eis
DEUT|13|3|non audies verba prophetae illius aut somniatoris quia temptat vos Dominus Deus vester ut palam fiat utrum diligatis eum an non in toto corde et in tota anima vestra
DEUT|13|4|Dominum Deum vestrum sequimini et ipsum timete mandata illius custodite et audite vocem eius ipsi servietis et ipsi adherebitis
DEUT|13|5|propheta autem ille aut fictor somniorum interficietur quia locutus est ut vos averteret a Domino Deo vestro qui eduxit vos de terra Aegypti et redemit de domo servitutis ut errare te faceret de via quam tibi praecepit Dominus Deus tuus et auferes malum de medio tui
DEUT|13|6|si tibi voluerit persuadere frater tuus filius matris tuae aut filius tuus vel filia sive uxor quae est in sinu tuo aut amicus quem diligis ut animam tuam clam dicens eamus et serviamus diis alienis quos ignoras tu et patres tui
DEUT|13|7|cunctarum in circuitu gentium quae iuxta vel procul sunt ab initio usque ad finem terrae
DEUT|13|8|non adquiescas ei nec audias neque parcat ei oculus tuus ut miserearis et occultes eum
DEUT|13|9|sed statim interficies sit primum manus tua super eum et post te omnis populus mittat manum
DEUT|13|10|lapidibus obrutus necabitur quia voluit te abstrahere a Domino Deo tuo qui eduxit te de terra Aegypti de domo servitutis
DEUT|13|11|ut omnis Israhel audiens timeat et nequaquam ultra faciat quippiam huius rei simile
DEUT|13|12|si audieris in una urbium tuarum quas Dominus Deus tuus dabit tibi ad habitandum dicentes aliquos
DEUT|13|13|egressi sunt filii Belial de medio tui et averterunt habitatores urbis tuae atque dixerunt eamus et serviamus diis alienis quos ignoratis
DEUT|13|14|quaere sollicite et diligenter rei veritate perspecta si inveneris certum esse quod dicitur et abominationem hanc opere perpetratam
DEUT|13|15|statim percuties habitatores urbis illius in ore gladii et delebis eam omniaque quae in illa sunt usque ad pecora
DEUT|13|16|quicquid etiam supellectilis fuerit congregabis in medium platearum eius et cum ipsa civitate succendes ita ut universa consumas Domino Deo tuo et sit tumulus sempiternus non aedificabitur amplius
DEUT|13|17|et non adherebit de illo anathemate quicquam in manu tua ut avertatur Dominus ab ira furoris sui et misereatur tui multiplicetque te sicut iuravit patribus tuis
DEUT|13|18|quando audieris vocem Domini Dei tui custodiens omnia praecepta eius quae ego praecipio tibi hodie ut facias quod placitum est in conspectu Domini Dei tui
DEUT|13|19|
DEUT|14|1|filii estote Domini Dei vestri non vos incidetis nec facietis calvitium super mortuo
DEUT|14|2|quoniam populus sanctus es Domino Deo tuo et te elegit ut sis ei in populum peculiarem de cunctis gentibus quae sunt super terram
DEUT|14|3|ne comedatis quae inmunda sunt
DEUT|14|4|hoc est animal quod comedere debetis bovem et ovem et capram
DEUT|14|5|cervum capream bubalum tragelaphum pygargon orygem camelopardalum
DEUT|14|6|omne animal quod in duas partes ungulam findit et ruminat comedetis
DEUT|14|7|de his autem quae ruminant et ungulam non findunt haec comedere non debetis camelum leporem choerogyllium quia ruminant et non dividunt ungulam inmunda erunt vobis
DEUT|14|8|sus quoque quoniam dividit ungulam et non ruminat inmunda erit carnibus eorum non vescemini et cadavera non tangetis
DEUT|14|9|haec comedetis ex omnibus quae morantur in aquis quae habent pinnulas et squamas comedite
DEUT|14|10|quae absque pinnulis et squamis sunt ne comedatis quia inmunda sunt
DEUT|14|11|omnes aves mundas comedite
DEUT|14|12|inmundas ne comedatis aquilam scilicet et grypem et alietum
DEUT|14|13|ixon et vulturem ac milvum iuxta genus suum
DEUT|14|14|et omne corvini generis
DEUT|14|15|strutionem ac noctuam et larum atque accipitrem iuxta genus suum
DEUT|14|16|herodium et cycnum et ibin
DEUT|14|17|ac mergulum porphirionem et nycticoracem
DEUT|14|18|onocrotalum et charadrium singula in genere suo upupam quoque et vespertilionem
DEUT|14|19|et omne quod reptat et pinnulas habet inmundum erit nec comedetur
DEUT|14|20|omne quod mundum est comedite
DEUT|14|21|quicquid morticinum est ne vescamini ex eo peregrino qui intra portas tuas est da ut comedat aut vende ei quia tu populus sanctus Domini Dei tui es non coques hedum in lacte matris suae
DEUT|14|22|decimam partem separabis de cunctis frugibus tuis quae nascuntur in terra per annos singulos
DEUT|14|23|et comedes in conspectu Domini Dei tui in loco quem elegerit ut in eo nomen illius invocetur decimam frumenti tui et vini et olei et primogenita de armentis et ovibus tuis ut discas timere Dominum Deum tuum omni tempore
DEUT|14|24|cum autem longior fuerit via et locus quem elegerit Dominus Deus tuus tibique benedixerit nec potueris ad eum haec cuncta portare
DEUT|14|25|vendes omnia et in pretium rediges portabisque manu tua et proficisceris ad locum quem elegerit Dominus Deus tuus
DEUT|14|26|et emes ex eadem pecunia quicquid tibi placuerit sive ex armentis sive ex ovibus vinum quoque et siceram et omne quod desiderat anima tua et comedes coram Domino Deo tuo et epulaberis tu et domus tua
DEUT|14|27|et Levita qui intra portas tuas est cave ne derelinquas eum quia non habet aliam partem in possessione tua
DEUT|14|28|anno tertio separabis aliam decimam ex omnibus quae nascuntur tibi eo tempore et repones intra ianuas tuas
DEUT|14|29|venietque Levites qui aliam non habet partem nec possessionem tecum et peregrinus et pupillus ac vidua qui intra portas tuas sunt et comedent et saturabuntur ut benedicat tibi Dominus Deus tuus in cunctis operibus manuum tuarum quae feceris
DEUT|15|1|septimo anno facies remissionem
DEUT|15|2|quae hoc ordine celebrabitur cui debetur aliquid ab amico vel proximo ac fratre suo repetere non poterit quia annus remissionis est Domini
DEUT|15|3|a peregrino et advena exiges civem et propinquum repetendi non habes potestatem
DEUT|15|4|et omnino indigens et mendicus non erit inter vos ut benedicat tibi Dominus in terra quam traditurus est tibi in possessionem
DEUT|15|5|si tamen audieris vocem Domini Dei tui et custodieris universa quae iussit et quae ego hodie praecipio tibi benedicet tibi ut pollicitus est
DEUT|15|6|fenerabis gentibus multis et ipse a nullo accipies mutuum dominaberis nationibus plurimis et tui nemo dominabitur
DEUT|15|7|si unus de fratribus tuis qui morantur intra portas civitatis tuae in terra quam Dominus Deus tuus daturus est tibi ad paupertatem venerit non obdurabis cor tuum nec contrahes manum
DEUT|15|8|sed aperies eam pauperi et dabis mutuum quod eum indigere perspexeris
DEUT|15|9|cave ne forte subripiat tibi impia cogitatio et dicas in corde tuo adpropinquat septimus annus remissionis et avertas oculos a paupere fratre tuo nolens ei quod postulat mutuum commodare ne clamet contra te ad Dominum et fiat tibi in peccatum
DEUT|15|10|sed dabis ei nec ages quippiam callide in eius necessitatibus sublevandis ut benedicat tibi Dominus Deus tuus in omni tempore et in cunctis ad quae manum miseris
DEUT|15|11|non deerunt pauperes in terra habitationis tuae idcirco ego praecipio tibi ut aperias manum fratri tuo egeno et pauperi qui tecum versatur in terra
DEUT|15|12|cum tibi venditus fuerit frater tuus hebraeus aut hebraea et sex annis servierit tibi in septimo anno dimittes eum liberum
DEUT|15|13|et quem libertate donaveris nequaquam vacuum abire patieris
DEUT|15|14|sed dabis viaticum de gregibus et de area et torculari tuo quibus Dominus Deus tuus benedixerit tibi
DEUT|15|15|memento quod et ipse servieris in terra Aegypti et liberaverit te Dominus Deus tuus et idcirco ego nunc praecipiam tibi
DEUT|15|16|sin autem dixerit nolo egredi eo quod diligat te et domum tuam et bene sibi apud te esse sentiat
DEUT|15|17|adsumes subulam et perforabis aurem eius in ianua domus tuae et serviet tibi usque in aeternum ancillae quoque similiter facies
DEUT|15|18|non avertes ab eis oculos tuos quando dimiseris eos liberos quoniam iuxta mercedem mercennarii per sex annos servivit tibi ut benedicat tibi Dominus Deus tuus in cunctis operibus quae agis
DEUT|15|19|de primogenitis quae nascuntur in armentis et ovibus tuis quicquid sexus est masculini sanctificabis Domino Deo tuo non operaberis in primogenito bovis et non tondebis primogenita ovium
DEUT|15|20|in conspectu Domini Dei tui comedes ea per annos singulos in loco quem elegerit Dominus tu et domus tua
DEUT|15|21|sin autem habuerit maculam et vel claudum fuerit vel caecum aut in aliqua parte deforme vel debile non immolabitur Domino Deo tuo
DEUT|15|22|sed intra portas urbis tuae comedes illud tam mundus quam inmundus similiter vescentur eis quasi caprea et cervo
DEUT|15|23|hoc solum observabis ut sanguinem eorum non comedas sed effundas in terram quasi aquam
DEUT|16|1|observa mensem novarum frugum et verni primum temporis ut facias phase Domino Deo tuo quoniam in isto mense eduxit te Dominus Deus tuus de Aegypto nocte
DEUT|16|2|immolabisque phase Domino Deo tuo de ovibus et de bubus in loco quem elegerit Dominus Deus tuus ut habitet nomen eius ibi
DEUT|16|3|non comedes in eo panem fermentatum septem diebus comedes absque fermento adflictionis panem quoniam in pavore egressus es de Aegypto ut memineris diei egressionis tuae de Aegypto omnibus diebus vitae tuae
DEUT|16|4|non apparebit fermentum in omnibus terminis tuis septem diebus et non manebit de carnibus eius quod immolatum est vesperi in die primo mane
DEUT|16|5|non poteris immolare phase in qualibet urbium tuarum quas Dominus Deus tuus daturus est tibi
DEUT|16|6|sed in loco quem elegerit Dominus Deus tuus ut habitet nomen eius ibi immolabis phase vesperi ad solis occasum quando egressus es de Aegypto
DEUT|16|7|et coques et comedes in loco quem elegerit Dominus Deus tuus maneque consurgens vades in tabernacula tua
DEUT|16|8|sex diebus comedes azyma et in die septimo quia collecta est Domini Dei tui non facies opus
DEUT|16|9|septem ebdomadas numerabis tibi ab ea die qua falcem in segetem miseris
DEUT|16|10|et celebrabis diem festum ebdomadarum Domino Deo tuo oblationem spontaneam manus tuae quam offeres iuxta benedictionem Domini Dei tui
DEUT|16|11|et epulaberis coram Domino Deo tuo tu et filius tuus et filia tua et servus tuus et ancilla et Levites qui est intra portas tuas et advena ac pupillus et vidua qui morantur vobiscum in loco quem elegerit Dominus Deus tuus ut habitet nomen eius ibi
DEUT|16|12|et recordaberis quoniam servus fueris in Aegypto custodiesque ac facies quae praecepta sunt
DEUT|16|13|sollemnitatem quoque tabernaculorum celebrabis per septem dies quando collegeris de area et torculari fruges tuas
DEUT|16|14|et epulaberis in festivitate tua tu et filius tuus et filia et servus tuus et ancilla Levites quoque et advena et pupillus ac vidua qui intra portas tuas sunt
DEUT|16|15|septem diebus Domino Deo tuo festa celebrabis in loco quem elegerit Dominus benedicetque tibi Dominus Deus tuus in cunctis frugibus tuis et in omni opere manuum tuarum erisque in laetitia
DEUT|16|16|tribus vicibus per annum apparebit omne masculinum tuum in conspectu Domini Dei tui in loco quem elegerit in sollemnitate azymorum et in sollemnitate ebdomadarum et in sollemnitate tabernaculorum non apparebit ante Dominum vacuus
DEUT|16|17|sed offeret unusquisque secundum quod habuerit iuxta benedictionem Domini Dei sui quam dederit ei
DEUT|16|18|iudices et magistros constitues in omnibus portis tuis quas Dominus Deus tuus dederit tibi per singulas tribus tuas ut iudicent populum iusto iudicio
DEUT|16|19|nec in alteram partem declinent non accipies personam nec munera quia munera excaecant oculos sapientium et mutant verba iustorum
DEUT|16|20|iuste quod iustum est persequeris ut vivas et possideas terram quam Dominus Deus tuus dederit tibi
DEUT|16|21|non plantabis lucum et omnem arborem iuxta altare Domini Dei tui
DEUT|16|22|nec facies tibi atque constitues statuam quae odit Dominus Deus tuus
DEUT|17|1|non immolabis Domino Deo tuo bovem et ovem in quo est macula aut quippiam vitii quia abominatio est Domini Dei tui
DEUT|17|2|cum repperti fuerint apud te intra unam portarum tuarum quas Dominus Deus tuus dabit tibi vir aut mulier qui faciant malum in conspectu Domini Dei tui et transgrediantur pactum illius
DEUT|17|3|ut vadant et serviant diis alienis et adorent eos solem et lunam et omnem militiam caeli quae non praecepi
DEUT|17|4|et hoc tibi fuerit nuntiatum audiensque inquisieris diligenter et verum esse reppereris et abominatio facta est in Israhel
DEUT|17|5|educes virum ac mulierem qui rem sceleratissimam perpetrarunt ad portas civitatis tuae et lapidibus obruentur
DEUT|17|6|in ore duorum aut trium testium peribit qui interficietur nemo occidatur uno contra se dicente testimonium
DEUT|17|7|manus testium prima interficiet eum et manus reliqui populi extrema mittetur ut auferas malum de medio tui
DEUT|17|8|si difficile et ambiguum apud te iudicium esse perspexeris inter sanguinem et sanguinem causam et causam lepram et non lepram et iudicum intra portas tuas videris verba variari surge et ascende ad locum quem elegerit Dominus Deus tuus
DEUT|17|9|veniesque ad sacerdotes levitici generis et ad iudicem qui fuerit illo tempore quaeresque ab eis qui indicabunt tibi iudicii veritatem
DEUT|17|10|et facies quodcumque dixerint qui praesunt loco quem elegerit Dominus et docuerint te
DEUT|17|11|iuxta legem eius sequeris sententiam eorum nec declinabis ad dextram vel ad sinistram
DEUT|17|12|qui autem superbierit nolens oboedire sacerdotis imperio qui eo tempore ministrat Domino Deo tuo et decreto iudicis morietur homo ille et auferes malum de Israhel
DEUT|17|13|cunctusque populus audiens timebit ut nullus deinceps intumescat superbia
DEUT|17|14|cum ingressus fueris terram quam Dominus Deus tuus dabit tibi et possederis eam habitaverisque in illa et dixeris constituam super me regem sicut habent omnes per circuitum nationes
DEUT|17|15|eum constitues quem Dominus Deus tuus elegerit de numero fratrum tuorum non poteris alterius gentis hominem regem facere qui non sit frater tuus
DEUT|17|16|cumque fuerit constitutus non multiplicabit sibi equos nec reducet populum in Aegyptum equitatus numero sublevatus praesertim cum Dominus praeceperit vobis ut nequaquam amplius per eandem viam revertamini
DEUT|17|17|non habebit uxores plurimas quae inliciant animum eius neque argenti et auri inmensa pondera
DEUT|17|18|postquam autem sederit in solio regni sui describet sibi deuteronomium legis huius in volumine accipiens exemplar a sacerdotibus leviticae tribus
DEUT|17|19|et habebit secum legetque illud omnibus diebus vitae suae ut discat timere Dominum Deum suum et custodire verba et caerimonias eius quae lege praecepta sunt
DEUT|17|20|nec elevetur cor eius in superbiam super fratres suos neque declinet in partem dextram vel sinistram ut longo tempore regnet ipse et filii eius super Israhel
DEUT|18|1|non habebunt sacerdotes et Levitae et omnes qui de eadem tribu sunt partem et hereditatem cum reliquo Israhel quia sacrificia Domini et oblationes eius comedent
DEUT|18|2|et nihil aliud accipient de possessione fratrum suorum Dominus enim ipse est hereditas eorum sicut locutus est illis
DEUT|18|3|hoc erit iudicium sacerdotum a populo et ab his qui offerunt victimas sive bovem sive ovem immolaverint dabunt sacerdoti armum ac ventriculum
DEUT|18|4|primitias frumenti vini et olei et lanarum partem ex ovium tonsione
DEUT|18|5|ipsum enim elegit Dominus Deus tuus de cunctis tribubus tuis ut stet et ministret nomini Domini ipse et filii eius in sempiternum
DEUT|18|6|si exierit Levites de una urbium tuarum ex omni Israhel in qua habitat et voluerit venire desiderans locum quem elegerit Dominus
DEUT|18|7|ministrabit in nomine Dei sui sicut omnes fratres eius Levitae qui stabunt eo tempore coram Domino
DEUT|18|8|partem ciborum eandem accipiet quam et ceteri excepto eo quod in urbe sua ex paterna ei successione debetur
DEUT|18|9|quando ingressus fueris terram quam Dominus Deus tuus dabit tibi cave ne imitari velis abominationes illarum gentium
DEUT|18|10|nec inveniatur in te qui lustret filium suum aut filiam ducens per ignem aut qui ariolos sciscitetur et observet somnia atque auguria ne sit maleficus
DEUT|18|11|ne incantator ne pythones consulat ne divinos et quaerat a mortuis veritatem
DEUT|18|12|omnia enim haec abominatur Dominus et propter istiusmodi scelera delebit eos in introitu tuo
DEUT|18|13|perfectus eris et absque macula cum Domino Deo tuo
DEUT|18|14|gentes istae quarum possidebis terram augures et divinos audiunt tu autem a Domino Deo tuo aliter institutus es
DEUT|18|15|prophetam de gente tua et de fratribus tuis sicut me suscitabit tibi Dominus Deus tuus ipsum audies
DEUT|18|16|ut petisti a Domino Deo tuo in Horeb quando contio congregata est atque dixisti ultra non audiam vocem Domini Dei mei et ignem hunc maximum amplius non videbo ne moriar
DEUT|18|17|et ait Dominus mihi bene omnia sunt locuti
DEUT|18|18|prophetam suscitabo eis de medio fratrum suorum similem tui et ponam verba mea in ore eius loqueturque ad eos omnia quae praecepero illi
DEUT|18|19|qui autem verba eius quae loquetur in nomine meo audire noluerit ego ultor existam
DEUT|18|20|propheta autem qui arrogantia depravatus voluerit loqui in nomine meo quae ego non praecepi illi ut diceret aut ex nomine alienorum deorum interficietur
DEUT|18|21|quod si tacita cogitatione responderis quomodo possum intellegere verbum quod non est locutus Dominus
DEUT|18|22|hoc habebis signum quod in nomine Domini propheta ille praedixerit et non evenerit hoc Dominus non locutus est sed per tumorem animi sui propheta confinxit et idcirco non timebis eum
DEUT|19|1|cum disperderit Dominus Deus tuus gentes quarum tibi traditurus est terram et possederis eam habitaverisque in urbibus eius et in aedibus
DEUT|19|2|tres civitates separabis tibi in medio terrae quam Dominus Deus tuus dabit tibi in possessionem
DEUT|19|3|sternens diligenter viam et in tres aequaliter partes totam terrae tuae provinciam divides ut habeat e vicino qui propter homicidium profugus est quo possit evadere
DEUT|19|4|haec erit lex homicidae fugientis cuius vita servanda est qui percusserit proximum suum nesciens et qui heri et nudius tertius nullum contra eum habuisse odium conprobatur
DEUT|19|5|sed abisse simpliciter cum eo in silvam ad ligna caedenda et in succisione lignorum securis fugerit manu ferrumque lapsum de manubrio amicum eius percusserit et occiderit hic ad unam supradictarum urbium confugiet et vivet
DEUT|19|6|ne forsitan proximus eius cuius effusus est sanguis dolore stimulatus persequatur et adprehendat eum si longior via fuerit et percutiat animam eius qui non est reus mortis quia nullum contra eum qui occisus est odium prius habuisse monstratur
DEUT|19|7|idcirco praecipio tibi ut tres civitates aequalis inter se spatii dividas
DEUT|19|8|cum autem dilataverit Dominus Deus tuus terminos tuos sicut iuravit patribus tuis et dederit tibi cunctam terram quam eis pollicitus est
DEUT|19|9|si tamen custodieris mandata eius et feceris quae hodie praecipio tibi ut diligas Dominum Deum tuum et ambules in viis eius omni tempore addes tibi tres alias civitates et supradictarum trium urbium numerum duplicabis
DEUT|19|10|ut non effundatur sanguis innoxius in medio terrae quam Dominus Deus tuus dabit tibi possidendam nec sis sanguinis reus
DEUT|19|11|si quis autem odio habens proximum suum insidiatus fuerit vitae eius surgensque percusserit illum et mortuus fuerit fugeritque ad unam de supradictis urbibus
DEUT|19|12|mittent seniores civitatis illius et arripient eum de loco effugii tradentque in manu proximi cuius sanguis effusus est et morietur
DEUT|19|13|nec misereberis eius et auferes innoxium sanguinem de Israhel ut bene sit tibi
DEUT|19|14|non adsumes et transferes terminos proximi tui quos fixerunt priores in possessione tua quam Dominus Deus tuus dabit tibi in terra quam acceperis possidendam
DEUT|19|15|non stabit testis unus contra aliquem quicquid illud peccati et facinoris fuerit sed in ore duorum aut trium testium stabit omne verbum
DEUT|19|16|si steterit testis mendax contra hominem accusans eum praevaricationis
DEUT|19|17|stabunt ambo quorum causa est ante Dominum in conspectu sacerdotum et iudicum qui fuerint in diebus illis
DEUT|19|18|cumque diligentissime perscrutantes invenerint falsum testem dixisse contra fratrem suum mendacium
DEUT|19|19|reddent ei sicut fratri suo facere cogitavit et auferes malum de medio tui
DEUT|19|20|ut audientes ceteri timorem habeant et nequaquam talia audeant facere
DEUT|19|21|non misereberis eius sed animam pro anima oculum pro oculo dentem pro dente manum pro manu pedem pro pede exiges
DEUT|20|1|si exieris ad bellum contra hostes tuos et videris equitatum et currus et maiorem quam tu habes adversarii exercitus multitudinem non timebis eos quia Dominus Deus tuus tecum est qui eduxit te de terra Aegypti
DEUT|20|2|adpropinquante autem iam proelio stabit sacerdos ante aciem et sic loquetur ad populum
DEUT|20|3|audi Israhel vos hodie contra inimicos vestros pugnam committitis non pertimescat cor vestrum nolite metuere nolite cedere nec formidetis eos
DEUT|20|4|quia Dominus Deus vester in medio vestri est et pro vobis contra adversarios dimicabit ut eruat vos de periculo
DEUT|20|5|duces quoque per singulas turmas audiente exercitu proclamabunt quis est homo qui aedificavit domum novam et non dedicavit eam vadat et revertatur in domum suam ne forte moriatur in bello et alius dedicet illam
DEUT|20|6|quis est homo qui plantavit vineam et necdum eam fecit esse communem et de qua vesci omnibus liceat vadat et revertatur in domum suam ne forte moriatur in bello et alius homo eius fungatur officio
DEUT|20|7|quis est homo qui despondit uxorem et non accepit eam vadat et revertatur in domum suam ne forte moriatur in bello et alius homo accipiat eam
DEUT|20|8|his dictis addent reliqua et loquentur ad populum quis est homo formidolosus et corde pavido vadat et revertatur in domum suam ne pavere faciat corda fratrum suorum sicut ipse timore perterritus est
DEUT|20|9|cumque siluerint exercitus duces et finem loquendi fecerint unusquisque suos ad bellandum cuneos praeparabit
DEUT|20|10|si quando accesseris ad expugnandam civitatem offeres ei primum pacem
DEUT|20|11|si receperit et aperuerit tibi portas cunctus populus qui in ea est salvabitur et serviet tibi sub tributo
DEUT|20|12|sin autem foedus inire noluerint et receperint contra te bellum obpugnabis eam
DEUT|20|13|cumque tradiderit Dominus Deus tuus illam in manu tua percuties omne quod in ea generis masculini est in ore gladii
DEUT|20|14|absque mulieribus et infantibus iumentis et ceteris quae in civitate sunt omnem praedam exercitui divides et comedes de spoliis hostium tuorum quae Dominus Deus tuus dederit tibi
DEUT|20|15|sic facies cunctis civitatibus quae a te procul valde sunt et non sunt de his urbibus quas in possessionem accepturus es
DEUT|20|16|de his autem civitatibus quae dabuntur tibi nullum omnino permittes vivere
DEUT|20|17|sed interficies in ore gladii Hettheum videlicet et Amorreum et Chananeum Ferezeum et Eveum et Iebuseum sicut praecepit tibi Dominus Deus tuus
DEUT|20|18|ne forte doceant vos facere cunctas abominationes quas ipsi operati sunt diis suis et peccetis in Dominum Deum vestrum
DEUT|20|19|quando obsederis civitatem multo tempore et munitionibus circumdederis ut expugnes eam non succides arbores de quibus vesci potest nec securibus per circuitum debes vastare regionem quoniam lignum est et non homo nec potest bellantium contra te augere numerum
DEUT|20|20|si qua autem ligna non sunt pomifera sed agrestia et in ceteros apta usus succide et extrue machinas donec capias civitatem quae contra te dimicat
DEUT|21|1|quando inventum fuerit in terra quam Dominus Deus tuus daturus est tibi hominis cadaver occisi et ignoratur caedis reus
DEUT|21|2|egredientur maiores natu et iudices tui et metientur a loco cadaveris singularum per circuitum spatia civitatum
DEUT|21|3|et quam viciniorem ceteris esse perspexerint seniores civitatis eius tollent vitulam de armento quae non traxit iugum nec terram scidit vomere
DEUT|21|4|et ducent eam ad vallem asperam atque saxosam quae numquam arata est nec sementem recepit et caedent in ea cervices vitulae
DEUT|21|5|accedentque sacerdotes filii Levi quos elegerit Dominus Deus tuus ut ministrent ei et benedicant in nomine eius et ad verbum eorum omne negotium et quicquid mundum vel inmundum est iudicetur
DEUT|21|6|et maiores natu civitatis illius ad interfectum lavabuntque manus suas super vitulam quae in valle percussa est
DEUT|21|7|et dicent manus nostrae non effuderunt hunc sanguinem nec oculi viderunt
DEUT|21|8|propitius esto populo tuo Israhel quem redemisti Domine et non reputes sanguinem innocentem in medio populi tui Israhel et auferetur ab eis reatus sanguinis
DEUT|21|9|tu autem alienus eris ab innocentis cruore qui fusus est cum feceris quod praecepit Dominus
DEUT|21|10|si egressus fueris ad pugnam contra inimicos tuos et tradiderit eos Dominus Deus tuus in manu tua captivosque duxeris
DEUT|21|11|et videris in numero captivorum mulierem pulchram et adamaveris eam voluerisque habere uxorem
DEUT|21|12|introduces in domum tuam quae radet caesariem et circumcidet ungues
DEUT|21|13|et deponet vestem in qua capta est sedensque in domo tua flebit patrem et matrem suam uno mense et postea intrabis ad eam dormiesque cum illa et erit uxor tua
DEUT|21|14|sin autem postea non sederit animo tuo dimittes eam liberam nec vendere poteris pecunia nec opprimere per potentiam quia humiliasti eam
DEUT|21|15|si habuerit homo uxores duas unam dilectam et alteram odiosam genuerintque ex eo liberos et fuerit filius odiosae primogenitus
DEUT|21|16|volueritque substantiam inter filios suos dividere non poterit filium dilectae facere primogenitum et praeferre filio odiosae
DEUT|21|17|sed filium odiosae agnoscet primogenitum dabitque ei de his quae habuerit cuncta duplicia iste est enim principium liberorum eius et huic debentur primogenita
DEUT|21|18|si genuerit homo filium contumacem et protervum qui non audiat patris aut matris imperium et coercitus oboedire contempserit
DEUT|21|19|adprehendent eum et ducent ad seniores civitatis illius et ad portam iudicii
DEUT|21|20|dicentque ad eos filius noster iste protervus et contumax est monita nostra audire contemnit comesationibus vacat et luxuriae atque conviviis
DEUT|21|21|lapidibus eum obruet populus civitatis et morietur ut auferatis malum de medio vestri et universus Israhel audiens pertimescat
DEUT|21|22|quando peccaverit homo quod morte plectendum est et adiudicatus morti adpensus fuerit in patibulo
DEUT|21|23|non permanebit cadaver eius in ligno sed in eadem die sepelietur quia maledictus a Deo est qui pendet in ligno et nequaquam contaminabis terram tuam quam Dominus Deus tuus dederit tibi in possessionem
DEUT|22|1|non videbis bovem fratris tui aut ovem errantem et praeteribis sed reduces fratri tuo
DEUT|22|2|etiam si non est propinquus tuus frater nec nosti eum duces in domum tuam et erunt apud te quamdiu quaerat ea frater tuus et recipiat
DEUT|22|3|similiter facies de asino et de vestimento et de omni re fratris tui quae perierit si inveneris eam ne neglegas quasi alienam
DEUT|22|4|si videris asinum fratris tui aut bovem cecidisse in via non despicies sed sublevabis cum eo
DEUT|22|5|non induetur mulier veste virili nec vir utetur veste feminea abominabilis enim apud Deum est qui facit haec
DEUT|22|6|si ambulans per viam in arbore vel in terra nidum avis inveneris et matrem pullis vel ovis desuper incubantem non tenebis eam cum filiis
DEUT|22|7|sed abire patieris captos tenens filios ut bene sit tibi et longo vivas tempore
DEUT|22|8|cum aedificaveris domum novam facies murum tecti per circuitum ne effundatur sanguis in domo tua et sis reus labente alio et in praeceps ruente
DEUT|22|9|non seres vineam tuam altero semine ne et sementis quam sevisti et quae nascuntur ex vinea pariter sanctificentur
DEUT|22|10|non arabis in bove simul et asino
DEUT|22|11|non indueris vestimento quod ex lana linoque contextum est
DEUT|22|12|funiculos in fimbriis facies per quattuor angulos pallii tui quo operieris
DEUT|22|13|si duxerit vir uxorem et postea eam odio habuerit
DEUT|22|14|quaesieritque occasiones quibus dimittat eam obiciens ei nomen pessimum et dixerit uxorem hanc accepi et ingressus ad eam non inveni virginem
DEUT|22|15|tollent eam pater et mater eius et ferent secum signa virginitatis eius ad seniores urbis qui in porta sunt
DEUT|22|16|et dicet pater filiam meam dedi huic uxorem quam quia odit
DEUT|22|17|inponet ei nomen pessimum ut dicat non inveni filiam tuam virginem et ecce haec sunt signa virginitatis filiae meae expandent vestimentum coram senibus civitatis
DEUT|22|18|adprehendentque senes urbis illius virum et verberabunt illum
DEUT|22|19|condemnantes insuper centum siclis argenti quos dabit patri puellae quoniam diffamavit nomen pessimum super virginem Israhel habebitque eam uxorem et non poterit dimittere omni tempore vitae suae
DEUT|22|20|quod si verum est quod obicit et non est in puella inventa virginitas
DEUT|22|21|eicient eam extra fores domus patris sui et lapidibus obruent viri civitatis eius et morietur quoniam fecit nefas in Israhel ut fornicaretur in domo patris sui et auferes malum de medio tui
DEUT|22|22|si dormierit vir cum uxore alterius uterque morientur id est adulter et adultera et auferes malum de Israhel
DEUT|22|23|si puellam virginem desponderit vir et invenerit eam aliquis in civitate et concubuerit cum illa
DEUT|22|24|educes utrumque ad portam civitatis illius et lapidibus obruentur puella quia non clamavit cum esset in civitate vir quia humiliavit uxorem proximi sui et auferes malum de medio tui
DEUT|22|25|sin autem in agro reppererit vir puellam quae desponsata est et adprehendens concubuerit cum illa ipse morietur solus
DEUT|22|26|puella nihil patietur nec est rea mortis quoniam sicut latro consurgit contra fratrem suum et occidit animam eius ita et puella perpessa est
DEUT|22|27|sola erat in agro clamavit et nullus adfuit qui liberaret eam
DEUT|22|28|si invenerit vir puellam virginem quae non habet sponsum et adprehendens concubuerit cum ea et res ad iudicium venerit
DEUT|22|29|dabit qui dormivit cum ea patri puellae quinquaginta siclos argenti et habebit eam uxorem quia humiliavit illam non poterit dimittere cunctis diebus vitae suae
DEUT|22|30|non accipiet homo uxorem patris sui nec revelabit operimentum eius
DEUT|23|1|non intrabit eunuchus adtritis vel amputatis testiculis et absciso veretro ecclesiam Domini
DEUT|23|2|non ingredietur mamzer hoc est de scorto natus in ecclesiam Domini usque ad decimam generationem
DEUT|23|3|Ammanites et Moabites etiam post decimam generationem non intrabunt ecclesiam Domini in aeternum
DEUT|23|4|quia noluerunt vobis occurrere cum pane et aqua in via quando egressi estis de Aegypto et quia conduxerunt contra te Balaam filium Beor de Mesopotamiam Syriae ut malediceret tibi
DEUT|23|5|et noluit Dominus Deus tuus audire Balaam vertitque maledictionem eius in benedictionem tuam eo quod diligeret te
DEUT|23|6|non facies cum eis pacem nec quaeres eis bona cunctis diebus vitae tuae in sempiternum
DEUT|23|7|non abominaberis Idumeum quia frater tuus est nec Aegyptium quia advena fuisti in terra eius
DEUT|23|8|qui nati fuerint ex eis tertia generatione intrabunt ecclesiam Domini
DEUT|23|9|quando egressus fueris adversus hostes tuos in pugnam custodies te ab omni re mala
DEUT|23|10|si fuerit inter vos homo qui nocturno pollutus sit somnio egredietur extra castra
DEUT|23|11|et non revertetur priusquam ad vesperam lavetur aqua et post solis occasum regredietur in castra
DEUT|23|12|habebis locum extra castra ad quem egrediaris ad requisita naturae
DEUT|23|13|gerens paxillum in balteo cumque sederis fodies per circuitum et egesta humo operies
DEUT|23|14|quo relevatus es Dominus enim Deus tuus ambulat in medio castrorum ut eruat te et tradat tibi inimicos tuos ut sint castra tua sancta et nihil in eis appareat foeditatis nec derelinquat te
DEUT|23|15|non trades servum domino suo qui ad te confugerit
DEUT|23|16|habitabit tecum in loco qui ei placuerit et in una urbium tuarum requiescet nec contristes eum
DEUT|23|17|non erit meretrix de filiabus Israhel neque scortator de filiis Israhel
DEUT|23|18|non offeres mercedem prostibuli nec pretium canis in domum Domini Dei tui quicquid illud est quod voverint quia abominatio est utrumque apud Dominum Deum tuum
DEUT|23|19|non fenerabis fratri tuo ad usuram pecuniam nec fruges nec quamlibet aliam rem
DEUT|23|20|sed alieno fratri autem tuo absque usura id quod indiget commodabis ut benedicat tibi Dominus Deus tuus in omni opere tuo in terra ad quam ingredieris possidendam
DEUT|23|21|cum voveris votum Domino Deo tuo non tardabis reddere quia requiret illud Dominus Deus tuus et si moratus fueris reputabit tibi in peccatum
DEUT|23|22|si nolueris polliceri absque peccato eris
DEUT|23|23|quod autem semel egressum est de labiis tuis observabis et facies sicut promisisti Domino Deo tuo et propria voluntate et ore tuo locutus es
DEUT|23|24|ingressus vineam proximi tui comede uvas quantum tibi placuerit foras autem ne efferas tecum
DEUT|23|25|si intraveris in segetem amici tui franges spicas et manu conteres falce autem non metes
DEUT|24|1|si acceperit homo uxorem et habuerit eam et non invenerit gratiam ante oculos eius propter aliquam foeditatem scribet libellum repudii et dabit in manu illius et dimittet eam de domo sua
DEUT|24|2|cumque egressa alterum maritum duxerit
DEUT|24|3|et ille quoque oderit eam dederitque ei libellum repudii et dimiserit de domo sua vel certe mortuus fuerit
DEUT|24|4|non poterit prior maritus recipere eam in uxorem quia polluta est et abominabilis facta est coram Domino ne peccare facias terram tuam quam Dominus Deus tuus tibi tradiderit possidendam
DEUT|24|5|cum acceperit homo nuper uxorem non procedet ad bellum nec ei quippiam necessitatis iniungetur publicae sed vacabit absque culpa domui suae ut uno anno laetetur cum uxore sua
DEUT|24|6|non accipies loco pignoris inferiorem et superiorem molam quia animam suam adposuit tibi
DEUT|24|7|si deprehensus fuerit homo sollicitans fratrem suum de filiis Israhel et vendito eo accipiens pretium interficietur et auferes malum de medio tui
DEUT|24|8|observa diligenter ne incurras in plagam leprae sed facies quaecumque docuerint te sacerdotes levitici generis iuxta id quod praecepi eis et imple sollicite
DEUT|24|9|mementote quae fecerit Dominus Deus vester Mariae in via cum egrederemini de Aegypto
DEUT|24|10|cum repetes a proximo tuo rem aliquam quam debet tibi non ingredieris domum eius ut pignus auferas
DEUT|24|11|sed stabis foris et ille tibi proferet quod habuerit
DEUT|24|12|sin autem pauper est non pernoctabit apud te pignus
DEUT|24|13|sed statim reddes ei ante solis occasum ut dormiens in vestimento suo benedicat tibi et habeas iustitiam coram Domino Deo tuo
DEUT|24|14|non negabis mercedem indigentis et pauperis fratris tui sive advenae qui tecum moratur in terra et intra portas tuas est
DEUT|24|15|sed eadem die reddes ei pretium laboris sui ante solis occasum quia pauper est et ex eo sustentat animam suam ne clamet contra te ad Dominum et reputetur tibi in peccatum
DEUT|24|16|non occidentur patres pro filiis nec filii pro patribus sed unusquisque pro suo peccato morietur
DEUT|24|17|non pervertes iudicium advenae et pupilli nec auferes pignoris loco viduae vestimentum
DEUT|24|18|memento quod servieris in Aegypto et eruerit te Dominus Deus tuus inde idcirco praecipio tibi ut facias hanc rem
DEUT|24|19|quando messueris segetem in agro tuo et oblitus manipulum reliqueris non reverteris ut tollas eum sed advenam et pupillum et viduam auferre patieris ut benedicat tibi Dominus Deus tuus in omni opere manuum tuarum
DEUT|24|20|si fruges colliges olivarum quicquid remanserit in arboribus non reverteris ut colligas sed relinques advenae pupillo ac viduae
DEUT|24|21|si vindemiaveris vineam tuam non colliges remanentes racemos sed cedent in usus advenae pupilli ac viduae
DEUT|24|22|memento quod et tu servieris in Aegypto et idcirco praecipiam tibi ut facias hanc rem
DEUT|25|1|si fuerit causa inter aliquos et interpellaverint iudices quem iustum esse perspexerint illi iustitiae palmam dabunt quem impium condemnabunt impietatis
DEUT|25|2|sin autem eum qui peccavit dignum viderint plagis prosternent et coram se facient verberari pro mensura peccati erit et plagarum modus
DEUT|25|3|ita dumtaxat ut quadragenarium numerum non excedant ne foede laceratus ante oculos tuos abeat frater tuus
DEUT|25|4|non ligabis os bovis terentis in area fruges tuas
DEUT|25|5|quando habitaverint fratres simul et unus ex eis absque liberis mortuus fuerit uxor defuncti non nubet alteri sed accipiet eam frater eius et suscitabit semen fratris sui
DEUT|25|6|et primogenitum ex ea filium nomine illius appellabit ut non deleatur nomen eius ex Israhel
DEUT|25|7|sin autem noluerit accipere uxorem fratris sui quae ei lege debetur perget mulier ad portam civitatis et interpellabit maiores natu dicetque non vult frater viri mei suscitare nomen fratris sui in Israhel nec me in coniugium sumere
DEUT|25|8|statimque accersiri eum facient et interrogabunt si responderit nolo eam uxorem accipere
DEUT|25|9|accedet mulier ad eum coram senioribus et tollet calciamentum de pede eius spuetque in faciem illius et dicet sic fit homini qui non aedificat domum fratris sui
DEUT|25|10|et vocabitur nomen illius in Israhel domus Disculciati
DEUT|25|11|si habuerint inter se iurgium viri et unus contra alterum rixari coeperit volensque uxor alterius eruere virum suum de manu fortioris miserit manum et adprehenderit verenda eius
DEUT|25|12|abscides manum illius nec flecteris super eam ulla misericordia
DEUT|25|13|non habebis in sacculo diversa pondera maius et minus
DEUT|25|14|nec erit in domo tua modius maior et minor
DEUT|25|15|pondus habebis iustum et verum et modius aequalis et verus erit tibi ut multo vivas tempore super terram quam Dominus Deus tuus dederit tibi
DEUT|25|16|abominatur enim Dominus eum qui facit haec et aversatur omnem iniustitiam
DEUT|25|17|memento quae fecerit tibi Amalech in via quando egrediebaris ex Aegypto
DEUT|25|18|quomodo occurrerit tibi et extremos agminis tui qui lassi residebant ceciderit quando tu eras fame et labore confectus et non timuerit Deum
DEUT|25|19|cum ergo Dominus Deus tuus dederit tibi requiem et subiecerit cunctas per circuitum nationes in terra quam tibi pollicitus est delebis nomen eius sub caelo cave ne obliviscaris
DEUT|26|1|cumque intraveris terram quam Dominus Deus tuus tibi daturus est possidendam et obtinueris eam atque habitaveris in illa
DEUT|26|2|tolles de cunctis frugibus primitias et pones in cartallo pergesque ad locum quem Dominus Deus tuus elegerit ut ibi invocetur nomen eius
DEUT|26|3|accedesque ad sacerdotem qui fuerit in diebus illis et dices ad eum profiteor hodie coram Domino Deo tuo quod ingressus sim terram pro qua iuravit patribus nostris ut daret eam nobis
DEUT|26|4|suscipiensque sacerdos cartallum de manu eius ponet ante altare Domini Dei tui
DEUT|26|5|et loqueris in conspectu Domini Dei tui Syrus persequebatur patrem meum qui descendit in Aegyptum et ibi peregrinatus est in paucissimo numero crevitque in gentem magnam et robustam et infinitae multitudinis
DEUT|26|6|adflixeruntque nos Aegyptii et persecuti sunt inponentes onera gravissima
DEUT|26|7|et clamavimus ad Dominum Deum patrum nostrorum qui exaudivit nos et respexit humilitatem nostram et laborem atque angustias
DEUT|26|8|et eduxit nos de Aegypto in manu forti et brachio extento in ingenti pavore in signis atque portentis
DEUT|26|9|et introduxit ad locum istum et tradidit nobis terram lacte et melle manantem
DEUT|26|10|et idcirco nunc offero primitias frugum terrae quam dedit Dominus mihi et dimittes eas in conspectu Domini Dei tui adorato Domino Deo tuo
DEUT|26|11|et epulaberis in omnibus bonis quae Dominus Deus tuus dederit tibi et domui tuae tu et Levites et advena qui tecum est
DEUT|26|12|quando conpleveris decimam cunctarum frugum tuarum anno decimarum tertio dabis Levitae et advenae et pupillo et viduae ut comedant intra portas tuas et saturentur
DEUT|26|13|loquerisque in conspectu Domini Dei tui abstuli quod sanctificatum est de domo mea et dedi illud Levitae et advenae pupillo et viduae sicut iussisti mihi non praeterivi mandata tua nec sum oblitus imperii
DEUT|26|14|non comedi ex eis in luctu meo nec separavi ea in qualibet inmunditia nec expendi ex his quicquam in re funebri oboedivi voci Domini Dei mei et feci omnia sicut praecepisti mihi
DEUT|26|15|respice de sanctuario tuo de excelso caelorum habitaculo et benedic populo tuo Israhel et terrae quam dedisti nobis sicut iurasti patribus nostris terrae lacte et melle mananti
DEUT|26|16|hodie Dominus Deus tuus praecepit tibi ut facias mandata haec atque iudicia et custodias et impleas ex toto corde tuo et ex tota anima tua
DEUT|26|17|Dominum elegisti hodie ut sit tibi Deus et ambules in viis eius et custodias caerimonias illius et mandata atque iudicia et oboedias eius imperio
DEUT|26|18|et Dominus elegit te hodie ut sis ei populus peculiaris sicut locutus est tibi et custodias omnia praecepta eius
DEUT|26|19|et faciat te excelsiorem cunctis gentibus quas creavit in laudem et nomen et gloriam suam ut sis populus sanctus Domini Dei tui sicut locutus est
DEUT|27|1|praecepit autem Moses et seniores Israhel populo dicentes custodite omne mandatum quod praecipio vobis hodie
DEUT|27|2|cumque transieritis Iordanem in terram quam Dominus Deus tuus dabit tibi eriges ingentes lapides et calce levigabis eos
DEUT|27|3|ut possis in eis scribere omnia verba legis huius Iordane transmisso ut introeas terram quam Dominus Deus tuus dabit tibi terram lacte et melle manantem sicut iuravit patribus tuis
DEUT|27|4|quando ergo transieritis Iordanem erige lapides quos ego hodie praecipio vobis in monte Hebal et levigabis calce
DEUT|27|5|et aedificabis ibi altare Domino Deo tuo de lapidibus quos ferrum non tetigit
DEUT|27|6|et de saxis informibus et inpolitis et offeres super eo holocausta Domino Deo tuo
DEUT|27|7|et immolabis hostias pacificas comedesque ibi et epulaberis coram Domino Deo tuo
DEUT|27|8|et scribes super lapides omnia verba legis huius plane et lucide
DEUT|27|9|dixeruntque Moses et sacerdotes levitici generis ad omnem Israhelem adtende et audi Israhel hodie factus es populus Domini Dei tui
DEUT|27|10|audies vocem eius et facies mandata atque iustitias quas ego praecipio tibi
DEUT|27|11|praecepitque Moses populo in die illo dicens
DEUT|27|12|hii stabunt ad benedicendum Domino super montem Garizim Iordane transmisso Symeon Levi Iudas Isachar Ioseph et Beniamin
DEUT|27|13|et e regione isti stabunt ad maledicendum in monte Hebal Ruben Gad et Aser Zabulon Dan et Nepthalim
DEUT|27|14|et pronuntiabunt Levitae dicentque ad omnes viros Israhel excelsa voce
DEUT|27|15|maledictus homo qui facit sculptile et conflatile abominationem Domini opus manuum artificum ponetque illud in abscondito et respondebit omnis populus et dicet amen
DEUT|27|16|maledictus qui non honorat patrem suum et matrem et dicet omnis populus amen
DEUT|27|17|maledictus qui transfert terminos proximi sui et dicet omnis populus amen
DEUT|27|18|maledictus qui errare facit caecum in itinere et dicet omnis populus amen
DEUT|27|19|maledictus qui pervertit iudicium advenae pupilli et viduae et dicet omnis populus amen
DEUT|27|20|maledictus qui dormit cum uxore patris sui et revelat operimentum lectuli eius et dicet omnis populus amen
DEUT|27|21|maledictus qui dormit cum omni iumento et dicet omnis populus amen
DEUT|27|22|maledictus qui dormit cum sorore sua filia patris sui sive matris suae et dicet omnis populus amen
DEUT|27|23|maledictus qui dormit cum socru sua et dicet omnis populus amen
DEUT|27|24|maledictus qui clam percusserit proximum suum et dicet omnis populus amen
DEUT|27|25|maledictus qui accipit munera ut percutiat animam sanguinis innocentis et dicet omnis populus amen
DEUT|27|26|maledictus qui non permanet in sermonibus legis huius nec eos opere perficit et dicet omnis populus amen
DEUT|28|1|sin autem audieris vocem Domini Dei tui ut facias atque custodias omnia mandata eius quae ego praecipio tibi hodie faciet te Dominus Deus tuus excelsiorem cunctis gentibus quae versantur in terra
DEUT|28|2|venientque super te universae benedictiones istae et adprehendent te si tamen praecepta eius audieris
DEUT|28|3|benedictus tu in civitate et benedictus in agro
DEUT|28|4|benedictus fructus ventris tui et fructus terrae tuae fructusque iumentorum tuorum greges armentorum et caulae ovium tuarum
DEUT|28|5|benedicta horrea tua et benedictae reliquiae tuae
DEUT|28|6|benedictus eris et ingrediens et egrediens
DEUT|28|7|dabit Dominus inimicos tuos qui consurgunt adversum te corruentes in conspectu tuo per unam viam venient contra te et per septem fugient a facie tua
DEUT|28|8|emittet Dominus benedictionem super cellaria tua et super omnia opera manuum tuarum benedicetque tibi in terra quam acceperis
DEUT|28|9|suscitabit te Dominus sibi in populum sanctum sicut iuravit tibi si custodieris mandata Domini Dei tui et ambulaveris in viis eius
DEUT|28|10|videbuntque omnes terrarum populi quod nomen Domini invocatum sit super te et timebunt te
DEUT|28|11|abundare te faciet Dominus omnibus bonis fructu uteri tui et fructu iumentorum tuorum fructu terrae tuae quam iuravit Dominus patribus tuis ut daret tibi
DEUT|28|12|aperiet Dominus thesaurum suum optimum caelum ut tribuat pluviam terrae tuae in tempore suo benedicet cunctis operibus manuum tuarum et fenerabis gentibus multis et ipse a nullo fenus accipies
DEUT|28|13|constituet te Dominus in caput et non in caudam et eris semper supra et non subter si audieris mandata Domini Dei tui quae ego praecipio tibi hodie et custodieris et feceris
DEUT|28|14|ac non declinaveris ab eis nec ad dextram nec ad sinistram nec secutus fueris deos alienos neque colueris eos
DEUT|28|15|quod si audire nolueris vocem Domini Dei tui ut custodias et facias omnia mandata eius et caerimonias quas ego praecipio tibi hodie venient super te omnes maledictiones istae et adprehendent te
DEUT|28|16|maledictus eris in civitate maledictus in agro
DEUT|28|17|maledictum horreum tuum et maledictae reliquiae tuae
DEUT|28|18|maledictus fructus ventris tui et fructus terrae tuae armenta boum tuorum et greges ovium tuarum
DEUT|28|19|maledictus eris ingrediens et maledictus egrediens
DEUT|28|20|mittet Dominus super te famem et esuriem et increpationem in omnia opera tua quae facies donec conterat te et perdat velociter propter adinventiones tuas pessimas in quibus reliquisti me
DEUT|28|21|adiungat Dominus tibi pestilentiam donec consumat te de terra ad quam ingredieris possidendam
DEUT|28|22|percutiat te Dominus egestate febri et frigore ardore et aestu et aere corrupto ac robigine et persequatur donec pereas
DEUT|28|23|sit caelum quod supra te est aeneum et terra quam calcas ferrea
DEUT|28|24|det Dominus imbrem terrae tuae pulverem et de caelo descendat super te cinis donec conteraris
DEUT|28|25|tradat te Dominus corruentem ante hostes tuos per unam viam egrediaris contra eos et per septem fugias et dispergaris per omnia regna terrae
DEUT|28|26|sitque cadaver tuum in escam cunctis volatilibus caeli et bestiis terrae et non sit qui abigat
DEUT|28|27|percutiat te Dominus ulcere Aegypti et parte corporis per quam stercora digeruntur scabie quoque et prurigine ita ut curari nequeas
DEUT|28|28|percutiat te Dominus amentia et caecitate ac furore mentis
DEUT|28|29|et palpes in meridie sicut palpare solet caecus in tenebris et non dirigas vias tuas omnique tempore calumniam sustineas et opprimaris violentia nec habeas qui liberet te
DEUT|28|30|uxorem accipias et alius dormiat cum ea domum aedifices et non habites in ea plantes vineam et non vindemies eam
DEUT|28|31|bos tuus immoletur coram te et non comedas ex eo asinus tuus rapiatur in conspectu tuo et non reddatur tibi oves tuae dentur inimicis tuis et non sit qui te adiuvet
DEUT|28|32|filii tui et filiae tuae tradantur alteri populo videntibus oculis tuis et deficientibus ad conspectum eorum tota die et non sit fortitudo in manu tua
DEUT|28|33|fructus terrae tuae et omnes labores tuos comedat populus quem ignoras et sis semper calumniam sustinens et oppressus cunctis diebus
DEUT|28|34|et stupens ad terrorem eorum quae videbunt oculi tui
DEUT|28|35|percutiat te Dominus ulcere pessimo in genibus et in suris sanarique non possis a planta pedis usque ad verticem tuum
DEUT|28|36|ducet Dominus te et regem tuum quem constitueris super te in gentem quam ignoras tu et patres tui et servies ibi diis alienis ligno et lapidi
DEUT|28|37|et eris perditus in proverbium ac fabulam omnibus populis ad quos te introduxerit Dominus
DEUT|28|38|sementem multam iacies in terram et modicum congregabis quia lucustae omnia devorabunt
DEUT|28|39|vineam plantabis et fodies et vinum non bibes nec colliges ex ea quippiam quoniam vastabitur vermibus
DEUT|28|40|olivas habebis in omnibus terminis tuis et non ungueris oleo quia defluent et peribunt
DEUT|28|41|filios generabis et filias et non frueris eis quoniam ducentur in captivitatem
DEUT|28|42|omnes arbores tuas et fruges terrae tuae robigo consumet
DEUT|28|43|advena qui tecum versatur in terra ascendet super te eritque sublimior tu autem descendes et eris inferior
DEUT|28|44|ipse fenerabit tibi et tu non fenerabis ei ipse erit in caput et tu eris in caudam
DEUT|28|45|et venient super te omnes maledictiones istae et persequentes adprehendent te donec intereas quia non audisti vocem Domini Dei tui nec servasti mandata eius et caerimonias quas praecepit tibi
DEUT|28|46|et erunt in te signa atque prodigia et in semine tuo usque in sempiternum
DEUT|28|47|eo quod non servieris Domino Deo tuo in gaudio cordisque laetitia propter rerum omnium abundantiam
DEUT|28|48|servies inimico tuo quem inmittet Dominus tibi in fame et siti et nuditate et omnium penuria et ponet iugum ferreum super cervicem tuam donec te conterat
DEUT|28|49|adducet Dominus super te gentem de longinquo et de extremis finibus terrae in similitudinem aquilae volantis cum impetu cuius linguam intellegere non possis
DEUT|28|50|gentem procacissimam quae non deferat seni nec misereatur parvulo
DEUT|28|51|et devoret fructum iumentorum tuorum ac fruges terrae tuae donec intereas et non relinquat tibi triticum vinum et oleum armenta boum et greges ovium donec te disperdat
DEUT|28|52|et conterat in cunctis urbibus tuis et destruantur muri tui firmi atque sublimes in quibus habebas fiduciam in omni terra tua obsideberis intra portas tuas in omni terra quam dabit tibi Dominus Deus tuus
DEUT|28|53|et comedes fructum uteri tui et carnes filiorum et filiarum tuarum quas dedit tibi Dominus Deus tuus in angustia et vastitate qua opprimet te hostis tuus
DEUT|28|54|homo delicatus in te et luxuriosus valde invidebit fratri suo et uxori quae cubat in sinu suo
DEUT|28|55|ne det eis de carnibus filiorum suorum quas comedet eo quod nihil habeat aliud in obsidione et penuria qua vastaverint te inimici tui intra omnes portas tuas
DEUT|28|56|tenera mulier et delicata quae super terram ingredi non valebat nec pedis vestigium figere propter mollitiem et teneritudinem nimiam invidebit viro suo qui cubat in sinu eius super filii et filiae carnibus
DEUT|28|57|et inluvie secundarum quae egrediuntur de medio feminum eius et super liberis qui eadem hora nati sunt comedent enim eos clam propter rerum omnium penuriam in obsidione et vastitate qua opprimet te inimicus tuus intra portas tuas
DEUT|28|58|nisi custodieris et feceris omnia verba legis huius quae scripta sunt in hoc volumine et timueris nomen eius gloriosum et terribile hoc est Dominum Deum tuum
DEUT|28|59|augebit Dominus plagas tuas et plagas seminis tui plagas magnas et perseverantes infirmitates pessimas et perpetuas
DEUT|28|60|et convertet in te omnes adflictiones Aegypti quas timuisti et adherebunt tibi
DEUT|28|61|insuper et universos languores et plagas quae non sunt scriptae in volumine legis huius inducet Dominus super te donec te conterat
DEUT|28|62|et remanebitis pauci numero qui prius eratis sicut astra caeli prae multitudine quoniam non audisti vocem Domini Dei tui
DEUT|28|63|et sicut ante laetatus est Dominus super vos bene vobis faciens vosque multiplicans sic laetabitur disperdens vos atque subvertens ut auferamini de terra ad quam ingredieris possidendam
DEUT|28|64|disperget te Dominus in omnes populos a summitate terrae usque ad terminos eius et servies ibi diis alienis quos et tu ignoras et patres tui lignis et lapidibus
DEUT|28|65|in gentibus quoque illis non quiesces neque erit requies vestigio pedis tui dabit enim tibi Dominus ibi cor pavidum et deficientes oculos et animam maerore consumptam
DEUT|28|66|et erit vita tua quasi pendens ante te timebis nocte et die et non credes vitae tuae
DEUT|28|67|mane dices quis mihi det vesperum et vespere quis mihi det mane propter cordis tui formidinem qua terreberis et propter ea quae tuis videbis oculis
DEUT|28|68|reducet te Dominus classibus in Aegyptum per viam de qua dixi tibi ut eam amplius non videres ibi venderis inimicis tuis in servos et ancillas et non erit qui emat
DEUT|29|1|haec sunt verba foederis quod praecepit Dominus Mosi ut feriret cum filiis Israhel in terra Moab praeter illud foedus quod cum eis pepigit in Horeb
DEUT|29|2|vocavitque Moses omnem Israhelem et dixit ad eos vos vidistis universa quae fecit Dominus coram vobis in terra Aegypti Pharaoni et omnibus servis eius universaeque terrae illius
DEUT|29|3|temptationes magnas quas viderunt oculi tui signa illa portentaque ingentia
DEUT|29|4|et non dedit Dominus vobis cor intellegens et oculos videntes et aures quae possint audire usque in praesentem diem
DEUT|29|5|adduxi vos quadraginta annis per desertum non sunt adtrita vestimenta vestra nec calciamenta pedum tuorum vetustate consumpta sunt
DEUT|29|6|panem non comedistis vinum et siceram non bibistis ut sciretis quia ego sum Dominus Deus vester
DEUT|29|7|et venistis ad locum hunc egressusque est Seon rex Esebon et Og rex Basan occurrens nobis ad pugnam et percussimus eos
DEUT|29|8|et tulimus terram eorum ac tradidimus possidendam Ruben et Gad et dimidiae tribui Manasse
DEUT|29|9|custodite ergo verba pacti huius et implete ea ut intellegatis universa quae facitis
DEUT|29|10|vos statis hodie cuncti coram Domino Deo vestro principes vestri ac tribus et maiores natu atque doctores omnis populus Israhel
DEUT|29|11|liberi et uxores vestrae et advena qui tecum moratur in castris exceptis lignorum caesoribus et his qui conportant aquas
DEUT|29|12|ut transeas in foedere Domini Dei tui et in iureiurando quod hodie Dominus Deus tuus percutit tecum
DEUT|29|13|ut suscitet te sibi in populum et ipse sit Deus tuus sicut locutus est tibi et sicut iuravit patribus tuis Abraham Isaac et Iacob
DEUT|29|14|nec vobis solis ego hoc foedus ferio et haec iuramenta confirmo
DEUT|29|15|sed cunctis praesentibus et absentibus
DEUT|29|16|vos enim nostis ut habitaverimus in terra Aegypti et quomodo transierimus per medium nationum quas transeuntes
DEUT|29|17|vidistis abominationes et sordes id est idola eorum lignum et lapidem argentum et aurum quae colebant
DEUT|29|18|ne forte sit inter vos vir aut mulier familia aut tribus cuius cor aversum est hodie a Domino Deo vestro ut vadat et serviat diis illarum gentium et sit inter vos radix germinans fel et amaritudinem
DEUT|29|19|cumque audierit verba iuramenti huius benedicat sibi in corde suo dicens pax erit mihi et ambulabo in pravitate cordis mei et adsumat ebria sitientem
DEUT|29|20|et Dominus non ignoscat ei sed tunc quam maxime furor eius fumet et zelus contra hominem illum et sedeant super eo omnia maledicta quae scripta sunt in hoc volumine et deleat nomen eius sub caelo
DEUT|29|21|et consumat eum in perditionem ex omnibus tribubus Israhel iuxta maledictiones quae in libro legis huius ac foederis continentur
DEUT|29|22|dicetque sequens generatio et filii qui nascentur deinceps et peregrini qui de longe venerint videntes plagas terrae illius et infirmitates quibus eam adflixerit Dominus
DEUT|29|23|sulphure et salis ardore conburens ita ut ultra non seratur nec virens quippiam germinet in exemplum subversionis Sodomae et Gomorrae Adamae et Seboim quas subvertit Dominus in ira et furore suo
DEUT|29|24|et dicent omnes gentes quare sic fecit Dominus terrae huic quae est haec ira furoris eius inmensa
DEUT|29|25|et respondebunt quia dereliquerunt pactum Domini quod pepigit cum patribus eorum quando eduxit eos de terra Aegypti
DEUT|29|26|et servierunt diis alienis et adoraverunt eos quos nesciebant et quibus non fuerant adtributi
DEUT|29|27|idcirco iratus est furor Domini contra terram istam ut induceret super eam omnia maledicta quae in hoc volumine scripta sunt
DEUT|29|28|et eiecit eos de terra sua in ira et furore et indignatione maxima proiecitque in terram alienam sicut hodie conprobatur
DEUT|29|29|abscondita Domino Deo nostro quae manifesta sunt nobis et filiis nostris usque in aeternum ut faciamus universa legis huius
DEUT|30|1|cum ergo venerint super te omnes sermones isti benedictio sive maledictio quam proposui in conspectu tuo et ductus paenitudine cordis tui in universis gentibus in quas disperserit te Dominus Deus tuus
DEUT|30|2|reversus fueris ad eum et oboedieris eius imperiis sicut ego hodie praecipio tibi cum filiis tuis in toto corde tuo et in tota anima tua
DEUT|30|3|reducet Dominus Deus tuus captivitatem tuam ac miserebitur tui et rursum congregabit te de cunctis populis in quos te ante dispersit
DEUT|30|4|si ad cardines caeli fueris dissipatus inde te retrahet Dominus Deus tuus
DEUT|30|5|et adsumet atque introducet in terram quam possederunt patres tui et obtinebis eam et benedicens tibi maioris numeri esse te faciet quam fuerunt patres tui
DEUT|30|6|circumcidet Dominus Deus tuus cor tuum et cor seminis tui ut diligas Dominum Deum tuum in toto corde tuo et in tota anima tua et possis vivere
DEUT|30|7|omnes autem maledictiones has convertet super inimicos tuos et eos qui oderunt te et persequuntur
DEUT|30|8|tu autem reverteris et audies vocem Domini Dei tui faciesque universa mandata quae ego praecipio tibi hodie
DEUT|30|9|et abundare te faciet Dominus Deus tuus in cunctis operibus manuum tuarum in subole uteri tui et in fructu iumentorum tuorum in ubertate terrae tuae et in rerum omnium largitate revertetur enim Dominus ut gaudeat super te in omnibus bonis sicut gavisus est in patribus tuis
DEUT|30|10|si tamen audieris vocem Domini Dei tui et custodieris praecepta eius et caerimonias quae in hac lege conscriptae sunt et revertaris ad Dominum Deum tuum in toto corde tuo et in tota anima tua
DEUT|30|11|mandatum hoc quod ego praecipio tibi hodie non supra te est neque procul positum
DEUT|30|12|nec in caelo situm ut possis dicere quis nostrum ad caelum valet conscendere ut deferat illud ad nos et audiamus atque opere conpleamus
DEUT|30|13|neque trans mare positum ut causeris et dicas quis e nobis transfretare poterit mare et illud ad nos usque deferre ut possimus audire et facere quod praeceptum est
DEUT|30|14|sed iuxta te est sermo valde in ore tuo et in corde tuo ut facias illum
DEUT|30|15|considera quod hodie proposuerim in conspectu tuo vitam et bonum et e contrario mortem et malum
DEUT|30|16|ut diligas Dominum Deum tuum et ambules in viis eius et custodias mandata illius et caerimonias atque iudicia et vivas ac multiplicet te benedicatque tibi in terra ad quam ingredieris possidendam
DEUT|30|17|sin autem aversum fuerit cor tuum et audire nolueris atque errore deceptus adoraveris deos alienos et servieris eis
DEUT|30|18|praedico tibi hodie quod pereas et parvo tempore moreris in terra ad quam Iordane transmisso ingredieris possidendam
DEUT|30|19|testes invoco hodie caelum et terram quod proposuerim vobis vitam et mortem bonum et malum benedictionem et maledictionem elige ergo vitam ut et tu vivas et semen tuum
DEUT|30|20|et diligas Dominum Deum tuum atque oboedias voci eius et illi adhereas ipse est enim vita tua et longitudo dierum tuorum ut habites in terra pro qua iuravit Dominus patribus tuis Abraham Isaac et Iacob ut daret eam illis
DEUT|31|1|abiit itaque Moses et locutus est omnia verba haec ad universum Israhel
DEUT|31|2|et dixit ad eos centum viginti annorum sum hodie non possum ultra egredi et ingredi praesertim cum et Dominus dixerit mihi non transibis Iordanem istum
DEUT|31|3|Dominus ergo Deus tuus transibit ante te ipse delebit omnes gentes has in conspectu tuo et possidebis eas et Iosue iste transibit ante te sicut locutus est Dominus
DEUT|31|4|facietque Dominus eis sicut fecit Seon et Og regibus Amorreorum et terrae eorum delebitque eos
DEUT|31|5|cum ergo et hos tradiderit vobis similiter facietis eis sicut praecepi vobis
DEUT|31|6|viriliter agite et confortamini nolite timere nec paveatis a conspectu eorum quia Dominus Deus tuus ipse est ductor tuus et non dimittet nec derelinquet te
DEUT|31|7|vocavitque Moses Iosue et dixit ei coram omni Israhel confortare et esto robustus tu enim introduces populum istum in terram quam daturum se patribus eorum iuravit Dominus et tu eam sorte divides
DEUT|31|8|et Dominus qui ductor vester est ipse erit tecum non dimittet nec derelinquet te noli timere nec paveas
DEUT|31|9|scripsit itaque Moses legem hanc et tradidit eam sacerdotibus filiis Levi qui portabant arcam foederis Domini et cunctis senioribus Israhelis
DEUT|31|10|praecepitque eis dicens post septem annos anno remissionis in sollemnitate tabernaculorum
DEUT|31|11|convenientibus cunctis ex Israhel ut appareant in conspectu Domini Dei tui in loco quem elegerit Dominus leges verba legis huius coram omni Israhel audientibus eis
DEUT|31|12|et in unum omni populo congregato tam viris quam mulieribus parvulis et advenis qui sunt intra portas tuas ut audientes discant et timeant Dominum Deum vestrum et custodiant impleantque omnes sermones legis huius
DEUT|31|13|filii quoque eorum qui nunc ignorant audire possint et timeant Dominum Deum suum cunctis diebus quibus versantur in terra ad quam vos Iordane transito pergitis obtinendam
DEUT|31|14|et ait Dominus ad Mosen ecce prope sunt dies mortis tuae voca Iosue et state in tabernaculo testimonii ut praecipiam ei abierunt ergo Moses et Iosue et steterunt in tabernaculo testimonii
DEUT|31|15|apparuitque Dominus ibi in columna nubis quae stetit in introitu tabernaculi
DEUT|31|16|dixitque Dominus ad Mosen ecce tu dormies cum patribus tuis et populus iste consurgens fornicabitur post deos alienos in terra ad quam ingredietur et habitabit in ea ibi derelinquet me et irritum faciet foedus quod pepigi cum eo
DEUT|31|17|et irascetur furor meus contra eum in die illo et derelinquam eum et abscondam faciem meam ab eo et erit in devorationem invenient eum omnia mala et adflictiones ita ut dicat in illo die vere quia non est Deus mecum invenerunt me haec mala
DEUT|31|18|ego autem abscondam et celabo faciem meam in die illo propter omnia mala quae fecit quia secutus est deos alienos
DEUT|31|19|nunc itaque scribite vobis canticum istud et docete filios Israhel ut memoriter teneant et ore decantent et sit mihi carmen istud pro testimonio inter filios Israhel
DEUT|31|20|introducam enim eum in terram pro qua iuravi patribus eius lacte et melle manantem cumque comederint et saturati crassique fuerint avertentur ad deos alienos et servient eis et detrahent mihi et irritum facient pactum meum
DEUT|31|21|postquam invenerint eum mala multa et adflictiones respondebit ei canticum istud pro testimonio quod nulla delebit oblivio ex ore seminis tui scio enim cogitationes eius quae facturus sit hodie antequam introducam eum in terram quam ei pollicitus sum
DEUT|31|22|scripsit ergo Moses canticum et docuit filios Israhel
DEUT|31|23|praecepitque Iosue filio Nun et ait confortare et esto robustus tu enim introduces filios Israhel in terram quam pollicitus sum et ego ero tecum
DEUT|31|24|postquam ergo scripsit Moses verba legis huius in volumine atque conplevit
DEUT|31|25|praecepit Levitis qui portabant arcam foederis Domini dicens
DEUT|31|26|tollite librum istum et ponite eum in latere arcae foederis Domini Dei vestri ut sit ibi contra te in testimonio
DEUT|31|27|ego enim scio contentionem tuam et cervicem tuam durissimam adhuc vivente me et ingrediente vobiscum semper contentiose egistis contra Dominum quanto magis cum mortuus fuero
DEUT|31|28|congregate ad me omnes maiores natu per tribus vestras atque doctores et loquar audientibus eis sermones istos et invocabo contra eos caelum et terram
DEUT|31|29|novi enim quod post mortem meam inique agetis et declinabitis cito de via quam praecepi vobis et occurrent vobis mala in extremo tempore quando feceritis malum in conspectu Domini ut inritetis eum per opera manuum vestrarum
DEUT|31|30|locutus est ergo Moses audiente universo coetu Israhel verba carminis huius et ad finem usque conplevit
DEUT|32|1|audite caeli quae loquor audiat terra verba oris mei
DEUT|32|2|concrescat in pluvia doctrina mea fluat ut ros eloquium meum quasi imber super herbam et quasi stillae super gramina
DEUT|32|3|quia nomen Domini invocabo date magnificentiam Deo nostro
DEUT|32|4|Dei perfecta sunt opera et omnes viae eius iudicia Deus fidelis et absque ulla iniquitate iustus et rectus
DEUT|32|5|peccaverunt ei non filii eius in sordibus generatio prava atque perversa
DEUT|32|6|haecine reddis Domino popule stulte et insipiens numquid non ipse est pater tuus qui possedit et fecit et creavit te
DEUT|32|7|memento dierum antiquorum cogita generationes singulas interroga patrem tuum et adnuntiabit tibi maiores tuos et dicent tibi
DEUT|32|8|quando dividebat Altissimus gentes quando separabat filios Adam constituit terminos populorum iuxta numerum filiorum Israhel
DEUT|32|9|pars autem Domini populus eius Iacob funiculus hereditatis eius
DEUT|32|10|invenit eum in terra deserta in loco horroris et vastae solitudinis circumduxit eum et docuit et custodivit quasi pupillam oculi sui
DEUT|32|11|sicut aquila provocans ad volandum pullos suos et super eos volitans expandit alas suas et adsumpsit eum atque portavit in umeris suis
DEUT|32|12|Dominus solus dux eius fuit et non erat cum eo deus alienus
DEUT|32|13|constituit eum super excelsam terram ut comederet fructus agrorum ut sugeret mel de petra oleumque de saxo durissimo
DEUT|32|14|butyrum de armento et lac de ovibus cum adipe agnorum et arietum filiorum Basan et hircos cum medulla tritici et sanguinem uvae biberet meracissimum
DEUT|32|15|incrassatus est dilectus et recalcitravit incrassatus inpinguatus dilatatus dereliquit Deum factorem suum et recessit a Deo salutari suo
DEUT|32|16|provocaverunt eum in diis alienis et in abominationibus ad iracundiam concitaverunt
DEUT|32|17|immolaverunt daemonibus et non Deo diis quos ignorabant novi recentesque venerunt quos non coluerunt patres eorum
DEUT|32|18|Deum qui te genuit dereliquisti et oblitus es Domini creatoris tui
DEUT|32|19|vidit Dominus et ad iracundiam concitatus est quia provocaverunt eum filii sui et filiae
DEUT|32|20|et ait abscondam faciem meam ab eis et considerabo novissima eorum generatio enim perversa est et infideles filii
DEUT|32|21|ipsi me provocaverunt in eo qui non erat Deus et inritaverunt in vanitatibus suis et ego provocabo eos in eo qui non est populus et in gente stulta inritabo illos
DEUT|32|22|ignis succensus est in furore meo et ardebit usque ad inferni novissima devorabitque terram cum germine suo et montium fundamenta conburet
DEUT|32|23|congregabo super eos mala et sagittas meas conplebo in eis
DEUT|32|24|consumentur fame et devorabunt eos aves morsu amarissimo dentes bestiarum inmittam in eos cum furore trahentium super terram atque serpentium
DEUT|32|25|foris vastabit eos gladius et intus pavor iuvenem simul ac virginem lactantem cum homine sene
DEUT|32|26|dixi ubinam sunt cessare faciam ex hominibus memoriam eorum
DEUT|32|27|sed propter iram inimicorum distuli ne forte superbirent hostes eorum et dicerent manus nostra excelsa et non Dominus fecit haec omnia
DEUT|32|28|gens absque consilio est et sine prudentia
DEUT|32|29|utinam saperent et intellegerent ac novissima providerent
DEUT|32|30|quomodo persequatur unus mille et duo fugent decem milia nonne ideo quia Deus suus vendidit eos et Dominus conclusit illos
DEUT|32|31|non enim est Deus noster ut deus eorum et inimici nostri sunt iudices
DEUT|32|32|de vinea Sodomorum vinea eorum et de suburbanis Gomorrae uva eorum uva fellis et botri amarissimi
DEUT|32|33|fel draconum vinum eorum et venenum aspidum insanabile
DEUT|32|34|nonne haec condita sunt apud me et signata in thesauris meis
DEUT|32|35|mea est ultio et ego retribuam in tempore ut labatur pes eorum iuxta est dies perditionis et adesse festinant tempora
DEUT|32|36|iudicabit Dominus populum suum et in servis suis miserebitur videbit quod infirmata sit manus et clausi quoque defecerint residuique consumpti sint
DEUT|32|37|et dicet ubi sunt dii eorum in quibus habebant fiduciam
DEUT|32|38|de quorum victimis comedebant adipes et bibebant vinum libaminum surgant et opitulentur vobis et in necessitate vos protegant
DEUT|32|39|videte quod ego sim solus et non sit alius deus praeter me ego occidam et ego vivere faciam percutiam et ego sanabo et non est qui de manu mea possit eruere
DEUT|32|40|levabo ad caelum manum meam et dicam vivo ego in aeternum
DEUT|32|41|si acuero ut fulgur gladium meum et arripuerit iudicium manus mea reddam ultionem hostibus meis et his qui oderunt me retribuam
DEUT|32|42|inebriabo sagittas meas sanguine et gladius meus devorabit carnes de cruore occisorum et de captivitate nudati inimicorum capitis
DEUT|32|43|laudate gentes populum eius quia sanguinem servorum suorum ulciscetur et vindictam retribuet in hostes eorum et propitius erit terrae populi sui
DEUT|32|44|venit ergo Moses et locutus est omnia verba cantici huius in auribus populi ipse et Iosue filius Nun
DEUT|32|45|conplevitque omnes sermones istos loquens ad universum Israhel
DEUT|32|46|et dixit ad eos ponite corda vestra in omnia verba quae ego testificor vobis hodie ut mandetis ea filiis vestris custodire et facere et implere universa quae scripta sunt legis huius
DEUT|32|47|quia non in cassum praecepta sunt vobis sed ut singuli in eis viverent quae facientes longo perseveretis tempore in terra ad quam Iordane transmisso ingredimini possidendam
DEUT|32|48|locutusque est Dominus ad Mosen in eadem die dicens
DEUT|32|49|ascende in montem istum Abarim id est transituum in montem Nebo qui est in terra Moab contra Hiericho et vide terram Chanaan quam ego tradam filiis Israhel obtinendam et morere in monte
DEUT|32|50|quem conscendens iungeris populis tuis sicut mortuus est Aaron frater tuus in monte Hor et adpositus populis suis
DEUT|32|51|quia praevaricati estis contra me in medio filiorum Israhel ad aquas Contradictionis in Cades deserti Sin et non sanctificastis me inter filios Israhel
DEUT|32|52|e contra videbis terram et non ingredieris in eam quam ego dabo filiis Israhel
DEUT|33|1|haec est benedictio qua benedixit Moses homo Dei filiis Israhel ante mortem suam
DEUT|33|2|et ait Dominus de Sina venit et de Seir ortus est nobis apparuit de monte Pharan et cum eo sanctorum milia in dextera eius ignea lex
DEUT|33|3|dilexit populos omnes sancti in manu illius sunt et qui adpropinquant pedibus eius accipient de doctrina illius
DEUT|33|4|legem praecepit nobis Moses hereditatem multitudinis Iacob
DEUT|33|5|erit apud rectissimum rex congregatis principibus populi cum tribubus Israhel
DEUT|33|6|vivat Ruben et non moriatur et sit parvus in numero
DEUT|33|7|haec est Iudae benedictio audi Domine vocem Iudae et ad populum suum introduc eum manus eius pugnabunt pro eo et adiutor illius contra adversarios eius erit
DEUT|33|8|Levi quoque ait perfectio tua et doctrina tua viro sancto tuo quem probasti in Temptatione et iudicasti ad aquas Contradictionis
DEUT|33|9|qui dixit patri suo et matri suae nescio vos et fratribus suis ignoro illos et nescierunt filios suos hii custodierunt eloquium tuum et pactum tuum servaverunt
DEUT|33|10|iudicia tua o Iacob et legem tuam o Israhel ponent thymiama in furore tuo et holocaustum super altare tuum
DEUT|33|11|benedic Domine fortitudini eius et opera manuum illius suscipe percute dorsa inimicorum eius et qui oderunt eum non consurgant
DEUT|33|12|et Beniamin ait amantissimus Domini habitabit confidenter in eo quasi in thalamo tota die morabitur et inter umeros illius requiescet
DEUT|33|13|Ioseph quoque ait de benedictione Domini terra eius de pomis caeli et rore atque abysso subiacente
DEUT|33|14|de pomis fructuum solis ac lunae
DEUT|33|15|de vertice antiquorum montium de pomis collium aeternorum
DEUT|33|16|et de frugibus terrae et plenitudine eius benedictio illius qui apparuit in rubo veniat super caput Ioseph et super verticem nazarei inter fratres suos
DEUT|33|17|quasi primogeniti tauri pulchritudo eius cornua rinocerotis cornua illius in ipsis ventilabit gentes usque ad terminos terrae hae sunt multitudines Ephraim et haec milia Manasse
DEUT|33|18|et Zabulon ait laetare Zabulon in exitu tuo et Isachar in tabernaculis tuis
DEUT|33|19|populos ad montem vocabunt ibi immolabunt victimas iustitiae qui inundationem maris quasi lac sugent et thesauros absconditos harenarum
DEUT|33|20|et Gad ait benedictus in latitudine Gad quasi leo requievit cepitque brachium et verticem
DEUT|33|21|et vidit principatum suum quod in parte sua doctor esset repositus qui fuit cum principibus populi et fecit iustitias Domini et iudicium suum cum Israhel
DEUT|33|22|Dan quoque ait Dan catulus leonis fluet largiter de Basan
DEUT|33|23|et Nepthalim dixit Nepthalim abundantia perfruetur et plenus erit benedictione Domini mare et meridiem possidebit
DEUT|33|24|Aser quoque ait benedictus in filiis Aser sit placens fratribus suis tinguat in oleo pedem suum
DEUT|33|25|ferrum et aes calciamentum eius sicut dies iuventutis tuae ita et senectus tua
DEUT|33|26|non est alius ut Deus rectissimi ascensor caeli auxiliator tuus magnificentia eius discurrunt nubes
DEUT|33|27|habitaculum eius sursum et subter brachia sempiterna eiciet a facie tua inimicum dicetque conterere
DEUT|33|28|habitabit Israhel confidenter et solus oculus Iacob in terra frumenti et vini caelique caligabunt rore
DEUT|33|29|beatus tu Israhel quis similis tui popule qui salvaris in Domino scutum auxilii tui et gladius gloriae tuae negabunt te inimici tui et tu eorum colla calcabis
DEUT|34|1|ascendit ergo Moses de campestribus Moab super montem Nebo in verticem Phasga contra Hiericho ostenditque ei Dominus omnem terram Galaad usque Dan
DEUT|34|2|et universum Nepthalim terramque Ephraim et Manasse et omnem terram usque ad mare Novissimum
DEUT|34|3|et australem partem et latitudinem campi Hiericho civitatis Palmarum usque Segor
DEUT|34|4|dixitque Dominus ad eum haec est terra pro qua iuravi Abraham Isaac et Iacob dicens semini tuo dabo eam vidisti eam oculis tuis et non transibis ad illam
DEUT|34|5|mortuusque est ibi Moses servus Domini in terra Moab iubente Domino
DEUT|34|6|et sepelivit eum in valle terrae Moab contra Phogor et non cognovit homo sepulchrum eius usque in praesentem diem
DEUT|34|7|Moses centum et viginti annorum erat quando mortuus est non caligavit oculus eius nec dentes illius moti sunt
DEUT|34|8|fleveruntque eum filii Israhel in campestribus Moab triginta diebus et conpleti sunt dies planctus lugentium Mosen
DEUT|34|9|Iosue vero filius Nun repletus est spiritu sapientiae quia Moses posuit super eum manus suas et oboedierunt ei filii Israhel feceruntque sicut praecepit Dominus Mosi
DEUT|34|10|et non surrexit propheta ultra in Israhel sicut Moses quem nosset Dominus facie ad faciem
DEUT|34|11|in omnibus signis atque portentis quae misit per eum ut faceret in terra Aegypti Pharaoni et omnibus servis eius universaeque terrae illius
DEUT|34|12|et cunctam manum robustam magnaque mirabilia quae fecit Moses coram universo Israhel
JOSH|1|1|et factum est ut post mortem Mosi servi Domini loqueretur Dominus ad Iosue filium Nun ministrum Mosi et diceret ei
JOSH|1|2|Moses servus meus mortuus est surge et transi Iordanem istum tu et omnis populus tecum in terram quam ego dabo filiis Israhel
JOSH|1|3|omnem locum quem calcaverit vestigium pedis vestri vobis tradam sicut locutus sum Mosi
JOSH|1|4|a deserto et Libano usque ad fluvium magnum Eufraten omnis terra Hettheorum usque ad mare Magnum contra solis occasum erit terminus vester
JOSH|1|5|nullus vobis poterit resistere cunctis diebus vitae tuae sicut fui cum Mose ero et tecum non dimittam nec derelinquam te
JOSH|1|6|confortare et esto robustus tu enim sorte divides populo huic terram pro qua iuravi patribus suis ut traderem eam illis
JOSH|1|7|confortare igitur et esto robustus valde ut custodias et facias omnem legem quam praecepit tibi Moses servus meus ne declines ab ea ad dextram vel ad sinistram ut intellegas cuncta quae agis
JOSH|1|8|non recedat volumen legis huius de ore tuo sed meditaberis in eo diebus ac noctibus ut custodias et facias omnia quae scripta sunt in eo tunc diriges viam tuam et intelleges eam
JOSH|1|9|ecce praecipio tibi confortare et esto robustus noli metuere et noli timere quoniam tecum est Dominus Deus tuus in omnibus ad quaecumque perrexeris
JOSH|1|10|praecepitque Iosue principibus populi dicens transite per medium castrorum et imperate populo ac dicite
JOSH|1|11|praeparate vobis cibaria quoniam post diem tertium transibitis Iordanem et intrabitis ad possidendam terram quam Dominus Deus vester daturus est vobis
JOSH|1|12|Rubenitis quoque et Gadditis et dimidiae tribui Manasse ait
JOSH|1|13|mementote sermonis quem praecepit vobis Moses famulus Domini dicens Dominus Deus vester dedit vobis requiem et omnem terram
JOSH|1|14|uxores vestrae et filii ac iumenta manebunt in terra quam tradidit vobis Moses trans Iordanem vos autem transite armati ante fratres vestros omnes fortes manu et pugnate pro eis
JOSH|1|15|donec det requiem Dominus fratribus vestris sicut et vobis dedit et possideant ipsi quoque terram quam Dominus Deus vester daturus est eis et sic revertemini in terram possessionis vestrae et habitabitis in ea quam vobis dedit Moses famulus Domini trans Iordanem contra solis ortum
JOSH|1|16|responderuntque ad Iosue atque dixerunt omnia quae praecepisti nobis faciemus et quocumque miseris ibimus
JOSH|1|17|sicut oboedivimus in cunctis Mosi ita oboediemus et tibi tantum sit Dominus Deus tecum sicut fuit cum Mose
JOSH|1|18|qui contradixerit ori tuo et non oboedierit cunctis sermonibus quos praeceperis ei moriatur tu tantum confortare et viriliter age
JOSH|2|1|misit ergo Iosue filius Nun de Setthim duos viros exploratores abscondito et dixit eis ite et considerate terram urbemque Hiericho qui pergentes ingressi sunt domum mulieris meretricis nomine Raab et quieverunt apud eam
JOSH|2|2|nuntiatumque est regi Hiericho et dictum ecce viri ingressi sunt huc per noctem de filiis Israhel ut explorarent terram
JOSH|2|3|misitque rex Hiericho ad Raab dicens educ viros qui venerunt ad te et ingressi sunt domum tuam exploratores quippe sunt et omnem terram considerare venerunt
JOSH|2|4|tollensque mulier viros abscondit et ait fateor venerunt ad me sed nesciebam unde essent
JOSH|2|5|cumque porta clauderetur in tenebris et illi pariter exierunt nescio quo abierunt persequimini cito et conprehendetis eos
JOSH|2|6|ipsa autem fecit ascendere viros in solarium domus suae operuitque eos lini stipula quae ibi erat
JOSH|2|7|hii autem qui missi fuerant secuti sunt eos per viam quae ducit ad vadum Iordanis illisque egressis statim porta clausa est
JOSH|2|8|necdum obdormierant qui latebant et ecce mulier ascendit ad eos et ait
JOSH|2|9|novi quod tradiderit Dominus vobis terram etenim inruit in nos terror vester et elanguerunt omnes habitatores terrae
JOSH|2|10|audivimus quod siccaverit Dominus aquas maris Rubri ad vestrum introitum quando egressi estis ex Aegypto et quae feceritis duobus Amorreorum regibus qui erant trans Iordanem Seon et Og quos interfecistis
JOSH|2|11|et haec audientes pertimuimus et elanguit cor nostrum nec remansit in nobis spiritus ad introitum vestrum Dominus enim Deus vester ipse est Deus in caelo sursum et in terra deorsum
JOSH|2|12|nunc ergo iurate mihi per Dominum ut quomodo ego feci vobiscum misericordiam ita et vos faciatis cum domo patris mei detisque mihi signum verum
JOSH|2|13|et salvetis patrem meum et matrem fratres ac sorores meas et omnia quae eorum sunt et eruatis animas nostras de morte
JOSH|2|14|qui responderunt ei anima nostra sit pro vobis in mortem si tamen non prodideris nos cumque tradiderit nobis Dominus terram faciemus in te misericordiam et veritatem
JOSH|2|15|dimisit ergo eos per funem de fenestra domus enim eius herebat muro
JOSH|2|16|dixitque ad eos ad montana conscendite ne forte occurrant vobis revertentes ibique latete diebus tribus donec redeant et sic ibitis per viam vestram
JOSH|2|17|qui dixerunt ad eam innoxii erimus a iuramento hoc quo adiurasti nos
JOSH|2|18|si ingredientibus nobis terram signum fuerit funiculus iste coccineus et ligaveris eum in fenestra per quam nos dimisisti et patrem tuum ac matrem fratresque et omnem cognationem tuam congregaveris in domum tuam
JOSH|2|19|qui ostium domus tuae egressus fuerit sanguis ipsius erit in caput eius et nos erimus alieni cunctorum autem sanguis qui tecum fuerint in domo redundabit in caput nostrum si eos aliquis tetigerit
JOSH|2|20|quod si nos prodere volueris et sermonem istum proferre in medium erimus mundi ab hoc iuramento quo adiurasti nos
JOSH|2|21|et illa respondit sicut locuti estis ita fiat dimittensque eos ut pergerent adpendit funiculum coccineum in fenestra
JOSH|2|22|illi vero ambulantes pervenerunt ad montana et manserunt ibi tres dies donec reverterentur qui fuerant persecuti quaerentes enim per omnem viam non reppererunt eos
JOSH|2|23|quibus urbem ingressis reversi sunt et descenderunt exploratores de monte et Iordane transmisso venerunt ad Iosue filium Nun narraveruntque ei omnia quae acciderant sibi
JOSH|2|24|atque dixerunt tradidit Dominus in manus nostras omnem terram hanc et timore prostrati sunt cuncti habitatores eius
JOSH|3|1|igitur Iosue de nocte consurgens movit castra egredientesque de Setthim venerunt ad Iordanem ipse et omnes filii Israhel et morati sunt ibi per tres dies
JOSH|3|2|quibus evolutis transierunt praecones per castrorum medium
JOSH|3|3|et clamare coeperunt quando videritis arcam foederis Domini Dei vestri et sacerdotes stirpis leviticae portantes eam vos quoque consurgite et sequimini praecedentes
JOSH|3|4|sitque inter vos et arcam spatium cubitorum duum milium ut procul videre possitis et nosse per quam viam ingrediamini quia prius non ambulastis per eam et cavete ne adpropinquetis ad arcam
JOSH|3|5|dixitque Iosue ad populum sanctificamini cras enim faciet Dominus inter vos mirabilia
JOSH|3|6|et ait ad sacerdotes tollite arcam foederis et praecedite populum qui iussa conplentes tulerunt et ambulaverunt ante eos
JOSH|3|7|dixitque Dominus ad Iosue hodie incipiam exaltare te coram omni Israhel ut sciant quod sicut cum Mosi fui ita et tecum sim
JOSH|3|8|tu autem praecipe sacerdotibus qui portant arcam foederis et dic eis cum ingressi fueritis partem aquae Iordanis state in ea
JOSH|3|9|dixitque Iosue ad filios Israhel accedite huc et audite verba Domini Dei vestri
JOSH|3|10|et rursum in hoc inquit scietis quod Dominus Deus vivens in medio vestri est et disperdat in conspectu vestro Chananeum Hettheum Eveum et Ferezeum Gergeseum quoque et Amorreum et Iebuseum
JOSH|3|11|ecce arca foederis Domini omnis terrae antecedet vos per Iordanem
JOSH|3|12|parate duodecim viros de tribubus Israhel singulos per singulas tribus
JOSH|3|13|et cum posuerint vestigia pedum suorum sacerdotes qui portant arcam Domini Dei universae terrae in aquis Iordanis aquae quae inferiores sunt decurrent atque deficient quae autem desuper veniunt in una mole consistent
JOSH|3|14|igitur egressus est populus de tabernaculis suis ut transirent Iordanem et sacerdotes qui portabant arcam foederis pergebant ante eum
JOSH|3|15|ingressisque eis Iordanem et pedibus eorum tinctis in parte aquae cum Iordanis autem ripas alvei sui tempore messis impleret
JOSH|3|16|steterunt aquae descendentes in uno loco et instar montis intumescentes apparebant procul ab urbe quae vocatur Adom usque ad locum Sarthan quae autem inferiores erant in mare Solitudinis quod nunc vocatur Mortuum descenderunt usquequo omnino deficerent
JOSH|3|17|populus autem incedebat contra Iordanem et sacerdotes qui portabant arcam foederis Domini stabant super siccam humum in medio Iordanis accincti omnisque populus per arentem alveum transiebat
JOSH|4|1|quibus transgressis dixit Dominus ad Iosue
JOSH|4|2|elige duodecim viros singulos per singulas tribus
JOSH|4|3|et praecipe eis ut tollant de medio Iordanis alveo ubi steterunt sacerdotum pedes duodecim durissimos lapides quos ponetis in loco castrorum ubi fixeritis hac nocte tentoria
JOSH|4|4|vocavitque Iosue duodecim viros quos elegerat de filiis Israhel singulos de tribubus singulis
JOSH|4|5|et ait ad eos ite ante arcam Domini Dei vestri ad Iordanis medium et portate singuli singulos lapides in umeris vestris iuxta numerum filiorum Israhel
JOSH|4|6|ut sit signum inter vos et quando interrogaverint vos filii vestri cras dicentes quid sibi volunt isti lapides
JOSH|4|7|respondebitis eis defecerunt aquae Iordanis ante arcam foederis Domini cum transiret eum idcirco positi sunt lapides isti in monumentum filiorum Israhel usque in aeternum
JOSH|4|8|fecerunt ergo filii Israhel sicut eis praecepit Iosue portantes de medio Iordanis alveo duodecim lapides ut ei Dominus imperarat iuxta numerum filiorum Israhel usque ad locum in quo castrametati sunt ibique posuerunt eos
JOSH|4|9|alios quoque duodecim lapides posuit Iosue in medio Iordanis alveo ubi steterunt sacerdotes qui portabant arcam foederis et sunt ibi usque in praesentem diem
JOSH|4|10|sacerdotes autem qui portabant arcam stabant in Iordanis medio donec omnia conplerentur quae Iosue ut loqueretur ad populum praeceperat Dominus et dixerat ei Moses festinavitque populus et transiit
JOSH|4|11|cumque transissent omnes transivit et arca Domini sacerdotesque pergebant ante populum
JOSH|4|12|filii quoque Ruben et Gad et dimidiae tribus Manasse armati praecedebant filios Israhel sicut eis praeceperat Moses
JOSH|4|13|et quadraginta pugnatorum milia per turmas et cuneos incedebant per plana atque campestria urbis Hiericho
JOSH|4|14|in illo die magnificavit Dominus Iosue coram omni Israhel ut timerent eum sicut timuerant Mosen dum adviveret
JOSH|4|15|dixitque ad eum
JOSH|4|16|praecipe sacerdotibus qui portant arcam foederis ut ascendant de Iordane
JOSH|4|17|qui praecepit eis dicens ascendite de Iordane
JOSH|4|18|cumque ascendissent portantes arcam foederis Domini et siccam humum calcare coepissent reversae sunt aquae in alveum suum et fluebant sicut ante consueverant
JOSH|4|19|populus autem ascendit de Iordane decimo mensis primi die et castrametati sunt in Galgalis contra orientalem plagam urbis Hiericho
JOSH|4|20|duodecim quoque lapides quos de Iordanis alveo sumpserant posuit Iosue in Galgalis
JOSH|4|21|et dixit ad filios Israhel quando interrogaverint filii vestri cras patres suos et dixerint eis quid sibi volunt isti lapides
JOSH|4|22|docebitis eos atque dicetis per arentem alveum transivit Israhel Iordanem istum
JOSH|4|23|siccante Domino Deo vestro aquas eius in conspectu vestro donec transiretis
JOSH|4|24|sicut fecerat prius in mari Rubro quod siccavit donec transiremus
JOSH|4|25|ut discant omnes terrarum populi fortissimam Domini manum et ut vos timeatis Dominum Deum vestrum omni tempore
JOSH|5|1|postquam ergo audierunt omnes reges Amorreorum qui habitabant trans Iordanem ad occidentalem plagam et cuncti reges Chanaan qui propinqua possidebant Magno mari loca quod siccasset Dominus fluenta Iordanis coram filiis Israhel donec transirent dissolutum est cor eorum et non remansit in eis spiritus timentium introitum filiorum Israhel
JOSH|5|2|eo tempore ait Dominus ad Iosue fac tibi cultros lapideos et circumcide secundo filios Israhel
JOSH|5|3|fecit quod iusserat Dominus et circumcidit filios Israhel in colle Praeputiorum
JOSH|5|4|haec autem causa est secundae circumcisionis omnis populus qui egressus est ex Aegypto generis masculini universi bellatores viri mortui sunt in deserto per longissimos viae circuitus
JOSH|5|5|qui omnes circumcisi erant populus autem qui natus est in deserto
JOSH|5|6|per quadraginta annos itineris latissimae solitudinis incircumcisus fuit donec consumerentur qui non audierant vocem Domini et quibus ante iuraverat ut ostenderet eis terram lacte et melle manantem
JOSH|5|7|horum filii in locum successerunt patrum et circumcisi sunt ab Iosue quia sicut nati fuerant in praeputio erant nec eos in via aliquis circumciderat
JOSH|5|8|postquam autem omnes circumcisi sunt manserunt in eodem castrorum loco donec sanarentur
JOSH|5|9|dixitque Dominus ad Iosue hodie abstuli obprobrium Aegypti a vobis vocatumque est nomen loci illius Galgala usque in praesentem diem
JOSH|5|10|manseruntque filii Israhel in Galgalis et fecerunt phase quartadecima die mensis ad vesperum in campestribus Hiericho
JOSH|5|11|et comederunt de frugibus terrae die altero azymos panes et pulentam eiusdem anni
JOSH|5|12|defecitque manna postquam comederunt de frugibus terrae nec usi sunt ultra illo cibo filii Israhel sed comederunt de frugibus praesentis anni terrae Chanaan
JOSH|5|13|cum autem esset Iosue in agro urbis Hiericho levavit oculos et vidit virum stantem contra se et evaginatum tenentem gladium perrexitque ad eum et ait noster es an adversariorum
JOSH|5|14|qui respondit nequaquam sed sum princeps exercitus Domini et nunc venio
JOSH|5|15|cecidit Iosue pronus in terram et adorans ait quid dominus meus loquitur ad servum suum
JOSH|5|16|solve inquit calciamentum de pedibus tuis locus enim in quo stas sanctus est fecitque Iosue ut sibi fuerat imperatum
JOSH|6|1|Hiericho autem clausa erat atque munita timore filiorum Israhel et nullus egredi audebat aut ingredi
JOSH|6|2|dixitque Dominus ad Iosue ecce dedi in manus tuas Hiericho et regem eius omnesque fortes viros
JOSH|6|3|circuite urbem cuncti bellatores semel per diem sic facietis sex diebus
JOSH|6|4|septimo autem die sacerdotes tollant septem bucinas quarum usus est in iobeleo et praecedant arcam foederis septiesque circuibitis civitatem et sacerdotes clangent bucinis
JOSH|6|5|cumque insonuerit vox tubae longior atque concisior et in auribus vestris increpuerit conclamabit omnis populus vociferatione maxima et muri funditus corruent civitatis ingredienturque singuli per locum contra quem steterint
JOSH|6|6|vocavit ergo Iosue filius Nun sacerdotes et dixit ad eos tollite arcam foederis et septem alii sacerdotes tollant septem iobeleorum bucinas et incedant ante arcam Domini
JOSH|6|7|ad populum quoque ait vadite et circuite civitatem armati praecedentes arcam Domini
JOSH|6|8|cumque Iosue verba finisset et septem sacerdotes septem bucinis clangerent ante arcam foederis Domini
JOSH|6|9|omnisque praecederet armatus exercitus reliquum vulgus arcam sequebatur ac bucinis omnia concrepabant
JOSH|6|10|praeceperat autem Iosue populo dicens non clamabitis nec audietur vox vestra neque ullus sermo ex ore vestro egredietur donec veniat dies in quo dicam vobis clamate et vociferamini
JOSH|6|11|circuivit ergo arca Domini civitatem semel per diem et reversa in castra mansit ibi
JOSH|6|12|igitur Iosue de nocte consurgente tulerunt sacerdotes arcam Domini
JOSH|6|13|et septem ex eis septem bucinas quarum in iobeleis usus est praecedebantque arcam Domini ambulantes atque clangentes et armatus populus ibat ante eos vulgus autem reliquum sequebatur arcam et bucinis personabat
JOSH|6|14|circumieruntque civitatem secundo die semel et reversi sunt in castra sic fecerunt sex diebus
JOSH|6|15|die autem septimo diluculo consurgentes circumierunt urbem sicut dispositum erat septies
JOSH|6|16|cumque septimo circuitu clangerent bucinis sacerdotes dixit Iosue ad omnem Israhel vociferamini tradidit enim vobis Dominus civitatem
JOSH|6|17|sitque civitas haec anathema et omnia quae in ea sunt Domino sola Raab meretrix vivat cum universis qui cum ea in domo sunt abscondit enim nuntios quos direximus
JOSH|6|18|vos autem cavete ne de his quae praecepta sunt quippiam contingatis et sitis praevaricationis rei et omnia castra Israhel sub peccato sint atque turbentur
JOSH|6|19|quicquid autem auri et argenti fuerit et vasorum aeneorum ac ferri Domino consecretur repositum in thesauris eius
JOSH|6|20|igitur omni vociferante populo et clangentibus tubis postquam in aures multitudinis vox sonitusque increpuit muri ilico corruerunt et ascendit unusquisque per locum qui contra se erat ceperuntque civitatem
JOSH|6|21|et interfecerunt omnia quae erant in ea a viro usque ad mulierem ab infante usque ad senem boves quoque et oves et asinos in ore gladii percusserunt
JOSH|6|22|duobus autem viris qui exploratores missi fuerant dixit Iosue ingredimini domum mulieris meretricis et producite eam omniaque quae illius sunt sicut illi iuramento firmastis
JOSH|6|23|ingressique iuvenes eduxerunt Raab et parentes eius fratres quoque et cunctam supellectilem ac cognationem illius et extra castra Israhel manere fecerunt
JOSH|6|24|urbem autem et omnia quae in ea sunt succenderunt absque argento et auro et vasis aeneis ac ferro quae in aerarium Domini consecrarunt
JOSH|6|25|Raab vero meretricem et domum patris eius atque omnia quae habebat fecit Iosue vivere et habitaverunt in medio Israhel usque in praesentem diem eo quod absconderit nuntios quos miserat ut explorarent Hiericho in tempore illo inprecatus est Iosue dicens
JOSH|6|26|maledictus vir coram Domino qui suscitaverit et aedificaverit civitatem Hiericho in primogenito suo fundamenta illius iaciat et in novissimo liberorum ponat portas eius
JOSH|6|27|fuit ergo Dominus cum Iosue et nomen eius in omni terra vulgatum est
JOSH|7|1|filii autem Israhel praevaricati sunt mandatum et usurpaverunt de anathemate nam Achan filius Charmi filii Zabdi filii Zare de tribu Iuda tulit aliquid de anathemate iratusque est Dominus contra filios Israhel
JOSH|7|2|cumque mitteret Iosue de Hiericho viros contra Ahi quae est iuxta Bethaven ad orientalem plagam oppidi Bethel dixit eis ascendite et explorate terram qui praecepta conplentes exploraverunt Ahi
JOSH|7|3|et reversi dixerunt ei non ascendat omnis populus sed duo vel tria milia virorum pergant et deleant civitatem quare omnis populus frustra vexatur contra hostes paucissimos
JOSH|7|4|ascenderunt ergo tria milia pugnatores qui statim terga vertentes
JOSH|7|5|percussi sunt a viris urbis Ahi et corruerunt ex eis triginta et sex homines persecutique sunt eos adversarii de porta usque Sabarim et ceciderunt per prona fugientes pertimuitque cor populi et instar aquae liquefactum est
JOSH|7|6|Iosue vero scidit vestimenta sua et cecidit pronus in terram coram arca Domini usque ad vesperum tam ipse quam omnes senes Israhel miseruntque pulverem super capita sua
JOSH|7|7|et dixit Iosue heu Domine Deus quid voluisti transducere populum istum Iordanem fluvium ut traderes nos in manus Amorrei et perderes utinam ut coepimus mansissemus trans Iordanem
JOSH|7|8|mi Domine Deus quid dicam videns Israhelem hostibus suis terga vertentem
JOSH|7|9|audient Chananei et omnes habitatores terrae ac pariter conglobati circumdabunt nos atque delebunt nomen nostrum de terra et quid facies magno nomini tuo
JOSH|7|10|dixitque Dominus ad Iosue surge cur iaces pronus in terra
JOSH|7|11|peccavit Israhel et praevaricatus est pactum meum tuleruntque de anathemate et furati sunt atque mentiti et absconderunt inter vasa sua
JOSH|7|12|nec poterit Israhel stare ante hostes suos eosque fugiet quia pollutus est anathemate non ero ultra vobiscum donec conteratis eum qui huius sceleris reus est
JOSH|7|13|surge sanctifica populum et dic eis sanctificamini in crastinum haec enim dicit Dominus Deus Israhel anathema in medio tui est Israhel non poteris stare coram hostibus tuis donec deleatur ex te qui hoc contaminatus est scelere
JOSH|7|14|accedetisque mane singuli per tribus vestras et quamcumque tribum sors invenerit accedet per cognationes suas et cognatio per domos domusque per viros
JOSH|7|15|et quicumque ille in hoc facinore fuerit deprehensus conburetur igni cum omni substantia sua quoniam praevaricatus est pactum Domini et fecit nefas in Israhel
JOSH|7|16|surgens itaque Iosue mane adplicavit Israhel per tribus suas et inventa est tribus Iuda
JOSH|7|17|quae cum iuxta familias suas esset oblata inventa est familia Zarai illam quoque per viros offerens repperit Zabdi
JOSH|7|18|cuius domum in singulos dividens viros invenit Achan filium Charmi filii Zabdi filii Zare de tribu Iuda
JOSH|7|19|et ait ad Achan fili mi da gloriam Domino Deo Israhel et confitere atque indica mihi quid feceris ne abscondas
JOSH|7|20|responditque Achan Iosue et dixit ei vere ego peccavi Domino Deo Israhel et sic et sic feci
JOSH|7|21|vidi enim inter spolia pallium coccineum valde bonum et ducentos siclos argenti regulamque auream quinquaginta siclorum et concupiscens abstuli et abscondi in terra contra medium tabernaculi mei argentumque fossa humo operui
JOSH|7|22|misit ergo Iosue ministros qui currentes ad tabernaculum illius reppererunt cuncta abscondita in eodem loco et argentum simul
JOSH|7|23|auferentesque de tentorio tulerunt ea ad Iosue et ad omnes filios Israhel proieceruntque ante Dominum
JOSH|7|24|tollens itaque Iosue Achan filium Zare argentumque et pallium et auream regulam filiosque eius et filias boves et asinos et oves ipsumque tabernaculum et cunctam supellectilem et omnis Israhel cum eo duxerunt eos ad vallem Achor
JOSH|7|25|ubi dixit Iosue quia turbasti nos exturbet te Dominus in die hac lapidavitque eum omnis Israhel et cuncta quae illius erant igne consumpta sunt
JOSH|7|26|congregaverunt quoque super eum acervum magnum lapidum qui permanet usque in praesentem diem et aversus est furor Domini ab eis vocatumque est nomen loci illius vallis Achor usque hodie
JOSH|8|1|dixit autem Dominus ad Iosue ne timeas neque formides tolle tecum omnem multitudinem pugnatorum et consurgens ascende in oppidum Ahi ecce tradidi in manu tua regem eius et populum urbemque et terram
JOSH|8|2|faciesque urbi Ahi et regi eius sicut fecisti Hiericho et regi illius praedam vero et omnia animantia diripietis vobis pone insidias urbi post eam
JOSH|8|3|surrexitque Iosue et omnis exercitus bellatorum cum eo ut ascenderent in Ahi et electa triginta milia virorum fortium misit nocte
JOSH|8|4|praecepitque eis dicens ponite insidias post civitatem nec longius recedatis et eritis omnes parati
JOSH|8|5|ego autem et reliqua multitudo quae mecum est accedemus ex adverso contra urbem cumque exierint contra nos sicut ante fecimus fugiemus et terga vertemus
JOSH|8|6|donec persequentes ab urbe longius protrahantur putabunt enim fugere nos sicut prius
JOSH|8|7|nobis ergo fugientibus et illis sequentibus consurgetis de insidiis et vastabitis civitatem tradetque eam Dominus Deus vester in manus vestras
JOSH|8|8|cumque ceperitis succendite eam sic omnia facietis ut iussi
JOSH|8|9|dimisitque eos et perrexerunt ad insidiarum locum sederuntque inter Bethel et Ahi ad occidentalem plagam urbis Ahi Iosue autem nocte illa in medio mansit populi
JOSH|8|10|surgensque diluculo recensuit socios et ascendit cum senioribus in fronte exercitus vallatus auxilio pugnatorum
JOSH|8|11|cumque venissent et ascendissent ex adverso civitatis steterunt ad septentrionalem urbis plagam inter quam et eos vallis media erat
JOSH|8|12|quinque milia autem viros elegerat et posuerat in insidiis inter Bethaven et Ahi ex occidentali parte eiusdem civitatis
JOSH|8|13|omnis vero reliquus exercitus ad aquilonem aciem dirigebat ita ut novissimi multitudinis occidentalem plagam urbis adtingerent abiit ergo Iosue nocte illa et stetit in vallis medio
JOSH|8|14|quod cum vidisset rex Ahi festinavit mane et egressus est cum omni exercitu civitatis direxitque aciem contra desertum ignorans quod post tergum laterent insidiae
JOSH|8|15|Iosue vero et omnis Israhel cesserunt loco simulantes metum et fugientes per viam solitudinis
JOSH|8|16|at illi vociferantes pariter et se mutuo cohortantes persecuti sunt eos cumque recessissent a civitate
JOSH|8|17|et ne unus quidem in urbe Ahi et Bethel remansisset qui non persequeretur Israhel sicut eruperant aperta oppida relinquentes
JOSH|8|18|dixit Dominus ad Iosue leva clypeum qui in manu tua est contra urbem Ahi quoniam tibi tradam eam
JOSH|8|19|cumque elevasset clypeum ex adverso civitatis insidiae quae latebant surrexerunt confestim et pergentes ad civitatem ceperunt et succenderunt eam
JOSH|8|20|viri autem civitatis qui persequebantur Iosue respicientes et videntes fumum urbis ad caelum usque conscendere non potuerunt ultra huc illucque diffugere praesertim cum hii qui simulaverant fugam et tendebant ad solitudinem contra persequentes fortissime restitissent
JOSH|8|21|vidensque Iosue et omnis Israhel quod capta esset civitas et fumus urbis ascenderet reversus percussit viros Ahi
JOSH|8|22|siquidem et illi qui ceperant et succenderant civitatem egressi ex urbe contra suos medios hostium ferire coeperunt cum ergo ex utraque parte adversarii caederentur ita ut nullus de tanta multitudine salvaretur
JOSH|8|23|regem quoque urbis Ahi adprehendere viventem et obtulerunt Iosue
JOSH|8|24|igitur omnibus interfectis qui Israhelem ad deserta tendentem fuerant persecuti et in eodem loco gladio corruentibus reversi filii Israhel percusserunt civitatem
JOSH|8|25|erant autem qui in eo die conciderant a viro usque ad mulierem duodecim milia hominum omnes urbis Ahi
JOSH|8|26|Iosue vero non contraxit manum quam in sublime porrexerat tenens clypeum donec interficerentur omnes habitatores Ahi
JOSH|8|27|iumenta autem et praedam civitatis diviserunt sibi filii Israhel sicut praeceperat Dominus Iosue
JOSH|8|28|qui succendit urbem et fecit eam tumulum sempiternum
JOSH|8|29|regem quoque eius suspendit in patibulo usque ad vesperum et solis occasum praecepitque et deposuerunt cadaver eius de cruce proieceruntque in ipso introitu civitatis congesto super eum magno acervo lapidum qui permanet usque in praesentem diem
JOSH|8|30|tunc aedificavit Iosue altare Domino Deo Israhel in monte Hebal
JOSH|8|31|sicut praeceperat Moses famulus Domini filiis Israhel et scriptum est in volumine legis Mosi altare de lapidibus inpolitis quos ferrum non tetigit et obtulit super eo holocausta Domino immolavitque pacificas victimas
JOSH|8|32|et scripsit super lapides deuteronomium legis Mosi quod ille digesserat coram filiis Israhel
JOSH|8|33|omnis autem populus et maiores natu ducesque ac iudices stabant ex utraque parte arcae in conspectu sacerdotum qui portabant arcam foederis Domini ut advena ita et indigena media eorum pars iuxta montem Garizim et media iuxta montem Hebal sicut praeceperat Moses famulus Domini et primum quidem benedixit populo Israhel
JOSH|8|34|post haec legit omnia verba benedictionis et maledictionis et cuncta quae scripta erant in legis volumine
JOSH|8|35|nihil ex his quae Moses iusserat reliquit intactum sed universa replicavit coram omni multitudine Israhel mulieribus ac parvulis et advenis qui inter eos morabantur
JOSH|9|1|quibus auditis cuncti reges trans Iordanem qui versabantur in montanis et in campestribus in maritimis ac litore maris Magni hii quoque qui habitabant iuxta Libanum Hettheus et Amorreus et Chananeus Ferezeus et Eveus et Iebuseus
JOSH|9|2|congregati sunt pariter ut pugnarent contra Iosue et Israhel uno animo eademque sententia
JOSH|9|3|at hii qui habitabant in Gabaon audientes cuncta quae fecerat Iosue Hiericho et Ahi
JOSH|9|4|et callide cogitantes tulerunt sibi cibaria saccos veteres asinis inponentes et utres vinarios scissos atque consutos
JOSH|9|5|calciamentaque perantiqua quae ad indicium vetustatis pittaciis consuta erant induti veteribus vestimentis panes quoque quos portabant ob viaticum duri erant et in frusta comminuti
JOSH|9|6|perrexeruntque ad Iosue qui tunc morabatur in castris Galgalae et dixerunt ei atque omni simul Israheli de terra longinqua venimus pacem vobiscum facere cupientes responderuntque viri Israhel ad eos atque dixerunt
JOSH|9|7|ne forsitan in terra quae nobis sorte debetur habitetis et non possimus foedus inire vobiscum
JOSH|9|8|at illi ad Iosue servi inquiunt tui sumus quibus Iosue quinam ait estis et unde venistis
JOSH|9|9|responderunt de terra longinqua valde venerunt servi tui in nomine Domini Dei tui audivimus enim famam potentiae eius cuncta quae fecit in Aegypto
JOSH|9|10|et duobus Amorreorum regibus trans Iordanem Seon regi Esebon et Og regi Basan qui erat in Astharoth
JOSH|9|11|dixeruntque nobis seniores et omnes habitatores terrae nostrae tollite in manibus cibaria ob longissimam viam et occurrite eis ac dicite servi vestri sumus foedus inite nobiscum
JOSH|9|12|en panes quando egressi sumus de domibus nostris ut veniremus ad vos calidos sumpsimus nunc sicci facti sunt et vetustate nimia comminuti
JOSH|9|13|utres vini novos implevimus nunc rupti sunt et soluti vestes et calciamenta quibus induimur et quae habemus in pedibus ob longitudinem largioris viae trita sunt et paene consumpta
JOSH|9|14|susceperunt igitur de cibariis eorum et os Domini non interrogaverunt
JOSH|9|15|fecitque Iosue cum eis pacem et inito foedere pollicitus est quod non occiderentur principes quoque multitudinis iuraverunt eis
JOSH|9|16|post dies autem tres initi foederis audierunt quod in vicino habitarent et inter eos futuri essent
JOSH|9|17|moveruntque castra filii Israhel et venerunt in civitates eorum die tertio quarum haec vocabula sunt Gabaon et Caphira et Beroth et Cariathiarim
JOSH|9|18|et non percusserunt eos eo quod iurassent eis principes multitudinis in nomine Domini Dei Israhel murmuravit itaque omne vulgus contra principes
JOSH|9|19|qui responderunt eis iuravimus illis in nomine Domini Dei Israhel et idcirco non possumus eos contingere
JOSH|9|20|sed hoc faciemus eis reserventur quidem ut vivant ne contra nos ira Domini concitetur si peieraverimus
JOSH|9|21|sed sic vivant ut in usus universae multitudinis ligna caedant aquasque conportent quibus haec loquentibus
JOSH|9|22|vocavit Gabaonitas Iosue et dixit eis cur nos decipere fraude voluistis ut diceretis procul valde habitamus a vobis cum in medio nostri sitis
JOSH|9|23|itaque sub maledictione eritis et non deficiet de stirpe vestra ligna caedens aquasque conportans in domum Dei mei
JOSH|9|24|qui responderunt nuntiatum est nobis servis tuis quae promisisset Dominus Deus tuus Mosi servo suo ut traderet vobis omnem terram et disperderet cunctos habitatores eius timuimus igitur valde et providimus animabus nostris vestro terrore conpulsi et hoc consilium inivimus
JOSH|9|25|nunc autem in manu tua sumus quod tibi bonum et rectum videtur fac nobis
JOSH|9|26|fecit ergo Iosue ut dixerat et liberavit eos de manibus filiorum Israhel ut non occiderentur
JOSH|9|27|decrevitque in illo die esse eos in ministerium cuncti populi et altaris Domini caedentes ligna et aquas conportantes usque in praesens tempus in loco quem Dominus elegisset
JOSH|10|1|quae cum audisset Adonisedec rex Hierusalem quod scilicet cepisset Iosue Ahi et subvertisset eam sicut enim fecerat Hiericho et regi eius sic fecit Ahi et regi illius et quod transfugissent Gabaonitae ad Israhel et essent foederati eorum
JOSH|10|2|timuit valde urbs enim magna erat Gabaon et una regalium civitatum et maior oppido Ahi omnesque bellatores eius fortissimi
JOSH|10|3|misit ergo Adonisedec rex Hierusalem ad Oham regem Hebron et ad Pharam regem Hieremoth ad Iaphie quoque regem Lachis et ad Dabir regem Eglon dicens
JOSH|10|4|ascendite ad me et ferte praesidium ut expugnemus Gabaon quare transfugerit ad Iosue et filios Israhel
JOSH|10|5|congregati igitur ascenderunt quinque reges Amorreorum rex Hierusalem rex Hebron rex Hieremoth rex Lachis rex Eglon simul cum exercitibus suis et castrametati sunt circa Gabaon obpugnantes eam
JOSH|10|6|habitatores autem Gabaon urbis obsessae miserunt ad Iosue qui tunc morabatur in castris apud Galgalam et dixerunt ei ne retrahas manus tuas ab auxilio servorum tuorum ascende cito et libera nos ferque praesidium convenerunt enim adversum nos omnes reges Amorreorum qui habitant in montanis
JOSH|10|7|ascenditque Iosue de Galgalis et omnis exercitus bellatorum cum eo viri fortissimi
JOSH|10|8|dixitque Dominus ad Iosue ne timeas eos in manus enim tuas tradidi illos nullus tibi ex eis resistere poterit
JOSH|10|9|inruit itaque Iosue super eos repente tota ascendens nocte de Galgalis
JOSH|10|10|et conturbavit eos Dominus a facie Israhel contrivitque plaga magna in Gabaon ac persecutus est per viam ascensus Bethoron et percussit usque Azeca et Maceda
JOSH|10|11|cumque fugerent filios Israhel et essent in descensu Bethoron Dominus misit super eos lapides magnos de caelo usque Azeca et mortui sunt multo plures lapidibus grandinis quam quos gladio percusserant filii Israhel
JOSH|10|12|tunc locutus est Iosue Domino in die qua tradidit Amorreum in conspectu filiorum Israhel dixitque coram eis sol contra Gabaon ne movearis et luna contra vallem Ahialon
JOSH|10|13|steteruntque sol et luna donec ulcisceretur se gens de inimicis suis nonne scriptum est hoc in libro Iustorum stetit itaque sol in medio caeli et non festinavit occumbere spatio unius diei
JOSH|10|14|non fuit ante et postea tam longa dies oboediente Domino voci hominis et pugnante pro Israhel
JOSH|10|15|reversusque est Iosue cum omni Israhel in castra Galgalae
JOSH|10|16|fugerant enim quinque reges et se absconderant in spelunca urbis Maceda
JOSH|10|17|nuntiatumque est Iosue quod inventi essent quinque reges latentes in spelunca Maceda
JOSH|10|18|qui praecepit sociis et ait volvite saxa ingentia ad os speluncae et ponite viros industrios qui clausos custodiant
JOSH|10|19|vos autem nolite stare sed persequimini hostes et extremos quosque fugientium caedite ne dimittatis eos urbium suarum intrare praesidia quos tradidit Dominus Deus in manus vestras
JOSH|10|20|caesis igitur adversariis plaga magna et usque ad internicionem paene consumptis hii qui Israhel effugere potuerunt ingressi sunt civitates munitas
JOSH|10|21|reversusque est omnis exercitus ad Iosue in Maceda ubi tunc erant castra sani et integro numero nullusque contra filios Israhel muttire ausus est
JOSH|10|22|praecepitque Iosue dicens aperite os speluncae et producite ad me quinque reges qui in ea latitant
JOSH|10|23|fecerunt ministri ut sibi fuerat imperatum et eduxerunt ad eum quinque reges de spelunca regem Hierusalem regem Hebron regem Hieremoth regem Lachis regem Eglon
JOSH|10|24|cumque educti essent ad eum vocavit omnes viros Israhel et ait ad principes exercitus qui secum erant ite et ponite pedes super colla regum istorum qui cum perrexissent et subiectorum pedibus colla calcarent
JOSH|10|25|rursum ait ad eos nolite timere nec paveatis confortamini et estote robusti sic enim faciet Dominus cunctis hostibus vestris adversum quos dimicatis
JOSH|10|26|percussitque Iosue et interfecit eos atque suspendit super quinque stipites fueruntque suspensi usque ad vesperum
JOSH|10|27|cumque occumberet sol praecepit sociis ut deponerent eos de patibulis qui depositos proiecerunt in speluncam in qua latuerant et posuerunt super os eius saxa ingentia quae permanent usque in praesens
JOSH|10|28|eodem die Macedam quoque cepit Iosue et percussit in ore gladii regemque illius interfecit et omnes habitatores eius non dimisit in ea saltim parvas reliquias fecitque regi Maceda sicut fecerat regi Hiericho
JOSH|10|29|transivit cum omni Israhel de Maceda in Lebna et pugnabat contra eam
JOSH|10|30|quam tradidit Dominus cum rege suo in manu Israhel percusseruntque urbem in ore gladii et omnes habitatores eius non dimiserunt in ea ullas reliquias feceruntque regi Lebna sicut fecerant regi Hiericho
JOSH|10|31|de Lebna transivit in Lachis et exercitu per gyrum disposito obpugnabat eam
JOSH|10|32|tradiditque Dominus Lachis in manu Israhel et cepit eam die altero atque percussit in ore gladii omnemque animam quae fuerat in ea sicut fecerat Lebna
JOSH|10|33|eo tempore ascendit Hiram rex Gazer ut auxiliaretur Lachis quem percussit Iosue cum omni populo eius usque ad internicionem
JOSH|10|34|transivitque de Lachis in Eglon et circumdedit
JOSH|10|35|atque expugnavit eam eadem die percussitque in ore gladii omnes animas quae erant in ea iuxta omnia quae fecerat Lachis
JOSH|10|36|ascendit quoque cum omni Israhele de Eglon in Hebron et pugnavit contra eam
JOSH|10|37|cepitque et percussit in ore gladii regem quoque eius et omnia oppida regionis illius universasque animas quae in ea fuerant commoratae non reliquit in ea ullas reliquias sicut fecerat Eglon sic fecit et Hebron cuncta quae in ea repperit consumens gladio
JOSH|10|38|inde reversus in Dabir
JOSH|10|39|cepit eam atque vastavit
JOSH|10|40|regem quoque eius et omnia per circuitum oppida percussit in ore gladii non dimisit in ea ullas reliquias sicut fecerat Hebron et Lebna et regibus earum sic fecit Dabir et regi illius
JOSH|10|41|percussit itaque Iosue omnem terram montanam et meridianam atque campestrem et Asedoth cum regibus suis non dimisit in ea ullas reliquias sed omne quod spirare poterat interfecit sicut praeceperat ei Dominus Deus Israhel
JOSH|10|42|a Cadesbarne usque Gazam omnem terram Gosen usque Gabaon
JOSH|10|43|universos reges et regiones eorum uno cepit impetu atque vastavit Dominus enim Deus Israhel pugnabat pro eo
JOSH|10|44|reversusque est cum omni Israhele ad locum castrorum in Galgala
JOSH|11|1|quae cum audisset Iabin rex Asor misit ad Iobab regem Madon et ad regem Someron atque ad regem Acsaph
JOSH|11|2|ad reges quoque aquilonis qui habitabant in montanis et in planitie contra meridiem Cheneroth in campestribus quoque et in regionibus Dor iuxta mare
JOSH|11|3|Chananeumque ab oriente et occidente et Amorreum atque Hettheum ac Ferezeum et Iebuseum in montanis Eveum quoque qui habitabat ad radices Hermon in terra Masphe
JOSH|11|4|egressique sunt omnes cum turmis suis populus multus nimis sicut harena quae est in litore maris equi quoque et currus inmensae multitudinis
JOSH|11|5|conveneruntque omnes reges isti in unum ad aquas Merom ut pugnarent contra Israhel
JOSH|11|6|dixitque Dominus ad Iosue ne timeas eos cras enim hac eadem hora ego tradam omnes istos vulnerandos in conspectu Israhel equos eorum subnervabis et currus igne conbures
JOSH|11|7|venitque Iosue et omnis exercitus cum eo adversum illos ad aquas Merom subito et inruerunt super eos
JOSH|11|8|tradiditque illos Dominus in manu Israhel qui percusserunt eos et persecuti sunt usque ad Sidonem magnam et aquas Maserefoth campumque Masphe qui est ad orientalem illius partem ita percussit omnes ut nullas dimitteret ex eis reliquias
JOSH|11|9|fecit sicut praeceperat ei Dominus equos eorum subnervavit currusque conbusit
JOSH|11|10|reversusque statim cepit Asor et regem eius percussit gladio Asor enim antiquitus inter omnia regna haec principatum tenebat
JOSH|11|11|percussitque omnes animas quae ibidem morabantur non dimisit in ea ullas reliquias sed usque ad internicionem universa vastavit ipsamque urbem permisit incendio
JOSH|11|12|et omnes per circuitum civitates regesque earum cepit percussit atque delevit sicut praeceperat ei Moses famulus Domini
JOSH|11|13|absque urbibus quae erant in collibus et in tumulis sitae ceteras succendit Israhel unam tantum Asor munitissimam flamma consumpsit
JOSH|11|14|omnemque praedam istarum urbium ac iumenta diviserunt sibi filii Israhel cunctis hominibus interfectis
JOSH|11|15|sicut praeceperat Dominus Mosi servo suo ita praecepit Moses Iosue et ille universa conplevit non praeteriit de universis mandatis ne unum quidem verbum quod iusserat Dominus Mosi
JOSH|11|16|cepit itaque Iosue omnem terram montanam et meridianam terramque Gosen et planitiem et occidentalem plagam montemque Israhel et campestria eius
JOSH|11|17|et partem montis quae ascendit Seir usque Baalgad per planitiem Libani subter montem Hermon omnes reges eorum cepit percussit occidit
JOSH|11|18|multo tempore pugnavit Iosue contra reges istos
JOSH|11|19|non fuit civitas quae se non traderet filiis Israhel praeter Eveum qui habitabat in Gabaon omnes bellando cepit
JOSH|11|20|Domini enim sententiae fuerat ut indurarentur corda eorum et pugnarent contra Israhel et caderent et non mererentur ullam clementiam ac perirent sicut praeceperat Dominus Mosi
JOSH|11|21|in tempore illo venit Iosue et interfecit Enacim de montanis Hebron et Dabir et Anab et de omni monte Iuda et Israhel urbesque eorum delevit
JOSH|11|22|non reliquit ullum de stirpe Enacim in terra filiorum Israhel absque civitatibus Gaza et Geth et Azoto in quibus solis relicti sunt
JOSH|11|23|cepit ergo Iosue omnem terram sicut locutus est Dominus ad Mosen et tradidit eam in possessionem filiis Israhel secundum partes et tribus suas quievitque terra a proeliis
JOSH|12|1|hii sunt reges quos percusserunt filii Israhel et possederunt terram eorum trans Iordanem ad solis ortum a torrente Arnon usque ad montem Hermon et omnem orientalem plagam quae respicit solitudinem
JOSH|12|2|Seon rex Amorreorum qui habitavit in Esebon dominatus est ab Aroer quae sita est super ripam torrentis Arnon et mediae partis in valle dimidiique Galaad usque ad torrentem Iaboc qui est terminus filiorum Ammon
JOSH|12|3|et a solitudine usque ad mare Cheneroth contra orientem et usque ad mare Deserti quod est mare Salsissimum ad orientalem plagam per viam quae ducit Bethesimoth et ab australi parte quae subiacent Asedothphasga
JOSH|12|4|terminus Og regis Basan de reliquiis Rafaim qui habitavit in Astharoth et in Edrain et dominatus est in monte Hermon et in Salacha atque in universa Basan usque ad terminos
JOSH|12|5|Gesuri et Machathi et dimidiae partis Galaad terminos Seon regis Esebon
JOSH|12|6|Moses famulus Domini et filii Israhel percusserunt eos tradiditque terram eorum Moses in possessionem Rubenitis et Gadditis et dimidiae tribui Manasse
JOSH|12|7|hii sunt reges terrae quos percussit Iosue et filii Israhel trans Iordanem ad occidentalem plagam a Baalgad in campo Libani usque ad montem cuius pars ascendit in Seir tradiditque eam Iosue in possessionem tribubus Israhel singulis partes suas
JOSH|12|8|tam in montanis quam in planis atque campestribus in Aseroth et solitudine ac meridie Hettheus fuit et Amorreus Chananeus et Ferezeus Eveus et Iebuseus
JOSH|12|9|rex Hiericho unus rex Ahi quae est ex latere Bethel unus
JOSH|12|10|rex Hierusalem unus rex Hebron unus
JOSH|12|11|rex Hierimoth unus rex Lachis unus
JOSH|12|12|rex Eglon unus rex Gazer unus
JOSH|12|13|rex Dabir unus rex Gader unus
JOSH|12|14|rex Herma unus rex Hered unus
JOSH|12|15|rex Lebna unus rex Odollam unus
JOSH|12|16|rex Maceda unus rex Bethel unus
JOSH|12|17|rex Thaffua unus rex Afer unus
JOSH|12|18|rex Afec unus rex Saron unus
JOSH|12|19|rex Madon unus rex Asor unus
JOSH|12|20|rex Someron unus rex Acsaph unus
JOSH|12|21|rex Thenach unus rex Mageddo unus
JOSH|12|22|rex Cades unus rex Iachanaem Chermeli unus
JOSH|12|23|rex Dor et provinciae Dor unus rex gentium Galgal unus
JOSH|12|24|rex Thersa unus omnes reges triginta et unus
JOSH|13|1|Iosue senex provectaeque aetatis erat et dixit Dominus ad eum senuisti et longevus es terraque latissima derelicta est quae necdum est sorte divisa
JOSH|13|2|omnis videlicet Galilea Philisthim et universa Gesuri
JOSH|13|3|a fluvio turbido qui inrigat Aegyptum usque ad terminos Accaron contra aquilonem terra Chanaan quae in quinque regulos Philisthim dividitur Gazeos Azotios Ascalonitas Gettheos et Accaronitas
JOSH|13|4|ad meridiem vero sunt Evei omnis terra Chanaan et Maara Sidoniorum usque Afeca et terminos Amorrei
JOSH|13|5|eiusque confinia Libani quoque regio contra orientem a Baalgad sub monte Hermon donec ingrediaris Emath
JOSH|13|6|omnium qui habitant in monte a Libano usque ad aquas Masrefoth universique Sidonii ego sum qui delebo eos a facie filiorum Israhel veniat ergo in parte hereditatis Israhel sicut praecepi tibi
JOSH|13|7|et nunc divide terram in possessionem novem tribubus et dimidiae tribui Manasse
JOSH|13|8|cum qua Ruben et Gad possederunt terram quam tradidit eis Moses famulus Domini trans fluenta Iordanis ad orientalem plagam
JOSH|13|9|ab Aroer quae sita est in ripa torrentis Arnon et in vallis medio universaque campestria Medaba usque Dibon
JOSH|13|10|et cunctas civitates Seon regis Amorrei qui regnavit in Esebon usque ad terminos filiorum Ammon
JOSH|13|11|et Galaad ac terminum Gesuri et Machathi omnemque montem Hermon et universam Basan usque Saleca
JOSH|13|12|omne regnum Og in Basan qui regnavit in Astharoth et Edraim ipse fuit de reliquiis Rafaim percussitque eos Moses atque delevit
JOSH|13|13|nolueruntque disperdere filii Israhel Gesuri et Machathi et habitaverunt in medio Israhel usque in praesentem diem
JOSH|13|14|tribui autem Levi non dedit possessionem sed sacrificia et victimae Domini Dei Israhel ipsa est eius hereditas sicut locutus est illi
JOSH|13|15|dedit ergo Moses possessionem tribui filiorum Ruben iuxta cognationes suas
JOSH|13|16|fuitque terminus eorum ab Aroer quae sita est in ripa torrentis Arnon et in valle eiusdem torrentis media universam planitiem quae ducit Medaba
JOSH|13|17|et Esebon cunctosque viculos earum qui sunt in campestribus Dibon quoque et Bamothbaal et oppidum Baalmaon
JOSH|13|18|Iessa et Cedmoth et Mepheeth
JOSH|13|19|Cariathaim et Sebama et Sarathasar in monte convallis
JOSH|13|20|Bethpheor et Asedothphasga et Bethaisimoth
JOSH|13|21|omnes urbes campestres universaque regna Seon regis Amorrei qui regnavit in Esebon quem percussit Moses cum principibus Madian Eveum et Recem et Sur et Ur et Rabee duces Seon habitatores terrae
JOSH|13|22|et Balaam filium Beor ariolum occiderunt filii Israhel gladio cum ceteris interfectis
JOSH|13|23|factusque est terminus filiorum Ruben Iordanis fluvius haec est possessio Rubenitarum per cognationes suas urbium et viculorum
JOSH|13|24|deditque Moses tribui Gad et filiis eius per cognationes suas possessionem cuius haec divisio est
JOSH|13|25|terminus Iazer et omnes civitates Galaad dimidiamque partem terrae filiorum Ammon usque ad Aroer quae est contra Rabba
JOSH|13|26|et ab Esebon usque Ramoth Masphe et Batanim et a Manaim usque ad terminos Dabir
JOSH|13|27|in valle quoque Betharaam et Bethnemra et Soccoth et Saphon reliquam partem regni Seon regis Esebon huius quoque Iordanis finis est usque ad extremam partem maris Chenereth trans Iordanem ad orientalem plagam
JOSH|13|28|haec est possessio filiorum Gad per familias suas civitates et villae earum
JOSH|13|29|dedit et dimidiae tribui Manasse filiisque eius iuxta cognationes suas possessionem
JOSH|13|30|cuius hoc principium est a Manaim universam Basan et cuncta regna Og regis Basan omnesque vicos Air qui sunt in Basan sexaginta oppida
JOSH|13|31|et dimidiam partem Galaad Astharoth et Edrai urbes regni Og in Basan filiis Machir filii Manasse dimidiae parti filiorum Machir iuxta cognationes suas
JOSH|13|32|hanc possessionem divisit Moses in campestribus Moab trans Iordanem contra Hiericho ad orientalem plagam
JOSH|13|33|tribui autem Levi non dedit possessionem quoniam Dominus Deus Israhel ipse est possessio eius ut locutus est illi
JOSH|14|1|hoc est quod possederunt filii Israhel in terra Chanaan quam dederunt eis Eleazar sacerdos et Iosue filius Nun et principes familiarum per tribus Israhel
JOSH|14|2|sorte omnia dividentes sicut praeceperat Dominus in manu Mosi novem tribubus et dimidiae tribui
JOSH|14|3|duabus enim tribubus et dimidiae dederat Moses trans Iordanem possessionem absque Levitis qui nihil terrae acceperunt inter fratres suos
JOSH|14|4|sed in eorum successerant locum filii Ioseph in duas divisi tribus Manasse et Ephraim nec acceperunt Levitae aliam in terra partem nisi urbes ad habitandum et suburbana earum ad alenda iumenta et pecora sua
JOSH|14|5|sicut praecepit Dominus Mosi ita fecerunt filii Israhel et diviserunt terram
JOSH|14|6|accesserunt itaque filii Iuda ad Iosue in Galgala locutusque est ad eum Chaleb filius Iepphonne Cenezeus nosti quid locutus sit Dominus ad Mosen hominem Dei de me et te in Cadesbarne
JOSH|14|7|quadraginta annorum eram quando me misit Moses famulus Domini de Cadesbarne ut considerarem terram nuntiavique ei quod mihi verum videbatur
JOSH|14|8|fratres autem mei qui ascenderant mecum dissolverunt cor populi et nihilominus ego secutus sum Dominum Deum meum
JOSH|14|9|iuravitque Moses in die illo dicens terram quam calcavit pes tuus erit possessio tua et filiorum tuorum in aeternum quia secutus es Dominum Deum meum
JOSH|14|10|concessit ergo Dominus vitam mihi sicut pollicitus est usque in praesentem diem quadraginta et quinque anni sunt ex quo locutus est Dominus verbum istud ad Mosen quando ambulabat Israhel per solitudinem hodie octoginta quinque annorum sum
JOSH|14|11|sic valens ut eo valebam tempore quando ad explorandum missus sum illius in me temporis fortitudo usque hodie perseverat tam ad bellandum quam ad gradiendum
JOSH|14|12|da ergo mihi montem istum quem pollicitus est Dominus te quoque audiente in quo Enacim sunt et urbes magnae atque munitae si forte sit Dominus mecum et potuero delere eos sicut promisit mihi
JOSH|14|13|benedixitque ei Iosue et tradidit Hebron in possessionem
JOSH|14|14|atque ex eo fuit Hebron Chaleb filio Iepphonne Cenezeo usque in praesentem diem quia secutus est Dominum Deum Israhel
JOSH|14|15|nomen Hebron antea vocabatur Cariatharbe Adam maximus ibi inter Enacim situs est et terra cessavit a proeliis
JOSH|15|1|igitur sors filiorum Iudae per cognationes suas ista fuit a termino Edom desertum Sin contra meridiem et usque ad extremam partem australis plagae
JOSH|15|2|initium eius a summitate maris Salsissimi et a lingua eius quae respicit meridiem
JOSH|15|3|egrediturque contra ascensum Scorpionis et pertransit in Sina ascenditque in Cadesbarne et pervenit in Esrom ascendens Addara et circumiens Caricaa
JOSH|15|4|atque inde pertransiens in Asemona et perveniens ad torrentem Aegypti eruntque termini eius mare Magnum hic erit finis meridianae plagae
JOSH|15|5|ab oriente vero erit initium mare Salsissimum usque ad extrema Iordanis et ea quae respiciunt aquilonem a lingua maris usque ad eundem Iordanem fluvium
JOSH|15|6|ascenditque terminus in Bethagla et transit ab aquilone in Betharaba ascendens ad lapidem Boem filii Ruben
JOSH|15|7|et tendens usque ad terminos Debera de valle Achor contra aquilonem respiciens Galgala quae est ex adverso ascensionis Adommim ab australi parte torrentis transitque aquas quae vocantur fons Solis et erunt exitus eius ad fontem Rogel
JOSH|15|8|ascenditque per convallem filii Ennom ex latere Iebusei ad meridiem haec est Hierusalem et inde se erigens ad verticem montis qui est contra Gehennom ad occidentem in summitate vallis Rafaim contra aquilonem
JOSH|15|9|pertransitque a vertice montis usque ad fontem aquae Nepthoa et pervenit usque ad vicos montis Ephron inclinaturque in Bala quae est Cariathiarim id est urbs Silvarum
JOSH|15|10|et circuit de Bala contra occidentem usque ad montem Seir transitque iuxta latus montis Iarim ad aquilonem in Cheslon et descendit in Bethsames transitque in Thamna
JOSH|15|11|et pervenit contra aquilonem partis Accaron ex latere inclinaturque Sechrona et transit montem Baala pervenitque in Iebnehel et maris Magni contra occidentem fine concluditur
JOSH|15|12|hii sunt termini filiorum Iuda per circuitum in cognationibus suis
JOSH|15|13|Chaleb vero filio Iepphonne dedit partem in medio filiorum Iuda sicut praeceperat ei Dominus Cariatharbe patris Enach ipsa est Hebron
JOSH|15|14|delevitque ex ea Chaleb tres filios Enach Sesai et Ahiman et Tholmai de stirpe Enach
JOSH|15|15|atque inde conscendens venit ad habitatores Dabir quae prius vocabatur Cariathsepher id est civitas Litterarum
JOSH|15|16|dixitque Chaleb qui percusserit Cariathsepher et ceperit eam dabo illi Axam filiam meam uxorem
JOSH|15|17|cepitque eam Othonihel filius Cenez frater Chaleb iunior deditque ei Axam filiam suam uxorem
JOSH|15|18|quae cum pergerent simul suasit viro ut peteret a patre suo agrum suspiravitque ut sedebat in asino cui Chaleb quid habes inquit
JOSH|15|19|at illa respondit da mihi benedictionem terram australem et arentem dedisti mihi iunge et inriguam dedit itaque ei Chaleb inriguum superius et inferius
JOSH|15|20|haec est possessio tribus filiorum Iuda per cognationes suas
JOSH|15|21|erantque civitates ab extremis partibus filiorum Iuda iuxta terminos Edom a meridie Cabsehel et Eder et Iagur
JOSH|15|22|et Cina et Dimona Adeda
JOSH|15|23|et Cedes et Asor Iethnan
JOSH|15|24|Zif et Thelem Baloth
JOSH|15|25|et Asor nova et Cariothesrom haec est Asor
JOSH|15|26|Aman Same et Molada
JOSH|15|27|et Asergadda et Asemon Bethfeleth
JOSH|15|28|et Asersual et Bersabee et Baziothia
JOSH|15|29|Bala et Hiim Esem
JOSH|15|30|et Heltholad Exiil et Harma
JOSH|15|31|Siceleg et Medemena et Sensenna
JOSH|15|32|Lebaoth et Selim et Aenremmon omnes civitates viginti novem et villae earum
JOSH|15|33|in campestribus vero Esthaul et Saraa et Asena
JOSH|15|34|et Azanoe et Aengannim Thaffua et Aenaim
JOSH|15|35|et Hierimoth Adulam Soccho et Azeca
JOSH|15|36|et Saraim Adithaim et Gedera et Giderothaim urbes quattuordecim et villae earum
JOSH|15|37|Sanan et Adesa et Magdalgad
JOSH|15|38|Delean et Mesfa et Iecthel
JOSH|15|39|Lachis et Bascath et Aglon
JOSH|15|40|Thebbon et Lehemas et Chethlis
JOSH|15|41|et Gideroth Bethdagon et Neema et Maceda civitates sedecim et villae earum
JOSH|15|42|Labana et Aether et Asan
JOSH|15|43|Ieptha et Esna et Nesib
JOSH|15|44|Ceila et Achzib et Maresa civitates novem et villae earum
JOSH|15|45|Accaron cum vicis et villulis suis
JOSH|15|46|ab Accaron usque ad mare omnia quae vergunt ad Azotum et viculos eius
JOSH|15|47|Azotus cum vicis et villulis suis Gaza cum viculis et villulis suis usque ad torrentem Aegypti mare Magnum terminus eius
JOSH|15|48|et in monte Samir et Iether et Soccho
JOSH|15|49|et Edenna Cariathsenna haec est Dabir
JOSH|15|50|Anab et Isthemo et Anim
JOSH|15|51|Gosen et Olon et Gilo civitates undecim et villae earum
JOSH|15|52|Arab et Roma et Esaan
JOSH|15|53|Ianum et Bethafua et Afeca
JOSH|15|54|Ammatha et Cariatharbe haec est Hebron et Sior civitates novem et villae earum
JOSH|15|55|Maon et Chermel et Zif et Iotae
JOSH|15|56|Iezrehel et Iucadam et Zanoe
JOSH|15|57|Accaim Gebaa et Thamna civitates decem et villae earum
JOSH|15|58|Alul et Bethsur et Gedor
JOSH|15|59|Mareth et Bethanoth et Elthecen civitates sex et villae earum
JOSH|15|60|Cariathbaal haec est Cariathiarim urbs Silvarum et Arebba civitates duae et villae earum
JOSH|15|61|in deserto Betharaba Meddin et Schacha
JOSH|15|62|Anepsan et civitas Salis et Engaddi civitates sex et villae earum
JOSH|15|63|Iebuseum autem habitatorem Hierusalem non potuerunt filii Iuda delere habitavitque Iebuseus cum filiis Iuda in Hierusalem usque in praesentem diem
JOSH|16|1|cecidit quoque sors filiorum Ioseph ab Iordane contra Hiericho et aquas eius ab oriente solitudo quae ascendit de Hiericho ad montana Bethel
JOSH|16|2|et egreditur de Bethel Luzam transitque terminum Archiatharoth
JOSH|16|3|et descendit ad occidentem iuxta terminum Ieflethi usque ad terminos Bethoron inferioris et Gazer finiunturque regiones eius mari Magno
JOSH|16|4|possederuntque filii Ioseph Manasse et Ephraim
JOSH|16|5|et factus est terminus filiorum Ephraim per cognationes suas et possessio eorum contra orientem Atharothaddar usque Bethoron superiorem
JOSH|16|6|egrediunturque confinia in mare Machmethath vero aquilonem respicit et circuit terminus contra orientem in Thanathselo et pertransit ab oriente Ianoe
JOSH|16|7|descenditque de Ianoe in Atharoth et Noaratha et pervenit in Hiericho et egreditur ad Iordanem
JOSH|16|8|de Taffua pertransitque contra mare in valle Harundineti suntque egressus eius in mare Salsissimum haec est possessio tribus filiorum Ephraim per familias suas
JOSH|16|9|urbesque quae separatae sunt filiis Ephraim in medio possessionis filiorum Manasse et villae earum
JOSH|16|10|et non interfecerunt filii Ephraim Chananeum qui habitabat in Gazer habitavitque Chananeus in medio Ephraim usque in diem hanc tributarius
JOSH|17|1|cecidit autem sors tribui Manasse ipse est enim primogenitus Ioseph Machir primogenito Manasse patri Galaad qui fuit vir pugnator habuitque possessionem Galaad et Basan
JOSH|17|2|et reliquis filiorum Manasse iuxta familias suas filiis Abiezer et filiis Elech et filiis Esrihel et filiis Sechem et filiis Epher et filiis Semida isti sunt filii Manasse filii Ioseph mares per cognationes suas
JOSH|17|3|Salphaad vero filio Epher filii Galaad filii Machir filii Manasse non erant filii sed solae filiae quarum ista sunt nomina Maala et Noa Egla et Melcha et Thersa
JOSH|17|4|veneruntque in conspectu Eleazari sacerdotis et Iosue filii Nun et principum dicentes Dominus praecepit per manum Mosi ut daretur nobis possessio in medio fratrum nostrorum deditque eis iuxta imperium Domini possessionem in medio fratrum patris earum
JOSH|17|5|et ceciderunt funiculi Manasse decem absque terra Galaad et Basan trans Iordanem
JOSH|17|6|filiae enim Manasse possederunt hereditatem in medio filiorum eius terra autem Galaad cecidit in sortem filiorum Manasse qui reliqui erant
JOSH|17|7|fuitque terminus Manasse ab Aser Machmathath quae respicit Sychem et egreditur ad dextram iuxta habitatores fontis Taffuae
JOSH|17|8|etenim in sorte Manasse ceciderat terra Taffuae quae est iuxta terminos Manasse filiorum Ephraim
JOSH|17|9|descenditque terminus vallis Harundineti in meridiem torrentis civitatum Ephraim quae in medio sunt urbium Manasse terminus Manasse ab aquilone torrentis et exitus eius pergit ad mare
JOSH|17|10|ita ut ab austro sit possessio Ephraim et ab aquilone Manasse et utramque claudat mare et coniungantur sibi in tribu Aser ab aquilone et in tribu Isachar ab oriente
JOSH|17|11|fuitque hereditas Manasse in Isachar et in Aser Bethsan et viculi eius et Ieblaam cum villulis suis et habitatores Dor cum oppidis suis habitatores quoque Hendor cum villulis suis similiterque habitatores Thanach cum villulis suis et habitatores Mageddo cum viculis suis et tertia pars urbis Nofeth
JOSH|17|12|nec potuerunt filii Manasse has subvertere civitates sed coepit Chananeus habitare in terra ista
JOSH|17|13|postquam autem convaluerunt filii Israhel subiecerunt Chananeos et fecerunt sibi tributarios nec interfecerunt eos
JOSH|17|14|locutique sunt filii Ioseph ad Iosue atque dixerunt quare dedisti mihi possessionem sortis et funiculi unius cum sim tantae multitudinis et benedixerit mihi Dominus
JOSH|17|15|ad quos Iosue ait si populus multus es ascende in silvam et succide tibi spatia in terra Ferezei et Rafaim quia angusta est tibi possessio montis Ephraim
JOSH|17|16|cui responderunt filii Ioseph non poterimus ad montana conscendere cum ferreis curribus utantur Chananei qui habitant in terra campestri in qua sitae sunt Bethsan cum viculis suis et Iezrahel mediam possidens vallem
JOSH|17|17|dixitque Iosue ad domum Ioseph Ephraim et Manasse populus multus es et magnae fortitudinis non habebis sortem unam
JOSH|17|18|sed transibis ad montem et succides tibi atque purgabis ad habitandum spatia et poteris ultra procedere cum subverteris Chananeum quem dicis ferreos habere currus et esse fortissimum
JOSH|18|1|congregatique sunt omnes filii Israhel in Silo ibique fixerunt tabernaculum testimonii et fuit eis terra subiecta
JOSH|18|2|remanserant autem filiorum Israhel septem tribus quae necdum acceperant possessiones suas
JOSH|18|3|ad quos Iosue ait usquequo marcetis ignavia et non intratis ad possidendam terram quam Dominus Deus patrum vestrorum dedit vobis
JOSH|18|4|eligite de singulis tribubus ternos viros ut mittam eos et pergant atque circumeant terram et describant eam iuxta numerum uniuscuiusque multitudinis referantque ad me quod descripserint
JOSH|18|5|dividite vobis terram in septem partes Iudas sit in terminis suis ab australi plaga et domus Ioseph ab aquilone
JOSH|18|6|mediam inter hos terram in septem partes describite et huc venietis ad me ut coram Domino Deo vestro mittam vobis hic sortem
JOSH|18|7|quia non est inter vos pars Levitarum sed sacerdotium Domini est eorum hereditas Gad autem et Ruben et dimidia tribus Manasse iam acceperant possessiones suas trans Iordanem ad orientalem plagam quas dedit eis Moses famulus Domini
JOSH|18|8|cumque surrexissent viri ut pergerent ad describendam terram praecepit eis Iosue dicens circuite terram et describite eam ac revertimini ad me ut hic coram Domino Deo in Silo mittam vobis sortem
JOSH|18|9|itaque perrexerunt et lustrantes eam in septem partes diviserunt scribentes in volumine reversique sunt ad Iosue in castra Silo
JOSH|18|10|qui misit sortes coram Domino in Silo divisitque terram filiis Israhel in septem partes
JOSH|18|11|et ascendit sors prima filiorum Beniamin per familias suas ut possiderent terram inter filios Iuda et filios Ioseph
JOSH|18|12|fuitque terminus eorum contra aquilonem ab Iordane pergens iuxta latus Hiericho septentrionalis plagae et inde contra occidentem ad montana conscendens et perveniens in solitudinem Bethaven
JOSH|18|13|atque pertransiens iuxta Luzam ad meridiem ipsa est Bethel descenditque in Atharothaddar in montem qui est ad meridiem Bethoron inferioris
JOSH|18|14|et inclinatur circumiens contra mare a meridie montis qui respicit Bethoron contra africum suntque exitus eius in Cariathbaal quae vocatur et Cariathiarim urbem filiorum Iuda haec est plaga contra mare et occidentem
JOSH|18|15|a meridie autem ex parte Cariathiarim egreditur terminus contra mare et pervenit usque ad fontem aquarum Nepthoa
JOSH|18|16|descenditque in partem montis qui respicit vallem filiorum Ennom et est contra septentrionalem plagam in extrema parte vallis Rafaim descenditque Gehennom id est vallis Ennom iuxta latus Iebusei ad austrum et pervenit ad fontem Rogel
JOSH|18|17|transiens ad aquilonem et egrediens ad Aensemes id est fontem Solis
JOSH|18|18|et pertransit usque ad tumulos qui sunt e regione ascensus Adommim descenditque ad Abenboen id est lapidem Boen filii Ruben et pertransit ex latere aquilonis ad campestria descenditque in planitiem
JOSH|18|19|et praetergreditur contra aquilonem Bethagla suntque exitus eius contra linguam maris Salsissimi ab aquilone in fine Iordanis ad australem plagam
JOSH|18|20|qui est terminus illius ab oriente haec est possessio filiorum Beniamin per terminos suos in circuitu et familias singulas
JOSH|18|21|fueruntque civitates eius Hiericho et Bethagla et vallis Casis
JOSH|18|22|Betharaba et Semaraim et Bethel
JOSH|18|23|Avim et Affara et Ofra
JOSH|18|24|villa Emona et Ofni et Gabee civitates duodecim et villae earum
JOSH|18|25|Gabaon et Rama et Beroth
JOSH|18|26|et Mesfe Cafera et Ammosa
JOSH|18|27|et Recem Iarafel et Tharala
JOSH|18|28|et Sela Eleph et Iebus quae est Hierusalem Gabaath et Cariath civitates quattuordecim et villae earum haec est possessio filiorum Beniamin iuxta familias suas
JOSH|19|1|et egressa est sors secunda filiorum Symeon per cognationes suas fuitque hereditas
JOSH|19|2|eorum in medio possessionis filiorum Iuda Bersabee et Sabee et Molada
JOSH|19|3|et Asersual Bala et Asem
JOSH|19|4|et Heltholath Bethul Arma
JOSH|19|5|et Seceleg et Bethmarchaboth Asersusa
JOSH|19|6|et Bethlebaoth et Saroen civitates tredecim et villae earum
JOSH|19|7|Ahin et Remmon et Athar et Asan civitates quattuor et villae earum
JOSH|19|8|omnes viculi per circuitum urbium istarum usque ad Balaath Berrameth contra australem plagam haec est hereditas filiorum Symeon iuxta cognationes suas
JOSH|19|9|in funiculo et possessione filiorum Iuda quia maior erat et idcirco possederunt filii Symeon in medio hereditatis eorum
JOSH|19|10|cecidit quoque sors tertia filiorum Zabulon per cognationes suas et factus est terminus possessionis eorum usque Sarith
JOSH|19|11|ascenditque de mari et Medala ac pervenit in Debbaseth usque ad torrentem qui est contra Iecennam
JOSH|19|12|et revertitur de Sarith contra orientem in fines Ceseleththabor et egreditur ad Dabereth ascenditque contra Iafie
JOSH|19|13|et inde pertransit ad orientalem plagam Getthefer Etthacasin et egreditur in Remmon Ampthar et Noa
JOSH|19|14|et circuit ad aquilonem et Nathon suntque egressus eius vallis Iepthahel
JOSH|19|15|et Catheth et Nehalal et Semron et Iedala et Bethleem civitates duodecim et villae earum
JOSH|19|16|haec est hereditas tribus filiorum Zabulon per cognationes suas urbes et viculi earum
JOSH|19|17|Isachar egressa est sors quarta per cognationes suas
JOSH|19|18|fuitque eius hereditas Hiezrahel et Chasaloth et Sunem
JOSH|19|19|et Afaraim Seon et Anaarath
JOSH|19|20|et Rabbith et Cesion Abes
JOSH|19|21|et Rameth et Engannim et Enadda et Bethfeses
JOSH|19|22|et pervenit terminus usque Thabor et Seesima et Bethsemes eruntque exitus eius Iordanes civitates sedecim et villae earum
JOSH|19|23|haec est possessio filiorum Isachar per cognationes suas urbes et viculi earum
JOSH|19|24|cecidit sors quinta tribui filiorum Aser per cognationes suas
JOSH|19|25|fuitque terminus eorum Alchath et Oali et Beten et Axab
JOSH|19|26|Elmelech et Amaad et Messal et pervenit usque ad Carmelum maris et Siorlabanath
JOSH|19|27|ac revertitur contra orientem Bethdagon et pertransit usque Zabulon et vallem Iepthahel contra aquilonem in Bethemech et Neihel egrediturque ad levam Chabul
JOSH|19|28|et Achran et Roob et Amon et Canae usque ad Sidonem magnam
JOSH|19|29|revertiturque in Orma usque ad civitatem munitissimam Tyrum et usque Osa eruntque exitus eius in mare de funiculo Acziba
JOSH|19|30|et Amma et Afec et Roob civitates viginti duae et villae earum
JOSH|19|31|haec est possessio filiorum Aser per cognationes suas urbes et viculi earum
JOSH|19|32|filiorum Nepthalim sexta pars cecidit per familias suas
JOSH|19|33|et coepit terminus de Heleb et Helon in Sananim et Adami quae est Neceb et Iebnahel usque Lecum et egressus eorum usque ad Iordanem
JOSH|19|34|revertiturque terminus contra occidentem in Aznoththabor atque inde egreditur in Ucoca et pertransit in Zabulon contra meridiem et in Aser contra occidentem et in Iuda ad Iordanem contra ortum solis
JOSH|19|35|civitates munitissimae Aseddim Ser et Ammath et Recchath Chenereth
JOSH|19|36|et Edema et Arama Asor
JOSH|19|37|et Cedes et Edrai Nasor
JOSH|19|38|et Ieron et Magdalel Horem et Bethanath et Bethsemes civitates decem et novem et villae earum
JOSH|19|39|haec est possessio tribus filiorum Nepthali per cognationes suas urbes et viculi earum
JOSH|19|40|tribui filiorum Dan per familias suas egressa est sors septima
JOSH|19|41|et fuit terminus possessionis eius Saraa et Esthaol et Ahirsemes id est civitas Solis
JOSH|19|42|Selebin et Ahialon et Iethela
JOSH|19|43|Helon et Themna et Acron
JOSH|19|44|Helthecen et Gebthon et Baalath
JOSH|19|45|Iud et Benebarach et Gethremmon
JOSH|19|46|aquae Hiercon et Areccon cum termino qui respicit Ioppen
JOSH|19|47|et ipso fine concluditur ascenderuntque filii Dan et pugnaverunt contra Lesem ceperuntque eam et percusserunt in ore gladii ac possederunt et habitaverunt in ea vocantes nomen eius Lesemdan ex nomine Dan patris sui
JOSH|19|48|haec est possessio tribus filiorum Dan per cognationes suas urbes et viculi earum
JOSH|19|49|cumque conplesset terram sorte dividere singulis per tribus suas dederunt filii Israhel possessionem Iosue filio Nun in medio sui
JOSH|19|50|iuxta praeceptum Domini urbem quam postulavit Thamnathseraa in monte Ephraim et aedificavit civitatem habitavitque in ea
JOSH|19|51|hae sunt possessiones quas sorte diviserunt Eleazar sacerdos et Iosue filius Nun et principes familiarum ac tribuum filiorum Israhel in Silo coram Domino ad ostium tabernaculi testimonii partitique sunt terram
JOSH|20|1|et locutus est Dominus ad Iosue dicens loquere filiis Israhel et dic eis
JOSH|20|2|separate urbes fugitivorum de quibus locutus sum ad vos per manum Mosi
JOSH|20|3|ut confugiat ad eas quicumque animam percusserit nescius et possit evadere iram proximi qui ultor est sanguinis
JOSH|20|4|cum ad unam harum confugerit civitatum stabitque ante portam civitatis et loquetur senioribus urbis illius ea quae se conprobent innocentem sicque suscipient eum et dabunt ei locum ad habitandum
JOSH|20|5|cumque ultor sanguinis eum fuerit persecutus non tradent in manus eius quia ignorans percussit proximum eius nec ante biduum triduumve eius probatur inimicus
JOSH|20|6|et habitabit in civitate illa donec stet ante iudicium causam reddens facti sui et moriatur sacerdos magnus qui fuerit in illo tempore tunc revertetur homicida et ingredietur civitatem et domum suam de qua fugerat
JOSH|20|7|decreveruntque Cedes in Galilea montis Nepthali et Sychem in monte Ephraim et Cariatharbe ipsa est Hebron in monte Iuda
JOSH|20|8|et trans Iordanem contra orientalem plagam Hiericho statuerunt Bosor quae sita est in campestri solitudine de tribu Ruben et Ramoth in Galaad de tribu Gad et Gaulon in Basan de tribu Manasse
JOSH|20|9|hae civitates constitutae sunt cunctis filiis Israhel et advenis qui habitant inter eos ut fugeret ad eas qui animam nescius percussisset et non moreretur in manu proximi effusum sanguinem vindicare cupientis donec staret ante populum expositurus causam suam
JOSH|21|1|accesseruntque principes familiarum Levi ad Eleazar sacerdotem et Iosue filium Nun et ad duces cognationum per singulas tribus filiorum Israhel
JOSH|21|2|locutique sunt ad eos in Silo terrae Chanaan atque dixerunt Dominus praecepit per manum Mosi ut darentur nobis urbes ad habitandum et suburbana earum ad alenda iumenta
JOSH|21|3|dederuntque filii Israhel de possessionibus suis iuxta imperium Domini civitates et suburbana earum
JOSH|21|4|egressaque est sors in familiam Caath filiorum Aaron sacerdotis de tribubus Iuda et Symeon et Beniamin civitates tredecim
JOSH|21|5|et reliquis filiorum Caath id est Levitis qui superflui erant de tribubus Ephraim et Dan et dimidia tribu Manasse civitates decem
JOSH|21|6|porro filiis Gerson egressa est sors ut acciperent de tribubus Isachar et Aser et Nepthalim dimidiaque tribu Manasse in Basan civitates numero tredecim
JOSH|21|7|et filiis Merari per cognationes suas de tribubus Ruben et Gad et Zabulon urbes duodecim
JOSH|21|8|dederuntque filii Israhel Levitis civitates et suburbana earum sicut praecepit Dominus per manum Mosi singulis sorte tribuentes
JOSH|21|9|de tribubus filiorum Iuda et Symeon dedit Iosue civitates quarum ista sunt nomina
JOSH|21|10|filiis Aaron per familias Caath levitici generis prima enim sors illis egressa est
JOSH|21|11|Cariatharbe patris Enach quae vocatur Hebron in monte Iuda et suburbana eius per circuitum
JOSH|21|12|agros vero et villas eius dederat Chaleb filio Iepphonne ad possidendum
JOSH|21|13|dedit ergo filiis Aaron sacerdotis Hebron confugii civitatem ac suburbana eius et Lebnam cum suburbanis suis
JOSH|21|14|et Iether et Isthimon
JOSH|21|15|et Helon Dabir
JOSH|21|16|et Ahin et Iethan et Bethsemes cum suburbanis suis civitates novem de tribubus ut dictum est duabus
JOSH|21|17|de tribu autem filiorum Beniamin Gabaon et Gabee
JOSH|21|18|et Anathoth et Almon cum suburbanis suis civitates quattuor
JOSH|21|19|omnes simul civitates filiorum Aaron sacerdotis tredecim cum suburbanis suis
JOSH|21|20|reliquis vero per familias filiorum Caath levitici generis haec est data possessio
JOSH|21|21|de tribu Ephraim urbs confugii Sychem cum suburbanis suis in monte Ephraim et Gazer
JOSH|21|22|et Cebsain et Bethoron cum suburbanis suis civitates quattuor
JOSH|21|23|de tribu quoque Dan Elthece et Gebbethon
JOSH|21|24|et Ahialon et Gethremmon cum suburbanis suis civitates quattuor
JOSH|21|25|porro de dimidia tribu Manasse Thanach et Gethremmon cum suburbanis suis civitates duae
JOSH|21|26|omnes civitates decem et suburbana earum datae sunt filiis Caath inferioris gradus
JOSH|21|27|filiis quoque Gerson levitici generis dedit de dimidia tribu Manasse confugii civitatem Gaulon in Basan et Bosram cum suburbanis suis civitates duas
JOSH|21|28|porro de tribu Isachar Cesion et Dabereth
JOSH|21|29|et Iaramoth et Engannim cum suburbanis suis civitates quattuor
JOSH|21|30|de tribu autem Aser Masal et Abdon
JOSH|21|31|et Elacoth et Roob cum suburbanis suis civitates quattuor
JOSH|21|32|de tribu quoque Nepthali civitatem confugii Cedes in Galilea et Ammothdor et Charthan cum suburbanis suis civitates tres
JOSH|21|33|omnes urbes familiarum Gerson tredecim cum suburbanis suis
JOSH|21|34|filiis autem Merari Levitis inferioris gradus per familias suas data est de tribu Zabulon Iechenam et Chartha
JOSH|21|35|et Damna et Nalol civitates quattuor cum suburbanis suis
JOSH|21|36|de tribu quoque Ruben ciuitates confugii Bosor in solitudine et Cedson et Misor et Ocho ciuitates quattuor cum suburbanis suis]
JOSH|21|37|et de tribu Gad civitates confugii Ramoth in Galaad et Manaim et Esebon et Iazer civitates quattuor cum suburbanis suis
JOSH|21|38|omnes urbes filiorum Merari per familias et cognationes suas duodecim
JOSH|21|39|itaque universae civitates Levitarum in medio possessionis filiorum Israhel fuerunt quadraginta octo
JOSH|21|40|cum suburbanis suis singulae per familias distributae
JOSH|21|41|deditque Dominus Israheli omnem terram quam traditurum se patribus eorum iuraverat et possederunt illam atque habitaverunt in ea
JOSH|21|42|dataque est ab eo pax in omnes per circuitum nationes nullusque eis hostium resistere ausus est sed cuncti in eorum dicionem redacti sunt
JOSH|21|43|ne unum quidem verbum quod illis praestaturum se esse promiserat irritum fuit sed rebus expleta sunt omnia
JOSH|22|1|eodem tempore vocavit Iosue Rubenitas et Gadditas et dimidiam tribum Manasse
JOSH|22|2|dixitque ad eos fecistis omnia quae vobis praecepit Moses famulus Domini mihi quoque in omnibus oboedistis
JOSH|22|3|nec reliquistis fratres vestros longo tempore usque in praesentem diem custodientes imperium Domini Dei vestri
JOSH|22|4|quia igitur dedit Dominus Deus vester fratribus vestris quietem ac pacem sicut pollicitus est revertimini et ite in tabernacula vestra et in terram possessionis quam tradidit vobis Moses famulus Domini trans Iordanem
JOSH|22|5|ita dumtaxat ut custodiatis adtente et opere conpleatis mandatum et legem quam praecepit vobis Moses servus Domini ut diligatis Dominum Deum vestrum et ambuletis in omnibus viis eius et observetis mandata illius adhereatisque ei ac serviatis in omni corde et in omni anima vestra
JOSH|22|6|benedixitque eis Iosue et dimisit eos qui reversi sunt in tabernacula sua
JOSH|22|7|tribui autem Manasse mediae possessionem Moses dederat in Basan et idcirco mediae quae superfuit dedit Iosue sortem inter ceteros fratres suos trans Iordanem ad occidentalem eius plagam cumque dimitteret eos in tabernacula sua et benedixisset illis
JOSH|22|8|dixit ad eos in multa substantia atque divitiis revertimini ad sedes vestras cum argento et auro aere ac ferro et veste multiplici dividite praedam hostium cum fratribus vestris
JOSH|22|9|reversique sunt et abierunt filii Ruben et filii Gad et dimidia tribus Manasse a filiis Israhel de Silo quae sita est in Chanaan ut intrarent Galaad terram possessionis suae quam obtinuerant iuxta imperium Domini in manu Mosi
JOSH|22|10|cumque venissent ad tumulos Iordanis in terra Chanaan aedificaverunt iuxta Iordanem altare infinitae magnitudinis
JOSH|22|11|quod cum audissent filii Israhel et ad eos certi nuntii detulissent aedificasse filios Ruben et Gad et dimidiae tribus Manasse altare in terra Chanaan super Iordanis tumulos contra filios Israhel
JOSH|22|12|convenerunt omnes in Silo ut ascenderent et dimicarent contra eos
JOSH|22|13|et interim miserunt ad illos in terram Galaad Finees filium Eleazar sacerdotem
JOSH|22|14|et decem principes cum eo singulos de tribubus singulis
JOSH|22|15|qui venerunt ad filios Ruben et Gad et dimidiae tribus Manasse in terram Galaad dixeruntque ad eos
JOSH|22|16|haec mandat omnis populus Domini quae est ista transgressio cur reliquistis Dominum Deum Israhel aedificantes altare sacrilegum et a cultu illius recedentes
JOSH|22|17|an parum vobis est quod peccastis in Beelphegor et usque in praesentem diem macula huius sceleris in nobis permanet multique de populo corruerunt
JOSH|22|18|et vos hodie reliquistis Dominum et cras in universum Israhel eius ira desaeviet
JOSH|22|19|quod si putatis inmundam esse terram possessionis vestrae transite ad terram in qua tabernaculum Domini est et habitate inter nos tantum ut a Domino et a nostro consortio non recedatis aedificato altari praeter altare Domini Dei vestri
JOSH|22|20|nonne Achan filius Zare praeteriit mandatum Domini et super omnem populum Israhel ira eius incubuit et ille erat unus homo atque utinam solus perisset in scelere suo
JOSH|22|21|responderuntque filii Ruben et Gad et dimidiae tribus Manasse principibus legationis Israhel
JOSH|22|22|fortissimus Deus Dominus fortissimus Deus Dominus ipse novit et Israhel simul intelleget si praevaricationis animo hoc altare construximus non custodiat nos sed puniat in praesenti
JOSH|22|23|et si ea mente fecimus ut holocausta et sacrificium et pacificas victimas super eo inponeremus ipse quaerat et iudicet
JOSH|22|24|et non ea magis cogitatione atque tractatu ut diceremus cras dicent filii vestri filiis nostris quid vobis et Domino Deo Israhel
JOSH|22|25|terminum posuit Dominus inter nos et vos o filii Ruben et filii Gad Iordanem fluvium et idcirco partem non habetis in Domino et per hanc occasionem avertent filii vestri filios nostros a timore Domini putavimus itaque melius
JOSH|22|26|et diximus extruamus nobis altare non in holocausta neque ad victimas offerendas
JOSH|22|27|sed in testimonium inter nos et vos et subolem nostram vestramque progeniem ut serviamus Domino et iuris nostri sit offerre holocausta et victimas et pacificas hostias et nequaquam dicant cras filii vestri filiis nostris non est vobis pars in Domino
JOSH|22|28|quod si voluerint dicere respondebunt eis ecce altare Domini quod fecerunt patres nostri non in holocausta neque in sacrificium sed in testimonium vestrum ac nostrum
JOSH|22|29|absit a nobis hoc scelus ut recedamus a Domino et eius vestigia relinquamus extructo altari ad holocausta et sacrificia et victimas offerendas praeter altare Domini Dei nostri quod extructum est ante tabernaculum eius
JOSH|22|30|quibus auditis Finees sacerdos et principes legationis Israhel qui erant cum eo placati sunt et verba filiorum Ruben et Gad et dimidiae tribus Manasse libentissime susceperunt
JOSH|22|31|dixitque Finees filius Eleazari sacerdos ad eos nunc scimus quod nobiscum sit Dominus quoniam alieni estis a praevaricatione hac et liberastis filios Israhel de manu Domini
JOSH|22|32|reversusque est cum principibus a filiis Ruben et Gad de terra Galaad finium Chanaan ad filios Israhel et rettulit eis
JOSH|22|33|placuitque sermo cunctis audientibus et laudaverunt Deum filii Israhel et nequaquam ultra dixerunt ut ascenderent contra eos atque pugnarent et delerent terram possessionis eorum
JOSH|22|34|vocaveruntque filii Ruben et filii Gad altare quod extruxerant Testimonium nostrum quod Dominus ipse sit Deus
JOSH|23|1|evoluto autem multo tempore postquam pacem Dominus dederat Israheli subiectis in gyro nationibus universis et Iosue iam longevo et persenilis aetatis
JOSH|23|2|vocavit Iosue omnem Israhelem maioresque natu et principes ac duces et magistros dixitque ad eos ego senui et progressioris aetatis sum
JOSH|23|3|vosque cernitis omnia quae fecerit Dominus Deus vester cunctis per circuitum nationibus quomodo pro vobis ipse pugnaverit
JOSH|23|4|et nunc quia vobis sorte divisit omnem terram ab orientali parte Iordanis usque ad mare Magnum multaeque adhuc supersunt nationes
JOSH|23|5|Dominus Deus vester disperdet eas et auferet a facie vestra et possidebitis terram sicut vobis pollicitus est
JOSH|23|6|tantum confortamini et estote solliciti ut custodiatis cuncta quae scripta sunt in volumine legis Mosi et non declinetis ab eis nec ad dextram nec ad sinistram
JOSH|23|7|ne postquam intraveritis ad gentes quae inter vos futurae sunt iuretis in nomine deorum earum et serviatis eis et adoretis illos
JOSH|23|8|sed adhereatis Domino Deo vestro quod fecistis usque in diem hanc
JOSH|23|9|et tunc auferet Dominus in conspectu vestro gentes magnas et robustissimas et nullus vobis resistere poterit
JOSH|23|10|unus e vobis persequetur hostium mille viros quia Dominus Deus vester pro vobis ipse pugnabit sicut pollicitus est
JOSH|23|11|hoc tantum diligentissime praecavete ut diligatis Dominum Deum vestrum
JOSH|23|12|quod si volueritis gentium harum quae inter vos habitant erroribus adherere et cum eis miscere conubia atque amicitias copulare
JOSH|23|13|iam nunc scitote quod Dominus Deus vester non eas deleat ante faciem vestram sed sint vobis in foveam ac laqueum et offendiculum ex latere vestro et sudes in oculis vestris donec vos auferat atque disperdat de terra hac optima quam tradidit vobis
JOSH|23|14|en ego hodie ingrediar viam universae terrae et toto animo cognoscetis quod de omnibus verbis quae se Dominus praestaturum nobis esse pollicitus est unum non praeterierit in cassum
JOSH|23|15|sicut ergo implevit opere quod promisit et prospera cuncta venerunt sic adducet super vos quicquid malorum comminatus est donec vos auferat atque disperdat de terra hac optima quam tradidit vobis
JOSH|23|16|eo quod praeterieritis pactum Domini Dei vestri quod pepigit vobiscum et servieritis diis alienis et adoraveritis eos cito atque velociter consurget in vos furor Domini et auferemini de terra hac optima quam tradidit vobis
JOSH|24|1|congregavitque Iosue omnes tribus Israhel in Sychem et vocavit maiores natu ac principes et iudices et magistros steteruntque in conspectu Domini
JOSH|24|2|et ad populum sic locutus est haec dicit Dominus Deus Israhel trans fluvium habitaverunt patres vestri ab initio Thare pater Abraham et Nahor servieruntque diis alienis
JOSH|24|3|tuli ergo patrem vestrum Abraham de Mesopotamiae finibus et adduxi eum in terram Chanaan multiplicavique semen eius
JOSH|24|4|et dedi ei Isaac illique rursum dedi Iacob et Esau e quibus Esau dedi montem Seir ad possidendum Iacob vero et filii eius descenderunt in Aegyptum
JOSH|24|5|misique Mosen et Aaron et percussi Aegyptum multis signis atque portentis
JOSH|24|6|eduxique vos et patres vestros de Aegypto et venistis ad mare persecutique sunt Aegyptii patres vestros cum curribus et equitatu usque ad mare Rubrum
JOSH|24|7|clamaverunt autem ad Dominum filii Israhel qui posuit tenebras inter vos et Aegyptios et adduxit super eos mare et operuit illos viderunt oculi vestri cuncta quae in Aegypto fecerim et habitastis in solitudine multo tempore
JOSH|24|8|et introduxi vos ad terram Amorrei qui habitabat trans Iordanem cumque pugnarent contra vos tradidi eos in manus vestras et possedistis terram eorum atque interfecistis illos
JOSH|24|9|surrexit autem Balac filius Sepphor rex Moab et pugnavit contra Israhelem misitque et vocavit Balaam filium Beor ut malediceret vobis
JOSH|24|10|et ego nolui audire eum sed e contrario per illum benedixi vobis et liberavi vos de manu eius
JOSH|24|11|transistisque Iordanem et venistis ad Hiericho pugnaveruntque contra vos viri civitatis eius Amorreus et Ferezeus et Chananeus et Hettheus et Gergeseus et Eveus et Iebuseus et tradidi illos in manus vestras
JOSH|24|12|misique ante vos crabrones et eieci eos de locis suis duos reges Amorreorum non in gladio et arcu tuo
JOSH|24|13|dedique vobis terram in qua non laborastis et urbes quas non aedificastis ut habitaretis in eis vineas et oliveta quae non plantastis
JOSH|24|14|nunc ergo timete Dominum et servite ei perfecto corde atque verissimo et auferte deos quibus servierunt patres vestri in Mesopotamia et in Aegypto ac servite Domino
JOSH|24|15|sin autem malum vobis videtur ut Domino serviatis optio vobis datur eligite hodie quod placet cui potissimum servire debeatis utrum diis quibus servierunt patres vestri in Mesopotamia an diis Amorreorum in quorum terra habitatis ego autem et domus mea serviemus Domino
JOSH|24|16|responditque populus et ait absit a nobis ut relinquamus Dominum et serviamus diis alienis
JOSH|24|17|Dominus Deus noster ipse eduxit nos et patres nostros de terra Aegypti de domo servitutis fecitque videntibus nobis signa ingentia et custodivit nos in omni via per quam ambulavimus et in cunctis populis per quos transivimus
JOSH|24|18|et eiecit universas gentes Amorreum habitatorem terrae quam nos intravimus serviemus igitur Domino quia ipse est Deus noster
JOSH|24|19|dixitque Iosue ad populum non poteritis servire Domino Deus enim sanctus et fortis aemulator est nec ignoscet sceleribus vestris atque peccatis
JOSH|24|20|si dimiseritis Dominum et servieritis diis alienis convertet se et adfliget vos atque subvertet postquam vobis praestiterit bona
JOSH|24|21|dixitque populus ad Iosue nequaquam ita ut loqueris erit sed Domino serviemus
JOSH|24|22|et Iosue ad populum testes inquit vos estis quia ipsi elegeritis vobis Dominum ut serviatis ei responderuntque testes
JOSH|24|23|nunc ergo ait auferte deos alienos de medio vestrum et inclinate corda vestra ad Dominum Deum Israhel
JOSH|24|24|dixitque populus ad Iosue Domino Deo nostro serviemus oboedientes praeceptis eius
JOSH|24|25|percussit igitur Iosue in die illo foedus et proposuit populo praecepta atque iudicia in Sychem
JOSH|24|26|scripsitque omnia verba haec in volumine legis Dei et tulit lapidem pergrandem posuitque eum subter quercum quae erat in sanctuario Domini
JOSH|24|27|et dixit ad omnem populum en lapis iste erit vobis in testimonium quod audierit omnia verba Domini quae locutus est vobis ne forte postea negare velitis et mentiri Domino Deo vestro
JOSH|24|28|dimisitque populum singulos in possessionem suam
JOSH|24|29|et post haec mortuus est Iosue filius Nun servus Domini centum decem annorum
JOSH|24|30|sepelieruntque eum in finibus possessionis suae in Thamnathsare quae sita est in monte Ephraim a septentrionali parte montis Gaas
JOSH|24|31|servivitque Israhel Domino cunctis diebus Iosue et seniorum qui longo vixerunt tempore post Iosue et qui noverant omnia opera Domini quae fecerat in Israhel
JOSH|24|32|ossa quoque Ioseph quae tulerant filii Israhel de Aegypto sepelierunt in Sychem in parte agri quem emerat Iacob a filiis Emmor patris Sychem centum novellis ovibus et fuit in possessione filiorum Ioseph
JOSH|24|33|Eleazar quoque filius Aaron mortuus est et sepelierunt eum in Gaab Finees filii eius quae data est ei in monte Ephraim
JUDG|1|1|post mortem Iosue consuluerunt filii Israhel Dominum dicentes quis ascendet ante nos contra Chananeum et erit dux belli
JUDG|1|2|dixitque Dominus Iudas ascendet ecce tradidi terram in manus eius
JUDG|1|3|et ait Iudas Symeoni fratri suo ascende mecum in sorte mea et pugna contra Chananeum ut et ego pergam tecum in sorte tua et abiit cum eo Symeon
JUDG|1|4|ascenditque Iudas et tradidit Dominus Chananeum ac Ferezeum in manus eorum et percusserunt in Bezec decem milia virorum
JUDG|1|5|inveneruntque Adonibezec in Bezec et pugnaverunt contra eum ac percusserunt Chananeum et Ferezeum
JUDG|1|6|fugit autem Adonibezec quem secuti conprehenderunt caesis summitatibus manuum eius ac pedum
JUDG|1|7|dixitque Adonibezec septuaginta reges amputatis manuum ac pedum summitatibus colligebant sub mensa mea ciborum reliquias sicut feci ita reddidit mihi Deus adduxeruntque eum in Hierusalem et ibi mortuus est
JUDG|1|8|obpugnantes ergo filii Iuda Hierusalem ceperunt eam et percusserunt in ore gladii tradentes cunctam incendio civitatem
JUDG|1|9|et postea descendentes pugnaverunt contra Chananeum qui habitabat in montanis et ad meridiem et in campestribus
JUDG|1|10|pergensque Iudas contra Chananeum qui habitabat in Hebron cui nomen fuit antiquitus Cariatharbe percussit Sisai et Ahiman et Tholmai
JUDG|1|11|atque inde profectus abiit ad habitatores Dabir cuius nomen vetus erat Cariathsepher id est civitas Litterarum
JUDG|1|12|dixitque Chaleb qui percusserit Cariathsepher et vastaverit eam dabo ei Axam filiam meam uxorem
JUDG|1|13|cumque cepisset eam Othonihel filius Cenez frater Chaleb minor dedit ei filiam suam coniugem
JUDG|1|14|quam pergentem in itinere monuit vir suus ut peteret a patre suo agrum quae cum suspirasset sedens asino dixit ei Chaleb quid habes
JUDG|1|15|at illa respondit da mihi benedictionem quia terram arentem dedisti mihi da et inriguam aquis dedit ergo ei Chaleb inriguum superius et inriguum inferius
JUDG|1|16|filii autem Cinei cognati Mosi ascenderunt de civitate Palmarum cum filiis Iuda in desertum sortis eius quod est ad meridiem Arad et habitaverunt cum eo
JUDG|1|17|abiit autem Iudas cum Symeone fratre suo et percusserunt simul Chananeum qui habitabat in Sephath et interfecerunt eum vocatumque est nomen urbis Horma id est anathema
JUDG|1|18|cepitque Iudas Gazam cum finibus suis et Ascalonem atque Accaron cum terminis suis
JUDG|1|19|fuitque Dominus cum Iuda et montana possedit nec potuit delere habitatores vallis quia falcatis curribus abundabant
JUDG|1|20|dederuntque Chaleb Hebron sicut dixerat Moses qui delevit ex ea tres filios Enach
JUDG|1|21|Iebuseum autem habitatorem Hierusalem non deleverunt filii Beniamin habitavitque Iebuseus cum filiis Beniamin in Hierusalem usque in praesentem diem
JUDG|1|22|domus quoque Ioseph ascendit in Bethel fuitque Dominus cum eis
JUDG|1|23|nam cum obsiderent urbem quae prius Luza vocabatur
JUDG|1|24|viderunt hominem egredientem de civitate dixeruntque ad eum ostende nobis introitum civitatis et faciemus tecum misericordiam
JUDG|1|25|qui cum ostendisset eis percusserunt urbem in ore gladii hominem autem illum et omnem cognationem eius dimiserunt
JUDG|1|26|qui dimissus abiit in terram Etthim et aedificavit ibi civitatem vocavitque eam Luzam quae ita appellatur usque in praesentem diem
JUDG|1|27|Manasses quoque non delevit Bethsan et Thanach cum viculis suis et habitatores Dor et Ieblaam et Mageddo cum viculis suis coepitque Chananeus habitare cum eis
JUDG|1|28|postquam autem confortatus est Israhel fecit eos tributarios et delere noluit
JUDG|1|29|Ephraim etiam non interfecit Chananeum qui habitabat in Gazer sed habitavit cum eo
JUDG|1|30|Zabulon non delevit habitatores Cetron et Naalon sed habitavit Chananeus in medio eius factusque est ei tributarius
JUDG|1|31|Aser quoque non delevit habitatores Achcho et Sidonis Alab et Achazib et Alba et Afec et Roob
JUDG|1|32|habitavitque in medio Chananei habitatoris illius terrae nec interfecit eum
JUDG|1|33|Nepthali non delevit habitatores Bethsemes et Bethanath et habitavit inter Chananeum habitatorem terrae fueruntque ei Bethsemitae et Bethanitae tributarii
JUDG|1|34|artavitque Amorreus filios Dan in monte nec dedit eis locum ut ad planiora descenderent
JUDG|1|35|habitavitque in monte Hares quod interpretatur testaceo in Ahilon et Salabim et adgravata est manus domus Ioseph factusque est ei tributarius
JUDG|1|36|fuit autem terminus Amorrei ab ascensu Scorpionis Petra et superiora loca
JUDG|2|1|ascenditque angelus Domini de Galgal ad locum Flentium et ait eduxi vos de Aegypto et introduxi in terram pro qua iuravi patribus vestris et pollicitus sum ut non facerem irritum pactum meum vobiscum in sempiternum
JUDG|2|2|ita dumtaxat ut non feriretis foedus cum habitatoribus terrae huius et aras eorum subverteretis et noluistis audire vocem meam cur hoc fecistis
JUDG|2|3|quam ob rem nolui delere eos a facie vestra ut habeatis hostes et dii eorum sint vobis in ruinam
JUDG|2|4|cumque loqueretur angelus Domini verba haec ad omnes filios Israhel elevaverunt vocem suam et fleverunt
JUDG|2|5|et vocatum est nomen loci illius Flentium sive Lacrimarum immolaveruntque ibi hostias Domino
JUDG|2|6|dimisit ergo Iosue populum et abierunt filii Israhel unusquisque in possessionem suam ut obtinerent eam
JUDG|2|7|servieruntque Domino cunctis diebus eius et seniorum qui longo post eum vixerunt tempore et noverant omnia opera Domini quae fecerat cum Israhel
JUDG|2|8|mortuus est autem Iosue filius Nun famulus Domini centum et decem annorum
JUDG|2|9|et sepelierunt eum in finibus possessionis suae in Thamnathsare in monte Ephraim a septentrionali plaga montis Gaas
JUDG|2|10|omnisque illa generatio congregata est ad patres suos et surrexerunt alii qui non noverant Dominum et opera quae fecerat cum Israhel
JUDG|2|11|feceruntque filii Israhel malum in conspectu Domini et servierunt Baalim
JUDG|2|12|ac dimiserunt Dominum Deum patrum suorum qui eduxerat eos de terra Aegypti et secuti sunt deos alienos deos quoque populorum qui habitabant in circuitu eorum et adoraverunt eos et ad iracundiam concitaverunt Dominum
JUDG|2|13|dimittentes eum et servientes Baal et Astharoth
JUDG|2|14|iratusque Dominus contra Israhel tradidit eos in manibus diripientium qui ceperunt eos et vendiderunt hostibus qui habitabant per gyrum nec potuerunt resistere adversariis suis
JUDG|2|15|sed quocumque pergere voluissent manus Domini erat super eos sicut locutus est et iuravit eis et vehementer adflicti sunt
JUDG|2|16|suscitavitque Dominus iudices qui liberarent eos de vastantium manibus sed nec illos audire voluerunt
JUDG|2|17|fornicantes cum diis alienis et adorantes eos cito deseruerunt viam per quam ingressi fuerant patres eorum et audientes mandata Domini omnia fecere contraria
JUDG|2|18|cumque Dominus iudices suscitaret in diebus eorum flectebatur misericordia et audiebat adflictorum gemitus et liberabat eos de caede vastantium
JUDG|2|19|postquam autem mortuus esset iudex revertebantur et multo maiora faciebant quam fecerant patres sui sequentes deos alienos et servientes eis et adorantes illos non dimiserunt adinventiones suas et viam durissimam per quam ambulare consueverant
JUDG|2|20|iratusque est furor Domini in Israhel et ait quia irritum fecit gens ista pactum meum quod pepigeram cum patribus eorum et vocem meam audire contempsit
JUDG|2|21|et ego non delebo gentes quas dimisit Iosue et mortuus est
JUDG|2|22|ut in ipsis experiar Israhel utrum custodiant viam Domini et ambulent in ea sicut custodierunt patres eorum an non
JUDG|2|23|dimisit ergo Dominus omnes has nationes et cito subvertere noluit nec tradidit in manibus Iosue
JUDG|3|1|hae sunt gentes quas Dominus dereliquit ut erudiret in eis Israhelem et omnes qui non noverant bella Chananeorum
JUDG|3|2|et postea discerent filii eorum certare cum hostibus et habere consuetudinem proeliandi
JUDG|3|3|quinque satrapas Philisthinorum omnemque Chananeum et Sidonium atque Eveum qui habitabat in monte Libano de monte Baalhermon usque ad introitum Emath
JUDG|3|4|dimisitque eos ut in ipsis experiretur Israhelem utrum audiret mandata Domini quae praeceperat patribus eorum per manum Mosi an non
JUDG|3|5|itaque filii Israhel habitaverunt in medio Chananei et Hetthei et Amorrei et Ferezei et Evei et Iebusei
JUDG|3|6|et duxerunt uxores filias eorum ipsique filias suas eorum filiis tradiderunt et servierunt diis eorum
JUDG|3|7|feceruntque malum in conspectu Domini et obliti sunt Dei sui servientes Baalim et Astharoth
JUDG|3|8|iratusque Dominus contra Israhel tradidit eos in manus Chusanrasathaim regis Mesopotamiae servieruntque ei octo annis
JUDG|3|9|et clamaverunt ad Dominum qui suscitavit eis salvatorem et liberavit eos Othonihel videlicet filium Cenez fratrem Chaleb minorem
JUDG|3|10|fuitque in eo spiritus Domini et iudicavit Israhel egressusque est ad pugnam et tradidit Dominus in manu eius Chusanrasathaim regem Syriae et oppressit eum
JUDG|3|11|quievitque terra quadraginta annis et mortuus est Othonihel filius Cenez
JUDG|3|12|addiderunt autem filii Israhel facere malum in conspectu Domini qui confortavit adversum eos Eglon regem Moab quia fecerunt malum in conspectu eius
JUDG|3|13|et copulavit ei filios Ammon et Amalech abiitque et percussit Israhel atque possedit urbem Palmarum
JUDG|3|14|servieruntque filii Israhel Eglon regi Moab decem et octo annis
JUDG|3|15|et postea clamaverunt ad Dominum qui suscitavit eis salvatorem vocabulo Ahoth filium Gera filii Iemini qui utraque manu utebatur pro dextera miseruntque filii Israhel per illum munera Eglon regi Moab
JUDG|3|16|qui fecit sibi gladium ancipitem habentem in medio capulum longitudinis palmae manus et accinctus est eo subter sagum in dextro femore
JUDG|3|17|obtulitque munera Eglon regi Moab erat autem Eglon crassus nimis
JUDG|3|18|cumque obtulisset ei munera prosecutus est socios qui cum eo venerant
JUDG|3|19|et reversus de Galgalis ubi erant idola dixit ad regem verbum secretum habeo ad te o rex et ille imperavit silentium egressisque omnibus qui circa eum erant
JUDG|3|20|ingressus est Ahoth ad eum sedebat autem in aestivo cenaculo solus dixitque verbum Dei habeo ad te qui statim surrexit de throno
JUDG|3|21|extenditque Ahoth manum sinistram et tulit sicam de dextro femore suo infixitque eam in ventre eius
JUDG|3|22|tam valide ut capulus ferrum sequeretur in vulnere ac pinguissimo adipe stringeretur nec eduxit gladium sed ita ut percusserat reliquit in corpore statimque per secreta naturae alvi stercora proruperunt
JUDG|3|23|Ahoth autem clausis diligentissime ostiis cenaculi et obfirmatis sera
JUDG|3|24|per posticam egressus est servique regis ingressi viderunt clausas fores cenaculi atque dixerunt forsitan purgat alvum in aestivo cubiculo
JUDG|3|25|expectantesque diu donec erubescerent et videntes quod nullus aperiret tulerunt clavem et aperientes invenerunt dominum suum iacentem in terra mortuum
JUDG|3|26|Ahoth autem dum illi turbarentur effugit et pertransiit locum Idolorum unde reversus fuerat venitque in Seirath
JUDG|3|27|et statim insonuit bucina in monte Ephraim descenderuntque cum eo filii Israhel ipso in fronte gradiente
JUDG|3|28|qui dixit ad eos sequimini me tradidit enim Dominus inimicos nostros Moabitas in manus nostras descenderuntque post eum et occupaverunt vada Iordanis quae transmittunt in Moab et non dimiserunt transire quemquam
JUDG|3|29|sed percusserunt Moabitas in tempore illo circiter decem milia omnes robustos et fortes viros nullus eorum evadere potuit
JUDG|3|30|humiliatusque est Moab die illo sub manu Israhel et quievit terra octoginta annis
JUDG|3|31|post hunc fuit Samgar filius Anath qui percussit de Philisthim sescentos viros vomere et ipse quoque defendit Israhel
JUDG|4|1|addideruntque filii Israhel facere malum in conspectu Domini post mortem Ahoth
JUDG|4|2|et tradidit illos Dominus in manu Iabin regis Chanaan qui regnavit in Asor habuitque ducem exercitus sui nomine Sisaram ipse autem habitabat in Aroseth gentium
JUDG|4|3|clamaveruntque filii Israhel ad Dominum nongentos enim habebat falcatos currus et per viginti annos vehementer oppresserat eos
JUDG|4|4|erat autem Debbora prophetis uxor Lapidoth quae iudicabat populum in illo tempore
JUDG|4|5|et sedebat sub palma quae nomine illius vocabatur inter Rama et Bethel in monte Ephraim ascendebantque ad eam filii Israhel in omne iudicium
JUDG|4|6|quae misit et vocavit Barac filium Abinoem de Cedes Nepthalim dixitque ad eum praecepit tibi Dominus Deus Israhel vade et duc exercitum in montem Thabor tollesque tecum decem milia pugnatorum de filiis Nepthalim et de filiis Zabulon
JUDG|4|7|ego autem ducam ad te in loco torrentis Cison Sisaram principem exercitus Iabin et currus eius atque omnem multitudinem et tradam eos in manu tua
JUDG|4|8|dixitque ad eam Barac si venis mecum vadam si nolueris venire non pergam
JUDG|4|9|quae dixit ad eum ibo quidem tecum sed in hac vice tibi victoria non reputabitur quia in manu mulieris tradetur Sisara surrexit itaque Debbora et perrexit cum Barac in Cedes
JUDG|4|10|qui accitis Zabulon et Nepthalim ascendit cum decem milibus pugnatorum habens Debboram in comitatu suo
JUDG|4|11|Aber autem Cineus recesserat quondam a ceteris Cineis fratribus suis filiis Obab cognati Mosi et tetenderat tabernacula usque ad vallem quae vocatur Sennim et erat iuxta Cedes
JUDG|4|12|nuntiatumque est Sisarae quod ascendisset Barac filius Abinoem in montem Thabor
JUDG|4|13|et congregavit nongentos falcatos currus omnemque exercitum de Aroseth gentium ad torrentem Cison
JUDG|4|14|dixitque Debbora ad Barac surge haec est enim dies in qua tradidit Dominus Sisaram in manus tuas en ipse ductor est tuus descendit itaque Barac de monte Thabor et decem milia pugnatorum cum eo
JUDG|4|15|perterruitque Dominus Sisaram et omnes currus eius universamque multitudinem in ore gladii ad conspectum Barac in tantum ut Sisara de curru desiliens pedibus fugeret
JUDG|4|16|et Barac persequeretur fugientes currus et exercitum usque ad Aroseth gentium et omnis hostium multitudo usque ad internicionem caderet
JUDG|4|17|Sisara autem fugiens pervenit ad tentorium Iahel uxoris Aber Cinei erat enim pax inter Iabin regem Asor et domum Aber Cinei
JUDG|4|18|egressa igitur Iahel in occursum Sisarae dixit ad eum intra ad me domine mi intra ne timeas qui ingressus tabernaculum eius et opertus ab ea pallio
JUDG|4|19|dixit ad eam da mihi obsecro paululum aquae quia valde sitio quae aperuit utrem lactis et dedit ei bibere et operuit illum
JUDG|4|20|dixitque Sisara ad eam sta ante ostium tabernaculi et cum venerit aliquis interrogans te et dicens numquid hic est aliquis respondebis nullus est
JUDG|4|21|tulit itaque Iahel uxor Aber clavum tabernaculi adsumens pariter malleum et ingressa abscondite et cum silentio posuit supra tempus capitis eius clavum percussumque malleo defixit in cerebrum usque ad terram qui soporem morti socians defecit et mortuus est
JUDG|4|22|et ecce Barac sequens Sisaram veniebat egressaque Iahel in occursum eius dixit ei veni et ostendam tibi virum quem quaeris qui cum intrasset ad eam vidit Sisaram iacentem mortuum et clavum infixum in tempore eius
JUDG|4|23|humiliavit ergo Deus in die illo Iabin regem Chanaan coram filiis Israhel
JUDG|4|24|qui crescebant cotidie et forti manu opprimebant Iabin regem Chanaan donec delerent eum
JUDG|5|1|cecineruntque Debbora et Barac filius Abinoem in die illo dicentes
JUDG|5|2|qui sponte obtulistis de Israhel animas vestras ad periculum benedicite Domino
JUDG|5|3|audite reges percipite auribus principes ego sum ego sum quae Domino canam psallam Domino Deo Israhel
JUDG|5|4|Domine cum exires de Seir et transires per regiones Edom terra mota est caelique ac nubes stillaverunt aquis
JUDG|5|5|montes fluxerunt a facie Domini et Sinai a facie Domini Dei Israhel
JUDG|5|6|in diebus Samgar filii Anath in diebus Iahel quieverunt semitae et qui ingrediebantur per eas ambulaverunt per calles devios
JUDG|5|7|cessaverunt fortes in Israhel et quieverunt donec surgeret Debbora surgeret mater in Israhel
JUDG|5|8|nova bella elegit Dominus et portas hostium ipse subvertit clypeus et hasta si apparuerint in quadraginta milibus Israhel
JUDG|5|9|cor meum diligit principes Israhel qui propria voluntate obtulistis vos discrimini benedicite Domino
JUDG|5|10|qui ascenditis super nitentes asinos et sedetis in iudicio et ambulatis in via loquimini
JUDG|5|11|ubi conlisi sunt currus et hostium est suffocatus exercitus ibi narrentur iustitiae Domini et clementia in fortes Israhel tunc descendit populus Domini ad portas et obtinuit principatum
JUDG|5|12|surge surge Debbora surge surge et loquere canticum surge Barac et adprehende captivos tuos fili Abinoem
JUDG|5|13|salvatae sunt reliquiae populi Dominus in fortibus dimicavit
JUDG|5|14|ex Ephraim delevit eos in Amalech et post eum ex Beniamin in populos tuos o Amalech de Machir principes descenderunt et de Zabulon qui exercitum ducerent ad bellandum
JUDG|5|15|duces Isachar fuere cum Debbora et Barac vestigia sunt secuti qui quasi in praeceps ac baratrum se discrimini dedit diviso contra se Ruben magnanimorum repperta contentio est
JUDG|5|16|quare habitas inter duos terminos ut audias sibilos gregum diviso contra se Ruben magnanimorum repperta contentio est
JUDG|5|17|Galaad trans Iordanem quiescebat et Dan vacabat navibus Aser habitabat in litore maris et in portibus morabatur
JUDG|5|18|Zabulon vero et Nepthalim obtulerunt animas suas morti in regione Merome
JUDG|5|19|venerunt reges et pugnaverunt pugnaverunt reges Chanaan in Thanach iuxta aquas Mageddo et tamen nihil tulere praedantes
JUDG|5|20|de caelo dimicatum est contra eos stellae manentes in ordine et cursu suo adversum Sisaram pugnaverunt
JUDG|5|21|torrens Cison traxit cadavera eorum torrens Cadumim torrens Cison conculca anima mea robustos
JUDG|5|22|ungulae equorum ceciderunt fugientibus impetu et per praeceps ruentibus fortissimis hostium
JUDG|5|23|maledicite terrae Meroz dixit angelus Domini maledicite habitatoribus eius quia non venerunt ad auxilium Domini in adiutorium fortissimorum eius
JUDG|5|24|benedicta inter mulieres Iahel uxor Aber Cinei benedicatur in tabernaculo suo
JUDG|5|25|aquam petenti lac dedit et in fiala principum obtulit butyrum
JUDG|5|26|sinistram manum misit ad clavum et dexteram ad fabrorum malleos percussitque Sisaram quaerens in capite vulneri locum et tempus valide perforans
JUDG|5|27|inter pedes eius ruit defecit et mortuus est ante pedes illius volvebatur et iacebat exanimis et miserabilis
JUDG|5|28|per fenestram prospiciens ululabat mater eius et de cenaculo loquebatur cur moratur regredi currus eius quare tardaverunt pedes quadrigarum illius
JUDG|5|29|una sapientior ceteris uxoribus eius haec socrui verba respondit
JUDG|5|30|forsitan nunc dividit spolia et pulcherrima feminarum eligitur ei vestes diversorum colorum Sisarae traduntur in praedam et supellex varia ad ornanda colla congeritur
JUDG|5|31|sic pereant omnes inimici tui Domine qui autem diligunt te sicut sol in ortu suo splendet ita rutilent
JUDG|5|32|quievitque terra per quadraginta annos
JUDG|6|1|fecerunt autem filii Israhel malum in conspectu Domini qui tradidit eos in manu Madian septem annis
JUDG|6|2|et oppressi sunt valde ab eis feceruntque sibi antra et speluncas in montibus et munitissima ad repugnandum loca
JUDG|6|3|cumque sevisset Israhel ascendebat Madian et Amalech et ceteri orientalium nationum
JUDG|6|4|et apud eos figentes tentoria sicut erant in herbis cuncta vastabant usque ad introitum Gazae nihilque omnino ad vitam pertinens relinquebant in Israhel non oves non boves non asinos
JUDG|6|5|ipsi enim et universi greges eorum veniebant cum tabernaculis et instar lucustarum universa conplebant innumera multitudo hominum et camelorum quicquid tetigerant devastantes
JUDG|6|6|humiliatusque est Israhel valde in conspectu Madian
JUDG|6|7|et clamavit ad Dominum postulans auxilium contra Madianitas
JUDG|6|8|qui misit ad eos virum prophetam et locutus est haec dicit Dominus Deus Israhel ego vos feci conscendere de Aegypto et eduxi de domo servitutis
JUDG|6|9|et liberavi de manu Aegyptiorum et omnium inimicorum qui adfligebant vos eiecique eos ad introitum vestrum et tradidi vobis terram eorum
JUDG|6|10|et dixi ego Dominus Deus vester ne timeatis deos Amorreorum in quorum terra habitatis et noluistis audire vocem meam
JUDG|6|11|venit autem angelus Domini et sedit sub quercu quae erat in Ephra et pertinebat ad Ioas patrem familiae Ezri cumque Gedeon filius eius excuteret atque purgaret frumenta in torculari ut fugeret Madian
JUDG|6|12|apparuit ei et ait Dominus tecum virorum fortissime
JUDG|6|13|dixitque ei Gedeon obsecro Domine si Dominus nobiscum est cur adprehenderunt nos haec omnia ubi sunt mirabilia eius quae narraverunt patres nostri atque dixerunt de Aegypto eduxit nos Dominus nunc autem dereliquit nos et tradidit in manibus Madian
JUDG|6|14|respexitque ad eum Dominus et ait vade in hac fortitudine tua et liberabis Israhel de manu Madian scito quod miserim te
JUDG|6|15|qui respondens ait obsecro Domine mi in quo liberabo Israhel ecce familia mea infima est in Manasse et ego minimus in domo patris mei
JUDG|6|16|dixitque ei Dominus ego ero tecum et percuties Madian quasi unum virum
JUDG|6|17|et ille si inveni inquit gratiam coram te da mihi signum quod tu sis qui loquaris ad me
JUDG|6|18|ne recedas hinc donec revertar ad te portans sacrificium et offerens tibi qui respondit ego praestolabor adventum tuum
JUDG|6|19|ingressus est itaque Gedeon et coxit hedum et de farinae modio azymos panes carnesque ponens in canistro et ius carnium mittens in ollam tulit omnia sub quercum et obtulit ei
JUDG|6|20|cui dixit angelus Domini tolle carnes et panes azymos et pone super petram illam et ius desuper funde cumque fecisset ita
JUDG|6|21|extendit angelus Domini summitatem virgae quam tenebat in manu et tetigit carnes et azymos panes ascenditque ignis de petra et carnes azymosque consumpsit angelus autem Domini evanuit ex oculis eius
JUDG|6|22|vidensque Gedeon quod esset angelus Domini ait heu mihi Domine Deus quia vidi angelum Domini facie ad faciem
JUDG|6|23|dixitque ei Dominus pax tecum ne timeas non morieris
JUDG|6|24|aedificavit ergo ibi Gedeon altare Domino vocavitque illud Domini pax usque in praesentem diem cum adhuc esset in Ephra quae est familiae Ezri
JUDG|6|25|nocte illa dixit Dominus ad eum tolle taurum patris tui et alterum taurum annorum septem destruesque aram Baal quae est patris tui et nemus quod circa aram est succide
JUDG|6|26|et aedificabis altare Domino Deo tuo in summitate petrae huius super quam sacrificium ante posuisti tollesque taurum secundum et offeres holocaustum super lignorum struem quae de nemore succideris
JUDG|6|27|adsumptis igitur Gedeon decem viris de servis suis fecit sicut praeceperat Dominus timens autem domum patris sui et homines illius civitatis per diem facere noluit sed omnia nocte conplevit
JUDG|6|28|cumque surrexissent viri oppidi eius mane viderunt destructam aram Baal lucumque succisum et taurum alterum inpositum super altare quod tunc aedificatum erat
JUDG|6|29|dixeruntque ad invicem quis hoc fecit cumque perquirerent auctorem facti dictum est Gedeon filius Ioas fecit haec omnia
JUDG|6|30|et dixerunt ad Ioas produc filium tuum ut moriatur quia destruxit aram Baal et succidit nemus
JUDG|6|31|quibus ille respondit numquid ultores estis Baal et pugnatis pro eo qui adversarius eius est moriatur antequam lux crastina veniat si deus est vindicet se de eo qui suffodit aram eius
JUDG|6|32|ex illo die vocatus est Gedeon Hierobbaal eo quod dixisset Ioas ulciscatur se de eo Baal qui suffodit altare eius
JUDG|6|33|igitur omnis Madian et Amalech et orientales populi congregati sunt simul et transeuntes Iordanem castrametati sunt in valle Iezrahel
JUDG|6|34|spiritus autem Domini induit Gedeon qui clangens bucina convocavit domum Abiezer ut sequeretur
JUDG|6|35|misitque nuntios in universum Manassen qui et ipse secutus est eum et alios nuntios in Aser et Zabulon et Nepthalim qui occurrerunt ei
JUDG|6|36|dixitque Gedeon ad Dominum si salvum facis per manum meam Israhel sicut locutus es
JUDG|6|37|ponam vellus hoc lanae in area si ros in solo vellere fuerit et in omni terra siccitas sciam quod per manum meam sicut locutus es liberabis Israhel
JUDG|6|38|factumque est ita et de nocte consurgens expresso vellere concam rore conplevit
JUDG|6|39|dixitque rursus ad Dominum ne irascatur furor tuus contra me si adhuc semel temptavero signum quaerens in vellere oro ut solum vellus siccum sit et omnis terra rore madens
JUDG|6|40|fecitque Dominus nocte illa ut postulaverat et fuit siccitas in solo vellere et ros in omni terra
JUDG|7|1|igitur Hierobbaal qui est et Gedeon de nocte consurgens et omnis populus cum eo venit ad fontem qui vocatur Arad erant autem castra Madian in valle ad septentrionalem plagam collis Excelsi
JUDG|7|2|dixitque Dominus ad Gedeon multus tecum est populus nec tradetur Madian in manus eius ne glorietur contra me Israhel et dicat meis viribus liberatus sum
JUDG|7|3|loquere ad populum et cunctis audientibus praedica qui formidolosus et timidus est revertatur recesseruntque de monte Galaad et reversa sunt ex populo viginti duo milia virorum et tantum decem milia remanserunt
JUDG|7|4|dixitque Dominus ad Gedeon adhuc populus multus est duc eos ad aquas et ibi probabo illos et de quo dixero tibi ut tecum vadat ipse pergat quem ire prohibuero revertatur
JUDG|7|5|cumque descendisset populus ad aquas dixit Dominus ad Gedeon qui lingua lambuerint aquas sicut solent canes lambere separabis eos seorsum qui autem curvatis genibus biberint in altera parte erunt
JUDG|7|6|fuit itaque numerus eorum qui manu ad os proiciente aquas lambuerant trecenti viri omnis autem reliqua multitudo flexo poplite biberat
JUDG|7|7|et ait Dominus ad Gedeon in trecentis viris qui lambuerunt aquas liberabo vos et tradam Madian in manu tua omnis autem reliqua multitudo revertatur in locum suum
JUDG|7|8|sumptis itaque pro numero cibariis et tubis omnem reliquam multitudinem abire praecepit ad tabernacula sua et ipse cum trecentis viris se certamini dedit castra autem Madian erant subter in valle
JUDG|7|9|eadem nocte dixit Dominus ad eum surge et descende in castra quia tradidi eos in manu tua
JUDG|7|10|sin autem solus ire formidas descendat tecum Phara puer tuus
JUDG|7|11|et cum audieris quid loquantur tunc confortabuntur manus tuae et securior ad hostium castra descendes descendit ergo ipse et Phara puer eius in partem castrorum ubi erant armatorum vigiliae
JUDG|7|12|Madian autem et Amalech et omnes orientales populi fusi iacebant in valle ut lucustarum multitudo cameli quoque innumerabiles erant sicut harena quae iacet in litoribus maris
JUDG|7|13|cumque venisset Gedeon narrabat aliquis somnium proximo suo et in hunc modum referebat quod viderat vidi somnium et videbatur mihi quasi subcinericius panis ex hordeo volvi et in Madian castra descendere cumque pervenisset ad tabernaculum percussit illud atque subvertit et terrae funditus coaequavit
JUDG|7|14|respondit is cui loquebatur non est hoc aliud nisi gladius Gedeonis filii Ioas viri Israhelitae tradidit Deus in manu eius Madian et omnia castra eius
JUDG|7|15|cumque audisset Gedeon somnium et interpretationem eius adoravit et reversus ad castra Israhel ait surgite tradidit enim Dominus in manus nostras castra Madian
JUDG|7|16|divisitque trecentos viros in tres partes et dedit tubas in manibus eorum lagoenasque vacuas ac lampadas in medio lagoenarum
JUDG|7|17|et dixit ad eos quod me facere videritis hoc facite ingrediar partem castrorum et quod fecero sectamini
JUDG|7|18|quando personaverit tuba in manu mea vos quoque per castrorum circuitum clangite et conclamate Domino et Gedeoni
JUDG|7|19|ingressusque est Gedeon et trecenti viri qui erant cum eo in parte castrorum incipientibus vigiliis noctis mediae et custodibus suscitatis coeperunt bucinis clangere et conplodere inter se lagoenas
JUDG|7|20|cumque per gyrum castrorum in tribus personarent locis et hydrias confregissent tenuerunt sinistris manibus lampadas et dextris sonantes tubas clamaveruntque gladius Domini et Gedeonis
JUDG|7|21|stantes singuli in loco suo per circuitum castrorum hostilium omnia itaque castra turbata sunt et vociferantes ululantesque fugerunt
JUDG|7|22|et nihilominus insistebant trecenti viri bucinis personantes inmisitque Dominus gladium in omnibus castris et mutua se caede truncabant
JUDG|7|23|fugientes usque Bethseta et crepidinem Abelmeula in Tebbath conclamantes autem viri Israhel de Nepthali et Aser et omni Manasse persequebantur Madian
JUDG|7|24|misitque Gedeon nuntios in omnem montem Ephraim dicens descendite in occursum Madian et occupate aquas usque Bethbera atque Iordanem clamavitque omnis Ephraim et praeoccupavit aquas atque Iordanem usque Bethbera
JUDG|7|25|adprehensosque duos viros Madian Oreb et Zeb interfecit Oreb in petra Oreb Zeb vero in torculari Zeb et persecuti sunt Madian capita Oreb et Zeb portantes ad Gedeon trans fluenta Iordanis
JUDG|8|1|dixeruntque ad eum viri Ephraim quid est hoc quod facere voluisti ut non nos vocares cum ad pugnam pergeres contra Madian iurgantes fortiter et prope vim inferentes
JUDG|8|2|quibus ille respondit quid enim tale facere potui quale vos fecistis nonne melior est racemus Ephraim vindemiis Abiezer
JUDG|8|3|in manus vestras tradidit Dominus principes Madian Oreb et Zeb quid tale facere potui quale vos fecistis quod cum locutus esset requievit spiritus eorum quo tumebant contra eum
JUDG|8|4|cumque venisset Gedeon ad Iordanem transivit eum cum trecentis viris qui secum erant et prae lassitudine fugientes persequi non poterant
JUDG|8|5|dixitque ad viros Soccoth date obsecro panes populo qui mecum est quia valde defecerunt ut possimus persequi Zebee et Salmana reges Madian
JUDG|8|6|responderunt principes Soccoth forsitan palmae manuum Zebee et Salmana in manu tua sunt et idcirco postulas ut demus exercitui tuo panes
JUDG|8|7|quibus ille ait cum ergo tradiderit Dominus Zebee et Salmana in manus meas conteram carnes vestras cum spinis tribulisque deserti
JUDG|8|8|et inde conscendens venit in Phanuhel locutusque est ad viros eius loci similia cui et illi responderunt sicut responderant viri Soccoth
JUDG|8|9|dixit itaque et eis cum reversus fuero victor in pace destruam turrem hanc
JUDG|8|10|Zebee autem et Salmana requiescebant cum omni exercitu suo quindecim milia enim viri remanserant ex omnibus turmis orientalium populorum caesis centum viginti milibus bellatorum et educentium gladium
JUDG|8|11|ascendensque Gedeon per viam eorum qui in tabernaculis morabantur ad orientalem partem Nobee et Iecbaa percussit castra hostium qui securi erant et nihil adversi suspicabantur
JUDG|8|12|fugeruntque Zebee et Salmana quos persequens Gedeon conprehendit turbato omni exercitu eorum
JUDG|8|13|revertensque de bello ante solis ortum
JUDG|8|14|adprehendit puerum de viris Soccoth interrogavitque eum nomina principum et seniorum Soccoth et descripsit septuaginta septem viros
JUDG|8|15|venitque ad Soccoth et dixit eis en Zebee et Salmana super quibus exprobrastis mihi dicentes forsitan manus Zebee et Salmana in manibus tuis sunt et idcirco postulas ut demus viris qui lassi sunt et defecerunt panes
JUDG|8|16|tulit ergo seniores civitatis et spinas deserti ac tribulos et contrivit cum eis atque comminuit viros Soccoth
JUDG|8|17|turrem quoque Phanuhel subvertit occisis habitatoribus civitatis
JUDG|8|18|dixitque ad Zebee et Salmana quales fuerunt viri quos occidistis in Thabor qui responderunt similes tui et unus ex eis quasi filius regis
JUDG|8|19|quibus ille ait fratres mei fuerunt filii matris meae vivit Dominus si servassetis eos non vos occiderem
JUDG|8|20|dixitque Ietther primogenito suo surge et interfice eos qui non eduxit gladium timebat enim quia adhuc puer erat
JUDG|8|21|dixeruntque Zebee et Salmana tu surge et inrue in nos quia iuxta aetatem robur est hominis surrexit Gedeon et interfecit Zebee et Salmana et tulit ornamenta ac bullas quibus colla regalium camelorum decorari solent
JUDG|8|22|dixeruntque omnes viri Israhel ad Gedeon dominare nostri tu et filius tuus et filius filii tui quia liberasti nos de manu Madian
JUDG|8|23|quibus ille ait non dominabor vestri nec dominabitur in vos filius meus sed dominabitur Dominus
JUDG|8|24|dixitque ad eos unam petitionem postulo a vobis date mihi inaures ex praeda vestra inaures enim aureas Ismahelitae habere consuerant
JUDG|8|25|qui responderunt libentissime dabimus expandentesque super terram pallium proiecerunt in eo inaures de praeda
JUDG|8|26|et fuit pondus postulatarum inaurium mille septingenti auri sicli absque ornamentis et monilibus et veste purpurea quibus Madian reges uti soliti erant et praeter torques aureos camelorum
JUDG|8|27|fecitque ex eo Gedeon ephod et posuit illud in civitate sua Ephra fornicatusque est omnis Israhel in eo et factum est Gedeoni et omni domui eius in ruinam
JUDG|8|28|humiliatus est autem Madian coram filiis Israhel nec potuerunt ultra elevare cervices sed quievit terra per quadraginta annos quibus praefuit Gedeon
JUDG|8|29|abiit itaque Hierobbaal filius Ioas et habitavit in domo sua
JUDG|8|30|habuitque septuaginta filios qui egressi sunt de femore eius eo quod plures haberet uxores
JUDG|8|31|concubina autem illius quam habebat in Sychem genuit ei filium nomine Abimelech
JUDG|8|32|mortuusque est Gedeon filius Ioas in senectute bona et sepultus in sepulchro Ioas patris sui in Ephra de familia Ezri
JUDG|8|33|postquam autem mortuus est Gedeon aversi sunt filii Israhel et fornicati cum Baalim percusseruntque cum Baal foedus ut esset eis in deum
JUDG|8|34|nec recordati sunt Domini Dei sui qui eruit eos de manu omnium inimicorum suorum per circuitum
JUDG|8|35|nec fecerunt misericordiam cum domo Hierobbaal Gedeon iuxta omnia bona quae fecerat Israheli
JUDG|9|1|abiit autem Abimelech filius Hierobbaal in Sychem ad fratres matris suae et locutus est ad eos et ad omnem cognationem domus patris matris suae dicens
JUDG|9|2|loquimini ad omnes viros Sychem quid vobis est melius ut dominentur vestri septuaginta viri omnes filii Hierobbaal an ut dominetur vobis unus vir simulque considerate quia os vestrum et caro vestra sum
JUDG|9|3|locutique sunt fratres matris eius de eo ad omnes viros Sychem universos sermones istos et inclinaverunt cor eorum post Abimelech dicentes frater noster est
JUDG|9|4|dederuntque illi septuaginta pondo argenti de fano Baalbrith qui conduxit sibi ex eo viros inopes et vagos secutique sunt eum
JUDG|9|5|et venit in domum patris sui Ephra et occidit fratres suos filios Hierobbaal septuaginta viros super lapidem unum remansitque Ioatham filius Hierobbaal minimus et absconditus est
JUDG|9|6|congregati sunt autem omnes viri Sychem et universae familiae urbis Mello abieruntque et constituerunt regem Abimelech iuxta quercum quae stabat in Sychem
JUDG|9|7|quod cum nuntiatum esset Ioatham ivit et stetit in vertice montis Garizim elevataque voce clamavit et dixit audite me viri Sychem ita audiat vos Deus
JUDG|9|8|ierunt ligna ut unguerent super se regem dixeruntque olivae impera nobis
JUDG|9|9|quae respondit numquid possum deserere pinguedinem meam qua et dii utuntur et homines et venire ut inter ligna promovear
JUDG|9|10|dixeruntque ligna ad arborem ficum veni et super nos regnum accipe
JUDG|9|11|quae respondit eis numquid possum deserere dulcedinem meam fructusque suavissimos et ire ut inter cetera ligna commovear
JUDG|9|12|locuta sunt quoque ligna ad vitem veni et impera nobis
JUDG|9|13|quae respondit numquid possum deserere vinum meum quod laetificat Deum et homines et inter ligna cetera commoveri
JUDG|9|14|dixeruntque omnia ligna ad ramnum veni et impera super nos
JUDG|9|15|quae respondit eis si vere me regem vobis constituitis venite et sub mea umbra requiescite sin autem non vultis egrediatur ignis de ramno et devoret cedros Libani
JUDG|9|16|nunc igitur si recte et absque peccato constituistis super vos regem Abimelech et bene egistis cum Hierobbaal et cum domo eius et reddidistis vicem beneficiis eius qui pugnavit pro vobis
JUDG|9|17|et animam suam dedit periculis ut erueret vos de manu Madian
JUDG|9|18|qui nunc surrexistis contra domum patris mei et interfecistis filios eius septuaginta viros super unum lapidem et constituistis regem Abimelech filium ancillae eius super habitatores Sychem eo quod frater vester sit
JUDG|9|19|si ergo recte et absque vitio egistis cum Hierobbaal et domo eius hodie laetamini in Abimelech et ille laetetur in vobis
JUDG|9|20|sin autem perverse egrediatur ignis ex eo et consumat habitatores Sychem et oppidum Mello egrediaturque ignis de viris Sychem et de oppido Mello et devoret Abimelech
JUDG|9|21|quae cum dixisset fugit et abiit in Bera habitavitque ibi metu Abimelech fratris sui
JUDG|9|22|regnavit itaque Abimelech super Israhel tribus annis
JUDG|9|23|misitque Deus spiritum pessimum inter Abimelech et habitatores Sychem qui coeperunt eum detestari
JUDG|9|24|et scelus interfectionis septuaginta filiorum Hierobbaal et effusionem sanguinis eorum conferre in Abimelech fratrem suum et in ceteros Sycimarum principes qui eum adiuverant
JUDG|9|25|posueruntque insidias adversum eum in montium summitate et dum illius praestolantur adventum exercebant latrocinia agentes praedas de praetereuntibus nuntiatumque est Abimelech
JUDG|9|26|venit autem Gaal filius Obed cum fratribus suis et transivit in Sycimam ad cuius adventum erecti habitatores Sychem
JUDG|9|27|egressi sunt in agros vastantes vineas uvasque calcantes et factis cantantium choris ingressi sunt fanum dei sui et inter epulas et pocula maledicebant Abimelech
JUDG|9|28|clamante Gaal filio Obed quis est Abimelech et quae est Sychem ut serviamus ei numquid non est filius Hierobbaal et constituit principem Zebul servum suum super viros Emmor patris Sychem cur igitur servimus ei
JUDG|9|29|utinam daret aliquis populum istum sub manu mea ut auferrem de medio Abimelech dictumque est Abimelech congrega exercitus multitudinem et veni
JUDG|9|30|Zebul enim princeps civitatis auditis sermonibus Gaal filii Obed iratus est valde
JUDG|9|31|et misit clam ad Abimelech nuntios dicens ecce Gaal filius Obed venit in Sycimam cum fratribus suis et obpugnat adversum te civitatem
JUDG|9|32|surge itaque nocte cum populo qui tecum est et latita in agro
JUDG|9|33|et primo mane oriente sole inrue super civitatem illo autem egrediente adversum te cum populo suo fac ei quod potueris
JUDG|9|34|surrexit itaque Abimelech cum omni exercitu suo nocte et tetendit insidias iuxta Sycimam in quattuor locis
JUDG|9|35|egressusque est Gaal filius Obed et stetit in introitu portae civitatis surrexit autem Abimelech et omnis exercitus cum eo de insidiarum loco
JUDG|9|36|cumque vidisset populum Gaal dixit ad Zebul ecce de montibus multitudo descendit cui ille respondit umbras montium vides quasi hominum capita et hoc errore deciperis
JUDG|9|37|rursumque Gaal ait ecce populus de umbilico terrae descendit et unus cuneus venit per viam quae respicit quercum
JUDG|9|38|cui dixit Zebul ubi est nunc os tuum quo loquebaris quis est Abimelech ut serviamus ei nonne iste est populus quem despiciebas egredere et pugna contra eum
JUDG|9|39|abiit ergo Gaal spectante Sycimarum populo et pugnavit contra Abimelech
JUDG|9|40|qui persecutus est eum fugientem et in urbem conpulit cecideruntque ex parte eius plurimi usque ad portam civitatis
JUDG|9|41|et Abimelech sedit in Ruma Zebul autem Gaal et socios eius expulit de urbe nec in ea passus est commorari
JUDG|9|42|sequenti ergo die egressus est populus in campum quod cum nuntiatum esset Abimelech
JUDG|9|43|tulit exercitum suum et divisit in tres turmas tendens insidias in agris vidensque quod egrederetur populus de civitate surrexit et inruit in eos
JUDG|9|44|cum cuneo suo obpugnans et obsidens civitatem duae autem turmae palantes per campum adversarios sequebantur
JUDG|9|45|porro Abimelech omni illo die obpugnabat urbem quam cepit interfectis habitatoribus eius ipsaque destructa ita ut sal in ea dispergeret
JUDG|9|46|quod cum audissent qui habitabant in turre Sycimorum ingressi sunt fanum dei sui Berith ubi foedus cum eo pepigerant et ex eo locus nomen acceperat qui erat valde munitus
JUDG|9|47|Abimelech quoque audiens viros turris Sycimorum pariter conglobatos
JUDG|9|48|ascendit in montem Selmon cum omni populo suo et arrepta securi praecidit arboris ramum inpositumque ferens umero dixit ad socios quod me vidistis facere cito facite
JUDG|9|49|igitur certatim ramos de arboribus praecidentes sequebantur ducem quos circumdantes praesidio succenderunt atque ita factum est ut fumo et igne mille hominum necarentur viri pariter ac mulieres habitatorum turris Sychem
JUDG|9|50|Abimelech autem inde proficiscens venit ad oppidum Thebes quod circumdans obsidebat exercitu
JUDG|9|51|erat autem turris excelsa in media civitate ad quam confugerant viri simul ac mulieres et omnes principes civitatis clausa firmissime ianua et super turris tectum stantes per propugnacula
JUDG|9|52|accedensque Abimelech iuxta turrem pugnabat fortiter et adpropinquans ostio ignem subponere nitebatur
JUDG|9|53|et ecce una mulier fragmen molae desuper iaciens inlisit capiti Abimelech et confregit cerebrum eius
JUDG|9|54|qui vocavit cito armigerum suum et ait ad eum evagina gladium tuum et percute me ne forte dicatur quod a femina interfectus sim qui iussa perficiens interfecit eum
JUDG|9|55|illoque mortuo omnes qui cum eo erant de Israhel reversi sunt in sedes suas
JUDG|9|56|et reddidit Deus malum quod fecerat Abimelech contra patrem suum interfectis septuaginta fratribus suis
JUDG|9|57|Sycimitis quoque quod operati erant retributum est et venit super eos maledictio Ioatham filii Hierobbaal
JUDG|10|1|post Abimelech surrexit dux in Israhel Thola filius Phoa patrui Abimelech vir de Isachar qui habitavit in Sanir montis Ephraim
JUDG|10|2|et iudicavit Israhel viginti et tribus annis mortuusque ac sepultus est in Sanir
JUDG|10|3|huic successit Iair Galaadites qui iudicavit Israhel per viginti et duos annos
JUDG|10|4|habens triginta filios sedentes super triginta pullos asinarum et principes triginta civitatum quae ex nomine eius appellatae sunt Avothiair id est oppida Iair usque in praesentem diem in terra Galaad
JUDG|10|5|mortuusque est Iair ac sepultus in loco cui est vocabulum Camon
JUDG|10|6|filii autem Israhel peccatis veteribus iungentes nova fecerunt malum in conspectu Domini et servierunt idolis Baalim et Astharoth et diis Syriae ac Sidonis et Moab et filiorum Ammon et Philisthim dimiseruntque Dominum et non colebant eum
JUDG|10|7|contra quos iratus tradidit eos in manu Philisthim et filiorum Ammon
JUDG|10|8|adflictique sunt et vehementer oppressi per annos decem et octo omnes qui habitabant trans Iordanem in terra Amorrei quae est in Galaad
JUDG|10|9|in tantum ut filii Ammon Iordane transmisso vastarent Iudam et Beniamin et Ephraim adflictusque est Israhel nimis
JUDG|10|10|et clamantes ad Dominum dixerunt peccavimus tibi quia dereliquimus Deum nostrum et servivimus Baalim
JUDG|10|11|quibus locutus est Dominus numquid non Aegyptii et Amorrei filiique Ammon et Philisthim
JUDG|10|12|Sidonii quoque et Amalech et Chanaan oppresserunt vos et clamastis ad me et erui vos de manu eorum
JUDG|10|13|et tamen reliquistis me et coluistis deos alienos idcirco non addam ut ultra vos liberem
JUDG|10|14|ite et invocate deos quos elegistis ipsi vos liberent in tempore angustiae
JUDG|10|15|dixeruntque filii Israhel ad Dominum peccavimus redde tu nobis quicquid tibi placet tantum nunc libera nos
JUDG|10|16|quae dicentes omnia de finibus suis alienorum deorum idola proiecerunt et servierunt Deo qui doluit super miseriis eorum
JUDG|10|17|itaque filii Ammon conclamantes in Galaad fixere tentoria contra quos congregati filii Israhel in Maspha castrametati sunt
JUDG|10|18|dixeruntque principes Galaad singuli ad proximos suos qui primus e nobis contra filios Ammon coeperit dimicare erit dux populi Galaad
JUDG|11|1|fuit illo tempore Iepthae Galaadites vir fortissimus atque pugnator filius meretricis mulieris qui natus est de Galaad
JUDG|11|2|habuit autem Galaad uxorem de qua suscepit filios qui postquam creverant eiecerunt Iepthae dicentes heres in domo patris nostri esse non poteris quia de altera matre generatus es
JUDG|11|3|quos ille fugiens atque devitans habitavit in terra Tob congregatique sunt ad eum viri inopes et latrocinantes et quasi principem sequebantur
JUDG|11|4|in illis diebus pugnabant filii Ammon contra Israhel
JUDG|11|5|quibus acriter instantibus perrexerunt maiores natu de Galaad ut tollerent in auxilium sui Iepthae de terra Tob
JUDG|11|6|dixeruntque ad eum veni et esto princeps noster et pugna contra filios Ammon
JUDG|11|7|quibus ille respondit nonne vos estis qui odistis me et eiecistis de domo patris mei et nunc venistis ad me necessitate conpulsi
JUDG|11|8|dixeruntque principes Galaad ad Iepthae ob hanc igitur causam nunc ad te venimus ut proficiscaris nobiscum et pugnes contra filios Ammon sisque dux omnium qui habitant in Galaad
JUDG|11|9|Iepthae quoque dixit eis si vere venistis ad me ut pugnem pro vobis contra filios Ammon tradideritque eos Dominus in manus meas ego ero princeps vester
JUDG|11|10|qui responderunt ei Dominus qui haec audit ipse mediator ac testis est quod nostra promissa faciamus
JUDG|11|11|abiit itaque Iepthae cum principibus Galaad fecitque eum omnis populus principem sui locutusque est Iepthae omnes sermones suos coram Domino in Maspha
JUDG|11|12|et misit nuntios ad regem filiorum Ammon qui ex persona sua dicerent quid mihi et tibi est quia venisti contra me ut vastares terram meam
JUDG|11|13|quibus ille respondit quia tulit Israhel terram meam quando ascendit de Aegypto a finibus Arnon usque Iaboc atque Iordanem nunc igitur cum pace redde mihi eam
JUDG|11|14|per quos rursum mandavit Iepthae et imperavit eis ut dicerent regi Ammon
JUDG|11|15|haec dicit Iepthae non tulit Israhel terram Moab nec terram filiorum Ammon
JUDG|11|16|sed quando de Aegypto conscenderunt ambulavit per solitudinem usque ad mare Rubrum et venit in Cades
JUDG|11|17|misitque nuntios ad regem Edom dicens dimitte ut transeam per terram tuam qui noluit adquiescere precibus eius misit quoque et ad regem Moab qui et ipse transitum praebere contempsit mansit itaque in Cades
JUDG|11|18|et circuivit ex latere terram Edom et terram Moab venitque contra orientalem plagam terrae Moab et castrametatus est trans Arnon nec voluit intrare terminos Moab Arnon quippe confinium est terrae Moab
JUDG|11|19|misit itaque Israhel nuntios ad Seon regem Amorreorum qui habitabat in Esebon et dixerunt ei dimitte ut transeam per terram tuam usque ad fluvium
JUDG|11|20|qui et ipse Israhel verba despiciens non dimisit eum transire per terminos suos sed infinita multitudine congregata egressus est contra eum in Iassa et fortiter resistebat
JUDG|11|21|tradiditque eum Dominus in manu Israhel cum omni exercitu suo qui percussit eum et possedit omnem terram Amorrei habitatoris regionis illius
JUDG|11|22|et universos fines eius de Arnon usque Iaboc et de solitudine usque ad Iordanem
JUDG|11|23|Dominus ergo Deus Israhel subvertit Amorreum pugnante contra illum populo suo Israhel et tu nunc vis possidere terram eius
JUDG|11|24|nonne ea quae possedit Chamos deus tuus tibi iure debentur quae autem Dominus Deus noster victor obtinuit in nostram cedent possessionem
JUDG|11|25|nisi forte melior es Balac filio Sepphor rege Moab aut docere potes quod iurgatus sit contra Israhel et pugnaverit contra eum
JUDG|11|26|quando habitavit in Esebon et viculis eius et in Aroer et villis illius vel in cunctis civitatibus iuxta Iordanem per trecentos annos quare tanto tempore nihil super hac repetitione temptastis
JUDG|11|27|igitur non ego pecco in te sed tu contra me male agis indicens mihi bella non iusta iudicet Dominus arbiter huius diei inter Israhel et inter filios Ammon
JUDG|11|28|noluitque adquiescere rex filiorum Ammon verbis Iepthae quae per nuntios mandaverat
JUDG|11|29|factus est ergo super Iepthae spiritus Domini et circumiens Galaad et Manasse Maspha quoque Galaad et inde transiens ad filios Ammon
JUDG|11|30|votum vovit Domino dicens si tradideris filios Ammon in manus meas
JUDG|11|31|quicumque primus fuerit egressus de foribus domus meae mihique occurrerit revertenti cum pace a filiis Ammon eum holocaustum offeram Domino
JUDG|11|32|transivitque Iepthae ad filios Ammon ut pugnaret contra eos quos tradidit Dominus in manus eius
JUDG|11|33|percussitque ab Aroer usque dum venias in Mennith viginti civitates et usque ad Abel quae est vineis consita plaga magna nimis humiliatique sunt filii Ammon a filiis Israhel
JUDG|11|34|revertenti autem Iepthae in Maspha domum suam occurrit unigenita filia cum tympanis et choris non enim habebat alios liberos
JUDG|11|35|qua visa scidit vestimenta sua et ait heu filia mi decepisti me et ipsa decepta es aperui enim os meum ad Dominum et aliud facere non potero
JUDG|11|36|cui illa respondit pater mi si aperuisti os tuum ad Dominum fac mihi quodcumque pollicitus es concessa tibi ultione atque victoria de hostibus tuis
JUDG|11|37|dixitque ad patrem hoc solum mihi praesta quod deprecor dimitte me ut duobus mensibus circumeam montes et plangam virginitatem meam cum sodalibus meis
JUDG|11|38|cui ille respondit vade et dimisit eam duobus mensibus cumque abisset cum sociis ac sodalibus suis flebat virginitatem suam in montibus
JUDG|11|39|expletisque duobus mensibus reversa est ad patrem suum et fecit ei sicut voverat quae ignorabat virum exinde mos increbuit in Israhel et consuetudo servata est
JUDG|11|40|ut post anni circulum conveniant in unum filiae Israhel et plangant filiam Iepthae Galaaditae diebus quattuor
JUDG|12|1|ecce autem in Ephraim orta seditio est nam transeuntes contra aquilonem dixerunt ad Iepthae quare vadens ad pugnam contra filios Ammon vocare nos noluisti ut pergeremus tecum igitur incendimus domum tuam
JUDG|12|2|quibus ille respondit disceptatio erat mihi et populo meo contra filios Ammon vehemens vocavique vos ut mihi praeberetis auxilium et facere noluistis
JUDG|12|3|quod cernens posui in manibus meis animam meam transivique ad filios Ammon et tradidit eos Dominus in manus meas quid commerui ut adversum me consurgatis in proelium
JUDG|12|4|vocatis itaque ad se cunctis viris Galaad pugnabat contra Ephraim percusseruntque viri Galaad Ephraim quia dixerat fugitivus est Galaad de Ephraim et habitat in medio Ephraim et Manasse
JUDG|12|5|occupaveruntque Galaaditae vada Iordanis per quae Ephraim reversurus erat cumque venisset ad ea de Ephraim numero fugiens atque dixisset obsecro ut me transire permittas dicebant ei Galaaditae numquid Ephrateus es quo dicente non sum
JUDG|12|6|interrogabant eum dic ergo sebboleth quod interpretatur spica qui respondebat tebboleth eadem littera spicam exprimere non valens statimque adprehensum iugulabant in ipso Iordanis transitu et ceciderunt in illo tempore de Ephraim quadraginta duo milia
JUDG|12|7|iudicavitque Iepthae Galaadites Israhel sex annis et mortuus est ac sepultus in civitate sua Galaad
JUDG|12|8|post hunc iudicavit Israhel Abessan de Bethleem
JUDG|12|9|qui habuit triginta filios et totidem filias quas emittens foras maritis dedit et eiusdem numeri filiis suis accepit uxores introducens in domum suam qui septem annis iudicavit Israhel
JUDG|12|10|mortuusque est ac sepultus in Bethleem
JUDG|12|11|cui successit Ahialon Zabulonites et iudicavit Israhelem decem annis
JUDG|12|12|mortuusque est ac sepultus in Zabulon
JUDG|12|13|post hunc iudicavit in Israhel Abdon filius Hellel Farathonites
JUDG|12|14|qui habuit quadraginta filios et triginta ex eis nepotes ascendentes super septuaginta pullos asinarum et iudicavit in Israhel octo annis
JUDG|12|15|mortuusque est ac sepultus in Farathon terrae Ephraim in monte Amalech
JUDG|13|1|rursumque filii Israhel fecerunt malum in conspectu Domini qui tradidit eos in manus Philisthinorum quadraginta annis
JUDG|13|2|erat autem vir quidam de Saraa et de stirpe Dan nomine Manue habens uxorem sterilem
JUDG|13|3|cui apparuit angelus Domini et dixit ad eam sterilis es et absque liberis sed concipies et paries filium
JUDG|13|4|cave ergo ne vinum bibas ac siceram ne inmundum quicquam comedas
JUDG|13|5|quia concipies et paries filium cuius non tanget caput novacula erit enim nazareus Dei ab infantia sua et ex matris utero et ipse incipiet liberare Israhel de manu Philisthinorum
JUDG|13|6|quae cum venisset ad maritum dixit ei vir Dei venit ad me habens vultum angelicum terribilis nimis quem cum interrogassem quis esset et unde venisset et quo nomine vocaretur noluit mihi dicere
JUDG|13|7|sed hoc respondit ecce concipies et paries filium cave ne vinum bibas et siceram et ne aliquo vescaris inmundo erit enim puer nazareus Dei ab infantia sua et ex utero matris usque ad diem mortis suae
JUDG|13|8|oravit itaque Manue Deum et ait obsecro Domine ut vir Dei quem misisti veniat iterum et doceat nos quid debeamus facere de puero qui nasciturus est
JUDG|13|9|exaudivitque Dominus precantem Manue et apparuit rursum angelus Domini uxori eius sedenti in agro Manue autem maritus eius non erat cum ea quae cum vidisset angelum
JUDG|13|10|festinavit et cucurrit ad virum suum nuntiavitque ei dicens ecce apparuit mihi vir quem ante videram
JUDG|13|11|qui surrexit et secutus est uxorem suam veniensque ad virum dixit ei tu es qui locutus es mulieri et ille respondit ego sum
JUDG|13|12|cui Manue quando inquit sermo tuus fuerit expletus quid vis ut faciat puer aut a quo se observare debebit
JUDG|13|13|dixitque angelus Domini ad Manue ab omnibus quae locutus sum uxori tuae abstineat se
JUDG|13|14|et quicquid ex vinea nascitur non comedat vinum et siceram non bibat nullo vescatur inmundo et quod ei praecepi impleat atque custodiat
JUDG|13|15|dixitque Manue ad angelum Domini obsecro te ut adquiescas precibus meis et faciamus tibi hedum de capris
JUDG|13|16|cui respondit angelus si me cogis non comedam panes tuos sin autem vis holocaustum facere offer illud Domino et nesciebat Manue quod angelus Dei esset
JUDG|13|17|dixitque ad eum quod est tibi nomen ut si sermo tuus fuerit expletus honoremus te
JUDG|13|18|cui ille respondit cur quaeris nomen meum quod est mirabile
JUDG|13|19|tulit itaque Manue hedum de capris et libamenta et posuit super petram offerens Domino qui facit mirabilia ipse autem et uxor eius intuebantur
JUDG|13|20|cumque ascenderet flamma altaris in caelum angelus Domini in flamma pariter ascendit quod cum vidisset Manue et uxor eius proni ceciderunt in terram
JUDG|13|21|et ultra non eis apparuit angelus Domini statimque intellexit Manue angelum esse Domini
JUDG|13|22|et dixit ad uxorem suam morte moriemur quia vidimus Deum
JUDG|13|23|cui respondit mulier si Dominus nos vellet occidere de manibus nostris holocaustum et libamenta non suscepisset nec ostendisset nobis haec omnia neque ea quae sunt ventura dixisset
JUDG|13|24|peperit itaque filium et vocavit nomen eius Samson crevitque puer et benedixit ei Dominus
JUDG|13|25|coepitque spiritus Domini esse cum eo in castris Dan inter Saraa et Esthaol
JUDG|14|1|descendit igitur Samson in Thamnatha vidensque ibi mulierem de filiabus Philisthim
JUDG|14|2|ascendit et nuntiavit patri suo et matri dicens vidi mulierem in Thamnatha de filiabus Philisthinorum quam quaeso ut mihi accipiatis uxorem
JUDG|14|3|cui dixerunt pater et mater sua numquid non est mulier in filiabus fratrum tuorum et in omni populo meo quia vis accipere uxorem de Philisthim qui incircumcisi sunt dixitque Samson ad patrem suum hanc mihi accipe quia placuit oculis meis
JUDG|14|4|parentes autem eius nesciebant quod res a Domino fieret et quaereret occasionem contra Philisthim eo enim tempore Philisthim dominabantur Israheli
JUDG|14|5|descendit itaque Samson cum patre suo et matre in Thamnatha cumque venissent ad vineas oppidi apparuit catulus leonis saevus rugiens et occurrit ei
JUDG|14|6|inruit autem spiritus Domini in Samson et dilaceravit leonem quasi hedum in frusta concerperet nihil omnino habens in manu et hoc patri et matri noluit indicare
JUDG|14|7|descenditque et locutus est mulieri quae placuerat oculis eius
JUDG|14|8|et post aliquot dies revertens ut acciperet eam declinavit ut videret cadaver leonis et ecce examen apium in ore leonis erat ac favus mellis
JUDG|14|9|quem cum sumpsisset in manibus comedebat in via veniensque ad patrem suum et matrem dedit eis partem qui et ipsi comederunt nec tamen eis voluit indicare quod mel de corpore leonis adsumpserat
JUDG|14|10|descendit itaque pater eius ad mulierem et fecit filio suo Samson convivium sic enim iuvenes facere consuerant
JUDG|14|11|cum igitur cives loci vidissent eum dederunt ei sodales triginta qui essent cum eo
JUDG|14|12|quibus locutus est Samson proponam vobis problema quod si solveritis mihi intra septem dies convivii dabo vobis triginta sindones et totidem tunicas
JUDG|14|13|sin autem non potueritis solvere vos dabitis mihi triginta sindones et eiusdem numeri tunicas qui responderunt ei propone problema ut audiamus
JUDG|14|14|dixitque eis de comedente exivit cibus et de forte est egressa dulcedo nec potuerunt per tres dies propositionem solvere
JUDG|14|15|cumque adesset dies septimus dixerunt ad uxorem Samson blandire viro tuo et suade ei ut indicet tibi quid significet problema quod si facere nolueris incendimus et te et domum patris tui an idcirco nos vocastis ad nuptias ut spoliaretis
JUDG|14|16|quae fundebat apud Samson lacrimas et querebatur dicens odisti me et non diligis idcirco problema quod proposuisti filiis populi mei non vis mihi exponere at ille respondit patri meo et matri nolui dicere et tibi indicare potero
JUDG|14|17|septem igitur diebus convivii flebat apud eum tandemque die septimo cum ei molesta esset exposuit quae statim indicavit civibus suis
JUDG|14|18|et illi dixerunt ei die septimo ante solis occubitum quid dulcius melle et quid leone fortius qui ait ad eos si non arassetis in vitula mea non invenissetis propositionem meam
JUDG|14|19|inruit itaque in eo spiritus Domini descenditque Ascalonem et percussit ibi triginta viros quorum ablatas vestes dedit his qui problema solverant iratusque nimis ascendit in domum patris sui
JUDG|14|20|uxor autem eius accepit maritum unum de amicis eius et pronubis
JUDG|15|1|post aliquantum autem temporis cum dies triticeae messis instarent venit Samson invisere volens uxorem suam et adtulit ei hedum de capris cumque cubiculum eius solito vellet intrare prohibuit eum pater illius dicens
JUDG|15|2|putavi quod odisses eam et ideo tradidi illam amico tuo sed habet sororem quae iunior et pulchrior illa est sit tibi pro ea uxor
JUDG|15|3|cui respondit Samson ab hac die non erit culpa in me contra Philistheos faciam enim vobis mala
JUDG|15|4|perrexitque et cepit trecentas vulpes caudasque earum iunxit ad caudas et faces ligavit in medio
JUDG|15|5|quas igne succendens dimisit ut huc illucque discurrerent quae statim perrexerunt in segetes Philisthinorum quibus succensis et conportatae iam fruges et adhuc stantes in stipula concrematae sunt in tantum ut vineas quoque et oliveta flamma consumeret
JUDG|15|6|dixeruntque Philisthim quis fecit hanc rem quibus dictum est Samson gener Thamnathei quia tulit uxorem eius et alteri tradidit haec operatus est ascenderuntque Philisthim et conbuserunt tam mulierem quam patrem eius
JUDG|15|7|quibus ait Samson licet haec feceritis tamen adhuc ex vobis expetam ultionem et tunc quiescam
JUDG|15|8|percussitque eos ingenti plaga ita ut stupentes suram femori inponerent et descendens habitavit in spelunca petrae Aetham
JUDG|15|9|igitur ascendentes Philisthim in terra Iuda castrametati sunt et in loco qui postea vocatus est Lehi id est Maxilla eorum est fusus exercitus
JUDG|15|10|dixeruntque ad eos de tribu Iuda cur ascendistis adversum nos qui responderunt ut ligemus Samson venimus et reddamus ei quae in nos operatus est
JUDG|15|11|descenderunt ergo tria milia virorum de Iuda ad specum silicis Aetham dixeruntque ad Samson nescis quod Philisthim imperent nobis quare hoc facere voluisti quibus ille ait sicut fecerunt mihi feci eis
JUDG|15|12|ligare inquiunt te venimus et tradere in manus Philisthinorum iurate respondit mihi quod non me occidatis
JUDG|15|13|dixerunt non te occidimus sed vinctum tradimus ligaveruntque eum duobus novis funibus et tulerunt de petra Aetham
JUDG|15|14|qui cum venisset ad locum Maxillae et Philisthim vociferantes occurrissent ei inruit spiritus Domini in eum et sicut solent ad odorem ignis lina consumi ita vincula quibus ligatus erat dissipata sunt et soluta
JUDG|15|15|inventamque maxillam id est mandibulam asini quae iacebat arripiens interfecit in ea mille viros
JUDG|15|16|et ait in maxilla asini in mandibula pulli asinarum delevi eos et percussi mille viros
JUDG|15|17|cumque haec canens verba conplesset proiecit mandibulam de manu et vocavit nomen loci illius Ramathlehi quod interpretatur elevatio Maxillae
JUDG|15|18|sitiensque valde clamavit ad Dominum et ait tu dedisti in manu servi tui salutem hanc maximam atque victoriam et en siti morior incidamque in manus incircumcisorum
JUDG|15|19|aperuit itaque Dominus molarem dentem in maxilla asini et egressae sunt ex eo aquae quibus haustis refocilavit spiritum et vires recepit idcirco appellatum est nomen loci illius Fons invocantis de maxilla usque in praesentem diem
JUDG|15|20|iudicavitque Israhel in diebus Philisthim viginti annis
JUDG|16|1|abiit quoque in Gazam et vidit ibi meretricem mulierem ingressusque est ad eam
JUDG|16|2|quod cum audissent Philisthim et percrebruisset apud eos intrasse urbem Samson circumdederunt eum positis in porta civitatis custodibus et ibi tota nocte cum silentio praestolantes ut facto mane exeuntem occiderent
JUDG|16|3|dormivit autem Samson usque ad noctis medium et inde consurgens adprehendit ambas portae fores cum postibus suis et sera inpositasque umeris portavit ad verticem montis qui respicit Hebron
JUDG|16|4|post haec amavit mulierem quae habitabat in valle Sorech et vocabatur Dalila
JUDG|16|5|veneruntque ad eam principes Philisthinorum atque dixerunt decipe eum et disce ab illo in quo tantam habeat fortitudinem et quomodo eum superare valeamus et vinctum adfligere quod si feceris dabimus tibi singuli mille centum argenteos
JUDG|16|6|locuta est ergo Dalila ad Samson dic mihi obsecro in quo sit tua maxima fortitudo et quid sit quo ligatus erumpere nequeas
JUDG|16|7|cui respondit Samson si septem nervicis funibus necdum siccis et adhuc humentibus ligatus fuero infirmus ero ut ceteri homines
JUDG|16|8|adtuleruntque ad eam satrapae Philisthinorum septem funes ut dixerat quibus vinxit eum
JUDG|16|9|latentibus apud se insidiis et in cubiculo finem rei expectantibus clamavitque ad eum Philisthim super te Samson qui rupit vincula quomodo si rumpat quis filum de stuppae tortum putamine cum odorem ignis acceperit et non est cognitum in quo esset fortitudo eius
JUDG|16|10|dixitque ad eum Dalila ecce inlusisti mihi et falsum locutus es saltim nunc indica quo ligari debeas
JUDG|16|11|cui ille respondit si ligatus fuero novis funibus qui numquam fuerunt in opere infirmus ero et aliorum hominum similis
JUDG|16|12|quibus rursum Dalila vinxit eum et clamavit Philisthim super te Samson in cubiculo insidiis praeparatis qui ita rupit vincula quasi fila telarum
JUDG|16|13|dixitque Dalila rursum ad eum usquequo decipis me et falsum loqueris ostende quo vinciri debeas si inquit septem crines capitis mei cum licio plexueris et clavum his circumligatum terrae fixeris infirmus ero
JUDG|16|14|quod cum fecisset Dalila dixit ad eum Philisthim super te Samson qui consurgens de somno extraxit clavum cum crinibus et licio
JUDG|16|15|dixitque ad eum Dalila quomodo dicis quod ames me cum animus tuus non sit mecum per tres vices mentitus es mihi et noluisti dicere in quo sit tua maxima fortitudo
JUDG|16|16|cumque molesta ei esset et per multos dies iugiter adhereret spatium ad quietem non tribuens defecit anima eius et ad mortem usque lassata est
JUDG|16|17|tunc aperiens veritatem rei dixit ad eam ferrum numquam ascendit super caput meum quia nazareus id est consecratus Deo sum de utero matris meae si rasum fuerit caput meum recedet a me fortitudo mea et deficiam eroque ut ceteri homines
JUDG|16|18|videns illa quod confessus ei esset omnem animum suum misit ad principes Philisthinorum atque mandavit ascendite adhuc semel quia nunc mihi aperuit cor suum qui ascenderunt adsumpta pecunia quam promiserant
JUDG|16|19|at illa dormire eum fecit super genua sua et in sinu suo reclinare caput vocavitque tonsorem et rasit septem crines eius et coepit abicere eum et a se repellere statim enim ab eo fortitudo discessit
JUDG|16|20|dixitque Philisthim super te Samson qui de somno consurgens dixit in animo suo egrediar sicut ante feci et me excutiam nesciens quod Dominus recessisset ab eo
JUDG|16|21|quem cum adprehendissent Philisthim statim eruerunt oculos eius et duxerunt Gazam vinctum catenis et clausum in carcere molere fecerunt
JUDG|16|22|iamque capilli eius renasci coeperant
JUDG|16|23|et principes Philisthinorum convenerunt in unum ut immolarent hostias magnificas Dagon deo suo et epularentur dicentes tradidit deus noster inimicum nostrum Samson in manus nostras
JUDG|16|24|quod etiam populus videns laudabat deum suum eademque dicebat tradidit deus noster in manus nostras adversarium qui delevit terram nostram et occidit plurimos
JUDG|16|25|laetantesque per convivia sumptis iam epulis praeceperunt ut vocaretur Samson et ante eos luderet qui adductus de carcere ludebat ante eos feceruntque eum stare inter duas columnas
JUDG|16|26|qui dixit puero regenti gressus suos dimitte me ut tangam columnas quibus omnis inminet domus ut recliner super eas et paululum requiescam
JUDG|16|27|domus autem plena erat virorum ac mulierum et erant ibi omnes principes Philisthinorum ac de tecto et solario circiter tria milia utriusque sexus spectabant ludentem Samson
JUDG|16|28|at ille invocato Domino ait Domine Deus memento mei et redde nunc mihi pristinam fortitudinem Deus meus ut ulciscar me de hostibus meis et pro amissione duorum luminum unam ultionem recipiam
JUDG|16|29|et adprehendens ambas columnas quibus innitebatur domus alteramque earum dextera et alteram leva tenens
JUDG|16|30|ait moriatur anima mea cum Philisthim concussisque fortiter columnis cecidit domus super omnes principes et ceteram multitudinem quae ibi erat multoque plures interfecit moriens quam ante vivus occiderat
JUDG|16|31|descendentes autem fratres eius et universa cognatio tulerunt corpus eius et sepelierunt inter Saraa et Esthaol in sepulchro patris Manue iudicavitque Israhel viginti annis
JUDG|17|1|fuit eo tempore vir quidam de monte Ephraim nomine Michas
JUDG|17|2|qui dixit matri suae mille centum argenteos quos separaveras tibi et super quibus me audiente iuraveras ecce ego habeo et apud me sunt cui illa respondit benedictus filius meus Domino
JUDG|17|3|reddidit ergo eos matri suae quae dixerat ei consecravi et vovi argentum hoc Domino ut de manu mea suscipiat filius meus et faciat sculptile atque conflatile et nunc trado illud tibi
JUDG|17|4|reddidit igitur matri suae quae tulit ducentos argenteos et dedit eos argentario ut faceret ex eis sculptile atque conflatile quod fuit in domo Micha
JUDG|17|5|qui aediculam quoque in ea Deo separavit et fecit ephod ac therafin id est vestem sacerdotalem et idola implevitque unius filiorum suorum manum et factus est ei sacerdos
JUDG|17|6|in diebus illis non erat rex in Israhel sed unusquisque quod sibi rectum videbatur hoc faciebat
JUDG|17|7|fuit quoque alter adulescens de Bethleem Iuda et cognatione eius eratque ipse Levites et habitabat ibi
JUDG|17|8|egressusque de civitate Bethleem peregrinari voluit ubicumque sibi commodum repperisset cumque venisset in monte Ephraim iter faciens et declinasset parumper in domum Micha
JUDG|17|9|interrogatus est ab eo unde venis qui respondit Levita sum de Bethleem Iuda et vado ut habitem ubi potuero et utile mihi esse perspexero
JUDG|17|10|mane inquit apud me et esto mihi parens ac sacerdos daboque tibi per annos singulos decem argenteos ac vestem duplicem et quae ad victum necessaria sunt
JUDG|17|11|adquievit et mansit apud hominem fuitque illi quasi unus de filiis
JUDG|17|12|implevitque Micha manum eius et habuit apud se puerum sacerdotem
JUDG|17|13|nunc scio dicens quod bene mihi faciat Deus habenti levitici generis sacerdotem
JUDG|18|1|in diebus illis non erat rex in Israhel et tribus Dan quaerebat possessionem sibi ut habitaret in ea usque ad illum enim diem inter ceteras tribus sortem non acceperat
JUDG|18|2|miserunt igitur filii Dan stirpis et familiae suae quinque viros fortissimos de Saraa et Esthaol ut explorarent terram et diligenter inspicerent dixeruntque eis ite et considerate terram qui cum pergentes venissent in montem Ephraim et intrassent domum Micha requieverunt ibi
JUDG|18|3|et agnoscentes vocem adulescentis Levitae utentesque illius diversorio dixerunt ad eum quis te huc adduxit quid hic agis quam ob causam huc venire voluisti
JUDG|18|4|qui respondit eis haec et haec praestitit mihi Michas et me mercede conduxit ut sim ei sacerdos
JUDG|18|5|rogaveruntque eum ut consuleret Dominum et scire possent an prospero itinere pergerent et res haberet effectum
JUDG|18|6|qui respondit eis ite cum pace Dominus respicit viam vestram et iter quo pergitis
JUDG|18|7|euntes itaque quinque viri venerunt Lais videruntque populum habitantem in ea absque ullo timore iuxta Sidoniorum consuetudinem securum et quietum nullo eis penitus resistente magnarumque opum et procul a Sidone atque a cunctis hominibus separatum
JUDG|18|8|reversique ad fratres suos in Saraa et Esthaol et quid egissent sciscitantibus responderunt
JUDG|18|9|surgite et ascendamus ad eos vidimus enim terram valde opulentam et uberem nolite neglegere nolite cessare eamus et possideamus eam nullus erit labor
JUDG|18|10|intrabimus ad securos in regionem latissimam tradetque nobis Dominus locum in quo nullius rei est penuria eorum quae gignuntur in terra
JUDG|18|11|profecti igitur sunt de cognatione Dan id est de Saraa et Esthaol sescenti viri accincti armis bellicis
JUDG|18|12|ascendentesque manserunt in Cariathiarim Iudae qui locus ex eo tempore castrorum Dan nomen accepit et est post tergum Cariathiarim
JUDG|18|13|inde transierunt in montem Ephraim cumque venissent ad domum Micha
JUDG|18|14|dixerunt quinque viri qui prius missi fuerant ad considerandam terram Lais ceteris fratribus suis nostis quod in domibus istis sit ephod et therafin et sculptile atque conflatile videte quid vobis placeat
JUDG|18|15|et cum paululum declinassent ingressi sunt domum adulescentis Levitae qui erat in domo Micha salutaveruntque eum verbis pacificis
JUDG|18|16|sescenti autem viri ita ut erant armati stabant ante ostium
JUDG|18|17|at illi qui ingressi fuerant domum iuvenis sculptile et ephod et therafin atque conflatile tollere nitebantur et sacerdos stabat ante ostium sescentis viris fortissimis haut procul expectantibus
JUDG|18|18|tulerunt igitur qui intraverant sculptile ephod et idola atque conflatile quibus dixit sacerdos quid facitis
JUDG|18|19|cui responderunt tace et pone digitum super os tuum venique nobiscum ut habeamus te patrem et sacerdotem quid tibi melius est ut sis sacerdos in domo unius viri an in una tribu et familia in Israhel
JUDG|18|20|quod cum audisset adquievit sermonibus eorum et tulit ephod et idola ac sculptile et cum eis profectus est
JUDG|18|21|qui cum pergerent et ante se ire fecissent parvulos et iumenta et omne quod erat pretiosum
JUDG|18|22|iamque a domo Michae essent procul viri qui habitabant in aedibus Michae conclamantes secuti sunt
JUDG|18|23|et post tergum clamare coeperunt qui cum respexissent dixerunt ad Micham quid tibi vis cur clamas
JUDG|18|24|qui respondit deos meos quos mihi feci tulistis et sacerdotem et omnia quae habeo et dicitis quid tibi est
JUDG|18|25|dixeruntque ei filii Dan cave ne ultra loquaris ad nos et veniant ad te viri animo concitati et ipse cum omni domo tua pereas
JUDG|18|26|et sic coepto itinere perrexerunt videns autem Micha quod fortiores se essent reversus est in domum suam
JUDG|18|27|sescenti autem viri tulerunt sacerdotem et quae supra diximus veneruntque in Lais ad populum quiescentem atque securum et percusserunt eos in ore gladii urbemque incendio tradiderunt
JUDG|18|28|nullo penitus ferente praesidium eo quod procul habitarent a Sidone et cum nullo hominum haberent quicquam societatis ac negotii erat autem civitas sita in regione Roob quam rursum extruentes habitaverunt in ea
JUDG|18|29|vocato nomine civitatis Dan iuxta vocabulum patris sui quem genuerat Israhel quae prius Lais dicebatur
JUDG|18|30|posueruntque sibi sculptile et Ionathan filium Gersan filii Mosi ac filios eius sacerdotes in tribu Dan usque ad diem captivitatis suae
JUDG|18|31|mansitque apud eos idolum Michae omni tempore quo fuit domus Dei in Silo in diebus illis non erat rex in Israhel
JUDG|19|1|fuit quidam vir Levites habitans in latere montis Ephraim qui accepit uxorem de Bethleem Iuda
JUDG|19|2|quae reliquit eum et reversa est in domum patris sui Bethleem mansitque apud eum quattuor mensibus
JUDG|19|3|secutusque est eam vir suus volens ei reconciliari atque blandiri et secum reducere habens in comitatu puerum et duos asinos quae suscepit eum et introduxit in domum patris sui quod cum audisset socer eius eumque vidisset occurrit ei laetus
JUDG|19|4|et amplexatus est hominem mansitque gener in domo soceri tribus diebus comedens cum eo et bibens familiariter
JUDG|19|5|die autem quarto de nocte consurgens proficisci voluit quem tenuit socer et ait ad eum gusta prius pauxillum panis et conforta stomachum et sic proficisceris
JUDG|19|6|sederuntque simul et comederunt ac biberunt dixitque pater puellae ad generum suum quaeso te ut hodie hic maneas pariterque laetemur
JUDG|19|7|at ille consurgens coepit velle proficisci et nihilominus obnixe eum socer tenuit et apud se fecit manere
JUDG|19|8|mane facto parabat Levites iter cui rursum socer oro te inquit ut paululum cibi capias et adsumptis viribus donec increscat dies postea proficiscaris comederunt ergo simul
JUDG|19|9|surrexitque adulescens ut pergeret cum uxore sua et puero cui rursum locutus est socer considera quod dies ad occasum declivior sit et propinquet ad vesperum mane apud me etiam hodie et duc laetum diem et cras proficisceris ut vadas in domum tuam
JUDG|19|10|noluit gener adquiescere sermonibus eius sed statim perrexit et venit contra Iebus quae altero nomine vocabatur Hierusalem ducens secum duos asinos onustos et concubinam
JUDG|19|11|iamque aderant iuxta Iebus et dies mutabatur in noctem dixitque puer ad dominum suum veni obsecro declinemus ad urbem Iebuseorum et maneamus in ea
JUDG|19|12|cui respondit dominus non ingrediar oppidum gentis alienae quae non est de filiis Israhel sed transibo usque Gabaa
JUDG|19|13|et cum illuc pervenero manebimus in ea aut certe in urbe Rama
JUDG|19|14|transierunt igitur Iebus et coeptum carpebant iter occubuitque eis sol iuxta Gabaa quae est in tribu Beniamin
JUDG|19|15|deverteruntque ad eam ut manerent ibi quo cum intrassent sedebant in platea civitatis et nullus eos recipere volebat hospitio
JUDG|19|16|et ecce apparuit homo senex revertens de agro et de opere suo vespere qui et ipse erat de monte Ephraim et peregrinus habitabat in Gabaa homines autem regionis illius erant filii Iemini
JUDG|19|17|elevatisque oculis vidit senex sedentem hominem cum sarcinulis suis in platea civitatis et dixit ad eum unde venis et quo vadis
JUDG|19|18|qui respondit ei profecti sumus de Bethleem Iuda et pergimus ad locum nostrum qui est in latere montis Ephraim unde ieramus Bethleem et nunc vadimus ad domum Dei nullusque nos sub tectum suum vult recipere
JUDG|19|19|habentes paleas et faenum in asinorum pabulum et panem ac vinum in meos et ancillae tuae usus et pueri qui mecum est nulla re indigemus nisi hospitio
JUDG|19|20|cui respondit senex pax tecum sit ego praebebo omnia quae necessaria sunt tantum quaeso ne in platea maneas
JUDG|19|21|introduxitque eum in domum suam et pabulum asinis praebuit ac postquam laverunt pedes suos recepit eos in convivium
JUDG|19|22|illis epulantibus et post laborem itineris cibo ac potu reficientibus corpora venerunt viri civitatis illius filii Belial id est absque iugo et circumdantes domum senis fores pulsare coeperunt clamantes ad dominum domus atque dicentes educ virum qui ingressus est domum tuam ut abutamur eo
JUDG|19|23|egressusque est ad eos senex et ait nolite fratres nolite facere malum hoc quia ingressus est homo hospitium meum et cessate ab hac stultitia
JUDG|19|24|habeo filiam virginem et hic homo habet concubinam educam eas ad vos ut humilietis eas et vestram libidinem conpleatis tantum obsecro ne scelus hoc contra naturam operemini in virum
JUDG|19|25|nolebant adquiescere sermonibus eius quod cernens homo eduxit ad eos concubinam suam et eis tradidit inludendam qua cum tota nocte abusi essent dimiserunt eam mane
JUDG|19|26|at mulier recedentibus tenebris venit ad ostium domus ubi manebat dominus suus et ibi corruit
JUDG|19|27|mane facto surrexit homo et aperuit ostium ut coeptam expleret viam et ecce concubina eius iacebat ante ostium sparsis in limine manibus
JUDG|19|28|cui ille putans eam quiescere loquebatur surge ut ambulemus qua nihil respondente intellegens quod erat tulit eam et inposuit asino reversusque est in domum suam
JUDG|19|29|quam cum esset ingressus arripuit gladium et cadaver uxoris cum ossibus suis in duodecim partes ac frusta concidens misit in omnes terminos Israhel
JUDG|19|30|quod cum vidissent singuli conclamabant numquam res talis facta est in Israhel ex eo die quo ascenderunt patres nostri de Aegypto usque in praesens tempus ferte sententiam et in commune decernite quid facto opus sit
JUDG|20|1|egressi sunt itaque omnes filii Israhel et pariter congregati quasi vir unus de Dan usque Bersabee et terra Galaad ad Dominum in Maspha
JUDG|20|2|omnesque anguli populorum et cunctae tribus Israhel in ecclesiam populi Dei convenerunt quadringenta milia peditum pugnatorum
JUDG|20|3|nec latuit filios Beniamin quod ascendissent filii Israhel in Maspha interrogatusque Levita maritus mulieris interfectae quomodo tantum scelus perpetratum esset
JUDG|20|4|respondit veni in Gabaa Beniamin cum uxore mea illucque deverti
JUDG|20|5|et ecce homines civitatis illius circumdederunt nocte domum in qua manebam volentes me occidere et uxorem meam incredibili libidinis furore vexantes denique mortua est
JUDG|20|6|quam arreptam in frusta concidi misique partes in omnes terminos possessionis vestrae quia numquam tantum nefas et tam grande piaculum factum est in Israhel
JUDG|20|7|adestis omnes filii Israhel decernite quid facere debeatis
JUDG|20|8|stansque omnis populus quasi unius hominis sermone respondit non recedemus in tabernacula nostra nec suam quisquam intrabit domum
JUDG|20|9|sed hoc contra Gabaa in commune faciemus
JUDG|20|10|decem viri eligantur e centum ex omnibus tribubus Israhel et centum de mille et mille de decem milibus ut conportent exercitui cibaria et possimus pugnantes contra Gabaa Beniamin reddere ei pro scelere quod meretur
JUDG|20|11|convenitque universus Israhel ad civitatem quasi unus homo eadem mente unoque consilio
JUDG|20|12|et miserunt nuntios ad omnem tribum Beniamin qui dicerent cur tantum nefas in vobis reppertum est
JUDG|20|13|tradite homines de Gabaa qui hoc flagitium perpetrarunt ut moriantur et auferatur malum de Israhel qui noluerunt fratrum suorum filiorum Israhel audire mandatum
JUDG|20|14|sed ex cunctis urbibus quae suae sortis erant convenerunt in Gabaa ut illis ferrent auxilium et contra universum Israhel populum dimicarent
JUDG|20|15|inventique sunt viginti quinque milia de Beniamin educentium gladium praeter habitatores Gabaa
JUDG|20|16|qui septingenti erant viri fortissimi ita sinistra ut dextra proeliantes et sic fundis ad certum iacientes lapides ut capillum quoque possent percutere et nequaquam in alteram partem ictus lapidis deferretur
JUDG|20|17|virorum quoque Israhel absque filiis Beniamin inventa sunt quadringenta milia educentium gladios et paratorum ad pugnam
JUDG|20|18|qui surgentes venerunt in domum Dei hoc est in Silo consulueruntque eum atque dixerunt quis erit in exercitu nostro princeps certaminis contra filios Beniamin quibus respondit Dominus Iudas sit dux vester
JUDG|20|19|statimque filii Israhel surgentes mane castrametati sunt iuxta Gabaa
JUDG|20|20|et inde procedentes ad pugnam contra Beniamin urbem obpugnare coeperunt
JUDG|20|21|egressique filii Beniamin de Gabaa occiderunt de filiis Israhel die illo viginti duo milia viros
JUDG|20|22|rursum filii Israhel et fortitudine et numero confidentes in eodem loco in quo prius certaverant aciem direxerunt
JUDG|20|23|ita tamen ut prius ascenderent et flerent coram Domino usque ad noctem consulerentque eum et dicerent debeo ultra procedere ad dimicandum contra filios Beniamin fratres meos an non quibus ille respondit ascendite ad eum et inite certamen
JUDG|20|24|cumque filii Israhel altero die contra Beniamin ad proelium processissent
JUDG|20|25|eruperunt filii Beniamin de portis Gabaa et occurrentes eis tanta in illos caede baccati sunt ut decem et octo milia virorum educentium gladium prosternerent
JUDG|20|26|quam ob rem omnes filii Israhel venerunt in domum Dei et sedentes flebant coram Domino ieiunaveruntque illo die usque ad vesperam et obtulerunt ei holocausta et pacificas victimas
JUDG|20|27|et super statu suo interrogaverunt eo tempore ibi erat arca foederis Dei
JUDG|20|28|et Finees filius Eleazari filii Aaron praepositus domus consuluerunt igitur Dominum atque dixerunt exire ultra debemus ad pugnam contra filios Beniamin fratres nostros an quiescere quibus ait Dominus ascendite cras enim tradam eos in manus vestras
JUDG|20|29|posueruntque filii Israhel insidias per circuitum urbis Gabaa
JUDG|20|30|et tertia vice sicut semel et bis contra Beniamin exercitum produxerunt
JUDG|20|31|sed et filii Beniamin audacter eruperunt de civitate et fugientes adversarios longius persecuti sunt ita ut vulnerarent ex eis sicut primo et secundo die et caederent per duas semitas terga vertentes quarum una ferebat in Bethel altera in Gabaa atque prosternerent triginta circiter viros
JUDG|20|32|putaverunt enim solito eos more cedere qui fugam arte simulantes iniere consilium ut abstraherent eos de civitate et quasi fugientes ad supradictas semitas perducerent
JUDG|20|33|omnes itaque filii Israhel surgentes de sedibus suis tetenderunt aciem in loco qui vocatur Baalthamar insidiae quoque quae circa urbem erant paulatim se aperire coeperunt
JUDG|20|34|et ab occidentali urbis parte procedere sed et alia decem milia virorum de universo Israhel habitatores urbis ad certamina provocabant ingravatumque est bellum contra filios Beniamin et non intellexerunt quod ex omni parte illis instaret interitus
JUDG|20|35|percussitque eos Dominus in conspectu filiorum Israhel et interfecerunt ex eis in illo die viginti quinque milia et centum viros omnes bellatores et educentes gladium
JUDG|20|36|filii autem Beniamin cum se inferiores esse vidissent coeperunt fugere quod cernentes filii Israhel dederunt eis ad fugiendum locum ut ad praeparatas insidias devenirent quas iuxta urbem posuerant
JUDG|20|37|qui cum repente de latibulis surrexissent et Beniamin terga caedentibus daret ingressi sunt civitatem et percusserunt eam in ore gladii
JUDG|20|38|signum autem dederant filii Israhel his quos in insidiis conlocaverant ut postquam urbem cepissent ignem accenderent et ascendente in altum fumo captam urbem demonstrarent
JUDG|20|39|quod cum cernerent filii Israhel in ipso certamine positi putaverunt enim filii Beniamin eos fugere et instantius sequebantur caesis de exercitu eorum triginta viris
JUDG|20|40|et viderent quasi columnam fumi de civitate conscendere Beniamin quoque retro aspiciens captam cerneret civitatem et flammas in sublime ferri
JUDG|20|41|qui prius simulaverant fugam versa facie fortius resistebant quod cum vidissent filii Beniamin in fugam versi sunt
JUDG|20|42|et ad viam deserti ire coeperunt illuc quoque eos adversariis persequentibus sed et hii qui urbem succenderant occurrerunt eis
JUDG|20|43|atque ita factum est ut ex utraque parte ab hostibus caederentur nec erat ulla morientium requies ceciderunt atque prostrati sunt ad orientalem plagam urbis Gabaa
JUDG|20|44|fuerunt autem qui in eodem loco interfecti sunt decem et octo milia virorum omnes robustissimi pugnatores
JUDG|20|45|quod cum vidissent qui remanserant de Beniamin fugerunt in solitudinem et pergebant ad petram cuius vocabulum est Remmon in illa quoque fuga palantes et in diversa tendentes occiderunt quinque milia viros et cum ultra tenderent persecuti sunt eos et interfecerunt etiam alios duo milia
JUDG|20|46|et sic factum est ut omnes qui ceciderant de Beniamin in diversis locis essent viginti quinque milia pugnatores ad bella promptissimi
JUDG|20|47|remanserunt itaque de omni numero Beniamin qui evadere potuerant et fugere in solitudinem sescenti viri sederuntque in petra Remmon mensibus quattuor
JUDG|20|48|regressi autem filii Israhel omnes reliquias civitatis a viris usque ad iumenta gladio percusserunt cunctasque urbes et viculos Beniamin vorax flamma consumpsit
JUDG|21|1|iuraverunt quoque filii Israhel in Maspha et dixerunt nullus nostrum dabit filiis Beniamin de filiabus suis uxorem
JUDG|21|2|veneruntque omnes ad domum Dei in Silo et in conspectu eius sedentes usque ad vesperam levaverunt vocem et magno ululatu coeperunt flere dicentes
JUDG|21|3|quare Domine Deus Israhel factum est hoc malum in populo tuo ut hodie una tribus auferretur ex nobis
JUDG|21|4|altera autem die diluculo consurgentes extruxerunt altare obtuleruntque ibi holocausta et pacificas victimas et dixerunt
JUDG|21|5|quis non ascendit in exercitu Domini de universis tribubus Israhel grandi enim se iuramento constrinxerant cum essent in Maspha interfici eos qui defuissent
JUDG|21|6|ductique paenitentia filii Israhel super fratre suo Beniamin coeperunt dicere ablata est una tribus de Israhel
JUDG|21|7|unde uxores accipient omnes enim in commune iuravimus non daturos nos his filias nostras
JUDG|21|8|idcirco dixerunt quis est de universis tribubus Israhel qui non ascendit ad Dominum in Maspha et ecce inventi sunt habitatores Iabisgalaad in illo exercitu non fuisse
JUDG|21|9|eo quoque tempore cum essent in Silo nullus ex eis ibi reppertus est
JUDG|21|10|miserunt itaque decem milia viros robustissimos et praeceperunt eis ite et percutite habitatores Iabisgalaad in ore gladii tam uxores quam parvulos eorum
JUDG|21|11|et hoc erit quod observare debetis omne generis masculini et mulieres quae cognoverunt viros interficite
JUDG|21|12|inventaeque sunt de Iabisgalaad quadringentae virgines quae nescierunt viri torum et adduxerunt eas in castra in Silo in terra Chanaan
JUDG|21|13|miseruntque nuntios ad filios Beniamin qui erant in petra Remmon et praeceperunt eis ut eos in pace susciperent
JUDG|21|14|veneruntque filii Beniamin in illo tempore et datae sunt eis uxores de filiabus Iabisgalaad alias autem non reppererunt quas simili modo traderent
JUDG|21|15|universusque Israhel valde doluit et egit paenitudinem super interfectione unius tribus ex Israhel
JUDG|21|16|dixeruntque maiores natu quid faciemus reliquis qui non acceperunt uxores omnes in Beniamin feminae conciderunt
JUDG|21|17|et magna nobis cura ingentique studio providendum est ne una tribus deleatur ex Israhel
JUDG|21|18|filias nostras eis dare non possumus constricti iuramento et maledictione qua diximus maledictus qui dederit de filiabus suis uxorem Beniamin
JUDG|21|19|ceperuntque consilium atque dixerunt ecce sollemnitas Domini est in Silo anniversaria quae sita est ad septentrionem urbis Bethel et ad orientalem plagam viae quae de Bethel tendit ad Sycimam et ad meridiem oppidi Lebona
JUDG|21|20|praeceperuntque filiis Beniamin atque dixerunt ite et latete in vineis
JUDG|21|21|cumque videritis filias Silo ad ducendos choros ex more procedere exite repente de vineis et rapite eas singuli uxores singulas et pergite in terram Beniamin
JUDG|21|22|cumque venerint patres earum ac fratres et adversum vos queri coeperint atque iurgari dicemus eis miseremini eorum non enim rapuerunt eas iure bellantium atque victorum sed rogantibus ut acciperent non dedistis et a vestra parte peccatum est
JUDG|21|23|feceruntque filii Beniamin ut sibi fuerat imperatum et iuxta numerum suum rapuerunt sibi de his quae ducebant choros uxores singulas abieruntque in possessionem suam aedificantes urbes et habitantes in eis
JUDG|21|24|filii quoque Israhel reversi sunt per tribus et familias in tabernacula sua in diebus illis non erat rex in Israhel sed unusquisque quod sibi rectum videbatur hoc faciebat
RUTH|1|1|in diebus unius iudicis quando iudices praeerant facta est fames in terra abiitque homo de Bethleem Iuda ut peregrinaretur in regione moabitide cum uxore sua ac duobus liberis
RUTH|1|2|ipse vocabatur Helimelech uxor eius Noemi e duobus filiis alter Maalon et alter Chellion Ephrathei de Bethleem Iuda ingressique regionem moabitidem morabantur ibi
RUTH|1|3|et mortuus est Helimelech maritus Noemi remansitque ipsa cum filiis
RUTH|1|4|qui acceperunt uxores moabitidas quarum una vocabatur Orpha altera Ruth manseruntque ibi decem annis
RUTH|1|5|et ambo mortui sunt Maalon videlicet et Chellion remansitque mulier orbata duobus liberis ac marito
RUTH|1|6|et surrexit ut in patriam pergeret cum utraque nuru sua de regione moabitide audierat enim quod respexisset Dominus populum suum et dedisset eis escas
RUTH|1|7|egressa est itaque de loco peregrinationis suae cum utraque nuru et iam in via posita revertendi in terram Iuda
RUTH|1|8|dixit ad eas ite in domum matris vestrae faciat Dominus vobiscum misericordiam sicut fecistis cum mortuis et mecum
RUTH|1|9|det vobis invenire requiem in domibus virorum quos sortiturae estis et osculata est eas quae elevata voce flere coeperunt
RUTH|1|10|et dicere tecum pergemus ad populum tuum
RUTH|1|11|quibus illa respondit revertimini filiae mi cur venitis mecum num ultra habeo filios in utero meo ut viros ex me sperare possitis
RUTH|1|12|revertimini filiae mi abite iam enim senectute confecta sum nec apta vinculo coniugali etiam si possem hac nocte concipere et parere filios
RUTH|1|13|si eos expectare velitis donec crescant et annos impleant pubertatis ante eritis vetulae quam nubatis nolite quaeso filiae mi quia vestra angustia me magis premit et egressa est manus Domini contra me
RUTH|1|14|elevata igitur voce rursum flere coeperunt Orpha osculata socrum est ac reversa Ruth adhesit socrui suae
RUTH|1|15|cui dixit Noemi en reversa est cognata tua ad populum suum et ad deos suos vade cum ea
RUTH|1|16|quae respondit ne adverseris mihi ut relinquam te et abeam quocumque perrexeris pergam ubi morata fueris et ego pariter morabor populus tuus populus meus et Deus tuus Deus meus
RUTH|1|17|quae te morientem terra susceperit in ea moriar ibique locum accipiam sepulturae haec mihi faciat Deus et haec addat si non sola mors me et te separaverit
RUTH|1|18|videns ergo Noemi quod obstinato Ruth animo decrevisset secum pergere adversari noluit nec ultra ad suos reditum persuadere
RUTH|1|19|profectaeque sunt simul et venerunt in Bethleem quibus urbem ingressis velox apud cunctos fama percrebuit dicebantque mulieres haec est illa Noemi
RUTH|1|20|quibus ait ne vocetis me Noemi id est pulchram sed vocate me Mara hoc est amaram quia valde me amaritudine replevit Omnipotens
RUTH|1|21|egressa sum plena et vacuam reduxit me Dominus cur igitur vocatis me Noemi quam humiliavit Dominus et adflixit Omnipotens
RUTH|1|22|venit ergo Noemi cum Ruth Moabitide nuru sua de terra peregrinationis suae ac reversa est in Bethleem quando primum hordea metebantur
RUTH|2|1|erat autem vir Helimelech consanguineus homo potens et magnarum opum nomine Booz
RUTH|2|2|dixitque Ruth Moabitis ad socrum suam si iubes vadam in agrum et colligam spicas quae metentium fugerint manus ubicumque clementis in me patris familias repperero gratiam cui illa respondit vade filia mi
RUTH|2|3|abiit itaque et colligebat spicas post terga metentium accidit autem ut ager ille haberet dominum Booz qui erat de cognatione Helimelech
RUTH|2|4|et ecce ipse veniebat de Bethleem dixitque messoribus Dominus vobiscum qui responderunt ei benedicat tibi Dominus
RUTH|2|5|dixitque Booz iuveni qui messoribus praeerat cuius est haec puella
RUTH|2|6|qui respondit haec est Moabitis quae venit cum Noemi de regione moabitide
RUTH|2|7|et rogavit ut spicas colligeret remanentes sequens messorum vestigia et de mane usque nunc stat in agro et ne ad momentum quidem domum reversa est
RUTH|2|8|et ait Booz ad Ruth audi filia ne vadas ad colligendum in alterum agrum nec recedas ab hoc loco sed iungere puellis meis
RUTH|2|9|et ubi messuerint sequere mandavi enim pueris meis ut nemo tibi molestus sit sed etiam si sitieris vade ad sarcinulas et bibe aquas de quibus et pueri bibunt
RUTH|2|10|quae cadens in faciem suam et adorans super terram dixit ad eum unde mihi hoc ut invenirem gratiam ante oculos tuos et nosse me dignareris peregrinam mulierem
RUTH|2|11|cui ille respondit nuntiata sunt mihi omnia quae feceris socrui tuae post mortem viri tui et quod dereliqueris parentes tuos et terram in qua nata es et veneris ad populum quem ante nesciebas
RUTH|2|12|reddat tibi Dominus pro opere tuo et plenam mercedem recipias a Domino Deo Israhel ad quem venisti et sub cuius confugisti alas
RUTH|2|13|quae ait inveni gratiam ante oculos tuos domine mi qui consolatus es me et locutus es ad cor ancillae tuae quae non sum similis unius puellarum tuarum
RUTH|2|14|dixitque ad eam Booz quando hora vescendi fuerit veni huc et comede panem et intingue buccellam tuam in aceto sedit itaque ad messorum latus et congessit pulentam sibi comeditque et saturata est et tulit reliquias
RUTH|2|15|atque inde surrexit ut spicas ex more colligeret praecepit autem Booz pueris suis dicens etiam si vobiscum metere voluerit ne prohibeatis eam
RUTH|2|16|et de vestris quoque manipulis proicite de industria et remanere permittite ut absque rubore colligat et colligentem nemo corripiat
RUTH|2|17|collegit ergo in agro usque ad vesperam et quae collegerat virga caedens et excutiens invenit hordei quasi oephi mensuram id est tres modios
RUTH|2|18|quos portans reversa est in civitatem et ostendit socrui suae insuper protulit et dedit ei de reliquiis cibi sui quo saturata fuerat
RUTH|2|19|dixitque ei socrus ubi hodie collegisti et ubi fecisti opus sit benedictus qui misertus est tui indicavitque ei apud quem esset operata et nomen dixit viri quod Booz vocaretur
RUTH|2|20|cui respondit Noemi benedictus sit a Domino quoniam eandem gratiam quam praebuerat vivis servavit et mortuis rursumque propinquus ait noster est homo
RUTH|2|21|et Ruth hoc quoque inquit praecepit mihi ut tamdiu messoribus eius iungerer donec omnes segetes meterentur
RUTH|2|22|cui dixit socrus melius est filia mi ut cum puellis eius exeas ad metendum ne in alieno agro quispiam resistat tibi
RUTH|2|23|iuncta est itaque puellis Booz et tamdiu cum eis messuit donec hordea et triticum in horreis conderentur
RUTH|3|1|postquam autem reversa est ad socrum suam audivit ab ea filia mi quaeram tibi requiem et providebo ut bene sit tibi
RUTH|3|2|Booz iste cuius puellis in agro iuncta es propinquus est noster et hac nocte aream hordei ventilat
RUTH|3|3|lava igitur et unguere et induere cultioribus vestimentis ac descende in aream non te videat homo donec esum potumque finierit
RUTH|3|4|quando autem ierit ad dormiendum nota locum in quo dormiat veniesque et discoperies pallium quo operitur a parte pedum et proicies te et ibi iacebis ipse autem dicet tibi quid agere debeas
RUTH|3|5|quae respondit quicquid praeceperis faciam
RUTH|3|6|descenditque in aream et fecit omnia quae sibi imperaverat socrus
RUTH|3|7|cumque comedisset Booz et bibisset et factus esset hilarior issetque ad dormiendum iuxta acervum manipulorum venit abscondite et discoperto a pedibus eius pallio se proiecit
RUTH|3|8|et ecce nocte iam media expavit homo et conturbatus est viditque mulierem iacentem ad pedes suos
RUTH|3|9|et ait illi quae es illaque respondit ego sum Ruth ancilla tua expande pallium tuum super famulam tuam quia propinquus es
RUTH|3|10|et ille benedicta inquit es Domino filia et priorem misericordiam posteriore superasti quia non es secuta iuvenes pauperes sive divites
RUTH|3|11|noli ergo metuere sed quicquid dixeris mihi faciam tibi scit enim omnis populus qui habitat intra portas urbis meae mulierem te esse virtutis
RUTH|3|12|nec abnuo me propinquum sed est alius me propinquior
RUTH|3|13|quiesce hac nocte et facto mane si te voluerit propinquitatis iure retinere bene res acta est sin autem ille noluerit ego te absque ulla dubitatione suscipiam vivit Dominus dormi usque mane
RUTH|3|14|dormivit itaque ad pedes eius usque ad noctis abscessum surrexitque antequam homines se cognoscerent mutuo et dixit Booz cave ne quis noverit quod huc veneris
RUTH|3|15|et rursum expande inquit palliolum tuum quo operiris et tene utraque manu qua extendente et tenente mensus est sex modios hordei et posuit super eam quae portans ingressa est civitatem
RUTH|3|16|et venit ad socrum suam quae dixit ei quid egisti filia narravitque ei omnia quae sibi fecisset homo
RUTH|3|17|et ait ecce sex modios hordei dedit mihi et ait nolo vacuam te reverti ad socrum tuam
RUTH|3|18|dixitque Noemi expecta filia donec videamus quem res exitum habeat neque enim cessabit homo nisi conpleverit quod locutus est
RUTH|4|1|ascendit ergo Booz ad portam et sedit ibi cumque vidisset propinquum praeterire de quo prius sermo habitus est dixit ad eum declina paulisper et sede hic vocans eum nomine suo qui devertit et sedit
RUTH|4|2|tollens autem Booz decem viros de senioribus civitatis dixit ad eos sedete hic
RUTH|4|3|quibus residentibus locutus est ad propinquum partem agri fratris nostri Helimelech vendit Noemi quae reversa est de regione moabitide
RUTH|4|4|quod audire te volui et tibi dicere coram cunctis sedentibus et maioribus natu de populo meo si vis possidere iure propinquitatis eme et posside sin autem tibi displicet hoc ipsum indica mihi ut sciam quid facere debeam nullus est enim propinquus excepto te qui prior es et me qui secundus sum at ille respondit ego agrum emam
RUTH|4|5|cui dixit Booz quando emeris agrum de manu mulieris Ruth quoque Moabitidem quae uxor defuncti fuit debes accipere ut suscites nomen propinqui tui in hereditate sua
RUTH|4|6|qui respondit cedo iure propinquitatis neque enim posteritatem familiae meae delere debeo tu meo utere privilegio quo me libenter carere profiteor
RUTH|4|7|hic autem erat mos antiquitus in Israhel inter propinquos et si quando alter alteri suo iure cedebat ut esset firma concessio solvebat homo calciamentum suum et dabat proximo suo hoc erat testimonium cessionis in Israhel
RUTH|4|8|dixit ergo propinquus Booz tolle calciamentum quod statim solvit de pede suo
RUTH|4|9|at ille maioribus natu et universo populo testes inquit vos estis hodie quod possederim omnia quae fuerunt Helimelech et Chellion et Maalon tradente Noemi
RUTH|4|10|et Ruth Moabitidem uxorem Maalon in coniugium sumpserim ut suscitem nomen defuncti in hereditate sua ne vocabulum eius de familia sua ac fratribus et populo deleatur vos inquam huius rei testes estis
RUTH|4|11|respondit omnis populus qui erat in porta et maiores natu nos testes sumus faciat Dominus hanc mulierem quae ingreditur domum tuam sicut Rachel et Liam quae aedificaverunt domum Israhel ut sit exemplum virtutis in Ephrata et habeat celebre nomen in Bethleem
RUTH|4|12|fiatque domus tua sicut domus Phares quem Thamar peperit Iudae de semine quod dederit Dominus tibi ex hac puella
RUTH|4|13|tulit itaque Booz Ruth et accepit uxorem ingressusque est ad eam et dedit illi Dominus ut conciperet et pareret filium
RUTH|4|14|dixeruntque mulieres ad Noemi benedictus Dominus qui non est passus ut deficeret successor familiae tuae et vocaretur nomen eius in Israhel
RUTH|4|15|et habeas qui consoletur animam tuam et enutriat senectutem de nuru enim tua natus est quae te diligit et multo tibi est melior quam si septem haberes filios
RUTH|4|16|susceptumque Noemi puerum posuit in sinu suo et nutricis ac gerulae officio fungebatur
RUTH|4|17|vicinae autem mulieres congratulantes ei et dicentes natus est filius Noemi vocaverunt nomen eius Obed hic est pater Isai patris David
RUTH|4|18|hae sunt generationes Phares Phares genuit Esrom
RUTH|4|19|Esrom genuit Aram Aram genuit Aminadab
RUTH|4|20|Aminadab genuit Naasson Naasson genuit Salma
RUTH|4|21|Salma genuit Booz Booz genuit Obed
1SAM|1|1|fuit vir unus de Ramathaimsophim de monte Ephraim et nomen eius Helcana filius Hieroam filii Heliu filii Thau filii Suph Ephratheus
1SAM|1|2|et habuit duas uxores nomen uni Anna et nomen secundae Fenenna fueruntque Fenennae filii Annae autem non erant liberi
1SAM|1|3|et ascendebat vir ille de civitate sua statutis diebus ut adoraret et sacrificaret Domino exercituum in Silo erant autem ibi duo filii Heli Ofni et Finees sacerdotes Domini
1SAM|1|4|venit ergo dies et immolavit Helcana deditque Fenennae uxori suae et cunctis filiis eius et filiabus partes
1SAM|1|5|Annae autem dedit partem unam tristis quia Annam diligebat Dominus autem concluserat vulvam eius
1SAM|1|6|adfligebat quoque eam aemula eius et vehementer angebat in tantum ut exprobraret quod conclusisset Dominus vulvam eius
1SAM|1|7|sicque faciebat per singulos annos cum redeunte tempore ascenderent templum Domini et sic provocabat eam porro illa flebat et non capiebat cibum
1SAM|1|8|dixit ergo ei Helcana vir suus Anna cur fles et quare non comedis et quam ob rem adfligitur cor tuum numquid non ego melior sum tibi quam decem filii
1SAM|1|9|surrexit autem Anna postquam comederat in Silo et biberat et Heli sacerdote sedente super sellam ante postes templi Domini
1SAM|1|10|cum esset amaro animo oravit Dominum flens largiter
1SAM|1|11|et votum vovit dicens Domine exercituum si respiciens videris adflictionem famulae tuae et recordatus mei fueris nec oblitus ancillae tuae dederisque servae tuae sexum virilem dabo eum Domino omnes dies vitae eius et novacula non ascendet super caput eius
1SAM|1|12|factum est ergo cum illa multiplicaret preces coram Domino ut Heli observaret os eius
1SAM|1|13|porro Anna loquebatur in corde suo tantumque labia illius movebantur et vox penitus non audiebatur aestimavit igitur eam Heli temulentam
1SAM|1|14|dixitque ei usquequo ebria eris digere paulisper vinum quo mades
1SAM|1|15|respondens Anna nequaquam inquit domine mi nam mulier infelix nimis ego sum vinumque et omne quod inebriare potest non bibi sed effudi animam meam in conspectu Domini
1SAM|1|16|ne reputes ancillam tuam quasi unam de filiabus Belial quia ex multitudine doloris et maeroris mei locuta sum usque in praesens
1SAM|1|17|tunc Heli ait ei vade in pace et Deus Israhel det tibi petitionem quam rogasti eum
1SAM|1|18|et illa dixit utinam inveniat ancilla tua gratiam in oculis tuis et abiit mulier in viam suam et comedit vultusque eius non sunt amplius in diversa mutati
1SAM|1|19|et surrexerunt mane et adoraverunt coram Domino reversique sunt et venerunt in domum suam Ramatha cognovit autem Helcana Annam uxorem suam et recordatus est eius Dominus
1SAM|1|20|et factum est post circulum dierum concepit Anna et peperit filium vocavitque nomen eius Samuhel eo quod a Domino postulasset eum
1SAM|1|21|ascendit autem vir Helcana et omnis domus eius ut immolaret Domino hostiam sollemnem et votum suum
1SAM|1|22|et Anna non ascendit dixit enim viro suo non vadam donec ablactetur infans et ducam eum et appareat ante conspectum Domini et maneat ibi iugiter
1SAM|1|23|et ait ei Helcana vir suus fac quod bonum tibi videtur et mane donec ablactes eum precorque ut impleat Dominus verbum suum mansit ergo mulier et lactavit filium suum donec amoveret eum a lacte
1SAM|1|24|et adduxit eum secum postquam ablactaverat in vitulis tribus et tribus modiis farinae et amphora vini et adduxit eum ad domum Domini in Silo puer autem erat adhuc infantulus
1SAM|1|25|et immolaverunt vitulum et obtulerunt puerum Heli
1SAM|1|26|et ait obsecro mi domine vivit anima tua domine ego sum illa mulier quae steti coram te hic orans Dominum
1SAM|1|27|pro puero isto oravi et dedit Dominus mihi petitionem meam quam postulavi eum
1SAM|1|28|idcirco et ego commodavi eum Domino cunctis diebus quibus fuerit accommodatus Domino et adoraverunt ibi Dominum et oravit Anna et ait
1SAM|2|1|exultavit cor meum in Domino exaltatum est cornu meum in Domino dilatatum est os meum super inimicos meos quia laetata sum in salutari tuo
1SAM|2|2|non est sanctus ut est Dominus neque enim est alius extra te et non est fortis sicut Deus noster
1SAM|2|3|nolite multiplicare loqui sublimia gloriantes recedant vetera de ore vestro quoniam Deus scientiarum Dominus est et ipsi praeparantur cogitationes
1SAM|2|4|arcus fortium superatus est et infirmi accincti sunt robore
1SAM|2|5|saturati prius pro pane se locaverunt et famelici saturati sunt donec sterilis peperit plurimos et quae multos habebat filios infirmata est
1SAM|2|6|Dominus mortificat et vivificat deducit ad infernum et reducit
1SAM|2|7|Dominus pauperem facit et ditat humiliat et sublevat
1SAM|2|8|suscitat de pulvere egenum et de stercore elevat pauperem ut sedeat cum principibus et solium gloriae teneat Domini enim sunt cardines terrae et posuit super eos orbem
1SAM|2|9|pedes sanctorum suorum servabit et impii in tenebris conticescent quia non in fortitudine roborabitur vir
1SAM|2|10|Dominum formidabunt adversarii eius super ipsos in caelis tonabit Dominus iudicabit fines terrae et dabit imperium regi suo et sublimabit cornu christi sui
1SAM|2|11|et abiit Helcana Ramatha in domum suam puer autem erat minister in conspectu Domini ante faciem Heli sacerdotis
1SAM|2|12|porro filii Heli filii Belial nescientes Dominum
1SAM|2|13|neque officium sacerdotum ad populum sed quicumque immolasset victimam veniebat puer sacerdotis dum coquerentur carnes et habebat fuscinulam tridentem in manu sua
1SAM|2|14|et mittebat eam in lebetem vel in caldariam aut in ollam sive in caccabum et omne quod levabat fuscinula tollebat sacerdos sibi sic faciebant universo Israheli venientium in Silo
1SAM|2|15|etiam antequam adolerent adipem veniebat puer sacerdotis et dicebat immolanti da mihi carnem ut coquam sacerdoti non enim accipiam a te carnem coctam sed crudam
1SAM|2|16|dicebatque illi immolans incendatur primum iuxta morem hodie adeps et tolle tibi quantumcumque desiderat anima tua qui respondens aiebat ei nequaquam nunc enim dabis alioquin tollam vi
1SAM|2|17|erat ergo peccatum puerorum grande nimis coram Domino quia detrahebant homines sacrificio Domini
1SAM|2|18|Samuhel autem ministrabat ante faciem Domini puer accinctus ephod lineo
1SAM|2|19|et tunicam parvam faciebat ei mater sua quam adferebat statutis diebus ascendens cum viro suo ut immolaret hostiam sollemnem
1SAM|2|20|et benedixit Heli Helcanae et uxori eius dixitque reddat Dominus tibi semen de muliere hac pro fenore quod commodasti Domino et abierunt in locum suum
1SAM|2|21|visitavit ergo Dominus Annam et concepit et peperit tres filios et duas filias et magnificatus est puer Samuhel apud Dominum
1SAM|2|22|Heli autem erat senex valde et audivit omnia quae faciebant filii sui universo Israheli et quomodo dormiebant cum mulieribus quae observabant ad ostium tabernaculi
1SAM|2|23|et dixit eis quare facitis res huiuscemodi quas ego audio res pessimas ab omni populo
1SAM|2|24|nolite filii mi non enim est bona fama quam ego audio ut transgredi faciatis populum Domini
1SAM|2|25|si peccaverit vir in virum placari ei potest Deus si autem in Domino peccaverit vir quis orabit pro eo et non audierunt vocem patris sui quia voluit Dominus occidere eos
1SAM|2|26|puer autem Samuhel proficiebat atque crescebat et placebat tam Deo quam hominibus
1SAM|2|27|venit autem vir Dei ad Heli et ait ad eum haec dicit Dominus numquid non aperte revelatus sum domui patris tui cum essent in Aegypto in domo Pharaonis
1SAM|2|28|et elegi eum ex omnibus tribubus Israhel mihi in sacerdotem ut ascenderet altare meum et adoleret mihi incensum et portaret ephod coram me et dedi domui patris tui omnia de sacrificiis filiorum Israhel
1SAM|2|29|quare calce abicitis victimam meam et munera mea quae praecepi ut offerrentur in templo et magis honorasti filios tuos quam me ut comederetis primitias omnis sacrificii Israhel populi mei
1SAM|2|30|propterea ait Dominus Deus Israhel loquens locutus sum ut domus tua et domus patris tui ministraret in conspectu meo usque in sempiternum nunc autem dicit Dominus absit hoc a me sed quicumque glorificaverit me glorificabo eum qui autem contemnunt me erunt ignobiles
1SAM|2|31|ecce dies veniunt et praecidam brachium tuum et brachium domus patris tui ut non sit senex in domo tua
1SAM|2|32|et videbis aemulum tuum in templo in universis prosperis Israhel et non erit senex in domo tua omnibus diebus
1SAM|2|33|verumtamen non auferam penitus virum ex te ab altari meo sed ut deficiant oculi tui et tabescat anima tua et pars magna domus tuae morietur cum ad virilem aetatem venerit
1SAM|2|34|hoc autem erit tibi signum quod venturum est duobus filiis tuis Ofni et Finees in die uno morientur ambo
1SAM|2|35|et suscitabo mihi sacerdotem fidelem qui iuxta cor meum et animam meam faciat et aedificabo ei domum fidelem et ambulabit coram christo meo cunctis diebus
1SAM|2|36|futurum est autem ut quicumque remanserit in domo tua veniat ut oretur pro eo et offerat nummum argenteum et tortam panis dicatque dimitte me obsecro ad unam partem sacerdotalem ut comedam buccellam panis
1SAM|3|1|puer autem Samuhel ministrabat Domino coram Heli et sermo Domini erat pretiosus in diebus illis non erat visio manifesta
1SAM|3|2|factum est ergo in die quadam Heli iacebat in loco suo et oculi eius caligaverant nec poterat videre
1SAM|3|3|lucerna Dei antequam extingueretur Samuhel autem dormiebat in templo Domini ubi erat arca Dei
1SAM|3|4|et vocavit Dominus Samuhel qui respondens ait ecce ego
1SAM|3|5|et cucurrit ad Heli et dixit ecce ego vocasti enim me qui dixit non vocavi revertere dormi et abiit et dormivit
1SAM|3|6|et adiecit Dominus vocare rursum Samuhel consurgensque Samuhel abiit ad Heli et dixit ecce ego quia vocasti me qui respondit non vocavi te fili mi revertere et dormi
1SAM|3|7|porro Samuhel necdum sciebat Dominum neque revelatus fuerat ei sermo Domini
1SAM|3|8|et adiecit Dominus et vocavit adhuc Samuhel tertio qui consurgens abiit ad Heli
1SAM|3|9|et ait ecce ego quia vocasti me intellexit igitur Heli quia Dominus vocaret puerum et ait ad Samuhel vade et dormi et si deinceps vocaverit te dices loquere Domine quia audit servus tuus abiit ergo Samuhel et dormivit in loco suo
1SAM|3|10|et venit Dominus et stetit et vocavit sicut vocaverat secundo Samuhel Samuhel et ait Samuhel loquere quia audit servus tuus
1SAM|3|11|et dixit Dominus ad Samuhel ecce ego facio verbum in Israhel quod quicumque audierit tinnient ambae aures eius
1SAM|3|12|in die illo suscitabo adversum Heli omnia quae locutus sum super domum eius incipiam et conplebo
1SAM|3|13|praedixi enim ei quod iudicaturus essem domum eius in aeternum propter iniquitatem eo quod noverat indigne agere filios suos et non corripuit eos
1SAM|3|14|idcirco iuravi domui Heli quod non expietur iniquitas domus eius victimis et muneribus usque in aeternum
1SAM|3|15|dormivit autem Samuhel usque mane aperuitque ostia domus Domini et Samuhel timebat indicare visionem Heli
1SAM|3|16|vocavit ergo Heli Samuhelem et dixit Samuhel fili mi qui respondens ait praesto sum
1SAM|3|17|et interrogavit eum quis est sermo quem locutus est ad te oro te ne celaveris me haec faciat tibi Deus et haec addat si absconderis a me sermonem ex omnibus verbis quae dicta sunt tibi
1SAM|3|18|indicavit itaque ei Samuhel universos sermones et non abscondit ab eo et ille respondit Dominus est quod bonum est in oculis suis faciat
1SAM|3|19|crevit autem Samuhel et Dominus erat cum eo et non cecidit ex omnibus verbis eius in terram
1SAM|3|20|et cognovit universus Israhel a Dan usque Bersabee quod fidelis Samuhel propheta esset Domini
1SAM|3|21|et addidit Dominus ut appareret in Silo quoniam revelatus fuerat Dominus Samuheli in Silo iuxta verbum Domini et evenit sermo Samuhelis universo Israheli
1SAM|4|1|egressus est namque Israhel obviam Philisthim in proelium et castrametatus est iuxta lapidem Adiutorii porro Philisthim venerunt in Afec
1SAM|4|2|et instruxerunt aciem contra Israhel inito autem certamine terga vertit Israhel Philistheis et caesa sunt in illo certamine passim per agros quasi quattuor milia virorum
1SAM|4|3|et reversus est populus ad castra dixeruntque maiores natu de Israhel quare percussit nos Dominus hodie coram Philisthim adferamus ad nos de Silo arcam foederis Domini et veniat in medium nostri ut salvet nos de manu inimicorum nostrorum
1SAM|4|4|misit ergo populus in Silo et tulerunt inde arcam foederis Domini exercituum sedentis super cherubin erantque duo filii Heli cum arca foederis Domini Ofni et Finees
1SAM|4|5|cumque venisset arca foederis Domini in castra vociferatus est omnis Israhel clamore grandi et personuit terra
1SAM|4|6|et audierunt Philisthim vocem clamoris dixeruntque quaenam haec est vox clamoris magni in castris Hebraeorum et cognoverunt quod arca Domini venisset in castra
1SAM|4|7|timueruntque Philisthim dicentes venit Deus in castra et ingemuerunt
1SAM|4|8|vae nobis non enim fuit tanta exultatio heri et nudius tertius vae nobis quis nos servabit de manu deorum sublimium istorum hii sunt dii qui percusserunt Aegyptum omni plaga in deserto
1SAM|4|9|confortamini et estote viri Philisthim ne serviatis Hebraeis sicut illi servierunt vobis confortamini et bellate
1SAM|4|10|pugnaverunt ergo Philisthim et caesus est Israhel et fugit unusquisque in tabernaculum suum et facta est plaga magna nimis et ceciderunt de Israhel triginta milia peditum
1SAM|4|11|et arca Dei capta est duoque filii Heli mortui sunt Ofni et Finees
1SAM|4|12|currens autem vir de Beniamin ex acie venit in Silo in die illo scissa veste et conspersus pulvere caput
1SAM|4|13|cumque ille venisset Heli sedebat super sellam contra viam aspectans erat enim cor eius pavens pro arca Domini vir autem ille postquam ingressus est nuntiavit urbi et ululavit omnis civitas
1SAM|4|14|et audivit Heli sonitum clamoris dixitque quis est hic sonitus tumultus huius at ille festinavit et venit et adnuntiavit Heli
1SAM|4|15|Heli autem erat nonaginta et octo annorum et oculi eius caligaverant et videre non poterat
1SAM|4|16|et dixit ad Heli ego sum qui veni de proelio et ego qui de acie fugi hodie cui ille ait quid actum est fili mi
1SAM|4|17|respondens autem qui nuntiabat fugit inquit Israhel coram Philisthim et ruina magna facta est in populo insuper et duo filii tui mortui sunt Ofni et Finees et arca Dei capta est
1SAM|4|18|cumque ille nominasset arcam Dei cecidit de sella retrorsum iuxta ostium et fractis cervicibus mortuus est senex enim erat vir et grandevus et ipse iudicavit Israhel quadraginta annis
1SAM|4|19|nurus autem eius uxor Finees praegnans erat vicinaque partui et audito nuntio quod capta esset arca Dei et mortuus socer suus et vir suus incurvavit se et peperit inruerant enim in eam dolores subiti
1SAM|4|20|in ipso autem momento mortis eius dixerunt ei quae stabant circa eam ne timeas quia filium peperisti quae non respondit eis neque animadvertit
1SAM|4|21|et vocavit puerum Hicabod dicens translata est gloria de Israhel quia capta est arca Dei et pro socero suo et pro viro suo
1SAM|4|22|et ait translata est gloria ab Israhel eo quod capta esset arca Dei
1SAM|5|1|Philisthim autem tulerunt arcam Dei et asportaverunt eam a lapide Adiutorii in Azotum
1SAM|5|2|tulerunt Philisthim arcam Dei et intulerunt eam in templum Dagon et statuerunt eam iuxta Dagon
1SAM|5|3|cumque surrexissent diluculo Azotii altera die ecce Dagon iacebat pronus in terram ante arcam Domini et tulerunt Dagon et restituerunt eum in loco suo
1SAM|5|4|rursumque mane die alio consurgentes invenerunt Dagon iacentem super faciem suam in terram coram arca Domini caput autem Dagon et duae palmae manuum eius abscisae erant super limen
1SAM|5|5|porro Dagon truncus solus remanserat in loco suo propter hanc causam non calcant sacerdotes Dagon et omnes qui ingrediuntur templum eius super limen Dagon in Azoto usque in hodiernum diem
1SAM|5|6|adgravata autem est manus Domini super Azotios et demolitus est eos et percussit in secretiori parte natium Azotum et fines eius
1SAM|5|7|videntes autem viri azotii huiuscemodi plagam dixerunt non maneat arca Dei Israhel apud nos quoniam dura est manus eius super nos et super Dagon deum nostrum
1SAM|5|8|et mittentes congregaverunt omnes satrapas Philisthinorum ad se et dixerunt quid faciemus de arca Dei Israhel responderuntque Getthei circumducatur arca Dei Israhel et circumduxerunt arcam Dei Israhel
1SAM|5|9|illis autem circumducentibus eam fiebat manus Dei per singulas civitates interfectionis magnae nimis et percutiebat viros uniuscuiusque urbis a parvo usque ad maiorem et conputrescebant prominentes extales eorum
1SAM|5|10|miserunt ergo arcam Dei in Accaron cumque venisset arca Dei in Accaron exclamaverunt Accaronitae dicentes adduxerunt ad nos arcam Dei Israhel ut interficiat nos et populum nostrum
1SAM|5|11|miserunt itaque et congregaverunt omnes satrapas Philisthinorum qui dixerunt dimittite arcam Dei Israhel et revertatur in locum suum et non interficiat nos cum populo nostro
1SAM|5|12|fiebat enim pavor mortis in singulis urbibus et gravissima valde manus Dei viri quoque qui mortui non fuerant percutiebantur in secretiori parte natium et ascendebat ululatus uniuscuiusque civitatis in caelum
1SAM|6|1|fuit ergo arca Domini in regione Philisthinorum septem mensibus
1SAM|6|2|et vocaverunt Philisthim sacerdotes et divinos dicentes quid faciemus de arca Dei indicate nobis quomodo remittemus eam in locum suum qui dixerunt
1SAM|6|3|si remittitis arcam Dei Israhel nolite dimittere eam vacuam sed quod debetis reddite ei pro peccato et tunc curabimini et scietis quare non recedat manus eius a vobis
1SAM|6|4|qui dixerunt quid est quod pro delicto reddere debeamus ei responderuntque illi
1SAM|6|5|iuxta numerum provinciarum Philisthim quinque anos aureos facietis et quinque mures aureos quia plaga una fuit omnibus vobis et satrapis vestris facietisque similitudines anorum vestrorum et similitudines murium qui demoliti sunt terram et dabitis Deo Israhel gloriam si forte relevet manum suam a vobis et a diis vestris et a terra vestra
1SAM|6|6|quare gravatis corda vestra sicut adgravavit Aegyptus et Pharao cor suum nonne postquam percussus est tunc dimisit eos et abierunt
1SAM|6|7|nunc ergo arripite et facite plaustrum novum unum et duas vaccas fetas quibus non est inpositum iugum iungite in plaustro et recludite vitulos earum domi
1SAM|6|8|tolletisque arcam Domini et ponetis in plaustro et vasa aurea quae exsolvistis ei pro delicto ponetis in capsella ad latus eius et dimittite eam ut vadat
1SAM|6|9|et aspicietis et si quidem per viam finium suorum ascenderit contra Bethsames ipse fecit nobis malum hoc grande sin autem minime sciemus quia nequaquam manus eius tetigit nos sed casu accidit
1SAM|6|10|fecerunt ergo illi hoc modo et tollentes duas vaccas quae lactabant vitulos iunxerunt ad plaustrum vitulosque earum concluserunt domi
1SAM|6|11|et posuerunt arcam Dei super plaustrum et capsellam quae habebat mures aureos et similitudinem anorum
1SAM|6|12|ibant autem in directum vaccae per viam quae ducit Bethsames et itinere uno gradiebantur pergentes et mugientes et non declinabant neque ad dextram neque ad sinistram sed et satrapae Philisthinorum sequebantur usque ad terminos Bethsames
1SAM|6|13|porro Bethsamitae metebant triticum in valle et elevantes oculos viderunt arcam et gavisi sunt cum vidissent
1SAM|6|14|et plaustrum venit in agrum Iosue Bethsamitae et stetit ibi erat autem ibi lapis magnus et conciderunt ligna plaustri vaccasque inposuerunt super ea holocaustum Domino
1SAM|6|15|Levitae autem deposuerunt arcam Dei et capsellam quae erat iuxta eam in qua erant vasa aurea et posuerunt super lapidem grandem viri autem bethsamitae obtulerunt holocausta et immolaverunt victimas in die illa Domino
1SAM|6|16|et quinque satrapae Philisthinorum viderunt et reversi sunt in Accaron in die illa
1SAM|6|17|hii sunt autem ani aurei quos reddiderunt Philisthim pro delicto Domino Azotus unum Gaza unum Ascalon unum Geth unum Accaron unum
1SAM|6|18|et mures aureos secundum numerum urbium Philisthim quinque provinciarum ab urbe murata usque ad villam quae erat absque muro et usque ad Abel magnum super quem posuerunt arcam Domini quae erat usque in illa die in agro Iosue Bethsamitis
1SAM|6|19|percussit autem de viris bethsamitibus eo quod vidissent arcam Domini et percussit de populo septuaginta viros et quinquaginta milia plebis luxitque populus quod percussisset Dominus plebem plaga magna
1SAM|6|20|et dixerunt viri bethsamitae quis poterit stare in conspectu Domini Dei sancti huius et ad quem ascendet a nobis
1SAM|6|21|miseruntque nuntios ad habitatores Cariathiarim dicentes reduxerunt Philisthim arcam Domini descendite et ducite eam ad vos
1SAM|7|1|venerunt ergo viri Cariathiarim et duxerunt arcam Domini et intulerunt eam in domum Abinadab in Gabaa Eleazarum autem filium eius sanctificaverunt ut custodiret arcam Domini
1SAM|7|2|et factum est ex qua die mansit arca in Cariathiarim multiplicati sunt dies erat quippe iam annus vicesimus et requievit omnis domus Israhel post Dominum
1SAM|7|3|ait autem Samuhel ad universam domum Israhel dicens si in toto corde vestro revertimini ad Dominum auferte deos alienos de medio vestrum et Astharoth et praeparate corda vestra Domino et servite ei soli et eruet vos de manu Philisthim
1SAM|7|4|abstulerunt ergo filii Israhel Baalim et Astharoth et servierunt Domino soli
1SAM|7|5|dixit autem Samuhel congregate universum Israhel in Masphat ut orem pro vobis Dominum
1SAM|7|6|et convenerunt in Masphat hauseruntque aquam et effuderunt in conspectu Domini et ieiunaverunt in die illa et dixerunt ibi peccavimus Domino iudicavitque Samuhel filios Israhel in Masphat
1SAM|7|7|et audierunt Philisthim quod congregati essent filii Israhel in Masphat et ascenderunt satrapae Philisthinorum ad Israhel quod cum audissent filii Israhel timuerunt a facie Philisthinorum
1SAM|7|8|dixeruntque ad Samuhel ne cesses pro nobis clamare ad Dominum Deum nostrum ut salvet nos de manu Philisthinorum
1SAM|7|9|tulit autem Samuhel agnum lactantem unum et obtulit illum holocaustum integrum Domino et clamavit Samuhel ad Dominum pro Israhel et exaudivit eum Dominus
1SAM|7|10|factum est ergo cum Samuhel offerret holocaustum Philistheos inire proelium contra Israhel intonuit autem Dominus fragore magno in die illa super Philisthim et exterruit eos et caesi sunt a filiis Israhel
1SAM|7|11|egressique viri Israhel de Masphat persecuti sunt Philistheos et percusserunt eos usque ad locum qui erat subter Bethchar
1SAM|7|12|tulit autem Samuhel lapidem unum et posuit eum inter Masphat et inter Sen et vocavit nomen eius lapis Adiutorii dixitque hucusque auxiliatus est nobis Dominus
1SAM|7|13|et humiliati sunt Philisthim nec adposuerunt ultra ut venirent in terminos Israhel facta est itaque manus Domini super Philistheos cunctis diebus Samuhel
1SAM|7|14|et redditae sunt urbes quas tulerant Philisthim ab Israhel Israheli ab Accaron usque Geth et terminos suos liberavit Israhel de manu Philisthinorum eratque pax inter Israhel et Amorreum
1SAM|7|15|iudicabat quoque Samuhel Israhel cunctis diebus vitae suae
1SAM|7|16|et ibat per singulos annos circumiens Bethel et Galgal et Masphat et iudicabat Israhelem in supradictis locis
1SAM|7|17|revertebaturque in Ramatha ibi enim erat domus eius et ibi iudicabat Israhelem aedificavit etiam ibi altare Domino
1SAM|8|1|factum est autem cum senuisset Samuhel posuit filios suos iudices Israhel
1SAM|8|2|fuitque nomen filii eius primogeniti Iohel et nomen secundi Abia iudicum in Bersabee
1SAM|8|3|et non ambulaverunt filii illius in viis eius sed declinaverunt post avaritiam acceperuntque munera et perverterunt iudicium
1SAM|8|4|congregati ergo universi maiores natu Israhel venerunt ad Samuhel in Ramatha
1SAM|8|5|dixeruntque ei ecce tu senuisti et filii tui non ambulant in viis tuis constitue nobis regem ut iudicet nos sicut universae habent nationes
1SAM|8|6|displicuitque sermo in oculis Samuhelis eo quod dixissent da nobis regem ut iudicet nos et oravit Samuhel Dominum
1SAM|8|7|dixit autem Dominus ad Samuhel audi vocem populi in omnibus quae loquuntur tibi non enim te abiecerunt sed me ne regnem super eos
1SAM|8|8|iuxta omnia opera sua quae fecerunt a die qua eduxi eos de Aegypto usque ad diem hanc sicut dereliquerunt me et servierunt diis alienis sic faciunt etiam tibi
1SAM|8|9|nunc ergo audi vocem eorum verumtamen contestare eos et praedic eis ius regis qui regnaturus est super eos
1SAM|8|10|dixit itaque Samuhel omnia verba Domini ad populum qui petierat a se regem
1SAM|8|11|et ait hoc erit ius regis qui imperaturus est vobis filios vestros tollet et ponet in curribus suis facietque sibi equites et praecursores quadrigarum suarum
1SAM|8|12|et constituet sibi tribunos et centuriones et aratores agrorum suorum et messores segetum et fabros armorum et curruum suorum
1SAM|8|13|filias quoque vestras faciet sibi unguentarias et focarias et panificas
1SAM|8|14|agros quoque vestros et vineas et oliveta optima tollet et dabit servis suis
1SAM|8|15|sed et segetes vestras et vinearum reditus addecimabit ut det eunuchis et famulis suis
1SAM|8|16|servos etiam vestros et ancillas et iuvenes optimos et asinos auferet et ponet in opere suo
1SAM|8|17|greges vestros addecimabit vosque eritis ei servi
1SAM|8|18|et clamabitis in die illa a facie regis vestri quem elegistis vobis et non exaudiet vos Dominus in die illa
1SAM|8|19|noluit autem populus audire vocem Samuhel sed dixerunt nequaquam rex enim erit super nos
1SAM|8|20|et erimus nos quoque sicut omnes gentes et iudicabit nos rex noster et egredietur ante nos et pugnabit bella nostra pro nobis
1SAM|8|21|et audivit Samuhel omnia verba populi et locutus est ea in auribus Domini
1SAM|8|22|dixit autem Dominus ad Samuhel audi vocem eorum et constitue super eos regem et ait Samuhel ad viros Israhel vadat unusquisque in civitatem suam
1SAM|9|1|et erat vir de Beniamin nomine Cis filius Abihel filii Seror filii Bechoreth filii Afia filii viri Iemini fortis robore
1SAM|9|2|et erat ei filius vocabulo Saul electus et bonus et non erat vir de filiis Israhel melior illo ab umero et sursum eminebat super omnem populum
1SAM|9|3|perierant autem asinae Cis patris Saul et dixit Cis ad Saul filium suum tolle tecum unum de pueris et consurgens vade et quaere asinas qui cum transissent per montem Ephraim
1SAM|9|4|et per terram Salisa et non invenissent transierunt etiam per terram Salim et non erant sed et per terram Iemini et minime reppererunt
1SAM|9|5|cum autem venissent in terram Suph dixit Saul ad puerum suum qui erat cum eo veni et revertamur ne forte dimiserit pater meus asinas et sollicitus sit pro nobis
1SAM|9|6|qui ait ei ecce est vir Dei in civitate hac vir nobilis omne quod loquitur absque ambiguitate venit nunc ergo eamus illuc si forte indicet nobis de via nostra propter quam venimus
1SAM|9|7|dixitque Saul ad puerum suum ecce ibimus quid feremus ad virum panis defecit in sitarciis nostris et sportulam non habemus ut demus homini Dei nec quicquam aliud
1SAM|9|8|rursum puer respondit Sauli et ait ecce inventa est in manu mea quarta pars stateris argenti demus homini Dei ut indicet nobis viam nostram
1SAM|9|9|olim in Israhel sic loquebatur unusquisque vadens consulere Deum venite et eamus ad videntem qui enim propheta dicitur hodie vocabatur olim videns
1SAM|9|10|et dixit Saul ad puerum suum optimus sermo tuus veni eamus et ierunt in civitatem in qua erat vir Dei
1SAM|9|11|cumque ascenderent clivum civitatis invenerunt puellas egredientes ad hauriendam aquam et dixerunt eis num hic est videns
1SAM|9|12|quae respondentes dixerunt illis hic est ecce ante te festina nunc hodie enim venit in civitate quia sacrificium est hodie populo in excelso
1SAM|9|13|ingredientes urbem statim invenietis eum antequam ascendat excelsum ad vescendum neque enim comesurus est populus donec ille veniat quia ipse benedicit hostiae et deinceps comedunt qui vocati sunt nunc ergo conscendite quia hodie repperietis eum
1SAM|9|14|et ascenderunt in civitatem cumque illi ambularent in medio urbis apparuit Samuhel egrediens obviam eis ut ascenderet in excelsum
1SAM|9|15|Dominus autem revelaverat auriculam Samuhel ante unam diem quam veniret Saul dicens
1SAM|9|16|hac ipsa quae nunc est hora cras mittam ad te virum de terra Beniamin et ungues eum ducem super populum meum Israhel et salvabit populum meum de manu Philisthinorum quia respexi populum meum venit enim clamor eorum ad me
1SAM|9|17|cumque aspexisset Samuhel Saulem Dominus ait ei ecce vir quem dixeram tibi iste dominabitur populo meo
1SAM|9|18|accessit autem Saul ad Samuhelem in medio portae et ait indica oro mihi ubi est domus videntis
1SAM|9|19|et respondit Samuhel Sauli dicens ego sum videns ascende ante me in excelsum ut comedatis mecum hodie et dimittam te mane et omnia quae sunt in corde tuo indicabo tibi
1SAM|9|20|et de asinis quas perdidisti nudius tertius ne sollicitus sis quia inventae sunt et cuius erunt optima quaeque Israhel nonne tibi et omni domui patris tui
1SAM|9|21|respondens autem Saul ait numquid non filius Iemini ego sum de minima tribu Israhel et cognatio mea novissima inter omnes familias de tribu Beniamin quare ergo locutus es mihi sermonem istum
1SAM|9|22|adsumens itaque Samuhel Saulem et puerum eius introduxit eos in triclinium et dedit eis locum in capite eorum qui fuerant invitati erant enim quasi triginta viri
1SAM|9|23|dixitque Samuhel coco da partem quam dedi tibi et praecepi ut reponeres seorsum apud te
1SAM|9|24|levavit autem cocus armum et posuit ante Saul dixitque Samuhel ecce quod remansit pone ante te et comede quia de industria servatum est tibi quando populum vocavi et comedit Saul cum Samuhel in die illa
1SAM|9|25|et descenderunt de excelso in oppidum et locutus est cum Saul in solario
1SAM|9|26|cumque mane surrexissent et iam dilucesceret vocavit Samuhel Saul in solarium dicens surge ut dimittam te et surrexit Saul egressique sunt ambo ipse videlicet et Samuhel
1SAM|9|27|cumque descenderent in extrema parte civitatis Samuhel dixit ad Saul dic puero ut antecedat nos et transeat tu autem subsiste paulisper ut indicem tibi verbum Domini
1SAM|10|1|tulit autem Samuhel lenticulam olei et effudit super caput eius et deosculatus eum ait ecce unxit te Dominus super hereditatem suam in principem
1SAM|10|2|cum abieris hodie a me invenies duos viros iuxta sepulchrum Rachel in finibus Beniamin in meridie dicentque tibi inventae sunt asinae ad quas ieras perquirendas et intermissis pater tuus asinis sollicitus est pro vobis et dicit quid faciam de filio meo
1SAM|10|3|cumque abieris inde et ultra transieris et veneris ad quercum Thabor invenient te ibi tres viri ascendentes ad Deum in Bethel unus portans tres hedos et alius tres tortas panis et alius portans lagoenam vini
1SAM|10|4|cumque te salutaverint dabunt tibi duos panes et accipies de manu eorum
1SAM|10|5|post haec venies in collem Domini ubi est statio Philisthinorum et cum ingressus fueris ibi urbem obviam habebis gregem prophetarum descendentium de excelso et ante eos psalterium et tympanum et tibiam et citharam ipsosque prophetantes
1SAM|10|6|et insiliet in te spiritus Domini et prophetabis cum eis et mutaberis in virum alium
1SAM|10|7|quando ergo evenerint signa haec omnia tibi fac quaecumque invenerit manus tua quia Dominus tecum est
1SAM|10|8|et descendes ante me in Galgala ego quippe descendam ad te ut offeras oblationem et immoles victimas pacificas septem diebus expectabis donec veniam ad te et ostendam tibi quae facias
1SAM|10|9|itaque cum avertisset umerum suum ut abiret a Samuhele inmutavit ei Deus cor aliud et venerunt omnia signa haec in die illa
1SAM|10|10|veneruntque ad praedictum collem et ecce cuneus prophetarum obvius ei et insilivit super eum spiritus Dei et prophetavit in medio eorum
1SAM|10|11|videntes autem omnes qui noverant eum heri et nudius tertius quod esset cum prophetis et prophetaret dixerunt ad invicem quaenam res accidit filio Cis num et Saul in prophetis
1SAM|10|12|responditque alius ad alterum dicens et quis pater eorum propterea versum est in proverbium num et Saul inter prophetas
1SAM|10|13|cessavit autem prophetare et venit ad excelsum
1SAM|10|14|dixitque patruus Saul ad eum et ad puerum eius quo abistis qui responderunt quaerere asinas quas cum non repperissemus venimus ad Samuhelem
1SAM|10|15|et dixit ei patruus suus indica mihi quid dixerit tibi Samuhel
1SAM|10|16|et ait Saul ad patruum suum indicavit nobis quia inventae essent asinae de sermone autem regni non indicavit ei quem locutus illi fuerat Samuhel
1SAM|10|17|et convocavit Samuhel populum ad Dominum in Maspha
1SAM|10|18|et ait ad filios Israhel haec dicit Dominus Deus Israhel ego eduxi Israhel de Aegypto et erui vos de manu Aegyptiorum et de manu omnium regum qui adfligebant vos
1SAM|10|19|vos autem hodie proiecistis Deum vestrum qui solus salvavit vos de universis malis et tribulationibus vestris et dixistis nequaquam sed regem constitue super nos nunc ergo state coram Domino per tribus vestras et per familias
1SAM|10|20|et adplicuit Samuhel omnes tribus Israhel et cecidit sors tribus Beniamin
1SAM|10|21|et adplicuit tribum Beniamin et cognationes eius et cecidit cognatio Metri et pervenit usque ad Saul filium Cis quaesierunt ergo eum et non est inventus
1SAM|10|22|et consuluerunt post haec Dominum utrumnam venturus esset illuc responditque Dominus ecce absconditus est domi
1SAM|10|23|cucurrerunt itaque et tulerunt eum inde stetitque in medio populi et altior fuit universo populo ab umero et sursum
1SAM|10|24|et ait Samuhel ad omnem populum certe videtis quem elegit Dominus quoniam non sit similis ei in omni populo et clamavit cunctus populus et ait vivat rex
1SAM|10|25|locutus est autem Samuhel ad populum legem regni et scripsit in libro et reposuit coram Domino et dimisit Samuhel omnem populum singulos in domum suam
1SAM|10|26|sed et Saul abiit in domum suam in Gabaath et abiit cum eo pars exercitus quorum tetigerat Deus corda
1SAM|10|27|filii vero Belial dixerunt num salvare nos poterit iste et despexerunt eum et non adtulerunt ei munera ille vero dissimulabat se audire
1SAM|11|1|ascendit autem Naas Ammonites et pugnare coepit adversus Iabesgalaad dixeruntque omnes viri Iabes ad Naas habeto nos foederatos et serviemus tibi
1SAM|11|2|et respondit ad eos Naas Ammonites in hoc feriam vobiscum foedus ut eruam omnium vestrum oculos dextros ponamque vos obprobrium in universo Israhel
1SAM|11|3|et dixerunt ad eum seniores Iabes concede nobis septem dies ut mittamus nuntios in universos terminos Israhel et si non fuerit qui defendat nos egrediemur ad te
1SAM|11|4|venerunt ergo nuntii in Gabaath Saulis et locuti sunt verba audiente populo et levavit omnis populus vocem suam et flevit
1SAM|11|5|et ecce Saul veniebat sequens boves de agro et ait quid habet populus quod plorat et narraverunt ei verba virorum Iabes
1SAM|11|6|et insilivit spiritus Domini in Saul cum audisset verba haec et iratus est furor eius nimis
1SAM|11|7|et adsumens utrumque bovem concidit in frusta misitque in omnes terminos Israhel per manum nuntiorum dicens quicumque non exierit secutusque fuerit Saul et Samuhelem sic fiet bubus eius invasit ergo timor Domini populum et egressi sunt quasi vir unus
1SAM|11|8|et recensuit eos in Bezec fueruntque filiorum Israhel trecenta milia virorum autem Iuda triginta milia
1SAM|11|9|et dixerunt nuntiis qui venerant sic dicetis viris qui sunt in Iabesgalaad cras erit vobis salus cum incaluerit sol venerunt ergo nuntii et adnuntiaverunt viris Iabes qui laetati sunt
1SAM|11|10|et dixerunt mane exibimus ad vos et facietis nobis omne quod placuerit vobis
1SAM|11|11|et factum est cum venisset dies crastinus constituit Saul populum in tres partes et ingressus est media castra in vigilia matutina et percussit Ammon usque dum incalesceret dies reliqui autem dispersi sunt ita ut non relinquerentur in eis duo pariter
1SAM|11|12|et ait populus ad Samuhel quis est iste qui dixit Saul non regnabit super nos date viros et interficiemus eos
1SAM|11|13|et ait Saul non occidetur quisquam in die hac quia hodie fecit Dominus salutem in Israhel
1SAM|11|14|dixit autem Samuhel ad populum venite et eamus in Galgala et innovemus ibi regnum
1SAM|11|15|et perrexit omnis populus in Galgala et fecerunt ibi regem Saul coram Domino in Galgala et immolaverunt ibi victimas pacificas coram Domino et laetatus est ibi Saul et cuncti viri Israhel nimis
1SAM|12|1|dixit autem Samuhel ad universum Israhel ecce audivi vocem vestram iuxta omnia quae locuti estis ad me et constitui super vos regem
1SAM|12|2|et nunc rex graditur ante vos ego autem senui et incanui porro filii mei vobiscum sunt itaque conversatus coram vobis ab adulescentia mea usque ad diem hanc ecce praesto sum
1SAM|12|3|loquimini de me coram Domino et coram christo eius utrum bovem cuiusquam tulerim an asinum si quempiam calumniatus sum si oppressi aliquem si de manu cuiusquam munus accepi et contemnam illud hodie restituamque vobis
1SAM|12|4|et dixerunt non es calumniatus nos neque oppressisti neque tulisti de manu alicuius quippiam
1SAM|12|5|dixitque ad eos testis Dominus adversus vos et testis christus eius in die hac quia non inveneritis in manu mea quippiam et dixerunt testis
1SAM|12|6|et ait Samuhel ad populum Dominus qui fecit Mosen et Aaron et eduxit patres nostros de terra Aegypti
1SAM|12|7|nunc ergo state ut iudicio contendam adversum vos coram Domino de omnibus misericordiis Domini quas fecit vobiscum et cum patribus vestris
1SAM|12|8|quomodo ingressus est Iacob in Aegyptum et clamaverunt patres vestri ad Dominum et misit Dominus Mosen et Aaron et eduxit patres vestros ex Aegypto et conlocavit eos in loco hoc
1SAM|12|9|qui obliti sunt Domini Dei sui et tradidit eos in manu Sisarae magistri militiae Asor et in manu Philisthinorum et in manu regis Moab et pugnaverunt adversum eos
1SAM|12|10|postea autem clamaverunt ad Dominum et dixerunt peccavimus quia dereliquimus Dominum et servivimus Baalim et Astharoth nunc ergo erue nos de manu inimicorum nostrorum et serviemus tibi
1SAM|12|11|et misit Dominus Hierobaal et Bedan et Ieptha et Samuhel et eruit vos de manu inimicorum vestrorum per circuitum et habitastis confidenter
1SAM|12|12|videntes autem quod Naas rex filiorum Ammon venisset adversum vos dixistis mihi nequaquam sed rex imperabit nobis cum Dominus Deus vester regnaret in vobis
1SAM|12|13|nunc ergo praesto est rex vester quem elegistis et petistis ecce dedit vobis Dominus regem
1SAM|12|14|si timueritis Dominum et servieritis ei et audieritis vocem eius et non exasperaveritis os Domini eritis et vos et rex qui imperat vobis sequentes Dominum Deum vestrum
1SAM|12|15|si autem non audieritis vocem Domini sed exasperaveritis sermonem Domini erit manus Domini super vos et super patres vestros
1SAM|12|16|sed et nunc state et videte rem istam grandem quam facturus est Dominus in conspectu vestro
1SAM|12|17|numquid non messis tritici est hodie invocabo Dominum et dabit voces et pluvias et scietis et videbitis quia grande malum feceritis vobis in conspectu Domini petentes super vos regem
1SAM|12|18|et clamavit Samuhel ad Dominum et dedit Dominus voces et pluviam in die illa
1SAM|12|19|et timuit omnis populus nimis Dominum et Samuhelem dixitque universus populus ad Samuhel ora pro servis tuis ad Dominum Deum tuum ut non moriamur addidimus enim universis peccatis nostris malum ut peteremus nobis regem
1SAM|12|20|dixit autem Samuhel ad populum nolite timere vos fecistis universum malum hoc verumtamen nolite recedere a tergo Domini et servite Domino in omni corde vestro
1SAM|12|21|et nolite declinare post vana quae non proderunt vobis neque eruent vos quia vana sunt
1SAM|12|22|et non derelinquet Dominus populum suum propter nomen suum magnum quia iuravit Dominus facere vos sibi populum
1SAM|12|23|absit autem a me hoc peccatum in Domino ut cessem orare pro vobis et docebo vos viam bonam et rectam
1SAM|12|24|igitur timete Dominum et servite ei in veritate et ex toto corde vestro vidistis enim magnifica quae in vobis gesserit
1SAM|12|25|quod si perseveraveritis in malitia et vos et rex vester pariter peribitis
1SAM|13|1|filius unius anni Saul cum regnare coepisset duobus autem annis regnavit super Israhel
1SAM|13|2|et elegit sibi Saul tria milia de Israhel et erant cum Saul duo milia in Machmas et in monte Bethel mille autem cum Ionathan in Gabaath Beniamin porro ceterum populum remisit unumquemque in tabernacula sua
1SAM|13|3|et percussit Ionathan stationem Philisthim quae erat in Gabaa quod cum audissent Philisthim Saul cecinit bucina in omni terra dicens audiant Hebraei
1SAM|13|4|et universus Israhel audivit huiuscemodi famam percussit Saul stationem Philisthinorum et erexit se Israhel adversum Philisthim clamavit ergo populus post Saul in Galgala
1SAM|13|5|et Philisthim congregati sunt ad proeliandum contra Israhel triginta milia curruum et sex milia equitum et reliquum vulgus sicut harena quae est in litore maris plurima et ascendentes castrametati sunt in Machmas ad orientem Bethaven
1SAM|13|6|quod cum vidissent viri Israhel se in arto sitos adflictus est enim populus absconderunt se in speluncis et in abditis in petris quoque et in antris et in cisternis
1SAM|13|7|Hebraei autem transierunt Iordanem terram Gad et Galaad cumque adhuc esset Saul in Galgal universus populus perterritus est qui sequebatur eum
1SAM|13|8|et expectavit septem diebus iuxta placitum Samuhel et non venit Samuhel in Galgala dilapsusque est populus ab eo
1SAM|13|9|ait ergo Saul adferte mihi holocaustum et pacifica et obtulit holocaustum
1SAM|13|10|cumque conplesset offerens holocaustum ecce Samuhel veniebat et egressus est Saul obviam ei ut salutaret eum
1SAM|13|11|locutusque est ad eum Samuhel quid fecisti respondit Saul quia vidi quod dilaberetur populus a me et tu non veneras iuxta placitos dies porro Philisthim congregati fuerant in Machmas
1SAM|13|12|dixi nunc descendent Philisthim ad me in Galgala et faciem Domini non placavi necessitate conpulsus obtuli holocaustum
1SAM|13|13|dixitque Samuhel ad Saul stulte egisti nec custodisti mandata Domini Dei tui quae praecepit tibi quod si non fecisses iam nunc praeparasset Dominus regnum tuum super Israhel in sempiternum
1SAM|13|14|sed nequaquam regnum tuum ultra consurget quaesivit sibi Dominus virum iuxta cor suum et praecepit ei Dominus ut esset dux super populum suum eo quod non servaveris quae praecepit Dominus
1SAM|13|15|surrexit autem Samuhel et ascendit de Galgalis in Gabaa Beniamin et recensuit Saul populum qui inventi fuerant cum eo quasi sescentos viros
1SAM|13|16|et Saul et Ionathan filius eius populusque qui inventus fuerat cum eis erat in Gabaa Beniamin porro Philisthim consederant in Machmas
1SAM|13|17|et egressi sunt ad praedandum de castris Philisthim tres cunei unus cuneus pergebat contra viam Ephra ad terram Saul
1SAM|13|18|porro alius ingrediebatur per viam Bethoron tertius autem verterat se ad iter termini inminentis valli Seboim contra desertum
1SAM|13|19|porro faber ferrarius non inveniebatur in omni terra Israhel caverant enim Philisthim ne forte facerent Hebraei gladium aut lanceam
1SAM|13|20|descendebat ergo omnis Israhel ad Philisthim ut exacueret unusquisque vomerem suum et ligonem et securim et sarculum
1SAM|13|21|retunsae itaque erant acies vomerum et ligonum et tridentum et securium usque ad stimulum corrigendum
1SAM|13|22|cumque venisset dies proelii non est inventus ensis et lancea in manu totius populi qui erat cum Saul et cum Ionathan excepto Saul et Ionathan filio eius
1SAM|13|23|egressa est autem statio Philisthim ut transcenderet in Machmas
1SAM|14|1|et accidit quadam die ut diceret Ionathan filius Saul ad adulescentem armigerum suum veni et transeamus ad stationem Philisthim quae est trans locum illum patri autem suo hoc ipsum non indicavit
1SAM|14|2|porro Saul morabatur in extrema parte Gabaa sub malogranato quae erat in Magron et erat populus cum eo quasi sescentorum virorum
1SAM|14|3|et Ahias filius Achitob fratris Ichabod filii Finees qui ortus fuerat ex Heli sacerdote Domini in Silo portabat ephod sed et populus ignorabat quod isset Ionathan
1SAM|14|4|erant autem inter ascensus per quos nitebatur Ionathan transire ad stationem Philisthinorum eminentes petrae ex utraque parte et quasi in modum dentium scopuli hinc inde praerupti nomen uni Boses et nomen alteri Sene
1SAM|14|5|unus scopulus prominens ad aquilonem ex adverso Machmas et alter a meridie contra Gabaa
1SAM|14|6|dixit autem Ionathan ad adulescentem armigerum suum veni transeamus ad stationem incircumcisorum horum si forte faciat Dominus pro nobis quia non est Domino difficile salvare vel in multitudine vel in paucis
1SAM|14|7|dixitque ei armiger suus fac omnia quae placent animo tuo perge quo cupis ero tecum ubicumque volueris
1SAM|14|8|et ait Ionathan ecce nos transimus ad viros istos cumque apparuerimus eis
1SAM|14|9|si taliter locuti fuerint ad nos manete donec veniamus ad vos stemus in loco nostro nec ascendamus ad eos
1SAM|14|10|si autem dixerint ascendite ad nos ascendamus quia tradidit eos Dominus in manibus nostris hoc erit nobis signum
1SAM|14|11|apparuit igitur uterque stationi Philisthinorum dixeruntque Philisthim en Hebraei egrediuntur de cavernis in quibus absconditi fuerant
1SAM|14|12|et locuti sunt viri de statione ad Ionathan et ad armigerum eius dixeruntque ascendite ad nos et ostendimus vobis rem et ait Ionathan ad armigerum suum ascendamus sequere me tradidit enim eos Dominus in manu Israhel
1SAM|14|13|ascendit autem Ionathan reptans manibus et pedibus et armiger eius post eum itaque alii cadebant ante Ionathan alios armiger eius interficiebat sequens eum
1SAM|14|14|et facta est plaga prima quam percussit Ionathan et armiger eius quasi viginti virorum in media parte iugeri quam par boum in die arare consuevit
1SAM|14|15|et factum est miraculum in castris per agros sed et omnis populus stationis eorum qui ierant ad praedandum obstipuit et conturbata est terra et accidit quasi miraculum a Deo
1SAM|14|16|et respexerunt speculatores Saul qui erant in Gabaa Beniamin et ecce multitudo prostrata et huc illucque diffugiens
1SAM|14|17|et ait Saul populo qui erat cum eo requirite et videte quis abierit ex nobis cumque requisissent reppertum est non adesse Ionathan et armigerum eius
1SAM|14|18|et ait Saul ad Ahiam adplica arcam Dei erat enim ibi arca Dei in die illa cum filiis Israhel
1SAM|14|19|cumque loqueretur Saul ad sacerdotem tumultus magnus exortus est in castris Philisthinorum crescebatque paulatim et clarius reboabat et ait Saul ad sacerdotem contrahe manum tuam
1SAM|14|20|conclamavit ergo Saul et omnis populus qui erat cum eo et venerunt usque ad locum certaminis et ecce versus fuerat gladius uniuscuiusque ad proximum suum et caedes magna nimis
1SAM|14|21|sed et Hebraei qui fuerant cum Philisthim heri et nudius tertius ascenderantque cum eis in castris reversi sunt ut essent cum Israhele qui erant cum Saul et Ionathan
1SAM|14|22|omnes quoque Israhelitae qui se absconderant in monte Ephraim audientes quod fugissent Philisthim sociaverunt se cum suis in proelio
1SAM|14|23|et salvavit Dominus in die illa Israhel pugna autem pervenit usque Bethaven
1SAM|14|24|et vir Israhel sociatus sibi est in die illa adiuravit autem Saul populum dicens maledictus vir qui comederit panem usque ad vesperam donec ulciscar de inimicis meis et non manducavit universus populus panem
1SAM|14|25|omneque terrae vulgus venit in saltum in quo erat mel super faciem agri
1SAM|14|26|ingressus est itaque populus saltum et apparuit fluens mel nullusque adplicuit manum ad os suum timebat enim populus iuramentum
1SAM|14|27|porro Ionathan non audierat cum adiuraret pater eius populum extenditque summitatem virgae quam habebat in manu et intinxit in favo mellis et convertit manum suam ad os suum et inluminati sunt oculi eius
1SAM|14|28|respondensque unus de populo ait iureiurando constrinxit pater tuus populum dicens maledictus qui comederit panem hodie defecerat autem populus
1SAM|14|29|dixitque Ionathan turbavit pater meus terram vidistis ipsi quia inluminati sunt oculi mei eo quod gustaverim paululum de melle isto
1SAM|14|30|quanto magis si comedisset populus de praeda inimicorum suorum quam repperit nonne maior facta fuisset plaga in Philisthim
1SAM|14|31|percusserunt ergo in die illa Philistheos a Machmis usque in Ahialon defatigatus est autem populus nimis
1SAM|14|32|et versus ad praedam tulit oves et boves et vitulos et mactaverunt in terra comeditque populus cum sanguine
1SAM|14|33|nuntiaverunt autem Saul dicentes quod populus peccasset Domino comedens cum sanguine qui ait praevaricati estis volvite ad me iam nunc saxum grande
1SAM|14|34|et dixit Saul dispergimini in vulgus et dicite eis ut adducat ad me unusquisque bovem suum et arietem et occidite super istud et vescimini et non peccabitis Domino comedentes cum sanguine adduxit itaque omnis populus unusquisque bovem in manu sua usque ad noctem et occiderunt ibi
1SAM|14|35|aedificavit autem Saul altare Domini tuncque primum coepit aedificare altare Domini
1SAM|14|36|et dixit Saul inruamus super Philisthim nocte et vastemus eos usque dum inlucescat mane nec relinquamus de eis virum dixitque populus omne quod bonum videtur in oculis tuis fac et ait sacerdos accedamus huc ad Deum
1SAM|14|37|et consuluit Saul Deum num persequar Philisthim si trades eos in manu Israhel et non respondit ei in die illa
1SAM|14|38|dixitque Saul adplicate huc universos angulos populi et scitote et videte per quem acciderit peccatum hoc hodie
1SAM|14|39|vivit Dominus salvator Israhel quia si per Ionathan filium meum factum est absque retractatione morietur ad quod nullus contradixit ei de omni populo
1SAM|14|40|et ait ad universum Israhel separamini vos in partem unam et ego cum Ionathan filio meo ero in parte una respondit populus ad Saul quod bonum videtur in oculis tuis fac
1SAM|14|41|et dixit Saul ad Dominum Deum Israhel da indicium et deprehensus est Ionathan et Saul populus autem exivit
1SAM|14|42|et ait Saul mittite sortem inter me et inter Ionathan filium meum et captus est Ionathan
1SAM|14|43|dixit autem Saul ad Ionathan indica mihi quid feceris et indicavit ei Ionathan et ait gustans gustavi in summitate virgae quae erat in manu mea paululum mellis et ecce ego morior
1SAM|14|44|et ait Saul haec faciat mihi Deus et haec addat quia morte morieris Ionathan
1SAM|14|45|dixitque populus ad Saul ergone Ionathan morietur qui fecit salutem hanc magnam in Israhel hoc nefas est vivit Dominus si ceciderit capillus de capite eius in terram quia cum Deo operatus est hodie liberavit ergo populus Ionathan ut non moreretur
1SAM|14|46|recessitque Saul nec persecutus est Philisthim porro Philisthim abierunt in loca sua
1SAM|14|47|at Saul confirmato regno super Israhel pugnabat per circuitum adversum omnes inimicos eius contra Moab et filios Ammon et Edom et reges Suba et Philistheos et quocumque se verterat superabat
1SAM|14|48|congregatoque exercitu percussit Amalech et eruit Israhel de manu vastatorum eius
1SAM|14|49|fuerunt autem filii Saul Ionathan et Iesui et Melchisua nomina duarum filiarum eius nomen primogenitae Merob et nomen minoris Michol
1SAM|14|50|et nomen uxoris Saul Ahinoem filia Ahimaas et nomina principum militiae eius Abner filius Ner patruelis Saul
1SAM|14|51|Cis fuerat pater Saul et Ner pater Abner filius Abihel
1SAM|14|52|erat autem bellum potens adversum Philistheos omnibus diebus Saul nam quemcumque viderat Saul virum fortem et aptum ad proelium sociabat eum sibi
1SAM|15|1|et dixit Samuhel ad Saul me misit Dominus ut unguerem te in regem super populum eius Israhel nunc ergo audi vocem Domini
1SAM|15|2|haec dicit Dominus exercituum recensui quaecumque fecit Amalech Israheli quomodo restitit ei in via cum ascenderet de Aegypto
1SAM|15|3|nunc igitur vade et percute Amalech et demolire universa eius non parcas ei sed interfice a viro usque ad mulierem et parvulum atque lactantem bovem et ovem camelum et asinum
1SAM|15|4|praecepit itaque Saul populo et recensuit eos quasi agnos ducenta milia peditum et decem milia virorum Iuda
1SAM|15|5|cumque venisset Saul usque ad civitatem Amalech tetendit insidias in torrente
1SAM|15|6|dixitque Saul Cineo abite recedite atque descendite ab Amalech ne forte involvam te cum eo tu enim fecisti misericordiam cum omnibus filiis Israhel cum ascenderent de Aegypto et recessit Cineus de medio Amalech
1SAM|15|7|percussitque Saul Amalech ab Evila donec venias Sur quae est e regione Aegypti
1SAM|15|8|et adprehendit Agag regem Amalech vivum omne autem vulgus interfecit in ore gladii
1SAM|15|9|et pepercit Saul et populus Agag et optimis gregibus ovium et armentorum et vestibus et arietibus et universis quae pulchra erant nec voluerunt disperdere ea quicquid vero vile fuit et reprobum hoc demoliti sunt
1SAM|15|10|factum est autem verbum Domini ad Samuhel dicens
1SAM|15|11|paenitet me quod constituerim Saul regem quia dereliquit me et verba mea opere non implevit contristatusque est Samuhel et clamavit ad Dominum tota nocte
1SAM|15|12|cumque de nocte surrexisset Samuhel ut iret ad Saul mane nuntiatum est Samuheli eo quod venisset Saul in Carmelum et erexisset sibi fornicem triumphalem et reversus transisset descendissetque in Galgala venit ergo Samuhel ad Saul et
1SAM|15|13|dixit ei Saul benedictus tu Domino implevi verbum Domini
1SAM|15|14|dixitque Samuhel et quae est haec vox gregum quae resonat in auribus meis et armentorum quam ego audio
1SAM|15|15|et ait Saul de Amalech adduxerunt ea pepercit enim populus melioribus ovibus et armentis ut immolarentur Domino Deo tuo reliqua vero occidimus
1SAM|15|16|dixit autem Samuhel ad Saul sine me et indicabo tibi quae locutus sit Dominus ad me nocte dixitque ei loquere
1SAM|15|17|et ait Samuhel nonne cum parvulus esses in oculis tuis caput in tribubus Israhel factus es unxitque te Dominus regem super Israhel
1SAM|15|18|et misit te Dominus in via et ait vade et interfice peccatores Amalech et pugnabis contra eos usque ad internicionem eorum
1SAM|15|19|quare ergo non audisti vocem Domini sed versus ad praedam es et fecisti malum in oculis Domini
1SAM|15|20|et ait Saul ad Samuhelem immo audivi vocem Domini et ambulavi in via per quam misit me Dominus et adduxi Agag regem Amalech et Amalech interfeci
1SAM|15|21|tulit autem populus de praeda oves et boves primitias eorum quae caesa sunt ut immolet Domino Deo suo in Galgalis
1SAM|15|22|et ait Samuhel numquid vult Dominus holocausta aut victimas et non potius ut oboediatur voci Domini melior est enim oboedientia quam victimae et auscultare magis quam offerre adipem arietum
1SAM|15|23|quoniam quasi peccatum ariolandi est repugnare et quasi scelus idolatriae nolle adquiescere pro eo ergo quod abiecisti sermonem Domini abiecit te ne sis rex
1SAM|15|24|dixitque Saul ad Samuhel peccavi quia praevaricatus sum sermonem Domini et verba tua timens populum et oboediens voci eorum
1SAM|15|25|sed nunc porta quaeso peccatum meum et revertere mecum ut adorem Dominum
1SAM|15|26|et ait Samuhel ad Saul non revertar tecum quia proiecisti sermonem Domini et proiecit te Dominus ne sis rex super Israhel
1SAM|15|27|et conversus est Samuhel ut abiret ille autem adprehendit summitatem pallii eius quae et scissa est
1SAM|15|28|et ait ad eum Samuhel scidit Dominus regnum Israhel a te hodie et tradidit illud proximo tuo meliori te
1SAM|15|29|porro Triumphator in Israhel non parcet et paenitudine non flectetur neque enim homo est ut agat paenitentiam
1SAM|15|30|at ille ait peccavi sed nunc honora me coram senibus populi mei et coram Israhel et revertere mecum ut adorem Dominum Deum tuum
1SAM|15|31|reversus ergo Samuhel secutus est Saulem et adoravit Saul Dominum
1SAM|15|32|dixitque Samuhel adducite ad me Agag regem Amalech et oblatus est ei Agag pinguissimus et dixit Agag sicine separat amara mors
1SAM|15|33|et ait Samuhel sicut fecit absque liberis mulieres gladius tuus sic absque liberis erit inter mulieres mater tua et in frusta concidit Samuhel Agag coram Domino in Galgalis
1SAM|15|34|abiit autem Samuhel in Ramatha Saul vero ascendit in domum suam in Gabaath
1SAM|15|35|et non vidit Samuhel ultra Saul usque ad diem mortis suae verumtamen lugebat Samuhel Saul quoniam Dominum paenitebat quod constituisset regem Saul super Israhel
1SAM|16|1|dixitque Dominus ad Samuhel usquequo tu luges Saul cum ego proiecerim eum ne regnet super Israhel imple cornu tuum oleo et veni ut mittam te ad Isai Bethleemitem providi enim in filiis eius mihi regem
1SAM|16|2|et ait Samuhel quomodo vadam audiet enim Saul et interficiet me et ait Dominus vitulum de armento tolles in manu tua et dices ad immolandum Domino veni
1SAM|16|3|et vocabis Isai ad victimam et ego ostendam tibi quid facias et ungues quemcumque monstravero tibi
1SAM|16|4|fecit ergo Samuhel sicut locutus est ei Dominus venitque in Bethleem et admirati sunt seniores civitatis occurrentes ei dixeruntque pacificus ingressus tuus
1SAM|16|5|et ait pacificus ad immolandum Domino veni sanctificamini et venite mecum ut immolem sanctificavit ergo Isai et filios eius et vocavit eos ad sacrificium
1SAM|16|6|cumque ingressi essent vidit Heliab et ait num coram Domino est christus eius
1SAM|16|7|et dixit Dominus ad Samuhel ne respicias vultum eius neque altitudinem staturae eius quoniam abieci eum nec iuxta intuitum hominis iudico homo enim videt ea quae parent Dominus autem intuetur cor
1SAM|16|8|et vocavit Isai Abinadab et adduxit eum coram Samuhel qui dixit nec hunc elegit Dominus
1SAM|16|9|adduxit autem Isai Samma de quo ait etiam hunc non elegit Dominus
1SAM|16|10|adduxit itaque Isai septem filios suos coram Samuhel et ait Samuhel ad Isai non elegit Dominus ex istis
1SAM|16|11|dixitque Samuhel ad Isai numquid iam conpleti sunt filii qui respondit adhuc reliquus est parvulus et pascit oves et ait Samuhel ad Isai mitte et adduc eum nec enim discumbemus priusquam ille huc venerit
1SAM|16|12|misit ergo et adduxit eum erat autem rufus et pulcher aspectu decoraque facie et ait Dominus surge ungue eum ipse est enim
1SAM|16|13|tulit igitur Samuhel cornu olei et unxit eum in medio fratrum eius et directus est spiritus Domini in David a die illa et in reliquum surgensque Samuhel abiit in Ramatha
1SAM|16|14|spiritus autem Domini recessit a Saul et exagitabat eum spiritus nequam a Domino
1SAM|16|15|dixeruntque servi Saul ad eum ecce spiritus Dei malus exagitat te
1SAM|16|16|iubeat dominus noster et servi tui qui coram te sunt quaerant hominem scientem psallere cithara ut quando arripuerit te spiritus Dei malus psallat manu sua et levius feras
1SAM|16|17|et ait Saul ad servos suos providete mihi aliquem bene psallentem et adducite eum ad me
1SAM|16|18|et respondens unus de pueris ait ecce vidi filium Isai Bethleemitem scientem psallere et fortissimum robore et virum bellicosum et prudentem in verbis et virum pulchrum et Dominus est cum eo
1SAM|16|19|misit ergo Saul nuntios ad Isai dicens mitte ad me David filium tuum qui est in pascuis
1SAM|16|20|tulitque Isai asinum plenum panibus et lagoenam vini et hedum de capris unum et misit per manum David filii sui Saul
1SAM|16|21|et venit David ad Saul et stetit coram eo at ille dilexit eum nimis et factus est eius armiger
1SAM|16|22|misitque Saul ad Isai dicens stet David in conspectu meo invenit enim gratiam in oculis meis
1SAM|16|23|igitur quandocumque spiritus Dei arripiebat Saul tollebat David citharam et percutiebat manu sua et refocilabatur Saul et levius habebat recedebat enim ab eo spiritus malus
1SAM|17|1|congregantes vero Philisthim agmina sua in proelium convenerunt in Soccho Iudae et castrametati sunt inter Soccho et Azeca in finibus Dommim
1SAM|17|2|porro Saul et viri Israhel congregati venerunt in valle Terebinthi et direxerunt aciem ad pugnandum contra Philisthim
1SAM|17|3|et Philisthim stabant super montem ex hac parte et Israhel stabat super montem ex altera parte vallisque erat inter eos
1SAM|17|4|et egressus est vir spurius de castris Philisthinorum nomine Goliath de Geth altitudinis sex cubitorum et palmo
1SAM|17|5|et cassis aerea super caput eius et lorica hamata induebatur porro pondus loricae eius quinque milia siclorum aeris
1SAM|17|6|et ocreas aereas habebat in cruribus et clypeus aereus tegebat umeros eius
1SAM|17|7|hastile autem hastae eius erat quasi liciatorium texentium ipsum autem ferrum hastae eius sescentos siclos habebat ferri et armiger eius antecedebat eum
1SAM|17|8|stansque clamabat adversum falangas Israhel et dicebat eis quare venitis parati ad proelium numquid ego non sum Philistheus et vos servi Saul eligite ex vobis virum et descendat ad singulare certamen
1SAM|17|9|si quiverit pugnare mecum et percusserit me erimus vobis servi si autem ego praevaluero et percussero eum vos servi eritis et servietis nobis
1SAM|17|10|et aiebat Philistheus ego exprobravi agminibus Israhelis hodie date mihi virum et ineat mecum singulare certamen
1SAM|17|11|audiens autem Saul et omnes viri israhelitae sermones Philisthei huiuscemodi stupebant et metuebant nimis
1SAM|17|12|David autem erat filius viri ephrathei de quo supra dictum est de Bethleem Iuda cui erat nomen Isai qui habebat octo filios et erat vir in diebus Saul senex et grandevus inter viros
1SAM|17|13|abierunt autem tres filii eius maiores post Saul in proelium et nomina trium filiorum eius qui perrexerant ad bellum Heliab primogenitus et secundus Abinadab tertiusque Samma
1SAM|17|14|David autem erat minimus tribus ergo maioribus secutis Saulem
1SAM|17|15|abiit David et reversus est a Saul ut pasceret gregem patris sui in Bethleem
1SAM|17|16|procedebat vero Philistheus mane et vespere et stabat quadraginta diebus
1SAM|17|17|dixit autem Isai ad David filium suum accipe fratribus tuis oephi pulentae et decem panes istos et curre in castra ad fratres tuos
1SAM|17|18|et decem formellas casei has deferes ad tribunum et fratres tuos visitabis si recte agant et cum quibus ordinati sint disce
1SAM|17|19|Saul autem et illi et omnes filii Israhel in valle Terebinthi pugnabant adversum Philisthim
1SAM|17|20|surrexit itaque David mane et commendavit gregem custodi et onustus abiit sicut praeceperat ei Isai et venit ad locum Magala et ad exercitum qui egressus ad pugnam vociferatus erat in certamine
1SAM|17|21|direxerat enim aciem Israhel sed et Philisthim ex adverso fuerant praeparati
1SAM|17|22|derelinquens ergo David vasa quae adtulerat sub manu custodis ad sarcinas cucurrit ad locum certaminis et interrogabat si omnia recte agerentur erga fratres suos
1SAM|17|23|cumque adhuc ille loqueretur eis apparuit vir ille spurius ascendens Goliath nomine Philistheus de Geth ex castris Philisthinorum et loquente eo haec eadem verba audivit David
1SAM|17|24|omnes autem Israhelitae cum vidissent virum fugerunt a facie eius timentes eum valde
1SAM|17|25|et dixit unus quispiam de Israhel num vidisti virum hunc qui ascendit ad exprobrandum enim Israheli ascendit virum ergo qui percusserit eum ditabit rex divitiis magnis et filiam suam dabit ei et domum patris eius faciet absque tributo in Israhel
1SAM|17|26|et ait David ad viros qui stabant secum dicens quid dabitur viro qui percusserit Philistheum hunc et tulerit obprobrium de Israhel quis est enim hic Philistheus incircumcisus qui exprobravit acies Dei viventis
1SAM|17|27|referebat autem ei populus eundem sermonem dicens haec dabuntur viro qui percusserit eum
1SAM|17|28|quod cum audisset Heliab frater eius maior loquente eo cum aliis iratus est contra David et ait quare venisti et quare dereliquisti pauculas oves illas in deserto ego novi superbiam tuam et nequitiam cordis tui quia ut videres proelium descendisti
1SAM|17|29|et dixit David quid feci numquid non verbum est
1SAM|17|30|et declinavit paululum ab eo ad alium dixitque eundem sermonem et respondit ei populus verbum sicut et prius
1SAM|17|31|audita sunt autem verba quae locutus est David et adnuntiata in conspectu Saul
1SAM|17|32|ad quem cum fuisset adductus locutus est ei non concidat cor cuiusquam in eo ego servus tuus vadam et pugnabo adversus Philistheum
1SAM|17|33|et ait Saul ad David non vales resistere Philistheo isti nec pugnare adversum eum quia puer es hic autem vir bellator ab adulescentia sua
1SAM|17|34|dixitque David ad Saul pascebat servus tuus patris sui gregem et veniebat leo vel ursus tollebatque arietem de medio gregis
1SAM|17|35|et sequebar eos et percutiebam eruebamque de ore eorum et illi consurgebant adversum me et adprehendebam mentum eorum et suffocabam interficiebamque eos
1SAM|17|36|nam et leonem et ursum interfeci ego servus tuus erit igitur et Philistheus hic incircumcisus quasi unus ex eis quia ausus est maledicere exercitum Dei viventis
1SAM|17|37|et ait David Dominus qui eruit me de manu leonis et de manu ursi ipse liberabit me de manu Philisthei huius dixit autem Saul ad David vade et Dominus tecum sit
1SAM|17|38|et induit Saul David vestimentis suis et inposuit galeam aeream super caput eius et vestivit eum lorica
1SAM|17|39|accinctus ergo David gladio eius super veste sua coepit temptare si armatus posset incedere non enim habebat consuetudinem dixitque David ad Saul non possum sic incedere quia nec usum habeo et deposuit ea
1SAM|17|40|et tulit baculum suum quem semper habebat in manibus et elegit sibi quinque limpidissimos lapides de torrente et misit eos in peram pastoralem quam habebat secum et fundam manu tulit et processit adversum Philistheum
1SAM|17|41|ibat autem Philistheus incedens et adpropinquans adversum David et armiger eius ante eum
1SAM|17|42|cumque inspexisset Philistheus et vidisset David despexit eum erat enim adulescens rufus et pulcher aspectu
1SAM|17|43|et dixit Philistheus ad David numquid ego canis sum quod tu venis ad me cum baculo et maledixit Philistheus David in diis suis
1SAM|17|44|dixitque ad David veni ad me et dabo carnes tuas volatilibus caeli et bestiis terrae
1SAM|17|45|dixit autem David ad Philistheum tu venis ad me cum gladio et hasta et clypeo ego autem venio ad te in nomine Domini exercituum Dei agminum Israhel quibus exprobrasti
1SAM|17|46|hodie et dabit te Dominus in manu mea et percutiam te et auferam caput tuum a te et dabo cadaver castrorum Philisthim hodie volatilibus caeli et bestiis terrae ut sciat omnis terra quia est Deus in Israhel
1SAM|17|47|et noverit universa ecclesia haec quia non in gladio nec in hasta salvat Dominus ipsius est enim bellum et tradet vos in manus nostras
1SAM|17|48|cum ergo surrexisset Philistheus et veniret et adpropinquaret contra David festinavit David et cucurrit ad pugnam ex adverso Philisthei
1SAM|17|49|et misit manum suam in peram tulitque unum lapidem et funda iecit et percussit Philistheum in fronte et infixus est lapis in fronte eius et cecidit in faciem suam super terram
1SAM|17|50|praevaluitque David adversus Philistheum in funda et in lapide percussumque Philistheum interfecit cumque gladium non haberet in manu David
1SAM|17|51|cucurrit et stetit super Philistheum et tulit gladium eius et eduxit de vagina sua et interfecit eum praeciditque caput eius videntes autem Philisthim quod mortuus esset fortissimus eorum fugerunt
1SAM|17|52|et consurgentes viri Israhel et Iuda vociferati sunt et persecuti Philistheos usque dum venirent in vallem et usque ad portas Accaron cecideruntque vulnerati de Philisthim in via Sarim usque ad Geth et usque Accaron
1SAM|17|53|et revertentes filii Israhel postquam persecuti fuerant Philistheos invaserunt castra eorum
1SAM|17|54|adsumens autem David caput Philisthei adtulit illud in Hierusalem arma vero eius posuit in tabernaculo suo
1SAM|17|55|eo autem tempore quo viderat Saul David egredientem contra Philistheum ait ad Abner principem militiae de qua stirpe descendit hic adulescens Abner dixitque Abner vivit anima tua rex si novi
1SAM|17|56|et ait rex interroga tu cuius filius sit iste puer
1SAM|17|57|cumque regressus esset David percusso Philistheo tulit eum Abner et introduxit coram Saul caput Philisthei habentem in manu
1SAM|17|58|et ait ad eum Saul de qua progenie es o adulescens dixitque David filius servi tui Isai Bethleemitae ego sum
1SAM|18|1|et factum est cum conplesset loqui ad Saul anima Ionathan conligata est animae David et dilexit eum Ionathan quasi animam suam
1SAM|18|2|tulitque eum Saul in die illa et non concessit ei ut reverteretur in domum patris sui
1SAM|18|3|inierunt autem Ionathan et David foedus diligebat enim eum quasi animam suam
1SAM|18|4|nam expoliavit se Ionathan tunicam qua erat vestitus et dedit eam David et reliqua vestimenta sua usque ad gladium et arcum suum et usque ad balteum
1SAM|18|5|egrediebatur quoque David ad omnia quaecumque misisset eum Saul et prudenter se agebat posuitque eum Saul super viros belli et acceptus erat in oculis universi populi maximeque in conspectu famulorum Saul
1SAM|18|6|porro cum reverteretur percusso Philistheo David egressae sunt mulieres de universis urbibus Israhel cantantes chorosque ducentes in occursum Saul regis in tympanis laetitiae et in sistris
1SAM|18|7|et praecinebant mulieres ludentes atque dicentes percussit Saul mille et David decem milia
1SAM|18|8|iratus est autem Saul nimis et displicuit in oculis eius iste sermo dixitque dederunt David decem milia et mihi dederunt mille quid ei superest nisi solum regnum
1SAM|18|9|non rectis ergo oculis Saul aspiciebat David ex die illa et deinceps
1SAM|18|10|post diem autem alteram invasit spiritus Dei malus Saul et prophetabat in medio domus suae David autem psallebat manu sua sicut per singulos dies tenebatque Saul lanceam
1SAM|18|11|et misit eam putans quod configere posset David cum pariete et declinavit David a facie eius secundo
1SAM|18|12|et timuit Saul David eo quod esset Dominus cum eo et a se recessisset
1SAM|18|13|amovit ergo eum Saul a se et fecit eum tribunum super mille viros et egrediebatur et intrabat in conspectu populi
1SAM|18|14|in omnibus quoque viis suis David prudenter agebat et Dominus erat cum eo
1SAM|18|15|vidit itaque Saul quod prudens esset nimis et coepit cavere eum
1SAM|18|16|omnis autem Israhel et Iuda diligebat David ipse enim egrediebatur et ingrediebatur ante eos
1SAM|18|17|dixit autem Saul ad David ecce filia mea maior Merob ipsam dabo tibi uxorem tantummodo esto vir fortis et proeliare bella Domini Saul autem reputabat dicens non sit manus mea in eo sed sit super illum manus Philisthinorum
1SAM|18|18|ait autem David ad Saul quis ego sum aut quae est vita mea aut cognatio patris mei in Israhel ut fiam gener regis
1SAM|18|19|factum est autem tempus cum deberet dari Merob filia Saul David data est Hadrihel Molathitae uxor
1SAM|18|20|dilexit autem Michol filia Saul altera David et nuntiatum est Saul et placuit ei
1SAM|18|21|dixitque Saul dabo eam illi ut fiat ei in scandalum et sit super eum manus Philisthinorum dixit ergo Saul ad David in duabus rebus gener meus eris hodie
1SAM|18|22|et mandavit Saul servis suis loquimini ad David clam me dicentes ecce places regi et omnes servi eius diligunt te nunc ergo esto gener regis
1SAM|18|23|et locuti sunt servi Saul in auribus David omnia verba haec et ait David num parum vobis videtur generum esse regis ego autem sum vir pauper et tenuis
1SAM|18|24|et renuntiaverunt servi Saul dicentes huiuscemodi verba locutus est David
1SAM|18|25|dixit autem Saul sic loquimini ad David non habet necesse rex sponsalia nisi tantum centum praeputia Philisthinorum ut fiat ultio de inimicis regis porro Saul cogitabat tradere David in manibus Philisthinorum
1SAM|18|26|cumque renuntiassent servi eius David verba quae diximus placuit sermo in oculis David ut fieret gener regis
1SAM|18|27|et post dies paucos surgens David abiit cum viris qui sub eo erant et percussis Philisthim ducentis viris adtulit praeputia eorum et adnumeravit ea regi ut esset gener eius dedit itaque ei Saul Michol filiam suam uxorem
1SAM|18|28|et vidit Saul et intellexit quia Dominus esset cum David Michol autem filia Saul diligebat eum
1SAM|18|29|et Saul magis coepit timere David factusque est Saul inimicus David cunctis diebus
1SAM|18|30|et egressi sunt principes Philisthinorum a principio autem egressionis eorum prudentius se gerebat David quam omnes servi Saul et celebre factum est nomen eius nimis
1SAM|19|1|locutus est autem Saul ad Ionathan filium suum et ad omnes servos suos ut occiderent David porro Ionathan filius Saul diligebat David valde
1SAM|19|2|et indicavit Ionathan David dicens quaerit Saul pater meus occidere te quapropter observa te quaeso mane et manebis clam et absconderis
1SAM|19|3|ego autem egrediens stabo iuxta patrem meum in agro ubicumque fueris et ego loquar de te ad patrem meum et quodcumque videro nuntiabo tibi
1SAM|19|4|locutus est ergo Ionathan de David bona ad Saul patrem suum dixitque ad eum ne pecces rex in servum tuum David quia non peccavit tibi et opera eius bona sunt tibi valde
1SAM|19|5|et posuit animam suam in manu sua et percussit Philistheum et fecit Dominus salutem magnam universo Israhel vidisti et laetatus es quare ergo peccas in sanguine innoxio interficiens David qui est absque culpa
1SAM|19|6|quod cum audisset Saul placatus voce Ionathae iuravit vivit Dominus quia non occidetur
1SAM|19|7|vocavit itaque Ionathan David et indicavit ei omnia verba haec et introduxit Ionathan David ad Saul et fuit ante eum sicut fuerat heri et nudius tertius
1SAM|19|8|motum est autem rursus bellum et egressus David pugnavit adversus Philisthim percussitque eos plaga magna et fugerunt a facie eius
1SAM|19|9|et factus est spiritus Domini malus in Saul sedebat autem in domo sua et tenebat lanceam porro David psallebat in manu sua
1SAM|19|10|nisusque est Saul configere lancea David in pariete et declinavit David a facie Saul lancea autem casso vulnere perlata est in parietem et David fugit et salvatus est nocte illa
1SAM|19|11|misit ergo Saul satellites suos in domum David ut custodirent eum et interficeretur mane quod cum adnuntiasset David Michol uxor sua dicens nisi salvaveris te nocte hac cras morieris
1SAM|19|12|deposuit eum per fenestram porro ille abiit et aufugit atque salvatus est
1SAM|19|13|tulit autem Michol statuam et posuit eam super lectum et pellem pilosam caprarum posuit ad caput eius et operuit eam vestimentis
1SAM|19|14|misit autem Saul apparitores qui raperent David et responsum est quod aegrotaret
1SAM|19|15|rursumque misit Saul nuntios ut viderent David dicens adferte eum ad me in lecto ut occidatur
1SAM|19|16|cumque venissent nuntii inventum est simulacrum super lectum et pellis caprarum ad caput eius
1SAM|19|17|dixitque Saul ad Michol quare sic inlusisti mihi et dimisisti inimicum meum ut fugeret et respondit Michol ad Saul quia ipse locutus est mihi dimitte me alioquin interficiam te
1SAM|19|18|David autem fugiens salvatus est et venit ad Samuhel in Ramatha et nuntiavit ei omnia quae fecerat sibi Saul et abierunt ipse et Samuhel et morati sunt in Nahioth
1SAM|19|19|nuntiatum est autem Sauli a dicentibus ecce David in Nahioth in Rama
1SAM|19|20|misit ergo Saul lictores ut raperent David qui cum vidissent cuneum prophetarum vaticinantium et Samuhel stantem super eos factus est etiam in illis spiritus Domini et prophetare coeperunt etiam ipsi
1SAM|19|21|quod cum nuntiatum esset Sauli misit alios nuntios prophetaverunt autem et illi et rursum Saul misit tertios nuntios qui et ipsi prophetaverunt
1SAM|19|22|abiit autem etiam ipse in Ramatha et venit usque ad cisternam magnam quae est in Soccho et interrogavit et dixit in quo loco sunt Samuhel et David dictumque est ei ecce in Nahioth sunt in Rama
1SAM|19|23|et abiit in Nahioth in Rama et factus est etiam super eum spiritus Dei et ambulabat ingrediens et prophetabat usque dum veniret in Nahioth in Rama
1SAM|19|24|et expoliavit se etiam ipse vestimentis suis et prophetavit cum ceteris coram Samuhel et cecidit nudus tota die illa et nocte unde et exivit proverbium num et Saul inter prophetas
1SAM|20|1|fugit autem David de Nahioth quae erat in Rama veniensque locutus est coram Ionathan quid feci quae est iniquitas mea et quod peccatum meum in patrem tuum quia quaerit animam meam
1SAM|20|2|qui dixit ei absit non morieris neque enim faciet pater meus quicquam grande vel parvum nisi prius indicaverit mihi hunc ergo celavit me pater meus sermonem tantummodo nequaquam erit istud
1SAM|20|3|et iuravit rursum David et ille ait scit profecto pater tuus quia inveni gratiam in oculis tuis et dicet nesciat hoc Ionathan ne forte tristetur quinimmo vivit Dominus et vivit anima tua quia uno tantum ut ita dicam gradu ego morsque dividimur
1SAM|20|4|et ait Ionathan ad David quodcumque dixerit mihi anima tua faciam tibi
1SAM|20|5|dixit autem David ad Ionathan ecce kalendae sunt crastino et ego ex more sedere soleo iuxta regem ad vescendum dimitte ergo me ut abscondar in agro usque ad vesperam diei tertiae
1SAM|20|6|si requisierit me pater tuus respondebis ei rogavit me David ut iret celeriter in Bethleem civitatem suam quia victimae sollemnes ibi sunt universis contribulibus eius
1SAM|20|7|si dixerit bene pax erit servo tuo si autem fuerit iratus scito quia conpleta est malitia eius
1SAM|20|8|fac ergo misericordiam in servum tuum quia foedus Domini me famulum tuum tecum inire fecisti si autem est in me aliqua iniquitas tu me interfice et ad patrem tuum ne introducas me
1SAM|20|9|et ait Ionathan absit hoc a te neque enim fieri potest ut si certo cognovero conpletam patris mei esse malitiam contra te non adnuntiem tibi
1SAM|20|10|responditque David ad Ionathan quis nuntiabit mihi si quid forte responderit tibi pater tuus dure
1SAM|20|11|et ait Ionathan ad David veni egrediamur in agrum cumque exissent ambo in agrum
1SAM|20|12|ait Ionathan ad David Domine Deus Israhel si investigavero sententiam patris mei crastino vel perendie et aliquid boni fuerit super David et non statim misero ad te et notum tibi fecero
1SAM|20|13|haec faciat Dominus Ionathan et haec augeat si autem perseveraverit patris mei malitia adversum te revelabo aurem tuam et dimittam te ut vadas in pace et sit Dominus tecum sicut fuit cum patre meo
1SAM|20|14|et si vixero facies mihi misericordiam Domini si vero mortuus fuero
1SAM|20|15|non auferas misericordiam tuam a domo mea usque in sempiternum quando eradicaverit Dominus inimicos David unumquemque de terra
1SAM|20|16|pepigit ergo foedus Ionathan cum domo David et requisivit Dominus de manu inimicorum David
1SAM|20|17|et addidit Ionathan deierare David eo quod diligeret illum sicut animam enim suam ita diligebat eum
1SAM|20|18|dixitque ad eum Ionathan cras kalendae sunt et requireris
1SAM|20|19|requiretur enim sessio tua usque perendie descendes ergo festinus et venies in locum ubi celandus es in die qua operari licet et sedebis iuxta lapidem cui est nomen Ezel
1SAM|20|20|et ego tres sagittas mittam iuxta eum et iaciam quasi exercens me ad signum
1SAM|20|21|mittam quoque et puerum dicens ei vade et adfer mihi sagittas
1SAM|20|22|si dixero puero ecce sagittae intra te sunt tolle eas tu veni ad me quia pax tibi est et nihil est mali vivit Dominus si autem sic locutus fuero puero ecce sagittae ultra te sunt vade quia dimisit te Dominus
1SAM|20|23|de verbo autem quod locuti fuimus ego et tu sit Dominus inter me et te usque in sempiternum
1SAM|20|24|absconditus est ergo David in agro et venerunt kalendae et sedit rex ad comedendum panem
1SAM|20|25|cumque sedisset rex super cathedram suam secundum consuetudinem quae erat iuxta parietem surrexit Ionathan et sedit Abner ex latere Saul vacuusque apparuit locus David
1SAM|20|26|et non est locutus Saul quicquam in die illa cogitabat enim quod forte evenisset ei ut non esset mundus nec purificatus
1SAM|20|27|cumque inluxisset dies secunda post kalendas rursum vacuus apparuit locus David dixitque Saul ad Ionathan filium suum cur non venit filius Isai nec heri nec hodie ad vescendum
1SAM|20|28|et respondit Ionathan Sauli rogavit me obnixe ut iret in Bethleem
1SAM|20|29|et ait dimitte me quoniam sacrificium sollemne est in civitate unus de fratribus meis accersivit me nunc ergo si inveni gratiam in oculis tuis vadam cito et videbo fratres meos ob hanc causam non venit ad mensam regis
1SAM|20|30|iratus autem Saul adversus Ionathan dixit ei fili mulieris virum ultro rapientis numquid ignoro quia diligis filium Isai in confusionem tuam et in confusionem ignominiosae matris tuae
1SAM|20|31|omnibus enim diebus quibus filius Isai vixerit super terram non stabilieris tu neque regnum tuum itaque iam nunc mitte et adduc eum ad me quia filius mortis est
1SAM|20|32|respondens autem Ionathan Sauli patri suo ait quare moritur quid fecit
1SAM|20|33|et arripuit Saul lanceam ut percuteret eum et intellexit Ionathan quod definitum esset patri suo ut interficeret David
1SAM|20|34|surrexit ergo Ionathan a mensa in ira furoris et non comedit in die kalendarum secunda panem contristatus est enim super David eo quod confudisset eum pater suus
1SAM|20|35|cumque inluxisset mane venit Ionathan in agrum iuxta placitum David et puer parvulus cum eo
1SAM|20|36|et ait ad puerum suum vade et adfer mihi sagittas quas ego iacio cumque puer cucurrisset iecit aliam sagittam trans puerum
1SAM|20|37|venit itaque puer ad locum iaculi quod miserat Ionathan et clamavit Ionathan post tergum pueri et ait ecce ibi est sagitta porro ultra te
1SAM|20|38|clamavitque Ionathan post tergum pueri festina velociter ne steteris collegit autem puer Ionathae sagittas et adtulit ad dominum suum
1SAM|20|39|et quid ageretur penitus ignorabat tantummodo enim Ionathan et David rem noverant
1SAM|20|40|dedit igitur Ionathan arma sua puero et dixit ei vade defer in civitatem
1SAM|20|41|cumque abisset puer surrexit David de loco qui vergebat ad austrum et cadens pronus in terram adoravit tertio et osculantes alterutrum fleverunt pariter David autem amplius
1SAM|20|42|dixit ergo Ionathan ad David vade in pace quaecumque iuravimus ambo in nomine Domini dicentes Dominus sit inter me et te et inter semen meum et semen tuum usque in sempiternum
1SAM|20|43|et surrexit et abiit sed et Ionathan ingressus est civitatem
1SAM|21|1|venit autem David in Nobe ad Ahimelech sacerdotem et obstipuit Ahimelech eo quod venisset David et dixit ei quare tu solus et nullus est tecum
1SAM|21|2|et ait David ad Ahimelech sacerdotem rex praecepit mihi sermonem et dixit nemo sciat rem propter quam a me missus es et cuiusmodi tibi praecepta dederim nam et pueris condixi in illum et illum locum
1SAM|21|3|nunc igitur si quid habes ad manum vel quinque panes da mihi aut quicquid inveneris
1SAM|21|4|et respondens sacerdos David ait ei non habeo panes laicos ad manum sed tantum panem sanctum si mundi sunt pueri maxime a mulieribus
1SAM|21|5|et respondit David sacerdoti et dixit ei equidem si de mulieribus agitur continuimus nos ab heri et nudius tertius quando egrediebamur et fuerunt vasa puerorum sancta porro via haec polluta est sed et ipsa hodie sanctificabitur in vasis
1SAM|21|6|dedit ergo ei sacerdos sanctificatum panem neque enim erat ibi panis nisi tantum panes propositionis qui sublati fuerant a facie Domini ut ponerentur panes calidi
1SAM|21|7|erat autem ibi vir de servis Saul in die illa intus in tabernaculo Domini et nomen eius Doec Idumeus potentissimus pastorum Saul
1SAM|21|8|dixit autem David ad Ahimelech si habes hic ad manum hastam aut gladium quia gladium meum et arma mea non tuli mecum sermo enim regis urguebat
1SAM|21|9|et dixit sacerdos gladius Goliath Philisthei quem percussisti in valle Terebinthi est involutus pallio post ephod si istum vis tollere tolle neque enim est alius hic absque eo et ait David non est huic alter similis da mihi eum
1SAM|21|10|surrexit itaque David et fugit in die illa a facie Saul et venit ad Achis regem Geth
1SAM|21|11|dixeruntque ei servi Achis numquid non iste est David rex terrae nonne huic cantabant per choros dicentes percussit Saul mille et David decem milia
1SAM|21|12|posuit autem David sermones istos in corde suo et extimuit valde a facie Achis regis Geth
1SAM|21|13|et inmutavit os suum coram eis et conlabebatur inter manus eorum et inpingebat in ostia portae defluebantque salivae eius in barbam
1SAM|21|14|et ait Achis ad servos suos vidistis hominem insanum quare adduxistis eum ad me
1SAM|21|15|an desunt nobis furiosi quod introduxistis istum ut fureret me praesente hicine ingredietur domum meam
1SAM|22|1|abiit ergo inde David et fugit in speluncam Odollam quod cum audissent fratres eius et omnis domus patris eius descenderunt ad eum illuc
1SAM|22|2|et convenerunt ad eum omnes qui erant in angustia constituti et oppressi aere alieno et amaro animo et factus est eorum princeps fueruntque cum eo quasi quadringenti viri
1SAM|22|3|et profectus est David inde in Maspha quae est Moab et dixit ad regem Moab maneat oro pater meus et mater mea vobiscum donec sciam quid faciat mihi Deus
1SAM|22|4|et reliquit eos ante faciem regis Moab manseruntque apud eum cunctis diebus quibus David fuit in praesidio
1SAM|22|5|dixitque Gad propheta ad David noli manere in praesidio proficiscere et vade in terram Iuda et profectus David venit in saltum Hareth
1SAM|22|6|et audivit Saul quod apparuisset David et viri qui erant cum eo Saul autem cum maneret in Gabaa et esset in nemore quod est in Rama hastam manu tenens cunctique socii eius circumstarent eum
1SAM|22|7|ait ad servos suos qui adsistebant ei audite filii Iemini numquid omnibus vobis dabit filius Isai agros et vineas et universos vos faciet tribunos et centuriones
1SAM|22|8|quoniam coniurastis omnes adversum me et non est qui mihi renuntiet maxime cum et filius meus foedus iunxerit cum filio Isai non est qui vicem meam doleat ex vobis nec qui adnuntiet mihi eo quod suscitaverit filius meus servum meum adversum me insidiantem mihi usque hodie
1SAM|22|9|respondens autem Doec Idumeus qui adsistebat et erat primus inter servos Saul vidi inquit filium Isai in Nobe apud Ahimelech filium Achitob
1SAM|22|10|qui consuluit pro eo Dominum et cibaria dedit ei sed et gladium Goliath Philisthei dedit illi
1SAM|22|11|misit ergo rex ad accersiendum Ahimelech filium Achitob sacerdotem et omnem domum patris eius sacerdotum qui erant in Nobe qui venerunt universi ad regem
1SAM|22|12|et ait Saul audi fili Achitob qui respondit praesto sum domine
1SAM|22|13|dixitque ad eum Saul quare coniurastis adversum me tu et filius Isai et dedisti ei panes et gladium et consuluisti pro eo Deum ut consurgeret adversum me insidiator usque hodie permanens
1SAM|22|14|respondensque Ahimelech regi ait et quis in omnibus servis tuis sicut David fidelis et gener regis et pergens ad imperium tuum et gloriosus in domo tua
1SAM|22|15|num hodie coepi consulere pro eo Deum absit hoc a me ne suspicetur rex adversus servum suum rem huiuscemodi in universa domo patris mei non enim scivit servus tuus quicquam super hoc negotio vel modicum vel grande
1SAM|22|16|dixitque rex morte morieris Ahimelech tu et omnis domus patris tui
1SAM|22|17|et ait rex emissariis qui circumstabant eum convertimini et interficite sacerdotes Domini nam manus eorum cum David est scientes quod fugisset non indicaverunt mihi noluerunt autem servi regis extendere manum suam in sacerdotes Domini
1SAM|22|18|et ait rex Doec convertere tu et inrue in sacerdotes conversusque Doec Idumeus inruit in sacerdotes et trucidavit in die illa octoginta quinque viros vestitos ephod lineo
1SAM|22|19|Nobe autem civitatem sacerdotum percussit in ore gladii viros et mulieres parvulos et lactantes bovem et asinum et ovem in ore gladii
1SAM|22|20|evadens autem unus filius Ahimelech filii Achitob cuius nomen erat Abiathar fugit ad David
1SAM|22|21|et adnuntiavit ei quod occidisset Saul sacerdotes Domini
1SAM|22|22|et ait David ad Abiathar sciebam in die illa quod cum ibi esset Doec Idumeus procul dubio adnuntiaret Saul ego sum reus omnium animarum patris tui
1SAM|22|23|mane mecum ne timeas si quis quaesierit animam meam quaeret et animam tuam mecumque servaberis
1SAM|23|1|et nuntiaverunt David dicentes ecce Philisthim obpugnant Ceila et diripiunt areas
1SAM|23|2|consuluit igitur David Dominum dicens num vadam et percutiam Philistheos istos et ait Dominus ad David vade et percuties Philistheos et salvabis Ceila
1SAM|23|3|et dixerunt viri qui erant cum David ad eum ecce nos hic in Iudaea consistentes timemus quanto magis si ierimus in Ceila adversum agmina Philisthinorum
1SAM|23|4|rursum ergo David consuluit Dominum qui respondens ei ait surge et vade in Ceila ego enim tradam Philistheos in manu tua
1SAM|23|5|abiit David et viri eius in Ceila et pugnavit adversum Philistheos et abegit iumenta eorum et percussit eos plaga magna et salvavit David habitatores Ceilae
1SAM|23|6|porro eo tempore quo fugiebat Abiathar filius Ahimelech ad David in Ceila ephod secum habens descenderat
1SAM|23|7|nuntiatum est autem Saul quod venisset David in Ceila et ait Saul tradidit eum Deus in manus meas conclususque est introgressus urbem in qua portae et serae
1SAM|23|8|et praecepit Saul omni populo ut ad pugnam descenderet in Ceila et obsideret David et viros eius
1SAM|23|9|quod cum rescisset David quia praepararet ei Saul clam malum dixit ad Abiathar sacerdotem adplica ephod
1SAM|23|10|et ait David Domine Deus Israhel audivit famam servus tuus quod disponat Saul venire ad Ceila ut evertat urbem propter me
1SAM|23|11|si tradent me viri Ceila in manus eius et si descendet Saul sicut audivit servus tuus Domine Deus Israhel indica servo tuo et ait Dominus descendet
1SAM|23|12|dixitque David si tradent viri Ceilae me et viros qui sunt mecum in manu Saul et dixit Dominus tradent
1SAM|23|13|surrexit ergo David et viri eius quasi sescenti et egressi de Ceila huc atque illuc vagabantur incerti nuntiatumque est Saul quod fugisset David de Ceila quam ob rem dissimulavit exire
1SAM|23|14|morabatur autem David in deserto in locis firmissimis mansitque in monte solitudinis Ziph quaerebat tamen eum Saul cunctis diebus et non tradidit eum Deus in manus eius
1SAM|23|15|et vidit David quod egressus esset Saul ut quaereret animam eius porro David erat in deserto Ziph in silva
1SAM|23|16|et surrexit Ionathan filius Saul et abiit ad David in silva et confortavit manus eius in Deo dixitque ei
1SAM|23|17|ne timeas neque enim inveniet te manus Saul patris mei et tu regnabis super Israhel et ego ero tibi secundus sed et Saul pater meus scit hoc
1SAM|23|18|percussit igitur uterque foedus coram Domino mansitque David in silva Ionathas autem reversus est in domum suam
1SAM|23|19|ascenderunt autem Ziphei ad Saul in Gabaa dicentes nonne David latitat apud nos in locis tutissimis silvae in colle Achilae quae est ad dexteram deserti
1SAM|23|20|nunc ergo sicut desideravit anima tua ut descenderes descende nostrum autem erit ut tradamus eum in manus regis
1SAM|23|21|dixitque Saul benedicti vos a Domino quia doluistis vicem meam
1SAM|23|22|abite oro et diligentius praeparate et curiosius agite et considerate locum ubi sit pes eius vel quis viderit eum ibi recogitat enim de me quod callide insidier ei
1SAM|23|23|considerate et videte omnia latibula eius in quibus absconditur et revertimini ad me ad rem certam ut vadam vobiscum quod si etiam in terra se abstruserit perscrutabor eum in cunctis milibus Iuda
1SAM|23|24|at illi surgentes abierunt in Ziph ante Saul David autem et viri eius erant in deserto Maon in campestribus ad dextram Iesimuth
1SAM|23|25|ivit ergo Saul et socii eius ad quaerendum et nuntiatum est David statimque descendit ad petram et versabatur in deserto Maon quod cum audisset Saul persecutus est David in deserto Maon
1SAM|23|26|et ibat Saul ad latus montis ex parte una David autem et viri eius erant in latere montis ex parte altera porro David desperabat se posse evadere a facie Saul itaque Saul et viri eius in modum coronae cingebant David et viros eius ut caperent eos
1SAM|23|27|et nuntius venit ad Saul dicens festina et veni quoniam infuderunt se Philisthim super terram
1SAM|23|28|reversus est ergo Saul desistens persequi David et perrexit in occursum Philisthinorum propter hoc vocaverunt locum illum petram Dividentem
1SAM|24|1|ascendit ergo David inde et habitavit in locis tutissimis Engaddi
1SAM|24|2|cumque reversus esset Saul postquam persecutus est Philistheos nuntiaverunt ei dicentes ecce David in deserto est Engaddi
1SAM|24|3|adsumens ergo Saul tria milia electorum virorum ex omni Israhel perrexit ad investigandum David et viros eius etiam super abruptissimas petras quae solis hibicibus perviae sunt
1SAM|24|4|et venit ad caulas quoque ovium quae se offerebant vianti eratque ibi spelunca quam ingressus est Saul ut purgaret ventrem porro David et viri eius in interiori parte speluncae latebant
1SAM|24|5|et dixerunt servi David ad eum ecce dies de qua locutus est Dominus ad te ego tradam tibi inimicum tuum ut facias ei sicut placuerit in oculis tuis surrexit ergo David et praecidit oram clamydis Saul silenter
1SAM|24|6|post haec percussit cor suum David eo quod abscidisset oram clamydis Saul
1SAM|24|7|dixitque ad viros suos propitius mihi sit Dominus ne faciam hanc rem domino meo christo Domini ut mittam manum meam in eum quoniam christus Domini est
1SAM|24|8|et confregit David viros suos sermonibus et non permisit eos ut consurgerent in Saul porro Saul exsurgens de spelunca pergebat coepto itinere
1SAM|24|9|surrexit autem et David post eum et egressus de spelunca clamavit post tergum Saul dicens domine mi rex et respexit Saul post se et inclinans se David pronus in terram adoravit
1SAM|24|10|dixitque ad Saul quare audis verba hominum loquentium David quaerit malum adversum te
1SAM|24|11|ecce hodie viderunt oculi tui quod tradiderit te Dominus in manu mea in spelunca et cogitavi ut occiderem te sed pepercit tibi oculus meus dixi enim non extendam manum meam in domino meo quia christus Domini est
1SAM|24|12|quin potius pater mi vide et cognosce oram clamydis tuae in manu mea quoniam cum praeciderem summitatem clamydis tuae nolui extendere manum meam in te animadverte et vide quoniam non est in manu mea malum neque iniquitas neque peccavi in te tu autem insidiaris animae meae ut auferas eam
1SAM|24|13|iudicet Dominus inter me et te et ulciscatur me Dominus ex te manus autem mea non sit in te
1SAM|24|14|sicut et in proverbio antiquo dicitur ab impiis egredietur impietas manus ergo mea non sit in te
1SAM|24|15|quem sequeris rex Israhel quem persequeris canem mortuum sequeris et pulicem unum
1SAM|24|16|sit Dominus iudex et iudicet inter me et te et videat et diiudicet causam meam et eruat me de manu tua
1SAM|24|17|cum autem conplesset David loquens sermones huiuscemodi ad Saul dixit Saul numquid vox haec tua est fili mi David et levavit Saul vocem suam et flevit
1SAM|24|18|dixitque ad David iustior tu es quam ego tu enim tribuisti mihi bona ego autem reddidi tibi mala
1SAM|24|19|et tu indicasti hodie quae feceris mihi bona quomodo tradiderit me Dominus in manu tua et non occideris me
1SAM|24|20|quis enim cum invenerit inimicum suum dimittet eum in via bona sed Dominus reddat tibi vicissitudinem hanc pro eo quod hodie operatus es in me
1SAM|24|21|et nunc quia scio quod certissime regnaturus sis et habiturus in manu tua regnum Israhel
1SAM|24|22|iura mihi in Domino ne deleas semen meum post me neque auferas nomen meum de domo patris mei
1SAM|24|23|et iuravit David Sauli abiit ergo Saul in domum suam et David et viri eius ascenderunt ad tutiora loca
1SAM|25|1|mortuus est autem Samuhel et congregatus est universus Israhel et planxerunt eum et sepelierunt in domo sua in Rama consurgensque David descendit in desertum Pharan
1SAM|25|2|erat autem vir quispiam in solitudine Maon et possessio eius in Carmelo et homo ille magnus nimis erantque ei oves tria milia et mille caprae et accidit ut tonderetur grex eius in Carmelo
1SAM|25|3|nomen autem viri illius erat Nabal et nomen uxoris eius Abigail eratque mulier illa prudentissima et speciosa porro vir eius durus et pessimus et malitiosus erat autem de genere Chaleb
1SAM|25|4|cum ergo audisset David in deserto quod tonderet Nabal gregem suum
1SAM|25|5|misit decem iuvenes et dixit eis ascendite in Carmelum et venietis ad Nabal et salutabitis eum ex nomine meo pacifice
1SAM|25|6|et dicetis sic fratribus meis et tibi pax et domui tuae pax et omnibus quaecumque habes sit pax
1SAM|25|7|audivi quod tonderent pastores tui qui erant nobiscum in deserto numquam eis molesti fuimus nec aliquando defuit eis quicquam de grege omni tempore quo fuerunt nobiscum in Carmelo
1SAM|25|8|interroga pueros tuos et indicabunt tibi nunc ergo inveniant pueri gratiam in oculis tuis in die enim bona venimus quodcumque invenerit manus tua da servis tuis et filio tuo David
1SAM|25|9|cumque venissent pueri David locuti sunt ad Nabal omnia verba haec ex nomine David et siluerunt
1SAM|25|10|respondens autem Nabal pueris David ait quis est David et quis est filius Isai hodie increverunt servi qui fugiunt dominos suos
1SAM|25|11|tollam ergo panes meos et aquas meas et carnes pecorum quae occidi tonsoribus meis et dabo viris quos nescio unde sint
1SAM|25|12|regressi sunt itaque pueri David per viam suam et reversi venerunt et nuntiaverunt ei omnia verba quae dixerat
1SAM|25|13|tunc David ait viris suis accingatur unusquisque gladio suo et accincti sunt singuli gladio suo accinctusque est et David ense suo et secuti sunt David quasi quadringenti viri porro ducenti remanserunt ad sarcinas
1SAM|25|14|Abigail autem uxori Nabal nuntiavit unus de pueris dicens ecce misit David nuntios de deserto ut benedicerent domino nostro et aversus est eos
1SAM|25|15|homines isti boni satis fuerunt nobis et non molesti nec quicquam aliquando periit omni tempore quo sumus conversati cum eis in deserto
1SAM|25|16|pro muro erant nobis tam in nocte quam in die omnibus diebus quibus pavimus apud eos greges
1SAM|25|17|quam ob rem considera et recogita quid facias quoniam conpleta est malitia adversum virum tuum et adversus domum tuam et ipse filius est Belial ita ut nemo ei possit loqui
1SAM|25|18|festinavit igitur Abigail et tulit ducentos panes et duos utres vini et quinque arietes coctos et quinque sata pulentae et centum ligaturas uvae passae et ducentas massas caricarum et inposuit super asinos
1SAM|25|19|dixitque pueris suis praecedite me ecce ego post tergum sequar vos viro autem suo Nabal non indicavit
1SAM|25|20|cum ergo ascendisset asinum et descenderet ad radices montis David et viri eius descendebant in occursum eius quibus et illa occurrit
1SAM|25|21|et ait David vere frustra servavi omnia quae huius erant in deserto et non periit quicquam de cunctis quae ad eum pertinebant et reddidit mihi malum pro bono
1SAM|25|22|haec faciat Deus inimicis David et haec addat si reliquero de omnibus quae ad eum pertinent usque mane mingentem ad parietem
1SAM|25|23|cum autem vidisset Abigail David festinavit et descendit de asino et procidit coram David super faciem suam et adoravit super terram
1SAM|25|24|et cecidit ad pedes eius et dixit in me sit domine mi haec iniquitas loquatur obsecro ancilla tua in auribus tuis et audi verba famulae tuae
1SAM|25|25|ne ponat oro dominus meus rex cor suum super virum istum iniquum Nabal quia secundum nomen suum stultus est et est stultitia cum eo ego autem ancilla tua non vidi pueros tuos domine mi quos misisti
1SAM|25|26|nunc ergo domine mi vivit Dominus et vivit anima tua qui prohibuit te ne venires in sanguine et salvavit manum tuam tibi et nunc fiant sicut Nabal inimici tui et qui quaerunt domino meo malum
1SAM|25|27|quapropter suscipe benedictionem hanc quam adtulit ancilla tua tibi domino meo et da pueris qui sequuntur te dominum meum
1SAM|25|28|aufer iniquitatem famulae tuae faciens enim faciet tibi Dominus domino meo domum fidelem quia proelia Domini domine mi tu proeliaris malitia ergo non inveniatur in te omnibus diebus vitae tuae
1SAM|25|29|si enim surrexerit aliquando homo persequens te et quaerens animam tuam erit anima domini mei custodita quasi in fasciculo viventium apud Dominum Deum tuum porro anima inimicorum tuorum rotabitur quasi in impetu et circulo fundae
1SAM|25|30|cum ergo fecerit tibi Dominus domino meo omnia quae locutus est bona de te et constituerit te ducem super Israhel
1SAM|25|31|non erit tibi hoc in singultum et in scrupulum cordis domino meo quod effuderis sanguinem innoxium aut ipse te ultus fueris et cum benefecerit Dominus domino meo recordaberis ancillae tuae
1SAM|25|32|et ait David ad Abigail benedictus Dominus Deus Israhel qui misit te hodie in occursum meum et benedictum eloquium tuum
1SAM|25|33|et benedicta tu quae prohibuisti me hodie ne irem ad sanguinem et ulciscerer me manu mea
1SAM|25|34|alioquin vivit Dominus Deus Israhel qui prohibuit me malum facere tibi nisi cito venisses in occursum mihi non remansisset Nabal usque ad lucem matutinam mingens ad parietem
1SAM|25|35|suscepit ergo David de manu eius omnia quae adtulerat ei dixitque ei vade pacifice in domum tuam ecce audivi vocem tuam et honoravi faciem tuam
1SAM|25|36|venit autem Abigail ad Nabal et ecce erat ei convivium in domo eius quasi convivium regis et cor Nabal iucundum erat enim ebrius nimis et non indicavit ei verbum pusillum aut grande usque in mane
1SAM|25|37|diluculo autem cum digessisset vinum Nabal indicavit ei uxor sua verba haec et emortuum est cor eius intrinsecus et factus est quasi lapis
1SAM|25|38|cumque pertransissent decem dies percussit Dominus Nabal et mortuus est
1SAM|25|39|quod cum audisset David mortuum Nabal ait benedictus Dominus qui iudicavit causam obprobrii mei de manu Nabal et servum suum custodivit a malo et malitiam Nabal reddidit Dominus in caput eius misit ergo David et locutus est ad Abigail ut sumeret eam sibi in uxorem
1SAM|25|40|et venerunt pueri David ad Abigail in Carmelum et locuti sunt ad eam dicentes David misit nos ad te ut accipiat te sibi in uxorem
1SAM|25|41|quae consurgens adoravit prona in terram et ait ecce famula tua sit in ancillam ut lavet pedes servorum domini mei
1SAM|25|42|et festinavit et surrexit Abigail et ascendit super asinum et quinque puellae ierunt cum ea pedisequae eius et secuta est nuntios David et facta est illi uxor
1SAM|25|43|sed et Ahinoem accepit David de Iezrahel et fuit utraque uxor eius
1SAM|25|44|Saul autem dedit Michol filiam suam uxorem David Falti filio Lais qui erat de Gallim
1SAM|26|1|et venerunt Ziphei ad Saul in Gabaa dicentes ecce David absconditus est in colle Achilae quae est ex adverso solitudinis
1SAM|26|2|et surrexit Saul et descendit in desertum Ziph et cum eo tria milia virorum de electis Israhel ut quaereret David in deserto Ziph
1SAM|26|3|et castrametatus est Saul in Gabaa Achilae quae erat ex adverso solitudinis in via David autem habitabat in deserto videns autem quod venisset Saul post se in desertum
1SAM|26|4|misit exploratores et didicit quod venisset certissime
1SAM|26|5|et surrexit David et venit ad locum ubi erat Saul cumque vidisset locum in quo dormiebat Saul et Abner filius Ner princeps militiae eius Saulem dormientem in tentorio et reliquum vulgus per circuitum eius
1SAM|26|6|ait David ad Ahimelech Cettheum et Abisai filium Sarviae fratrem Ioab dicens quis descendet mecum ad Saul in castra dixitque Abisai ego descendam tecum
1SAM|26|7|venerunt ergo David et Abisai ad populum nocte et invenerunt Saul iacentem et dormientem in tentorio et hastam fixam in terra ad caput eius Abner autem et populum dormientes in circuitu eius
1SAM|26|8|dixitque Abisai ad David conclusit Deus hodie inimicum tuum in manus tuas nunc ergo perfodiam eum lancea in terra semel et secundo opus non erit
1SAM|26|9|et dixit David ad Abisai ne interficias eum quis enim extendit manum suam in christum Domini et innocens erit
1SAM|26|10|et dixit David vivit Dominus quia nisi Dominus percusserit eum aut dies eius venerit ut moriatur aut in proelium descendens perierit
1SAM|26|11|propitius mihi sit Dominus ne extendam manum meam in christum Domini nunc igitur tolle hastam quae est ad caput eius et scyphum aquae et abeamus
1SAM|26|12|tulit ergo David hastam et scyphum aquae qui erat ad caput Saul et abierunt et non erat quisquam qui videret et intellegeret et vigilaret sed omnes dormiebant quia sopor Domini inruerat super eos
1SAM|26|13|cumque transisset David ex adverso et stetisset in vertice montis de longe et esset grande intervallum inter eos
1SAM|26|14|clamavit David ad populum et ad Abner filium Ner dicens nonne respondebis Abner et respondens Abner ait quis es tu qui clamas et inquietas regem
1SAM|26|15|et ait David ad Abner numquid non vir tu es et quis alius similis tui in Israhel quare ergo non custodisti dominum tuum regem ingressus est enim unus de turba ut interficeret regem dominum tuum
1SAM|26|16|non est bonum hoc quod fecisti vivit Dominus quoniam filii mortis estis vos qui non custodistis dominum vestrum christum Domini nunc ergo vide ubi sit hasta regis et ubi scyphus aquae qui erat ad caput eius
1SAM|26|17|cognovit autem Saul vocem David et dixit num vox tua est haec fili mi David et David vox mea domine mi rex
1SAM|26|18|et ait quam ob causam dominus meus persequitur servum suum quid feci aut quod est in manu mea malum
1SAM|26|19|nunc ergo audi oro domine mi rex verba servi tui si Dominus incitat te adversum me odoretur sacrificium si autem filii hominum maledicti sunt in conspectu Domini qui eiecerunt me hodie ut non habitem in hereditate Domini dicentes vade servi diis alienis
1SAM|26|20|et nunc non effundatur sanguis meus in terra coram Domino quia egressus est rex Israhel ut quaerat pulicem unum sicut persequitur perdix in montibus
1SAM|26|21|et ait Saul peccavi revertere fili mi David nequaquam enim ultra male tibi faciam eo quod pretiosa fuerit anima mea in oculis tuis hodie apparet quod stulte egerim et ignoraverim multa nimis
1SAM|26|22|et respondens David ait ecce hasta regis transeat unus de pueris et tollat eam
1SAM|26|23|Dominus autem retribuet unicuique secundum iustitiam suam et fidem tradidit enim te Dominus hodie in manu mea et nolui levare manum meam in christum Domini
1SAM|26|24|et sicuti magnificata est anima tua hodie in oculis meis sic magnificetur anima mea in oculis Domini et liberet me de omni angustia
1SAM|26|25|ait ergo Saul ad David benedictus tu fili mi David et quidem faciens facies et potens poteris abiit autem David in viam suam et Saul reversus est in locum suum
1SAM|27|1|et ait David in corde suo aliquando incidam in uno die in manu Saul nonne melius est ut fugiam et salver in terra Philisthinorum ut desperet Saul cessetque me quaerere in cunctis finibus Israhel fugiam ergo manus eius
1SAM|27|2|et surrexit David et abiit ipse et sescenti viri cum eo ad Achis filium Mahoc regem Geth
1SAM|27|3|et habitavit David cum Achis in Geth ipse et viri eius vir et domus eius David et duae uxores eius Ahinoem Iezrahelites et Abigail uxor Nabal Carmeli
1SAM|27|4|et nuntiatum est Saul quod fugisset David in Geth et non addidit ultra ut quaereret eum
1SAM|27|5|dixit autem David ad Achis si inveni gratiam in oculis tuis detur mihi locus in una urbium regionis huius ut habitem ibi cur enim manet servus tuus in civitate regis tecum
1SAM|27|6|dedit itaque ei Achis in die illa Siceleg propter quam causam facta est Siceleg regum Iuda usque in diem hanc
1SAM|27|7|fuit autem numerus dierum quibus habitavit David in regione Philisthinorum quattuor mensuum
1SAM|27|8|et ascendit David et viri eius et agebant praedas de Gesuri et de Gedri et de Amalechitis hii enim pagi habitabantur in terra antiquitus euntibus Sur usque ad terram Aegypti
1SAM|27|9|et percutiebat David omnem terram nec relinquebat viventem virum et mulierem tollensque oves et boves et asinos et camelos et vestes revertebatur et veniebat ad Achis
1SAM|27|10|dicebat autem ei Achis in quem inruisti hodie respondebatque David contra meridiem Iudae et contra meridiem Hiramel et contra meridiem Ceni
1SAM|27|11|virum et mulierem non vivificabat David nec adducebat in Geth dicens ne forte loquantur adversum nos haec fecit David et hoc erat decretum illi omnibus diebus quibus habitavit in regione Philisthinorum
1SAM|27|12|credidit ergo Achis David dicens multa mala operatus est contra populum suum Israhel erit igitur mihi servus sempiternus
1SAM|28|1|factum est autem in diebus illis congregaverunt Philisthim agmina sua ut praepararentur ad bellum contra Israhel dixitque Achis ad David sciens nunc scito quoniam mecum egredieris in castris tu et viri tui
1SAM|28|2|dixitque David ad Achis nunc scies quae facturus est servus tuus et ait Achis ad David et ego custodem capitis mei ponam te cunctis diebus
1SAM|28|3|Samuhel autem mortuus est planxitque eum omnis Israhel et sepelierunt eum in Rama urbe sua et Saul abstulit magos et ariolos de terra
1SAM|28|4|congregatique sunt Philisthim et venerunt et castrametati sunt in Sunam congregavit autem et Saul universum Israhel et venit in Gelboe
1SAM|28|5|et vidit Saul castra Philisthim et timuit et expavit cor eius nimis
1SAM|28|6|consuluitque Dominum et non respondit ei neque per somnia neque per sacerdotes neque per prophetas
1SAM|28|7|dixitque Saul servis suis quaerite mihi mulierem habentem pythonem et vadam ad eam et sciscitabor per illam et dixerunt servi eius ad eum est mulier habens pythonem in Aendor
1SAM|28|8|mutavit ergo habitum suum vestitusque est aliis vestimentis abiit ipse et duo viri cum eo veneruntque ad mulierem nocte et ait divina mihi in pythone et suscita mihi quem dixero tibi
1SAM|28|9|et ait mulier ad eum ecce tu nosti quanta fecerit Saul et quomodo eraserit magos et ariolos de terra quare ergo insidiaris animae meae ut occidar
1SAM|28|10|et iuravit ei Saul in Domino dicens vivit Dominus quia non veniet tibi quicquam mali propter hanc rem
1SAM|28|11|dixitque ei mulier quem suscitabo tibi qui ait Samuhelem suscita mihi
1SAM|28|12|cum autem vidisset mulier Samuhelem exclamavit voce magna et dixit ad Saul quare inposuisti mihi tu es enim Saul
1SAM|28|13|dixitque ei rex noli timere quid vidisti et ait mulier ad Saul deos vidi ascendentes de terra
1SAM|28|14|dixitque ei qualis est forma eius quae ait vir senex ascendit et ipse amictus est pallio intellexit Saul quod Samuhel esset et inclinavit se super faciem suam in terra et adoravit
1SAM|28|15|dixit autem Samuhel ad Saul quare inquietasti me ut suscitarer et ait Saul coartor nimis siquidem Philisthim pugnant adversum me et Deus recessit a me et exaudire me noluit neque in manu prophetarum neque per somnia vocavi ergo te ut ostenderes mihi quid faciam
1SAM|28|16|et ait Samuhel quid interrogas me cum Dominus recesserit a te et transierit ad aemulum tuum
1SAM|28|17|faciet enim Dominus tibi sicut locutus est in manu mea et scindet regnum de manu tua et dabit illud proximo tuo David
1SAM|28|18|quia non oboedisti voci Domini neque fecisti iram furoris eius in Amalech idcirco quod pateris fecit tibi Dominus hodie
1SAM|28|19|et dabit Dominus etiam Israhel tecum in manu Philisthim cras autem tu et filii tui mecum eritis sed et castra Israhel tradet Dominus in manu Philisthim
1SAM|28|20|statimque Saul cecidit porrectus in terram extimuerat enim verba Samuhel et robur non erat in eo quia non comederat panem tota die illa
1SAM|28|21|ingressa est itaque mulier ad Saul et ait conturbatus enim erat valde dixitque ad eum ecce oboedivit ancilla tua voci tuae et posui animam meam in manu mea et audivi sermones tuos quos locutus es ad me
1SAM|28|22|nunc igitur audi et tu vocem ancillae tuae ut ponam coram te buccellam panis et comedens convalescas ut possis iter facere
1SAM|28|23|qui rennuit et ait non comedam coegerunt autem eum servi sui et mulier et tandem audita voce eorum surrexit de terra et sedit super lectum
1SAM|28|24|mulier autem illa habebat vitulum pascualem in domo et festinavit et occidit eum tollensque farinam miscuit eam et coxit azyma
1SAM|28|25|et posuit ante Saul et ante servos eius qui cum comedissent surrexerunt et ambulaverunt per totam noctem illam
1SAM|29|1|congregata sunt ergo Philisthim universa agmina in Afec sed et Israhel castrametatus est super fontem qui erat in Iezrahel
1SAM|29|2|et satrapae quidem Philisthim incedebant in centuriis et milibus David autem et viri eius erant in novissimo agmine cum Achis
1SAM|29|3|dixeruntque principes Philisthim quid sibi volunt Hebraei isti et ait Achis ad principes Philisthim num ignoratis David qui fuit servus Saul regis Israhel et est apud me multis diebus vel annis et non inveni in eo quicquam ex die qua transfugit ad me usque ad diem hanc
1SAM|29|4|irati sunt autem adversus eum principes Philisthim et dixerunt ei revertatur vir et sedeat in loco suo in quo constituisti eum et non descendat nobiscum in proelium ne fiat nobis adversarius cum proeliari coeperimus quomodo enim aliter placare poterit dominum suum nisi in capitibus nostris
1SAM|29|5|nonne iste est David cui cantabant in choro dicentes percussit Saul in milibus suis et David in decem milibus suis
1SAM|29|6|vocavit ergo Achis David et ait ei vivit Dominus quia rectus es tu et bonus in conspectu meo et exitus tuus et introitus tuus mecum est in castris et non inveni in te quicquam mali ex die qua venisti ad me usque ad diem hanc sed satrapis non places
1SAM|29|7|revertere ergo et vade in pace et non offendes oculos satraparum Philisthim
1SAM|29|8|dixitque David ad Achis quid enim feci et quid invenisti in me servo tuo a die qua fui in conspectu tuo usque in diem hanc ut non veniam et pugnem contra inimicos domini mei regis
1SAM|29|9|respondens autem Achis locutus est ad David scio quia bonus es tu in oculis meis sicut angelus Dei sed principes Philisthim dixerunt non ascendet nobiscum in proelium
1SAM|29|10|igitur consurge mane tu et servi domini tui qui venerunt tecum et cum de nocte surrexeritis et coeperit dilucescere pergite
1SAM|29|11|surrexit itaque de nocte David ipse et viri eius ut proficiscerentur mane et reverterentur ad terram Philisthim Philisthim autem ascenderunt in Iezrahel
1SAM|30|1|cumque venissent David et viri eius in Siceleg die tertia Amalechitae impetum fecerant ex parte australi in Siceleg et percusserant Siceleg et succenderant eam igni
1SAM|30|2|et captivas duxerant mulieres ex ea et a minimo usque ad magnum et non interfecerant quemquam sed secum duxerant et pergebant in itinere suo
1SAM|30|3|cum ergo venisset David et viri eius ad civitatem et invenissent eam succensam igni et uxores suas et filios suos et filias ductas esse captivas
1SAM|30|4|levaverunt David et populus qui erat cum eo voces suas et planxerunt donec deficerent in eis lacrimae
1SAM|30|5|siquidem et duae uxores David captivae ductae fuerant Ahinoem Iezrahelites et Abigail uxor Nabal Carmeli
1SAM|30|6|et contristatus est David valde volebat enim eum populus lapidare quia amara erat anima uniuscuiusque viri super filiis suis et filiabus confortatus est autem David in Domino Deo suo
1SAM|30|7|et ait ad Abiathar sacerdotem filium Ahimelech adplica ad me ephod et adplicuit Abiathar ephod ad David
1SAM|30|8|et consuluit David Dominum dicens persequar an non latrunculos hos et conprehendam eos dixitque ei persequere absque dubio enim conprehendes eos et excuties praedam
1SAM|30|9|abiit ergo David ipse et sescenti viri qui erant cum eo et venerunt usque ad torrentem Besor et lassi quidam substiterunt
1SAM|30|10|persecutus est autem David ipse et quadringenti viri substiterant enim ducenti qui lassi transire non poterant torrentem Besor
1SAM|30|11|et invenerunt virum aegyptium in agro et adduxerunt eum ad David dederuntque ei panem ut comederet et ut biberet aquam
1SAM|30|12|sed et fragmen massae caricarum et duas ligaturas uvae passae quae cum comedisset reversus est spiritus eius et refocilatus est non enim comederat panem neque biberat aquam tribus diebus et tribus noctibus
1SAM|30|13|dixit itaque ei David cuius es tu vel unde quo pergis qui ait ei puer aegyptius ego sum servus viri amalechitae dereliquit autem me dominus meus quia aegrotare coepi nudius tertius
1SAM|30|14|siquidem nos erupimus ad australem partem Cerethi et contra Iudam et ad meridiem Chaleb et Siceleg succendimus igni
1SAM|30|15|dixitque ei David potes me ducere ad istum cuneum qui ait iura mihi per Deum quod non occidas me et non tradas me in manu domini mei et ducam te ad cuneum istum
1SAM|30|16|qui cum duxisset eum ecce illi discumbebant super faciem universae terrae comedentes et bibentes et quasi festum celebrantes diem pro cuncta praeda et spoliis quae ceperant de terra Philisthim et de terra Iuda
1SAM|30|17|et percussit eos David a vespere usque ad vesperam alterius diei et non evasit ex eis quisquam nisi quadringenti viri adulescentes qui ascenderant camelos et fugerant
1SAM|30|18|eruit ergo David omnia quae tulerant Amalechitae et duas uxores suas eruit
1SAM|30|19|nec defuit quicquam a parvo usque ad magnum tam de filiis quam de filiabus et de spoliis et quaecumque rapuerant omnia reduxit David
1SAM|30|20|et tulit universos greges et armenta et minavit ante faciem suam dixeruntque haec est praeda David
1SAM|30|21|venit autem David ad ducentos viros qui lassi substiterant nec sequi potuerant David et residere eos iusserat in torrente Besor qui egressi sunt obviam David et populo qui erat cum eo accedens autem David ad populum salutavit eos pacifice
1SAM|30|22|respondensque omnis vir pessimus et iniquus de viris qui ierant cum David dixit quia non venerunt nobiscum non dabimus eis quicquam de praeda quam eruimus sed sufficiat unicuique uxor sua et filii quos cum acceperint recedant
1SAM|30|23|dixit autem David non sic facietis fratres mei de his quae tradidit Dominus nobis et custodivit nos et dedit latrunculos qui eruperant adversum nos in manu nostra
1SAM|30|24|nec audiet vos quisquam super sermone hoc aequa enim pars erit descendentis ad proelium et remanentis ad sarcinas et similiter divident
1SAM|30|25|et factum est hoc ex die illa et deinceps constitutum et praefinitum et quasi lex in Israhel usque ad diem hanc
1SAM|30|26|venit ergo David in Siceleg et misit dona de praeda senioribus Iuda proximis suis dicens accipite benedictionem de praeda hostium Domini
1SAM|30|27|his qui erant in Bethel et qui in Ramoth ad meridiem et qui in Iether
1SAM|30|28|et qui in Aroer et qui in Sefamoth et qui in Esthama
1SAM|30|29|et qui in Rachal et qui in urbibus Ierameli et qui in urbibus Ceni
1SAM|30|30|et qui in Arama et qui in lacu Asan et qui in Athac
1SAM|30|31|et qui in Hebron et reliquis qui erant in his locis in quibus commoratus fuerat David ipse et viri eius
1SAM|31|1|Philisthim autem pugnabant adversum Israhel et fugerunt viri Israhel ante faciem Philisthim et ceciderunt interfecti in monte Gelboe
1SAM|31|2|inrueruntque Philisthim in Saul et filios eius et percusserunt Ionathan et Abinadab et Melchisue filios Saul
1SAM|31|3|totumque pondus proelii versum est in Saul et consecuti sunt eum viri sagittarii et vulneratus est vehementer a sagittariis
1SAM|31|4|dixitque Saul ad armigerum suum evagina gladium tuum et percute me ne forte veniant incircumcisi isti et interficiant me inludentes mihi et noluit armiger eius fuerat enim nimio timore perterritus arripuit itaque Saul gladium et inruit super eum
1SAM|31|5|quod cum vidisset armiger eius videlicet quod mortuus esset Saul inruit etiam ipse super gladium suum et mortuus est cum eo
1SAM|31|6|mortuus est ergo Saul et tres filii eius et armiger illius et universi viri eius in die illa pariter
1SAM|31|7|videntes autem viri Israhel qui erant trans vallem et trans Iordanem quod fugissent viri israhelitae et quod mortuus esset Saul et filii eius reliquerunt civitates suas et fugerunt veneruntque Philisthim et habitaverunt ibi
1SAM|31|8|facta autem die altera venerunt Philisthim ut spoliarent interfectos et invenerunt Saul et tres filios eius iacentes in monte Gelboe
1SAM|31|9|et praeciderunt caput Saul et expoliaverunt eum armis et miserunt in terram Philisthinorum per circuitum ut adnuntiaretur in templo idolorum et in populis
1SAM|31|10|et posuerunt arma eius in templo Astharoth corpus vero eius suspenderunt in muro Bethsan
1SAM|31|11|quod cum audissent habitatores Iabesgalaad quaecumque fecerant Philisthim Saul
1SAM|31|12|surrexerunt omnes viri fortissimi et ambulaverunt tota nocte et tulerunt cadaver Saul et cadavera filiorum eius de muro Bethsan veneruntque Iabes et conbuserunt ea ibi
1SAM|31|13|et tulerunt ossa eorum et sepelierunt in nemore Iabes et ieiunaverunt septem diebus
2SAM|1|1|factum est autem postquam mortuus est Saul ut David reverteretur a caede Amalech et maneret in Siceleg dies duos
2SAM|1|2|in die autem tertia apparuit homo veniens de castris Saul veste conscissa et pulvere aspersus caput et ut venit ad David cecidit super faciem suam et adoravit
2SAM|1|3|dixitque ad eum David unde venis qui ait ad eum de castris Israhel fugi
2SAM|1|4|et dixit ad eum David quod est verbum quod factum est indica mihi qui ait fugit populus e proelio et multi corruentes e populo mortui sunt sed et Saul et Ionathan filius eius interierunt
2SAM|1|5|dixitque David ad adulescentem qui nuntiabat unde scis quia mortuus est Saul et Ionathan filius eius
2SAM|1|6|ait adulescens qui narrabat ei casu veni in montem Gelboe et Saul incumbebat super hastam suam porro currus et equites adpropinquabant ei
2SAM|1|7|et conversus post tergum suum vidensque me vocavit cui cum respondissem adsum
2SAM|1|8|dixit mihi quisnam es tu et aio ad eum Amalechites sum
2SAM|1|9|et locutus est mihi sta super me et interfice me quoniam tenent me angustiae et adhuc tota anima in me est
2SAM|1|10|stansque super eum occidi illum sciebam enim quod vivere non poterat post ruinam et tuli diadema quod erat in capite eius et armillam de brachio illius et adtuli ad te dominum meum huc
2SAM|1|11|adprehendens autem David vestimenta sua scidit omnesque viri qui erant cum eo
2SAM|1|12|et planxerunt et fleverunt et ieiunaverunt usque ad vesperam super Saul et super Ionathan filium eius et super populum Domini et super domum Israhel quod corruissent gladio
2SAM|1|13|dixitque David ad iuvenem qui nuntiaverat ei unde es qui respondit filius hominis advenae amalechitae ego sum
2SAM|1|14|et ait ad eum David quare non timuisti mittere manum tuam ut occideres christum Domini
2SAM|1|15|vocansque David unum de pueris ait accedens inrue in eum qui percussit illum et mortuus est
2SAM|1|16|et ait ad eum David sanguis tuus super caput tuum os enim tuum locutum est adversum te dicens ego interfeci christum Domini
2SAM|1|17|planxit autem David planctum huiuscemodi super Saul et super Ionathan filium eius
2SAM|1|18|et praecepit ut docerent filios Iuda arcum sicut scriptum est in libro Iustorum
2SAM|1|19|incliti Israhel super montes tuos interfecti sunt quomodo ceciderunt fortes
2SAM|1|20|nolite adnuntiare in Geth neque adnuntietis in conpetis Ascalonis ne forte laetentur filiae Philisthim ne exultent filiae incircumcisorum
2SAM|1|21|montes Gelboe nec ros nec pluviae veniant super vos neque sint agri primitiarum quia ibi abiectus est clypeus fortium clypeus Saul quasi non esset unctus oleo
2SAM|1|22|a sanguine interfectorum ab adipe fortium sagitta Ionathan numquam rediit retrorsum et gladius Saul non est reversus inanis
2SAM|1|23|Saul et Ionathan amabiles et decori in vita sua in morte quoque non sunt divisi aquilis velociores leonibus fortiores
2SAM|1|24|filiae Israhel super Saul flete qui vestiebat vos coccino in deliciis qui praebebat ornamenta aurea cultui vestro
2SAM|1|25|quomodo ceciderunt fortes in proelio Ionathan in excelsis tuis occisus est
2SAM|1|26|doleo super te frater mi Ionathan decore nimis et amabilis super amorem mulierum
2SAM|1|27|quomodo ceciderunt robusti et perierunt arma bellica
2SAM|2|1|igitur post haec consuluit David Dominum dicens num ascendam in unam de civitatibus Iuda et ait Dominus ad eum ascende dixitque David quo ascendam et respondit ei in Hebron
2SAM|2|2|ascendit ergo David et duae uxores eius Ahinoem Iezrahelites et Abigail uxor Nabal Carmeli
2SAM|2|3|sed et viros qui erant cum eo duxit David singulos cum domo sua et manserunt in oppidis Hebron
2SAM|2|4|veneruntque viri Iuda et unxerunt ibi David ut regnaret super domum Iuda et nuntiatum est David quod viri Iabesgalaad sepelissent Saul
2SAM|2|5|misit ergo David nuntios ad viros Iabesgalaad dixitque ad eos benedicti vos Domino qui fecistis misericordiam hanc cum domino vestro Saul et sepelistis eum
2SAM|2|6|et nunc retribuet quidem vobis Dominus misericordiam et veritatem sed et ego reddam gratiam eo quod feceritis verbum istud
2SAM|2|7|confortentur manus vestrae et estote filii fortitudinis licet enim mortuus sit dominus vester Saul tamen me unxit domus Iuda regem sibi
2SAM|2|8|Abner autem filius Ner princeps exercitus Saul tulit Hisboseth filium Saul et circumduxit eum per Castra
2SAM|2|9|regemque constituit super Galaad et super Gesuri et super Iezrahel et super Ephraim et super Beniamin et super Israhel universum
2SAM|2|10|quadraginta annorum erat Hisboseth filius Saul cum regnare coepisset super Israhel et duobus annis regnavit sola autem domus Iuda sequebatur David
2SAM|2|11|et fuit numerus dierum quos commoratus est David imperans in Hebron super domum Iuda septem annorum et sex mensuum
2SAM|2|12|egressusque Abner filius Ner et pueri Hisboseth filii Saul de Castris in Gabaon
2SAM|2|13|porro Ioab filius Sarviae et pueri David egressi sunt et occurrerunt eis iuxta piscinam Gabaon et cum in unum convenissent e regione sederunt hii ex una parte piscinae et illi ex altera
2SAM|2|14|dixitque Abner ad Ioab surgant pueri et ludant coram nobis et respondit Ioab surgant
2SAM|2|15|surrexerunt ergo et transierunt numero duodecim de Beniamin ex parte Hisboseth filii Saul et duodecim de pueris David
2SAM|2|16|adprehensoque unusquisque capite conparis sui defixit gladium in latus contrarii et ceciderunt simul vocatumque est nomen loci illius ager Robustorum in Gabaon
2SAM|2|17|et ortum est bellum durum satis in die illa fugatusque est Abner et viri Israhel a pueris David
2SAM|2|18|erant autem ibi tres filii Sarviae Ioab et Abisai et Asahel porro Asahel cursor velocissimus fuit quasi unus ex capreis quae morantur in silvis
2SAM|2|19|persequebatur autem Asahel Abner et non declinavit ad dexteram sive ad sinistram omittens persequi Abner
2SAM|2|20|respexit itaque Abner post tergum suum et ait tune es Asahel qui respondit ego sum
2SAM|2|21|dixitque ei Abner vade ad dextram sive ad sinistram et adprehende unum de adulescentibus et tolle tibi spolia eius noluit autem Asahel omittere quin urgueret eum
2SAM|2|22|rursumque locutus est Abner ad Asahel recede noli me sequi ne conpellar confodere te in terra et levare non potero faciem meam ad Ioab fratrem tuum
2SAM|2|23|qui audire contempsit et noluit declinare percussit ergo eum Abner aversa hasta in inguine et transfodit et mortuus est in eodem loco omnesque qui transiebant per locum in quo ceciderat Asahel et mortuus erat subsistebant
2SAM|2|24|persequentibus autem Ioab et Abisai fugientem Abner sol occubuit et venerunt usque ad collem Aquaeductus qui est ex adverso vallis et itineris deserti in Gabaon
2SAM|2|25|congregatique sunt filii Beniamin ad Abner et conglobati in unum cuneum steterunt in summitate tumuli unius
2SAM|2|26|et exclamavit Abner ad Ioab et ait num usque ad internicionem tuus mucro desaeviet an ignoras quod periculosa sit desperatio usquequo non dicis populo ut omittat persequi fratres suos
2SAM|2|27|et ait Ioab vivit Dominus si locutus fuisses mane recessisset populus persequens fratrem suum
2SAM|2|28|insonuit ergo Ioab bucina et stetit omnis exercitus nec persecuti sunt ultra Israhel neque iniere certamen
2SAM|2|29|Abner autem et viri eius abierunt per campestria tota nocte illa et transierunt Iordanem et lustrata omni Bethoron venerunt ad Castra
2SAM|2|30|porro Ioab reversus omisso Abner congregavit omnem populum et defuerunt de pueris David decem et novem viri excepto Asahele
2SAM|2|31|servi autem David percusserunt de Beniamin et de viris qui erant cum Abner trecentos sexaginta qui et mortui sunt
2SAM|2|32|tuleruntque Asahel et sepelierunt eum in sepulchro patris sui in Bethleem et ambulaverunt tota nocte Ioab et viri qui erant cum eo et in ipso crepusculo pervenerunt in Hebron
2SAM|3|1|facta est ergo longa concertatio inter domum Saul et inter domum David David proficiens et semper se ipso robustior domus autem Saul decrescens cotidie
2SAM|3|2|nati quoque sunt filii David in Hebron fuitque primogenitus eius Amnon de Ahinoem Iezrahelitide
2SAM|3|3|et post eum Chelaab de Abigail uxore Nabal Carmeli porro tertius Absalom filius Maacha filiae Tholomai regis Gessur
2SAM|3|4|quartus autem Adonias filius Aggith et quintus Safathia filius Abital
2SAM|3|5|sextus quoque Iethraam de Agla uxore David hii nati sunt David in Hebron
2SAM|3|6|cum ergo esset proelium inter domum Saul et domum David Abner filius Ner regebat domum Saul
2SAM|3|7|fuerat autem Sauli concubina nomine Respha filia Ahia dixitque Hisboseth ad Abner
2SAM|3|8|quare ingressus es ad concubinam patris mei qui iratus nimis propter verba Hisboseth ait numquid caput canis ego sum adversum Iuda hodie qui fecerim misericordiam super domum Saul patris tui et super fratres et proximos eius et non tradidi te in manu David et tu requisisti in me quod argueres pro muliere hodie
2SAM|3|9|haec faciat Deus Abner et haec addat ei nisi quomodo iuravit Dominus David sic faciam cum eo
2SAM|3|10|ut transferatur regnum de domo Saul et elevetur thronus David super Israhel et super Iudam a Dan usque Bersabee
2SAM|3|11|et non potuit respondere ei quicquam quia metuebat illum
2SAM|3|12|misit ergo Abner nuntios ad David pro se dicentes cuius est terra et loquerentur fac mecum amicitias et erit manus mea tecum et reducam ad te universum Israhel
2SAM|3|13|qui ait optime ego faciam tecum amicitias sed unam rem peto a te dicens non videbis faciem meam antequam adduxeris Michol filiam Saul et sic venies et videbis me
2SAM|3|14|misit autem David nuntios ad Hisboseth filium Saul dicens redde uxorem meam Michol quam despondi mihi centum praeputiis Philisthim
2SAM|3|15|misit ergo Hisboseth et tulit eam a viro suo Faltihel filio Lais
2SAM|3|16|sequebaturque eam vir suus plorans usque Baurim et dixit ad eum Abner vade revertere qui reversus est
2SAM|3|17|sermonem quoque intulit Abner ad seniores Israhel dicens tam heri quam nudius tertius quaerebatis David ut regnaret super vos
2SAM|3|18|nunc ergo facite quoniam Dominus locutus est ad David dicens in manu servi mei David salvabo populum meum Israhel de manu Philisthim et omnium inimicorum eius
2SAM|3|19|locutus est autem Abner etiam ad Beniamin et abiit ut loqueretur ad David in Hebron omnia quae placuerant Israhel et universo Beniamin
2SAM|3|20|venitque ad David in Hebron cum viginti viris et fecit David Abner et viris eius qui venerant cum eo convivium
2SAM|3|21|et dixit Abner ad David surgam ut congregem ad te dominum meum regem omnem Israhel et ineam tecum foedus et imperes omnibus sicut desiderat anima tua cum ergo deduxisset David Abner et ille isset in pace
2SAM|3|22|statim pueri David et Ioab venerunt caesis latronibus cum praeda magna nimis Abner autem non erat cum David in Hebron quia iam dimiserat eum et profectus fuerat in pace
2SAM|3|23|et Ioab et omnis exercitus qui erat cum eo postea venerant nuntiatum est itaque Ioab a narrantibus venit Abner filius Ner ad regem et dimisit eum et abiit in pace
2SAM|3|24|et ingressus est Ioab ad regem et ait quid fecisti ecce venit Abner ad te quare dimisisti eum et abiit et recessit
2SAM|3|25|ignoras Abner filium Ner quoniam ad hoc venit ut deciperet te et sciret exitum tuum et introitum tuum et nosset omnia quae agis
2SAM|3|26|egressus itaque Ioab a David misit nuntios post Abner et reduxit eum a cisterna Sira ignorante David
2SAM|3|27|cumque redisset Abner in Hebron seorsum abduxit eum Ioab ad medium portae ut loqueretur ei in dolo et percussit illum ibi in inguine et mortuus est in ultionem sanguinis Asahel fratris eius
2SAM|3|28|quod cum audisset David rem iam gestam ait mundus ego sum et regnum meum apud Dominum usque in sempiternum a sanguine Abner filii Ner
2SAM|3|29|et veniat super caput Ioab et super omnem domum patris eius nec deficiat de domo Ioab fluxum seminis sustinens et leprosus tenens fusum et cadens gladio et indigens pane
2SAM|3|30|igitur Ioab et Abisai frater eius interfecerunt Abner eo quod occidisset Asahel fratrem eorum in Gabaon in proelio
2SAM|3|31|dixit autem David ad Ioab et ad omnem populum qui erat cum eo scindite vestimenta vestra et accingimini saccis et plangite ante exequias Abner porro rex David sequebatur feretrum
2SAM|3|32|cumque sepelissent Abner in Hebron levavit rex vocem suam et flevit super tumulum Abner flevit autem et omnis populus
2SAM|3|33|plangensque rex Abner ait nequaquam ut mori solent ignavi mortuus est Abner
2SAM|3|34|manus tuae non sunt ligatae et pedes tui non sunt conpedibus adgravati sed sicut solent cadere coram filiis iniquitatis corruisti congeminansque omnis populus flevit super eum
2SAM|3|35|cumque venisset universa multitudo cibum capere cum David clara adhuc die iuravit David dicens haec faciat mihi Deus et haec addat si ante occasum solis gustavero panem vel aliud quicquam
2SAM|3|36|omnisque populus audivit et placuerunt eis cuncta quae fecit rex in conspectu totius populi
2SAM|3|37|et cognovit omne vulgus et universus Israhel in die illa quoniam non actum fuisset a rege ut occideretur Abner filius Ner
2SAM|3|38|dixit quoque rex ad servos suos num ignoratis quoniam princeps et maximus cecidit hodie in Israhel
2SAM|3|39|ego autem adhuc delicatus et unctus rex porro viri isti filii Sarviae duri mihi sunt retribuat Dominus facienti malum iuxta malitiam suam
2SAM|4|1|audivit autem filius Saul quod cecidisset Abner in Hebron et dissolutae sunt manus eius omnisque Israhel perturbatus est
2SAM|4|2|duo autem viri principes latronum erant filio Saul nomen uni Baana et nomen alteri Rechab filii Remmon Berothitae de filiis Beniamin siquidem et Beroth reputata est in Beniamin
2SAM|4|3|et fugerunt Berothitae in Getthaim fueruntque ibi advenae usque in tempus illud
2SAM|4|4|erat autem Ionathan filio Saul filius debilis pedibus quinquennis enim fuit quando venit nuntius de Saul et Ionathan ex Iezrahel tollens itaque eum nutrix sua fugit cumque festinaret ut fugeret cecidit et claudus effectus est habuitque vocabulum Mifiboseth
2SAM|4|5|venientes igitur filii Remmon Berothitae Rechab et Baana ingressi sunt fervente die domum Hisboseth qui dormiebat super stratum suum meridie
2SAM|4|6|ingressi sunt autem domum adsumentes spicas tritici et percusserunt eum in inguine Rechab et Baana frater eius et fugerunt
2SAM|4|7|cum autem ingressi fuissent domum ille dormiebat super lectulum suum in conclavi et percutientes interfecerunt eum sublatoque capite eius abierunt per viam deserti tota nocte
2SAM|4|8|et adtulerunt caput Hisboseth ad David in Hebron dixeruntque ad regem ecce caput Hisboseth filii Saul inimici tui qui quaerebat animam tuam et dedit Dominus domino meo regi ultiones hodie de Saul et de semine eius
2SAM|4|9|respondens autem David Rechab et Baana fratri eius filiis Remmon Berothei dixit ad eos vivit Dominus qui eruit animam meam de omni angustia
2SAM|4|10|quoniam eum qui adnuntiaverat mihi et dixerat mortuus est Saul qui putabat se prospera nuntiare tenui et occidi in Siceleg cui oportebat me dare mercedem pro nuntio
2SAM|4|11|quanto magis nunc cum homines impii interfecerint virum innoxium in domo sua super lectulum suum non quaeram sanguinem eius de manu vestra et auferam vos de terra
2SAM|4|12|praecepit itaque David pueris et interfecerunt eos praecidentesque manus et pedes eorum suspenderunt eos super piscinam in Hebron caput autem Hisboseth tulerunt et sepelierunt in sepulchro Abner in Hebron
2SAM|5|1|et venerunt universae tribus Israhel ad David in Hebron dicentes ecce nos os tuum et caro tua sumus
2SAM|5|2|sed et heri et nudius tertius cum esset Saul rex super nos tu eras educens et reducens Israhel dixit autem Dominus ad te tu pasces populum meum Israhel et tu eris dux super Israhel
2SAM|5|3|venerunt quoque et senes de Israhel ad regem in Hebron et percussit cum eis rex David foedus in Hebron coram Domino unxeruntque David in regem super Israhel
2SAM|5|4|filius triginta annorum erat David cum regnare coepisset et quadraginta annis regnavit
2SAM|5|5|in Hebron regnavit super Iudam septem annis et sex mensibus in Hierusalem autem regnavit triginta tribus annis super omnem Israhel et Iudam
2SAM|5|6|et abiit rex et omnes viri qui erant cum eo in Hierusalem ad Iebuseum habitatorem terrae dictumque est ad David ab eis non ingredieris huc nisi abstuleris caecos et claudos dicentes non ingredietur David huc
2SAM|5|7|cepit autem David arcem Sion haec est civitas David
2SAM|5|8|proposuerat enim in die illa praemium qui percussisset Iebuseum et tetigisset domatum fistulas et claudos et caecos odientes animam David idcirco dicitur in proverbio caecus et claudus non intrabunt templum
2SAM|5|9|habitavit autem David in arce et vocavit eam civitatem David et aedificavit per gyrum a Mello et intrinsecus
2SAM|5|10|et ingrediebatur proficiens atque succrescens et Dominus Deus exercituum erat cum eo
2SAM|5|11|misit quoque Hiram rex Tyri nuntios ad David et ligna cedrina et artifices lignorum artificesque lapidum ad parietes et aedificaverunt domum David
2SAM|5|12|et cognovit David quoniam confirmasset eum Dominus regem super Israhel et quoniam exaltasset regnum eius super populum suum Israhel
2SAM|5|13|accepit ergo adhuc concubinas et uxores de Hierusalem postquam venerat de Hebron natique sunt David et alii filii et filiae
2SAM|5|14|et haec nomina eorum qui nati sunt ei in Hierusalem Samua et Sobab et Nathan et Salomon
2SAM|5|15|et Ibaar et Helisua et Nepheg
2SAM|5|16|et Iafia et Helisama et Helida et Helifeleth
2SAM|5|17|audierunt vero Philisthim quod unxissent David regem super Israhel et ascenderunt universi ut quaererent David quod cum audisset David descendit in praesidium
2SAM|5|18|Philisthim autem venientes diffusi sunt in valle Raphaim
2SAM|5|19|et consuluit David Dominum dicens si ascendam ad Philisthim et si dabis eos in manu mea et dixit Dominus ad David ascende quia tradens dabo Philisthim in manu tua
2SAM|5|20|venit ergo David in Baalpharasim et percussit eos ibi et dixit divisit Dominus inimicos meos coram me sicut dividuntur aquae propterea vocatum est nomen loci illius Baalpharasim
2SAM|5|21|et reliquerunt ibi sculptilia sua quae tulit David et viri eius
2SAM|5|22|et addiderunt adhuc Philisthim ut ascenderent et diffusi sunt in valle Raphaim
2SAM|5|23|consuluit autem David Dominum qui respondit non ascendas sed gyra post tergum eorum et venies ad eos ex adverso pirorum
2SAM|5|24|et cum audieris sonitum gradientis in cacumine pirorum tunc inibis proelium quia tunc egredietur Dominus ante faciem tuam ut percutiat castra Philisthim
2SAM|5|25|fecit itaque David sicut ei praeceperat Dominus et percussit Philisthim de Gabee usque dum venias Gezer
2SAM|6|1|congregavit autem rursum David omnes electos ex Israhel triginta milia
2SAM|6|2|surrexitque et abiit et universus populus qui erat cum eo de viris Iuda ut adducerent arcam Dei super quam invocatum est nomen Domini exercituum sedentis in cherubin super eam
2SAM|6|3|et inposuerunt arcam Domini super plaustrum novum tuleruntque eam de domo Abinadab qui erat in Gabaa Oza autem et Haio filii Abinadab minabant plaustrum novum
2SAM|6|4|cumque tulissent eam de domo Abinadab qui erat in Gabaa custodiens arcam Dei Haio praecedebat arcam
2SAM|6|5|David autem et omnis Israhel ludebant coram Domino in omnibus lignis fabrefactis et citharis et lyris et tympanis et sistris et cymbalis
2SAM|6|6|postquam autem venerunt ad aream Nachon extendit manum Oza ad arcam Dei et tenuit eam quoniam calcitrabant boves
2SAM|6|7|iratusque est indignatione Dominus contra Ozam et percussit eum super temeritate qui mortuus est ibi iuxta arcam Dei
2SAM|6|8|contristatus autem est David eo quod percussisset Dominus Ozam et vocatum est nomen loci illius Percussio Oza usque in diem hanc
2SAM|6|9|et extimuit David Dominum in die illa dicens quomodo ingredietur ad me arca Domini
2SAM|6|10|et noluit devertere ad se arcam Domini in civitate David sed devertit eam in domo Obededom Getthei
2SAM|6|11|et habitavit arca Domini in domo Obededom Getthei tribus mensibus et benedixit Dominus Obededom et omnem domum eius
2SAM|6|12|nuntiatumque est regi David benedixit Dominus Obededom et omnia eius propter arcam Dei abiit ergo David et adduxit arcam Dei de domo Obededom in civitatem David cum gaudio
2SAM|6|13|cumque transcendissent qui portabant arcam Domini sex passus immolabat bovem et arietem
2SAM|6|14|et David saltabat totis viribus ante Dominum porro David erat accinctus ephod lineo
2SAM|6|15|et David et omnis domus Israhel ducebant arcam testamenti Domini in iubilo et in clangore bucinae
2SAM|6|16|cumque intrasset arca Domini civitatem David Michol filia Saul prospiciens per fenestram vidit regem David subsilientem atque saltantem coram Domino et despexit eum in corde suo
2SAM|6|17|et introduxerunt arcam Domini et posuerunt eam in loco suo in medio tabernaculi quod tetenderat ei David et obtulit David holocausta coram Domino et pacifica
2SAM|6|18|cumque conplesset offerens holocaustum et pacifica benedixit populo in nomine Domini exercituum
2SAM|6|19|et partitus est multitudini universae Israhel tam viro quam mulieri singulis collyridam panis unam et assaturam bubulae carnis unam et similam frixam oleo et abiit omnis populus unusquisque in domum suam
2SAM|6|20|reversusque est et David ut benediceret domui suae et egressa Michol filia Saul in occursum David ait quam gloriosus fuit hodie rex Israhel discoperiens se ante ancillas servorum suorum et nudatus est quasi si nudetur unus de scurris
2SAM|6|21|dixitque David ad Michol ante Dominum qui elegit me potius quam patrem tuum et quam omnem domum eius et praecepit mihi ut essem dux super populum Domini Israhel
2SAM|6|22|et ludam et vilior fiam plus quam factus sum et ero humilis in oculis meis et cum ancillis de quibus locuta es gloriosior apparebo
2SAM|6|23|igitur Michol filiae Saul non est natus filius usque ad diem mortis suae
2SAM|7|1|factum est autem cum sedisset rex in domo sua et Dominus dedisset ei requiem undique ab universis inimicis suis
2SAM|7|2|dixit ad Nathan prophetam videsne quod ego habitem in domo cedrina et arca Dei posita sit in medio pellium
2SAM|7|3|dixitque Nathan ad regem omne quod est in corde tuo vade fac quia Dominus tecum est
2SAM|7|4|factum est autem in nocte illa et ecce sermo Domini ad Nathan dicens
2SAM|7|5|vade et loquere ad servum meum David haec dicit Dominus numquid tu aedificabis mihi domum ad habitandum
2SAM|7|6|neque enim habitavi in domo ex die qua eduxi filios Israhel de terra Aegypti usque in diem hanc sed ambulans ambulabam in tabernaculo et in tentorio
2SAM|7|7|per cuncta loca quae transivi cum omnibus filiis Israhel numquid loquens locutus sum ad unam de tribubus Israhel cui praecepi ut pasceret populum meum Israhel dicens quare non aedificastis mihi domum cedrinam
2SAM|7|8|et nunc haec dices servo meo David haec dicit Dominus exercituum ego tuli te de pascuis sequentem greges ut esses dux super populum meum Israhel
2SAM|7|9|et fui tecum in omnibus ubicumque ambulasti et interfeci universos inimicos tuos a facie tua fecique tibi nomen grande iuxta nomen magnorum qui sunt in terra
2SAM|7|10|et ponam locum populo meo Israhel et plantabo eum et habitabit sub eo et non turbabitur amplius nec addent filii iniquitatis ut adfligant eum sicut prius
2SAM|7|11|ex die qua constitui iudices super populum meum Israhel et requiem dabo tibi ab omnibus inimicis tuis praedicitque tibi Dominus quod domum faciat tibi Dominus
2SAM|7|12|cumque conpleti fuerint dies tui et dormieris cum patribus tuis suscitabo semen tuum post te quod egredietur de utero tuo et firmabo regnum eius
2SAM|7|13|ipse aedificabit domum nomini meo et stabiliam thronum regni eius usque in sempiternum
2SAM|7|14|ego ero ei in patrem et ipse erit mihi in filium qui si inique aliquid gesserit arguam eum in virga virorum et in plagis filiorum hominum
2SAM|7|15|misericordiam autem meam non auferam ab eo sicut abstuli a Saul quem amovi a facie tua
2SAM|7|16|et fidelis erit domus tua et regnum tuum usque in aeternum ante faciem tuam et thronus tuus erit firmus iugiter
2SAM|7|17|secundum omnia verba haec et iuxta universam visionem istam sic locutus est Nathan ad David
2SAM|7|18|ingressus est autem rex David et sedit coram Domino et dixit quis ego sum Domine Deus et quae domus mea quia adduxisti me hucusque
2SAM|7|19|sed et hoc parum visum est in conspectu tuo Domine Deus nisi loquereris etiam de domo servi tui in longinquum ista est enim lex Adam Domine Deus
2SAM|7|20|quid ergo addere poterit adhuc David ut loquatur ad te tu enim scis servum tuum Domine Deus
2SAM|7|21|propter verbum tuum et secundum cor tuum fecisti omnia magnalia haec ita ut notum faceres servo tuo
2SAM|7|22|idcirco magnificatus es Domine Deus quia non est similis tui neque est deus extra te in omnibus quae audivimus auribus nostris
2SAM|7|23|quae est autem ut populus tuus Israhel gens in terra propter quam ivit Deus ut redimeret eam sibi in populum et poneret sibi nomen faceretque eis magnalia et horribilia super terram a facie populi tui quem redemisti tibi ex Aegypto gentem et deum eius
2SAM|7|24|et firmasti tibi populum tuum Israhel in populum sempiternum et tu Domine factus es eis in Deum
2SAM|7|25|nunc ergo Domine Deus verbum quod locutus es super servum tuum et super domum eius suscita in sempiternum et fac sicut locutus es
2SAM|7|26|et magnificetur nomen tuum usque in sempiternum atque dicatur Dominus exercituum Deus super Israhel et domus servi tui David erit stabilita coram Domino
2SAM|7|27|quia tu Domine exercituum Deus Israhel revelasti aurem servi tui dicens domum aedificabo tibi propterea invenit servus tuus cor suum ut oraret te oratione hac
2SAM|7|28|nunc ergo Domine Deus tu es Deus et verba tua erunt vera locutus es enim ad servum tuum bona haec
2SAM|7|29|incipe igitur et benedic domui servi tui ut sit in sempiternum coram te quia tu Domine Deus locutus es et benedictione tua benedicetur domus servi tui in sempiternum
2SAM|8|1|factum est autem post haec percussit David Philisthim et humiliavit eos et tulit David frenum tributi de manu Philisthim
2SAM|8|2|et percussit Moab et mensus est eos funiculo coaequans terrae mensus est autem duos funiculos unum ad occidendum et unum ad vivificandum factusque est Moab David serviens sub tributo
2SAM|8|3|et percussit David Adadezer filium Roob regem Soba quando profectus est ut dominaretur super flumen Eufraten
2SAM|8|4|et captis David ex parte eius mille septingentis equitibus et viginti milibus peditum subnervavit omnes iugales curruum dereliquit autem ex eis centum currus
2SAM|8|5|venit quoque Syria Damasci ut praesidium ferret Adadezer regi Soba et percussit David de Syria viginti duo milia virorum
2SAM|8|6|et posuit David praesidium in Syria Damasci factaque est Syria David serviens sub tributo servavit Dominus David in omnibus ad quaecumque profectus est
2SAM|8|7|et tulit David arma aurea quae habebant servi Adadezer et detulit ea in Hierusalem
2SAM|8|8|et de Bete et de Beroth civitatibus Adadezer tulit rex David aes multum nimis
2SAM|8|9|audivit autem Thou rex Emath quod percussisset David omne robur Adadezer
2SAM|8|10|et misit Thou Ioram filium suum ad regem David ut salutaret eum congratulans et gratias ageret eo quod expugnasset Adadezer et percussisset eum hostis quippe erat Thou Adadezer et in manu eius erant vasa argentea et vasa aurea et vasa aerea
2SAM|8|11|quae et ipsa sanctificavit rex David Domino cum argento et auro quae sanctificaverat de universis gentibus quas subegerat
2SAM|8|12|de Syria et Moab et filiis Ammon et Philisthim et Amalech et de manubiis Adadezer filii Roob regis Soba
2SAM|8|13|fecit quoque sibi David nomen cum reverteretur capta Syria in valle Salinarum caesis duodecim milibus
2SAM|8|14|et posuit in Idumea custodes statuitque praesidium et facta est universa Idumea serviens David et servavit Dominus David in omnibus ad quaecumque profectus est
2SAM|8|15|et regnavit David super omnem Israhel faciebat quoque David iudicium et iustitiam omni populo suo
2SAM|8|16|Ioab autem filius Sarviae erat super exercitum porro Iosaphat filius Ahilud erat a commentariis
2SAM|8|17|et Sadoc filius Achitob et Ahimelech filius Abiathar sacerdotes et Saraias scriba
2SAM|8|18|Banaias autem filius Ioiada super Cherethi et Felethi filii autem David sacerdotes erant
2SAM|9|1|et dixit David putasne est aliquis qui remanserit de domo Saul ut faciam cum eo misericordiam propter Ionathan
2SAM|9|2|erat autem de domo Saul servus nomine Siba quem cum vocasset rex ad se dixit ei tune es Siba et ille respondit ego sum servus tuus
2SAM|9|3|et ait rex num superest aliquis de domo Saul ut faciam cum eo misericordiam Dei dixitque Siba regi superest filius Ionathan debilis pedibus
2SAM|9|4|ubi inquit est et Siba ad regem ecce ait in domo est Machir filii Amihel in Lodabar
2SAM|9|5|misit ergo rex David et tulit eum de domo Machir filii Amihel de Lodabar
2SAM|9|6|cum autem venisset Mifiboseth filius Ionathan filii Saul ad David corruit in faciem suam et adoravit dixitque David Mifiboseth qui respondit adsum servus tuus
2SAM|9|7|et ait ei David ne timeas quia faciens faciam in te misericordiam propter Ionathan patrem tuum et restituam tibi omnes agros Saul patris tui et tu comedes panem in mensa mea semper
2SAM|9|8|qui adorans eum dixit quis ego sum servus tuus quoniam respexisti super canem mortuum similem mei
2SAM|9|9|vocavit itaque rex Sibam puerum Saul et dixit ei omnia quaecumque fuerunt Saul et universam domum eius dedi filio domini tui
2SAM|9|10|operare igitur ei terram tu et filii tui et servi tui et inferes filio domini tui cibos ut alatur Mifiboseth autem filius domini tui comedet semper panem super mensam meam erant autem Sibae quindecim filii et viginti servi
2SAM|9|11|dixitque Siba ad regem sicut iussisti domine mi rex servo tuo sic faciet servus tuus et Mifiboseth comedet super mensam tuam quasi unus de filiis regis
2SAM|9|12|habebat autem Mifiboseth filium parvulum nomine Micha omnis vero cognatio domus Siba serviebat Mifiboseth
2SAM|9|13|porro Mifiboseth habitabat in Hierusalem quia de mensa regis iugiter vescebatur et erat claudus utroque pede
2SAM|10|1|factum est autem post haec ut moreretur rex filiorum Ammon et regnaret Anon filius eius pro eo
2SAM|10|2|dixitque David faciam misericordiam cum Anon filio Naas sicut fecit pater eius mecum misericordiam misit ergo David consolans eum per servos suos super patris interitu cum autem venissent servi David in terram filiorum Ammon
2SAM|10|3|dixerunt principes filiorum Ammon ad Anon dominum suum putas quod propter honorem patris tui David miserit ad te consolatores et non ideo ut investigaret et exploraret civitatem et everteret eam misit David servos suos ad te
2SAM|10|4|tulit itaque Anon servos David rasitque dimidiam partem barbae eorum et praecidit vestes eorum medias usque ad nates et dimisit eos
2SAM|10|5|quod cum nuntiatum esset David misit in occursum eorum erant enim viri confusi turpiter valde et mandavit eis David manete Hiericho donec crescat barba vestra et tunc revertimini
2SAM|10|6|videntes autem filii Ammon quod iniuriam fecissent David miserunt et conduxerunt mercede Syrum Roob et Syrum Soba viginti milia peditum et a rege Maacha mille viros et ab Histob duodecim milia virorum
2SAM|10|7|quod cum audisset David misit Ioab et omnem exercitum bellatorum
2SAM|10|8|egressi sunt ergo filii Ammon et direxerunt aciem ante ipsum introitum portae Syrus autem Soba et Roob et Histob et Maacha seorsum erant in campo
2SAM|10|9|videns igitur Ioab quod praeparatum esset adversum se proelium et ex adverso et post tergum elegit ex omnibus electis Israhel et instruxit aciem contra Syrum
2SAM|10|10|reliquam autem partem populi tradidit Abisai fratri suo qui direxit aciem adversum filios Ammon
2SAM|10|11|et ait Ioab si praevaluerint adversum me Syri eris mihi in adiutorium si autem filii Ammon praevaluerint adversum te auxiliabor tibi
2SAM|10|12|esto vir fortis et pugnemus pro populo nostro et civitate Dei nostri Dominus autem faciet quod bonum est in conspectu suo
2SAM|10|13|iniit itaque Ioab et populus qui erat cum eo certamen contra Syros qui statim fugerunt a facie eius
2SAM|10|14|filii autem Ammon videntes quod fugissent Syri fugerunt et ipsi a facie Abisai et ingressi sunt civitatem reversusque est Ioab a filiis Ammon et venit Hierusalem
2SAM|10|15|videntes igitur Syri quoniam corruissent coram Israhel congregati sunt pariter
2SAM|10|16|misitque Adadezer et eduxit Syros qui erant trans Fluvium et adduxit exercitum eorum Sobach autem magister militiae Adadezer erat princeps eorum
2SAM|10|17|quod cum nuntiatum esset David contraxit omnem Israhelem et transivit Iordanem venitque in Helema et direxerunt aciem Syri ex adverso David et pugnaverunt contra eum
2SAM|10|18|fugeruntque Syri a facie Israhel et occidit David de Syris septingentos currus et quadraginta milia equitum et Sobach principem militiae percussit qui statim mortuus est
2SAM|10|19|videntes autem universi reges qui erant in praesidio Adadezer victos se ab Israhel fecerunt pacem cum Israhel et servierunt eis timueruntque Syri auxilium praebere filiis Ammon
2SAM|11|1|factum est ergo vertente anno eo tempore quo solent reges ad bella procedere misit David Ioab et servos suos cum eo et universum Israhel et vastaverunt filios Ammon et obsederunt Rabba David autem remansit in Hierusalem
2SAM|11|2|dum haec agerentur accidit ut surgeret David de stratu suo post meridiem et deambularet in solario domus regiae viditque mulierem se lavantem ex adverso super solarium suum erat autem mulier pulchra valde
2SAM|11|3|misit ergo rex et requisivit quae esset mulier nuntiatumque ei est quod ipsa esset Bethsabee filia Heliam uxor Uriae Hetthei
2SAM|11|4|missis itaque David nuntiis tulit eam quae cum ingressa esset ad illum dormivit cum ea statimque sanctificata est ab inmunditia sua
2SAM|11|5|et reversa est domum suam concepto fetu mittensque nuntiavit David et ait concepi
2SAM|11|6|misit autem David ad Ioab dicens mitte ad me Uriam Hettheum misitque Ioab Uriam ad David
2SAM|11|7|et venit Urias ad David quaesivitque David quam recte ageret Ioab et populus et quomodo administraretur bellum
2SAM|11|8|et dixit David ad Uriam vade in domum tuam et lava pedes tuos egressus est Urias de domo regis secutusque est eum cibus regius
2SAM|11|9|dormivit autem Urias ante portam domus regiae cum aliis servis domini sui et non descendit ad domum suam
2SAM|11|10|nuntiatumque est David a dicentibus non ivit Urias ad domum suam et ait David ad Uriam numquid non de via venisti quare non descendisti ad domum tuam
2SAM|11|11|et ait Urias ad David arca et Israhel et Iuda habitant in papilionibus et dominus meus Ioab et servi domini mei super faciem terrae manent et ego ingrediar domum meam ut comedam et bibam et dormiam cum uxore mea per salutem tuam et per salutem animae tuae quod non faciam rem hanc
2SAM|11|12|ait ergo David ad Uriam mane hic etiam hodie et cras dimittam te mansit Urias in Hierusalem die illa et altera
2SAM|11|13|et vocavit eum David ut comederet coram se et biberet et inebriavit eum qui egressus vespere dormivit in stratu suo cum servis domini sui et in domum suam non descendit
2SAM|11|14|factum est ergo mane et scripsit David epistulam ad Ioab misitque per manum Uriae
2SAM|11|15|scribens in epistula ponite Uriam ex adverso belli ubi fortissimum proelium est et derelinquite eum ut percussus intereat
2SAM|11|16|igitur cum Ioab obsideret urbem posuit Uriam in loco quo sciebat viros esse fortissimos
2SAM|11|17|egressique viri de civitate bellabant adversum Ioab et ceciderunt de populo servorum David et mortuus est etiam Urias Hettheus
2SAM|11|18|misit itaque Ioab et nuntiavit David omnia verba proelii
2SAM|11|19|praecepitque nuntio dicens cum conpleveris universos sermones belli ad regem
2SAM|11|20|si eum videris indignari et dixerit quare accessistis ad murum ut proeliaremini an ignorabatis quod multa desuper ex muro tela mittantur
2SAM|11|21|quis percussit Abimelech filium Hieroboseth nonne mulier misit super eum fragmen molae de muro et interfecit eum in Thebes quare iuxta murum accessistis dices etiam servus tuus Urias Hettheus occubuit
2SAM|11|22|abiit ergo nuntius et venit et narravit David omnia quae ei praeceperat Ioab
2SAM|11|23|et dixit nuntius ad David praevaluerunt adversum nos viri et egressi sunt ad nos in agrum nos autem facto impetu persecuti eos sumus usque ad portam civitatis
2SAM|11|24|et direxerunt iacula sagittarii ad servos tuos ex muro desuper mortuique sunt de servis regis quin etiam servus tuus Urias Hettheus mortuus est
2SAM|11|25|et dixit David ad nuntium haec dices Ioab non te frangat ista res varius enim eventus est proelii et nunc hunc nunc illum consumit gladius conforta bellatores tuos adversum urbem ut destruas eam et exhortare eos
2SAM|11|26|audivit autem uxor Uriae quod mortuus esset Urias vir suus et planxit eum
2SAM|11|27|transactoque luctu misit David et introduxit eam domum suam et facta est ei uxor peperitque ei filium et displicuit verbum hoc quod fecerat David coram Domino
2SAM|12|1|misit ergo Dominus Nathan ad David qui cum venisset ad eum dixit ei duo viri erant in civitate una unus dives et alter pauper
2SAM|12|2|dives habebat oves et boves plurimos valde
2SAM|12|3|pauper autem nihil habebat omnino praeter ovem unam parvulam quam emerat et nutrierat et quae creverat apud eum cum filiis eius simul de pane illius comedens et de calice eius bibens et in sinu illius dormiens eratque illi sicut filia
2SAM|12|4|cum autem peregrinus quidam venisset ad divitem parcens ille sumere de ovibus et de bubus suis ut exhiberet convivium peregrino illi qui venerat ad se tulit ovem viri pauperis et praeparavit cibos homini qui venerat ad se
2SAM|12|5|iratus autem indignatione David adversus hominem illum nimis dixit ad Nathan vivit Dominus quoniam filius mortis est vir qui fecit hoc
2SAM|12|6|ovem reddet in quadruplum eo quod fecerit verbum istud et non pepercerit
2SAM|12|7|dixit autem Nathan ad David tu es ille vir haec dicit Dominus Deus Israhel ego unxi te in regem super Israhel et ego erui te de manu Saul
2SAM|12|8|et dedi tibi domum domini tui et uxores domini tui in sinu tuo dedique tibi domum Israhel et Iuda et si parva sunt ista adiciam tibi multo maiora
2SAM|12|9|quare ergo contempsisti verbum Domini ut faceres malum in conspectu meo Uriam Hettheum percussisti gladio et uxorem illius accepisti uxorem et interfecisti eum gladio filiorum Ammon
2SAM|12|10|quam ob rem non recedet gladius de domo tua usque in sempiternum eo quod despexeris me et tuleris uxorem Uriae Hetthei ut esset uxor tua
2SAM|12|11|itaque haec dicit Dominus ecce ego suscitabo super te malum de domo tua et tollam uxores tuas in oculis tuis et dabo proximo tuo et dormiet cum uxoribus tuis in oculis solis huius
2SAM|12|12|tu enim fecisti abscondite ego vero faciam verbum istud in conspectu omnis Israhel et in conspectu solis
2SAM|12|13|et dixit David ad Nathan peccavi Domino dixitque Nathan ad David Dominus quoque transtulit peccatum tuum non morieris
2SAM|12|14|verumtamen quoniam blasphemare fecisti inimicos Domini propter verbum hoc filius qui natus est tibi morte morietur
2SAM|12|15|et reversus est Nathan domum suam percussitque Dominus parvulum quem pepererat uxor Uriae David et desperatus est
2SAM|12|16|deprecatusque est David Dominum pro parvulo et ieiunavit David ieiunio et ingressus seorsum iacuit super terram
2SAM|12|17|venerunt autem seniores domus eius cogentes eum ut surgeret de terra qui noluit neque comedit cum eis cibum
2SAM|12|18|accidit autem die septima ut moreretur infans timueruntque servi David nuntiare ei quod mortuus esset parvulus dixerunt enim ecce cum parvulus adhuc viveret loquebamur ad eum et non audiebat vocem nostram quanto magis si dixerimus mortuus est puer se adfliget
2SAM|12|19|cum ergo vidisset David servos suos musitantes intellexit quod mortuus esset infantulus dixitque ad servos suos num mortuus est puer qui responderunt ei mortuus est
2SAM|12|20|surrexit igitur David de terra et lotus unctusque est cumque mutasset vestem ingressus est domum Domini et adoravit et venit in domum suam petivitque ut ponerent ei panem et comedit
2SAM|12|21|dixerunt autem ei servi sui quis est sermo quem fecisti propter infantem cum adhuc viveret ieiunasti et flebas mortuo autem puero surrexisti et comedisti panem
2SAM|12|22|qui ait propter infantem dum adhuc viveret ieiunavi et flevi dicebam enim quis scit si forte donet eum mihi Dominus et vivet infans
2SAM|12|23|nunc autem quia mortuus est quare ieiuno numquid potero revocare eum amplius ego vadam magis ad eum ille vero non revertetur ad me
2SAM|12|24|et consolatus est David Bethsabee uxorem suam ingressusque ad eam dormivit cum ea quae genuit filium et vocavit nomen eius Salomon et Dominus dilexit eum
2SAM|12|25|misitque in manu Nathan prophetae et vocavit nomen eius Amabilis Domino eo quod diligeret eum Dominus
2SAM|12|26|igitur pugnabat Ioab contra Rabbath filiorum Ammon et expugnabat urbem regiam
2SAM|12|27|misitque Ioab nuntios ad David dicens dimicavi adversum Rabbath et capienda est urbs Aquarum
2SAM|12|28|nunc igitur congrega reliquam partem populi et obside civitatem et cape eam ne cum a me vastata fuerit urbs nomini meo adscribatur victoria
2SAM|12|29|congregavit itaque David omnem populum et profectus est adversum Rabbath cumque dimicasset cepit eam
2SAM|12|30|et tulit diadema regis eorum de capite eius pondo auri talentum habens gemmas pretiosissimas et inpositum est super caput David sed et praedam civitatis asportavit multam valde
2SAM|12|31|populum quoque eius adducens serravit et circumegit super eos ferrata carpenta divisitque cultris et transduxit in typo laterum sic fecit universis civitatibus filiorum Ammon et reversus est David et omnis exercitus Hierusalem
2SAM|13|1|factum est autem post haec ut Absalom filii David sororem speciosissimam vocabulo Thamar adamaret Amnon filius David
2SAM|13|2|et deperiret eam valde ita ut aegrotaret propter amorem eius quia cum esset virgo difficile ei videbatur ut quippiam inhoneste ageret cum ea
2SAM|13|3|erat autem Amnonis amicus nomine Ionadab filius Semaa fratris David vir prudens valde
2SAM|13|4|qui dixit ad eum quare sic adtenuaris macie fili regis per singulos dies cur non indicas mihi dixitque ei Amnon Thamar sororem Absalom fratris mei amo
2SAM|13|5|cui respondit Ionadab cuba super lectulum tuum et languorem simula cumque venerit pater tuus ut visitet te dic ei veniat oro Thamar soror mea ut det mihi cibum et faciat pulmentum ut comedam de manu eius
2SAM|13|6|accubuit itaque Amnon et quasi aegrotare coepit cumque venisset rex ad visitandum eum ait Amnon ad regem veniat obsecro Thamar soror mea ut faciat in oculis meis duas sorbitiunculas et cibum capiam de manu eius
2SAM|13|7|misit ergo David ad Thamar domum dicens veni in domum Amnon fratris tui et fac ei pulmentum
2SAM|13|8|venitque Thamar in domum Amnon fratris sui ille autem iacebat quae tollens farinam commiscuit et liquefaciens in oculis eius coxit sorbitiunculas
2SAM|13|9|tollensque quod coxerat effudit et posuit coram eo et noluit comedere dixitque Amnon eicite universos a me cumque eiecissent omnes
2SAM|13|10|dixit Amnon ad Thamar infer cibum in conclave ut vescar de manu tua tulit ergo Thamar sorbitiunculas quas fecerat et intulit ad Amnon fratrem suum in conclave
2SAM|13|11|cumque obtulisset ei cibum adprehendit eam et ait veni cuba mecum soror mea
2SAM|13|12|quae respondit ei noli frater mi noli opprimere me neque enim hoc fas est in Israhel noli facere stultitiam hanc
2SAM|13|13|et ego enim ferre non potero obprobrium meum et tu eris quasi unus de insipientibus in Israhel quin potius loquere ad regem et non negabit me tibi
2SAM|13|14|noluit autem adquiescere precibus eius sed praevalens viribus oppressit eam et cubavit cum illa
2SAM|13|15|et exosam eam habuit Amnon magno odio nimis ita ut maius esset odium quo oderat eam amore quo ante dilexerat dixitque ei Amnon surge vade
2SAM|13|16|quae respondit ei maius est hoc malum quod nunc agis adversum me quam quod ante fecisti expellens me et noluit audire eam
2SAM|13|17|sed vocato puero qui ministrabat ei dixit eice hanc a me foras et claude ostium post eam
2SAM|13|18|quae induta erat talari tunica huiuscemodi enim filiae regis virgines vestibus utebantur eiecit itaque eam minister illius foras clausitque fores post eam
2SAM|13|19|quae aspergens cinerem capiti suo scissa talari tunica inpositisque manibus super caput suum ibat ingrediens et clamans
2SAM|13|20|dixit autem ei Absalom frater suus num Amnon frater tuus concubuit tecum sed nunc soror tace frater tuus est neque adfligas cor tuum pro re hac mansit itaque Thamar contabescens in domo Absalom fratris sui
2SAM|13|21|cum autem audisset rex David verba haec contristatus est valde
2SAM|13|22|porro non est locutus Absalom ad Amnon nec malum nec bonum oderat enim Absalom Amnon eo quod violasset Thamar sororem suam
2SAM|13|23|factum est autem post tempus biennii ut tonderentur oves Absalom in Baalasor quae est iuxta Ephraim et vocavit Absalom omnes filios regis
2SAM|13|24|venitque ad regem et ait ad eum ecce tondentur oves servi tui veniat oro rex cum servis suis ad servum suum
2SAM|13|25|dixitque rex ad Absalom noli fili mi noli rogare ut veniamus omnes et gravemus te cum autem cogeret eum et noluisset ire benedixit ei
2SAM|13|26|et ait Absalom si non vis venire veniat obsecro nobiscum saltem Amnon frater meus dixitque ad eum rex non est necesse ut vadat tecum
2SAM|13|27|coegit itaque eum Absalom et dimisit cum eo Amnon et universos filios regis
2SAM|13|28|praeceperat autem Absalom pueris suis dicens observate cum temulentus fuerit Amnon vino et dixero vobis percutite eum et interficite nolite timere ego enim sum qui praecepi vobis roboramini et estote viri fortes
2SAM|13|29|fecerunt ergo pueri Absalom adversum Amnon sicut praeceperat eis Absalom surgentesque omnes filii regis ascenderunt singuli mulas suas et fugerunt
2SAM|13|30|cumque adhuc pergerent in itinere fama praevenit ad David dicens percussit Absalom omnes filios regis et non remansit ex eis saltem unus
2SAM|13|31|surrexit itaque rex et scidit vestimenta sua et cecidit super terram et omnes servi ipsius qui adsistebant ei sciderunt vestimenta sua
2SAM|13|32|respondens autem Ionadab filius Samaa fratris David dixit ne aestimet dominus meus quod omnes pueri filii regis occisi sint Amnon solus mortuus est quoniam in ore Absalom erat positus ex die qua oppressit Thamar sororem eius
2SAM|13|33|nunc ergo ne ponat dominus meus rex super cor suum verbum istud dicens omnes filii regis occisi sunt quoniam Amnon solus mortuus est
2SAM|13|34|fugit autem Absalom et levavit puer speculator oculos suos et aspexit et ecce populus multus veniebat per iter devium ex latere montis
2SAM|13|35|dixit autem Ionadab ad regem ecce filii regis adsunt iuxta verbum servi tui sic factum est
2SAM|13|36|cumque cessasset loqui apparuerunt et filii regis et intrantes levaverunt vocem suam et fleverunt sed et rex et omnes servi eius fleverunt ploratu magno nimis
2SAM|13|37|porro Absalom fugiens abiit ad Tholomai filium Amiur regem Gessur luxit ergo David filium suum cunctis diebus
2SAM|13|38|Absalom autem cum fugisset et venisset in Gessur fuit ibi tribus annis
2SAM|13|39|cessavitque David rex persequi Absalom eo quod consolatus esset super Amnon interitu
2SAM|14|1|intellegens autem Ioab filius Sarviae quod cor regis versum esset ad Absalom
2SAM|14|2|misit Thecuam et tulit inde mulierem sapientem dixitque ad eam lugere te simula et induere veste lugubri et ne unguaris oleo ut sis quasi mulier plurimo iam tempore lugens mortuum
2SAM|14|3|et ingredieris ad regem et loqueris ad eum sermones huiuscemodi posuit autem Ioab verba in ore eius
2SAM|14|4|itaque cum ingressa fuisset mulier thecuites ad regem cecidit coram eo super terram et adoravit et dixit serva me rex
2SAM|14|5|et ait ad eam rex quid causae habes quae respondit heu mulier vidua ego sum mortuus est enim vir meus
2SAM|14|6|et ancillae tuae erant duo filii qui rixati sunt adversum se in agro nullusque erat qui eos prohibere posset et percussit alter alterum et interfecit eum
2SAM|14|7|et ecce consurgens universa cognatio adversum ancillam tuam dicit trade eum qui percussit fratrem suum ut occidamus eum pro anima fratris sui quem interfecit et deleamus heredem et quaerunt extinguere scintillam meam quae relicta est ut non supersit viro meo nomen et reliquiae super terram
2SAM|14|8|et ait rex ad mulierem vade in domum tuam et ego iubebo pro te
2SAM|14|9|dixitque mulier thecuites ad regem in me domine mi rex iniquitas et in domum patris mei rex autem et thronus eius sit innocens
2SAM|14|10|et ait rex qui contradixerit tibi adduc eum ad me et ultra non addet ut tangat te
2SAM|14|11|quae ait recordetur rex Domini Dei sui ut non multiplicentur proximi sanguinis ad ulciscendum et nequaquam interficient filium meum qui ait vivit Dominus quia non cadet de capillis filii tui super terram
2SAM|14|12|dixit ergo mulier loquatur ancilla tua ad dominum meum regem verbum et ait loquere
2SAM|14|13|dixitque mulier quare cogitasti istiusmodi rem contra populum Dei et locutus est rex verbum istud ut peccet et non reducat eiectum suum
2SAM|14|14|omnes morimur et quasi aquae delabimur in terram quae non revertuntur nec vult perire Deus animam sed retractat cogitans ne penitus pereat qui abiectus est
2SAM|14|15|nunc igitur veni ut loquar ad regem dominum meum verbum hoc praesente populo et dixit ancilla tua loquar ad regem si quo modo faciat rex verbum ancillae suae
2SAM|14|16|et audivit rex ut liberaret ancillam suam de manu omnium qui volebant delere me et filium meum simul de hereditate Dei
2SAM|14|17|dicat ergo ancilla tua ut fiat verbum domini mei regis quasi sacrificium sicut enim angelus Dei sic est dominus meus rex ut nec benedictione nec maledictione moveatur unde et Dominus Deus tuus est tecum
2SAM|14|18|et respondens rex dixit ad mulierem ne abscondas a me verbum quod te interrogo dixitque mulier loquere domine mi rex
2SAM|14|19|et ait rex numquid manus Ioab tecum est in omnibus istis respondit mulier et ait per salutem animae tuae domine mi rex nec ad dextram nec ad sinistram est ex omnibus his quae locutus est dominus meus rex servus enim tuus Ioab ipse praecepit mihi et ipse posuit in os ancillae tuae omnia verba haec
2SAM|14|20|ut verterem figuram sermonis huius servus tuus Ioab praecepit istud tu autem domine mi sapiens es sicut habet sapientiam angelus Dei ut intellegas omnia super terram
2SAM|14|21|et ait rex ad Ioab ecce placatus feci verbum tuum vade igitur et revoca puerum Absalom
2SAM|14|22|cadensque Ioab super faciem suam in terram adoravit et benedixit regi et dixit Ioab hodie intellexit servus tuus quia inveni gratiam in oculis tuis domine mi rex fecisti enim sermonem servi tui
2SAM|14|23|surrexit ergo Ioab et abiit in Gessur et adduxit Absalom in Hierusalem
2SAM|14|24|dixit autem rex revertatur in domum suam et faciem meam non videat reversus est itaque Absalom in domum suam et faciem regis non vidit
2SAM|14|25|porro sicut Absalom vir non erat pulcher in omni Israhel et decorus nimis a vestigio pedis usque ad verticem non erat in eo ulla macula
2SAM|14|26|et quando tondebatur capillum semel autem in anno tondebatur quia gravabat eum caesaries ponderabat capillos capitis sui ducentis siclis pondere publico
2SAM|14|27|nati sunt autem Absalom filii tres et filia una nomine Thamar eleganti forma
2SAM|14|28|mansitque Absalom Hierusalem duobus annis et faciem regis non vidit
2SAM|14|29|misit itaque ad Ioab ut mitteret eum ad regem qui noluit venire ad eum cumque secundo misisset et ille noluisset venire
2SAM|14|30|dixit servis suis scitis agrum Ioab iuxta agrum meum habentem messem hordei ite igitur et succendite eum igni succenderunt ergo servi Absalom segetem igni
2SAM|14|31|surrexitque Ioab et venit ad Absalom in domum eius et dixit quare succenderunt servi tui segetem meam igni
2SAM|14|32|et respondit Absalom ad Ioab misi ad te obsecrans ut venires ad me et mitterem te ad regem ut diceres ei quare veni de Gessur melius mihi erat ibi esse obsecro ergo ut videam faciem regis quod si memor est iniquitatis meae interficiat me
2SAM|14|33|ingressus Ioab ad regem nuntiavit ei vocatusque Absalom intravit ad regem et adoravit super faciem terrae coram eo osculatusque est rex Absalom
2SAM|15|1|igitur post haec fecit sibi Absalom currum et equites et quinquaginta viros qui praecederent eum
2SAM|15|2|et mane consurgens Absalom stabat iuxta introitum portae et omnem virum qui habebat negotium ut veniret ad regis iudicium vocabat Absalom ad se et dicebat de qua civitate es tu qui respondens aiebat ex una tribu Israhel ego sum servus tuus
2SAM|15|3|respondebatque ei Absalom videntur mihi sermones tui boni et iusti sed non est qui te audiat constitutus a rege dicebatque Absalom
2SAM|15|4|quis me constituat iudicem super terram ut ad me veniant omnes qui habent negotium et iuste iudicem
2SAM|15|5|sed et cum accederet ad eum homo ut salutaret illum extendebat manum suam et adprehendens osculabatur eum
2SAM|15|6|faciebatque hoc omni Israhel qui veniebat ad iudicium ut audiretur a rege et sollicitabat corda virorum Israhel
2SAM|15|7|post quattuor autem annos dixit Absalom ad regem vadam et reddam vota mea quae vovi Domino in Hebron
2SAM|15|8|vovens enim vovit servus tuus cum esset in Gessur Syriae dicens si reduxerit me Dominus in Hierusalem sacrificabo Domino
2SAM|15|9|dixitque ei rex vade in pace et surrexit et abiit in Hebron
2SAM|15|10|misit autem Absalom exploratores in universas tribus Israhel dicens statim ut audieritis clangorem bucinae dicite regnavit Absalom in Hebron
2SAM|15|11|porro cum Absalom ierunt ducenti viri de Hierusalem vocati euntes simplici corde et causam penitus ignorantes
2SAM|15|12|accersivit quoque Absalom Ahitofel Gilonitem consiliarium David de civitate sua Gilo cum immolaret victimas et facta est coniuratio valida populusque concurrens augebatur cum Absalom
2SAM|15|13|venit igitur nuntius ad David dicens toto corde universus Israhel sequitur Absalom
2SAM|15|14|et ait David servis suis qui erant cum eo in Hierusalem surgite fugiamus neque enim erit nobis effugium a facie Absalom festinate egredi ne forte veniens occupet nos et inpellat super nos ruinam et percutiat civitatem in ore gladii
2SAM|15|15|dixeruntque servi regis ad eum omnia quaecumque praeceperit dominus noster rex libenter exsequimur servi tui
2SAM|15|16|egressus est ergo rex et universa domus eius pedibus suis et dereliquit rex decem mulieres concubinas ad custodiendam domum
2SAM|15|17|egressusque rex et omnis Israhel pedibus suis stetit procul a domo
2SAM|15|18|et universi servi eius ambulabant iuxta eum et legiones Cherethi et Felethi et omnes Getthei sescenti viri qui secuti eum fuerant de Geth praecedebant regem
2SAM|15|19|dixit autem rex ad Ethai Gettheum cur venis nobiscum revertere et habita cum rege quia peregrinus es et egressus de loco tuo
2SAM|15|20|heri venisti et hodie inpelleris nobiscum egredi ego autem vadam quo iturus sum revertere et reduc tecum fratres tuos ostendisti gratiam et fidem
2SAM|15|21|et respondit Ethai regi dicens vivit Dominus et vivit dominus meus rex quoniam in quocumque loco fueris domine mi rex sive in morte sive in vita ibi erit servus tuus
2SAM|15|22|et ait David Ethai veni et transi et transivit Ethai Gettheus et omnes viri qui cum eo erant et reliqua multitudo
2SAM|15|23|omnesque flebant voce magna et universus populus transiebat rex quoque transgrediebatur torrentem Cedron et cunctus populus incedebat contra viam quae respicit ad desertum
2SAM|15|24|venit autem et Sadoc et universi Levitae cum eo portantes arcam foederis Dei et deposuerunt arcam Dei et ascendit Abiathar donec expletus est omnis populus qui egressus fuerat de civitate
2SAM|15|25|et dixit rex ad Sadoc reporta arcam Dei in urbem si invenero gratiam in oculis Domini reducet me et ostendet mihi eam et tabernaculum suum
2SAM|15|26|si autem dixerit non places praesto sum faciat quod bonum est coram se
2SAM|15|27|et dixit rex ad Sadoc sacerdotem o videns revertere in civitatem in pace et Achimaas filius tuus et Ionathan filius Abiathar duo filii vestri sint vobiscum
2SAM|15|28|ecce ego abscondar in campestribus deserti donec veniat sermo a vobis indicans mihi
2SAM|15|29|reportaverunt igitur Sadoc et Abiathar arcam Dei Hierusalem et manserunt ibi
2SAM|15|30|porro David ascendebat clivum Olivarum scandens et flens operto capite et nudis pedibus incedens sed et omnis populus qui erat cum eo operto capite ascendebat plorans
2SAM|15|31|nuntiatum est autem David quod et Ahitofel esset in coniuratione cum Absalom dixitque David infatua quaeso consilium Ahitofel Domine
2SAM|15|32|cumque ascenderet David summitatem montis in quo adoraturus erat Dominum ecce occurrit ei Husai Arachites scissa veste et terra pleno capite
2SAM|15|33|et dixit ei David si veneris mecum eris mihi oneri
2SAM|15|34|si autem in civitatem revertaris et dixeris Absalom servus tuus sum rex sicut fui servus patris tui sic ero servus tuus dissipabis consilium Ahitofel
2SAM|15|35|habes autem tecum Sadoc et Abiathar sacerdotes et omne verbum quodcumque audieris de domo regis indicabis Sadoc et Abiathar sacerdotibus
2SAM|15|36|sunt autem cum eis duo filii eorum Achimaas Sadoc et Ionathan Abiathar et mittetis per eos ad me omne verbum quod audieritis
2SAM|15|37|veniente ergo Husai amico David in civitatem Absalom quoque ingressus est Hierusalem
2SAM|16|1|cumque David transisset paululum montis verticem apparuit Siba puer Mifiboseth in occursum eius cum duobus asinis qui onerati erant ducentis panibus et centum alligaturis uvae passae et centum massis palatarum et utribus vini
2SAM|16|2|et dixit rex Sibae quid sibi volunt haec responditque Siba asini domestici regis ut sedeant et panes et palatae ad vescendum pueris tuis vinum autem ut bibat si quis defecerit in deserto
2SAM|16|3|et ait rex ubi est filius domini tui responditque Siba regi remansit in Hierusalem dicens hodie restituet mihi domus Israhel regnum patris mei
2SAM|16|4|et ait rex Sibae tua sint omnia quae fuerunt Mifiboseth dixitque Siba adoro inveniam gratiam coram te domine mi rex
2SAM|16|5|venit ergo rex David usque Baurim et ecce egrediebatur inde vir de cognatione domus Saul nomine Semei filius Gera procedebat egrediens et maledicebat
2SAM|16|6|mittebatque lapides contra David et contra universos servos regis David omnis autem populus et universi bellatores a dextro et sinistro latere regis incedebant
2SAM|16|7|ita autem loquebatur Semei cum malediceret regi egredere egredere vir sanguinum et vir Belial
2SAM|16|8|reddidit tibi Dominus universum sanguinem domus Saul quoniam invasisti regnum pro eo et dedit Dominus regnum in manu Absalom filii tui et ecce premunt te mala tua quoniam vir sanguinum es
2SAM|16|9|dixit autem Abisai filius Sarviae regi quare maledicit canis hic moriturus domino meo regi vadam et amputabo caput eius
2SAM|16|10|et ait rex quid mihi et vobis filii Sarviae dimittite eum maledicat Dominus enim praecepit ei ut malediceret David et quis est qui audeat dicere quare sic fecerit
2SAM|16|11|et ait rex Abisai et universis servis suis ecce filius meus qui egressus est de utero meo quaerit animam meam quanto magis nunc filius Iemini dimittite eum ut maledicat iuxta praeceptum Domini
2SAM|16|12|si forte respiciat Dominus adflictionem meam et reddat mihi bonum pro maledictione hac hodierna
2SAM|16|13|ambulabat itaque David et socii eius per viam cum eo Semei autem per iugum montis ex latere contra illum gradiebatur maledicens et mittens lapides adversum eum terramque spargens
2SAM|16|14|venit itaque rex et universus populus cum eo lassus et refocilati sunt ibi
2SAM|16|15|Absalom autem et omnis populus Israhel ingressi sunt Hierusalem sed et Ahitofel cum eo
2SAM|16|16|cum autem venisset Husai Arachites amicus David ad Absalom locutus est ad eum salve rex salve rex
2SAM|16|17|ad quem Absalom haec est inquit gratia tua ad amicum tuum quare non isti cum amico tuo
2SAM|16|18|responditque Husai ad Absalom nequaquam quia illius ero quem elegit Dominus et omnis hic populus et universus Israhel et cum eo manebo
2SAM|16|19|sed ut et hoc inferam cui ego serviturus sum nonne filio regis sicut parui patri tuo sic parebo et tibi
2SAM|16|20|dixit autem Absalom ad Ahitofel inite consilium quid agere debeamus
2SAM|16|21|et ait Ahitofel ad Absalom ingredere ad concubinas patris tui quas dimisit ad custodiendam domum ut cum audierit omnis Israhel quod foedaveris patrem tuum roborentur manus eorum tecum
2SAM|16|22|tetenderunt igitur Absalom tabernaculum in solario ingressusque est ad concubinas patris sui coram universo Israhel
2SAM|16|23|consilium autem Ahitofel quod dabat in diebus illis quasi si quis consuleret Deum sic erat omne consilium Ahitofel et cum esset cum David et cum esset cum Absalom
2SAM|17|1|dixit igitur Ahitofel ad Absalom eligam mihi duodecim milia virorum et consurgens persequar David hac nocte
2SAM|17|2|et inruens super eum quippe qui lassus est et solutis manibus percutiam eum cumque fugerit omnis populus qui cum eo est percutiam regem desolatum
2SAM|17|3|et reducam universum populum quomodo omnis reverti solet unum enim virum tu quaeris et omnis populus erit in pace
2SAM|17|4|placuitque sermo eius Absalom et cunctis maioribus natu Israhel
2SAM|17|5|ait autem Absalom vocate et Husai Arachiten et audiamus quid etiam ipse dicat
2SAM|17|6|cumque venisset Husai ad Absalom ait Absalom ad eum huiuscemodi sermonem locutus est Ahitofel facere debemus an non quod das consilium
2SAM|17|7|et dixit Husai ad Absalom non bonum consilium quod dedit Ahitofel hac vice
2SAM|17|8|et rursum intulit Husai tu nosti patrem tuum et viros qui cum eo sunt esse fortissimos et amaro animo veluti si ursa raptis catulis in saltu saeviat sed et pater tuus vir bellator est nec morabitur cum populo
2SAM|17|9|forsitan nunc latitat in foveis aut in uno quo voluerit loco et cum ceciderit unus quilibet in principio audiet quicumque audierit et dicet facta est plaga in populo qui sequebatur Absalom
2SAM|17|10|et fortissimus quoque cuius cor est quasi leonis pavore solvetur scit enim omnis populus Israhel fortem esse patrem tuum et robustos omnes qui cum eo sunt
2SAM|17|11|sed hoc mihi videtur rectum esse consilium congregetur ad te universus Israhel a Dan usque Bersabee quasi harena maris innumerabilis et tu eris in medio eorum
2SAM|17|12|et inruemus super eum in quocumque loco fuerit inventus et operiemus eum sicut cadere solet ros super terram et non relinquemus de viris qui cum eo sunt ne unum quidem
2SAM|17|13|quod si urbem aliquam fuerit ingressus circumdabit omnis Israhel civitati illi funes et trahemus eam in torrentem ut non repperiatur nec calculus quidem ex ea
2SAM|17|14|dixitque Absalom et omnis vir Israhel melius consilium Husai Arachitae consilio Ahitofel Domini autem nutu dissipatum est consilium Ahitofel utile ut induceret Dominus super Absalom malum
2SAM|17|15|et ait Husai Sadoc et Abiathar sacerdotibus hoc et hoc modo consilium dedit Ahitofel Absalom et senibus Israhel et ego tale et tale dedi consilium
2SAM|17|16|nunc ergo mittite cito et nuntiate David dicentes ne moremini nocte hac in campestribus deserti sed absque dilatione transgredere ne forte absorbeatur rex et omnis populus qui cum eo est
2SAM|17|17|Ionathan autem et Achimaas stabant iuxta fontem Rogel abiit ancilla et nuntiavit eis et illi profecti sunt ut referrent ad regem David nuntium non enim poterant videri aut introire civitatem
2SAM|17|18|vidit autem eos quidam puer et indicavit Absalom illi vero concito gradu ingressi sunt domum cuiusdam viri in Baurim qui habebat puteum in vestibulo suo et descenderunt in eum
2SAM|17|19|tulit autem mulier et expandit velamen super os putei quasi siccans ptisanas et sic res latuit
2SAM|17|20|cumque venissent servi Absalom ad mulierem in domum dixerunt ubi est Achimaas et Ionathan et respondit eis mulier transierunt gustata paululum aqua at hii qui quaerebant cum non repperissent reversi sunt Hierusalem
2SAM|17|21|cumque abissent ascenderunt illi de puteo et pergentes nuntiaverunt regi David atque dixerunt surgite transite cito fluvium quoniam huiuscemodi dedit consilium contra vos Ahitofel
2SAM|17|22|surrexit ergo David et omnis populus qui erat cum eo et transierunt Iordanem donec dilucesceret et ne unus quidem residuus fuit qui non transisset fluvium
2SAM|17|23|porro Ahitofel videns quod non fuisset factum consilium suum stravit asinum suum et surrexit et abiit in domum suam et in civitatem suam et disposita domo sua suspendio interiit et sepultus est in sepulchro patris sui
2SAM|17|24|David autem venit in Castra et Absalom transivit Iordanem ipse et omnis vir Israhel cum eo
2SAM|17|25|Amasam vero constituit Absalom pro Ioab super exercitum Amasa autem erat filius viri qui vocabatur Iethra de Hiesreli qui ingressus est ad Abigail filiam Naas sororem Sarviae quae fuit mater Ioab
2SAM|17|26|et castrametatus est Israhel cum Absalom in terra Galaad
2SAM|17|27|cumque venisset David in Castra Sobi filius Naas de Rabbath filiorum Ammon et Machir filius Ammihel de Lodabar et Berzellai Galaadites de Rogelim
2SAM|17|28|obtulerunt ei stratoria et tappetia et vasa fictilia frumentum et hordeum et farinam pulentam et fabam et lentem frixum cicer
2SAM|17|29|et mel et butyrum oves et pingues vitulos dederuntque David et populo qui cum eo erat ad vescendum suspicati enim sunt populum fame et siti fatigari in deserto
2SAM|18|1|igitur considerato David populo suo constituit super eum tribunos et centuriones
2SAM|18|2|et dedit populi tertiam partem sub manu Ioab et tertiam in manu Abisai filii Sarviae fratris Ioab et tertiam sub manu Ethai qui erat de Geth dixitque rex ad populum egrediar et ego vobiscum
2SAM|18|3|et respondit populus non exibis sive enim fugerimus non magnopere ad eos de nobis pertinebit sive media pars ceciderit e nobis non satis curabunt quia tu unus pro decem milibus conputaris melius est igitur ut sis nobis in urbe praesidio
2SAM|18|4|ad quos rex ait quod vobis rectum videtur hoc faciam stetit ergo rex iuxta portam egrediebaturque populus per turmas suas centeni et milleni
2SAM|18|5|et praecepit rex Ioab et Abisai et Ethai dicens servate mihi puerum Absalom et omnis populus audiebat praecipientem regem cunctis principibus pro Absalom
2SAM|18|6|itaque egressus est populus in campum contra Israhel et factum est proelium in saltu Ephraim
2SAM|18|7|et caesus est ibi populus Israhel ab exercitu David factaque est ibi plaga magna in die illa viginti milium
2SAM|18|8|fuit autem ibi proelium dispersum super faciem omnis terrae et multo plures erant quos saltus consumpserat de populo quam hii quos voraverat gladius in die illa
2SAM|18|9|accidit autem ut occurreret Absalom servis David sedens mulo cumque ingressus fuisset mulus subter condensam quercum et magnam adhesit caput eius quercui et illo suspenso inter caelum et terram mulus cui sederat pertransivit
2SAM|18|10|vidit autem hoc quispiam et nuntiavit Ioab dicens vidi Absalom pendere de quercu
2SAM|18|11|et ait Ioab viro qui nuntiaverat ei si vidisti quare non confodisti eum cum terra et ego dedissem tibi decem argenti siclos et unum balteum
2SAM|18|12|qui dixit ad Ioab si adpenderes in manibus meis mille argenteos nequaquam mitterem manum meam in filium regis audientibus enim nobis praecepit rex tibi et Abisai et Ethai dicens custodite mihi puerum Absalom
2SAM|18|13|sed et si fecissem contra animam meam audacter nequaquam hoc regem latere potuisset et tu stares ex adverso
2SAM|18|14|et ait Ioab non sicut tu vis sed adgrediar eum coram te tulit ergo tres lanceas in manu sua et infixit eas in corde Absalom cumque adhuc palpitaret herens in quercu
2SAM|18|15|cucurrerunt decem iuvenes armigeri Ioab et percutientes interfecerunt eum
2SAM|18|16|cecinit autem Ioab bucina et retinuit populum ne persequeretur fugientem Israhel volens parcere multitudini
2SAM|18|17|et tulerunt Absalom et proiecerunt eum in saltu in foveam grandem et conportaverunt super eum acervum lapidum magnum nimis omnis autem Israhel fugit in tabernacula sua
2SAM|18|18|porro Absalom erexerat sibi cum adhuc viveret titulum qui est in valle Regis dixerat enim non habeo filium et hoc erit monumentum nominis mei vocavitque titulum nomine suo et appellatur manus Absalom usque ad hanc diem
2SAM|18|19|Achimaas autem filius Sadoc ait curram et nuntiabo regi quia iudicium fecerit ei Dominus de manu inimicorum eius
2SAM|18|20|ad quem Ioab dixit non eris nuntius in hac die sed nuntiabis in alia hodie nolo te nuntiare filius enim regis est mortuus
2SAM|18|21|et ait Ioab Chusi vade et nuntia regi quae vidisti adoravit Chusi Ioab et cucurrit
2SAM|18|22|rursum autem Achimaas filius Sadoc dixit ad Ioab quid inpedit si etiam ego curram post Chusi dixitque Ioab quid vis currere fili mi non eris boni nuntii baiulus
2SAM|18|23|qui respondit quid enim si cucurrero et ait ei curre currens ergo Achimaas per viam conpendii transivit Chusi
2SAM|18|24|David autem sedebat inter duas portas speculator vero qui erat in fastigio portae super murum elevans oculos vidit hominem currentem solum
2SAM|18|25|et exclamans indicavit regi dixitque rex si solus est bonus est nuntius in ore eius properante autem illo et accedente propius
2SAM|18|26|vidit speculator hominem alterum currentem et vociferans in culmine ait apparet mihi homo currens solus dixitque rex et iste bonus est nuntius
2SAM|18|27|speculator autem contemplor ait cursum prioris quasi cursum Achimaas filii Sadoc et ait rex vir bonus est et nuntium portans bonum venit
2SAM|18|28|clamans autem Achimaas dixit ad regem salve et adorans regem coram eo pronus in terram ait benedictus Dominus Deus tuus qui conclusit homines qui levaverunt manus suas contra dominum meum regem
2SAM|18|29|et ait rex estne pax puero Absalom dixitque Achimaas vidi tumultum magnum cum mitteret Ioab servus tuus o rex me servum tuum nescio aliud
2SAM|18|30|ad quem rex transi ait et sta hic cumque ille transisset et staret
2SAM|18|31|apparuit Chusi et veniens ait bonum adporto nuntium domine mi rex iudicavit enim pro te Dominus hodie de manu omnium qui surrexerunt contra te
2SAM|18|32|dixit autem rex ad Chusi estne pax puero Absalom cui respondens Chusi fiant inquit sicut puer inimici domini mei regis et universi qui consurgunt adversum eum in malum
2SAM|18|33|contristatus itaque rex ascendit cenaculum portae et flevit et sic loquebatur vadens fili mi Absalom fili mi Absalom quis mihi tribuat ut ego moriar pro te Absalom fili mi fili mi
2SAM|19|1|nuntiatum est autem Ioab quod rex fleret et lugeret filium suum
2SAM|19|2|et versa est victoria in die illa in luctum omni populo audivit enim populus in die illa dici dolet rex super filio suo
2SAM|19|3|et declinabat populus in die illa ingredi civitatem quomodo declinare solet populus versus et fugiens de proelio
2SAM|19|4|porro rex operuit caput suum et clamabat voce magna fili mi Absalom Absalom fili mi fili mi
2SAM|19|5|ingressus ergo Ioab ad regem in domo dixit confudisti hodie vultus omnium servorum tuorum qui salvam fecerunt animam tuam et animam filiorum tuorum et filiarum tuarum et animam uxorum tuarum et animam concubinarum tuarum
2SAM|19|6|diligis odientes te et odio habes diligentes te et ostendisti hodie quia non curas de ducibus tuis et de servis tuis et vere cognovi modo quia si Absalom viveret et nos omnes occubuissemus tunc placeret tibi
2SAM|19|7|nunc igitur surge et procede et adloquens satisfac servis tuis iuro enim tibi per Dominum quod si non exieris ne unus quidem remansurus sit tecum nocte hac et peius erit hoc tibi quam omnia mala quae venerunt super te ab adulescentia tua usque in praesens
2SAM|19|8|surrexit ergo rex et sedit in porta et omni populo nuntiatum est quod rex sederet in porta venitque universa multitudo coram rege Israhel autem fugit in tabernacula sua
2SAM|19|9|omnis quoque populus certabat in cunctis tribubus Israhel dicens rex liberavit nos de manu inimicorum nostrorum ipse salvavit nos de manu Philisthinorum et nunc fugit de terra propter Absalom
2SAM|19|10|Absalom autem quem unximus super nos mortuus est in bello usquequo siletis et non reducitis regem
2SAM|19|11|rex vero David misit ad Sadoc et ad Abiathar sacerdotes dicens loquimini ad maiores natu Iuda dicentes cur venitis novissimi ad reducendum regem in domum suam sermo autem omnis Israhel pervenerat ad regem in domo eius
2SAM|19|12|fratres mei vos os meum et caro mea vos quare novissimi reducitis regem
2SAM|19|13|et Amasae dicite nonne os meum es et caro mea haec faciat mihi Deus et haec addat si non magister militiae fueris coram me omni tempore pro Ioab
2SAM|19|14|et inclinavit cor omnium virorum Iuda quasi viri unius miseruntque ad regem dicentes revertere tu et omnes servi tui
2SAM|19|15|et reversus est rex et venit usque ad Iordanem et Iuda venit in Galgala ut occurreret regi et transduceret eum Iordanem
2SAM|19|16|festinavit autem Semei filius Gera filii Iemini de Baurim et descendit cum viris Iuda in occursum regis David
2SAM|19|17|cum mille viris de Beniamin et Siba puer de domo Saul et quindecim filii eius ac viginti servi erant cum eo et inrumpentes Iordanem ante regem
2SAM|19|18|transierunt vada ut transducerent domum regis et facerent iuxta iussionem eius Semei autem filius Gera prostratus coram rege cum iam transisset Iordanem
2SAM|19|19|dixit ad eum ne reputes mihi domine mi iniquitatem neque memineris iniuriam servi tui in die qua egressus es domine mi rex de Hierusalem neque ponas rex in corde tuo
2SAM|19|20|agnosco enim servus tuus peccatum meum et idcirco hodie primus veni de omni domo Ioseph descendique in occursum domini mei regis
2SAM|19|21|respondens vero Abisai filius Sarviae dixit numquid pro his verbis non occidetur Semei quia maledixit christo Domini
2SAM|19|22|et ait David quid mihi et vobis filii Sarviae cur efficimini mihi hodie in Satan ergone hodie interficietur vir in Israhel an ignoro hodie me factum regem super Israhel
2SAM|19|23|et ait rex Semei non morieris iuravitque ei
2SAM|19|24|Mifiboseth quoque filius Saul descendit in occursum regis inlotis pedibus et intonsa barba vestesque suas non laverat a die qua egressus fuerat rex usque ad diem reversionis eius in pace
2SAM|19|25|cumque Hierusalem occurrisset regi dixit ei rex quare non venisti mecum Mifiboseth
2SAM|19|26|qui respondens ait domine mi rex servus meus contempsit me dixi ei ego famulus tuus ut sterneret mihi asinum et ascendens abirem cum rege claudus enim sum servus tuus
2SAM|19|27|insuper et accusavit me servum tuum ad te dominum meum regem tu autem domine mi rex sicut angelus Dei fac quod placitum est tibi
2SAM|19|28|neque enim fuit domus patris mei nisi morti obnoxia domino meo regi tu autem posuisti me servum tuum inter convivas mensae tuae quid igitur habeo iustae querellae aut quid possum ultra vociferari ad regem
2SAM|19|29|ait ergo ei rex quid ultra loqueris fixum est quod locutus sum tu et Siba dividite possessiones
2SAM|19|30|responditque Mifiboseth regi etiam cuncta accipiat postquam reversus est dominus meus rex pacifice in domum suam
2SAM|19|31|Berzellai quoque Galaadites descendens de Rogelim transduxit regem Iordanem paratus etiam ultra fluvium prosequi eum
2SAM|19|32|erat autem Berzellai Galaadites senex valde id est octogenarius et ipse praebuit alimenta regi cum moraretur in Castris fuit quippe vir dives nimis
2SAM|19|33|dixit itaque rex ad Berzellai veni mecum ut requiescas secure mecum in Hierusalem
2SAM|19|34|et ait Berzellai ad regem quot sunt dies annorum vitae meae ut ascendam cum rege Hierusalem
2SAM|19|35|octogenarius sum hodie numquid vigent sensus mei ad discernendum suave aut amarum aut delectare potest servum tuum cibus et potus vel audire ultra possum vocem cantorum atque cantricum quare servus tuus fit oneri domino meo regi
2SAM|19|36|paululum procedam famulus tuus ab Iordane tecum nec indigeo hac vicissitudine
2SAM|19|37|sed obsecro ut revertar servus tuus et moriar in civitate mea iuxta sepulchrum patris mei et matris meae est autem servus tuus Chamaam ipse vadat tecum domine mi rex et fac ei quod tibi bonum videtur
2SAM|19|38|dixitque rex mecum transeat Chamaam et ego faciam ei quicquid tibi placuerit et omne quod petieris a me inpetrabis
2SAM|19|39|cumque transisset universus populus et rex Iordanem osculatus est rex Berzellai et benedixit ei et ille reversus est in locum suum
2SAM|19|40|transivit ergo rex in Galgalam et Chamaam cum eo omnis autem populus Iuda transduxerat regem et media tantum pars adfuerat de populo Israhel
2SAM|19|41|itaque omnes viri Israhel concurrentes ad regem dixerunt ei quare te furati sunt fratres nostri viri Iuda et transduxerunt regem et domum eius Iordanem omnesque viros David cum eo
2SAM|19|42|et respondit omnis vir Iuda ad viros Israhel quia propior mihi est rex cur irasceris super hac re numquid comedimus aliquid ex rege aut munera nobis data sunt
2SAM|19|43|et respondit vir Israhel ad viros Iuda et ait decem partibus maior ego sum apud regem magisque ad me pertinet David quam ad te cur mihi fecisti iniuriam et non mihi nuntiatum est priori ut reducerem regem meum durius autem responderunt viri Iuda viris Israhel
2SAM|20|1|accidit quoque ut ibi esset vir Belial nomine Seba filius Bochri vir iemineus et cecinit bucina et ait non est nobis pars in David neque hereditas in filio Isai vir in tabernacula tua Israhel
2SAM|20|2|et separatus est omnis Israhel a David secutusque est Seba filium Bochri viri autem Iuda adheserunt regi suo a Iordane usque Hierusalem
2SAM|20|3|cumque venisset rex in domum suam Hierusalem tulit decem mulieres concubinas quas dereliquerat ad custodiendam domum et tradidit eas in custodiam alimenta eis praebens et non est ingressus ad eas sed erant clausae usque ad diem mortis suae in viduitate viventes
2SAM|20|4|dixit autem rex Amasae convoca mihi omnes viros Iuda in diem tertium et tu adesto praesens
2SAM|20|5|abiit ergo Amasa ut convocaret Iudam et moratus est extra placitum quod ei constituerat
2SAM|20|6|ait autem David ad Abisai nunc magis adflicturus est nos Seba filius Bochri quam Absalom tolle igitur servos domini tui et persequere eum ne forte inveniat civitates munitas et effugiat nos
2SAM|20|7|egressi sunt ergo cum eo viri Ioab Cherethi quoque et Felethi et omnes robusti exierunt de Hierusalem ad persequendum Seba filium Bochri
2SAM|20|8|cumque illi essent iuxta lapidem grandem qui est in Gabaon Amasa veniens occurrit eis porro Ioab vestitus erat tunica stricta ad mensuram habitus sui et desuper accinctus gladio dependente usque ad ilia in vagina qui fabrefactus levi motu egredi poterat et percutere
2SAM|20|9|dixit itaque Ioab ad Amasa salve mi frater et tenuit manu dextra mentum Amasae quasi osculans eum
2SAM|20|10|porro Amasa non observavit gladium quem habebat Ioab qui percussit eum in latere et effudit intestina eius in terram nec secundum vulnus adposuit Ioab autem et Abisai frater eius persecuti sunt Seba filium Bochri
2SAM|20|11|interea quidam viri cum stetissent iuxta cadaver Amasae de sociis Ioab dixerunt ecce qui esse voluit pro Ioab comes David pro Ioab
2SAM|20|12|Amasa autem conspersus sanguine iacebat in media via vidit hoc quidam vir quod subsisteret omnis populus ad videndum eum et amovit Amasam de via in agrum operuitque eum vestimento ne subsisterent transeuntes propter eum
2SAM|20|13|amoto igitur illo de via transiebat omnis vir sequens Ioab ad persequendum Seba filium Bochri
2SAM|20|14|porro ille transierat per omnes tribus Israhel in Abelam et in Bethmacha omnesque electi congregati fuerant ad eum
2SAM|20|15|venerunt itaque et obpugnabant eum in Abela et in Bethmacha et circumdederunt munitionibus civitatem et obsessa est urbs omnis autem turba quae erat cum Ioab moliebatur destruere muros
2SAM|20|16|et exclamavit mulier sapiens de civitate audite audite dicite Ioab adpropinqua huc et loquar tecum
2SAM|20|17|qui cum accessisset ad eam ait illi tu es Ioab et ille respondit ego ad quem sic locuta est audi sermones ancillae tuae qui respondit audio
2SAM|20|18|rursumque illa sermo inquit dicebatur in veteri proverbio qui interrogant interrogent in Abela et sic perficiebant
2SAM|20|19|nonne ego sum quae respondeo veritatem Israhel et tu quaeris subruere civitatem et evertere matrem in Israhel quare praecipitas hereditatem Domini
2SAM|20|20|respondensque Ioab ait absit absit hoc a me non praecipito neque demolior
2SAM|20|21|non se sic habet res sed homo de monte Ephraim Seba filius Bochri cognomine levavit manum contra regem David tradite illum solum et recedemus a civitate et ait mulier ad Ioab ecce caput eius mittetur ad te per murum
2SAM|20|22|ingressa est ergo ad omnem populum et locuta est eis sapienter qui abscisum caput Seba filii Bochri proiecerunt ad Ioab et ille cecinit tuba et recesserunt ab urbe unusquisque in tabernacula sua Ioab autem reversus est Hierusalem ad regem
2SAM|20|23|fuit ergo Ioab super omnem exercitum Israhel Banaias autem filius Ioiadae super Cheretheos et Feletheos
2SAM|20|24|Aduram vero super tributa porro Iosaphat filius Ahilud a commentariis
2SAM|20|25|Sia autem scriba Sadoc vero et Abiathar sacerdotes
2SAM|20|26|Hira autem Hiaiarites erat sacerdos David
2SAM|21|1|facta est quoque fames in diebus David tribus annis iugiter et consuluit David oraculum Domini dixitque Dominus propter Saul et domum eius et sanguinem quia occidit Gabaonitas
2SAM|21|2|vocatis ergo Gabaonitis rex dixit ad eos porro Gabaonitae non sunt de filiis Israhel sed reliquiae Amorreorum filii quippe Israhel iuraverant eis et voluit Saul percutere eos zelo quasi pro filiis Israhel et Iuda
2SAM|21|3|dixit ergo David ad Gabaonitas quid faciam vobis et quod erit vestri piaculum ut benedicatis hereditati Domini
2SAM|21|4|dixeruntque ei Gabaonitae non est nobis super argento et auro quaestio contra Saul et contra domum eius neque volumus ut interficiatur homo de Israhel ad quos ait quid ergo vultis ut faciam vobis
2SAM|21|5|qui dixerunt regi virum qui adtrivit nos et oppressit inique ita delere debemus ut ne unus quidem residuus sit de stirpe eius in cunctis finibus Israhel
2SAM|21|6|dentur nobis septem viri de filiis eius et crucifigamus eos Domino in Gabaath Saul quondam electi Domini et ait rex ego dabo
2SAM|21|7|pepercitque rex Mifiboseth filio Ionathan filii Saul propter iusiurandum Domini quod fuerat inter David et inter Ionathan filium Saul
2SAM|21|8|tulit itaque rex duos filios Respha filiae Ahia quos peperit Saul Armoni et Mifiboseth et quinque filios Michol filiae Saul quos genuerat Hadriheli filio Berzellai qui fuit de Molathi
2SAM|21|9|et dedit eos in manu Gabaonitarum qui crucifixerunt illos in monte coram Domino et ceciderunt hii septem simul occisi in diebus messis primis incipiente messione hordei
2SAM|21|10|tollens autem Respha filia Ahia cilicium substravit sibi super petram ab initio messis donec stillaret aqua super eos de caelo et non dimisit aves lacerare eos per diem neque bestias per noctem
2SAM|21|11|et nuntiata sunt David quae fecerat Respha filia Ahia concubina Saul
2SAM|21|12|et abiit David et tulit ossa Saul et ossa Ionathan filii eius a viris Iabesgalaad qui furati fuerant ea de platea Bethsan in qua suspenderant eos Philisthim cum interfecissent Saul in Gelboe
2SAM|21|13|et asportavit inde ossa Saul et ossa Ionathan filii eius et colligentes ossa eorum qui adfixi fuerant
2SAM|21|14|sepelierunt ea cum ossibus Saul et Ionathan filii eius in terra Beniamin in latere in sepulchro Cis patris eius feceruntque omnia quae praeceperat rex et repropitiatus est Deus terrae post haec
2SAM|21|15|factum est autem rursum proelium Philisthinorum adversum Israhel et descendit David et servi eius cum eo et pugnabant contra Philisthim deficiente autem David
2SAM|21|16|Iesbidenob qui fuit de genere Arafa cuius ferrum hastae trecentas uncias adpendebat et accinctus erat ense novo nisus est percutere David
2SAM|21|17|praesidioque ei fuit Abisai filius Sarviae et percussum Philistheum interfecit tunc iuraverunt viri David dicentes non egredieris nobiscum in bellum ne extinguas lucernam Israhel
2SAM|21|18|secundum quoque fuit bellum in Gob contra Philistheos tunc percussit Sobbochai de Usathi Seph de stirpe Arafa
2SAM|21|19|tertium quoque fuit bellum in Gob contra Philistheos in quo percussit Adeodatus filius Saltus polymitarius bethleemites Goliath Gettheum cuius hastile hastae erat quasi liciatorium texentium
2SAM|21|20|quartum bellum fuit in Geth in quo vir excelsus qui senos in manibus pedibusque habebat digitos id est viginti et quattuor et erat de origine Arafa
2SAM|21|21|blasphemavit Israhel percussit autem eum Ionathan filius Sammaa fratris David
2SAM|21|22|hii quattuor nati sunt de Arafa in Geth et ceciderunt in manu David et servorum eius
2SAM|22|1|locutus est autem David Domino verba carminis huius in die qua liberavit eum Dominus de manu omnium inimicorum suorum et de manu Saul
2SAM|22|2|et ait Dominus petra mea et robur meum et salvator meus
2SAM|22|3|Deus meus fortis meus sperabo in eum scutum meum et cornu salutis meae elevator meus et refugium meum salvator meus de iniquitate liberabis me
2SAM|22|4|laudabilem invocabo Dominum et ab inimicis meis salvus ero
2SAM|22|5|quia circumdederunt me contritiones mortis torrentes Belial terruerunt me
2SAM|22|6|funes inferi circumdederunt me praevenerunt me laquei mortis
2SAM|22|7|in tribulatione mea invocabo Dominum et ad Deum meum clamabo et exaudiet de templo suo vocem meam et clamor meus veniet ad aures eius
2SAM|22|8|commota est et contremuit terra fundamenta montium concussa sunt et conquassata quoniam iratus est
2SAM|22|9|ascendit fumus de naribus eius et ignis de ore eius voravit carbones incensi sunt ab eo
2SAM|22|10|et inclinavit caelos et descendit et caligo sub pedibus eius
2SAM|22|11|et ascendit super cherubin et volavit et lapsus est super pinnas venti
2SAM|22|12|posuit tenebras in circuitu suo latibulum cribrans aquas de nubibus caelorum
2SAM|22|13|prae fulgore in conspectu eius succensi sunt carbones ignis
2SAM|22|14|tonabit de caelis Dominus et Excelsus dabit vocem suam
2SAM|22|15|misit sagittas et dissipavit eos fulgur et consumpsit eos
2SAM|22|16|et apparuerunt effusiones maris et revelata sunt fundamenta orbis ab increpatione Domini ab inspiratione spiritus furoris eius
2SAM|22|17|misit de excelso et adsumpsit me extraxit me de aquis multis
2SAM|22|18|liberavit me ab inimico meo potentissimo ab his qui oderant me quoniam robustiores me erant
2SAM|22|19|praevenit me in die adflictionis meae et factus est Dominus firmamentum meum
2SAM|22|20|et eduxit me in latitudinem liberavit me quia placuit ei
2SAM|22|21|retribuet mihi Dominus secundum iustitiam meam et secundum munditiam manuum mearum reddet mihi
2SAM|22|22|quia custodivi vias Domini et non egi impie a Deo meo
2SAM|22|23|omnia enim iudicia eius in conspectu meo et praecepta eius non amovi a me
2SAM|22|24|et ero perfectus cum eo et custodiam me ab iniquitate mea
2SAM|22|25|et restituet Dominus mihi secundum iustitiam meam et secundum munditiam manuum mearum in conspectu oculorum suorum
2SAM|22|26|cum sancto sanctus eris et cum robusto perfectus
2SAM|22|27|cum electo electus eris et cum perverso perverteris
2SAM|22|28|et populum pauperem salvum facies oculisque tuis excelsos humiliabis
2SAM|22|29|quia tu lucerna mea Domine et Domine inluminabis tenebras meas
2SAM|22|30|in te enim curram accinctus in Deo meo transiliam murum
2SAM|22|31|Deus inmaculata via eius eloquium Domini igne examinatum scutum est omnium sperantium in se
2SAM|22|32|quis est deus praeter Dominum et quis fortis praeter Deum nostrum
2SAM|22|33|Deus qui accingit me fortitudine et conplanavit perfectam viam meam
2SAM|22|34|coaequans pedes meos cervis et super excelsa mea statuens me
2SAM|22|35|docens manus meas ad proelium et conponens quasi arcum aereum brachia mea
2SAM|22|36|dedisti mihi clypeum salutis tuae et mansuetudo mea multiplicavit me
2SAM|22|37|dilatabis gressus meos subtus me et non deficient tali mei
2SAM|22|38|persequar inimicos meos et conteram et non revertar donec consumam eos
2SAM|22|39|consumam eos et confringam ut non consurgant cadent sub pedibus meis
2SAM|22|40|accinxisti me fortitudine ad proelium incurvabis resistentes mihi sub me
2SAM|22|41|inimicos meos dedisti mihi dorsum odientes me et disperdam eos
2SAM|22|42|clamabunt et non erit qui salvet ad Dominum et non exaudiet eos
2SAM|22|43|delebo eos ut pulverem terrae quasi lutum platearum comminuam eos atque conpingam
2SAM|22|44|salvabis me a contradictionibus populi mei custodies in caput gentium populus quem ignoro serviet mihi
2SAM|22|45|filii alieni resistent mihi auditu auris oboedient mihi
2SAM|22|46|filii alieni defluxerunt et contrahentur in angustiis suis
2SAM|22|47|vivit Dominus et benedictus Deus meus et exaltabitur Deus fortis salutis meae
2SAM|22|48|Deus qui das vindictas mihi et deicis populos sub me
2SAM|22|49|qui educis me ab inimicis meis et a resistentibus mihi elevas me a viro iniquo liberabis me
2SAM|22|50|propterea confitebor tibi Domine in gentibus et nomini tuo cantabo
2SAM|22|51|magnificanti salutes regis sui et facienti misericordiam christo suo David et semini eius in sempiternum
2SAM|23|1|haec autem sunt verba novissima quae dixit David filius Isai dixit vir cui constitutum est de christo Dei Iacob egregius psalta Israhel
2SAM|23|2|spiritus Domini locutus est per me et sermo eius per linguam meam
2SAM|23|3|dixit Deus Israhel mihi locutus est Fortis Israhel dominator hominum iustus dominator in timore Dei
2SAM|23|4|sicut lux aurorae oriente sole mane absque nubibus rutilat et sicut pluviis germinat herba de terra
2SAM|23|5|nec tanta est domus mea apud Deum ut pactum aeternum iniret mecum firmum in omnibus atque munitum cuncta enim salus mea et omnis voluntas nec est quicquam ex ea quod non germinet
2SAM|23|6|praevaricatores autem quasi spinae evellentur universi quae non tolluntur manibus
2SAM|23|7|et si quis tangere voluerit eas armabitur ferro et ligno lanceato igneque succensae conburentur usque ad nihilum
2SAM|23|8|haec nomina fortium David Sedens in cathedra sapientissimus princeps inter tres ipse est quasi tenerrimus ligni vermiculus qui octingentos interfecit impetu uno
2SAM|23|9|post hunc Eleazar filius patrui eius Ahoi inter tres fortes qui erant cum David quando exprobraverunt Philisthim et congregati sunt illuc in proelium
2SAM|23|10|cumque ascendissent viri Israhel ipse stetit et percussit Philistheos donec deficeret manus eius et obrigesceret cum gladio fecitque Dominus salutem magnam in die illa et populus qui fugerat reversus est ad caesorum spolia detrahenda
2SAM|23|11|et post hunc Semma filius Age de Arari et congregati sunt Philisthim in statione erat quippe ibi ager plenus lente cumque fugisset populus a facie Philisthim
2SAM|23|12|stetit ille in medio agri et tuitus est eum percussitque Philistheos et fecit Dominus salutem magnam
2SAM|23|13|necnon ante descenderant tres qui erant principes inter triginta et venerant tempore messis ad David in speluncam Odollam castra autem Philisthim erant posita in valle Gigantum
2SAM|23|14|et David erat in praesidio porro statio Philisthinorum tunc erat in Bethleem
2SAM|23|15|desideravit igitur David et ait si quis mihi daret potum aquae de cisterna quae est in Bethleem iuxta portam
2SAM|23|16|inruperunt ergo tres fortes castra Philisthinorum et hauserunt aquam de cisterna Bethleem quae erat iuxta portam et adtulerunt ad David at ille noluit bibere sed libavit illam Domino
2SAM|23|17|dicens propitius mihi sit Dominus ne faciam hoc num sanguinem hominum istorum qui profecti sunt et animarum periculum bibam noluit ergo bibere haec fecerunt tres robustissimi
2SAM|23|18|Abisai quoque frater Ioab filius Sarviae princeps erat de tribus ipse est qui elevavit hastam suam contra trecentos quos interfecit nominatus in tribus
2SAM|23|19|et inter tres nobilior eratque eorum princeps sed usque ad tres primos non pervenerat
2SAM|23|20|et Banaias filius Ioiada viri fortissimi magnorum operum de Capsehel ipse percussit duos leones Moab et ipse descendit et percussit leonem in media cisterna diebus nivis
2SAM|23|21|ipse quoque interfecit virum aegyptium virum dignum spectaculo habentem in manu hastam itaque cum descendisset ad eum in virga vi extorsit hastam de manu Aegyptii et interfecit eum hasta sua
2SAM|23|22|haec fecit Banaias filius Ioiadae
2SAM|23|23|et ipse nominatus inter tres robustos qui erant inter triginta nobiliores verumtamen usque ad tres non pervenerat fecitque eum David sibi auricularium a secreto
2SAM|23|24|Asahel frater Ioab inter triginta Eleanan filius patrui eius de Bethleem
2SAM|23|25|Semma de Arari Helica de Arodi
2SAM|23|26|Helas de Felthi Hira filius Aces de Thecua
2SAM|23|27|Abiezer de Anathoth Mobonnai de Usathi
2SAM|23|28|Selmon Aohites Maharai Netophathites
2SAM|23|29|Heled filius Banaa et ipse Netophathites Hithai filius Ribai de Gebeeth filiorum Beniamin
2SAM|23|30|Banahi Aufrathonites Heddai de torrente Gaas
2SAM|23|31|Abialbon Arbathites Azmaveth de Beromi
2SAM|23|32|Eliaba de Salboni filii Iasen Ionathan
2SAM|23|33|Semma de Horodi Haiam filius Sarar Arorites
2SAM|23|34|Elifeleth filius Aasbai filii Maachathi Heliam filius Ahitofel Gelonites
2SAM|23|35|Esrai de Carmelo Farai de Arbi
2SAM|23|36|Igaal filius Nathan de Soba Bonni de Gaddi
2SAM|23|37|Selech de Ammoni Naharai Berothites armiger Ioab filii Sarviae
2SAM|23|38|Hira Hiethrites Gareb et ipse Hiethrites
2SAM|23|39|Urias Hettheus omnes triginta septem
2SAM|24|1|et addidit furor Domini irasci contra Israhel commovitque David in eis dicentem vade numera Israhel et Iudam
2SAM|24|2|dixitque rex ad Ioab principem exercitus sui perambula omnes tribus Israhel a Dan usque Bersabee et numerate populum ut sciam numerum eius
2SAM|24|3|dixitque Ioab regi adaugeat Dominus Deus tuus ad populum quantus nunc est iterumque centuplicet in conspectu domini mei regis sed quid sibi dominus meus rex vult in re huiuscemodi
2SAM|24|4|obtinuit autem sermo regis verba Ioab et principum exercitus egressusque est Ioab et principes militum a facie regis ut numerarent populum Israhel
2SAM|24|5|cumque pertransissent Iordanem venerunt in Aroer ad dextram urbis quae est in valle Gad
2SAM|24|6|et per Iazer transierunt in Galaad et in terram inferiorem Hodsi et venerunt in Dan silvestria circumeuntesque iuxta Sidonem
2SAM|24|7|transierunt propter moenia Tyri et omnem terram Hevei et Chananei veneruntque ad meridiem Iuda in Bersabee
2SAM|24|8|et lustrata universa terra adfuerunt post novem menses et viginti dies in Hierusalem
2SAM|24|9|dedit ergo Ioab numerum descriptionis populi regi et inventa sunt de Israhel octingenta milia virorum fortium qui educerent gladium et de Iuda quingenta milia pugnatorum
2SAM|24|10|percussit autem cor David eum postquam numeratus est populus et dixit David ad Dominum peccavi valde in hoc facto sed precor Domine ut transferas iniquitatem servi tui quia stulte egi nimis
2SAM|24|11|surrexit itaque David mane et sermo Domini factus est ad Gad propheten et videntem David dicens
2SAM|24|12|vade et loquere ad David haec dicit Dominus trium tibi datur optio elige unum quod volueris ex his ut faciam tibi
2SAM|24|13|cumque venisset Gad ad David nuntiavit ei dicens aut septem annis veniet tibi fames in terra tua aut tribus mensibus fugies adversarios tuos et illi persequentur aut certe tribus diebus erit pestilentia in terra tua nunc ergo delibera et vide quem respondeam ei qui me misit sermonem
2SAM|24|14|dixit autem David ad Gad artor nimis sed melius est ut incidam in manu Domini multae enim misericordiae eius sunt quam in manu hominis
2SAM|24|15|inmisitque Dominus pestilentiam in Israhel de mane usque ad tempus constitutum et mortui sunt ex populo a Dan usque Bersabee septuaginta milia virorum
2SAM|24|16|cumque extendisset manum angelus Dei super Hierusalem ut disperderet eam misertus est Dominus super adflictione et ait angelo percutienti populum sufficit nunc contine manum tuam erat autem angelus Domini iuxta aream Areuna Iebusei
2SAM|24|17|dixitque David ad Dominum cum vidisset angelum caedentem populum ego sum qui peccavi ego inique egi isti qui oves sunt quid fecerunt vertatur obsecro manus tua contra me et contra domum patris mei
2SAM|24|18|venit autem Gad ad David in die illa et dixit ei ascende constitue Domino altare in area Areuna Iebusei
2SAM|24|19|et ascendit David iuxta sermonem Gad quem praeceperat ei Dominus
2SAM|24|20|conspiciensque Areuna animadvertit regem et servos eius transire ad se
2SAM|24|21|et egressus adoravit regem prono vultu in terra et ait quid causae est ut veniat dominus meus rex ad servum suum cui David ait ut emam a te aream et aedificem altare Domino et cesset interfectio quae grassatur in populo
2SAM|24|22|et ait Areuna ad David accipiat et offerat dominus meus rex sicut ei placet habes boves in holocaustum et plaustrum et iuga boum in usum lignorum
2SAM|24|23|omnia dedit Areuna rex regi dixitque Areuna ad regem Dominus Deus tuus suscipiat votum tuum
2SAM|24|24|cui respondens rex ait nequaquam ut vis sed emam pretio a te et non offeram Domino Deo meo holocausta gratuita emit ergo David aream et boves argenti siclis quinquaginta
2SAM|24|25|et aedificavit ibi David altare Domino et obtulit holocausta et pacifica et repropitiatus est Dominus terrae et cohibita est plaga ab Israhel
1KGS|1|1|et rex David senuerat habebatque aetatis plurimos dies cumque operiretur vestibus non calefiebat
1KGS|1|2|dixerunt ergo ei servi sui quaeramus domino nostro regi adulescentulam virginem et stet coram rege et foveat eum dormiatque in sinu tuo et calefaciat dominum nostrum regem
1KGS|1|3|quaesierunt igitur adulescentulam speciosam in omnibus finibus Israhel et invenerunt Abisag Sunamitin et adduxerunt eam ad regem
1KGS|1|4|erat autem puella pulchra nimis dormiebatque cum rege et ministrabat ei rex vero non cognovit eam
1KGS|1|5|Adonias autem filius Aggith elevabatur dicens ego regnabo fecitque sibi currum et equites et quinquaginta viros qui ante eum currerent
1KGS|1|6|nec corripuit eum pater suus aliquando dicens quare hoc fecisti erat autem et ipse pulcher valde secundus natu post Absalom
1KGS|1|7|et sermo ei cum Ioab filio Sarviae et cum Abiathar sacerdote qui adiuvabant partes Adoniae
1KGS|1|8|Sadoc vero sacerdos et Banaias filius Ioiadae et Nathan propheta et Semei et Rhei et robur exercitus David non erat cum Adonia
1KGS|1|9|immolatis ergo Adonias arietibus et vitulis et universis pinguibus iuxta lapidem Zoheleth qui erat vicinus fonti Rogel vocavit universos fratres suos filios regis et omnes viros Iuda servos regis
1KGS|1|10|Nathan autem prophetam et Banaiam et robustos quosque et Salomonem fratrem suum non vocavit
1KGS|1|11|dixit itaque Nathan ad Bethsabee matrem Salomonis num audisti quod regnaverit Adonias filius Aggith et dominus noster David hoc ignorat
1KGS|1|12|nunc ergo veni accipe a me consilium et salva animam tuam filiique tui Salomonis
1KGS|1|13|vade et ingredere ad regem David et dic ei nonne tu domine mi rex iurasti mihi ancillae tuae dicens quod Salomon filius tuus regnabit post me et ipse sedebit in solio meo quare ergo regnavit Adonias
1KGS|1|14|et adhuc ibi te loquente cum rege ego veniam post te et conplebo sermones tuos
1KGS|1|15|ingressa est itaque Bethsabee ad regem in cubiculo rex autem senuerat nimis et Abisag Sunamitis ministrabat ei
1KGS|1|16|inclinavit se Bethsabee et adoravit regem ad quam rex quid tibi inquit vis
1KGS|1|17|quae respondens ait domine mi tu iurasti per Dominum Deum tuum ancillae tuae Salomon filius tuus regnabit post me et ipse sedebit in solio meo
1KGS|1|18|et ecce nunc Adonias regnavit te domine mi rex ignorante
1KGS|1|19|mactavit boves et pinguia quaeque et arietes plurimos et vocavit omnes filios regis Abiathar quoque sacerdotem et Ioab principem militiae Salomonem autem servum tuum non vocavit
1KGS|1|20|verumtamen domine mi rex in te oculi respiciunt totius Israhel ut indices eis qui sedere debeat in solio tuo domine mi rex post te
1KGS|1|21|eritque cum dormierit dominus meus rex cum patribus suis erimus ego et filius meus Salomon peccatores
1KGS|1|22|adhuc illa loquente cum rege Nathan prophetes venit
1KGS|1|23|et nuntiaverunt regi dicentes adest Nathan propheta cumque introisset ante conspectum regis et adorasset eum pronus in terram
1KGS|1|24|dixit Nathan domine mi rex tu dixisti Adonias regnet post me et ipse sedeat super thronum meum
1KGS|1|25|quia descendit hodie et immolavit boves et pinguia et arietes plurimos et vocavit universos filios regis et principes exercitus Abiathar quoque sacerdotem illisque vescentibus et bibentibus coram eo et dicentibus vivat rex Adonias
1KGS|1|26|me servum tuum et Sadoc sacerdotem et Banaiam filium Ioiadae et Salomonem famulum tuum non vocavit
1KGS|1|27|numquid a domino meo rege exivit hoc verbum et mihi non indicasti servo tuo qui sessurus esset super thronum domini mei regis post eum
1KGS|1|28|et respondit rex David dicens vocate ad me Bethsabee quae cum fuisset ingressa coram rege et stetisset ante eum
1KGS|1|29|iuravit rex et ait vivit Dominus qui eruit animam meam de omni angustia
1KGS|1|30|quia sicut iuravi tibi per Dominum Deum Israhel dicens Salomon filius tuus regnabit post me et ipse sedebit super solium meum pro me sic faciam hodie
1KGS|1|31|submissoque Bethsabee in terram vultu adoravit regem dicens vivat dominus meus rex David in aeternum
1KGS|1|32|dixit quoque rex David vocate mihi Sadoc sacerdotem et Nathan propheten et Banaiam filium Ioiadae qui cum ingressi fuissent coram rege
1KGS|1|33|dixit ad eos tollite vobiscum servos domini vestri et inponite Salomonem filium meum super mulam meam et ducite eum in Gion
1KGS|1|34|et unguat eum ibi Sadoc sacerdos et Nathan propheta in regem super Israhel et canetis bucina atque dicetis vivat rex Salomon
1KGS|1|35|et ascendetis post eum et veniet et sedebit super solium meum et ipse regnabit pro me illique praecipiam ut sit dux super Israhel et super Iudam
1KGS|1|36|et respondit Banaias filius Ioiadae regi dicens amen sic loquatur Dominus Deus domini mei regis
1KGS|1|37|quomodo fuit Dominus cum domino meo rege sic sit cum Salomone et sublimius faciat solium eius a solio domini mei regis David
1KGS|1|38|descendit ergo Sadoc sacerdos et Nathan propheta et Banaias filius Ioiadae et Cherethi et Felethi et inposuerunt Salomonem super mulam regis David et adduxerunt eum in Gion
1KGS|1|39|sumpsitque Sadoc sacerdos cornu olei de tabernaculo et unxit Salomonem et cecinerunt bucina et dixit omnis populus vivat rex Salomon
1KGS|1|40|et ascendit universa multitudo post eum et populus canentium tibiis et laetantium gaudio magno et insonuit terra ad clamorem eorum
1KGS|1|41|audivit autem Adonias et omnes qui invitati fuerant ab eo iamque convivium finitum erat sed et Ioab audita voce tubae ait quid sibi vult clamor civitatis tumultuantis
1KGS|1|42|adhuc illo loquente Ionathan filius Abiathar sacerdotis venit cui dixit Adonias ingredere quia vir fortis es et bona nuntians
1KGS|1|43|responditque Ionathan Adoniae nequaquam dominus enim noster rex David regem constituit Salomonem
1KGS|1|44|misitque cum eo Sadoc sacerdotem et Nathan prophetam et Banaiam filium Ioiadae et Cherethi et Felethi et inposuerunt eum super mulam regis
1KGS|1|45|unxeruntque eum Sadoc sacerdos et Nathan propheta regem in Gion et ascenderunt inde laetantes et insonuit civitas haec est vox quam audistis
1KGS|1|46|sed et Salomon sedit super solio regni
1KGS|1|47|et ingressi servi regis benedixerunt domino nostro regi David dicentes amplificet Deus nomen Salomonis super nomen tuum et magnificet thronum eius super thronum tuum et adoravit rex in lectulo suo
1KGS|1|48|insuper et haec locutus est benedictus Dominus Deus Israhel qui dedit hodie sedentem in solio meo videntibus oculis meis
1KGS|1|49|territi sunt ergo et surrexerunt omnes qui invitati fuerant ab Adonia et ivit unusquisque in viam suam
1KGS|1|50|Adonias autem timens Salomonem surrexit et abiit tenuitque cornu altaris
1KGS|1|51|et nuntiaverunt Salomoni dicentes ecce Adonias timens regem Salomonem tenuit cornu altaris dicens iuret mihi hodie rex Salomon quod non interficiat servum suum gladio
1KGS|1|52|dixitque Salomon si fuerit vir bonus non cadet ne unus quidem capillus eius in terram sin autem malum inventum fuerit in eo morietur
1KGS|1|53|misit ergo rex Salomon et eduxit eum ab altari et ingressus adoravit regem Salomonem dixitque ei Salomon vade in domum tuam
1KGS|2|1|adpropinquaverant autem dies David ut moreretur praecepitque Salomoni filio suo dicens
1KGS|2|2|ego ingredior viam universae terrae confortare et esto vir
1KGS|2|3|et observa custodias Domini Dei tui ut ambules in viis eius et custodias caerimonias eius et praecepta eius et iudicia et testimonia sicut scriptum est in lege Mosi ut intellegas universa quae facis et quocumque te verteris
1KGS|2|4|ut confirmet Dominus sermones suos quos locutus est de me dicens si custodierint filii tui viam suam et ambulaverint coram me in veritate in omni corde suo et in omni anima sua non auferetur tibi vir de solio Israhel
1KGS|2|5|tu quoque nosti quae fecerit mihi Ioab filius Sarviae quae fecerit duobus principibus exercitus Israhel Abner filio Ner et Amasa filio Iether quos occidit et effudit sanguinem belli in pace et posuit cruorem proelii in balteo suo qui erat circa lumbos eius et in calciamento suo quod erat in pedibus eius
1KGS|2|6|facies ergo iuxta sapientiam tuam et non deduces canitiem eius pacifice ad inferos
1KGS|2|7|sed et filiis Berzellai Galaaditis reddes gratiam eruntque comedentes in mensa tua occurrerunt enim mihi quando fugiebam a facie Absalom fratris tui
1KGS|2|8|habes quoque apud te Semei filium Gera filii Iemini de Baurim qui maledixit mihi maledictione pessima quando ibam ad Castra sed quia descendit mihi in occursum cum transirem Iordanem et iuravi ei per Dominum dicens non te interficiam gladio
1KGS|2|9|tu noli pati esse eum innoxium vir autem sapiens es et scies quae facias ei deducesque canos eius cum sanguine ad infernum
1KGS|2|10|dormivit igitur David cum patribus suis et sepultus est in civitate David
1KGS|2|11|dies autem quibus regnavit David super Israhel quadraginta anni sunt in Hebron regnavit septem annis in Hierusalem triginta tribus
1KGS|2|12|Salomon autem sedit super thronum David patris sui et firmatum est regnum eius nimis
1KGS|2|13|et ingressus est Adonias filius Aggith ad Bethsabee matrem Salomonis quae dixit ei pacificusne ingressus tuus qui respondit pacificus
1KGS|2|14|addiditque sermo mihi est ad te cui ait loquere et ille
1KGS|2|15|tu inquit nosti quia meum erat regnum et me proposuerat omnis Israhel sibi in regem sed translatum est regnum et factum est fratris mei a Domino enim constitutum est ei
1KGS|2|16|nunc ergo petitionem unam deprecor a te ne confundas faciem meam quae dixit ad eum loquere
1KGS|2|17|et ille ait precor ut dicas Salomoni regi neque enim negare tibi quicquam potest ut det mihi Abisag Sunamitin uxorem
1KGS|2|18|et ait Bethsabee bene ego loquar pro te regi
1KGS|2|19|venit ergo Bethsabee ad regem Salomonem ut loqueretur ei pro Adonia et surrexit rex in occursum eius adoravitque eam et sedit super thronum suum positus quoque est thronus matri regis quae sedit ad dexteram eius
1KGS|2|20|dixitque ei petitionem unam parvulam ego deprecor a te ne confundas faciem meam dixit ei rex pete mater mi neque enim fas est ut avertam faciem tuam
1KGS|2|21|quae ait detur Abisag Sunamitis Adoniae fratri tuo uxor
1KGS|2|22|responditque rex Salomon et dixit matri suae quare postulas Abisag Sunamitin Adoniae postula ei et regnum ipse est enim frater meus maior me et habet Abiathar sacerdotem et Ioab filium Sarviae
1KGS|2|23|iuravit itaque rex Salomon per Dominum dicens haec faciat mihi Deus et haec addat quia contra animam suam locutus est Adonias verbum hoc
1KGS|2|24|et nunc vivit Dominus qui firmavit me et conlocavit super solium David patris mei et qui fecit mihi domum sicut locutus est quia hodie occidetur Adonias
1KGS|2|25|misitque rex Salomon per manum Banaiae filii Ioiadae qui interfecit eum et mortuus est
1KGS|2|26|Abiathar quoque sacerdoti dixit rex vade in Anathot ad agrum tuum es quidem vir mortis sed hodie te non interficiam quia portasti arcam Domini Dei coram David patre meo et sustinuisti laborem in omnibus in quibus laboravit pater meus
1KGS|2|27|eiecit ergo Salomon Abiathar ut non esset sacerdos Domini ut impleretur sermo Domini quem locutus est super domum Heli in Silo
1KGS|2|28|venit autem nuntius ad Ioab quod Ioab declinasset post Adoniam et post Absalom non declinasset fugit ergo Ioab in tabernaculum Domini et adprehendit cornu altaris
1KGS|2|29|nuntiatumque est regi Salomoni quod fugisset Ioab in tabernaculum Domini et esset iuxta altare misitque Salomon Banaiam filium Ioiadae dicens vade interfice eum
1KGS|2|30|venit Banaias ad tabernaculum Domini et dixit ei haec dicit rex egredere qui ait non egrediar sed hic moriar renuntiavit Banaias regi sermonem dicens haec locutus est Ioab et haec respondit mihi
1KGS|2|31|dixitque ei rex fac sicut locutus est et interfice eum et sepeli et amovebis sanguinem innocentem qui effusus est a Ioab a me et a domo patris mei
1KGS|2|32|et reddat Dominus sanguinem eius super caput eius quia interfecit duos viros iustos melioresque se et occidit eos gladio patre meo David ignorante Abner filium Ner principem militiae Israhel et Amasa filium Iether principem exercitus Iuda
1KGS|2|33|et revertetur sanguis illorum in caput Ioab et in caput seminis eius in sempiternum David autem et semini eius et domui et throno illius sit pax usque in aeternum a Domino
1KGS|2|34|ascendit itaque Banaias filius Ioiadae et adgressus eum interfecit sepultusque est in domo sua in deserto
1KGS|2|35|et constituit rex Banaiam filium Ioiadae pro eo super exercitum et Sadoc sacerdotem posuit pro Abiathar
1KGS|2|36|misit quoque rex et vocavit Semei dixitque ei aedifica tibi domum in Hierusalem et habita ibi et non egredieris inde huc atque illuc
1KGS|2|37|quacumque autem die egressus fueris et transieris torrentem Cedron scito te interficiendum sanguis tuus erit super caput tuum
1KGS|2|38|dixitque Semei regi bonus sermo sicut locutus est dominus meus rex sic faciet servus tuus habitavit itaque Semei in Hierusalem diebus multis
1KGS|2|39|factum est autem post annos tres ut fugerent servi Semei ad Achis filium Maacha regem Geth nuntiatumque est Semei quod servi eius essent in Geth
1KGS|2|40|et surrexit Semei et stravit asinum suum ivitque in Geth ad Achis ad requirendos servos suos et adduxit eos de Geth
1KGS|2|41|nuntiatum est autem Salomoni quod isset Semei in Geth de Hierusalem et redisset
1KGS|2|42|et mittens vocavit eum dixitque illi nonne testificatus sum tibi per Dominum et praedixi tibi quacumque die egressus ieris huc et illuc scito te esse moriturum et respondisti mihi bonus sermo audivi
1KGS|2|43|quare ergo non custodisti iusiurandum Domini et praeceptum quod praeceperam tibi
1KGS|2|44|dixitque rex ad Semei tu nosti omne malum cuius tibi conscium est cor tuum quod fecisti David patri meo reddidit Dominus malitiam tuam in caput tuum
1KGS|2|45|et rex Salomon benedictus et thronus David erit stabilis coram Domino usque in sempiternum
1KGS|2|46|iussit itaque rex Banaiae filio Ioiadae qui egressus percussit eum et mortuus est
1KGS|3|1|confirmatum est igitur regnum in manu Salomonis et adfinitate coniunctus est Pharaoni regi Aegypti accepit namque filiam eius et adduxit in civitatem David donec conpleret aedificans domum suam et domum Domini et murum Hierusalem per circuitum
1KGS|3|2|et tamen populus immolabat in excelsis non enim aedificatum erat templum nomini Domini usque in die illo
1KGS|3|3|dilexit autem Salomon Dominum ambulans in praeceptis David patris sui excepto quod in excelsis immolabat et accendebat thymiama
1KGS|3|4|abiit itaque in Gabaon ut immolaret ibi illud quippe erat excelsum maximum mille hostias in holocaustum obtulit Salomon super altare illud in Gabaon
1KGS|3|5|apparuit Dominus Salomoni per somnium nocte dicens postula quod vis ut dem tibi
1KGS|3|6|et ait Salomon tu fecisti cum servo tuo David patre meo misericordiam magnam sicut ambulavit in conspectu tuo in veritate et iustitia et recto corde tecum custodisti ei misericordiam tuam grandem et dedisti ei filium sedentem super thronum eius sicut et hodie
1KGS|3|7|et nunc Domine Deus tu regnare fecisti servum tuum pro David patre meo ego autem sum puer parvus et ignorans egressum et introitum meum
1KGS|3|8|et servus tuus in medio est populi quem elegisti populi infiniti qui numerari et supputari non potest prae multitudine
1KGS|3|9|dabis ergo servo tuo cor docile ut iudicare possit populum tuum et discernere inter malum et bonum quis enim potest iudicare populum istum populum tuum hunc multum
1KGS|3|10|placuit ergo sermo coram Domino quod Salomon rem huiuscemodi postulasset
1KGS|3|11|et dixit Deus Salomoni quia postulasti verbum hoc et non petisti tibi dies multos nec divitias aut animam inimicorum tuorum sed postulasti tibi sapientiam ad discernendum iudicium
1KGS|3|12|ecce feci tibi secundum sermones tuos et dedi tibi cor sapiens et intellegens in tantum ut nullus ante te similis tui fuerit nec post te surrecturus sit
1KGS|3|13|sed et haec quae non postulasti dedi tibi divitias scilicet et gloriam ut nemo fuerit similis tui in regibus cunctis retro diebus
1KGS|3|14|si autem ambulaveris in viis meis et custodieris praecepta mea et mandata mea sicut ambulavit pater tuus longos faciam dies tuos
1KGS|3|15|igitur evigilavit Salomon et intellexit quod esset somnium cumque venisset Hierusalem stetit coram arca foederis Domini et obtulit holocausta et fecit victimas pacificas et grande convivium universis famulis suis
1KGS|3|16|tunc venerunt duae mulieres meretrices ad regem steteruntque coram eo
1KGS|3|17|quarum una ait obsecro mi domine ego et mulier haec habitabamus in domo una et peperi apud eam in cubiculo
1KGS|3|18|tertia vero die postquam ego peperi peperit et haec et eramus simul nullusque alius in domo nobiscum exceptis nobis duabus
1KGS|3|19|mortuus est autem filius mulieris huius nocte dormiens quippe oppressit eum
1KGS|3|20|et consurgens intempesta nocte silentio tulit filium meum de latere meo ancillae tuae dormientis et conlocavit in sinu suo suum autem filium qui erat mortuus posuit in sinu meo
1KGS|3|21|cumque surrexissem mane ut darem lac filio meo apparuit mortuus quem diligentius intuens clara luce deprehendi non esse meum quem genueram
1KGS|3|22|responditque altera mulier non est ita sed filius tuus mortuus est meus autem vivit e contrario illa dicebat mentiris filius quippe meus vivit et filius tuus mortuus est atque in hunc modum contendebant coram rege
1KGS|3|23|tunc rex ait haec dicit filius meus vivit et filius tuus mortuus est et ista respondit non sed filius tuus mortuus est et filius meus vivit
1KGS|3|24|dixit ergo rex adferte mihi gladium cumque adtulissent gladium coram rege
1KGS|3|25|dividite inquit infantem vivum in duas partes et date dimidiam partem uni et dimidiam partem alteri
1KGS|3|26|dixit autem mulier cuius filius erat vivus ad regem commota sunt quippe viscera eius super filio suo obsecro domine date illi infantem vivum et nolite interficere eum contra illa dicebat nec mihi nec tibi sit dividatur
1KGS|3|27|respondens rex ait date huic infantem vivum et non occidatur haec est mater eius
1KGS|3|28|audivit itaque omnis Israhel iudicium quod iudicasset rex et timuerunt regem videntes sapientiam Dei esse in eo ad faciendum iudicium
1KGS|4|1|erat autem rex Salomon regnans super omnem Israhel
1KGS|4|2|et hii principes quos habebat Azarias filius Sadoc sacerdos
1KGS|4|3|Helioreph et Ahia filii Sesa scribae Iosaphat filius Ahilud a commentariis
1KGS|4|4|Banaias filius Ioiadae super exercitum Sadoc autem et Abiathar sacerdotes
1KGS|4|5|Azarias filius Nathan super eos qui adsistebant regi Zabud filius Nathan sacerdos amicus regis
1KGS|4|6|et Ahisar praepositus domus et Adoniram filius Abda super tributa
1KGS|4|7|habebat autem Salomon duodecim praefectos super omnem Israhel qui praebebant annonam regi et domui eius per singulos enim menses in anno singuli necessaria ministrabant
1KGS|4|8|et haec nomina eorum Benhur in monte Ephraim
1KGS|4|9|Bendecar in Macces et in Salebbim et in Bethsemes et Helon Bethanan
1KGS|4|10|Benesed in Araboth ipsius erat Soccho et omnis terra Epher
1KGS|4|11|Benabinadab cuius omnis Nepthad Dor Tapheth filiam Salomonis habebat uxorem
1KGS|4|12|Bana filius Ahilud regebat Thanac et Mageddo et universam Bethsan quae est iuxta Sarthana subter Hiezrahel a Bethsan usque Abelmeula e regione Iecmaan
1KGS|4|13|Bengaber in Ramoth Galaad habebat Avothiair filii Manasse in Galaad ipse praeerat in omni regione Argob quae est in Basan sexaginta civitatibus magnis atque muratis quae habebant seras aereas
1KGS|4|14|Ahinadab filius Addo praeerat in Manaim
1KGS|4|15|Ahimaas in Nepthali sed et ipse habebat Basmath filiam Salomonis in coniugio
1KGS|4|16|Baana filius Usi in Aser et in Balod
1KGS|4|17|Iosaphat filius Pharue in Isachar
1KGS|4|18|Semei filius Hela in Beniamin
1KGS|4|19|Gaber filius Uri in terra Galaad in terra Seon regis Amorrei et Og regis Basan super omnia quae erant in illa terra
1KGS|4|20|Iuda et Israhel innumerabiles sicut harena maris in multitudine comedentes et bibentes atque laetantes
1KGS|4|21|Salomon autem erat in dicione sua habens omnia regna sicut a flumine terrae Philisthim usque ad terminum Aegypti offerentium sibi munera et servientium ei cunctis diebus vitae eius
1KGS|4|22|erat autem cibus Salomonis per dies singulos triginta chori similae et sexaginta chori farinae
1KGS|4|23|decem boves pingues et viginti boves pascuales et centum arietes excepta venatione cervorum caprearum atque bubalorum et avium altilium
1KGS|4|24|ipse enim obtinebat omnem regionem quae erat trans flumen quasi a Thapsa usque Gazam et cunctos reges illarum regionum et habebat pacem ex omni parte in circuitu
1KGS|4|25|habitabatque Iudas et Israhel absque timore ullo unusquisque sub vite sua et sub ficu sua a Dan usque Bersabee cunctis diebus Salomonis
1KGS|4|26|et habebat Salomon quadraginta milia praesepia equorum currulium et duodecim milia equestrium
1KGS|4|27|nutriebantque eos supradicti regis praefecti sed et necessaria mensae regis Salomonis cum ingenti cura praebebant in tempore suo
1KGS|4|28|hordeum quoque et paleas equorum et iumentorum deferebant in locum ubi erat rex iuxta constitutum sibi
1KGS|4|29|dedit quoque Deus sapientiam Salomoni et prudentiam multam nimis et latitudinem cordis quasi harenam quae est in litore maris
1KGS|4|30|et praecedebat sapientia Salomonis sapientiam omnium Orientalium et Aegyptiorum
1KGS|4|31|et erat sapientior cunctis hominibus sapientior Aethan Ezraita et Heman et Chalcal et Dorda filiis Maol et erat nominatus in universis gentibus per circuitum
1KGS|4|32|locutus est quoque Salomon tria milia parabolas et fuerunt carmina eius quinque et mille
1KGS|4|33|et disputavit super lignis a cedro quae est in Libano usque ad hysopum quae egreditur de pariete et disseruit de iumentis et volucribus et reptilibus et piscibus
1KGS|4|34|et veniebant de cunctis populis ad audiendam sapientiam Salomonis et ab universis regibus terrae qui audiebant sapientiam eius
1KGS|5|1|misit quoque Hiram rex Tyri servos suos ad Salomonem audivit enim quod ipsum unxissent regem pro patre eius quia amicus fuerat Hiram David omni tempore
1KGS|5|2|misit autem et Salomon ad Hiram dicens
1KGS|5|3|tu scis voluntatem David patris mei et quia non potuerit aedificare domum nomini Domini Dei sui propter bella inminentia per circuitum donec daret Dominus eos sub vestigio pedum eius
1KGS|5|4|nunc autem requiem dedit Deus meus mihi per circuitum non est Satan neque occursus malus
1KGS|5|5|quam ob rem cogito aedificare templum nomini Domini Dei mei sicut locutus est Dominus David patri meo dicens filius tuus quem dabo pro te super solium tuum ipse aedificabit domum nomini meo
1KGS|5|6|praecipe igitur ut praecidant mihi cedros de Libano et servi mei sint cum servis tuis mercedem autem servorum tuorum dabo tibi quamcumque praeceperis scis enim quoniam non est in populo meo vir qui noverit ligna caedere sicut Sidonii
1KGS|5|7|cum ergo audisset Hiram verba Salomonis laetatus est valde et ait benedictus Dominus hodie qui dedit David filium sapientissimum super populum hunc plurimum
1KGS|5|8|et misit Hiram ad Salomonem dicens audivi quaecumque mandasti mihi ego faciam omnem voluntatem tuam in lignis cedrinis et abiegnis
1KGS|5|9|servi mei deponent ea de Libano ad mare et ego conponam ea in ratibus in mari usque ad locum quem significaveris mihi et adplicabo ea ibi et tu tolles ea praebebisque necessaria mihi ut detur cibus domui meae
1KGS|5|10|itaque Hiram dabat Salomoni ligna cedrina et ligna abiegna iuxta omnem voluntatem eius
1KGS|5|11|Salomon autem praebebat Hiram viginti milia chororum tritici in cibum domui eius et viginti choros purissimi olei haec tribuebat Salomon Hiram per annos singulos
1KGS|5|12|dedit quoque Dominus sapientiam Salomoni sicut locutus est ei et erat pax inter Hiram et Salomonem et percusserunt foedus ambo
1KGS|5|13|legitque rex Salomon operas de omni Israhel et erat indictio triginta milia virorum
1KGS|5|14|mittebatque eos in Libanum decem milia per menses singulos vicissim ita ut duobus mensibus essent in domibus suis et Adoniram erat super huiuscemodi indictione
1KGS|5|15|fuerunt itaque Salomoni septuaginta milia eorum qui onera portabant et octoginta milia latomorum in monte
1KGS|5|16|absque praepositis qui praeerant singulis operibus numero trium milium et trecentorum praecipientium populo et his qui faciebant opus
1KGS|5|17|praecepitque rex ut tollerent lapides grandes lapides pretiosos in fundamentum templi et quadrarent eos
1KGS|5|18|quos dolaverunt cementarii Salomonis et cementarii Hiram porro Biblii praeparaverunt ligna et lapides ad aedificandam domum
1KGS|6|1|factum est igitur quadringentesimo et octogesimo anno egressionis filiorum Israhel de terra Aegypti in anno quarto mense zio ipse est mensis secundus regis Salomonis super Israhel aedificare coepit domum Domino
1KGS|6|2|domus autem quam aedificabat rex Salomon Domino habebat sexaginta cubitos in longitudine et viginti cubitos in latitudine et triginta cubitos in altitudine
1KGS|6|3|et porticus erat ante templum viginti cubitorum longitudinis iuxta mensuram latitudinis templi et habebat decem cubitos latitudinis ante faciem templi
1KGS|6|4|fecitque in templo fenestras obliquas
1KGS|6|5|et aedificavit super parietem templi tabulata per gyrum in parietibus domus per circuitum templi et oraculi et fecit latera in circuitu
1KGS|6|6|tabulatum quod subter erat quinque cubitos habebat latitudinis et medium tabulatum sex cubitorum latitudinis et tertium tabulatum septem habens cubitos latitudinis trabes autem posuit in domo per circuitum forinsecus ut non hererent muris templi
1KGS|6|7|domus autem cum aedificaretur lapidibus dedolatis atque perfectis aedificata est et malleus et securis et omne ferramentum non sunt audita in domo cum aedificaretur
1KGS|6|8|ostium lateris medii in parte erat domus dexterae et per cocleam ascendebant in medium cenaculum et a medio in tertium
1KGS|6|9|et aedificavit domum et consummavit eam texit quoque domum laquearibus cedrinis
1KGS|6|10|et aedificavit tabulatum super omnem domum quinque cubitis altitudinis et operuit domum lignis cedrinis
1KGS|6|11|et factus est sermo Domini ad Salomonem dicens
1KGS|6|12|domus haec quam aedificas si ambulaveris in praeceptis meis et iudicia mea feceris et custodieris omnia mandata mea gradiens per ea firmabo sermonem meum tibi quem locutus sum ad David patrem tuum
1KGS|6|13|et habitabo in medio filiorum Israhel et non derelinquam populum meum Israhel
1KGS|6|14|igitur aedificavit Salomon domum et consummavit eam
1KGS|6|15|et aedificavit parietes domus intrinsecus tabulatis cedrinis a pavimento domus usque ad summitatem parietum et usque ad laquearia operuit lignis intrinsecus et texit pavimentum domus tabulis abiegnis
1KGS|6|16|aedificavitque viginti cubitorum ad posteriorem partem templi tabulata cedrina a pavimento usque ad superiora et fecit interiorem domum oraculi in sanctum sanctorum
1KGS|6|17|porro quadraginta cubitorum erat ipsum templum pro foribus oraculi
1KGS|6|18|et cedro omnis domus intrinsecus vestiebatur habens tornaturas suas et iuncturas fabrefactas et celaturas eminentes omnia cedrinis tabulis vestiebantur nec omnino lapis apparere poterat in pariete
1KGS|6|19|oraculum autem in medio domus in interiori parte fecerat ut poneret ibi arcam foederis Domini
1KGS|6|20|porro oraculum habebat viginti cubitos longitudinis et viginti cubitos latitudinis et viginti cubitos altitudinis et operuit illud atque vestivit auro purissimo sed et altare vestivit cedro
1KGS|6|21|domum quoque ante oraculum operuit auro purissimo et adfixit lamminas clavis aureis
1KGS|6|22|nihilque erat in templo quod non auro tegeretur sed et totum altare oraculi texit auro
1KGS|6|23|et fecit in oraculo duo cherubin de lignis olivarum decem cubitorum altitudinis
1KGS|6|24|quinque cubitorum ala cherub una et quinque cubitorum ala cherub altera id est decem cubitos habentes a summitate alae usque ad alae alterius summitatem
1KGS|6|25|decem quoque cubitorum erat cherub secundus mensura pari et opus unum erat in duobus cherubin
1KGS|6|26|id est altitudinem habebat unus cherub decem cubitorum et similiter cherub secundus
1KGS|6|27|posuitque cherubin in medio templi interioris extendebant autem alas suas cherubin et tangebat ala una parietem et ala cherub secundi tangebat parietem alterum alae autem alterae in media parte templi se invicem contingebant
1KGS|6|28|texit quoque cherubin auro
1KGS|6|29|et omnes parietes templi per circuitum scalpsit variis celaturis et torno et fecit in eis cherubin et palmas et picturas varias quasi prominentes de pariete et egredientes
1KGS|6|30|sed et pavimentum domus texit auro intrinsecus et extrinsecus
1KGS|6|31|et in ingressu oraculi fecit ostiola de lignis olivarum postesque angulorum quinque
1KGS|6|32|et duo ostia de lignis olivarum et scalpsit in eis picturam cherubin et palmarum species et anaglyfa valde prominentia et texit ea auro et operuit tam cherubin quam palmas et cetera auro
1KGS|6|33|fecitque in introitum templi postes de lignis olivarum quadrangulatos
1KGS|6|34|et duo ostia de lignis abiegnis altrinsecus et utrumque ostium duplex erat et se invicem tenens aperiebatur
1KGS|6|35|et scalpsit cherubin et palmas et celaturas valde eminentes operuitque omnia lamminis aureis opere quadro ad regulam
1KGS|6|36|et aedificavit atrium interius tribus ordinibus lapidum politorum et uno ordine lignorum cedri
1KGS|6|37|anno quarto fundata est domus Domini in mense zio
1KGS|6|38|et in anno undecimo mense bul ipse est mensis octavus perfecta est domus in omni opere suo et in universis utensilibus aedificavitque eam annis septem
1KGS|7|1|domum autem suam aedificavit Salomon tredecim annis et ad perfectum usque perduxit
1KGS|7|2|aedificavit quoque domum saltus Libani centum cubitorum longitudinis et quinquaginta cubitorum latitudinis et triginta cubitorum altitudinis et quattuor deambulacra inter columnas cedrinas ligna quippe cedrina exciderat in columnas
1KGS|7|3|et tabulatis cedrinis vestivit totam cameram quae quadraginta quinque columnis sustentabatur unus autem ordo habebat columnas quindecim
1KGS|7|4|contra se invicem positas
1KGS|7|5|et e regione se respicientes aequali spatio inter columnas et super columnas quadrangulata ligna in cunctis aequalia
1KGS|7|6|et porticum columnarum fecit quinquaginta cubitorum longitudinis et triginta cubitorum latitudinis et alteram porticum in facie maioris porticus et columnas et epistylia super columnas
1KGS|7|7|porticum quoque solii in qua tribunal est fecit et texit lignis cedrinis a pavimento usque ad summitatem
1KGS|7|8|et domuncula in qua sedetur ad iudicandum erat in media porticu simili opere domum quoque fecit filiae Pharaonis quam uxorem duxerat Salomon tali opere quali et hanc porticum
1KGS|7|9|omnia lapidibus pretiosis qui ad normam quandam atque mensuram tam intrinsecus quam extrinsecus serrati erant a fundamento usque ad summitatem parietum et intrinsecus usque ad atrium maius
1KGS|7|10|fundamenta autem de lapidibus pretiosis lapidibus magnis decem sive octo cubitorum
1KGS|7|11|et desuper lapides pretiosi aequalis mensurae secti erant similiterque de cedro
1KGS|7|12|et atrium maius rotundum trium ordinum de lapidibus sectis et unius ordinis dolata cedro necnon et in atrio domus Domini interiori et in porticu domus
1KGS|7|13|misit quoque rex Salomon et tulit Hiram de Tyro
1KGS|7|14|filium mulieris viduae de tribu Nepthali patre Tyrio artificem aerarium et plenum sapientia et intellegentia et doctrina ad faciendum omne opus ex aere qui cum venisset ad regem Salomonem fecit omne opus eius
1KGS|7|15|et finxit duas columnas aereas decem et octo cubitorum altitudinis columnam unam et linea duodecim cubitorum ambiebat columnam utramque
1KGS|7|16|duo quoque capitella fecit quae ponerentur super capita columnarum fusili aere quinque cubitorum altitudinis capitellum unum et quinque cubitorum altitudinis capitellum alterum
1KGS|7|17|et quasi in modum retis et catenarum sibi invicem miro opere contextarum utrumque capitellum columnarum fusile erat septena versuum retiacula in capitello uno et septena retiacula in capitello altero
1KGS|7|18|et perfecit columnas et duos ordines per circuitum retiaculorum singulorum ut tegerent capitella quae erant super summitatem malogranatorum eodem modo fecit et capitello secundo
1KGS|7|19|capitella autem quae erant super capita columnarum quasi opere lilii fabricata erant in porticu quattuor cubitorum
1KGS|7|20|et rursum alia capitella in summitate columnarum desuper iuxta mensuram columnae contra retiacula malogranatorum autem ducenti ordines erant in circuitu capitelli secundi
1KGS|7|21|et statuit duas columnas in porticum templi cumque statuisset columnam dexteram vocavit eam nomine Iachin similiter erexit columnam secundam et vocavit nomen eius Booz
1KGS|7|22|et super capita columnarum opus in modum lilii posuit perfectumque est opus columnarum
1KGS|7|23|fecit quoque mare fusile decem cubitorum a labio usque ad labium rotundum in circuitu quinque cubitorum altitudo eius et resticula triginta cubitorum cingebat illud per circuitum
1KGS|7|24|et scalptura subter labium circumibat illud decem cubitis ambiens mare duo ordines scalpturarum histriatarum erant fusiles
1KGS|7|25|et stabat super duodecim boves e quibus tres respiciebant ad aquilonem et tres ad occidentem et tres ad meridiem et tres ad orientem et mare super eos desuper erat quorum posteriora universa intrinsecus latitabant
1KGS|7|26|grossitudo autem luteris trium unciarum erat labiumque eius quasi labium calicis et folium repandi lilii duo milia batos capiebat
1KGS|7|27|et fecit bases decem aereas quattuor cubitorum longitudinis bases singulas et quattuor cubitorum latitudinis et trium cubitorum altitudinis
1KGS|7|28|et ipsum opus basium interrasile erat et scalpturae inter iuncturas
1KGS|7|29|et inter coronulas et plectas leones et boves et cherubin et in iuncturis similiter desuper et subter leones et boves quasi lora ex aere dependentia
1KGS|7|30|et quattuor rotae per bases singulas et axes aerei et per quattuor partes quasi umeruli subter luterem fusiles contra se invicem respectantes
1KGS|7|31|os quoque luteris intrinsecus erat in capitis summitate et quod forinsecus apparebat unius cubiti erat totum rotundum pariterque habebat unum cubitum et dimidium in angulis autem columnarum variae celaturae erant et media intercolumnia quadrata non rotunda
1KGS|7|32|quattuor quoque rotae quae per quattuor angulos basis erant coherebant subter basi una rota habebat altitudinis cubitum et semis
1KGS|7|33|tales autem rotae erant quales solent in curru fieri et axes earum et radii et canti et modioli omnia fusilia
1KGS|7|34|nam et umeruli illi quattuor per singulos angulos basis unius ex ipsa basi fusiles et coniuncti erant
1KGS|7|35|in summitate autem basis erat quaedam rotunditas dimidii cubiti ita fabrefacta ut luter desuper possit inponi habens celaturas suas et scalpturas varias ex semet ipso
1KGS|7|36|scalpsit quoque in tabulatis illis quae erant ex aere et in angulis cherubin et leones et palmas quasi in similitudinem stantis hominis ut non celata sed adposita per circuitum viderentur
1KGS|7|37|in hunc modum fecit decem bases fusura una et mensura scalpturaque consimili
1KGS|7|38|fecit quoque decem luteres aereos quadraginta batos capiebat luter unus eratque quattuor cubitorum singulosque luteres per singulas id est decem bases posuit
1KGS|7|39|et constituit decem bases quinque ad dexteram partem templi et quinque ad sinistram mare autem posuit ad dexteram partem templi contra orientem ad meridiem
1KGS|7|40|fecit ergo Hiram lebetas et scutras et amulas et perfecit omne opus regis Salomonis in templo Domini
1KGS|7|41|columnas duas et funiculos capitulorum super capitella columnarum duos et retiacula duo ut operirent duos funiculos qui erant super capita columnarum
1KGS|7|42|et malogranata quadringenta in duobus retiaculis duos versus malogranatorum in retiaculis singulis ad operiendos funiculos capitellorum qui erant super capita columnarum
1KGS|7|43|et bases decem et luteres decem super bases
1KGS|7|44|et mare unum et boves duodecim subter mare
1KGS|7|45|et lebetas et scutras et amulas omnia vasa quae fecit Hiram regi Salomoni in domo Domini de aurichalco erant
1KGS|7|46|in campestri regione Iordanis fudit ea rex in argillosa terra inter Socchoth et Sarthan
1KGS|7|47|et posuit Salomon omnia vasa propter multitudinem autem nimiam non erat pondus aeris
1KGS|7|48|fecitque Salomon omnia vasa in domo Domini altare aureum et mensam super quam ponerentur panes propositionis auream
1KGS|7|49|et candelabra aurea quinque ad dexteram et quinque ad sinistram contra oraculum ex auro primo et quasi lilii flores et lucernas desuper aureas et forcipes aureos
1KGS|7|50|et hydrias et fuscinulas et fialas et mortariola et turibula de auro purissimo et cardines ostiorum domus interioris sancti sanctorum et ostiorum domus templi ex auro erant
1KGS|7|51|et perfecit omne opus quod faciebat Salomon in domo Domini et intulit quae sanctificaverat David pater suus argentum et aurum et vasa reposuitque in thesauris domus Domini
1KGS|8|1|tunc congregavit omnes maiores natu Israhel cum principibus tribuum et duces familiarum filiorum Israhel ad regem Salomonem in Hierusalem ut deferrent arcam foederis Domini de civitate David id est de Sion
1KGS|8|2|convenitque ad regem Salomonem universus Israhel in mense hethanim in sollemni die ipse est mensis septimus
1KGS|8|3|veneruntque cuncti senes ex Israhel et tulerunt sacerdotes arcam
1KGS|8|4|et portaverunt arcam Domini et tabernaculum foederis et omnia vasa sanctuarii quae erant in tabernaculo et ferebant ea sacerdotes et Levitae
1KGS|8|5|rex autem Salomon et omnis multitudo Israhel quae convenerat ad eum gradiebatur cum illo ante arcam et immolabant oves et boves absque aestimatione et numero
1KGS|8|6|et intulerunt sacerdotes arcam foederis Domini in locum suum in oraculum templi in sanctum sanctorum subter alas cherubin
1KGS|8|7|siquidem cherubin expandebant alas super locum arcae et protegebant arcam et vectes eius desuper
1KGS|8|8|cumque eminerent vectes et apparerent summitates eorum foris sanctuarium ante oraculum non apparebant ultra extrinsecus qui et fuerunt ibi usque in praesentem diem
1KGS|8|9|in arca autem non est aliud nisi duae tabulae lapideae quas posuerat in ea Moses in Horeb quando pepigit foedus Dominus cum filiis Israhel cum egrederentur de terra Aegypti
1KGS|8|10|factum est autem cum exissent sacerdotes de sanctuario nebula implevit domum Domini
1KGS|8|11|et non poterant sacerdotes stare et ministrare propter nebulam impleverat enim gloria Domini domum Domini
1KGS|8|12|tunc ait Salomon Dominus dixit ut habitaret in nebula
1KGS|8|13|aedificans aedificavi domum in habitaculum tuum firmissimum solium tuum in sempiternum
1KGS|8|14|convertitque rex faciem suam et benedixit omni ecclesiae Israhel omnis enim ecclesia Israhel stabat
1KGS|8|15|et ait benedictus Dominus Deus Israhel qui locutus est ore suo ad David patrem meum et in manibus eius perfecit dicens
1KGS|8|16|a die qua eduxi populum meum Israhel de Aegypto non elegi civitatem de universis tribubus Israhel ut aedificaretur domus et esset nomen meum ibi sed elegi David ut esset super populum meum Israhel
1KGS|8|17|voluitque David pater meus aedificare domum nomini Domini Dei Israhel
1KGS|8|18|et ait Dominus ad David patrem meum quod cogitasti in corde tuo aedificare domum nomini meo bene fecisti hoc ipsum mente tractans
1KGS|8|19|verumtamen tu non aedificabis domum sed filius tuus qui egredietur de renibus tuis ipse aedificabit domum nomini meo
1KGS|8|20|confirmavit Dominus sermonem suum quem locutus est stetique pro David patre meo et sedi super thronum Israhel sicut locutus est Dominus et aedificavi domum nomini Domini Dei Israhel
1KGS|8|21|et constitui ibi locum arcae in qua foedus est Domini quod percussit cum patribus nostris quando egressi sunt de terra Aegypti
1KGS|8|22|stetit autem Salomon ante altare Domini in conspectu ecclesiae Israhel et expandit manus suas in caelum
1KGS|8|23|et ait Domine Deus Israhel non est similis tui Deus in caelo desuper et super terra deorsum qui custodis pactum et misericordiam servis tuis qui ambulant coram te in toto corde suo
1KGS|8|24|qui custodisti servo tuo David patri meo quae locutus es ei ore locutus es et manibus perfecisti ut et haec dies probat
1KGS|8|25|nunc igitur Domine Deus Israhel conserva famulo tuo David patri meo quae locutus es ei dicens non auferetur de te vir coram me qui sedeat super thronum Israhel ita tamen si custodierint filii tui viam suam ut ambulent coram me sicut tu ambulasti in conspectu meo
1KGS|8|26|et nunc Deus Israhel firmentur verba tua quae locutus es servo tuo David patri meo
1KGS|8|27|ergone putandum est quod vere Deus habitet super terram si enim caelum et caeli caelorum te capere non possunt quanto magis domus haec quam aedificavi
1KGS|8|28|sed respice ad orationem servi tui et ad preces eius Domine Deus meus audi hymnum et orationem quam servus tuus orat coram te hodie
1KGS|8|29|ut sint oculi tui aperti super domum hanc nocte et die super domum de qua dixisti erit nomen meum ibi ut exaudias orationem qua orat te servus tuus in loco isto
1KGS|8|30|ut exaudias deprecationem servi tui et populi tui Israhel quodcumque oraverint in loco isto et exaudies in loco habitaculi tui in caelo et cum exaudieris propitius eris
1KGS|8|31|si peccaverit homo in proximum suum et habuerit aliquod iuramentum quo teneatur adstrictus et venerit propter iuramentum coram altari tuo in domum tuam
1KGS|8|32|tu exaudies in caelo et facies et iudicabis servos tuos condemnans impium et reddens viam suam super caput eius iustificansque iustum et retribuens ei secundum iustitiam suam
1KGS|8|33|si fugerit populus tuus Israhel inimicos suos quia peccaturus est tibi et agentes paenitentiam et confitentes nomini tuo venerint et oraverint et deprecati te fuerint in domo hac
1KGS|8|34|exaudi in caelo et dimitte peccatum populi tui Israhel et reduces eos in terram quam dedisti patribus eorum
1KGS|8|35|si clausum fuerit caelum et non pluerit propter peccata eorum et orantes in loco isto paenitentiam egerint nomini tuo et a peccatis suis conversi fuerint propter adflictionem suam
1KGS|8|36|exaudi eos in caelo et dimitte peccata servorum tuorum et populi tui Israhel et ostende eis viam bonam per quam ambulent et da pluviam super terram tuam quam dedisti populo tuo in possessionem
1KGS|8|37|fames si oborta fuerit in terra aut pestilentia aut corruptus aer aurugo lucusta rubigo et adflixerit eum et inimicus eius portas obsidens omnis plaga universa infirmitas
1KGS|8|38|cuncta devotatio et inprecatio quae acciderit omni homini de populo tuo Israhel si quis cognoverit plagam cordis sui et expanderit manus suas in domo hac
1KGS|8|39|tu audies in caelo in loco habitationis tuae et repropitiaberis et facies ut des unicuique secundum omnes vias suas sicut videris cor eius quia tu nosti solus cor omnium filiorum hominum
1KGS|8|40|ut timeant te cunctis diebus quibus vivunt super faciem terrae quam dedisti patribus nostris
1KGS|8|41|insuper et alienigena qui non est de populo tuo Israhel cum venerit de terra longinqua propter nomen tuum audietur enim nomen tuum magnum et manus tua fortis et brachium tuum
1KGS|8|42|extentum ubique cum venerit ergo et oraverit in loco hoc
1KGS|8|43|tu exaudies in caelo in firmamento habitaculi tui et facies omnia pro quibus invocaverit te alienigena ut discant universi populi terrarum nomen tuum timere sicut populus tuus Israhel et probent quia nomen tuum invocatum est super domum hanc quam aedificavi
1KGS|8|44|si egressus fuerit populus tuus ad bellum contra inimicos suos per viam quocumque miseris eos orabunt te contra viam civitatis quam elegisti et contra domum quam aedificavi nomini tuo
1KGS|8|45|et exaudies in caelo orationem eorum et preces eorum et facies iudicium eorum
1KGS|8|46|quod si peccaverint tibi non est enim homo qui non peccet et iratus tradideris eos inimicis suis et capti ducti fuerint in terram inimicorum longe vel prope
1KGS|8|47|et egerint paenitentiam in corde suo in loco captivitatis et conversi deprecati te fuerint in captivitate sua dicentes peccavimus inique egimus impie gessimus
1KGS|8|48|et reversi fuerint ad te in universo corde suo et tota anima sua in terra inimicorum suorum ad quam captivi ducti sunt et oraverint te contra viam terrae suae quam dedisti patribus eorum et civitatis quam elegisti et templi quod aedificavi nomini tuo
1KGS|8|49|exaudies in caelo in firmamento solii tui orationem eorum et preces et facies iudicium eorum
1KGS|8|50|et propitiaberis populo tuo qui peccavit tibi et omnibus iniquitatibus eorum quibus praevaricati sunt in te et dabis misericordiam coram eis qui eos captivos habuerint ut misereantur eis
1KGS|8|51|populus enim tuus est et hereditas tua quos eduxisti de terra Aegypti de medio fornacis ferreae
1KGS|8|52|ut sint oculi tui aperti ad deprecationem servi tui et populi tui Israhel et exaudias eos in universis pro quibus invocaverint te
1KGS|8|53|tu enim separasti eos tibi in hereditatem de universis populis terrae sicut locutus es per Mosen servum tuum quando eduxisti patres nostros de Aegypto Domine Deus
1KGS|8|54|factum est autem cum conplesset Salomon orans Dominum omnem orationem et deprecationem hanc surrexit de conspectu altaris Domini utrumque enim genu in terram fixerat et manus expanderat ad caelum
1KGS|8|55|stetit ergo et benedixit omni ecclesiae Israhel voce magna dicens
1KGS|8|56|benedictus Dominus qui dedit requiem populo suo Israhel iuxta omnia quae locutus est non cecidit ne unus quidem sermo ex omnibus bonis quae locutus est per Mosen servum suum
1KGS|8|57|sit Dominus Deus noster nobiscum sicut fuit cum patribus nostris non derelinquens nos neque proiciens
1KGS|8|58|sed inclinet corda nostra ad se ut ambulemus in universis viis eius et custodiamus mandata eius et caerimonias et iudicia quaecumque mandavit patribus nostris
1KGS|8|59|et sint sermones mei isti quibus deprecatus sum coram Domino adpropinquantes Domino Deo nostro die et nocte ut faciat iudicium servo suo et populo suo Israhel per singulos dies
1KGS|8|60|et sciant omnes populi terrae quia Dominus ipse est Deus et non est ultra absque eo
1KGS|8|61|sit quoque cor nostrum perfectum cum Domino Deo nostro ut ambulemus in decretis eius et custodiamus mandata eius sicut et hodie
1KGS|8|62|igitur rex et omnis Israhel cum eo immolabant victimas coram Domino
1KGS|8|63|mactavitque Salomon hostias pacificas quas immolavit Domino boum viginti duo milia ovium centum viginti milia et dedicaverunt templum Domini rex et filii Israhel
1KGS|8|64|in die illa sanctificavit rex medium atrii quod erat ante domum Domini fecit quippe ibi holocaustum et sacrificium et adipem pacificorum quia altare aereum quod erat coram Domino minus erat et capere non poterat holocausta et sacrificium et adipem pacificorum
1KGS|8|65|fecit ergo Salomon in tempore illo festivitatem celebrem et omnis Israhel cum eo multitudo magna ab introitu Emath usque ad rivum Aegypti coram Domino Deo nostro septem diebus et septem diebus id est quattuordecim diebus
1KGS|8|66|et in die octava dimisit populos qui benedicentes regi profecti sunt in tabernacula sua laetantes et alacri corde super omnibus bonis quae fecerat Dominus David servo suo et Israhel populo suo
1KGS|9|1|factum est autem cum perfecisset Salomon aedificium domus Domini et aedificium regis et omne quod optaverat et voluerat facere
1KGS|9|2|apparuit Dominus ei secundo sicut apparuerat ei in Gabaon
1KGS|9|3|dixitque Dominus ad eum exaudivi orationem tuam et deprecationem tuam qua deprecatus es coram me sanctificavi domum hanc quam aedificasti ut ponerem nomen meum ibi in sempiternum et erunt oculi mei et cor meum ibi cunctis diebus
1KGS|9|4|tu quoque si ambulaveris coram me sicut ambulavit pater tuus in simplicitate cordis et in aequitate et feceris omnia quae praecepi tibi et legitima mea et iudicia mea servaveris
1KGS|9|5|ponam thronum regni tui super Israhel in sempiternum sicut locutus sum David patri tuo dicens non auferetur de genere tuo vir de solio Israhel
1KGS|9|6|si autem aversione aversi fueritis vos et filii vestri non sequentes me nec custodientes mandata mea et caerimonias quas proposui vobis sed abieritis et colueritis deos alienos et adoraveritis eos
1KGS|9|7|auferam Israhel de superficie terrae quam dedi eis et templum quod sanctificavi nomini meo proiciam a conspectu meo eritque Israhel in proverbium et in fabulam cunctis populis
1KGS|9|8|et domus haec erit in exemplum omnis qui transierit per eam stupebit et sibilabit et dicet quare fecit Dominus sic terrae huic et domui huic
1KGS|9|9|et respondebunt quia dereliquerunt Dominum Deum suum qui eduxit patres eorum de terra Aegypti et secuti sunt deos alienos et adoraverunt eos et coluerunt idcirco induxit Dominus super eos omne malum hoc
1KGS|9|10|expletis autem annis viginti postquam aedificaverat Salomon duas domos id est domum Domini et domum regis
1KGS|9|11|Hiram rege Tyri praebente Salomoni ligna cedrina et abiegna et aurum iuxta omne quod opus habuerat tunc dedit Salomon Hiram viginti oppida in terra Galileae
1KGS|9|12|egressusque est Hiram de Tyro ut videret oppida quae dederat ei Salomon et non placuerunt ei
1KGS|9|13|et ait haecine sunt civitates quas dedisti mihi frater et appellavit eas terram Chabul usque in diem hanc
1KGS|9|14|misit quoque Hiram ad regem centum viginti talenta auri
1KGS|9|15|haec est summa expensarum quam obtulit rex Salomon ad aedificandam domum Domini et domum suam et Mello et murum Hierusalem et Eser et Mageddo et Gazer
1KGS|9|16|Pharao rex Aegypti ascendit et cepit Gazer succenditque eam igni et Chananeum qui habitabat in civitate interfecit et dedit eam in dote filiae suae uxori Salomonis
1KGS|9|17|aedificavit ergo Salomon Gazer et Bethoron inferiorem
1KGS|9|18|et Baalath et Palmyram in terra solitudinis
1KGS|9|19|et omnes vicos qui ad se pertinebant et erant absque muro munivit et civitates curruum et civitates equitum et quodcumque ei placuit ut aedificaret in Hierusalem et in Libano et in omni terra potestatis suae
1KGS|9|20|universum populum qui remanserat de Amorreis et Hettheis et Ferezeis et Eveis et Iebuseis qui non sunt de filiis Israhel
1KGS|9|21|horum filios qui remanserant in terra quos scilicet non potuerant filii Israhel exterminare fecit Salomon tributarios usque ad diem hanc
1KGS|9|22|de filiis autem Israhel non constituit Salomon servire quemquam sed erant viri bellatores et ministri eius et principes et duces et praefecti curruum et equorum
1KGS|9|23|erant autem principes super omnia opera Salomonis praepositi quingenti quinquaginta qui habebant subiectum populum et statutis operibus imperabant
1KGS|9|24|filia autem Pharaonis ascendit de civitate David in domum suam quam aedificaverat ei tunc aedificavit Mello
1KGS|9|25|offerebat quoque Salomon tribus vicibus per annos singulos holocausta et pacificas victimas super altare quod aedificaverat Domino et adolebat thymiama coram Domino perfectumque est templum
1KGS|9|26|classem quoque fecit rex Salomon in Asiongaber quae est iuxta Ahilam in litore maris Rubri in terra Idumea
1KGS|9|27|misitque Hiram in classe illa servos suos viros nauticos et gnaros maris cum servis Salomonis
1KGS|9|28|qui cum venissent in Ophir sumptum inde aurum quadringentorum viginti talentorum detulerunt ad regem Salomonem
1KGS|10|1|sed et regina Saba audita fama Salomonis in nomine Domini venit temptare eum in enigmatibus
1KGS|10|2|et ingressa Hierusalem multo comitatu et divitiis camelis portantibus aromata et aurum infinitum nimis et gemmas pretiosas venit ad Salomonem et locuta est ei universa quae habebat in corde suo
1KGS|10|3|et docuit eam Salomon omnia verba quae proposuerat non fuit sermo qui regem posset latere et non responderet ei
1KGS|10|4|videns autem regina Saba omnem sapientiam Salomonis et domum quam aedificaverat
1KGS|10|5|et cibos mensae eius et habitacula servorum et ordinem ministrantium vestesque eorum et pincernas et holocausta quae offerebat in domo Domini non habebat ultra spiritum
1KGS|10|6|dixitque ad regem verus est sermo quem audivi in terra mea
1KGS|10|7|super sermonibus tuis et super sapientia tua et non credebam narrantibus mihi donec ipsa veni et vidi oculis meis et probavi quod media pars mihi nuntiata non fuerit maior est sapientia et opera tua quam rumor quem audivi
1KGS|10|8|beati viri tui et beati servi tui hii qui stant coram te semper et audiunt sapientiam tuam
1KGS|10|9|sit Dominus Deus tuus benedictus cui placuisti et posuit te super thronum Israhel eo quod dilexerit Dominus Israhel in sempiternum et constituit te regem ut faceres iudicium et iustitiam
1KGS|10|10|dedit ergo regi centum viginti talenta auri et aromata multa nimis et gemmas pretiosas non sunt adlata ultra aromata tam multa quam ea quae dedit regina Saba regi Salomoni
1KGS|10|11|sed et classis Hiram quae portabat aurum de Ophir adtulit ex Ophir ligna thyina multa nimis et gemmas pretiosas
1KGS|10|12|fecitque rex de lignis thyinis fulchra domus Domini et domus regiae et citharas lyrasque cantoribus non sunt adlata huiuscemodi ligna thyina neque visa usque in praesentem diem
1KGS|10|13|rex autem Salomon dedit reginae Saba omnia quae voluit et petivit ab eo exceptis his quae ultro obtulerat ei munere regio quae reversa est et abiit in terram suam cum servis suis
1KGS|10|14|erat autem pondus auri quod adferebatur Salomoni per annos singulos sescentorum sexaginta sex talentorum auri
1KGS|10|15|excepto eo quod offerebant viri qui super vectigalia erant et negotiatores universique scruta vendentes et omnes reges Arabiae ducesque terrae
1KGS|10|16|fecit quoque rex Salomon ducenta scuta de auro puro sescentos auri siclos dedit in lamminas scuti unius
1KGS|10|17|et trecentas peltas ex auro probato trecentae minae auri unam peltam vestiebant posuitque ea rex in domo silvae Libani
1KGS|10|18|fecit etiam rex Salomon thronum de ebore grandem et vestivit eum auro fulvo nimis
1KGS|10|19|qui habebat sex gradus et summitas throni rotunda erat in parte posteriori et duae manus hinc atque inde tenentes sedile et duo leones stabant iuxta manus singulas
1KGS|10|20|et duodecim leunculi stantes super sex gradus hinc atque inde non est factum tale opus in universis regnis
1KGS|10|21|sed et omnia vasa de quibus potabat rex Salomon erant aurea et universa supellex domus saltus Libani de auro purissimo non erat argentum nec alicuius pretii putabatur in diebus Salomonis
1KGS|10|22|quia classis regis per mare cum classe Hiram semel per tres annos ibat in Tharsis deferens inde aurum et argentum dentes elefantorum et simias et pavos
1KGS|10|23|magnificatus est ergo rex Salomon super omnes reges terrae divitiis et sapientia
1KGS|10|24|et universa terra desiderabat vultum Salomonis ut audiret sapientiam eius quam dederat Deus in corde eius
1KGS|10|25|et singuli deferebant ei munera vasa argentea et aurea vestes et arma bellica aromata quoque et equos et mulos per annos singulos
1KGS|10|26|congregavitque Salomon currus et equites et facti sunt ei mille quadringenti currus et duodecim milia equitum et disposuit eos per civitates munitas et cum rege in Hierusalem
1KGS|10|27|fecitque ut tanta esset abundantia argenti in Hierusalem quanta lapidum et cedrorum praebuit multitudinem quasi sycomoros quae nascuntur in campestribus
1KGS|10|28|et educebantur equi Salomoni de Aegypto et de Coa negotiatores enim regis emebant de Coa et statuto pretio perducebant
1KGS|10|29|egrediebatur autem quadriga ex Aegypto sescentis siclis argenti et equus centum quinquaginta atque in hunc modum cuncti reges Hettheorum et Syriae equos venundabant
1KGS|11|1|rex autem Salomon amavit mulieres alienigenas multas filiam quoque Pharaonis et Moabitidas et Ammanitidas Idumeas et Sidonias et Chettheas
1KGS|11|2|de gentibus super quibus dixit Dominus filiis Israhel non ingrediemini ad eas neque de illis ingredientur ad vestras certissimo enim avertent corda vestra ut sequamini deos earum his itaque copulatus est Salomon ardentissimo amore
1KGS|11|3|fueruntque ei uxores quasi reginae septingentae et concubinae trecentae et averterunt mulieres cor eius
1KGS|11|4|cumque iam esset senex depravatum est per mulieres cor eius ut sequeretur deos alienos nec erat cor eius perfectum cum Domino Deo suo sicut cor David patris eius
1KGS|11|5|sed colebat Salomon Astharthen deam Sidoniorum et Moloch idolum Ammanitarum
1KGS|11|6|fecitque Salomon quod non placuerat coram Domino et non adimplevit ut sequeretur Dominum sicut pater eius
1KGS|11|7|tunc aedificavit Salomon fanum Chamos idolo Moab in monte qui est contra Hierusalem et Moloch idolo filiorum Ammon
1KGS|11|8|atque in hunc modum fecit universis uxoribus suis alienigenis quae adolebant tura et immolabant diis suis
1KGS|11|9|igitur iratus est Dominus Salomoni quod aversa esset mens eius a Domino Deo Israhel qui apparuerat ei secundo
1KGS|11|10|et praeceperat de verbo hoc ne sequeretur deos alienos et non custodivit quae mandavit ei Dominus
1KGS|11|11|dixit itaque Dominus Salomoni quia habuisti hoc apud te et non custodisti pactum meum et praecepta mea quae mandavi tibi disrumpens scindam regnum tuum et dabo illud servo tuo
1KGS|11|12|verumtamen in diebus tuis non faciam propter David patrem tuum de manu filii tui scindam illud
1KGS|11|13|nec totum regnum auferam sed tribum unam dabo filio tuo propter David servum meum et Hierusalem quam elegi
1KGS|11|14|suscitavit autem Dominus adversarium Salomoni Adad Idumeum de semine regio qui erat in Edom
1KGS|11|15|cum enim esset David in Idumea et ascendisset Ioab princeps militiae ad sepeliendos eos qui fuerant interfecti et occidisset omne masculinum in Idumea
1KGS|11|16|sex enim mensibus ibi moratus est Ioab et omnis Israhel donec interimerent omne masculinum in Idumea
1KGS|11|17|fugit Adad ipse et viri idumei de servis patris eius cum eo ut ingrederetur Aegyptum erat autem Adad puer parvulus
1KGS|11|18|cumque surrexissent de Madian venerunt in Pharan tuleruntque secum viros de Pharan et introierunt Aegyptum ad Pharaonem regem Aegypti qui dedit ei domum et cibos constituit et terram delegavit
1KGS|11|19|et invenit Adad gratiam coram Pharao valde in tantum ut daret ei uxorem sororem uxoris suae germanam Tafnes reginae
1KGS|11|20|genuitque ei soror Tafnes Genebath filium et nutrivit eum Tafnes in domo Pharaonis eratque Genebath habitans apud Pharaonem cum filiis eius
1KGS|11|21|cumque audisset Adad in Aegypto dormisse David cum patribus suis et mortuum esse Ioab principem militiae dixit Pharaoni dimitte me ut vadam in terram meam
1KGS|11|22|dixitque ei Pharao qua enim re apud me indiges ut quaeras ire ad terram tuam at ille respondit nulla sed obsecro ut dimittas me
1KGS|11|23|suscitavit quoque ei Deus adversarium Razon filium Heliada qui fugerat Adadezer regem Soba dominum suum
1KGS|11|24|et congregavit contra eum viros et factus est princeps latronum cum interficeret eos David abieruntque Damascum et habitaverunt ibi et constituerunt eum regem in Damasco
1KGS|11|25|eratque adversarius Israhel cunctis diebus Salomonis et hoc est malum Adad et odium contra Israhel regnavitque in Syria
1KGS|11|26|Hieroboam quoque filius Nabath Ephratheus de Sareda cuius mater erat nomine Sarva mulier vidua servus Salomonis levavit manum contra regem
1KGS|11|27|et haec causa rebellionis adversus eum quia Salomon aedificavit Mello et coaequavit voraginem civitatis David patris sui
1KGS|11|28|erat autem Hieroboam vir fortis et potens vidensque Salomon adulescentem bonae indolis et industrium constituerat eum praefectum super tributa universae domus Ioseph
1KGS|11|29|factum est igitur in tempore illo ut Hieroboam egrederetur de Hierusalem et inveniret eum Ahias Silonites propheta in via opertus pallio novo erant autem duo tantum in agro
1KGS|11|30|adprehendensque Ahia pallium suum novum quo opertus erat scidit in duodecim partes
1KGS|11|31|et ait ad Hieroboam tolle tibi decem scissuras haec enim dicit Dominus Deus Israhel ecce ego scindam regnum de manu Salomonis et dabo tibi decem tribus
1KGS|11|32|porro una tribus remanebit ei propter servum meum David et Hierusalem civitatem quam elegi ex omnibus tribubus Israhel
1KGS|11|33|eo quod dereliquerint me et adoraverint Astharoth deam Sidoniorum et Chamos deum Moab et Melchom deum filiorum Ammon et non ambulaverint in viis meis ut facerent iustitiam coram me et praecepta mea et iudicia sicut David pater eius
1KGS|11|34|nec auferam omne regnum de manu eius sed ducem ponam eum cunctis diebus vitae suae propter David servum meum quem elegi qui custodivit mandata mea et praecepta mea
1KGS|11|35|auferam autem regnum de manu filii eius et dabo tibi decem tribus
1KGS|11|36|filio autem eius dabo tribum unam ut remaneat lucerna David servo meo cunctis diebus coram me in Hierusalem civitatem quam elegi ut esset nomen meum ibi
1KGS|11|37|te autem adsumam et regnabis super omnia quae desiderat anima tua erisque rex super Israhel
1KGS|11|38|si igitur audieris omnia quae praecepero tibi et ambulaveris in viis meis et feceris quod rectum est coram me custodiens mandata mea et praecepta mea sicut fecit David servus meus ero tecum et aedificabo tibi domum fidelem quomodo aedificavi David et tradam tibi Israhel
1KGS|11|39|et adfligam semen David super hoc verumtamen non cunctis diebus
1KGS|11|40|voluit ergo Salomon interficere Hieroboam qui surrexit et aufugit in Aegyptum ad Susac regem Aegypti et fuit in Aegypto usque ad mortem Salomonis
1KGS|11|41|reliquum autem verborum Salomonis et omnia quae fecit et sapientia eius ecce universa scripta sunt in libro verborum Salomonis
1KGS|11|42|dies autem quos regnavit Salomon in Hierusalem super omnem Israhel quadraginta anni sunt
1KGS|11|43|dormivitque Salomon cum patribus suis et sepultus est in civitate David patris sui regnavitque Roboam filius eius pro eo
1KGS|12|1|venit autem Roboam in Sychem illuc enim congregatus erat omnis Israhel ad constituendum eum regem
1KGS|12|2|at Hieroboam filius Nabath cum adhuc esset in Aegypto profugus a facie regis Salomonis audita morte eius reversus est de Aegypto
1KGS|12|3|miseruntque et vocaverunt eum venit ergo Hieroboam et omnis multitudo Israhel et locuti sunt ad Roboam dicentes
1KGS|12|4|pater tuus durissimum iugum inposuit nobis tu itaque nunc inminue paululum de imperio patris tui durissimo et de iugo gravissimo quod inposuit nobis et serviemus tibi
1KGS|12|5|qui ait eis ite usque ad tertium diem et revertimini ad me cumque abisset populus
1KGS|12|6|iniit consilium rex Roboam cum senibus qui adsistebant coram Salomone patre eius dum adviveret et ait quod mihi datis consilium ut respondeam populo
1KGS|12|7|qui dixerunt ei si hodie oboedieris populo huic et servieris et petitioni eorum cesseris locutusque fueris ad eos verba lenia erunt tibi servi cunctis diebus
1KGS|12|8|qui dereliquit consilium senum quod dederant ei et adhibuit adulescentes qui nutriti fuerant cum eo et adsistebant illi
1KGS|12|9|dixitque ad eos quod mihi datis consilium ut respondeam populo huic qui dixerunt mihi levius fac iugum quod inposuit pater tuus super nos
1KGS|12|10|et dixerunt ei iuvenes qui nutriti fuerant cum eo sic loquere populo huic qui locuti sunt ad te dicentes pater tuus adgravavit iugum nostrum tu releva nos sic loqueris ad eos minimus digitus meus grossior est dorso patris mei
1KGS|12|11|et nunc pater meus posuit super vos iugum grave ego autem addam super iugum vestrum pater meus cecidit vos flagellis ego autem caedam scorpionibus
1KGS|12|12|venit ergo Hieroboam et omnis populus ad Roboam die tertia sicut locutus fuerat rex dicens revertimini ad me die tertia
1KGS|12|13|responditque rex populo dura derelicto consilio seniorum quod ei dederant
1KGS|12|14|et locutus est eis secundum consilium iuvenum dicens pater meus adgravavit iugum vestrum ego autem addam iugo vestro pater meus cecidit vos flagellis et ego caedam scorpionibus
1KGS|12|15|et non adquievit rex populo quoniam aversatus eum fuerat Dominus ut suscitaret verbum suum quod locutus fuerat in manu Ahiae Silonitae ad Hieroboam filium Nabath
1KGS|12|16|videns itaque populus quod noluisset eos audire rex respondit ei dicens quae nobis pars in David vel quae hereditas in filio Isai in tabernacula tua Israhel nunc vide domum tuam David et abiit Israhel in tabernacula sua
1KGS|12|17|super filios autem Israhel quicumque habitabant in civitatibus Iuda regnavit Roboam
1KGS|12|18|misit igitur rex Roboam Aduram qui erat super tributum et lapidavit eum omnis Israhel et mortuus est porro rex Roboam festinus ascendit currum et fugit in Hierusalem
1KGS|12|19|recessitque Israhel a domo David usque in praesentem diem
1KGS|12|20|factum est autem cum audisset omnis Israhel quod reversus esset Hieroboam miserunt et vocaverunt eum congregato coetu et constituerunt regem super omnem Israhel nec secutus est quisquam domum David praeter tribum Iuda solam
1KGS|12|21|venit autem Roboam Hierusalem et congregavit universam domum Iuda et tribum Beniamin centum octoginta milia electorum virorum et bellatorum ut pugnaret contra domum Israhel et reduceret regnum Roboam filio Salomonis
1KGS|12|22|factus est vero sermo Domini ad Semeiam virum Dei dicens
1KGS|12|23|loquere ad Roboam filium Salomonis regem Iuda et ad omnem domum Iuda et Beniamin et reliquos de populo dicens
1KGS|12|24|haec dicit Dominus non ascendetis nec bellabitis contra fratres vestros filios Israhel revertatur vir in domum suam a me enim factum est verbum hoc audierunt sermonem Domini et reversi sunt de itinere sicut eis praeceperat Dominus
1KGS|12|25|aedificavit autem Hieroboam Sychem in monte Ephraim et habitavit ibi et egressus inde aedificavit Phanuhel
1KGS|12|26|dixitque Hieroboam in corde suo nunc revertetur regnum ad domum David
1KGS|12|27|si ascenderit populus iste ut faciat sacrificia in domo Domini in Hierusalem et convertetur cor populi huius ad dominum suum Roboam regem Iuda interficientque me et revertentur ad eum
1KGS|12|28|et excogitato consilio fecit duos vitulos aureos et dixit eis nolite ultra ascendere Hierusalem ecce dii tui Israhel qui eduxerunt te de terra Aegypti
1KGS|12|29|posuitque unum in Bethel et alterum in Dan
1KGS|12|30|et factum est verbum hoc in peccatum ibat enim populus ad adorandum vitulum usque in Dan
1KGS|12|31|et fecit fana in excelsis et sacerdotes de extremis populi qui non erant de filiis Levi
1KGS|12|32|constituitque diem sollemnem in mense octavo quintadecima die mensis in similitudinem sollemnitatis quae celebratur in Iuda et ascendens altare similiter fecit in Bethel ut immolaret vitulis quos fabricatus erat constituitque in Bethel sacerdotes excelsorum quae fecerat
1KGS|12|33|et ascendit super altare quod extruxerat in Bethel quintadecima die mensis octavi quem finxerat de corde suo et fecit sollemnitatem filiis Israhel et ascendit super altare ut adoleret incensum
1KGS|13|1|et ecce vir Dei venit de Iuda in sermone Domini in Bethel Hieroboam stante super altare et tus iaciente
1KGS|13|2|et exclamavit contra altare in sermone Domini et ait altare altare haec dicit Dominus ecce filius nascetur domui David Iosias nomine et immolabit super te sacerdotes excelsorum qui nunc in te tura succendunt et ossa hominum incendet super te
1KGS|13|3|deditque in die illa signum dicens hoc erit signum quod locutus est Dominus ecce altare scinditur et effunditur cinis qui in eo est
1KGS|13|4|cumque audisset rex sermonem hominis Dei quem inclamaverat contra altare in Bethel extendit manum suam de altari dicens adprehendite eum et exaruit manus eius quam extenderat contra eum nec valuit retrahere eam ad se
1KGS|13|5|altare quoque scissum est et effusus cinis de altari iuxta signum quod praedixerat vir Dei in sermone Domini
1KGS|13|6|et ait rex ad virum Dei deprecare faciem Domini Dei tui et ora pro me ut restituatur manus mea mihi oravit vir Dei faciem Domini et reversa est manus regis ad eum et facta est sicut prius fuerat
1KGS|13|7|locutus est autem rex ad virum Dei veni mecum domum ut prandeas et dabo tibi munera
1KGS|13|8|responditque vir Dei ad regem si dederis mihi mediam partem domus tuae non veniam tecum nec comedam panem neque bibam aquam in loco isto
1KGS|13|9|sic enim mandatum est mihi in sermone Domini praecipientis non comedes panem neque bibes aquam nec reverteris per viam qua venisti
1KGS|13|10|abiit ergo per aliam viam et non est reversus per iter quo venerat in Bethel
1KGS|13|11|prophetes autem quidam senex habitabat in Bethel ad quem venit filius suus et narravit ei omnia opera quae fecerat vir Dei illa die in Bethel et verba quae locutus fuerat ad regem et narraverunt patri suo
1KGS|13|12|et dixit eis pater eorum per quam viam abiit ostenderunt ei filii sui viam per quam abierat vir Dei qui venerat de Iuda
1KGS|13|13|et ait filiis suis sternite mihi asinum qui cum stravissent ascendit
1KGS|13|14|et abiit post virum Dei et invenit eum sedentem subtus terebinthum et ait illi tune es vir Dei qui venisti de Iuda respondit ille ego sum
1KGS|13|15|dixit ad eum veni mecum domum ut comedas panem
1KGS|13|16|qui ait non possum reverti neque venire tecum nec comedam panem nec bibam aquam in loco isto
1KGS|13|17|quia locutus est Dominus ad me in sermone Domini dicens non comedes panem et non bibes ibi aquam nec reverteris per viam qua ieris
1KGS|13|18|qui ait illi et ego propheta sum similis tui et angelus locutus est mihi in sermone Domini dicens reduc eum tecum in domum tuam et comedat panem et bibat aquam fefellit eum
1KGS|13|19|et reduxit secum comedit ergo panem in domo eius et bibit aquam
1KGS|13|20|cumque sederent ad mensam factus est sermo Domini ad prophetam qui reduxerat eum
1KGS|13|21|et exclamavit ad virum Dei qui venerat de Iuda dicens haec dicit Dominus quia inoboediens fuisti ori Domini et non custodisti mandatum quod praecepit tibi Dominus Deus tuus
1KGS|13|22|et reversus es et comedisti panem et bibisti aquam in loco in quo praecepit tibi ne comederes panem neque biberes aquam non inferetur cadaver tuum in sepulchrum patrum tuorum
1KGS|13|23|cumque comedisset et bibisset stravit asinum prophetae quem reduxerat
1KGS|13|24|qui cum abisset invenit eum leo in via et occidit et erat cadaver eius proiectum in itinere asinus autem stabat iuxta illum et leo stabat iuxta cadaver
1KGS|13|25|et ecce viri transeuntes viderunt cadaver proiectum in via et leonem stantem iuxta cadaver et venerunt et divulgaverunt in civitate in qua prophetes senex ille habitabat
1KGS|13|26|quod cum audisset propheta ille qui reduxerat eum de via ait vir Dei est qui inoboediens fuit ori Domini et tradidit eum Dominus leoni et confregit eum et occidit iuxta verbum Domini quod locutus est ei
1KGS|13|27|dixitque ad filios suos sternite mihi asinum qui cum stravissent
1KGS|13|28|et ille abisset invenit cadaver eius proiectum in via et asinum et leonem stantes iuxta cadaver non comedit leo de cadavere nec laesit asinum
1KGS|13|29|tulit ergo prophetes cadaver viri Dei et posuit illud super asinum et reversus intulit in civitatem prophetae senis ut plangerent eum
1KGS|13|30|et posuit cadaver eius in sepulchro suo et planxerunt eum heu frater
1KGS|13|31|cumque planxissent eum dixit ad filios suos cum mortuus fuero sepelite me in sepulchro in quo vir Dei sepultus est iuxta ossa eius ponite ossa mea
1KGS|13|32|profecto enim veniet sermo quem praedixit in sermone Domini contra altare quod est in Bethel et contra omnia fana excelsorum quae sunt in urbibus Samariae
1KGS|13|33|post verba haec non est reversus Hieroboam de via sua pessima sed e contrario fecit de novissimis populi sacerdotes excelsorum quicumque volebat implebat manum suam et fiebat sacerdos excelsorum
1KGS|13|34|et propter hanc causam peccavit domus Hieroboam et eversa est et deleta de superficie terrae
1KGS|14|1|in tempore illo aegrotavit Abia filius Hieroboam
1KGS|14|2|dixitque Hieroboam uxori suae surge et commuta habitum ne cognoscaris quod sis uxor Hieroboam et vade in Silo ubi est Ahia propheta qui locutus est mihi quod regnaturus essem super populum hunc
1KGS|14|3|tolle quoque in manu tua decem panes et crustula et vas mellis et vade ad illum ipse indicabit tibi quid eventurum sit huic puero
1KGS|14|4|fecit ut dixerat uxor Hieroboam et consurgens abiit in Silo et venit in domum Ahia at ille non poterat videre quia caligaverant oculi eius prae senectute
1KGS|14|5|dixit autem Dominus ad Ahiam ecce uxor Hieroboam ingreditur ut consulat te super filio suo qui aegrotat haec et haec loqueris ei cum ergo illa intraret et dissimularet se esse quae erat
1KGS|14|6|audivit Ahias sonitum pedum eius introeuntis per ostium et ait ingredere uxor Hieroboam quare aliam esse te simulas ego autem missus sum ad te durus nuntius
1KGS|14|7|vade et dic Hieroboam haec dicit Dominus Deus Israhel quia exaltavi te de medio populi et dedi te ducem super populum meum Israhel
1KGS|14|8|et scidi regnum domus David et dedi illud tibi et non fuisti sicut servus meus David qui custodivit mandata mea et secutus est me in toto corde suo faciens quod placitum esset in conspectu meo
1KGS|14|9|sed operatus es male super omnes qui fuerunt ante te et fecisti tibi deos alienos et conflatiles ut me ad iracundiam provocares me autem proiecisti post corpus tuum
1KGS|14|10|idcirco ecce ego inducam mala super domum Hieroboam et percutiam de Hieroboam mingentem ad parietem et clausum et novissimum in Israhel et mundabo reliquias domus Hieroboam sicut mundari solet fimus usque ad purum
1KGS|14|11|qui mortui fuerint de Hieroboam in civitate comedent eos canes qui autem mortui fuerint in agro vorabunt eos aves caeli quia Dominus locutus est
1KGS|14|12|tu igitur surge et vade in domum tuam et in ipso introitu pedum tuorum in urbem morietur puer
1KGS|14|13|et planget eum omnis Israhel et sepeliet iste enim solus infertur de Hieroboam in sepulchrum quia inventus est super eo sermo bonus ad Dominum Deum Israhel in domo Hieroboam
1KGS|14|14|constituet autem sibi Dominus regem super Israhel qui percutiat domum Hieroboam in hac die et in hoc tempore
1KGS|14|15|et percutiet Dominus Israhel sicut moveri solet harundo in aqua et evellet Israhel de terra bona hac quam dedit patribus eorum et ventilabit eos trans Flumen quia fecerunt sibi lucos ut inritarent Dominum
1KGS|14|16|et tradet Dominus Israhel propter peccata Hieroboam qui peccavit et peccare fecit Israhel
1KGS|14|17|surrexit itaque uxor Hieroboam et abiit et venit in Thersa cumque illa ingrederetur limen domus puer mortuus est
1KGS|14|18|et sepelierunt eum et planxit illum omnis Israhel iuxta sermonem Domini quem locutus est in manu servi sui Ahiae prophetae
1KGS|14|19|reliqua autem verborum Hieroboam quomodo pugnaverit et quomodo regnaverit ecce scripta sunt in libro verborum dierum regum Israhel
1KGS|14|20|dies autem quibus regnavit Hieroboam viginti duo anni sunt et dormivit cum patribus suis regnavitque Nadab filius eius pro eo
1KGS|14|21|porro Roboam filius Salomonis regnavit in Iuda quadraginta et unius anni erat Roboam cum regnare coepisset et decem et septem annis regnavit in Hierusalem civitatem quam elegit Dominus ut poneret nomen suum ibi ex omnibus tribubus Israhel nomen autem matris eius Naama Ammanites
1KGS|14|22|et fecit Iudas malum coram Domino et inritaverunt eum super omnibus quae fecerant patres eorum in peccatis suis quae peccaverant
1KGS|14|23|aedificaverunt enim et ipsi sibi aras et statuas et lucos super omnem collem excelsum et subter omnem arborem frondosam
1KGS|14|24|sed et effeminati fuerunt in terra feceruntque omnes abominationes gentium quas adtrivit Dominus ante faciem filiorum Israhel
1KGS|14|25|in quinto autem anno regni Roboam ascendit Sesac rex Aegypti in Hierusalem
1KGS|14|26|et tulit thesauros domus Domini et thesauros regios et universa diripuit scuta quoque aurea quae fecerat Salomon
1KGS|14|27|pro quibus fecit rex Roboam scuta aerea et tradidit ea in manu ducum scutariorum et eorum qui excubabant ante ostium domus regis
1KGS|14|28|cumque ingrederetur rex in domum Domini portabant ea qui praeeundi habebant officium et postea reportabant ad armamentarium scutariorum
1KGS|14|29|reliqua autem sermonum Roboam et omnium quae fecit ecce scripta sunt in libro verborum dierum regum Iuda
1KGS|14|30|fuitque bellum inter Roboam et Hieroboam cunctis diebus
1KGS|14|31|dormivit itaque Roboam cum patribus suis et sepultus est cum eis in civitate David nomen autem matris eius Naama Ammanites et regnavit Abiam filius eius pro eo
1KGS|15|1|igitur in octavodecimo anno regni Hieroboam filii Nabath regnavit Abiam super Iudam
1KGS|15|2|tribus annis regnavit in Hierusalem nomen matris eius Maacha filia Absalom
1KGS|15|3|ambulavitque in omnibus peccatis patris sui quae fecerat ante eum nec erat cor eius perfectum cum Domino Deo suo sicut cor David patris eius
1KGS|15|4|sed propter David dedit ei Dominus Deus suus lucernam in Hierusalem ut suscitaret filium eius post eum et staret Hierusalem
1KGS|15|5|eo quod fecisset David rectum in oculis Domini et non declinasset ab omnibus quae praeceperat ei cunctis diebus vitae suae excepto sermone Uriae Hetthei
1KGS|15|6|attamen bellum fuit inter Roboam et inter Hieroboam omni tempore vitae eius
1KGS|15|7|reliqua autem sermonum Abiam et omnia quae fecit nonne haec scripta sunt in libro verborum dierum regum Iuda fuitque proelium inter Abiam et inter Hieroboam
1KGS|15|8|et dormivit Abiam cum patribus suis et sepelierunt eum in civitate David regnavitque Asa filius eius pro eo
1KGS|15|9|in anno ergo vicesimo Hieroboam regis Israhel regnavit Asa rex Iuda
1KGS|15|10|et quadraginta uno anno regnavit in Hierusalem nomen matris eius Maacha filia Absalom
1KGS|15|11|et fecit Asa rectum ante conspectum Domini sicut David pater eius
1KGS|15|12|et abstulit effeminatos de terra purgavitque universas sordes idolorum quae fecerant patres eius
1KGS|15|13|insuper et Maacham matrem suam amovit ne esset princeps in sacris Priapi et in luco eius quem consecraverat subvertitque specum eius et confregit simulacrum turpissimum et conbusit in torrente Cedron
1KGS|15|14|excelsa autem non abstulit verumtamen cor Asa perfectum erat cum Deo cunctis diebus suis
1KGS|15|15|et intulit ea quae sanctificaverat pater suus et voverat in domum Domini argentum et aurum et vasa
1KGS|15|16|bellum autem erat inter Asa et Baasa regem Israhel cunctis diebus eorum
1KGS|15|17|ascendit quoque Baasa rex Israhel in Iudam et aedificavit Rama ut non possit quispiam egredi vel ingredi de parte Asa regis Iudae
1KGS|15|18|tollens itaque Asa omne argentum et aurum quod remanserat in thesauris domus Domini et in thesauris domus regiae dedit illud in manu servorum suorum et misit ad Benadad filium Tabremmon filii Ezion regem Syriae qui habitabat in Damasco dicens
1KGS|15|19|foedus est inter me et te et inter patrem meum et patrem tuum ideo misi tibi munera argentum et aurum et peto ut venias et irritum facias foedus quod habes cum Baasa rege Israhel et recedat a me
1KGS|15|20|adquiescens Benadad regi Asa misit principes exercitus sui in civitates Israhel et percusserunt Ahion et Dan et Abel domum Maacha et universam Cenneroth omnem scilicet terram Nepthalim
1KGS|15|21|quod cum audisset Baasa intermisit aedificare Rama et reversus est in Thersa
1KGS|15|22|rex autem Asa nuntium misit in omnem Iudam nemo sit excusatus et tulerunt lapides Rama et ligna eius quibus aedificaverat Baasa et extruxit de eis rex Asa Gaba Beniamin et Maspha
1KGS|15|23|reliqua autem omnium sermonum Asa et universae fortitudines eius et cuncta quae fecit et civitates quas extruxit nonne haec scripta sunt in libro verborum dierum regum Iuda verumtamen in tempore senectutis suae doluit pedes
1KGS|15|24|et dormivit cum patribus suis et sepultus est cum eis in civitate David patris sui regnavitque Iosaphat filius eius pro eo
1KGS|15|25|Nadab vero filius Hieroboam regnavit super Israhel anno secundo Asa regis Iuda regnavitque super Israhel duobus annis
1KGS|15|26|et fecit quod malum est in conspectu Domini et ambulavit in viis patris sui et in peccatis eius quibus peccare fecit Israhel
1KGS|15|27|insidiatus est autem ei Baasa filius Ahia de domo Isachar et percussit eum in Gebbethon quae est urbs Philisthinorum siquidem Nadab et omnis Israhel obsidebant Gebbethon
1KGS|15|28|interfecit igitur illum Baasa in anno tertio Asa regis Iuda et regnavit pro eo
1KGS|15|29|cumque regnasset percussit omnem domum Hieroboam non dimisit ne unam quidem animam de semine eius donec deleret eum iuxta verbum Domini quod locutus fuerat in manu servi sui Ahiae Silonitis
1KGS|15|30|propter peccata Hieroboam quae peccaverat et quibus peccare fecerat Israhel et propter delictum quo inritaverat Dominum Deum Israhel
1KGS|15|31|reliqua autem sermonum Nadab et omnia quae operatus est nonne haec scripta sunt in libro verborum dierum regum Israhel
1KGS|15|32|fuitque bellum inter Asa et Baasa regem Israhel cunctis diebus eorum
1KGS|15|33|anno tertio Asa regis Iuda regnavit Baasa filius Ahia super omnem Israhel in Thersa viginti quattuor annis
1KGS|15|34|et fecit malum coram Domino ambulavitque in via Hieroboam et in peccatis eius quibus peccare fecit Israhel
1KGS|16|1|factus est autem sermo Domini ad Hieu filium Anani contra Baasa dicens
1KGS|16|2|pro eo quod exaltavi te de pulvere et posui ducem super populum meum Israhel tu autem ambulasti in via Hieroboam et peccare fecisti populum meum Israhel ut me inritares in peccatis eorum
1KGS|16|3|ecce ego demetam posteriora Baasa et posteriora domus eius et faciam domum tuam sicut domum Hieroboam filii Nabath
1KGS|16|4|qui mortuus fuerit de Baasa in civitate comedent eum canes et qui mortuus fuerit ex eo in regione comedent eum volucres caeli
1KGS|16|5|reliqua autem sermonum Baasa et quaecumque fecit et proelia eius nonne haec scripta sunt in libro verborum dierum regum Israhel
1KGS|16|6|dormivit ergo Baasa cum patribus suis sepultusque est in Thersa et regnavit Hela filius eius pro eo
1KGS|16|7|cum autem in manu Hieu filii Anani prophetae verbum Domini factum esset contra Baasa et contra domum eius et contra omne malum quod fecerat coram Domino ad inritandum eum in operibus manuum suarum ut fieret sicut domus Hieroboam ob hanc causam occidit eum
1KGS|16|8|anno vicesimo sexto Asa regis Iuda regnavit Hela filius Baasa super Israhel in Thersa duobus annis
1KGS|16|9|et rebellavit contra eum servus suus Zamri dux mediae partis equitum erat autem Hela in Thersa bibens et temulentus in domo Arsa praefecti Thersa
1KGS|16|10|inruens ergo Zamri percussit et occidit eum anno vicesimo septimo Asa regis Iuda et regnavit pro eo
1KGS|16|11|cumque regnasset et sedisset super solium eius percussit omnem domum Baasa et non dereliquit ex eo mingentem ad parietem et propinquos et amicos eius
1KGS|16|12|delevitque Zamri omnem domum Baasa iuxta verbum Domini quod locutus fuerat ad Baasa in manu Hieu prophetae
1KGS|16|13|propter universa peccata Baasa et peccata Hela filii eius qui peccaverunt et peccare fecerunt Israhel provocantes Dominum Deum Israhel in vanitatibus suis
1KGS|16|14|reliqua autem sermonum Hela et omnia quae fecit nonne haec scripta sunt in libro verborum dierum regum Israhel
1KGS|16|15|anno vicesimo et septimo Asa regis Iuda regnavit Zamri septem diebus in Thersa porro exercitus obsidebat Gebbethon urbem Philisthinorum
1KGS|16|16|cumque audisset rebellasse Zamri et occidisse regem fecit sibi regem omnis Israhel Amri qui erat princeps militiae super Israhel in die illa in castris
1KGS|16|17|ascendit ergo Amri et omnis Israhel cum eo de Gebbethon et obsidebant Thersa
1KGS|16|18|videns autem Zamri quod expugnanda esset civitas ingressus est palatium et succendit secum domum regiam et mortuus est
1KGS|16|19|in peccatis suis quae peccaverat faciens malum coram Domino et ambulans in via Hieroboam et in peccato eius quo fecit peccare Israhel
1KGS|16|20|reliqua autem sermonum Zamri et insidiarum eius et tyrannidis nonne haec scripta sunt in libro verborum dierum regum Israhel
1KGS|16|21|tunc divisus est populus Israhel in duas partes media pars populi sequebatur Thebni filium Gineth ut constitueret eum regem et media pars Amri
1KGS|16|22|praevaluit autem populus qui erat cum Amri populo qui sequebatur Thebni filium Gineth mortuusque est Thebni et regnavit Amri
1KGS|16|23|anno tricesimo primo Asa regis Iuda regnavit Amri super Israhel duodecim annis in Thersa regnavit sex annis
1KGS|16|24|emitque montem Samariae a Somer duobus talentis argenti et aedificavit eam et vocavit nomen civitatis quam extruxerat nomine Somer domini montis Samariae
1KGS|16|25|fecit autem Amri malum in conspectu Domini et operatus est nequiter super omnes qui fuerant ante eum
1KGS|16|26|ambulavitque in omni via Hieroboam filii Nabath et in peccatis eius quibus peccare fecerat Israhel ut inritaret Dominum Deum Israhel in vanitatibus suis
1KGS|16|27|reliqua autem sermonum Amri et proelia eius quae gessit nonne haec scripta sunt in libro verborum dierum regum Israhel
1KGS|16|28|et dormivit Amri cum patribus suis et sepultus est in Samaria regnavitque Ahab filius eius pro eo
1KGS|16|29|Ahab vero filius Amri regnavit super Israhel anno tricesimo octavo Asa regis Iuda et regnavit Ahab filius Amri super Israhel in Samaria viginti et duobus annis
1KGS|16|30|et fecit Ahab filius Amri malum in conspectu Domini super omnes qui fuerunt ante eum
1KGS|16|31|nec suffecit ei ut ambularet in peccatis Hieroboam filii Nabath insuper duxit uxorem Hiezabel filiam Ethbaal regis Sidoniorum et abiit et servivit Baal et adoravit eum
1KGS|16|32|et posuit aram Baal in templo Baal quod aedificaverat in Samaria
1KGS|16|33|et plantavit lucum et addidit Ahab in opere suo inritans Dominum Deum Israhel super omnes reges Israhel qui fuerant ante eum
1KGS|16|34|in diebus eius aedificavit Ahiel de Bethel Hiericho in Abiram primitivo suo fundavit eam et in Segub novissimo suo posuit portas eius iuxta verbum Domini quod locutus fuerat in manu Iosue filii Nun
1KGS|17|1|et dixit Helias Thesbites de habitatoribus Galaad ad Ahab vivit Dominus Deus Israhel in cuius conspectu sto si erit annis his ros et pluvia nisi iuxta oris mei verba
1KGS|17|2|et factum est verbum Domini ad eum dicens
1KGS|17|3|recede hinc et vade contra orientem et abscondere in torrente Charith qui est contra Iordanem
1KGS|17|4|et ibi de torrente bibes corvisque praecepi ut pascant te ibi
1KGS|17|5|abiit ergo et fecit iuxta verbum Domini cumque abisset sedit in torrente Charith qui est contra Iordanem
1KGS|17|6|corvi quoque deferebant panem et carnes mane similiter panem et carnes vesperi et bibebat de torrente
1KGS|17|7|post dies autem siccatus est torrens non enim pluerat super terram
1KGS|17|8|factus est igitur sermo Domini ad eum dicens
1KGS|17|9|surge et vade in Sareptha Sidoniorum et manebis ibi praecepi enim ibi mulieri viduae ut pascat te
1KGS|17|10|surrexit et abiit Sareptham cumque venisset ad portam civitatis apparuit ei mulier vidua colligens ligna et vocavit eam dixitque da mihi paululum aquae in vase ut bibam
1KGS|17|11|cumque illa pergeret ut adferret clamavit post tergum eius dicens adfer mihi obsecro et buccellam panis in manu tua
1KGS|17|12|quae respondit vivit Dominus Deus tuus quia non habeo panem nisi quantum pugillus capere potest farinae in hydria et paululum olei in lecytho en colligo duo ligna ut ingrediar et faciam illud mihi et filio meo ut comedamus et moriamur
1KGS|17|13|ad quam Helias ait noli timere sed vade et fac sicut dixisti verumtamen mihi primum fac de ipsa farinula subcinericium panem parvulum et adfer ad me tibi autem et filio tuo facies postea
1KGS|17|14|haec autem dicit Dominus Deus Israhel hydria farinae non deficiet nec lecythus olei minuetur usque ad diem in qua daturus est Dominus pluviam super faciem terrae
1KGS|17|15|quae abiit et fecit iuxta verbum Heliae et comedit ipse et illa et domus eius et ex illa die
1KGS|17|16|hydria farinae non defecit et lecythus olei non est inminutus iuxta verbum Domini quod locutus fuerat in manu Heliae
1KGS|17|17|factum est autem post verba haec aegrotavit filius mulieris matris familiae et erat languor fortis nimis ita ut non remaneret in eo halitus
1KGS|17|18|dixit ergo ad Heliam quid mihi et tibi vir Dei ingressus es ad me ut rememorarentur iniquitates meae et interficeres filium meum
1KGS|17|19|et ait ad eam da mihi filium tuum tulitque eum de sinu illius et portavit in cenaculum ubi ipse manebat et posuit super lectulum suum
1KGS|17|20|et clamavit ad Dominum et dixit Domine Deus meus etiamne viduam apud quam ego utcumque sustentor adflixisti ut interficeres filium eius
1KGS|17|21|et expandit se atque mensus est super puerum tribus vicibus clamavitque ad Dominum et ait Domine Deus meus revertatur oro anima pueri huius in viscera eius
1KGS|17|22|exaudivit Dominus vocem Heliae et reversa est anima pueri intra eum et revixit
1KGS|17|23|tulitque Helias puerum et deposuit eum de cenaculo in inferiorem domum et tradidit matri suae et ait illi en vivit filius tuus
1KGS|17|24|dixitque mulier ad Heliam nunc in isto cognovi quoniam vir Dei es tu et verbum Domini in ore tuo verum est
1KGS|18|1|post dies multos verbum Domini factum est ad Heliam in anno tertio dicens vade et ostende te Ahab ut dem pluviam super faciem terrae
1KGS|18|2|ivit ergo Helias ut ostenderet se Ahab erat autem fames vehemens in Samaria
1KGS|18|3|vocavitque Ahab Abdiam dispensatorem domus suae Abdias autem timebat Dominum valde
1KGS|18|4|nam cum interficeret Hiezabel prophetas Domini tulit ille centum prophetas et abscondit eos quinquagenos in speluncis et pavit eos pane et aqua
1KGS|18|5|dixit ergo Ahab ad Abdiam vade in terram ad universos fontes aquarum et in cunctas valles si forte invenire possimus herbam et salvare equos et mulos et non penitus iumenta intereant
1KGS|18|6|diviseruntque sibi regiones ut circuirent eas Ahab ibat per viam unam et Abdias per viam alteram seorsum
1KGS|18|7|cumque esset Abdias in via Helias occurrit ei qui cum cognovisset eum cecidit super faciem suam et ait num tu es domine mi Helias
1KGS|18|8|cui ille respondit ego vade dic domino tuo adest Helias
1KGS|18|9|et ille quid peccavi inquit quoniam trades me servum tuum in manu Ahab ut interficiat me
1KGS|18|10|vivit Dominus Deus tuus non est gens aut regnum quo non miserit dominus meus te requirens et respondentibus cunctis non est hic adiuravit regna singula et gentes eo quod minime repperireris
1KGS|18|11|et nunc dicis mihi vade et dic domino tuo adest Helias
1KGS|18|12|cumque recessero a te spiritus Domini asportabit te in locum quem ego ignoro ingressus nuntiabo Ahab et non inveniet te et interficiet me servus autem tuus timet Dominum ab infantia sua
1KGS|18|13|numquid non indicatum est tibi domino meo quid fecerim cum interficeret Hiezabel prophetas Domini quod absconderim de prophetis Domini centum viros quinquagenos et quinquagenos in speluncis et paverim eos pane et aqua
1KGS|18|14|et nunc tu dicis vade et dic domino tuo adest Helias ut interficiat me
1KGS|18|15|dixit Helias vivit Dominus exercituum ante cuius vultum sto quia hodie apparebo ei
1KGS|18|16|abiit ergo Abdias in occursum Ahab et indicavit ei venitque Ahab in occursum Heliae
1KGS|18|17|et cum vidisset eum ait tune es ille qui conturbas Israhel
1KGS|18|18|et ille ait non turbavi Israhel sed tu et domus patris tui qui dereliquistis mandata Domini et secuti estis Baalim
1KGS|18|19|verumtamen nunc mitte et congrega ad me universum Israhel in monte Carmeli et prophetas Baal quadringentos quinquaginta prophetasque lucorum quadringentos qui comedunt de mensa Hiezabel
1KGS|18|20|misit Ahab ad omnes filios Israhel et congregavit prophetas in monte Carmeli
1KGS|18|21|accedens autem Helias ad omnem populum ait usquequo claudicatis in duas partes si Dominus est Deus sequimini eum si autem Baal sequimini illum et non respondit ei populus verbum
1KGS|18|22|et ait rursum Helias ad populum ego remansi propheta Domini solus prophetae autem Baal quadringenti et quinquaginta viri sunt
1KGS|18|23|dentur nobis duo boves et illi eligant bovem unum et in frusta caedentes ponant super ligna ignem autem non subponant et ego faciam bovem alterum et inponam super ligna ignemque non subponam
1KGS|18|24|invocate nomina deorum vestrorum et ego invocabo nomen Domini et deus qui exaudierit per ignem ipse sit Deus respondens omnis populus ait optima propositio
1KGS|18|25|dixit ergo Helias prophetis Baal eligite vobis bovem unum et facite primi quia vos plures estis et invocate nomina deorum vestrorum ignemque non subponatis
1KGS|18|26|qui cum tulissent bovem quem dederat eis fecerunt et invocabant nomen Baal de mane usque ad meridiem dicentes Baal exaudi nos et non erat vox nec qui responderet transiliebantque altare quod fecerant
1KGS|18|27|cumque esset iam meridies inludebat eis Helias dicens clamate voce maiore deus enim est et forsitan loquitur aut in diversorio est aut in itinere aut certe dormit ut excitetur
1KGS|18|28|clamabant ergo voce magna et incidebant se iuxta ritum suum cultris et lanceolis donec perfunderentur sanguine
1KGS|18|29|postquam autem transiit meridies et illis prophetantibus venerat tempus quo sacrificium offerri solet nec audiebatur vox neque aliquis respondebat nec adtendebat orantes
1KGS|18|30|dixit Helias omni populo venite ad me et accedente ad se populo curavit altare Domini quod destructum fuerat
1KGS|18|31|et tulit duodecim lapides iuxta numerum tribuum filiorum Iacob ad quem factus est sermo Domini dicens Israhel erit nomen tuum
1KGS|18|32|et aedificavit lapidibus altare in nomine Domini fecitque aquaeductum quasi per duas aratiunculas in circuitu altaris
1KGS|18|33|et conposuit ligna divisitque per membra bovem et posuit super ligna
1KGS|18|34|et ait implete quattuor hydrias aqua et fundite super holocaustum et super ligna rursumque dixit etiam secundo hoc facite qui cum fecissent et secundo ait etiam tertio id ipsum facite feceruntque et tertio
1KGS|18|35|et currebant aquae circa altare et fossa aquaeductus repleta est
1KGS|18|36|cumque iam tempus esset ut offerretur holocaustum accedens Helias propheta ait Domine Deus Abraham Isaac et Israhel hodie ostende quia tu es Deus Israhel et ego servus tuus et iuxta praeceptum tuum feci omnia verba haec
1KGS|18|37|exaudi me Domine exaudi me ut discat populus iste quia tu es Dominus Deus et tu convertisti cor eorum iterum
1KGS|18|38|cecidit autem ignis Domini et voravit holocaustum et ligna et lapides pulverem quoque et aquam quae erat in aquaeductu lambens
1KGS|18|39|quod cum vidisset omnis populus cecidit in faciem suam et ait Dominus ipse est Deus Dominus ipse est Deus
1KGS|18|40|dixitque Helias ad eos adprehendite prophetas Baal et ne unus quidem fugiat ex eis quos cum conprehendissent duxit eos Helias ad torrentem Cison et interfecit eos ibi
1KGS|18|41|et ait Helias ad Ahab ascende comede et bibe quia sonus multae pluviae est
1KGS|18|42|ascendit Ahab ut comederet et biberet Helias autem ascendit in vertice Carmeli et pronus in terram posuit faciem inter genua sua
1KGS|18|43|et dixit ad puerum suum ascende et prospice contra mare qui cum ascendisset et contemplatus esset ait non est quicquam et rursum ait illi revertere septem vicibus
1KGS|18|44|in septima autem vice ecce nubicula parva quasi vestigium hominis ascendebat de mari qui ait ascende et dic Ahab iunge et descende ne occupet te pluvia
1KGS|18|45|cumque se verterent huc atque illuc ecce caeli contenebrati sunt et nubes et ventus et facta est pluvia grandis ascendens itaque Ahab abiit in Hiezrahel
1KGS|18|46|et manus Domini facta est super Heliam accinctisque lumbis currebat ante Ahab donec veniret in Hiezrahel
1KGS|19|1|nuntiavit autem Ahab Hiezabel omnia quae fecerat Helias et quomodo occidisset universos prophetas gladio
1KGS|19|2|misitque Hiezabel nuntium ad Heliam dicens haec mihi faciant dii et haec addant nisi hac hora cras posuero animam tuam sicut animam unius ex illis
1KGS|19|3|timuit ergo Helias et surgens abiit quocumque eum ferebat voluntas venitque in Bersabee Iuda et dimisit ibi puerum suum
1KGS|19|4|et perrexit in desertum via unius diei cumque venisset et sederet subter unam iuniperum petivit animae suae ut moreretur et ait sufficit mihi Domine tolle animam meam neque enim melior sum quam patres mei
1KGS|19|5|proiecitque se et obdormivit in umbra iuniperi et ecce angelus tetigit eum et dixit illi surge comede
1KGS|19|6|respexit et ecce ad caput suum subcinericius panis et vas aquae comedit ergo et bibit et rursum obdormivit
1KGS|19|7|reversusque est angelus Domini secundo et tetigit eum dixitque illi surge comede grandis enim tibi restat via
1KGS|19|8|qui cum surrexisset comedit et bibit et ambulavit in fortitudine cibi illius quadraginta diebus et quadraginta noctibus usque ad montem Dei Horeb
1KGS|19|9|cumque venisset illuc mansit in spelunca et ecce sermo Domini ad eum dixitque illi quid hic agis Helia
1KGS|19|10|at ille respondit zelo zelatus sum pro Domino Deo exercituum quia dereliquerunt pactum Domini filii Israhel altaria tua destruxerunt et prophetas tuos occiderunt gladio et derelictus sum ego solus et quaerunt animam meam ut auferant eam
1KGS|19|11|et ait ei egredere et sta in monte coram Domino et ecce Dominus transit et spiritus grandis et fortis subvertens montes et conterens petras ante Dominum non in spiritu Dominus et post spiritum commotio non in commotione Dominus
1KGS|19|12|et post commotionem ignis non in igne Dominus et post ignem sibilus aurae tenuis
1KGS|19|13|quod cum audisset Helias operuit vultum suum pallio et egressus stetit in ostio speluncae et ecce vox ad eum dicens quid agis hic Helia
1KGS|19|14|et ille respondit zelo zelatus sum pro Domino Deo exercituum quia dereliquerunt pactum tuum filii Israhel altaria tua destruxerunt et prophetas tuos occiderunt gladio et derelictus sum ego solus et quaerunt animam meam ut auferant eam
1KGS|19|15|et ait Dominus ad eum vade et revertere in viam tuam per desertum in Damascum cumque perveneris ungues Azahel regem super Syriam
1KGS|19|16|et Hieu filium Namsi ungues regem super Israhel Heliseum autem filium Saphat qui est de Abelmaula ungues prophetam pro te
1KGS|19|17|et erit quicumque fugerit gladium Azahel occidet eum Hieu et qui fugerit gladium Hieu interficiet eum Heliseus
1KGS|19|18|et derelinquam mihi in Israhel septem milia universorum genua quae non sunt incurvata Baal et omne os quod non adoravit eum osculans manum
1KGS|19|19|profectus ergo inde repperit Heliseum filium Saphat arantem duodecim iugis boum et ipse in duodecim arantibus unus erat cumque venisset Helias ad eum misit pallium suum super illum
1KGS|19|20|qui statim relictis bubus cucurrit post Heliam et ait osculer oro te patrem meum et matrem meam et sic sequar te dixitque ei vade et revertere quod enim meum erat feci tibi
1KGS|19|21|reversus autem ab eo tulit par boum et mactavit illud et in aratro boum coxit carnes et dedit populo et comederunt consurgensque abiit et secutus est Heliam et ministrabat ei
1KGS|20|1|porro Benadad rex Syriae congregavit omnem exercitum suum et triginta et duos reges secum et equos et currus et ascendens pugnabat contra Samariam et obsidebat eam
1KGS|20|2|mittensque nuntios ad Ahab regem Israhel in civitatem
1KGS|20|3|ait haec dicit Benadad argentum tuum et aurum tuum meum est et uxores tuae et filii tui optimi mei sunt
1KGS|20|4|responditque rex Israhel iuxta verbum tuum domine mi rex tuus sum ego et omnia mea
1KGS|20|5|revertentesque nuntii dixerunt haec dicit Benadad qui misit nos ad te argentum tuum et aurum tuum et uxores tuas et filios tuos dabis mihi
1KGS|20|6|cras igitur hac eadem hora mittam servos meos ad te et scrutabuntur domum tuam et domum servorum tuorum et omne quod eis placuerit ponent in manibus suis et auferent
1KGS|20|7|vocavit autem rex Israhel omnes seniores terrae et ait animadvertite et videte quoniam insidietur nobis misit enim ad me pro uxoribus meis et filiis et pro argento et auro et non abnui
1KGS|20|8|dixeruntque omnes maiores natu et universus populus ad eum non audias neque adquiescas illi
1KGS|20|9|respondit itaque nuntiis Benadad dicite domino meo regi omnia propter quae misisti ad me servum tuum initio faciam hanc autem rem facere non possum
1KGS|20|10|reversique nuntii rettulerunt ei qui remisit et ait haec faciant mihi dii et haec addant si suffecerit pulvis Samariae pugillis omnis populi qui sequitur me
1KGS|20|11|et respondens rex Israhel ait dicite ei ne glorietur accinctus aeque ut discinctus
1KGS|20|12|factum est autem cum audisset verbum istud bibebat ipse et reges in umbraculis et ait servis suis circumdate civitatem et circumdederunt eam
1KGS|20|13|et ecce propheta unus accedens ad Ahab regem Israhel ait haec dicit Dominus certe vidisti omnem multitudinem hanc nimiam ecce ego tradam eam in manu tua hodie ut scias quia ego sum Dominus
1KGS|20|14|et ait Ahab per quem dixitque ei haec dicit Dominus per pedisequos principum provinciarum et ait quis incipiet proeliari et ille dixit tu
1KGS|20|15|recensuit ergo pueros principum provinciarum et repperit numerum ducentorum triginta duum et post eos recensuit populum omnes filios Israhel septem milia
1KGS|20|16|et egressi sunt meridie Benadad autem bibebat temulentus in umbraculo suo et reges triginta duo cum eo qui ad auxilium eius venerant
1KGS|20|17|egressi sunt autem pueri principum provinciarum in prima fronte misit itaque Benadad qui nuntiaverunt ei dicentes viri egressi sunt de Samaria
1KGS|20|18|at ille sive ait pro pace veniunt adprehendite eos vivos sive ut proelientur vivos eos capite
1KGS|20|19|egressi sunt ergo pueri principum provinciarum ac reliquus exercitus sequebatur
1KGS|20|20|et percussit unusquisque virum qui contra se venerat fugeruntque Syri et persecutus est eos Israhel fugit quoque Benadad rex Syriae in equo cum equitibus
1KGS|20|21|necnon et egressus rex Israhel percussit equos et currus et percussit Syriam plaga magna
1KGS|20|22|accedens autem propheta ad regem Israhel dixit ei vade et confortare et scito et vide quid facias sequenti enim anno rex Syriae ascendet contra te
1KGS|20|23|servi vero regis Syriae dixerunt ei dii montium sunt dii eorum ideo superaverunt nos sed melius est ut pugnemus contra eos in campestribus et obtinebimus eos
1KGS|20|24|tu ergo verbum hoc fac amove reges singulos ab exercitu suo et pone principes pro eis
1KGS|20|25|et instaura numerum militum qui ceciderunt de tuis et equos secundum equos pristinos et currus secundum currus quos ante habuisti et pugnabimus contra eos in campestribus et videbis quod obtinebimus eos credidit consilio eorum et fecit ita
1KGS|20|26|igitur postquam annus transierat recensuit Benadad Syros et ascendit in Afec ut pugnaret contra Israhel
1KGS|20|27|porro filii Israhel recensiti sunt et acceptis cibariis profecti ex adverso castraque metati contra eos quasi duo parvi greges caprarum Syri autem repleverunt terram
1KGS|20|28|et accedens unus vir Dei dixit ad regem Israhel haec dicit Dominus quia dixerunt Syri deus montium est Dominus et non est deus vallium dabo omnem multitudinem grandem hanc in manu tua et scietis quia ego Dominus
1KGS|20|29|dirigebant septem diebus ex adverso hii atque illi acies septima autem die commissum est bellum percusseruntque filii Israhel de Syris centum milia peditum in die una
1KGS|20|30|fugerunt autem qui remanserant in Afec in civitatem et cecidit murus super viginti septem milia hominum qui remanserant porro Benadad fugiens ingressus est civitatem in cubiculum quod erat intra cubiculum
1KGS|20|31|dixeruntque ei servi sui ecce audivimus quod reges domus Israhel clementes sint ponamus itaque saccos in lumbis nostris et funiculos in capitibus nostris et egrediamur ad regem Israhel forsitan salvabit animas nostras
1KGS|20|32|accinxerunt saccis lumbos suos et posuerunt funes in capitibus veneruntque ad regem Israhel et dixerunt servus tuus Benadad dicit vivat oro te anima mea et ille ait si adhuc vivit frater meus est
1KGS|20|33|quod acceperunt viri pro omine et festinantes rapuerunt verbum ex ore eius atque dixerunt frater tuus Benadad et dixit eis ite et adducite eum egressus est ergo ad eum Benadad et levavit eum in currum suum
1KGS|20|34|qui dixit ei civitates quas tulit pater meus a patre tuo reddam et plateas fac tibi in Damasco sicut fecit pater meus in Samaria et ego foederatus recedam a te pepigit ergo foedus et dimisit eum
1KGS|20|35|tunc vir quidam de filiis prophetarum dixit ad socium suum in sermone Domini percute me at ille noluit percutere
1KGS|20|36|cui ait quia noluisti audire vocem Domini ecce recedes a me et percutiet te leo cumque paululum recessisset ab eo invenit eum leo atque percussit
1KGS|20|37|sed et alterum conveniens virum dixit ad eum percute me qui percussit eum et vulneravit
1KGS|20|38|abiit ergo propheta et occurrit regi in via et mutavit aspersione pulveris os et oculos suos
1KGS|20|39|cumque rex transiret clamavit ad regem et ait servus tuus egressus est ad proeliandum comminus cumque fugisset vir unus adduxit eum quidam ad me et ait custodi virum istum qui si lapsus fuerit erit anima tua pro anima eius aut talentum argenti adpendes
1KGS|20|40|dum autem ego turbatus huc illucque me verterem subito non conparuit et ait rex Israhel ad eum hoc est iudicium tuum quod ipse decrevisti
1KGS|20|41|at ille statim abstersit pulverem de facie sua et cognovit eum rex Israhel quod esset de prophetis
1KGS|20|42|qui ait ad eum haec dicit Dominus quia dimisisti virum dignum morte de manu tua erit anima tua pro anima eius et populus tuus pro populo eius
1KGS|20|43|reversus est igitur rex Israhel in domum suam audire contemnens et furibundus venit Samariam
1KGS|21|1|post verba autem haec vinea erat Naboth Hiezrahelitae qui erat in Hiezrahel iuxta palatium Ahab regis Samariae
1KGS|21|2|locutus est ergo Ahab ad Naboth dicens da mihi vineam tuam ut faciam mihi hortum holerum quia vicina est et prope domum meam daboque tibi pro ea vineam meliorem aut si tibi commodius putas argenti pretium quanto digna est
1KGS|21|3|cui respondit Naboth propitius mihi sit Dominus ne dem hereditatem patrum meorum tibi
1KGS|21|4|venit ergo Ahab in domum suam indignans et frendens super verbo quod locutus fuerat ad eum Naboth Hiezrahelites dicens non do tibi hereditatem patrum meorum et proiciens se in lectulum suum avertit faciem ad parietem et non comedit panem
1KGS|21|5|ingressa est autem ad eum Hiezabel uxor sua dixitque ei quid est hoc unde anima tua contristata est et quare non comedis panem
1KGS|21|6|qui respondit ei locutus sum Naboth Hiezrahelitae et dixi ei da mihi vineam tuam accepta pecunia aut si tibi placet dabo tibi vineam pro ea et ille ait non do tibi vineam meam
1KGS|21|7|dixit ergo ad eum Hiezabel uxor eius grandis auctoritatis es et bene regis regnum Israhel surge et comede panem et aequo esto animo ego dabo tibi vineam Naboth Hiezrahelitae
1KGS|21|8|scripsit itaque litteras ex nomine Ahab et signavit eas anulo eius et misit ad maiores natu et ad optimates qui erant in civitate eius et habitabant cum Naboth
1KGS|21|9|litterarum autem erat ista sententia praedicate ieiunium et sedere facite Naboth inter primos populi
1KGS|21|10|et submittite duos viros filios Belial contra eum et falsum testimonium dicant benedixit Deum et regem et educite eum et lapidate sicque moriatur
1KGS|21|11|fecerunt ergo cives eius maiores natu et optimates qui habitabant cum eo in urbe sicut praeceperat eis Hiezabel et sicut scriptum erat in litteris quas miserat ad eos
1KGS|21|12|praedicaverunt ieiunium et sedere fecerunt Naboth inter primos populi
1KGS|21|13|et adductis duobus viris filiis diaboli fecerunt eos sedere contra eum at illi scilicet ut viri diabolici dixerunt contra eum testimonium coram multitudine benedixit Naboth Deo et regi quam ob rem eduxerunt eum extra civitatem et lapidibus interfecerunt
1KGS|21|14|miseruntque ad Hiezabel dicentes lapidatus est Naboth et mortuus est
1KGS|21|15|factum est autem cum audisset Hiezabel lapidatum Naboth et mortuum locuta est ad Ahab surge posside vineam Naboth Hiezrahelitae qui noluit tibi adquiescere et dare eam accepta pecunia non enim vivit Naboth sed mortuus est
1KGS|21|16|quod cum audisset Ahab mortuum videlicet Naboth surrexit et descendebat in vineam Naboth Hiezrahelitae ut possideret eam
1KGS|21|17|factus est igitur sermo Domini ad Heliam Thesbiten dicens
1KGS|21|18|surge et descende in occursum Ahab regis Israhel qui est in Samaria ecce ad vineam Naboth descendit ut possideat eam
1KGS|21|19|et loqueris ad eum dicens haec dicit Dominus occidisti insuper et possedisti et post haec addes haec dicit Dominus in loco hoc in quo linxerunt canes sanguinem Naboth lambent tuum quoque sanguinem
1KGS|21|20|et ait Ahab ad Heliam num invenisti me inimice mee qui dixit inveni eo quod venundatus sis ut faceres malum in conspectu Domini
1KGS|21|21|ecce ego inducam super te malum et demetam posteriora tua et interficiam de Ahab mingentem ad parietem et clausum et ultimum in Israhel
1KGS|21|22|et dabo domum tuam sicut domum Hieroboam filii Nabath et sicut domum Baasa filii Ahia quia egisti ut me ad iracundiam provocares et peccare fecisti Israhel
1KGS|21|23|sed et de Hiezabel locutus est Dominus dicens canes comedent Hiezabel in agro Hiezrahel
1KGS|21|24|si mortuus fuerit Ahab in civitate comedent eum canes si autem mortuus fuerit in agro comedent eum volucres caeli
1KGS|21|25|igitur non fuit alter talis ut Ahab qui venundatus est ut faceret malum in conspectu Domini concitavit enim eum Hiezabel uxor sua
1KGS|21|26|et abominabilis effectus est in tantum ut sequeretur idola quae fecerant Amorrei quos consumpsit Dominus a facie filiorum Israhel
1KGS|21|27|itaque cum audisset Ahab sermones istos scidit vestem suam et operuit cilicio carnem suam ieiunavitque et dormivit in sacco et ambulabat dimisso capite
1KGS|21|28|factus est autem sermo Domini ad Heliam Thesbiten dicens
1KGS|21|29|nonne vidisti humiliatum Ahab coram me quia igitur humiliatus est mei causa non inducam malum in diebus eius sed in diebus filii sui inferam malum domui eius
1KGS|22|1|transierunt igitur tres anni absque bello inter Syriam et Israhel
1KGS|22|2|in anno autem tertio descendit Iosaphat rex Iuda ad regem Israhel
1KGS|22|3|dixitque rex Israhel ad servos suos ignoratis quod nostra sit Ramoth Galaad et neglegimus tollere eam de manu regis Syriae
1KGS|22|4|et ait ad Iosaphat veniesne mecum ad proeliandum in Ramoth Galaad
1KGS|22|5|dixitque Iosaphat ad regem Israhel sicut ego sum ita et tu populus meus et populus tuus unum sunt et equites mei et equites tui dixitque Iosaphat ad regem Israhel quaere oro te hodie sermonem Domini
1KGS|22|6|congregavit ergo rex Israhel prophetas quadringentos circiter viros et ait ad eos ire debeo in Ramoth Galaad ad bellandum an quiescere qui responderunt ascende et dabit Dominus in manu regis
1KGS|22|7|dixit autem Iosaphat non est hic propheta Domini quispiam ut interrogemus per eum
1KGS|22|8|et ait rex Israhel ad Iosaphat remansit vir unus per quem possimus interrogare Dominum sed ego odi eum quia non prophetat mihi bonum sed malum Micheas filius Hiemla cui Iosaphat ait ne loquaris ita rex
1KGS|22|9|vocavit ergo rex Israhel eunuchum quendam et dixit ei festina adducere Micheam filium Hiemla
1KGS|22|10|rex autem Israhel et Iosaphat rex Iuda sedebat unusquisque in solio suo vestiti cultu regio in area iuxta ostium portae Samariae et universi prophetae prophetabant in conspectu eorum
1KGS|22|11|fecit quoque sibi Sedecias filius Chanaan cornua ferrea et ait haec dicit Dominus his ventilabis Syriam donec deleas eam
1KGS|22|12|omnesque prophetae similiter prophetabant dicentes ascende in Ramoth Galaad et vade prospere et tradet Dominus in manu regis
1KGS|22|13|nuntius vero qui ierat ut vocaret Micheam locutus est ad eum dicens ecce sermones prophetarum ore uno bona regi praedicant sit ergo et sermo tuus similis eorum et loquere bona
1KGS|22|14|cui Micheas ait vivit Dominus quia quodcumque dixerit mihi Dominus hoc loquar
1KGS|22|15|venit itaque ad regem et ait illi rex Michea ire debemus in Ramoth Galaad ad proeliandum an cessare cui ille respondit ascende et vade prospere et tradet Dominus in manu regis
1KGS|22|16|dixit autem rex ad eum iterum atque iterum adiuro te ut non loquaris mihi nisi quod verum est in nomine Domini
1KGS|22|17|et ille ait vidi cunctum Israhel dispersum in montibus quasi oves non habentes pastorem et ait Dominus non habent dominum isti revertatur unusquisque in domum suam in pace
1KGS|22|18|dixit ergo rex Israhel ad Iosaphat numquid non dixi tibi quia non prophetat mihi bonum sed semper malum
1KGS|22|19|ille vero addens ait propterea audi sermonem Domini vidi Dominum sedentem super solium suum et omnem exercitum caeli adsistentem ei a dextris et a sinistris
1KGS|22|20|et ait Dominus quis decipiet Ahab regem Israhel ut ascendat et cadat in Ramoth Galaad et dixit unus verba huiuscemodi et alius aliter
1KGS|22|21|egressus est autem spiritus et stetit coram Domino et ait ego decipiam illum cui locutus est Dominus in quo
1KGS|22|22|et ille ait egrediar et ero spiritus mendax in ore omnium prophetarum eius et dixit Dominus decipies et praevalebis egredere et fac ita
1KGS|22|23|nunc igitur ecce dedit Dominus spiritum mendacii in ore omnium prophetarum tuorum qui hic sunt et Dominus locutus est contra te malum
1KGS|22|24|accessit autem Sedecias filius Chanaan et percussit Micheam in maxillam et dixit mene ergo dimisit spiritus Domini et locutus est tibi
1KGS|22|25|et ait Micheas visurus es in die illa quando ingredieris cubiculum intra cubiculum ut abscondaris
1KGS|22|26|et ait rex Israhel tollite Micheam et maneat apud Amon principem civitatis et apud Ioas filium Ammelech
1KGS|22|27|et dicite eis haec dicit rex mittite virum istum in carcerem et sustentate eum pane tribulationis et aqua angustiae donec revertar in pace
1KGS|22|28|dixitque Micheas si reversus fueris in pace non est locutus Dominus in me et ait audite populi omnes
1KGS|22|29|ascendit itaque rex Israhel et Iosaphat rex Iuda in Ramoth Galaad
1KGS|22|30|dixitque rex Israhel ad Iosaphat sume arma et ingredere proelium et induere vestibus tuis porro rex Israhel mutavit habitum et ingressus est bellum
1KGS|22|31|rex autem Syriae praeceperat principibus curruum triginta duobus dicens non pugnabitis contra minorem et maiorem quempiam nisi contra regem Israhel solum
1KGS|22|32|cum ergo vidissent principes curruum Iosaphat suspicati sunt quod ipse esset rex Israhel et impetu facto pugnabant contra eum et exclamavit Iosaphat
1KGS|22|33|intellexeruntque principes curruum quod non esset rex Israhel et cessaverunt ab eo
1KGS|22|34|unus autem quidam tetendit arcum in incertum sagittam dirigens et casu percussit regem Israhel inter pulmonem et stomachum at ille dixit aurigae suo verte manum tuam et eice me de exercitu quia graviter vulneratus sum
1KGS|22|35|commissum est ergo proelium in die illa et rex Israhel stabat in curru suo contra Syros et mortuus est vesperi fluebat autem sanguis plagae in sinum currus
1KGS|22|36|et praeco personuit in universo exercitu antequam sol occumberet dicens unusquisque revertatur in civitatem et in terram suam
1KGS|22|37|mortuus est autem rex et perlatus est Samariam sepelieruntque regem in Samaria
1KGS|22|38|et laverunt currum in piscina Samariae et linxerunt canes sanguinem eius et habenas laverunt iuxta verbum Domini quod locutus fuerat
1KGS|22|39|reliqua vero sermonum Ahab et universa quae fecit et domus eburneae quam aedificavit cunctarumque urbium quas extruxit nonne scripta sunt haec in libro verborum dierum regum Israhel
1KGS|22|40|dormivit ergo Ahab cum patribus suis et regnavit Ohozias filius eius pro eo
1KGS|22|41|Iosaphat filius Asa regnare coeperat super Iudam anno quarto Ahab regis Israhel
1KGS|22|42|triginta quinque annorum erat cum regnare coepisset et viginti et quinque annos regnavit in Hierusalem nomen matris eius Azuba filia Salai
1KGS|22|43|et ambulavit in omni via Asa patris sui et non declinavit ex ea fecitque quod rectum est in conspectu Domini
1KGS|22|44|verumtamen excelsa non abstulit adhuc enim populus sacrificabat et adolebat incensum in excelsis
1KGS|22|45|pacemque habuit Iosaphat cum rege Israhel
1KGS|22|46|reliqua autem verborum Iosaphat et opera eius quae gessit et proelia nonne haec scripta sunt in libro verborum dierum regum Iuda
1KGS|22|47|sed et reliquias effeminatorum qui remanserant in diebus Asa patris eius abstulit de terra
1KGS|22|48|nec erat tunc rex constitutus in Edom
1KGS|22|49|rex vero Iosaphat fecerat classes in mari quae navigarent in Ophir propter aurum et ire non potuerunt quia confractae sunt in Asiongaber
1KGS|22|50|tunc ait Ohozias filius Ahab ad Iosaphat vadant servi mei cum servis tuis in navibus et noluit Iosaphat
1KGS|22|51|dormivitque cum patribus suis et sepultus est cum eis in civitate David patris sui regnavitque Ioram filius eius pro eo
1KGS|22|52|Ohozias autem filius Ahab regnare coeperat super Israhel in Samaria anno septimodecimo Iosaphat regis Iuda regnavitque super Israhel duobus annis
1KGS|22|53|et fecit malum in conspectu Domini et ambulavit in via patris sui et matris suae et in via Hieroboam filii Nabath qui peccare fecit Israhel
1KGS|22|54|servivit quoque Baal et adoravit eum et inritavit Dominum Deum Israhel iuxta omnia quae fecerat pater eius
2KGS|1|1|praevaricatus est autem Moab in Israhel postquam mortuus est Ahab
2KGS|1|2|ceciditque Ohozias per cancellos cenaculi sui quod habebat in Samaria et aegrotavit misitque nuntios dicens ad eos ite consulite Beelzebub deum Accaron utrum vivere queam de infirmitate mea hac
2KGS|1|3|angelus autem Domini locutus est ad Heliam Thesbiten surge ascende in occursum nuntiorum regis Samariae et dices ad eos numquid non est Deus in Israhel ut eatis ad consulendum Beelzebub deum Accaron
2KGS|1|4|quam ob rem haec dicit Dominus de lectulo super quem ascendisti non descendes sed morte morieris et abiit Helias
2KGS|1|5|reversique sunt nuntii ad Ohoziam qui dixit eis quare reversi estis
2KGS|1|6|at illi responderunt ei vir occurrit nobis et dixit ad nos ite revertimini ad regem qui misit vos et dicetis ei haec dicit Dominus numquid quia non erat Deus in Israhel mittis ut consulatur Beelzebub deus Accaron idcirco de lectulo super quem ascendisti non descendes sed morte morieris
2KGS|1|7|qui dixit eis cuius figurae et habitu est vir qui occurrit vobis et locutus est verba haec
2KGS|1|8|at illi dixerunt vir pilosus et zona pellicia accinctis renibus qui ait Helias Thesbites est
2KGS|1|9|misitque ad eum quinquagenarium principem et quinquaginta qui erant sub eo qui ascendit ad eum sedentique in vertice montis ait homo Dei rex praecepit ut descendas
2KGS|1|10|respondensque Helias dixit quinquagenario si homo Dei sum descendat ignis e caelo et devoret te et quinquaginta tuos descendit itaque ignis e caelo et devoravit eum et quinquaginta qui erant cum eo
2KGS|1|11|rursum misit ad eum principem quinquagenarium alterum et quinquaginta cum eo qui locutus est illi homo Dei haec dicit rex festina descende
2KGS|1|12|respondens Helias ait si homo Dei ego sum descendat ignis e caelo et devoret te et quinquaginta tuos descendit ergo ignis Dei e caelo et devoravit illum et quinquaginta eius
2KGS|1|13|iterum misit principem quinquagenarium tertium et quinquaginta qui erant cum eo qui cum venisset curvavit genua contra Heliam et precatus est eum et ait homo Dei noli despicere animam meam et animam servorum tuorum qui mecum sunt
2KGS|1|14|ecce descendit ignis de caelo et devoravit duos principes quinquagenarios primos et quinquagenos qui cum eis erant sed nunc obsecro ut miserearis animae meae
2KGS|1|15|locutus est autem angelus Domini ad Heliam dicens descende cum eo ne timeas surrexit igitur et descendit cum eo ad regem
2KGS|1|16|et locutus est ei haec dicit Dominus quia misisti nuntios ad consulendum Beelzebub deum Accaron quasi non esset Deus in Israhel a quo possis interrogare sermonem ideo de lectulo super quem ascendisti non descendes sed morte morieris
2KGS|1|17|mortuus est ergo iuxta sermonem Domini quem locutus est Helias et regnavit Ioram frater eius pro eo anno secundo Ioram filii Iosaphat regis Iudae non enim habebat filium
2KGS|1|18|reliqua autem verborum Ohoziae quae operatus est nonne haec scripta sunt in libro sermonum dierum regum Israhel
2KGS|2|1|factum est autem cum levare vellet Dominus Heliam per turbinem in caelum ibant Helias et Heliseus de Galgalis
2KGS|2|2|dixitque Helias ad Heliseum sede hic quia Dominus misit me usque Bethel cui ait Heliseus vivit Dominus et vivit anima tua quia non derelinquam te cumque descendissent Bethel
2KGS|2|3|egressi sunt filii prophetarum qui erant Bethel ad Heliseum et dixerunt ei numquid nosti quia hodie Dominus tollat dominum tuum a te qui respondit et ego novi silete
2KGS|2|4|dixit autem Helias ad Heliseum sede hic quia Dominus misit me in Hiericho et ille ait vivit Dominus et vivit anima tua quia non derelinquam te cumque venissent Hierichum
2KGS|2|5|accesserunt filii prophetarum qui erant in Hiericho ad Heliseum et dixerunt ei numquid nosti quia hodie Dominus tollet dominum tuum a te et ait et ego novi silete
2KGS|2|6|dixit autem ei Helias sede hic quia Dominus misit me ad Iordanem qui ait vivit Dominus et vivit anima tua quia non derelinquam te ierunt igitur ambo pariter
2KGS|2|7|et quinquaginta viri de filiis prophetarum secuti sunt qui et steterunt e contra longe illi autem ambo stabant super Iordanem
2KGS|2|8|tulitque Helias pallium suum et involvit illud et percussit aquas quae divisae sunt in utramque partem et transierunt ambo per siccum
2KGS|2|9|cumque transissent Helias dixit ad Heliseum postula quod vis ut faciam tibi antequam tollar a te dixitque Heliseus obsecro ut fiat duplex spiritus tuus in me
2KGS|2|10|qui respondit rem difficilem postulasti attamen si videris me quando tollor a te erit quod petisti si autem non videris non erit
2KGS|2|11|cumque pergerent et incedentes sermocinarentur ecce currus igneus et equi ignei diviserunt utrumque et ascendit Helias per turbinem in caelum
2KGS|2|12|Heliseus autem videbat et clamabat pater mi pater mi currus Israhel et auriga eius et non vidit eum amplius adprehenditque vestimenta sua et scidit illa in duas partes
2KGS|2|13|et levavit pallium Heliae quod ceciderat ei reversusque stetit super ripam Iordanis
2KGS|2|14|et pallio Heliae quod ceciderat ei percussit aquas et dixit ubi est Deus Heliae etiam nunc percussitque aquas et divisae sunt huc atque illuc et transiit Heliseus
2KGS|2|15|videntes autem filii prophetarum qui erant in Hiericho de contra dixerunt requievit spiritus Heliae super Heliseum et venientes in occursum eius adoraverunt eum proni in terram
2KGS|2|16|dixeruntque illi ecce cum servis tuis sunt quinquaginta viri fortes qui possint ire et quaerere dominum tuum ne forte tulerit eum spiritus Domini et proiecerit in uno montium aut in una vallium qui ait nolite mittere
2KGS|2|17|coegeruntque eum donec adquiesceret et diceret mittite et miserunt quinquaginta viros qui cum quaesissent tribus diebus non invenerunt
2KGS|2|18|et reversi sunt ad eum at ille habitabat in Hiericho dixitque eis numquid non dixi vobis nolite ire
2KGS|2|19|dixerunt quoque viri civitatis ad Heliseum ecce habitatio civitatis huius optima est sicut tu ipse domine perspicis sed aquae pessimae sunt et terra sterilis
2KGS|2|20|at ille ait adferte mihi vas novum et mittite in illud sal qui cum adtulissent
2KGS|2|21|egressus ad fontem aquarum misit in eum sal et ait haec dicit Dominus sanavi aquas has et non erit ultra in eis mors neque sterilitas
2KGS|2|22|sanatae sunt ergo aquae usque ad diem hanc iuxta verbum Helisei quod locutus est
2KGS|2|23|ascendit autem inde Bethel cumque ascenderet per viam pueri parvi egressi sunt de civitate et inludebant ei dicentes ascende calve ascende calve
2KGS|2|24|qui cum se respexisset vidit eos et maledixit eis in nomine Domini egressique sunt duo ursi de saltu et laceraverunt ex eis quadraginta duos pueros
2KGS|2|25|abiit autem inde in montem Carmeli et inde reversus est Samariam
2KGS|3|1|Ioram vero filius Ahab regnavit super Israhel in Samaria anno octavodecimo Iosaphat regis Iudae regnavitque duodecim annis
2KGS|3|2|et fecit malum coram Domino sed non sicut pater suus et mater tulit enim statuas Baal quas fecerat pater eius
2KGS|3|3|verumtamen in peccatis Hieroboam filii Nabath qui peccare fecit Israhel adhesit nec recessit ab eis
2KGS|3|4|porro Mesa rex Moab nutriebat pecora multa et solvebat regi Israhel centum milia agnorum et centum milia arietum cum velleribus suis
2KGS|3|5|cumque mortuus fuisset Ahab praevaricatus est foedus quod habebat cum rege Israhel
2KGS|3|6|egressus est igitur rex Ioram in die illa de Samaria et recensuit universum Israhel
2KGS|3|7|misitque ad Iosaphat regem Iuda dicens rex Moab recessit a me veni mecum contra Moab ad proelium qui respondit ascendam qui meus est tuus est populus meus populus tuus equi mei equi tui
2KGS|3|8|dixitque per quam viam ascendemus at ille respondit per desertum Idumeae
2KGS|3|9|perrexerunt igitur rex Israhel et rex Iuda et rex Edom et circumierunt per viam septem dierum nec erat aqua exercitui et iumentis quae sequebantur eos
2KGS|3|10|dixitque rex Israhel eheu eheu eheu congregavit nos Dominus tres reges ut traderet in manu Moab
2KGS|3|11|et ait Iosaphat estne hic propheta Domini ut deprecemur Dominum per eum et respondit unus de servis regis Israhel est hic Heliseus filius Saphat qui fundebat aquam super manus Heliae
2KGS|3|12|et ait Iosaphat est apud eum sermo Domini descenditque ad eum rex Israhel et Iosaphat et rex Edom
2KGS|3|13|dixit autem Heliseus ad regem Israhel quid mihi et tibi est vade ad prophetas patris tui et matris tuae et ait illi rex Israhel quare congregavit Dominus tres reges hos ut traderet eos in manu Moab
2KGS|3|14|dixit autem Heliseus vivit Dominus exercituum in cuius conspectu sto quod si non vultum Iosaphat regis Iudae erubescerem ne adtendissem quidem te nec respexissem
2KGS|3|15|nunc autem adducite mihi psalten cumque caneret psaltes facta est super eum manus Domini et ait
2KGS|3|16|haec dicit Dominus facite alveum torrentis huius fossas et fossas
2KGS|3|17|haec enim dicit Dominus non videbitis ventum neque pluviam et alveus iste replebitur aquis et bibetis vos et familiae vestrae et iumenta vestra
2KGS|3|18|parumque hoc est in conspectu Domini insuper tradet etiam Moab in manu vestra
2KGS|3|19|et percutietis omnem civitatem munitam et omnem urbem electam et universum lignum fructiferum succidetis cunctosque fontes aquarum obturabitis et omnem agrum egregium operietis lapidibus
2KGS|3|20|factum est igitur mane quando sacrificium offerri solet et ecce aquae veniebant per viam Edom et repleta est terra aquis
2KGS|3|21|universi autem Moabitae audientes quod ascendissent reges ut pugnarent adversum eos convocaverunt omnes qui accincti erant balteo desuper et steterunt in terminis
2KGS|3|22|primoque mane surgentes et orto iam sole ex adverso aquarum viderunt Moabitae contra aquas rubras quasi sanguinem
2KGS|3|23|dixeruntque sanguis est gladii pugnaverunt reges contra se et caesi sunt mutuo nunc perge ad praedam Moab
2KGS|3|24|perrexeruntque in castra Israhel porro consurgens Israhel percussit Moab at illi fugerunt coram eis venerunt igitur qui vicerant et percusserunt Moab
2KGS|3|25|et civitates destruxerunt et omnem agrum optimum mittentes singuli lapides repleverunt et universos fontes aquarum obturaverunt et omnia ligna fructifera succiderunt ita ut muri tantum fictiles remanerent et circumdata est civitas a fundibalariis et magna ex parte percussa
2KGS|3|26|quod cum vidisset rex Moab praevaluisse scilicet hostes tulit secum septingentos viros educentes gladium ut inrumperet ad regem Edom et non potuerunt
2KGS|3|27|arripiensque filium suum primogenitum qui regnaturus erat pro eo obtulit holocaustum super murum et facta est indignatio magna in Israhel statimque recesserunt ab eo et reversi sunt in terram suam
2KGS|4|1|mulier autem quaedam de uxoribus prophetarum clamabat ad Heliseum dicens servus tuus vir meus mortuus est et tu nosti quia servus tuus fuit timens Dominum et ecce creditor venit ut tollat duos filios meos ad serviendum sibi
2KGS|4|2|cui dixit Heliseus quid vis ut faciam tibi dic mihi quid habes in domo tua at illa respondit non habeo ancilla tua quicquam in domo mea nisi parum olei quo unguear
2KGS|4|3|cui ait vade pete mutuo ab omnibus vicinis tuis vasa vacua non pauca
2KGS|4|4|et ingredere et claude ostium cum intrinsecus fueris tu et filii tui et mitte inde in omnia vasa haec et cum plena fuerint tolles
2KGS|4|5|ivit itaque mulier et clusit ostium super se et super filios suos illi offerebant vasa et illa infundebat
2KGS|4|6|cumque plena fuissent vasa dixit ad filium suum adfer mihi adhuc vas et ille respondit non habeo stetitque oleum
2KGS|4|7|venit autem illa et indicavit homini Dei et ille vade inquit vende oleum et redde creditori tuo tu autem et filii tui vivite de reliquo
2KGS|4|8|facta est autem quaedam dies et transiebat Heliseus per Sunam erat autem ibi mulier magna quae tenuit eum ut comederet panem cumque frequenter inde transiret devertebat ad eam ut comederet panem
2KGS|4|9|quae dixit ad virum suum animadverto quod vir Dei sanctus est iste qui transit per nos frequenter
2KGS|4|10|faciamus ergo cenaculum parvum et ponamus ei in eo lectulum et mensam et sellam et candelabrum ut cum venerit ad nos maneat ibi
2KGS|4|11|facta est igitur dies quaedam et veniens devertit in cenaculum et requievit ibi
2KGS|4|12|dixitque ad Giezi puerum suum voca Sunamitin istam qui cum vocasset eam et illa stetisset coram eo
2KGS|4|13|dixit ad puerum loquere ad eam ecce sedule in omnibus ministrasti nobis quid vis ut faciam tibi numquid habes negotium et vis ut loquar regi sive principi militiae quae respondit in medio populi mei habito
2KGS|4|14|et ait quid ergo vult ut faciam ei dixitque Giezi ne quaeras filium enim non habet et vir eius senex est
2KGS|4|15|praecepit itaque ut vocaret eam quae cum vocata fuisset et stetisset ad ostium
2KGS|4|16|dixit ad eam in tempore isto et in hac eadem hora si vita comes fuerit habebis in utero filium at illa respondit noli quaeso domine mi vir Dei noli mentiri ancillae tuae
2KGS|4|17|et concepit mulier et peperit filium in tempore et in hora eadem quam dixerat Heliseus
2KGS|4|18|crevit autem puer et cum esset quaedam dies et egressus isset ad patrem suum ad messores
2KGS|4|19|ait patri suo caput meum caput meum at ille dixit puero tolle et duc eum ad matrem suam
2KGS|4|20|qui cum tulisset et adduxisset eum ad matrem suam posuit eum illa super genua sua usque ad meridiem et mortuus est
2KGS|4|21|ascendit autem et conlocavit eum super lectulum hominis Dei et clusit ostium et egressa
2KGS|4|22|vocavit virum suum et ait mitte mecum obsecro unum de pueris et asinam ut excurram usque ad hominem Dei et revertar
2KGS|4|23|qui ait illi quam ob causam vadis ad eum hodie non sunt kalendae neque sabbatum quae respondit vale
2KGS|4|24|stravitque asinam et praecepit puero mina et propera ne mihi moram facias in eundo et hoc age quod praecipio tibi
2KGS|4|25|profecta est igitur et venit ad virum Dei in montem Carmeli cumque vidisset eam vir Dei de contra ait ad Giezi puerum suum ecce Sunamitis illa
2KGS|4|26|vade ergo in occursum eius et dic ei rectene agitur circa te et circa virum tuum et circa filium tuum quae respondit recte
2KGS|4|27|cumque venisset ad virum Dei in monte adprehendit pedes eius et accessit Giezi ut amoveret eam et ait homo Dei dimitte illam anima enim eius in amaritudine est et Dominus celavit me et non indicavit mihi
2KGS|4|28|quae dixit illi numquid petivi filium a domino meo numquid non dixi tibi ne inludas me
2KGS|4|29|et ille ait ad Giezi accinge lumbos tuos et tolle baculum meum in manu tua et vade si occurrerit tibi homo non salutes eum et si salutaverit te quispiam non respondeas illi et pones baculum meum super faciem pueri
2KGS|4|30|porro mater pueri ait vivit Dominus et vivit anima tua non dimittam te surrexit ergo et secutus est eam
2KGS|4|31|Giezi autem praecesserat eos et posuerat baculum super faciem pueri et non erat vox neque sensus reversusque est in occursum eius et nuntiavit ei dicens non surrexit puer
2KGS|4|32|ingressus est ergo Heliseus domum et ecce puer mortuus iacebat in lectulo eius
2KGS|4|33|ingressusque clusit ostium super se et puerum et oravit ad Dominum
2KGS|4|34|et ascendit et incubuit super puerum posuitque os suum super os eius et oculos suos super oculos eius et manus suas super manus eius et incurvavit se super eum et calefacta est caro pueri
2KGS|4|35|at ille reversus deambulavit in domo semel huc et illuc et ascendit et incubuit super eum et oscitavit puer septies aperuitque oculos
2KGS|4|36|et ille vocavit Giezi et dixit ei voca Sunamitin hanc quae vocata ingressa est ad eum qui ait tolle filium tuum
2KGS|4|37|venit illa et corruit ad pedes eius et adoravit super terram tulitque filium suum et egressa est
2KGS|4|38|et Heliseus reversus est in Galgala erat autem fames in terra et filii prophetarum habitabant coram eo dixitque uni de pueris suis pone ollam grandem et coque pulmentum filiis prophetarum
2KGS|4|39|et egressus est unus in agrum ut colligeret herbas agrestes invenitque quasi vitem silvestrem et collegit ex ea colocyntidas agri et implevit pallium suum et reversus concidit in ollam pulmenti nesciebat enim quid esset
2KGS|4|40|infuderunt ergo sociis ut comederent cumque gustassent de coctione exclamaverunt dicentes mors in olla vir Dei et non potuerunt comedere
2KGS|4|41|at ille adferte inquit farinam et misit in ollam et ait infunde turbae et comedat et non fuit amplius quicquam amaritudinis in olla
2KGS|4|42|vir autem quidam venit de Balsalisa deferens viro Dei panes primitiarum et viginti panes hordiacios et frumentum novum in pera sua at ille dixit da populo ut comedat
2KGS|4|43|responditque ei minister eius quantum est hoc ut adponam coram centum viris rursum ille da ait populo ut comedat haec enim dicit Dominus comedent et supererit
2KGS|4|44|posuit itaque coram eis qui comederunt et superfuit iuxta verbum Domini
2KGS|5|1|Naaman princeps militiae regis Syriae erat vir magnus apud dominum suum et honoratus per illum enim dedit Dominus salutem Syriae erat autem vir fortis et dives sed leprosus
2KGS|5|2|porro de Syria egressi fuerant latrunculi et captivam duxerant de terra Israhel puellam parvulam quae erat in obsequio uxoris Naaman
2KGS|5|3|quae ait ad dominam suam utinam fuisset dominus meus ad prophetam qui est in Samaria profecto curasset eum a lepra quam habet
2KGS|5|4|ingressus est itaque Naaman ad dominum suum et nuntiavit ei dicens sic et sic locuta est puella de terra Israhel
2KGS|5|5|dixitque ei rex Syriae vade et mittam litteras ad regem Israhel qui cum profectus esset et tulisset secum decem talenta argenti et sex milia aureos et decem mutatoria vestimentorum
2KGS|5|6|detulit litteras ad regem Israhel in haec verba cum acceperis epistulam hanc scito quod miserim ad te Naaman servum meum ut cures eum a lepra sua
2KGS|5|7|cumque legisset rex Israhel litteras scidit vestimenta sua et ait numquid Deus sum ut occidere possim et vivificare quia iste misit ad me ut curem hominem a lepra sua animadvertite et videte quod occasiones quaerat adversum me
2KGS|5|8|quod cum audisset Heliseus vir Dei scidisse videlicet regem Israhel vestimenta sua misit ad eum dicens quare scidisti vestimenta tua veniat ad me et sciat esse prophetam in Israhel
2KGS|5|9|venit ergo Naaman cum equis et curribus et stetit ad ostium domus Helisei
2KGS|5|10|misitque ad eum Heliseus nuntium dicens vade et lavare septies in Iordane et recipiet sanitatem caro tua atque mundaberis
2KGS|5|11|iratus Naaman recedebat dicens putabam quod egrederetur ad me et stans invocaret nomen Domini Dei sui et tangeret manu sua locum leprae et curaret me
2KGS|5|12|numquid non meliores sunt Abana et Pharphar fluvii Damasci omnibus aquis Israhel ut laver in eis et munder cum ergo vertisset se et abiret indignans
2KGS|5|13|accesserunt ad eum servi sui et locuti sunt ei pater si rem grandem dixisset tibi propheta certe facere debueras quanto magis quia nunc dixit tibi lavare et mundaberis
2KGS|5|14|descendit et lavit in Iordane septies iuxta sermonem viri Dei et restituta est caro eius sicut caro pueri parvuli et mundatus est
2KGS|5|15|reversusque ad virum Dei cum universo comitatu suo venit et stetit coram eo et ait vere scio quod non sit Deus in universa terra nisi tantum in Israhel obsecro itaque ut accipias benedictionem a servo tuo
2KGS|5|16|at ille respondit vivit Dominus ante quem sto quia non accipiam cumque vim faceret penitus non adquievit
2KGS|5|17|dixitque Naaman ut vis sed obsecro concede mihi servo tuo ut tollam onus duorum burdonum de terra non enim faciet ultra servus tuus holocaustum aut victimam diis alienis nisi Domino
2KGS|5|18|hoc autem solum est de quo depreceris Dominum pro servo tuo quando ingreditur dominus meus templum Remmon ut adoret et illo innitente super manum meam si adoravero in templo Remmon adorante me in eodem loco ut ignoscat mihi Dominus servo tuo pro hac re
2KGS|5|19|qui dixit ei vade in pace abiit ergo ab eo electo terrae tempore
2KGS|5|20|dixitque Giezi puer viri Dei pepercit dominus meus Naaman Syro isti ut non acciperet ab eo quae adtulit vivit Dominus quia curram post eum et accipiam ab eo aliquid
2KGS|5|21|et secutus est Giezi post tergum Naaman quem cum vidisset ille currentem ad se desilivit de curru in occursum eius et ait rectene sunt omnia
2KGS|5|22|et ille ait recte dominus meus misit me dicens modo venerunt ad me duo adulescentes de monte Ephraim ex filiis prophetarum da eis talentum argenti et vestes mutatorias duplices
2KGS|5|23|dixitque Naaman melius est ut accipias duo talenta et coegit eum ligavitque duo talenta argenti in duobus saccis et duplicia vestimenta et inposuit duobus pueris suis qui et portaverunt coram eo
2KGS|5|24|cumque venisset iam vesperi tulit de manu eorum et reposuit in domo dimisitque viros et abierunt
2KGS|5|25|ipse autem ingressus stetit coram domino suo et dixit Heliseus unde venis Giezi qui respondit non ivit servus tuus quoquam
2KGS|5|26|at ille nonne ait cor meum in praesenti erat quando reversus est homo de curru suo in occursum tui nunc igitur accepisti argentum et accepisti vestes ut emas oliveta et vineta et oves et boves et servos et ancillas
2KGS|5|27|sed et lepra Naaman adherebit tibi et semini tuo in sempiternum et egressus est ab eo leprosus quasi nix
2KGS|6|1|dixerunt autem filii prophetarum ad Heliseum ecce locus in quo habitamus coram te angustus est nobis
2KGS|6|2|eamus usque ad Iordanem et tollant singuli de silva materias singulas ut aedificemus nobis ibi locum ad habitandum qui dixit ite
2KGS|6|3|et ait unus ex illis veni ergo et tu cum servis tuis respondit ego veniam
2KGS|6|4|et abiit cum eis cumque venissent ad Iordanem caedebant ligna
2KGS|6|5|accidit autem ut cum unus materiem succidisset caderet ferrum securis in aquam exclamavitque ille et ait eheu eheu eheu domine mi et hoc ipsum mutuo acceperam
2KGS|6|6|dixit autem homo Dei ubi cecidit at ille monstravit ei locum praecidit ergo lignum et misit illuc natavitque ferrum
2KGS|6|7|et ait tolle qui extendit manum et tulit illud
2KGS|6|8|rex autem Syriae pugnabat contra Israhel consiliumque iniit cum servis suis dicens in loco illo et illo ponamus insidias
2KGS|6|9|misit itaque vir Dei ad regem Israhel dicens cave ne transeas in loco illo quia ibi Syri in insidiis sunt
2KGS|6|10|misit rex Israhel ad locum quem dixerat ei vir Dei et praeoccupavit eum et observavit se ibi non semel neque bis
2KGS|6|11|conturbatumque est cor regis Syriae pro hac re et convocatis servis suis ait quare non indicastis mihi quis proditor mei sit apud regem Israhel
2KGS|6|12|dixitque unus servorum eius nequaquam domine mi rex sed Heliseus propheta qui est in Israhel indicat regi Israhel omnia verba quaecumque locutus fueris in conclavi tuo
2KGS|6|13|dixit eis ite et videte ubi sit ut mittam et capiam eum adnuntiaveruntque ei dicentes ecce in Dothan
2KGS|6|14|misit ergo illuc equos et currus et robur exercitus qui cum venissent nocte circumdederunt civitatem
2KGS|6|15|consurgens autem diluculo minister viri Dei egressus est viditque exercitum in circuitu civitatis et equos et currus nuntiavitque ei dicens eheu eheu domine mi quid faciemus
2KGS|6|16|at ille respondit noli timere plures enim nobiscum sunt quam cum illis
2KGS|6|17|cumque orasset Heliseus ait Domine aperi oculos huius ut videat et aperuit Dominus oculos pueri et vidit et ecce mons plenus equorum et curruum igneorum in circuitu Helisei
2KGS|6|18|hostes vero descenderunt ad eum porro Heliseus oravit Dominum dicens percute obsecro gentem hanc caecitate percussitque eos Dominus ne viderent iuxta verbum Helisei
2KGS|6|19|dixit autem ad eos Heliseus non est haec via nec ista est civitas sequimini me et ostendam vobis virum quem quaeritis duxit ergo eos in Samariam
2KGS|6|20|cumque ingressi fuissent in Samaria dixit Heliseus Domine aperi oculos istorum ut videant aperuitque Dominus oculos eorum et viderunt esse se in medio Samariae
2KGS|6|21|dixitque rex Israhel ad Heliseum cum vidisset eos numquid percutiam eos pater mi
2KGS|6|22|at ille ait non percuties neque enim cepisti eos gladio et arcu tuo ut percutias pone panem et aquam coram eis ut comedant et bibant et vadant ad dominum suum
2KGS|6|23|adpositaque est eis ciborum magna praeparatio et comederunt et biberunt et dimisit eos abieruntque ad dominum suum et ultra non venerunt latrones Syriae in terram Israhel
2KGS|6|24|factum est autem post haec congregavit Benadad rex Syriae universum exercitum suum et ascendit et obsidebat Samariam
2KGS|6|25|factaque est fames magna in Samaria et tamdiu obsessa est donec venundaretur caput asini octoginta argenteis et quarta pars cabi stercoris columbarum quinque argenteis
2KGS|6|26|cumque rex Israhel transiret per murum mulier exclamavit ad eum dicens salva me domine mi rex
2KGS|6|27|qui ait non te salvet Dominus unde salvare te possum de area an de torculari dixitque ad eam rex quid tibi vis quae respondit
2KGS|6|28|mulier ista dixit mihi da filium tuum ut comedamus eum hodie et filium meum comedemus cras
2KGS|6|29|coximus ergo filium meum et comedimus dixique ei die altera da filium tuum ut comedamus eum quae abscondit filium suum
2KGS|6|30|quod cum audisset rex scidit vestimenta sua et transiebat super murum viditque omnis populus cilicium quo vestitus erat ad carnem intrinsecus
2KGS|6|31|et ait haec mihi faciat Deus et haec addat si steterit caput Helisei filii Saphat super eum hodie
2KGS|6|32|Heliseus autem sedebat in domo sua et senes sedebant cum eo praemisit itaque virum et antequam veniret nuntius ille dixit ad senes numquid scitis quod miserit filius homicidae hic ut praecidatur caput meum videte ergo cum venerit nuntius cludite ostium et non sinatis eum introire ecce enim sonitus pedum domini eius post eum est
2KGS|6|33|et adhuc illo loquente eis apparuit nuntius qui veniebat ad eum et ait ecce tantum malum a Domino est quid amplius expectabo a Domino
2KGS|7|1|dixit autem Heliseus audite verbum Domini haec dicit Dominus in tempore hoc cras modius similae uno statere erit et duo modii hordei statere uno in porta Samariae
2KGS|7|2|respondens unus de ducibus super cuius manum rex incumbebat homini Dei ait si Dominus fecerit etiam cataractas in caelo numquid poterit esse quod loqueris qui ait videbis oculis tuis et inde non comedes
2KGS|7|3|quattuor ergo viri erant leprosi iuxta introitum portae qui dixerunt ad invicem quid hic esse volumus donec moriamur
2KGS|7|4|sive ingredi voluerimus civitatem fame moriemur sive manserimus hic moriendum nobis est venite igitur et transfugiamus ad castra Syriae si pepercerint nobis vivemus si autem occidere voluerint nihilominus moriemur
2KGS|7|5|surrexerunt igitur vesperi ut venirent ad castra Syriae cumque venissent ad principium castrorum Syriae nullum ibidem reppererunt
2KGS|7|6|siquidem Dominus sonitum audiri fecerat in castris Syriae curruum et equorum et exercitus plurimi dixeruntque ad invicem ecce mercede conduxit adversum nos rex Israhel reges Hettheorum et Aegyptiorum et venerunt super nos
2KGS|7|7|surrexerunt ergo et fugerunt in tenebris et dereliquerunt tentoria sua et equos et asinos in castris fugeruntque animas tantum suas salvare cupientes
2KGS|7|8|igitur cum venissent leprosi illi ad principium castrorum ingressi sunt unum tabernaculum et comederunt et biberunt tuleruntque inde argentum et aurum et vestes et abierunt et absconderunt et rursum reversi sunt ad aliud tabernaculum et inde similiter auferentes absconderunt
2KGS|7|9|dixeruntque ad invicem non recte facimus haec enim dies boni nuntii est si tacuerimus et noluerimus nuntiare usque mane sceleris arguemur venite eamus et nuntiemus in aula regis
2KGS|7|10|cumque venissent ad portam civitatis narraverunt eis dicentes ivimus ad castra Syriae et nullum ibidem repperimus hominum nisi equos et asinos alligatos et fixa tentoria
2KGS|7|11|ierunt ergo portarii et nuntiaverunt in palatio regis intrinsecus
2KGS|7|12|qui surrexit nocte et ait ad servos suos dico vobis quid fecerint nobis Syri sciunt quia fame laboramus et idcirco egressi sunt de castris et latitant in agris dicentes cum egressi fuerint de civitate capiemus eos viventes et tunc civitatem ingredi poterimus
2KGS|7|13|respondit autem unus servorum eius tollamus quinque equos qui remanserunt in urbe quia ipsi tantum sunt in universa multitudine Israhel alii enim consumpti sunt et mittentes explorare poterimus
2KGS|7|14|adduxerunt ergo duos equos misitque rex ad castra Syrorum dicens ite videte
2KGS|7|15|qui abierunt post eos usque ad Iordanem ecce autem omnis via plena erat vestibus et vasis quae proiecerant Syri cum turbarentur reversique nuntii indicaverunt regi
2KGS|7|16|et egressus populus diripuit castra Syriae factusque est modius similae statere uno et duo modii hordei statere uno iuxta verbum Domini
2KGS|7|17|porro rex ducem illum in cuius manu incubuerat constituit ad portam quem conculcavit turba in introitu et mortuus est iuxta quod locutus fuerat vir Dei quando descenderat rex ad eum
2KGS|7|18|factumque est secundum sermonem viri Dei quem dixerat regi quando ait duo modii hordei statere uno erunt et modius similae statere uno hoc eodem tempore cras in porta Samariae
2KGS|7|19|quando responderat dux ille viro Dei et dixerat etiam si Dominus fecerit cataractas in caelo numquid fieri poterit quod loqueris et dixit ei videbis oculis tuis et inde non comedes
2KGS|7|20|evenit ergo ei sicut praedictum erat et conculcavit eum populus in porta et mortuus est
2KGS|8|1|Heliseus autem locutus est ad mulierem cuius vivere fecerat filium dicens surge vade tu et domus tua et peregrinare ubicumque reppereris vocavit enim Dominus famem et veniet super terram septem annis
2KGS|8|2|quae surrexit et fecit iuxta verbum hominis Dei et vadens cum domo sua peregrinata est in terra Philisthim diebus multis
2KGS|8|3|cumque finiti essent anni septem reversa est mulier de terra Philisthim et egressa est ut interpellaret regem pro domo sua et agris suis
2KGS|8|4|rex autem loquebatur cum Giezi puero viri Dei dicens narra mihi omnia magnalia quae fecit Heliseus
2KGS|8|5|cumque ille narraret regi quomodo mortuum suscitasset apparuit mulier cuius vivificaverat filium clamans ad regem pro domo sua et pro agris suis dixitque Giezi domine mi rex haec est mulier et hic filius eius quem suscitavit Heliseus
2KGS|8|6|et interrogavit rex mulierem quae narravit ei deditque ei rex eunuchum unum dicens restitue ei omnia quae sua sunt et universos reditus agrorum a die qua reliquit terram usque ad praesens
2KGS|8|7|venit quoque Heliseus Damascum et Benadad rex Syriae aegrotabat nuntiaveruntque ei dicentes venit vir Dei huc
2KGS|8|8|et ait rex ad Azahel tolle tecum munera et vade in occursum viri Dei et consule Dominum per eum dicens si evadere potero de infirmitate mea hac
2KGS|8|9|ivit igitur Azahel in occursum eius habens secum munera et omnia bona Damasci onera quadraginta camelorum cumque stetisset coram eo ait filius tuus Benadad rex Syriae misit me ad te dicens si sanari potero de infirmitate mea hac
2KGS|8|10|dixitque ei Heliseus vade dic ei sanaberis porro ostendit mihi Dominus quia morte morietur
2KGS|8|11|stetitque cum eo et conturbatus est usque ad suffusionem vultus flevitque vir Dei
2KGS|8|12|cui Azahel ait quare dominus meus flet at ille respondit quia scio quae facturus sis filiis Israhel mala civitates eorum munitas igne succendes et iuvenes eorum interficies gladio et parvulos eorum elides et praegnantes divides
2KGS|8|13|dixitque Azahel quid enim sum servus tuus canis ut faciam rem istam magnam et ait Heliseus ostendit mihi Dominus te regem Syriae fore
2KGS|8|14|qui cum recessisset ab Heliseo venit ad dominum suum qui ait ei quid tibi dixit Heliseus at ille respondit dixit mihi recipiet sanitatem
2KGS|8|15|cumque venisset dies altera tulit sagulum et infudit aqua et expandit super faciem eius quo mortuo regnavit Azahel pro eo
2KGS|8|16|anno quinto Ioram filii Ahab regis Israhel et Iosaphat regis Iuda regnavit Ioram filius Iosaphat rex Iuda
2KGS|8|17|triginta duorum erat annorum cum regnare coepisset et octo annis regnavit in Hierusalem
2KGS|8|18|ambulavitque in viis regum Israhel sicut ambulaverat domus Ahab filia enim Ahab erat uxor eius et fecit quod malum est coram Domino
2KGS|8|19|noluit autem Dominus disperdere Iudam propter David servum suum sicut promiserat ei ut daret illi lucernam et filiis eius cunctis diebus
2KGS|8|20|in diebus eius recessit Edom ne esset sub Iuda et constituit sibi regem
2KGS|8|21|venitque Ioram Seira et omnis currus cum eo et surrexit nocte percussitque Idumeos qui eum circumdederant et principes curruum populus autem fugit in tabernacula sua
2KGS|8|22|recessit ergo Edom ne esset sub Iuda usque ad diem hanc tunc recessit et Lobna in tempore illo
2KGS|8|23|reliqua autem sermonum Ioram et universa quae fecit nonne haec scripta sunt in libro verborum dierum regum Iuda
2KGS|8|24|et dormivit Ioram cum patribus suis sepultusque est cum eis in civitate David et regnavit Ahazias filius eius pro eo
2KGS|8|25|anno duodecimo Ioram filii Ahab regis Israhel regnavit Ahazias filius Ioram regis Iudae
2KGS|8|26|viginti duorum annorum erat Ahazias cum regnare coepisset et uno anno regnavit in Hierusalem nomen matris eius Athalia filia Amri regis Israhel
2KGS|8|27|et ambulavit in viis domus Ahab et fecit quod malum est coram Domino sicut domus Ahab gener enim domus Ahab fuit
2KGS|8|28|abiit quoque cum Ioram filio Ahab ad proeliandum contra Azahel regem Syriae in Ramoth Galaad et vulneraverunt Syri Ioram
2KGS|8|29|qui reversus est ut curaretur in Hiezrahel quia vulneraverant eum Syri in Rama proeliantem contra Azahel regem Syriae porro Ahazias filius Ioram rex Iuda descendit invisere Ioram filium Ahab in Hiezrahel quia aegrotabat
2KGS|9|1|Heliseus autem prophetes vocavit unum de filiis prophetarum et ait illi accinge lumbos tuos et tolle lenticulam olei hanc in manu tua et vade in Ramoth Galaad
2KGS|9|2|cumque veneris illuc videbis Hieu filium Iosaphat filii Namsi et ingressus suscitabis eum de medio fratrum suorum et introduces interius cubiculum
2KGS|9|3|tenensque lenticulam olei fundes super caput eius et dices haec dicit Dominus unxi te regem super Israhel aperiesque ostium et fugies et non ibi subsistes
2KGS|9|4|abiit ergo adulescens puer prophetae Ramoth Galaad
2KGS|9|5|et ingressus est ecce autem principes exercitus sedebant et ait verbum mihi ad te princeps dixitque Hieu ad quem ex omnibus nobis at ille dixit ad te o princeps
2KGS|9|6|et surrexit et ingressus est cubiculum at ille fudit oleum super caput eius et ait haec dicit Dominus Deus Israhel unxi te regem super populum Domini Israhel
2KGS|9|7|et percuties domum Ahab domini tui ut ulciscar sanguinem servorum meorum prophetarum et sanguinem omnium servorum Domini de manu Hiezabel
2KGS|9|8|perdamque omnem domum Ahab et interficiam de Ahab mingentem ad parietem et clausum et novissimum in Israhel
2KGS|9|9|et dabo domum Ahab sicut domum Hieroboam filii Nabath et sicut domum Baasa filii Ahia
2KGS|9|10|Hiezabel quoque comedent canes in agro Hiezrahel nec erit qui sepeliat eam aperuitque ostium et fugit
2KGS|9|11|Hieu autem egressus est ad servos domini sui qui dixerunt ei rectene sunt omnia quid venit insanus iste ad te qui ait eis nostis hominem et quid locutus sit
2KGS|9|12|at illi responderunt falsum est sed magis narra nobis qui ait eis haec et haec locutus est mihi et ait haec dicit Dominus unxi te regem super Israhel
2KGS|9|13|festinaverunt itaque et unusquisque tollens pallium suum posuerunt sub pedibus eius in similitudinem tribunalis et cecinerunt tuba atque dixerunt regnavit Hieu
2KGS|9|14|coniuravit ergo Hieu filius Iosaphat filii Namsi contra Ioram porro Ioram obsederat Ramoth Galaad ipse et omnis Israhel contra Azahel regem Syriae
2KGS|9|15|et reversus fuerat ut curaretur in Hiezrahel propter vulnera quia percusserant eum Syri proeliantem contra Azahel regem Syriae dixitque Hieu si placet vobis nemo egrediatur profugus de civitate ne vadat et nuntiet in Hiezrahel
2KGS|9|16|et ascendit et profectus est in Hiezrahel Ioram enim aegrotabat ibi et Ahazia rex Iuda descenderat ad visitandum Ioram
2KGS|9|17|igitur speculator qui stabat super turrem Hiezrahel vidit globum Hieu venientis et ait video ego globum dixitque Ioram tolle currum et mitte in occursum eorum et dicat vadens rectene sunt omnia
2KGS|9|18|abiit igitur qui ascenderat currum in occursum eius et ait haec dicit rex pacata sunt omnia dixitque ei Hieu quid tibi et paci transi et sequere me nuntiavit quoque speculator dicens venit nuntius ad eos et non revertitur
2KGS|9|19|misit etiam currum equorum secundum venitque ad eos et ait haec dicit rex num pax est et ait Hieu quid tibi et paci transi et sequere me
2KGS|9|20|nuntiavit autem speculator dicens venit usque ad eos et non revertitur est autem incessus quasi incessus Hieu filii Namsi praeceps enim graditur
2KGS|9|21|et ait Ioram iunge currum iunxeruntque currum eius et egressus est Ioram rex Israhel et Ahazias rex Iuda singuli in curribus suis egressique sunt in occursum Hieu et invenerunt eum in agro Naboth Hiezrahelitis
2KGS|9|22|cumque vidisset Ioram Hieu dixit pax est Hieu at ille respondit quae pax adhuc fornicationes Hiezabel matris tuae et veneficia eius multa vigent
2KGS|9|23|convertit autem Ioram manum suam et fugiens ait ad Ahaziam insidiae Ahazia
2KGS|9|24|porro Hieu tetendit arcum manu et percussit Ioram inter scapulas et egressa est sagitta per cor eius statimque corruit in curru suo
2KGS|9|25|dixitque Hieu ad Baddacer ducem tolle proice eum in agro Naboth Hiezrahelitae memini enim quando ego et tu sedentes in curru sequebamur Ahab patrem huius quod Dominus onus hoc levaverit super eum dicens
2KGS|9|26|si non pro sanguine Naboth et pro sanguine filiorum eius quem vidi heri ait Dominus reddam tibi in agro isto dicit Dominus nunc igitur tolle proice eum in agro iuxta verbum Domini
2KGS|9|27|Ahazias autem rex Iuda videns hoc fugit per viam domus horti persecutusque est eum Hieu et ait etiam hunc percutite in curru suo in ascensu Gaber qui est iuxta Ieblaam qui fugit in Mageddo et mortuus est ibi
2KGS|9|28|et inposuerunt eum servi eius super currum suum et tulerunt Hierusalem sepelieruntque in sepulchro cum patribus suis in civitate David
2KGS|9|29|anno undecimo Ioram filii Ahab rege Ahazia super Iudam
2KGS|9|30|venit Hieu Hiezrahel porro Hiezabel introitu eius audito depinxit oculos suos stibio et ornavit caput suum et respexit per fenestram
2KGS|9|31|ingredientem Hieu per portam et ait numquid pax esse potest Zamri qui interfecit dominum suum
2KGS|9|32|levavitque Hieu faciem suam ad fenestram et ait quae est ista et inclinaverunt se ad eum duo vel tres eunuchi
2KGS|9|33|at ille dixit eis praecipitate eam deorsum et praecipitaverunt eam aspersusque est sanguine paries et equorum ungulae qui conculcaverunt eam
2KGS|9|34|cumque ingressus esset et comederet bibissetque ait ite videte maledictam illam et sepelite eam quia filia regis est
2KGS|9|35|cumque issent ut sepelirent eam non invenerunt nisi calvariam et pedes et summas manus
2KGS|9|36|reversique nuntiaverunt ei et ait Hieu sermo Domini est quem locutus est per servum suum Heliam Thesbiten dicens in agro Hiezrahel comedent canes carnes Hiezabel
2KGS|9|37|et erunt carnes Hiezabel sicut stercus super faciem terrae in agro Hiezrahel ita ut praetereuntes dicant haecine est illa Hiezabel
2KGS|10|1|erant autem Ahab septuaginta filii in Samaria scripsit ergo Hieu litteras et misit in Samariam ad optimates civitatis et ad maiores natu et ad nutricios Ahab dicens
2KGS|10|2|statim ut acceperitis litteras has qui habetis filios domini vestri et currus et equos et civitates firmas et arma
2KGS|10|3|eligite meliorem et eum qui vobis placuerit de filiis domini vestri et ponite eum super solium patris sui et pugnate pro domo domini vestri
2KGS|10|4|timuerunt illi vehementer et dixerunt ecce duo reges non potuerunt stare coram eo et quomodo nos valebimus resistere
2KGS|10|5|miserunt ergo praepositus domus et praefectus civitatis et maiores natu et nutricii ad Hieu dicentes servi tui sumus quaecumque iusseris faciemus nec constituemus regem quodcumque tibi placet fac
2KGS|10|6|rescripsit autem eis litteras secundo dicens si mei estis et oboeditis mihi tollite capita filiorum domini vestri et venite ad me hac eadem hora cras in Hiezrahel porro filii regis septuaginta viri apud optimates civitatis nutriebantur
2KGS|10|7|cumque venissent litterae ad eos tulerunt filios regis et occiderunt septuaginta viros et posuerunt capita eorum in cofinis et miserunt ad eum in Hiezrahel
2KGS|10|8|venit autem nuntius et indicavit ei dicens adtulerunt capita filiorum regis qui respondit ponite ea duos acervos iuxta introitum portae usque mane
2KGS|10|9|cumque diluxisset egressus est et stans dixit ad omnem populum iusti estis si ego coniuravi contra dominum meum et interfeci eum quis percussit omnes hos
2KGS|10|10|videte ergo nunc quoniam non cecidit de sermonibus Domini in terram quos locutus est Dominus super domum Ahab et Dominus fecit quod locutus est in manu servi sui Heliae
2KGS|10|11|percussit igitur Hieu omnes qui reliqui erant de domo Ahab in Hiezrahel et universos optimates eius et notos et sacerdotes donec non remanerent ex eo reliquiae
2KGS|10|12|et surrexit et venit in Samariam cumque venisset ad Camaram pastorum in via
2KGS|10|13|invenit fratres Ahaziae regis Iuda dixitque ad eos quinam estis vos at illi responderunt fratres Ahaziae sumus et descendimus ad salutandos filios regis et filios reginae
2KGS|10|14|qui ait conprehendite eos vivos quos cum conprehendissent vivos iugulaverunt eos in cisterna iuxta Camaram quadraginta duos viros et non reliquit ex eis quemquam
2KGS|10|15|cumque abisset inde invenit Ionadab filium Rechab in occursum sibi et benedixit ei et ait ad eum numquid est cor tuum rectum sicut cor meum cum corde tuo et ait Ionadab est si est inquit da manum tuam qui dedit manum suam at ille levavit eum ad se in curru
2KGS|10|16|dixitque ad eum veni mecum et vide zelum meum pro Domino et inpositum currui suo
2KGS|10|17|duxit in Samariam et percussit omnes qui reliqui fuerant de Ahab in Samaria usque ad unum iuxta verbum Domini quod locutus est per Heliam
2KGS|10|18|congregavit ergo Hieu omnem populum et dixit ad eos Ahab coluit Baal parum ego autem colam eum amplius
2KGS|10|19|nunc igitur omnes prophetas Baal et universos servos eius et cunctos sacerdotes ipsius vocate ad me nullus sit qui non veniat sacrificium enim grande est mihi Baal quicumque defuerit non vivet porro Hieu faciebat hoc insidiose ut disperderet cultores Baal
2KGS|10|20|dixit sanctificate diem sollemnem Baal vocavitque
2KGS|10|21|et misit in universos terminos Israhel et venerunt cuncti servi Baal non fuit residuus ne unus quidem qui non veniret et ingressi sunt templum Baal et repleta est domus Baal a summo usque ad summum
2KGS|10|22|dixitque his qui erant super vestes proferte vestimenta universis servis Baal et protulerunt eis vestes
2KGS|10|23|ingressusque Hieu et Ionadab filius Rechab templum Baal et ait cultoribus Baal perquirite et videte ne quis forte vobiscum sit de servis Domini sed ut sint soli servi Baal
2KGS|10|24|ingressi sunt igitur ut facerent victimas et holocausta Hieu autem praeparaverat sibi foris octoginta viros et dixerat eis quicumque fugerit de hominibus his quos ego adduxero in manus vestras anima eius erit pro anima illius
2KGS|10|25|factum est ergo cum conpletum esset holocaustum praecepit Hieu militibus et ducibus suis ingredimini et percutite eos nullus evadat percusseruntque eos ore gladii et proiecerunt milites et duces et ierunt in civitatem templi Baal
2KGS|10|26|et protulerunt statuam de fano Baal et conbuserunt
2KGS|10|27|et comminuerunt eam destruxerunt quoque aedem Baal et fecerunt pro ea latrinas usque ad diem hanc
2KGS|10|28|delevit itaque Hieu Baal de Israhel
2KGS|10|29|verumtamen a peccatis Hieroboam filii Nabath qui peccare fecerat Israhel non recessit nec dereliquit vitulos aureos qui erant in Bethel et in Dan
2KGS|10|30|dixit autem Dominus ad Hieu quia studiose fecisti quod rectum erat et placebat in oculis meis et omnia quae erant in corde meo fecisti contra domum Ahab filii tui usque ad quartam generationem sedebunt super thronum Israhel
2KGS|10|31|porro Hieu non custodivit ut ambularet in lege Domini Dei Israhel in toto corde suo non enim recessit a peccatis Hieroboam qui peccare fecerat Israhel
2KGS|10|32|in diebus illis coepit Dominus taedere super Israhel percussitque eos Azahel in universis finibus Israhel
2KGS|10|33|a Iordane contra orientalem plagam omnem terram Galaad et Gad et Ruben et Manasse ab Aroer quae est super torrentem Arnon et Galaad et Basan
2KGS|10|34|reliqua autem verborum Hieu et universa quae fecit et fortitudo eius nonne haec scripta sunt in libro verborum dierum regum Israhel
2KGS|10|35|et dormivit Hieu cum patribus suis sepelieruntque eum in Samaria et regnavit Ioachaz filius eius pro eo
2KGS|10|36|dies autem quos regnavit Hieu super Israhel viginti et octo anni sunt in Samaria
2KGS|11|1|Athalia vero mater Ahaziae videns mortuum filium suum surrexit et interfecit omne semen regium
2KGS|11|2|tollens autem Iosaba filia regis Ioram soror Ahaziae Ioas filium Ahaziae furata est eum de medio filiorum regis qui interficiebantur et nutricem eius de triclinio et abscondit eum a facie Athaliae ut non interficeretur
2KGS|11|3|eratque cum ea in domo Domini clam sex annis porro Athalia regnavit super terram
2KGS|11|4|anno autem septimo misit Ioiada et adsumens centuriones et milites introduxit ad se in templum Domini pepigitque cum eis foedus et adiurans eos in domo Domini ostendit eis filium regis
2KGS|11|5|et praecepit illis dicens iste sermo quem facere debetis
2KGS|11|6|tertia pars vestrum introeat sabbato et observet excubitum domus regis tertia autem pars sit ad portam Sir et tertia pars ad portam quae est post habitaculum scutariorum et custodietis excubitum domus Messa
2KGS|11|7|duae vero partes e vobis omnes egredientes sabbato custodiant excubias domus Domini circum regem
2KGS|11|8|et vallabitis eum habentes arma in manibus vestris si quis autem ingressus fuerit septum templi interficiatur eritisque cum rege introeunte et egrediente
2KGS|11|9|et fecerunt centuriones iuxta omnia quae praeceperat eis Ioiada sacerdos et adsumentes singuli viros suos qui ingrediebantur sabbatum cum his qui egrediebantur e sabbato venerunt ad Ioiada sacerdotem
2KGS|11|10|qui dedit eis hastas et arma regis David quae erant in domo Domini
2KGS|11|11|et steterunt singuli habentes arma in manu sua a parte templi dextra usque ad partem sinistram altaris et aedis circum regem
2KGS|11|12|produxitque filium regis et posuit super eum diadema et testimonium feceruntque eum regem et unxerunt et plaudentes manu dixerunt vivat rex
2KGS|11|13|audivit Athalia vocem currentis populi et ingressa ad turbas in templum Domini
2KGS|11|14|vidit regem stantem super tribunal iuxta morem et cantores et tubas propter eum omnemque populum terrae laetantem et canentem tubis et scidit vestimenta sua clamavitque coniuratio coniuratio
2KGS|11|15|praecepit autem Ioiada centurionibus qui erant super exercitum et ait eis educite eam extra consepta templi et quicumque secutus eam fuerit feriatur gladio dixerat enim sacerdos non occidatur in templo Domini
2KGS|11|16|inposueruntque ei manus et inpegerunt eam per viam introitus equorum iuxta palatium et interfecta est ibi
2KGS|11|17|pepigit igitur Ioiada foedus inter Dominum et inter regem et inter populum ut esset populus Domini et inter regem et populum
2KGS|11|18|ingressusque est omnis populus terrae templum Baal et destruxerunt aras eius et imagines contriverunt valide Matthan quoque sacerdotem Baal occiderunt coram altari et posuit sacerdos custodias in domo Domini
2KGS|11|19|tulitque centuriones et Cherethi et Felethi legiones et omnem populum terrae deduxeruntque regem de domo Domini et venerunt per viam portae scutariorum in palatium et sedit super thronum regum
2KGS|11|20|laetatusque est omnis populus terrae et civitas conquievit Athalia autem occisa est gladio in domo regis
2KGS|11|21|septemque annorum erat Ioas cum regnare coepisset
2KGS|12|1|anno septimo Hieu regnavit Ioas quadraginta annis regnavit in Hierusalem nomen matris eius Sebia de Bersabee
2KGS|12|2|fecitque Ioas rectum coram Domino cunctis diebus quibus docuit eum Ioiada sacerdos
2KGS|12|3|verumtamen excelsa non abstulit adhuc populus immolabat et adolebat in excelsis incensum
2KGS|12|4|dixitque Ioas ad sacerdotes omnem pecuniam sanctorum quae inlata fuerit in templum Domini a praetereuntibus quae offertur pro pretio animae et quam sponte et arbitrio cordis sui inferunt in templum Domini
2KGS|12|5|accipiant illam sacerdotes iuxta ordinem suum et instaurent sarta tecta domus si quid necessarium viderint instauratione
2KGS|12|6|igitur usque ad vicesimum tertium annum regis Ioas non instauraverunt sacerdotes sarta tecta templi
2KGS|12|7|vocavitque rex Ioas Ioiada pontificem et sacerdotes dicens eis quare sarta tecta non instaurastis templi nolite ergo amplius accipere pecuniam iuxta ordinem vestrum sed ad instaurationem templi reddite eam
2KGS|12|8|prohibitique sunt sacerdotes ultra accipere pecuniam a populo et instaurare sarta tecta domus
2KGS|12|9|et tulit Ioiada pontifex gazofilacium unum aperuitque foramen desuper et posuit illud iuxta altare ad dexteram ingredientium domum Domini mittebantque in eo sacerdotes qui custodiebant ostia omnem pecuniam quae deferebatur ad templum Domini
2KGS|12|10|cumque viderent nimiam pecuniam esse in gazofilacio ascendebat scriba regis et pontifex effundebantque et numerabant pecuniam quae inveniebatur in domo Domini
2KGS|12|11|et dabant eam iuxta numerum atque mensuram in manu eorum qui praeerant cementariis domus Domini qui inpendebant eam in fabris lignorum et in cementariis his qui operabantur in domo Domini
2KGS|12|12|et sarta tecta faciebant et in his qui caedebant saxa et ut emerent ligna et lapides qui excidebantur ita ut impleretur instauratio domus Domini in universis quae indigebant expensa ad muniendam domum
2KGS|12|13|verumtamen non fiebant ex eadem pecunia hydriae templi Domini et fuscinulae et turibula et tubae omne vas aureum et argenteum de pecunia quae inferebatur in templum Domini
2KGS|12|14|his enim qui faciebant opus dabatur ut instauraretur templum Domini
2KGS|12|15|et non fiebat ratio his hominibus qui accipiebant pecuniam ut distribuerent eam artificibus sed in fide tractabant eam
2KGS|12|16|pecuniam vero pro delicto et pecuniam pro peccatis non inferebant in templum Domini quia sacerdotum erat
2KGS|12|17|tunc ascendit Azahel rex Syriae et pugnabat contra Geth cepitque eam et direxit faciem suam ut ascenderet in Hierusalem
2KGS|12|18|quam ob rem tulit Ioas rex Iuda omnia sanctificata quae consecraverant Iosaphat et Ioram et Ahazia patres eius reges Iuda et quae ipse obtulerat et universum argentum quod inveniri potuit in thesauris templi Domini et in palatio regis misitque Azaheli regi Syriae et recessit ab Hierusalem
2KGS|12|19|reliqua autem sermonum Ioas et universa quae fecit nonne haec scripta sunt in libro verborum dierum regum Iuda
2KGS|12|20|surrexerunt autem servi eius et coniuraverunt inter se percusseruntque Ioas in domo Mello in descensu Sela
2KGS|12|21|Iozachar namque filius Semath et Iozabad filius Somer servi eius percusserunt eum et mortuus est et sepelierunt eum cum patribus suis in civitate David regnavitque Amasias filius eius pro eo
2KGS|13|1|anno vicesimo tertio Ioas filii Ahaziae regis Iudae regnavit Ioachaz filius Hieu super Israhel in Samaria decem et septem annis
2KGS|13|2|et fecit malum coram Domino secutusque est peccata Hieroboam filii Nabath qui peccare fecit Israhel non declinavit ab eis
2KGS|13|3|iratusque est furor Domini contra Israhel et tradidit eos in manu Azahelis regis Syriae et in manu Benadad filii Azahel cunctis diebus
2KGS|13|4|deprecatus est autem Ioachaz faciem Domini et audivit eum Dominus vidit enim angustiam Israhel qua adtriverat eos rex Syriae
2KGS|13|5|et dedit Dominus Israheli salvatorem et liberatus est de manu Syriae habitaveruntque filii Israhel in tabernaculis suis sicut heri et nudius tertius
2KGS|13|6|verumtamen non recesserunt a peccatis domus Hieroboam qui peccare fecit Israhel in ipsis ambulaverunt siquidem et lucus permansit in Samaria
2KGS|13|7|et non sunt derelicti Ioachaz de populo nisi quinquaginta equites et decem currus et decem milia peditum interfecerat enim eos rex Syriae et redegerat quasi pulverem in tritura areae
2KGS|13|8|reliqua autem sermonum Ioachaz et universa quae fecit sed et fortitudo eius nonne haec scripta sunt in libro sermonum dierum regum Israhel
2KGS|13|9|dormivitque Ioachaz cum patribus suis et sepelierunt eum in Samaria regnavitque Ioas filius eius pro eo
2KGS|13|10|anno tricesimo septimo Ioas regis Iuda regnavit Ioas filius Ioachaz super Israhel in Samaria sedecim annis
2KGS|13|11|et fecit quod malum est in conspectu Domini non declinavit ab omnibus peccatis Hieroboam filii Nabath qui peccare fecit Israhel in ipsis ambulavit
2KGS|13|12|reliqua autem sermonum Ioas et universa quae fecit sed et fortitudo eius quomodo pugnaverit contra Amasiam regem Iuda nonne haec scripta sunt in libro sermonum regum Israhel
2KGS|13|13|et dormivit Ioas cum patribus suis Hieroboam autem sedit super solium eius porro Ioas sepultus est in Samaria cum regibus Israhel
2KGS|13|14|Heliseus autem aegrotabat infirmitate qua et mortuus est descenditque ad eum Ioas rex Israhel et flebat coram eo dicebatque pater mi pater mi currus Israhel et auriga eius
2KGS|13|15|et ait illi Heliseus adfer arcum et sagittas cumque adtulisset ad eum arcum et sagittas
2KGS|13|16|dixit ad regem Israhel pone manum tuam super arcum et cum posuisset ille manum suam superposuit Heliseus manus suas manibus regis
2KGS|13|17|et ait aperi fenestram orientalem cumque aperuisset dixit Heliseus iace sagittam et iecit et ait Heliseus sagitta salutis Domini et sagitta salutis contra Syriam percutiesque Syriam in Afec donec consumas eam
2KGS|13|18|et ait tolle sagittas qui cum tulisset rursum dixit ei percute iaculo terram et cum percussisset tribus vicibus et stetisset
2KGS|13|19|iratus est contra eum vir Dei et ait si percussisses quinquies aut sexies sive septies percussisses Syriam usque ad consummationem nunc autem tribus vicibus percuties eam
2KGS|13|20|mortuus est ergo Heliseus et sepelierunt eum latrunculi quoque de Moab venerunt in terra in ipso anno
2KGS|13|21|quidam autem sepelientes hominem viderunt latrunculos et proiecerunt cadaver in sepulchro Helisei quod ambulavit et tetigit ossa Helisei et revixit homo et stetit super pedes suos
2KGS|13|22|igitur Azahel rex Syriae adflixit Israhel cunctis diebus Ioachaz
2KGS|13|23|et misertus est Dominus eorum et reversus est ad eos propter pactum suum quod habebat cum Abraham Isaac et Iacob et noluit disperdere eos neque proicere penitus usque in praesens tempus
2KGS|13|24|mortuus est autem Azahel rex Syriae et regnavit Benadad filius eius pro eo
2KGS|13|25|porro Ioas filius Ioachaz tulit urbes de manu Benadad filii Azahel quas tulerat de manu Ioachaz patris sui iure proelii tribus vicibus percussit eum Ioas et reddidit civitates Israheli
2KGS|14|1|anno secundo Ioas filii Ioachaz regis Israhel regnavit Amasias filius Ioas regis Iuda
2KGS|14|2|viginti quinque annorum erat cum regnare coepisset viginti autem et novem annis regnavit in Hierusalem nomen matris eius Ioaden de Hierusalem
2KGS|14|3|et fecit rectum coram Domino verumtamen non ut David pater eius iuxta omnia quae fecit Ioas pater suus fecit
2KGS|14|4|nisi hoc tantum quod excelsa non abstulit adhuc enim populus immolabat et adolebat in excelsis
2KGS|14|5|cumque obtinuisset regnum percussit servos suos qui interfecerant regem patrem suum
2KGS|14|6|filios autem eorum qui occiderant non occidit iuxta quod scriptum est in libro legis Mosi sicut praecepit Dominus dicens non morientur patres pro filiis neque filii morientur pro patribus sed unusquisque in peccato suo morietur
2KGS|14|7|ipse percussit Edom in valle Salinarum decem milia et adprehendit Petram in proelio vocavitque nomen eius Iecethel usque in praesentem diem
2KGS|14|8|tunc misit Amasias nuntios ad Ioas filium Ioachaz filii Hieu regis Israhel dicens veni et videamus nos
2KGS|14|9|remisitque Ioas rex Israhel ad Amasiam regem Iuda dicens carduus Libani misit ad cedrum quae est in Libano dicens da filiam tuam filio meo uxorem transieruntque bestiae saltus quae sunt in Libano et conculcaverunt carduum
2KGS|14|10|percutiens invaluisti super Edom et sublevavit te cor tuum contentus esto gloria et sede in domo tua quare provocas malum ut cadas tu et Iuda tecum
2KGS|14|11|et non adquievit Amasias ascenditque Ioas rex Israhel et viderunt se ipse et Amasias rex Iuda in Bethsames oppido Iudae
2KGS|14|12|percussusque est Iuda coram Israhel et fugerunt unusquisque in tabernacula sua
2KGS|14|13|Amasiam vero regem Iuda filium Ioas filii Ahaziae cepit Ioas rex Israhel in Bethsames et adduxit eum in Hierusalem et interrupit murum Hierusalem a porta Ephraim usque ad portam Anguli quadringentis cubitis
2KGS|14|14|tulitque omne aurum et argentum et universa vasa quae inventa sunt in domo Domini et in thesauris regis et obsides et reversus est Samariam
2KGS|14|15|reliqua autem verborum Ioas quae fecit et fortitudo eius qua pugnavit contra Amasiam regem Iuda nonne haec scripta sunt in libro sermonum dierum regum Israhel
2KGS|14|16|dormivitque Ioas cum patribus suis et sepultus est in Samaria cum regibus Israhel et regnavit Hieroboam filius eius pro eo
2KGS|14|17|vixit autem Amasias filius Ioas rex Iuda postquam mortuus est Ioas filius Ioachaz regis Israhel viginti quinque annis
2KGS|14|18|reliqua autem sermonum Amasiae nonne haec scripta sunt in libro sermonum dierum regum Iuda
2KGS|14|19|factaque est contra eum coniuratio in Hierusalem at ille fugit in Lachis miseruntque post eum in Lachis et interfecerunt eum ibi
2KGS|14|20|et asportaverunt in equis sepultusque est in Hierusalem cum patribus suis in civitate David
2KGS|14|21|tulit autem universus populus Iudae Azariam annos natum sedecim et constituerunt eum regem pro patre eius Amasia
2KGS|14|22|ipse aedificavit Ahilam et restituit eam Iudae postquam dormivit rex cum patribus suis
2KGS|14|23|anno quintodecimo Amasiae filii Ioas regis Iuda regnavit Hieroboam filius Ioas regis Israhel in Samaria quadraginta et uno anno
2KGS|14|24|et fecit quod malum est coram Domino non recessit ab omnibus peccatis Hieroboam filii Nabath qui peccare fecit Israhel
2KGS|14|25|ipse restituit terminos Israhel ab introitu Emath usque ad mare Solitudinis iuxta sermonem Domini Dei Israhel quem locutus est per servum suum Ionam filium Amathi prophetam qui erat de Geth quae est in Opher
2KGS|14|26|vidit enim Dominus adflictionem Israhel amaram nimis et quod consumpti essent usque ad clausos carcere et extremos et non esset qui auxiliaretur Israhel
2KGS|14|27|nec locutus est Dominus ut deleret nomen Israhel sub caelo sed salvavit eos in manu Hieroboam filii Ioas
2KGS|14|28|reliqua autem sermonum Hieroboam et universa quae fecit et fortitudo eius qua proeliatus est et quomodo restituit Damascum et Emath Iudae in Israhel nonne haec scripta sunt in libro sermonum dierum regum Israhel
2KGS|14|29|dormivitque Hieroboam cum patribus suis regibus Israhel et regnavit Zaccharias filius eius pro eo
2KGS|15|1|anno vicesimo septimo Hieroboam regis Israhel regnavit Azarias filius Amasiae regis Iudae
2KGS|15|2|sedecim annorum erat cum regnare coepisset et quinquaginta duobus annis regnavit in Hierusalem nomen matris eius Iecelia de Hierusalem
2KGS|15|3|fecitque quod erat placitum coram Domino iuxta omnia quae fecit Amasias pater eius
2KGS|15|4|verumtamen excelsa non est demolitus adhuc populus sacrificabat et adolebat incensum in excelsis
2KGS|15|5|percussit autem Dominus regem et fuit leprosus usque in diem mortis suae et habitabat in domo libera seorsum Ioatham vero filius regis gubernabat palatium et iudicabat populum terrae
2KGS|15|6|reliqua autem sermonum Azariae et universa quae fecit nonne haec scripta sunt in libro verborum dierum regum Iuda
2KGS|15|7|et dormivit Azarias cum patribus suis sepelieruntque eum cum maioribus suis in civitate David et regnavit Ioatham filius eius pro eo
2KGS|15|8|anno tricesimo octavo Azariae regis Iudae regnavit Zaccharias filius Hieroboam super Israhel in Samaria sex mensibus
2KGS|15|9|et fecit quod malum est coram Domino sicut fecerant patres eius non recessit a peccatis Hieroboam filii Nabath qui peccare fecit Israhel
2KGS|15|10|coniuravit autem contra eum Sellum filius Iabes percussitque eum palam et interfecit regnavitque pro eo
2KGS|15|11|reliqua autem verborum Zacchariae nonne haec scripta sunt in libro sermonum dierum regum Israhel
2KGS|15|12|ipse est sermo Domini quem locutus est ad Hieu dicens filii usque ad quartam generationem sedebunt de te super thronum Israhel factumque est ita
2KGS|15|13|Sellum filius Iabes regnavit tricesimo nono anno Azariae regis Iudae regnavit autem uno mense in Samaria
2KGS|15|14|et ascendit Manahem filius Gaddi de Thersa venitque Samariam et percussit Sellum filium Iabes in Samaria et interfecit eum regnavitque pro eo
2KGS|15|15|reliqua autem verborum Sellum et coniuratio eius per quam tetendit insidias nonne haec scripta sunt in libro sermonum dierum regum Israhel
2KGS|15|16|tunc percussit Manahem Thapsam et omnes qui erant in ea et terminos eius de Thersa noluerant enim aperire ei et interfecit omnes praegnantes eius et scidit eas
2KGS|15|17|anno tricesimo nono Azariae regis Iuda regnavit Manahem filius Gaddi super Israhel decem annis in Samaria
2KGS|15|18|fecitque quod erat malum coram Domino non recessit a peccatis Hieroboam filii Nabath qui peccare fecit Israhel cunctis diebus eius
2KGS|15|19|veniebat Phul rex Assyriorum in terram et dabat Manahem Phul mille talenta argenti ut esset ei in auxilio et firmaret regnum eius
2KGS|15|20|indixitque Manahem argentum super Israhel cunctis potentibus et divitibus ut daret regi Assyriorum quinquaginta siclos argenti per singulos reversusque est rex Assyriorum et non est moratus in terra
2KGS|15|21|reliqua autem sermonum Manahem et universa quae fecit nonne haec scripta sunt in libro sermonum dierum regum Israhel
2KGS|15|22|et dormivit Manahem cum patribus suis regnavitque Phaceia filius eius pro eo
2KGS|15|23|anno quinquagesimo Azariae regis Iudae regnavit Phaceia filius Manahem super Israhel in Samaria biennio
2KGS|15|24|et fecit quod erat malum coram Domino non recessit a peccatis Hieroboam filii Nabath qui peccare fecit Israhel
2KGS|15|25|coniuravit autem adversum eum Phacee filius Romeliae dux eius et percussit eum in Samaria in turre domus regiae iuxta Argob et iuxta Ari et cum eo quinquaginta viros de filiis Galaaditarum et interfecit eum regnavitque pro eo
2KGS|15|26|reliqua autem sermonum Phaceia et universa quae fecit nonne haec scripta sunt in libro sermonum dierum regum Israhel
2KGS|15|27|anno quinquagesimo secundo Azariae regis Iudae regnavit Phacee filius Romeliae super Israhel in Samaria viginti annis
2KGS|15|28|et fecit quod malum erat coram Domino non recessit a peccatis Hieroboam filii Nabath qui peccare fecit Israhel
2KGS|15|29|in diebus Phacee regis Israhel venit Theglathfalassar rex Assur et cepit Aiom et Abel domum Maacha et Ianoe et Cedes et Asor et Galaad et Galileam universam terram Nepthalim et transtulit eos in Assyrios
2KGS|15|30|coniuravit autem et tetendit insidias Osee filius Hela contra Phacee filium Romeliae et percussit eum et interfecit regnavitque pro eo vicesimo anno Ioatham filii Oziae
2KGS|15|31|reliqua autem sermonum Phacee et universa quae fecit nonne haec scripta sunt in libro sermonum dierum regum Israhel
2KGS|15|32|anno secundo Phacee filii Romeliae regis Israhel regnavit Ioatham filius Oziae regis Iuda
2KGS|15|33|viginti quinque annorum erat cum regnare coepisset et sedecim annis regnavit in Hierusalem nomen matris eius Hierusa filia Sadoc
2KGS|15|34|fecitque quod erat placitum coram Domino iuxta omnia quae fecerat Ozias pater suus operatus est
2KGS|15|35|verumtamen excelsa non abstulit adhuc populus immolabat et adolebat incensum in excelsis ipse aedificavit portam domus Domini sublimissimam
2KGS|15|36|reliqua autem sermonum Ioatham et universa quae fecit nonne haec scripta sunt in libro verborum dierum regum Iuda
2KGS|15|37|in diebus illis coepit Dominus mittere in Iudam Rasin regem Syriae et Phacee filium Romeliae
2KGS|15|38|et dormivit Ioatham cum patribus suis sepultusque est cum eis in civitate David patris sui et regnavit Ahaz filius eius pro eo
2KGS|16|1|anno septimodecimo Phacee filii Romeliae regnavit Ahaz filius Ioatham regis Iuda
2KGS|16|2|viginti annorum erat Ahaz cum regnare coepisset et sedecim annis regnavit in Hierusalem non fecit quod erat placitum in conspectu Domini Dei sui sicut David pater eius
2KGS|16|3|sed ambulavit in via regum Israhel insuper et filium suum consecravit transferens per ignem secundum idola gentium quae dissipavit Dominus coram filiis Israhel
2KGS|16|4|immolabat quoque victimas et adolebat incensum in excelsis et in collibus et sub omni ligno frondoso
2KGS|16|5|tunc ascendit Rasin rex Syriae et Phacee filius Romeliae rex Israhel in Hierusalem ad proeliandum cumque obsiderent Ahaz non valuerunt superare eum
2KGS|16|6|in tempore illo restituit Rasin rex Syriae Ahilam Syriae et eiecit Iudaeos de Ahilam et Idumei venerunt in Ahilam et habitaverunt ibi usque in diem hanc
2KGS|16|7|misit autem Ahaz nuntios ad Theglathfalassar regem Assyriorum dicens servus tuus et filius tuus ego sum ascende et salvum me fac de manu regis Syriae et de manu regis Israhel qui consurrexerunt adversum me
2KGS|16|8|et cum collegisset argentum et aurum quod invenire potuit in domo Domini et in thesauris regis misit regi Assyriorum munera
2KGS|16|9|qui et adquievit voluntati eius ascendit enim rex Assyriorum in Damascum et vastavit eam et transtulit habitatores eius Cyrenen Rasin autem interfecit
2KGS|16|10|perrexitque rex Ahaz in occursum Theglathfalassar regis Assyriorum in Damascum cumque vidisset altare Damasci misit rex Ahaz ad Uriam sacerdotem exemplar eius et similitudinem iuxta omne opus eius
2KGS|16|11|extruxitque Urias sacerdos altare iuxta omnia quae praeceperat rex Ahaz de Damasco ita fecit Urias sacerdos donec veniret rex Ahaz de Damasco
2KGS|16|12|cumque venisset rex de Damasco vidit altare et veneratus est illud ascenditque et immolavit holocausta et sacrificium suum
2KGS|16|13|et libavit libamina et fudit sanguinem pacificorum quae obtulerat super altare
2KGS|16|14|porro altare aeneum quod erat coram Domino transtulit de facie templi et de loco altaris et de loco templi Domini posuitque illud ex latere altaris ad aquilonem
2KGS|16|15|praecepit quoque rex Ahaz Uriae sacerdoti dicens super altare maius offer holocaustum matutinum et sacrificium vespertinum et holocaustum regis et sacrificium eius et holocaustum universi populi terrae et sacrificia eorum et libamina eorum et omnem sanguinem holocausti et universum sanguinem victimae super illud effundes altare vero aeneum erit paratum ad voluntatem meam
2KGS|16|16|fecit igitur Urias sacerdos iuxta omnia quae praeceperat rex Ahaz
2KGS|16|17|tulit autem rex Ahaz celatas bases et luterem qui erat desuper et mare deposuit de bubus aeneis qui sustentabant illud et posuit super pavimentum stratum lapide
2KGS|16|18|Musach quoque sabbati quod aedificaverat in templo et ingressum regis exterius convertit in templo Domini propter regem Assyriorum
2KGS|16|19|reliqua autem verborum Ahaz quae fecit nonne haec scripta sunt in libro sermonum dierum regum Iuda
2KGS|16|20|dormivitque Ahaz cum patribus suis et sepultus est cum eis in civitate David et regnavit Ezechias filius eius pro eo
2KGS|17|1|anno duodecimo Ahaz regis Iuda regnavit Osee filius Hela in Samaria super Israhel novem annis
2KGS|17|2|fecitque malum coram Domino sed non sicut reges Israhel qui ante eum fuerant
2KGS|17|3|contra hunc ascendit Salmanassar rex Assyriorum et factus est ei Osee servus reddebatque illi tributa
2KGS|17|4|cumque deprehendisset rex Assyriorum Osee quod rebellare nitens misisset nuntios ad Sua regem Aegypti ne praestaret tributa regi Assyriorum sicut singulis annis solitus erat obsedit eum et vinctum misit in carcerem
2KGS|17|5|pervagatusque est omnem terram et ascendens Samariam obsedit eam tribus annis
2KGS|17|6|anno autem nono Osee cepit rex Assyriorum Samariam et transtulit Israhel in Assyrios posuitque eos in Ala et in Habor iuxta fluvium Gozan in civitatibus Medorum
2KGS|17|7|factum est enim cum peccassent filii Israhel Domino Deo suo qui eduxerat eos de terra Aegypti de manu Pharaonis regis Aegypti coluerunt deos alienos
2KGS|17|8|et ambulaverunt iuxta ritum gentium quas consumpserat Dominus in conspectu filiorum Israhel et regum Israhel quia similiter fecerant
2KGS|17|9|et operuerunt filii Israhel verbis non rectis Dominum Deum suum et aedificaverunt sibi excelsa in cunctis urbibus suis a turre custodum usque ad civitatem munitam
2KGS|17|10|feceruntque sibi statuas et lucos in omni colle sublimi et subter omne lignum nemorosum
2KGS|17|11|et adolebant ibi incensum super aras in more gentium quas transtulerat Dominus a facie eorum feceruntque verba pessima inritantes Dominum
2KGS|17|12|et coluerunt inmunditias de quibus praecepit Dominus eis ne facerent verbum hoc
2KGS|17|13|et testificatus est Dominus in Israhel et in Iuda per manum omnium prophetarum et videntum dicens revertimini a viis vestris pessimis et custodite praecepta mea et caerimonias iuxta omnem legem quam praecepi patribus vestris et sicut misi ad vos in manu servorum meorum prophetarum
2KGS|17|14|qui non audierunt sed induraverunt cervicem suam iuxta cervicem patrum suorum qui noluerunt oboedire Domino Deo suo
2KGS|17|15|et abiecerunt legitima eius et pactum quod pepigit cum patribus eorum et testificationes quibus contestatus est eos secutique sunt vanitates et vane egerunt et secuti sunt gentes quae erant per circuitum eorum super quibus praeceperat Dominus eis ut non facerent sicut et illae faciebant
2KGS|17|16|et dereliquerunt omnia praecepta Domini Dei sui feceruntque sibi conflatiles duos vitulos et lucos et adoraverunt universam militiam caeli servieruntque Baal
2KGS|17|17|et consecrabant ei filios suos et filias suas per ignem et divinationibus inserviebant et auguriis et tradiderunt se ut facerent malum coram Domino et inritarent eum
2KGS|17|18|iratusque est Dominus vehementer Israhel et abstulit eos de conspectu suo et non remansit nisi tribus Iuda tantummodo
2KGS|17|19|sed nec ipse Iuda custodivit mandata Domini Dei sui verum ambulavit in erroribus Israhel quos operatus fuerat
2KGS|17|20|proiecitque Dominus omne semen Israhel et adflixit eos et tradidit in manu diripientium donec proiceret eos a facie sua
2KGS|17|21|ex eo iam tempore quo scissus est Israhel a domo David et constituerunt sibi regem Hieroboam filium Nabath separavit enim Hieroboam Israhel a Domino et peccare eos fecit peccatum magnum
2KGS|17|22|et ambulaverunt filii Israhel in universis peccatis Hieroboam quae fecerat non recesserunt ab eis
2KGS|17|23|usquequo auferret Dominus Israhel a facie sua sicut locutus fuerat in manu omnium servorum suorum prophetarum translatusque est Israhel de terra sua in Assyrios usque in diem hanc
2KGS|17|24|adduxit autem rex Assyriorum de Babylone et de Chutha et de Haiath et de Emath et de Sepharvaim et conlocavit eos in civitatibus Samariae pro filiis Israhel qui possederunt Samariam et habitaverunt in urbibus eius
2KGS|17|25|cumque ibi habitare coepissent non timebant Dominum et inmisit eis Dominus leones qui interficiebant eos
2KGS|17|26|nuntiatumque est regi Assyriorum et dictum gentes quas transtulisti et habitare fecisti in civitatibus Samariae ignorant legitima Dei terrae et inmisit in eos Dominus leones et ecce interficiunt eos eo quod ignorent ritum Dei terrae
2KGS|17|27|praecepit autem rex Assyriorum dicens ducite illuc unum de sacerdotibus quos inde captivos adduxistis et vadat et habitet cum eis et doceat eos legitima Dei terrae
2KGS|17|28|igitur cum venisset unus de sacerdotibus his qui captivi ducti fuerant de Samaria habitavit in Bethel et docebat eos quomodo colerent Dominum
2KGS|17|29|et unaquaeque gens fabricata est deum suum posueruntque eos in fanis excelsis quae fecerant Samaritae gens et gens in urbibus suis in quibus habitabant
2KGS|17|30|viri enim babylonii fecerunt Socchothbenoth viri autem chutheni fecerunt Nergel et viri de Emath fecerunt Asima
2KGS|17|31|porro Evei fecerunt Nebaaz et Tharthac hii autem qui erant de Sepharvaim conburebant filios suos igni Adramelech et Anamelech diis Sepharvaim
2KGS|17|32|et nihilominus colebant Dominum fecerunt autem sibi de novissimis sacerdotes excelsorum et ponebant eos in fanis sublimibus
2KGS|17|33|et cum Dominum colerent diis quoque suis serviebant iuxta consuetudinem gentium de quibus translati fuerant Samariam
2KGS|17|34|usque in praesentem diem morem sequuntur antiquum non timent Dominum neque custodiunt caerimonias eius et iudicia et legem et mandatum quod praeceperat Dominus filiis Iacob quem cognominavit Israhel
2KGS|17|35|et percusserat cum eis pactum et mandaverat eis dicens nolite timere deos alienos et non adoretis eos neque colatis et non immoletis eis
2KGS|17|36|sed Dominum Deum vestrum qui eduxit vos de terra Aegypti in fortitudine magna et in brachio extento ipsum timete illum adorate et ipsi immolate
2KGS|17|37|caerimonias quoque et iudicia et legem et mandatum quod scripsit vobis custodite ut faciatis cunctis diebus et non timeatis deos alienos
2KGS|17|38|et pactum quod percussi vobiscum nolite oblivisci nec colatis deos alienos
2KGS|17|39|sed Dominum Deum vestrum timete et ipse eruet vos de manu omnium inimicorum vestrorum
2KGS|17|40|illi vero non audierunt sed iuxta consuetudinem suam pristinam perpetrabant
2KGS|17|41|fuerunt igitur gentes istae timentes quidem Dominum sed nihilominus et idolis suis servientes nam et filii eorum et nepotes sicut fecerunt parentes sui ita faciunt usque in praesentem diem
2KGS|18|1|anno tertio Osee filii Hela regis Israhel regnavit Ezechias filius Ahaz regis Iuda
2KGS|18|2|viginti quinque annorum erat cum regnare coepisset et viginti et novem annis regnavit in Hierusalem nomen matris eius Abi filia Zacchariae
2KGS|18|3|fecitque quod erat bonum coram Domino iuxta omnia quae fecerat David pater suus
2KGS|18|4|ipse dissipavit excelsa et contrivit statuas et succidit lucos confregitque serpentem aeneum quem fecerat Moses siquidem usque ad illud tempus filii Israhel adolebant ei incensum vocavitque eum Naasthan
2KGS|18|5|in Domino Deo Israhel speravit itaque post eum non fuit similis ei de cunctis regibus Iuda sed neque in his qui ante eum fuerunt
2KGS|18|6|et adhesit Domino et non recessit a vestigiis eius fecitque mandata eius quae praeceperat Dominus Mosi
2KGS|18|7|unde et erat Dominus cum eo et in cunctis ad quae procedebat sapienter se agebat rebellavit quoque contra regem Assyriorum et non servivit ei
2KGS|18|8|ipse percussit Philistheos usque Gazam et omnes terminos eorum a turre custodum usque ad civitatem muratam
2KGS|18|9|anno quarto regis Ezechiae qui erat annus septimus Osee filii Hela regis Israhel ascendit Salmanassar rex Assyriorum Samariam et obpugnavit eam
2KGS|18|10|et cepit nam post annos tres anno sexto Ezechiae id est nono anno Osee regis Israhel capta est Samaria
2KGS|18|11|et transtulit rex Assyriorum Israhel in Assyrios conlocavitque eos in Ala et in Habor fluviis Gozan in civitatibus Medorum
2KGS|18|12|quia non audierunt vocem Domini Dei sui sed praetergressi sunt pactum eius omnia quae praeceperat Moses servus Domini non audierunt neque fecerunt
2KGS|18|13|anno quartodecimo regis Ezechiae ascendit Sennacherib rex Assyriorum ad universas civitates Iuda munitas et cepit eas
2KGS|18|14|tunc misit Ezechias rex Iuda nuntios ad regem Assyriorum Lachis dicens peccavi recede a me et omne quod inposueris mihi feram indixit itaque rex Assyriorum Ezechiae regi Iudae trecenta talenta argenti et triginta talenta auri
2KGS|18|15|deditque Ezechias omne argentum quod reppertum fuerat in domo Domini et in thesauris regis
2KGS|18|16|in tempore illo confregit Ezechias valvas templi Domini et lamminas auri quas ipse adfixerat et dedit eas regi Assyriorum
2KGS|18|17|misit autem rex Assyriorum Tharthan et Rabsaris et Rabsacen de Lachis ad regem Ezechiam cum manu valida Hierusalem qui cum ascendissent venerunt in Hierusalem et steterunt iuxta aquaeductum piscinae superioris quae est in via agri Fullonis
2KGS|18|18|vocaveruntque regem egressus est autem ad eos Eliachim filius Helciae praepositus domus et Sobna scriba et Ioahe filius Asaph a commentariis
2KGS|18|19|dixitque ad eos Rabsaces loquimini Ezechiae haec dicit rex magnus rex Assyriorum quae est ista fiducia qua niteris
2KGS|18|20|forsitan inisti consilium ut praepares te ad proelium in quo confidis ut audeas rebellare
2KGS|18|21|an speras in baculo harundineo atque confracto Aegypto super quem si incubuerit homo comminutus ingreditur manum eius et perforabit eam sic est Pharao rex Aegypti omnibus qui confidunt in se
2KGS|18|22|quod si dixeritis mihi in Domino Deo nostro habemus fiduciam nonne iste est cuius abstulit Ezechias excelsa et altaria et praecepit Iudae et Hierusalem ante altare hoc adorabitis in Hierusalem
2KGS|18|23|nunc igitur transite ad dominum meum regem Assyriorum et dabo vobis duo milia equorum et videte an habere valeatis ascensores eorum
2KGS|18|24|et quomodo potestis resistere ante unum satrapam de servis domini mei minimis an fiduciam habes in Aegypto propter currus et equites
2KGS|18|25|numquid sine Domini voluntate ascendi ad locum istum ut demolirer eum Dominus dixit mihi ascende ad terram hanc et demolire eam
2KGS|18|26|dixerunt autem Eliachim filius Helciae et Sobna et Ioahe Rabsaci precamur ut loquaris nobis servis tuis syriace siquidem intellegimus hanc linguam et non loquaris nobis iudaice audiente populo qui est super murum
2KGS|18|27|responditque eis Rabsaces numquid ad dominum tuum et ad te misit me dominus meus ut loquerer sermones hos et non ad viros qui sedent super murum ut comedant stercora sua et bibant urinam suam vobiscum
2KGS|18|28|stetit itaque Rabsaces et clamavit voce magna iudaice et ait audite verba regis magni regis Assyriorum
2KGS|18|29|haec dicit rex non vos seducat Ezechias non enim poterit eruere vos de manu mea
2KGS|18|30|neque fiduciam vobis tribuat super Domino dicens eruens liberabit nos Dominus et non tradetur civitas haec in manu regis Assyriorum
2KGS|18|31|nolite audire Ezechiam haec enim dicit rex Assyriorum facite mecum quod vobis est utile et egredimini ad me et comedet unusquisque de vinea sua et de ficu sua et bibetis aquas de cisternis vestris
2KGS|18|32|donec veniam et transferam vos in terram quae similis terrae vestrae est in terram fructiferam et fertilem vini terram panis et vinearum terram olivarum et olei ac mellis et vivetis et non moriemini nolite audire Ezechiam qui vos decipit dicens Dominus liberabit nos
2KGS|18|33|numquid liberaverunt dii gentium terram suam de manu regis Assyriorum
2KGS|18|34|ubi est deus Emath et Arfad ubi est deus Sepharvaim Ana et Ava numquid liberaverunt Samariam de manu mea
2KGS|18|35|quinam illi sunt in universis diis terrarum qui eruerunt regionem suam de manu mea ut possit eruere Dominus Hierusalem de manu mea
2KGS|18|36|tacuit itaque populus et non respondit ei quicquam siquidem praeceptum regis acceperant ut non responderent ei
2KGS|18|37|venitque Eliachim filius Helciae praepositus domus et Sobna scriba et Ioahe filius Asaph a commentariis ad Ezechiam scissis vestibus et nuntiaverunt ei verba Rabsacis
2KGS|19|1|quae cum audisset rex Ezechias scidit vestimenta sua et opertus est sacco ingressusque est domum Domini
2KGS|19|2|et misit Eliachim praepositum domus et Sobnam scribam et senes de sacerdotibus opertos saccis ad Esaiam prophetam filium Amos
2KGS|19|3|qui dixerunt haec dicit Ezechias dies tribulationis et increpationis et blasphemiae dies iste venerunt filii usque ad partum et vires non habet parturiens
2KGS|19|4|si forte audiat Dominus Deus tuus universa verba Rabsacis quem misit rex Assyriorum dominus suus ut exprobraret Deum viventem et argueret verbis quae audivit Dominus Deus tuus et fac orationem pro reliquiis quae reppertae sunt
2KGS|19|5|venerunt ergo servi regis Ezechiae ad Esaiam
2KGS|19|6|dixitque eis Esaias haec dicetis domino vestro haec dicit Dominus noli timere a facie sermonum quos audisti quibus blasphemaverunt pueri regis Assyriorum me
2KGS|19|7|ecce ego inmittam ei spiritum et audiet nuntium et revertetur in terram suam et deiciam eum gladio in terra sua
2KGS|19|8|reversus est igitur Rabsaces et invenit regem Assyriorum expugnantem Lobnam audierat enim quod recessisset de Lachis
2KGS|19|9|cumque audisset de Tharaca rege Aethiopiae dicentes ecce egressus est ut pugnet adversum te et iret contra eum misit nuntios ad Ezechiam dicens
2KGS|19|10|haec dicite Ezechiae regi Iudae non te seducat Deus tuus in quo habes fiduciam neque dicas non tradetur Hierusalem in manu regis Assyriorum
2KGS|19|11|tu enim ipse audisti quae fecerint reges Assyriorum universis terris quomodo vastaverint eas num ergo solus poteris liberari
2KGS|19|12|numquid liberaverunt dii gentium singulos quos vastaverunt patres mei Gozan videlicet et Aran et Reseph et filios Eden qui erant in Thelassar
2KGS|19|13|ubi est rex Emath et rex Arfad et rex civitatis Sepharvaim Ana et Ava
2KGS|19|14|itaque cum accepisset Ezechias litteras de manu nuntiorum et legisset eas ascendit in domum Domini et expandit eas coram Domino
2KGS|19|15|et oravit in conspectu eius dicens Domine Deus Israhel qui sedes super cherubin tu es Deus solus regum omnium terrae tu fecisti caelum et terram
2KGS|19|16|inclina aurem tuam et audi aperi Domine oculos tuos et vide et audi omnia verba Sennacherib qui misit ut exprobraret nobis Deum viventem
2KGS|19|17|vere Domine dissipaverunt reges Assyriorum gentes et terras omnium
2KGS|19|18|et miserunt deos eorum in ignem non enim erant dii sed opera manuum hominum e ligno et lapide et perdiderunt eos
2KGS|19|19|nunc igitur Domine Deus noster salvos nos fac de manu eius ut sciant omnia regna terrae quia tu es Dominus Deus solus
2KGS|19|20|misit autem Esaias filius Amos ad Ezechiam dicens haec dicit Dominus Deus Israhel quae deprecatus es me super Sennacherib rege Assyriorum audivi
2KGS|19|21|iste est sermo quem locutus est Dominus de eo sprevit te et subsannavit virgo filia Sion post tergum tuum caput movit filia Hierusalem
2KGS|19|22|cui exprobrasti et quem blasphemasti contra quem exaltasti vocem et elevasti in excelsum oculos tuos contra Sanctum Israhel
2KGS|19|23|per manum servorum tuorum exprobrasti Domino et dixisti in multitudine curruum meorum ascendi excelsa montium in summitate Libani et succidi sublimes cedros eius electas abietes eius et ingressus sum usque ad terminos eius saltum Carmeli eius
2KGS|19|24|ego succidi et bibi aquas alienas et siccavi vestigiis pedum meorum omnes aquas clausas
2KGS|19|25|numquid non audisti quid ab initio fecerim ex diebus antiquis plasmavi illud et nunc adduxi eruntque in ruinam collium pugnantium civitates munitae
2KGS|19|26|et qui sedent in eis humiles manu contremuerunt et confusi sunt facti sunt quasi faenum agri et virens herba tectorum quae arefacta est antequam veniret ad maturitatem
2KGS|19|27|habitaculum tuum et egressum tuum et viam tuam ego praescivi et furorem tuum contra me
2KGS|19|28|insanisti in me et superbia tua ascendit in aures meas ponam itaque circulum in naribus tuis et camum in labris tuis et reducam te in viam per quam venisti
2KGS|19|29|tibi autem Ezechia hoc erit signum comede hoc anno quod reppereris in secundo autem anno quae sponte nascuntur porro in anno tertio seminate et metite plantate vineas et comedite fructum earum
2KGS|19|30|et quodcumque reliquum fuerit de domo Iuda mittet radicem deorsum et faciet fructum sursum
2KGS|19|31|de Hierusalem quippe egredientur reliquiae et quod salvetur de monte Sion zelus Domini exercituum faciet hoc
2KGS|19|32|quam ob rem haec dicit Dominus de rege Assyriorum non ingredietur urbem hanc nec mittet in eam sagittam nec occupabit eam clypeus nec circumdabit eam munitio
2KGS|19|33|per viam qua venit revertetur et civitatem hanc non ingredietur dicit Dominus
2KGS|19|34|protegamque urbem hanc et salvabo eam propter me et propter David servum meum
2KGS|19|35|factum est igitur in nocte illa venit angelus Domini et percussit castra Assyriorum centum octoginta quinque milia cumque diluculo surrexisset vidit omnia corpora mortuorum et recedens abiit
2KGS|19|36|et reversus est Sennacherib rex Assyriorum et mansit in Nineve
2KGS|19|37|cumque adoraret in templo Neserach deum suum Adramelech et Sarasar filii eius percusserunt eum gladio fugeruntque in terram Armeniorum et regnavit Eseraddon filius eius pro eo
2KGS|20|1|in diebus illis aegrotavit Ezechias usque ad mortem et venit ad eum Esaias filius Amos prophetes dixitque ei haec dicit Dominus Deus praecipe domui tuae morieris enim et non vives
2KGS|20|2|qui convertit faciem suam ad parietem et oravit Dominum dicens
2KGS|20|3|obsecro Domine memento quomodo ambulaverim coram te in veritate et in corde perfecto et quod placitum est coram te fecerim flevit itaque Ezechias fletu magno
2KGS|20|4|et antequam egrederetur Esaias mediam partem atrii factus est sermo Domini ad eum dicens
2KGS|20|5|revertere et dic Ezechiae duci populi mei haec dicit Dominus Deus David patris tui audivi orationem tuam vidi lacrimam tuam et ecce sanavi te die tertio ascendes templum Domini
2KGS|20|6|et addam diebus tuis quindecim annos sed et de manu regis Assyriorum liberabo te et civitatem hanc et protegam urbem istam propter me et propter David servum meum
2KGS|20|7|dixitque Esaias adferte massam ficorum quam cum adtulissent et posuissent super ulcus eius curatus est
2KGS|20|8|dixerat autem Ezechias ad Esaiam quod erit signum quia Dominus me sanabit et quia ascensurus sum die tertio templum Domini
2KGS|20|9|cui ait Esaias hoc erit signum a Domino quod facturus sit Dominus sermonem quem locutus est vis ut accedat umbra decem lineis an ut revertatur totidem gradibus
2KGS|20|10|et ait Ezechias facile est umbram crescere decem lineis nec hoc volo ut fiat sed ut revertatur retrorsum decem gradibus
2KGS|20|11|invocavit itaque Esaias propheta Dominum et reduxit umbram per lineas quibus iam descenderat in horologio Ahaz retrorsum decem gradibus
2KGS|20|12|in tempore illo misit Berodach Baladan filius Baladan rex Babyloniorum litteras et munera ad Ezechiam audierat enim quod aegrotasset Ezechias
2KGS|20|13|laetatus est autem in adventum eorum Ezechias et ostendit eis domum aromatum et aurum et argentum et pigmenta varia unguenta quoque et domum vasorum suorum et omnia quae habere potuerat in thesauris suis non fuit quod non monstraret eis Ezechias in domo sua et in omni potestate sua
2KGS|20|14|venit autem Esaias propheta ad regem Ezechiam dixitque ei quid dixerunt viri isti aut unde venerunt ad te cui ait Ezechias de terra longinqua venerunt de Babylone
2KGS|20|15|at ille respondit quid viderunt in domo tua ait Ezechias omnia quae sunt in domo mea viderunt nihil est quod non monstraverim eis in thesauris meis
2KGS|20|16|dixit itaque Esaias Ezechiae audi sermonem Domini
2KGS|20|17|ecce dies venient et auferentur omnia quae sunt in domo tua et quae condiderunt patres tui usque in diem hanc in Babylone non remanebit quicquam ait Dominus
2KGS|20|18|sed et de filiis tuis qui egredientur ex te quos generabis tollentur et erunt eunuchi in palatio regis Babylonis
2KGS|20|19|dixit Ezechias ad Esaiam bonus sermo Domini quem locutus est sit pax et veritas in diebus meis
2KGS|20|20|reliqua autem sermonum Ezechiae et omnis fortitudo eius et quomodo fecerit piscinam et aquaeductum et introduxerit aquas in civitatem nonne haec scripta sunt in libro sermonum dierum regum Iuda
2KGS|20|21|dormivitque Ezechias cum patribus suis et regnavit Manasses filius eius pro eo
2KGS|21|1|duodecim annorum erat Manasses cum regnare coepisset et quinquaginta quinque annis regnavit in Hierusalem nomen matris eius Aphsiba
2KGS|21|2|fecitque malum in conspectu Domini iuxta idola gentium quas delevit Dominus a facie filiorum Israhel
2KGS|21|3|conversusque est et aedificavit excelsa quae dissipaverat Ezechias pater eius et erexit aras Baal et fecit lucos sicut fecerat Ahab rex Israhel et adoravit omnem militiam caeli et coluit eam
2KGS|21|4|extruxitque aras in domo Domini de qua dixit Dominus in Hierusalem ponam nomen meum
2KGS|21|5|et extruxit altaria universae militiae caeli in duobus atriis templi Domini
2KGS|21|6|et transduxit filium suum per ignem et ariolatus est et observavit auguria et fecit pythones et aruspices multiplicavit ut faceret malum coram Domino et inritaret eum
2KGS|21|7|posuit quoque idolum luci quem fecerat in templo Domini super quo locutus est Dominus ad David et ad Salomonem filium eius in templo hoc et in Hierusalem quam elegi de cunctis tribubus Israhel ponam nomen meum in sempiternum
2KGS|21|8|et ultra non faciam commoveri pedem Israhel de terra quam dedi patribus eorum sic tamen si custodierint opere omnia quae praecepi eis et universam legem quam mandavit eis servus meus Moses
2KGS|21|9|illi vero non audierunt sed seducti sunt a Manasse ut facerent malum super gentes quas contrivit Dominus a facie filiorum Israhel
2KGS|21|10|locutusque est Dominus in manu servorum suorum prophetarum dicens
2KGS|21|11|quia fecit Manasses rex Iuda abominationes istas pessimas super omnia quae fecerunt Amorrei ante eum et peccare fecit etiam Iudam in inmunditiis suis
2KGS|21|12|propterea haec dicit Dominus Deus Israhel ecce ego inducam mala super Hierusalem et Iudam ut quicumque audierit tinniant ambae aures eius
2KGS|21|13|et extendam super Hierusalem funiculum Samariae et pondus domus Ahab et delebo Hierusalem sicut deleri solent tabulae delens vertam et ducam crebrius stilum super faciem eius
2KGS|21|14|dimittam vero reliquias hereditatis meae et tradam eas in manu inimicorum eius eruntque in vastitate et rapina cunctis adversariis suis
2KGS|21|15|eo quod fecerint malum coram me et perseveraverint inritantes me ex die qua egressi sunt patres eorum ex Aegypto usque ad diem hanc
2KGS|21|16|insuper et sanguinem innoxium fudit Manasses multum nimis donec impleret Hierusalem usque ad os absque peccatis suis quibus peccare fecit Iudam ut faceret malum coram Domino
2KGS|21|17|reliqua autem sermonum Manasse et universa quae fecit et peccatum eius quod peccavit nonne haec scripta sunt in libro sermonum dierum regum Iuda
2KGS|21|18|dormivitque Manasses cum patribus suis et sepultus est in horto domus suae in horto Aza et regnavit Amon filius eius pro eo
2KGS|21|19|viginti et duo annorum erat Amon cum regnare coepisset duobusque annis regnavit in Hierusalem nomen matris eius Mesallemeth filia Arus de Iethba
2KGS|21|20|fecitque malum in conspectu Domini sicut fecerat Manasses pater eius
2KGS|21|21|et ambulavit in omni via per quam ambulaverat pater eius servivitque inmunditiis quibus servierat pater suus et adoravit eas
2KGS|21|22|et dereliquit Dominum Deum patrum suorum et non ambulavit in via Domini
2KGS|21|23|tetenderuntque ei insidias servi sui et interfecerunt regem in domo sua
2KGS|21|24|percussit autem populus terrae omnes qui coniuraverant contra regem Amon et constituerunt sibi regem Iosiam filium eius pro eo
2KGS|21|25|reliqua autem sermonum Amon quae fecit nonne haec scripta sunt in libro sermonum dierum regum Iuda
2KGS|21|26|sepelieruntque eum in sepulchro suo in horto Aza et regnavit Iosias filius eius pro eo
2KGS|22|1|octo annorum erat Iosias cum regnare coepisset et triginta uno anno regnavit in Hierusalem nomen matris eius Idida filia Phadaia de Besecath
2KGS|22|2|fecitque quod placitum erat coram Domino et ambulavit per omnes vias David patris sui non declinavit ad dextram sive ad sinistram
2KGS|22|3|anno autem octavodecimo regis Iosiae misit rex Saphan filium Aslia filii Mesullam scribam templi Domini dicens ei
2KGS|22|4|vade ad Helciam sacerdotem magnum ut confletur pecunia quae inlata est in templum Domini quam collegerunt ianitores a populo
2KGS|22|5|deturque fabris per praepositos in domo Domini qui et distribuent eam his qui operantur in templo Domini ad instauranda sarta tecta templi
2KGS|22|6|tignariis videlicet et cementariis et his qui interrupta conponunt et ut emantur ligna et lapides de lapidicinis ad instaurandum templum
2KGS|22|7|verumtamen non supputetur eis argentum quod accipiunt sed in potestate habeant et in fide
2KGS|22|8|dixit autem Helcias pontifex ad Saphan scribam librum legis repperi in domo Domini deditque Helcias volumen Saphan qui et legit illud
2KGS|22|9|venit quoque Saphan scriba ad regem et renuntiavit ei quod praeceperat et ait conflaverunt servi tui pecuniam quae repperta est in domo Domini et dederunt ut distribueretur fabris a praefectis operum templi Domini
2KGS|22|10|narravitque Saphan scriba regi dicens librum dedit mihi Helcias sacerdos quem cum legisset Saphan coram rege
2KGS|22|11|et audisset rex verba libri legis Domini scidit vestimenta sua
2KGS|22|12|et praecepit Helciae sacerdoti et Ahicham filio Saphan et Achobor filio Micha et Saphan scribae et Asaiae servo regis dicens
2KGS|22|13|ite et consulite Dominum super me et super populo et super omni Iuda de verbis voluminis istius quod inventum est magna enim ira Domini succensa est contra nos quia non audierunt patres nostri verba libri huius ut facerent omne quod scriptum est nobis
2KGS|22|14|ierunt itaque Helcias sacerdos et Ahicham et Achobor et Saphan et Asaia ad Oldam propheten uxorem Sellum filii Thecue filii Araas custodis vestium quae habitabat in Hierusalem in secunda locutique sunt ad eam
2KGS|22|15|et illa respondit eis haec dicit Dominus Deus Israhel dicite viro qui misit vos ad me
2KGS|22|16|haec dicit Dominus ecce ego adducam mala super locum hunc et super habitatores eius omnia verba legis quae legit rex Iuda
2KGS|22|17|quia dereliquerunt me et sacrificaverunt diis alienis inritantes me in cunctis operibus manuum suarum et succendetur indignatio mea in loco hoc et non extinguetur
2KGS|22|18|regi autem Iuda qui misit vos ut consuleretis Dominum sic dicetis haec dicit Dominus Deus Israhel pro eo quod audisti verba voluminis
2KGS|22|19|et perterritum est cor tuum et humiliatus es coram Domino auditis sermonibus contra locum istum et habitatores eius quo videlicet fierent in stuporem et in maledictum et scidisti vestimenta tua et flevisti coram me et ego audivi ait Dominus
2KGS|22|20|idcirco colligam te ad patres tuos et colligeris ad sepulchrum tuum in pace ut non videant oculi tui omnia mala quae inducturus sum super locum istum
2KGS|23|1|et renuntiaverunt regi quod dixerat qui misit et congregati sunt ad eum omnes senes Iuda et Hierusalem
2KGS|23|2|ascenditque rex templum Domini et omnes viri Iuda universique qui habitant in Hierusalem cum eo sacerdotes et prophetae et omnis populus a parvo usque ad magnum legitque cunctis audientibus omnia verba libri foederis qui inventus est in domo Domini
2KGS|23|3|stetitque rex super gradum et percussit foedus coram Domino ut ambularent post Dominum et custodirent praecepta eius et testimonia et caerimonias in omni corde et in tota anima et suscitarent verba foederis huius quae scripta erant in libro illo adquievitque populus pacto
2KGS|23|4|et praecepit rex Helciae pontifici et sacerdotibus secundi ordinis et ianitoribus ut proicerent de templo Domini omnia vasa quae facta fuerant Baal et in luco et universae militiae caeli et conbusit ea foris Hierusalem in convalle Cedron et tulit pulverem eorum in Bethel
2KGS|23|5|et delevit aruspices quos posuerant reges Iuda ad sacrificandum in excelsis per civitates Iuda et in circuitu Hierusalem et eos qui adolebant incensum Baal et soli et lunae et duodecim signis et omni militiae caeli
2KGS|23|6|et efferri fecit lucum de domo Domini foras Hierusalem in convalle Cedron et conbusit eum ibi et redegit in pulverem et proiecit super sepulchrum vulgi
2KGS|23|7|destruxit quoque aediculas effeminatorum quae erant in domo Domini pro quibus mulieres texebant quasi domunculas luci
2KGS|23|8|congregavitque omnes sacerdotes de civitatibus Iuda et contaminavit excelsa ubi sacrificabant sacerdotes de Gabaa usque Bersabee et destruxit aras portarum in introitu ostii Iosue principis civitatis quod erat ad sinistram portae civitatis
2KGS|23|9|verumtamen non ascendebant sacerdotes excelsorum ad altare Domini in Hierusalem sed tantum comedebant azyma in medio fratrum suorum
2KGS|23|10|contaminavit quoque Thafeth quod est in convalle filii Ennom ut nemo consecraret filium suum aut filiam per ignem Moloch
2KGS|23|11|abstulit quoque equos quos dederant reges Iudae soli in introitu templi Domini iuxta exedram Nathanmelech eunuchi qui erat in Farurim currus autem solis conbusit igni
2KGS|23|12|altaria quoque quae erant super tecta cenaculi Ahaz quae fecerant reges Iuda et altaria quae fecerat Manasses in duobus atriis templi Domini destruxit rex et cucurrit inde et dispersit cinerem eorum in torrentem Cedron
2KGS|23|13|excelsa quoque quae erant in Hierusalem ad dexteram partem montis Offensionis quae aedificaverat Salomon rex Israhel Astharoth idolo Sidoniorum et Chamos offensioni Moab et Melchom abominationi filiorum Ammon polluit rex
2KGS|23|14|et contrivit statuas et succidit lucos replevitque loca eorum ossibus mortuorum
2KGS|23|15|insuper et altare quod erat in Bethel excelsum quod fecerat Hieroboam filius Nabath qui peccare fecit Israhel et altare illud et excelsum destruxit atque conbusit et comminuit in pulverem succenditque etiam lucum
2KGS|23|16|et conversus Iosias vidit ibi sepulchra quae erant in monte misitque et tulit ossa de sepulchris et conbusit ea super altare et polluit illud iuxta verbum Domini quod locutus est vir Dei qui praedixerat verba haec
2KGS|23|17|et ait quis est titulus ille quem video responderuntque ei cives illius urbis sepulchrum est hominis Dei qui venit de Iuda et praedixit verba haec quae fecisti super altare Bethel
2KGS|23|18|et ait dimittite eum nemo commoveat ossa eius et intacta manserunt ossa illius cum ossibus prophetae qui venerat de Samaria
2KGS|23|19|insuper et omnia fana excelsorum quae erant in civitatibus Samariae quae fecerant reges Israhel ad inritandum Dominum abstulit Iosias et fecit eis secundum omnia opera quae fecerat in Bethel
2KGS|23|20|et occidit universos sacerdotes excelsorum qui erant ibi super altaria et conbusit ossa humana super ea reversusque est Hierusalem
2KGS|23|21|et praecepit omni populo dicens facite phase Domino Deo vestro secundum quod scriptum est in libro foederis huius
2KGS|23|22|nec enim factum est phase tale a diebus iudicum qui iudicaverunt Israhel et omnium dierum regum Israhel et regum Iuda
2KGS|23|23|sicut in octavodecimo anno regis Iosiae factum est phase istud Domino in Hierusalem
2KGS|23|24|sed et pythones et ariolos et figuras idolorum et inmunditias abominationesque quae fuerant in terra Iuda et in Hierusalem abstulit Iosias ut statueret verba legis quae scripta sunt in libro quem invenit Helcias sacerdos in templo Domini
2KGS|23|25|similis illi non fuit ante eum rex qui reverteretur ad Dominum in omni corde suo et in tota anima sua et in universa virtute sua iuxta omnem legem Mosi neque post eum surrexit similis illi
2KGS|23|26|verumtamen non est aversus Dominus ab ira furoris sui magni quo iratus est furor eius contra Iudam propter inritationes quibus provocaverat eum Manasses
2KGS|23|27|dixit itaque Dominus etiam Iudam auferam a facie mea sicut abstuli Israhel et proiciam civitatem hanc quam elegi Hierusalem et domum de qua dixi erit nomen meum ibi
2KGS|23|28|reliqua autem verba Iosiae et universa quae fecit nonne haec scripta sunt in libro verborum dierum regum Iuda
2KGS|23|29|in diebus eius ascendit Pharao Necho rex Aegypti contra regem Assyriorum ad flumen Eufraten et abiit Iosias rex in occursum eius et occisus est in Mageddo cum vidisset eum
2KGS|23|30|et portaverunt eum servi sui mortuum de Mageddo et pertulerunt in Hierusalem et sepelierunt eum in sepulchro suo tulitque populus terrae Ioahaz filium Iosiae et unxerunt eum et constituerunt eum regem pro patre suo
2KGS|23|31|viginti trium annorum erat Ioahaz cum regnare coepisset et tribus mensibus regnavit in Hierusalem nomen matris eius Amithal filia Hieremiae de Lobna
2KGS|23|32|et fecit malum coram Domino iuxta omnia quae fecerant patres eius
2KGS|23|33|vinxitque eum Pharao Necho in Rebla quae est in terra Emath ne regnaret in Hierusalem et inposuit multam terrae centum talentis argenti et talento auri
2KGS|23|34|regemque constituit Pharao Necho Eliachim filium Iosiae pro Iosia patre eius vertitque nomen eius Ioiachim porro Ioahaz tulit et duxit in Aegyptum
2KGS|23|35|argentum autem et aurum dedit Ioiachim Pharaoni cum indixisset terrae per singulos ut conferretur iuxta praeceptum Pharaonis et unumquemque secundum vires suas exegit tam argentum quam aurum de populo terrae ut daret Pharaoni Necho
2KGS|23|36|viginti quinque annorum erat Ioiachim cum regnare coepisset et undecim annis regnavit in Hierusalem nomen matris eius Zebida filia Phadaia de Ruma
2KGS|23|37|et fecit malum coram Domino iuxta omnia quae fecerant patres eius
2KGS|24|1|in diebus eius ascendit Nabuchodonosor rex Babylonis et factus est ei Ioiachim servus tribus annis et rursum rebellavit contra eum
2KGS|24|2|inmisitque ei Dominus latrunculos Chaldeorum et latrunculos Syriae latrunculos Moab et latrunculos filiorum Ammon et inmisit eos in Iudam ut disperderent eum iuxta verbum Domini quod locutus erat per servos suos prophetas
2KGS|24|3|factum est autem hoc per verbum Domini contra Iudam ut auferret eum coram se propter peccata Manasse universa quae fecit
2KGS|24|4|et propter sanguinem innoxium quem effudit et implevit Hierusalem cruore innocentium et ob hanc rem noluit Dominus propitiari
2KGS|24|5|reliqua autem sermonum Ioiachim et universa quae fecit nonne haec scripta sunt in libro sermonum dierum regum Iuda et dormivit Ioiachim cum patribus suis
2KGS|24|6|regnavitque Ioiachin filius eius pro eo
2KGS|24|7|et ultra non addidit rex Aegypti ut egrederetur de terra sua tulerat enim rex Babylonis a rivo Aegypti usque ad fluvium Eufraten omnia quae fuerant regis Aegypti
2KGS|24|8|decem et octo annorum erat Ioiachin cum regnare coepisset et tribus mensibus regnavit in Hierusalem nomen matris eius Naestha filia Helnathan de Hierusalem
2KGS|24|9|et fecit malum coram Domino iuxta omnia quae fecerat pater eius
2KGS|24|10|in tempore illo ascenderunt servi Nabuchodonosor regis Babylonis in Hierusalem et circumdata est urbs munitionibus
2KGS|24|11|venitque Nabuchodonosor rex Babylonis ad civitatem cum servi eius obpugnarent eam
2KGS|24|12|egressusque est Ioiachin rex Iuda ad regem Babylonis ipse et mater eius et servi eius et principes eius et eunuchi eius et suscepit eum rex Babylonis anno octavo regni sui
2KGS|24|13|et protulit inde omnes thesauros domus Domini et thesauros domus regiae et concidit universa vasa aurea quae fecerat Salomon rex Israhel in templo Domini iuxta verbum Domini
2KGS|24|14|et transtulit omnem Hierusalem et universos principes et omnes fortes exercitus decem milia in captivitatem et omnem artificem et clusorem nihilque relictum est exceptis pauperibus populi terrae
2KGS|24|15|transtulit quoque Ioiachin in Babylonem et matrem regis et uxores regis et eunuchos eius et iudices terrae duxit in captivitatem de Hierusalem in Babylonem
2KGS|24|16|et omnes viros robustos septem milia et artifices et clusores mille omnes viros fortes et bellatores duxitque eos rex Babylonis captivos in Babylonem
2KGS|24|17|et constituit Matthaniam patruum eius pro eo inposuitque nomen ei Sedeciam
2KGS|24|18|vicesimum et primum annum aetatis habebat Sedecias cum regnare coepisset et undecim annis regnavit in Hierusalem nomen matris eius erat Amithal filia Hieremiae de Lobna
2KGS|24|19|et fecit malum coram Domino iuxta omnia quae fecerat Ioiachim
2KGS|24|20|irascebatur enim Dominus contra Hierusalem et contra Iudam donec proiceret eos a facie sua recessitque Sedecias a rege Babylonis
2KGS|25|1|factum est autem anno nono regni eius mense decimo decima die mensis venit Nabuchodonosor rex Babylonis ipse et omnis exercitus eius in Hierusalem et circumdederunt eam et extruxerunt in circuitu eius munitiones
2KGS|25|2|et clausa est civitas atque vallata usque ad undecimum annum regis Sedeciae
2KGS|25|3|nona die mensis praevaluitque fames in civitate nec erat panis populo terrae
2KGS|25|4|et interrupta est civitas et omnes viri bellatores nocte fugerunt per viam portae quae est inter duplicem murum ad hortum regis porro Chaldei obsidebant in circuitu civitatem fugit itaque per viam quae ducit ad campestria solitudinis
2KGS|25|5|et persecutus est exercitus Chaldeorum regem conprehenditque eum in planitie Hiericho et omnes bellatores qui erant cum eo dispersi sunt et reliquerunt eum
2KGS|25|6|adprehensum ergo regem duxerunt ad regem Babylonis in Reblatha qui locutus est cum eo iudicium
2KGS|25|7|filios autem Sedeciae occidit coram eo et oculos eius effodit vinxitque eum catenis et adduxit in Babylonem
2KGS|25|8|mense quinto septima die mensis ipse est annus nonusdecimus regis Babylonis venit Nabuzardan princeps exercitus servus regis Babylonis Hierusalem
2KGS|25|9|et succendit domum Domini et domum regis et domos Hierusalem omnemque domum conbusit igni
2KGS|25|10|et muros Hierusalem in circuitu destruxit omnis exercitus Chaldeorum qui erat cum principe militum
2KGS|25|11|reliquam autem populi partem qui remanserat in civitate et perfugas qui transfugerant ad regem Babylonis et reliquum vulgus transtulit Nabuzardan princeps militiae
2KGS|25|12|et de pauperibus terrae reliquit vinitores et agricolas
2KGS|25|13|columnas autem aereas quae erant in templo Domini et bases et mare aereum quod erat in domo Domini confregerunt Chaldei et transtulerunt aes omnium in Babylonem
2KGS|25|14|ollas quoque aereas et trullas et tridentes et scyphos et omnia vasa aerea in quibus ministrabant tulerunt
2KGS|25|15|necnon turibula et fialas quae aurea aurea et quae argentea argentea tulit princeps militiae
2KGS|25|16|id est columnas duas mare unum et bases quas fecerat Salomon in templo Domini non erat pondus aeris omnium vasorum
2KGS|25|17|decem et octo cubitos altitudinis habebat columna una et capitellum aereum super se altitudinis trium cubitorum et reticulum et malogranata super capitellum columnae omnia aerea similem et columna secunda habebat ornatum
2KGS|25|18|tulit quoque princeps militiae Seraian sacerdotem primum et Sophoniam sacerdotem secundum et tres ianitores
2KGS|25|19|et de civitate eunuchum unum qui erat praefectus super viros bellatores et quinque viros de his qui steterant coram rege quos repperit in civitate et Sopher principem exercitus qui probabat tirones de populo terrae et sex viros e vulgo qui inventi fuerant in civitate
2KGS|25|20|quos tollens Nabuzardan princeps militum duxit ad regem Babylonis in Reblatha
2KGS|25|21|percussitque eos rex Babylonis et interfecit in Reblatha in terra Emath et translatus est Iuda de terra sua
2KGS|25|22|populo autem qui relictus erat in terra Iuda quem dimiserat Nabuchodonosor rex Babylonis praefecit Godoliam filium Ahicham filii Saphan
2KGS|25|23|quod cum audissent omnes duces militum ipsi et viri qui erant cum eis videlicet quod constituisset rex Babylonis Godoliam venerunt ad Godoliam in Maspha Ismahel filius Nathaniae et Iohanan filius Caree et Sareia filius Thenaameth Nethophathites et Iezonias filius Maachathi ipsi et socii eorum
2KGS|25|24|iuravitque eis Godolias et sociis eorum dicens nolite timere servire Chaldeis manete in terra et servite regi Babylonis et bene erit vobis
2KGS|25|25|factum est autem in mense septimo venit Ismahel filius Nathaniae filii Elisama de semine regio et decem viri cum eo percusseruntque Godoliam qui mortuus est sed et Iudaeos et Chaldeos qui erant cum eo in Maspha
2KGS|25|26|consurgens autem omnis populus a parvo usque ad magnum et principes militum venerunt in Aegyptum timentes Chaldeos
2KGS|25|27|factum est vero anno tricesimo septimo transmigrationis Ioiachin regis Iudae mense duodecimo vicesima septima die mensis sublevavit Evilmerodach rex Babylonis anno quo regnare coeperat caput Ioiachin regis Iuda de carcere
2KGS|25|28|et locutus est ei benigna et posuit thronum eius super thronum regum qui erant cum eo in Babylone
2KGS|25|29|et mutavit vestes eius quas habuerat in carcere et comedebat panem semper in conspectu eius cunctis diebus vitae suae
2KGS|25|30|annonam quoque constituit ei absque intermissione quae et dabatur ei a rege per singulos dies omnibus diebus vitae suae
1CHR|1|1|Adam Seth Enos
1CHR|1|2|Cainan Malelehel Iared
1CHR|1|3|Enoch Matusale Lamech
1CHR|1|4|Noe Sem Ham et Iafeth
1CHR|1|5|filii Iafeth Gomer Magog Madai et Iavan Thubal Mosoch Thiras
1CHR|1|6|porro filii Gomer Aschenez et Rifath et Thogorma
1CHR|1|7|filii autem Iavan Elisa et Tharsis Cetthim et Dodanim
1CHR|1|8|filii Ham Chus et Mesraim Phut et Chanaan
1CHR|1|9|filii autem Chus Saba et Evila Sabatha et Rechma et Sabathaca porro filii Rechma Saba et Dadan
1CHR|1|10|Chus autem genuit Nemrod iste coepit esse potens in terra
1CHR|1|11|Mesraim vero genuit Ludim et Anamim et Laabim et Nepthuim
1CHR|1|12|Phethrosim quoque et Chasluim de quibus egressi sunt Philisthim et Capthurim
1CHR|1|13|Chanaan vero genuit Sidonem primogenitum et Heth
1CHR|1|14|Iebuseum quoque et Amorreum et Gergeseum
1CHR|1|15|Evheumque et Aruceum et Asineum
1CHR|1|16|Aradium quoque et Samareum et Ematheum
1CHR|1|17|filii Sem Aelam et Assur et Arfaxad et Lud et Aram et Us et Hul et Gothor et Mosoch
1CHR|1|18|Arfaxad autem genuit Sala qui et ipse genuit Heber
1CHR|1|19|porro Heber nati sunt duo filii nomen uni Phaleg quia in diebus eius divisa est terra et nomen fratris eius Iectan
1CHR|1|20|Iectan autem genuit Helmodad et Saleph et Asermoth et Iare
1CHR|1|21|Aduram quoque et Uzal et Decla
1CHR|1|22|Ebal etiam et Abimahel et Saba necnon
1CHR|1|23|et Ophir et Evila et Iobab omnes isti filii Iectan
1CHR|1|24|Sem Arfaxad Sale
1CHR|1|25|Heber Phaleg Raau
1CHR|1|26|Serug Nahor Thare
1CHR|1|27|Abram iste est Abraham
1CHR|1|28|filii autem Abraham Isaac et Ismahel
1CHR|1|29|et hae generationes eorum primogenitus Ismahelis Nabaioth et Cedar et Adbeel et Mabsam
1CHR|1|30|Masma et Duma Massa Adad et Thema
1CHR|1|31|Iathur Naphis Cedma hii sunt filii Ismahelis
1CHR|1|32|filii autem Cetthurae concubinae Abraham quos genuit Zamram Iecsan Madan Madian Iesboc Sue porro filii Iecsan Saba et Dadan
1CHR|1|33|filii autem Madian Epha et Apher et Enoch et Abida et Eldaa omnes hii filii Cetthurae
1CHR|1|34|generavit autem Abraham Isaac cuius fuerunt filii Esau et Israhel
1CHR|1|35|filii Esau Eliphaz Rauhel Iaus Ialam Core
1CHR|1|36|filii Eliphaz Theman Omer Sepphu Gethem Cenez Thamna Amalech
1CHR|1|37|filii Rauhel Naath Zara Samma Maza
1CHR|1|38|filii Seir Lothan Sobal Sebeon Ana Dison Eser Disan
1CHR|1|39|filii Lothan Horri Humam soror autem Lothan fuit Thamna
1CHR|1|40|filii Sobal Alian et Manaath et Ebal et Sepphi et Onam filii Sebeon Aia et Ana filii Ana Dison
1CHR|1|41|filii Dison Amaran et Eseban et Iethran et Charan
1CHR|1|42|filii Eser Balaan et Zaban et Iacan filii Dison Us et Aran
1CHR|1|43|isti sunt reges qui imperaverunt in terra Edom antequam esset rex super filios Israhel Bale filius Beor et nomen civitatis eius Denaba
1CHR|1|44|mortuus est autem Bale et regnavit pro eo Iobab filius Zare de Bosra
1CHR|1|45|cumque et Iobab fuisset mortuus regnavit pro eo Husam de terra Themanorum
1CHR|1|46|obiit quoque et Husam et regnavit pro eo Adad filius Badad qui percussit Madian in terra Moab et nomen civitatis eius Avith
1CHR|1|47|cumque et Adad fuisset mortuus regnavit pro eo Semla de Masreca
1CHR|1|48|sed et Semla mortuus est et regnavit pro eo Saul de Rooboth quae iuxta amnem sita est
1CHR|1|49|mortuo quoque Saul regnavit pro eo Baalanan filius Achobor
1CHR|1|50|sed et hic mortuus est et regnavit pro eo Adad cuius urbis fuit nomen Phou et appellata est uxor eius Mehetabel filia Matred filiae Mezaab
1CHR|1|51|Adad autem mortuo duces pro regibus in Edom esse coeperunt dux Thamna dux Alva dux Ietheth
1CHR|1|52|dux Oolibama dux Hela dux Phinon
1CHR|1|53|dux Cenez dux Theman dux Mabsar
1CHR|1|54|dux Magdihel dux Iram hii duces Edom
1CHR|2|1|filii autem Israhel Ruben Symeon Levi Iuda Isachar et Zabulon
1CHR|2|2|Dan Ioseph Beniamin Nepthali Gad Aser
1CHR|2|3|filii Iuda Her Aunan Sela tres nati sunt ei de filia Sue Chananitidis fuit autem Her primogenitus Iuda malus coram Domino et occidit eum
1CHR|2|4|Thamar autem nurus eius peperit ei Phares et Zara omnes ergo filii Iuda quinque
1CHR|2|5|filii autem Phares Esrom et Hamul
1CHR|2|6|filii quoque Zarae Zamri et Ethan et Eman Chalchal quoque et Darda simul quinque
1CHR|2|7|filii Carmi Achar qui turbavit Israhel et peccavit in furto anathematis
1CHR|2|8|filii Ethan Azarias
1CHR|2|9|filii autem Esrom qui nati sunt ei Ieremahel et Ram et Chalubi
1CHR|2|10|porro Ram genuit Aminadab Aminadab autem genuit Naasson principem filiorum Iuda
1CHR|2|11|Naasson quoque genuit Salma de quo ortus est Boez
1CHR|2|12|Boez vero genuit Obed qui et ipse genuit Isai
1CHR|2|13|Isai autem genuit primogenitum Heliab secundum Abinadab tertium Samaa
1CHR|2|14|quartum Nathanahel quintum Raddai
1CHR|2|15|sextum Asom septimum David
1CHR|2|16|quorum sorores fuerunt Sarvia et Abigail filii Sarviae Abisai Ioab et Asahel tres
1CHR|2|17|Abigail autem genuit Amasa cuius pater fuit Iether Ismahelites
1CHR|2|18|Chaleb vero filius Esrom accepit uxorem nomine Azuba de qua genuit Ierioth fueruntque filii eius Iesar et Sobab et Ardon
1CHR|2|19|cumque mortua fuisset Azuba accepit uxorem Chaleb Ephrath quae peperit ei Ur
1CHR|2|20|porro Ur genuit Uri et Uri genuit Beselehel
1CHR|2|21|post haec ingressus est Esrom ad filiam Machir patris Galaad et accepit eam cum esset annorum sexaginta quae peperit ei Segub
1CHR|2|22|sed et Segub genuit Iair et possedit viginti tres civitates in terra Galaad
1CHR|2|23|cepitque Gessur et Aram oppida Iair et Canath et viculos eius sexaginta civitatum omnes isti filii Machir patris Galaad
1CHR|2|24|cum autem mortuus esset Esrom ingressus est Chaleb ad Ephrata habuit quoque Esrom uxorem Abia quae peperit ei Assur patrem Thecue
1CHR|2|25|nati sunt autem filii Hieramehel primogeniti Esrom Ram primogenitus eius et Buna et Aran et Asom et Ahia
1CHR|2|26|duxit quoque uxorem alteram Hieramehel nomine Atara quae fuit mater Onam
1CHR|2|27|sed et filii Ram primogeniti Hieramehel fuerunt Moos et Iamin et Achar
1CHR|2|28|Onam autem habuit filios Semmei et Iada filii autem Semmei Nadab et Abisur
1CHR|2|29|nomen vero uxoris Abisur Abiail quae peperit Ahobban et Molid
1CHR|2|30|filii autem Nadab fuerunt Saled et Apphaim mortuus est autem Saled absque liberis
1CHR|2|31|filius vero Apphaim Iesi qui Iesi genuit Sesan porro Sesan genuit Oholi
1CHR|2|32|filii autem Iada fratris Semmei Iether et Ionathan sed et Iether mortuus est absque liberis
1CHR|2|33|porro Ionathan genuit Phaleth et Ziza isti fuerunt filii Hieramehel
1CHR|2|34|Sesan autem non habuit filios sed filias et servum aegyptium nomine Ieraa
1CHR|2|35|deditque ei filiam suam uxorem quae peperit ei Eththei
1CHR|2|36|Eththei autem genuit Nathan et Nathan genuit Zabad
1CHR|2|37|Zabad quoque genuit Ophlal et Ophlal genuit Obed
1CHR|2|38|Obed genuit Ieu Ieu genuit Azariam
1CHR|2|39|Azarias genuit Helles Helles genuit Elasa
1CHR|2|40|Elasa genuit Sisamoi Sisamoi genuit Sellum
1CHR|2|41|Sellum genuit Icamian Icamian genuit Elisama
1CHR|2|42|filii autem Chaleb fratris Hieramehel Mosa primogenitus eius ipse est pater Ziph et filii Maresa patris Hebron
1CHR|2|43|porro filii Hebron Core et Thapphu et Recem et Samma
1CHR|2|44|Samma autem genuit Raam patrem Iercaam et Recem genuit Semmei
1CHR|2|45|filius Semmei Maon et Maon pater Bethsur
1CHR|2|46|Epha autem concubina Chaleb peperit Arran et Musa et Gezez porro Arran genuit Gezez
1CHR|2|47|filii Iadai Regom et Iotham et Gesum et Phaleth et Epha et Saaph
1CHR|2|48|concubina Chaleb Maacha peperit Saber et Tharana
1CHR|2|49|genuit autem Saaph pater Madmena Sue patrem Machbena et patrem Gabaa filia vero Chaleb fuit Achsa
1CHR|2|50|hii erant filii Chaleb filii Ur primogeniti Ephrata Sobal pater Cariathiarim
1CHR|2|51|Salma pater Bethleem Ariph pater Bethgader
1CHR|2|52|fuerunt autem filii Sobal patris Cariathiarim qui videbat dimidium requietionum
1CHR|2|53|et de cognatione Cariathiarim Iethrei et Apphutei et Semathei et Maserei ex his egressi sunt Saraitae et Esthaolitae
1CHR|2|54|filii Salma Bethleem et Netophathi coronae domus Ioab et dimidium requietionis Sarai
1CHR|2|55|cognationes quoque scribarum habitantium in Iabis canentes atque resonantes et in tabernaculis commorantes hii sunt Cinei qui venerunt de calore patris domus Rechab
1CHR|3|1|David vero hos habuit filios qui ei nati sunt in Hebron primogenitum Amnon ex Achinaam Iezrahelitide secundum Danihel de Abigail Carmelitide
1CHR|3|2|tertium Absalom filium Maacha filiae Tholmei regis Gessur quartum Adoniam filium Aggith
1CHR|3|3|quintum Saphatiam ex Abital sextum Iethraam de Egla uxore sua
1CHR|3|4|sex ergo nati sunt ei in Hebron ubi regnavit septem annis et sex mensibus triginta autem et tribus annis regnavit in Hierusalem
1CHR|3|5|porro in Hierusalem nati sunt ei filii Samaa et Sobab et Nathan et Salomon quattuor de Bethsabee filia Amihel
1CHR|3|6|Iebaar quoque et Elisama
1CHR|3|7|et Eliphalet et Noge et Napheg et Iaphie
1CHR|3|8|necnon Elisama et Heliade et Eliphalet novem
1CHR|3|9|omnes hii filii David absque filiis concubinarum habuerunt sororem Thamar
1CHR|3|10|filius autem Salomonis Roboam cuius Abia filius genuit Asa de hoc quoque natus est Iosaphat
1CHR|3|11|pater Ioram qui Ioram genuit Ohoziam ex quo ortus est Ioas
1CHR|3|12|et huius Amasias filius genuit Azariam porro Azariae filius Ioatham
1CHR|3|13|procreavit Achaz patrem Ezechiae de quo natus est Manasses
1CHR|3|14|sed et Manasses genuit Amon patrem Iosiae
1CHR|3|15|filii autem Iosiae fuerunt primogenitus Iohanan secundus Ioacim tertius Sedecias quartus Sellum
1CHR|3|16|de Ioacim natus est Iechonias et Sedecias
1CHR|3|17|filii Iechoniae fuerunt Asir Salathihel
1CHR|3|18|Melchiram Phadaia Sennaser et Iecemia Sama et Nadabia
1CHR|3|19|de Phadaia orti sunt Zorobabel et Semei Zorobabel genuit Mosollam Ananiam et Salomith sororem eorum
1CHR|3|20|Asabamque et Ohol et Barachiam et Asadiam Iosabesed quinque
1CHR|3|21|filius autem Ananiae Phaltias pater Ieseiae cuius filius Raphaia huius quoque filius Arnam de quo natus est Obdia cuius filius fuit Sechenia
1CHR|3|22|filius Secheniae Semeia cuius filii Attus et Iegal et Baria et Naaria et Saphat sex numero
1CHR|3|23|filius Naariae Helioenai et Ezechias et Ezricam tres
1CHR|3|24|filii Helioenai Oduia et Heliasub et Pheleia et Accub et Iohanan et Dalaia et Anani septem
1CHR|4|1|filii Iuda Phares Esrom et Carmi et Ur et Subal
1CHR|4|2|Reaia vero filius Subal genuit Ieth de quo nati sunt Ahimai et Laed hae cognationes Sarathi
1CHR|4|3|ista quoque stirps Hetam Iezrahel et Iesema et Iedebos nomenque sororis eorum Asalelphuni
1CHR|4|4|Phunihel autem pater Gedor et Ezer pater Osa isti sunt filii Ur primogeniti Ephrata patris Bethleem
1CHR|4|5|Asur vero patris Thecue erant duae uxores Halaa et Naara
1CHR|4|6|peperit autem ei Naara Oozam et Epher et Themani et Asthari isti sunt filii Naara
1CHR|4|7|porro filii Halaa Sereth Isaar et Ethnan
1CHR|4|8|Cos autem genuit Anob et Sobaba et cognationem Aral filii Arum
1CHR|4|9|fuit autem Iabes inclitus prae fratribus suis et mater eius vocavit nomen illius Iabes dicens quia peperi eum in dolore
1CHR|4|10|invocavit vero Iabes Deum Israhel dicens si benedicens benedixeris mihi et dilataveris terminos meos et fuerit manus tua mecum et feceris me a malitia non opprimi et praestitit Deus quae precatus est
1CHR|4|11|Chaleb autem frater Suaa genuit Machir qui fuit pater Esthon
1CHR|4|12|porro Esthon genuit Bethrapha et Phesse et Thena patrem urbis Naas hii sunt viri Recha
1CHR|4|13|filii autem Cenez Othonihel et Saraia porro filii Othonihel Athath
1CHR|4|14|et Maonathi genuit Ophra Saraias autem genuit Ioab patrem vallis Artificum ibi quippe artifices erant
1CHR|4|15|filii vero Chaleb filii Iephonne Hir et Hela et Nahem filiique Hela et Cenez
1CHR|4|16|filii quoque Iallelel Ziph et Zipha Thiria et Asrahel
1CHR|4|17|et filii Ezra Iether et Mered et Epher et Ialon genuitque Mariam et Sammai et Iesba patrem Esthamo
1CHR|4|18|uxor quoque eius Iudaia peperit Iared patrem Gedor et Heber patrem Soccho et Hicuthihel patrem Zano hii autem filii Beththiae filiae Pharaonis quam accepit Mered
1CHR|4|19|et filii uxoris Odaiae sororis Naham patris Ceila Garmi et Esthamo qui fuit de Machathi
1CHR|4|20|filii quoque Simon Amnon et Rena filius Anan et Thilon et filii Iesi Zoeth et Benzoeth
1CHR|4|21|filii Sela filii Iuda Her pater Lecha et Laada pater Maresa et cognationes Domus operantium byssum in domo Iuramenti
1CHR|4|22|et Qui stare fecit solem virique Mendacii et Securus et Incendens qui principes fuerunt in Moab et qui reversi sunt in Leem haec autem verba vetera
1CHR|4|23|hii sunt figuli habitantes in plantationibus et in praesepibus apud regem in operibus eius commoratique sunt ibi
1CHR|4|24|filii Symeon Namuhel et Iamin Iarib Zara Saul
1CHR|4|25|Sellum filius eius Mabsam filius eius Masma filius eius
1CHR|4|26|filii Masma Amuhel filius eius Zacchur filius eius Semei filius eius
1CHR|4|27|filii Semei sedecim et filiae sex fratres autem eius non habuerunt filios multos et universa cognatio non potuit adaequare summam filiorum Iuda
1CHR|4|28|habitaverunt autem in Bersabee et Molada et Asarsual
1CHR|4|29|et in Ballaa et in Asom et in Tholad
1CHR|4|30|et in Bathuhel et in Orma et in Siceleg
1CHR|4|31|et in Bethmarchaboth et in Asarsusim et in Bethberai et in Saarim hae civitates eorum usque ad regem David
1CHR|4|32|villae quoque eorum Etham et Aen et Remmon et Thochen et Asan civitates quinque
1CHR|4|33|et universi viculi eorum per circuitum civitatum istarum usque ad Baal haec est habitatio eorum et sedum distributio
1CHR|4|34|Masobab quoque et Iemlech et Iosa filius Amasiae
1CHR|4|35|et Iohel et Ieu filius Iosabiae filii Saraiae filii Asihel
1CHR|4|36|et Helioenai et Iacoba et Isuaia et Asaia et Adihel et Isimihel et Banaia
1CHR|4|37|Ziza quoque filius Sephei filii Allon filii Idaia filii Semri filii Samaia
1CHR|4|38|isti sunt nominati principes in cognationibus suis et in domo adfinitatum suarum multiplicati sunt vehementer
1CHR|4|39|et profecti sunt ut ingrederentur in Gador usque ad orientem vallis et ut quaererent pascua gregibus suis
1CHR|4|40|inveneruntque pascuas uberes et valde bonas et terram latissimam et quietam et fertilem in qua ante habitaverunt de stirpe Ham
1CHR|4|41|hii ergo venerunt quos supra descripsimus nominatim in diebus Ezechiae regis Iuda et percusserunt tabernacula eorum et habitatores qui inventi fuerant ibi et deleverunt eos usque in praesentem diem habitaveruntque pro eis quoniam uberrimas ibidem pascuas reppererunt
1CHR|4|42|de filiis quoque Symeon abierunt in montem Seir viri quingenti habentes principes Phaltiam et Nahariam et Raphaiam et Ozihel filios Iesi
1CHR|4|43|et percusserunt reliquias quae evadere potuerant Amalechitarum et habitaverunt ibi pro eis usque ad diem hanc
1CHR|5|1|filii quoque Ruben primogeniti Israhel ipse quippe fuit primogenitus eius sed cum violasset torum patris sui data sunt primogenita eius filiis Ioseph filii Israhel et non est ille reputatus in primogenitum
1CHR|5|2|porro Iudas qui erat fortissimus inter fratres suos de stirpe eius principes germinati sunt primogenita autem reputata sunt Ioseph
1CHR|5|3|filii ergo Ruben primogeniti Israhel Enoch et Phallu Esrom et Charmi
1CHR|5|4|filii Iohel Samaia filius eius Gog filius eius Semei filius eius
1CHR|5|5|Micha filius eius Reeia filius eius Baal filius eius
1CHR|5|6|Beera filius eius quem captivum duxit Theglathphalnasar rex Assyriorum et fuit princeps in tribu Ruben
1CHR|5|7|fratres autem eius et universa cognatio quando numerabantur per familias suas habuerunt principes Ieihel et Zacchariam
1CHR|5|8|porro Bala filius Azaz filii Samma filii Iohel ipse habitavit in Aroer usque ad Nebo et Beelmeon
1CHR|5|9|contra orientalem quoque plagam habitavit usque ad introitum heremi et flumen Eufraten multum quippe iumentorum numerum possidebat in terra Galaad
1CHR|5|10|in diebus autem Saul proeliati sunt contra Agareos et interfecerunt illos habitaveruntque pro eis in tabernaculis eorum in omni plaga quae respicit ad orientem Galaad
1CHR|5|11|filii vero Gad e regione eorum habitaverunt in terra Basan usque Selcha
1CHR|5|12|Iohel in capite et Saphan secundus Ianai autem et Saphat in Basan
1CHR|5|13|fratres vero eorum secundum domos cognationum suarum Michahel et Mosollam et Sebe et Iori et Iachan et Zie et Heber septem
1CHR|5|14|hii filii Abiahil filii Uri filii Iaro filii Galaad filii Michahel filii Iesesi filii Ieddo filii Buz
1CHR|5|15|fratres quoque filii Abdihel filii Guni princeps domus in familiis suis
1CHR|5|16|et habitaverunt in Galaad et in Basan et in viculis eius et in cunctis suburbanis Saron usque ad terminos
1CHR|5|17|omnes hii numerati sunt in diebus Ioatham regis Iuda et in diebus Hieroboam regis Israhel
1CHR|5|18|filii Ruben et Gad et dimidiae tribus Manasse viri bellatores scuta portantes et gladios et tendentes arcum eruditique ad proelia quadraginta quattuor milia et septingenti sexaginta procedentes ad pugnam
1CHR|5|19|dimicaverunt contra Agarenos Iturei vero et Naphei et Nodab
1CHR|5|20|praebuerunt eis auxilium traditique sunt in manus eorum Agareni et universi qui fuerant cum eis quia Deum invocaverunt cum proeliarentur et exaudivit eos eo quod credidissent in eum
1CHR|5|21|ceperuntque omnia quae possederant camelorum quinquaginta milia et ovium ducenta quinquaginta milia asinos duo milia et animas hominum centum milia
1CHR|5|22|vulnerati autem multi corruerunt fuit enim bellum Domini habitaveruntque pro eis usque ad transmigrationem
1CHR|5|23|filii quoque dimidiae tribus Manasse possederunt terram a finibus Basan usque Baalhermon et Sanir et montem Hermon ingens quippe numerus erat
1CHR|5|24|et hii fuerunt principes domus cognationis eorum Epher et Iesi et Helihel Ezrihel et Hieremia et Odoia et Iedihel viri fortissimi et potentes et nominati duces in familiis suis
1CHR|5|25|reliquerunt autem Deum patrum suorum et fornicati sunt post deos populorum terrae quos abstulit Dominus coram eis
1CHR|5|26|et suscitavit Deus Israhel spiritum Ful regis Assyriorum et spiritum Theglathphalnasar regis Assur et transtulit Ruben et Gad et dimidium tribus Manasse et adduxit eos in Alae et Abor et Ara et fluvium Gozan usque ad diem hanc
1CHR|6|1|filii Levi Gersom Caath Merari
1CHR|6|2|filii Caath Amram Isaar Hebron et Ozihel
1CHR|6|3|filii Amram Aaron Moses et Maria filii Aaron Nadab et Abiu Eleazar et Ithamar
1CHR|6|4|Eleazar genuit Finees et Finees genuit Abisue
1CHR|6|5|Abisue vero genuit Bocci et Bocci genuit Ozi
1CHR|6|6|Ozi genuit Zaraiam et Zaraias genuit Meraioth
1CHR|6|7|porro Meraioth genuit Amariam et Amarias genuit Ahitob
1CHR|6|8|Ahitob genuit Sadoc Sadoc genuit Achimaas
1CHR|6|9|Achimaas genuit Azariam Azarias genuit Iohanan
1CHR|6|10|Iohanan genuit Azariam ipse est qui sacerdotio functus est in domo quam aedificavit Salomon in Hierusalem
1CHR|6|11|genuit autem Azarias Amariam et Amarias genuit Ahitob
1CHR|6|12|Ahitob genuit Sadoc et Sadoc genuit Sellum
1CHR|6|13|Sellum genuit Helciam et Helcias genuit Azariam
1CHR|6|14|Azarias genuit Saraiam et Saraias genuit Iosedec
1CHR|6|15|porro Iosedec egressus est quando transtulit Dominus Iudam et Hierusalem per manus Nabuchodonosor
1CHR|6|16|filii ergo Levi Gersom Caath et Merari
1CHR|6|17|et haec nomina filiorum Gersom Lobeni et Semei
1CHR|6|18|filii Caath Amram et Isaar et Hebron et Ozihel
1CHR|6|19|filii Merari Mooli et Musi hae autem cognationes Levi secundum familias eorum
1CHR|6|20|Gersom Lobeni filius eius Iaath filius eius Zamma filius eius
1CHR|6|21|Ioaa filius eius Addo filius eius Zara filius eius Iethrai filius eius
1CHR|6|22|filii Caath Aminadab filius eius Core filius eius Asir filius eius
1CHR|6|23|Helcana filius eius Abiasaph filius eius Asir filius eius
1CHR|6|24|Thaath filius eius Urihel filius eius Ozias filius eius Saul filius eius
1CHR|6|25|filii Helcana Amasai et Ahimoth
1CHR|6|26|Helcana filii Helcana Sophai filius eius Naath filius eius
1CHR|6|27|Heliab filius eius Hieroam filius eius Helcana filius eius
1CHR|6|28|filii Samuhel primogenitus Vasseni et Abia
1CHR|6|29|filii autem Merari Mooli Lobeni filius eius Semei filius eius Oza filius eius
1CHR|6|30|Samaa filius eius Aggia filius eius Asaia filius eius
1CHR|6|31|isti sunt quos constituit David super cantores domus Domini ex quo conlocata est arca
1CHR|6|32|et ministrabant coram tabernaculo testimonii canentes donec aedificaret Salomon domum Domini in Hierusalem stabant autem iuxta ordinem suum in ministerio
1CHR|6|33|hii vero sunt qui adsistebant cum filiis suis de filiis Caath Heman cantor filius Iohel filii Samuhel
1CHR|6|34|filii Helcana filii Hieroam filii Helihel filii Thou
1CHR|6|35|filii Suph filii Helcana filii Maath filii Amasai
1CHR|6|36|filii Helcana filii Iohel filii Azariae filii Sophoniae
1CHR|6|37|filii Thaath filii Asir filii Abiasaph filii Core
1CHR|6|38|filii Isaar filii Caath filii Levi filii Israhel
1CHR|6|39|et fratres eius Asaph qui stabat a dextris eius Asaph filius Barachiae filii Samaa
1CHR|6|40|filii Michahel filii Basiae filii Melchiae
1CHR|6|41|filii Athnai filii Zara filii Adaia
1CHR|6|42|filii Ethan filii Zamma filii Semei
1CHR|6|43|filii Ieth filii Gersom filii Levi
1CHR|6|44|filii autem Merari fratres eorum ad sinistram Ethan filius Cusi filii Abdi filii Maloch
1CHR|6|45|filii Asabiae filii Amasiae filii Helciae
1CHR|6|46|filii Amasai filii Bonni filii Somer
1CHR|6|47|filii Mooli filii Musi filii Merari filii Levi
1CHR|6|48|fratres quoque eorum Levitae qui ordinati sunt in cunctum ministerium tabernaculi domus Domini
1CHR|6|49|Aaron vero et filii eius adolebant incensum super altare holocausti et super altare thymiamatis in omne opus sancti sanctorum et ut precarentur pro Israhel iuxta omnia quae praecepit Moses servus Dei
1CHR|6|50|hii sunt autem filii Aaron Eleazar filius eius Finees filius eius Abisue filius eius
1CHR|6|51|Bocci filius eius Ozi filius eius Zaraia filius eius
1CHR|6|52|Meraioth filius eius Amaria filius eius Ahitob filius eius
1CHR|6|53|Sadoc filius eius Achimaas filius eius
1CHR|6|54|et haec habitacula eorum per vicos atque confinia filiorum scilicet Aaron iuxta cognationes Caathitarum ipsis enim sorte contigerat
1CHR|6|55|dederunt igitur eis Hebron in terra Iuda et suburbana eius per circuitum
1CHR|6|56|agros autem civitatis et villas Chaleb filio Iephonne
1CHR|6|57|porro filiis Aaron dederunt civitates ad confugiendum Hebron et Lobna et suburbana eius
1CHR|6|58|Iether quoque et Esthmo cum suburbanis suis sed et Helon et Dabir cum suburbanis suis
1CHR|6|59|Asan quoque et Bethsemes et suburbana eorum
1CHR|6|60|de tribu autem Beniamin Gabee et suburbana eius et Almath cum suburbanis suis Anathoth quoque cum suburbanis suis omnes civitates tredecim per cognationes suas
1CHR|6|61|filiis autem Caath residuis de cognatione sua dederunt ex dimidia tribu Manasse in possessionem urbes decem
1CHR|6|62|porro filiis Gersom per cognationes suas de tribu Isachar et de tribu Aser et de tribu Nepthali et de tribu Manasse in Basan urbes tredecim
1CHR|6|63|filiis autem Merari per cognationes suas de tribu Ruben et de tribu Gad et de tribu Zabulon dederunt sorte civitates duodecim
1CHR|6|64|dederunt quoque filii Israhel Levitis civitates et suburbana earum
1CHR|6|65|dederuntque per sortem ex tribu filiorum Iuda et ex tribu filiorum Symeon et ex tribu filiorum Beniamin urbes has quas vocaverunt nominibus suis
1CHR|6|66|et his qui erant ex cognatione filiorum Caath fueruntque civitates in terminis eorum de tribu Ephraim
1CHR|6|67|dederunt ergo eis urbes ad confugiendum Sychem cum suburbanis suis in monte Ephraim et Gazer cum suburbanis suis
1CHR|6|68|Hicmaam quoque cum suburbanis suis et Bethoron similiter
1CHR|6|69|necnon et Helon cum suburbanis suis et Gethremmon in eundem modum
1CHR|6|70|porro ex dimidia tribu Manasse Aner et suburbana eius Balaam et suburbana eius his videlicet qui de cognatione filiorum Caath reliqui erant
1CHR|6|71|filiis autem Gersom de cognatione dimidiae tribus Manasse Gaulon in Basan et suburbana eius et Astharoth cum suburbanis suis
1CHR|6|72|de tribu Isachar Cedes et suburbana eius et Dabereth cum suburbanis suis
1CHR|6|73|Ramoth quoque et suburbana illius et Anem cum suburbanis suis
1CHR|6|74|de tribu vero Aser Masal cum suburbanis suis et Abdon similiter
1CHR|6|75|Acac quoque et suburbana eius et Roob cum suburbanis suis
1CHR|6|76|porro de tribu Nepthali Cedes in Galilea et suburbana eius Amon cum suburbanis suis et Cariathaim et suburbana eius
1CHR|6|77|filiis autem Merari residuis de tribu Zabulon Remmono et suburbana eius et Thabor cum suburbanis suis
1CHR|6|78|trans Iordanem quoque ex adverso Hiericho contra orientem Iordanis de tribu Ruben Bosor in solitudine cum suburbanis suis et Iasa cum suburbanis suis
1CHR|6|79|Cademoth quoque et suburbana eius et Miphaath cum suburbanis suis
1CHR|6|80|necnon de tribu Gad Ramoth in Galaad et suburbana eius et Manaim cum suburbanis suis
1CHR|6|81|sed et Esbon cum suburbanis eius et Iezer cum suburbanis suis
1CHR|7|1|porro filii Isachar Thola et Phua Iasub et Samaron quattuor
1CHR|7|2|filii Thola Ozi et Raphaia et Ierihel et Iemai et Iebsem et Samuhel principes per domos cognationum suarum de stirpe Thola viri fortissimi numerati sunt in diebus David viginti duo milia sescenti
1CHR|7|3|filii Ozi Iezraia de quo nati sunt Michahel et Obadia et Iohel et Iesia quinque omnes principes
1CHR|7|4|cumque eis per familias et populos suos accincti ad proelium viri fortissimi triginta sex milia multas enim habuere uxores et filios
1CHR|7|5|fratresque eorum per omnem cognationem Isachar robustissimi ad pugnandum octoginta septem milia numerati sunt
1CHR|7|6|Beniamin Bale et Bochor et Iadihel tres
1CHR|7|7|filii Bale Esbon et Ozi et Ozihel et Ierimoth et Urai quinque principes familiarum et ad pugnandum robustissimi numerus autem eorum viginti duo milia et triginta quattuor
1CHR|7|8|porro filii Bochor Zamira et Ioas et Eliezer et Helioenai et Amri et Ierimoth et Abia et Anathoth et Almathan omnes hii filii Bochor
1CHR|7|9|numerati sunt autem per familias suas principes cognationum ad bella fortissimi viginti milia et ducenti
1CHR|7|10|porro filii Iadihel Balan filii autem Balan Hieus et Beniamin et Ahoth et Chanana et Iothan et Tharsis et Haisaar
1CHR|7|11|omnes hii filii Iadihel principes cognationum suarum viri fortissimi decem et septem milia et ducenti ad proelium procedentes
1CHR|7|12|Sephan quoque et Apham filii Hir et Asim filii Aer
1CHR|7|13|filii autem Nepthali Iasihel et Guni et Asar et Sellum filii Balaa
1CHR|7|14|porro filius Manasse Esrihel concubinaque eius syra peperit Machir patrem Galaad
1CHR|7|15|Machir autem accepit uxores filiis suis Happhim et Sepham et habuit sororem nomine Maacha nomen autem secundi Salphaad nataeque sunt Salphaad filiae
1CHR|7|16|et peperit Maacha uxor Machir filium vocavitque nomen eius Phares porro nomen fratris eius Sares et filii eius Ulam et Recem
1CHR|7|17|filius autem Ulam Badan hii sunt filii Galaad filii Machir filii Manasse
1CHR|7|18|soror autem eius Regina peperit virum Decorum et Abiezer et Moola
1CHR|7|19|erant autem filii Semida Ahin et Sechem et Leci et Aniam
1CHR|7|20|filii autem Ephraim Suthala Bareth filius eius Thaath filius eius Elada filius eius Thaath filius eius et huius filius Zabad
1CHR|7|21|et huius filius Suthala et huius filius Ezer et Elad occiderunt autem eos viri Geth indigenae quia descenderant ut invaderent possessiones eorum
1CHR|7|22|luxit igitur Ephraim pater eorum multis diebus et venerunt fratres eius ut consolarentur eum
1CHR|7|23|ingressusque est ad uxorem suam quae concepit et peperit filium et vocavit nomen eius Beria eo quod in malis domus eius ortus esset
1CHR|7|24|filia autem eius fuit Sara quae aedificavit Bethoron inferiorem et superiorem et Ozensara
1CHR|7|25|porro filius eius Rapha et Reseph et Thale de quo natus est Thaan
1CHR|7|26|qui genuit Laadan huius quoque filius Ammiud genuit Elisama
1CHR|7|27|de quo ortus est Nun qui habuit filium Iosue
1CHR|7|28|possessio autem eorum et habitatio Bethel cum filiabus suis et contra orientem Noran ad occidentalem plagam Gazer et filiae eius Sychem quoque cum filiabus suis usque Aza et filias eius
1CHR|7|29|iuxta filios quoque Manasse Bethsan et filias eius Thanach et filias eius Mageddo et filias eius Dor et filias eius in his habitaverunt filii Ioseph filii Israhel
1CHR|7|30|filii Aser Iomna et Iesua et Isui et Baria et Sara soror eorum
1CHR|7|31|filii autem Baria Heber et Melchihel ipse est pater Barzaith
1CHR|7|32|Heber autem genuit Iephlat et Somer et Otham et Suaa sororem eorum
1CHR|7|33|filii Iephlat Phosech et Chamaal et Asoth hii filii Iephlat
1CHR|7|34|porro filii Somer Ahi et Roaga et Iaba et Aram
1CHR|7|35|filii autem Helem fratris eius Supha et Iemna et Selles et Amal
1CHR|7|36|filii Supha Sue Arnaphed et Sual et Beri et Iamra
1CHR|7|37|Bosor et Od et Samma et Salusa et Iethran et Bera
1CHR|7|38|filii Iether Iephonne et Phaspha et Ara
1CHR|7|39|filii autem Olla Aree et Anihel et Resia
1CHR|7|40|omnes hii filii Aser principes cognationum electi atque fortissimi duces ducum numerus autem eorum aetatis quae apta esset ad bellum viginti sex milia
1CHR|8|1|Beniamin autem genuit Bale primogenitum suum Asbal secundum Ohora tertium
1CHR|8|2|Nuaha quartum et Rapha quintum
1CHR|8|3|fueruntque filii Bale Addaor et Gera et Abiud
1CHR|8|4|Abisue quoque et Neman et Ahoe
1CHR|8|5|sed et Gera et Sephuphan et Uram
1CHR|8|6|hii sunt filii Aod principes cognationum habitantium in Gabaa qui translati sunt in Manath
1CHR|8|7|Nooman autem et Achia et Gera ipse transtulit eos et genuit Oza et Ahiud
1CHR|8|8|porro Saarim genuit in regione Moab postquam dimisit Usim et Bara uxores suas
1CHR|8|9|genuit autem de Edes uxore sua Iobab et Sebia et Mosa et Molchom
1CHR|8|10|Iehus quoque et Sechia et Marma hii sunt filii eius principes in familiis suis
1CHR|8|11|Meusim vero genuit Abitob et Elphaal
1CHR|8|12|porro filii Elphaal Heber et Misaam et Samad hic aedificavit Ono et Lod et filias eius
1CHR|8|13|Bara autem et Samma principes cognationum habitantium in Aialon hii fugaverunt habitatores Geth
1CHR|8|14|et Haio et Sesac et Ierimoth
1CHR|8|15|et Zabadia et Arod et Eder
1CHR|8|16|Michahel quoque et Iespha et Ioaa filii Baria
1CHR|8|17|et Zabadia et Mosollam et Ezeci et Heber
1CHR|8|18|et Iesamari et Iezlia et Iobab filii Elphaal
1CHR|8|19|et Iacim et Zechri et Zabdi
1CHR|8|20|et Helioenai et Selethai et Helihel
1CHR|8|21|et Adaia et Baraia et Samarath filii Semei
1CHR|8|22|et Iesphan et Heber et Helihel
1CHR|8|23|et Abdon et Zechri et Hanan
1CHR|8|24|et Anania et Ailam et Anathothia
1CHR|8|25|et Iephdaia et Phanuhel filii Sesac
1CHR|8|26|et Samsari et Sooria et Otholia
1CHR|8|27|et Iersia et Helia et Zechri filii Ieroam
1CHR|8|28|hii patriarchae et cognationum principes qui habitaverunt in Hierusalem
1CHR|8|29|in Gabaon autem habitaverunt Abigabaon et nomen uxoris eius Maacha
1CHR|8|30|filiusque eius primogenitus Abdon et Sur et Cis et Baal et Nadab
1CHR|8|31|Gedor quoque et Ahio et Zacher
1CHR|8|32|et Macelloth genuit Samaa habitaveruntque ex adverso fratrum suorum in Hierusalem cum fratribus suis
1CHR|8|33|Ner autem genuit Cis et Cis genuit Saul porro Saul genuit Ionathan et Melchisuae et Abinadab et Esbaal
1CHR|8|34|filius autem Ionathan Meribbaal et Meribbaal genuit Micha
1CHR|8|35|filii Micha Phithon et Melech et Thara et Ahaz
1CHR|8|36|et Ahaz genuit Ioada et Ioada genuit Almoth et Azmoth et Zamari porro Zamari genuit Mosa
1CHR|8|37|et Mosa genuit Baana cuius filius fuit Rapha de quo ortus est Elasa qui genuit Asel
1CHR|8|38|porro Asel sex filii fuere his nominibus Ezricam Bochru Ismahel Saria Abadia Anan omnes hii filii Asel
1CHR|8|39|filii autem Esec fratris eius Ulam primogenitus et Us secundus et Eliphalet tertius
1CHR|8|40|fueruntque filii Ulam viri robustissimi et magno robore tendentes arcum et multos habentes filios ac nepotes usque ad centum quinquaginta omnes hii filii Beniamin
1CHR|9|1|universus ergo Israhel dinumeratus est et summa eorum scripta est in libro regum Israhel et Iuda translatique sunt in Babylonem propter delictum suum
1CHR|9|2|qui autem habitaverunt primi in possessionibus et in urbibus suis Israhel et sacerdotes Levitae et Nathinnei
1CHR|9|3|commorati sunt in Hierusalem de filiis Iuda et de filiis Beniamin de filiis quoque Ephraim et Manasse
1CHR|9|4|Othei filius Amiud filius Emri filii Omrai filii Bonni de filiis Phares filii Iuda
1CHR|9|5|et de Siloni Asaia primogenitus et filii eius
1CHR|9|6|de filiis autem Zara Ieuhel et fratres eorum sescenti nonaginta
1CHR|9|7|porro de filiis Beniamin Salo filius Mosollam filii Oduia filii Asana
1CHR|9|8|et Iobania filius Hieroam et Hela filius Ozi filii Mochori et Mosollam filius Saphatiae filii Rahuhel filii Iebaniae
1CHR|9|9|et fratres eorum per familias suas nongenti quinquaginta sex omnes hii principes cognationum per domos patrum suorum
1CHR|9|10|de sacerdotibus autem Iedaia Ioiarib et Iachin
1CHR|9|11|Azarias quoque filius Helciae filii Mosollam filii Sadoc filii Maraioth filii Ahitob pontifex domus Dei
1CHR|9|12|porro Adaias filius Hieroam filii Phasor filii Melchia et Masaia filius Adihel filii Iezra filii Mosollam filii Mosollamoth filii Emmer
1CHR|9|13|fratres quoque eorum principes per familias suas mille septingenti sexaginta fortissimi robore ad faciendum opus ministerii in domo Dei
1CHR|9|14|de Levitis autem Semeia filius Assub filii Ezricam filii Asebiu de filiis Merari
1CHR|9|15|Bacbacar quoque carpentarius et Galal et Mathania filius Micha filii Zechri filii Asaph
1CHR|9|16|et Obdia filius Semeiae filii Galal filii Idithun et Barachia filius Asa filii Helcana qui habitavit in atriis Netophathi
1CHR|9|17|ianitores autem Sellum et Acub et Telmon et Ahiman et frater eorum Sellum princeps
1CHR|9|18|usque ad illud tempus in porta Regis ad orientem observabant per vices suas de filiis Levi
1CHR|9|19|Sellum vero filius Core filii Abiasaph filii Core cum fratribus suis et domo patris sui hii sunt Coritae super opera ministerii custodes vestibulorum tabernaculi et familiae eorum per vices castrorum Domini custodientes introitum
1CHR|9|20|Finees autem filius Eleazar erat dux eorum coram Domino
1CHR|9|21|porro Zaccharias filius Mosollamia ianitor portae tabernaculi testimonii
1CHR|9|22|omnes hii electi in ostiarios per portas ducenti duodecim et descripti in villis propriis quos constituerunt David et Samuhel videns in fide sua
1CHR|9|23|tam ipsos quam filios eorum in ostiis domus Domini et in tabernaculo vicibus suis
1CHR|9|24|per quattuor ventos erant ostiarii id est ad orientem et ad occidentem ad aquilonem et ad austrum
1CHR|9|25|fratres autem eorum in viculis morabantur et veniebant in sabbatis suis de tempore usque ad tempus
1CHR|9|26|his quattuor Levitis creditus erat omnis numerus ianitorum et erant super exedras et thesauros domus Domini
1CHR|9|27|per gyrum quoque templi Domini morabantur in custodiis suis ut cum tempus fuisset ipsi mane aperirent fores
1CHR|9|28|de horum grege erant et super vasa ministerii ad numerum enim et inferebantur vasa et efferebantur
1CHR|9|29|de ipsis et qui credita habebant utensilia sanctuarii praeerant similae et vino et oleo et turi et aromatibus
1CHR|9|30|filii autem sacerdotum unguenta ex aromatibus conficiebant
1CHR|9|31|et Matthathias Levites primogenitus Sellum Coritae praefectus erat eorum quae in sartagine frigebantur
1CHR|9|32|porro de filiis Caath fratribus eorum super panes erant propositionis ut semper novos per singula sabbata praepararent
1CHR|9|33|hii sunt principes cantorum per familias Levitarum qui in exedris morabantur ita ut die et nocte iugiter suo ministerio deservirent
1CHR|9|34|capita Levitarum per familias suas principes manserunt in Hierusalem
1CHR|9|35|in Gabaon autem commorati sunt pater Gabaon Iaihel et nomen uxoris eius Maacha
1CHR|9|36|filius primogenitus eius Abdon et Sur et Cis et Baal et Ner et Nadab
1CHR|9|37|Gedor quoque et Ahio et Zaccharias et Macelloth
1CHR|9|38|porro Macelloth genuit Semmaam isti habitaverunt e regione fratrum suorum in Hierusalem cum fratribus suis
1CHR|9|39|Ner autem genuit Cis et Cis genuit Saul et Saul genuit Ionathan et Melchisuae et Abinadab et Esbaal
1CHR|9|40|filius autem Ionathan Meribbaal et Meribbaal genuit Micha
1CHR|9|41|porro filii Micha Phiton et Malech et Thara
1CHR|9|42|Ahaz autem genuit Iara et Iara genuit Alamath et Azmoth et Zamri et Zamri genuit Mosa
1CHR|9|43|Mosa vero genuit Baana cuius filius Raphaia genuit Elasa de quo ortus est Esel
1CHR|9|44|porro Esel sex filios habuit his nominibus Ezricam Bochru Ismahel Saria Obdia Anan hii filii Esel
1CHR|10|1|Philisthim autem pugnabant contra Israhel fugeruntque viri Israhel Palestinos et ceciderunt vulnerati in monte Gelboe
1CHR|10|2|cumque adpropinquassent Philisthei persequentes Saul et filios eius percusserunt Ionathan et Abinadab et Melchisuae filios Saul
1CHR|10|3|et adgravatum est proelium contra Saul inveneruntque eum sagittarii et vulneraverunt iaculis
1CHR|10|4|et dixit Saul ad armigerum suum evagina gladium tuum et interfice me ne forte veniant incircumcisi isti et inludant mihi noluit autem armiger eius hoc facere timore perterritus arripuit igitur Saul ensem et inruit in eum
1CHR|10|5|quod cum vidisset armiger eius videlicet mortuum esse Saul inruit etiam ipse in gladium suum et mortuus est
1CHR|10|6|interiit ergo Saul et tres filii eius et omnis domus illius pariter concidit
1CHR|10|7|quod cum vidissent viri Israhel qui habitabant in campestribus fugerunt et Saul ac filiis eius mortuis dereliquerunt urbes suas et huc illucque dispersi sunt veneruntque Philisthim et habitaverunt in eis
1CHR|10|8|die igitur altero detrahentes Philisthim spolia caesorum invenerunt Saul et filios eius iacentes in monte Gelboe
1CHR|10|9|cumque spoliassent eum et amputassent caput armisque nudassent miserunt in terram suam ut circumferretur et ostenderetur idolorum templis et populis
1CHR|10|10|arma autem eius consecraverunt in fano dei sui et caput adfixerunt in templo Dagon
1CHR|10|11|hoc cum audissent viri Iabesgalaad omnia scilicet quae Philisthim fecerunt super Saul
1CHR|10|12|consurrexerunt singuli virorum fortium et tulerunt cadavera Saul et filiorum eius adtuleruntque ea in Iabes et sepelierunt ossa eorum subter quercum quae erat in Iabes et ieiunaverunt septem diebus
1CHR|10|13|mortuus est ergo Saul propter iniquitates suas eo quod praevaricatus sit mandatum Domini quod praeceperat et non custodierit illud sed insuper etiam pythonissam consuluerit
1CHR|10|14|nec speraverit in Domino propter quod et interfecit eum et transtulit regnum eius ad David filium Isai
1CHR|11|1|congregatus est igitur omnis Israhel ad David in Hebron dicens os tuum sumus et caro tua
1CHR|11|2|heri quoque et nudius tertius cum adhuc regnaret Saul tu eras qui educebas et introducebas Israhel tibi enim dixit Dominus Deus tuus tu pasces populum meum Israhel et tu eris princeps super eum
1CHR|11|3|venerunt ergo omnes maiores natu Israhel ad regem in Hebron et iniit David cum eis foedus coram Domino unxeruntque eum regem super Israhel iuxta sermonem Domini quem locutus est in manu Samuhel
1CHR|11|4|abiit quoque David et omnis Israhel in Hierusalem haec est Iebus ubi erant Iebusei habitatores terrae
1CHR|11|5|dixeruntque qui habitabant in Iebus ad David non ingredieris huc porro David cepit arcem Sion quae est civitas David
1CHR|11|6|dixitque omnis qui percusserit Iebuseum in primis erit princeps et dux ascendit igitur primus Ioab filius Sarviae et factus est princeps
1CHR|11|7|habitavit autem David in arce et idcirco appellata est civitas David
1CHR|11|8|aedificavitque urbem in circuitu a Mello usque ad gyrum Ioab autem reliqua urbis extruxit
1CHR|11|9|proficiebatque David vadens et crescens et Dominus exercituum erat cum eo
1CHR|11|10|hii principes virorum fortium David qui adiuverunt eum ut rex fieret super omnem Israhel iuxta verbum Domini quod locutus est ad Israhel
1CHR|11|11|et iste numerus robustorum David Iesbaam filius Achamoni princeps inter triginta iste levavit hastam suam super trecentos vulneratos una vice
1CHR|11|12|et post eum Eleazar filius patrui eius Ahoites qui erat inter tres potentes
1CHR|11|13|iste fuit cum David in Aphesdommim quando Philisthim congregati sunt ad locum illum in proelium et erat ager regionis illius plenus hordeo fugeratque populus a facie Philisthinorum
1CHR|11|14|hic stetit in medio agri et defendit eum cumque percussisset Philistheos dedit Dominus salutem magnam populo suo
1CHR|11|15|descenderunt autem tres de triginta principibus ad petram in qua erat David ad speluncam Odollam quando Philisthim fuerant castrametati in valle Raphaim
1CHR|11|16|porro David erat in praesidio et statio Philisthinorum in Bethleem
1CHR|11|17|desideravit igitur David et dixit o si quis daret mihi aquam de cisterna Bethleem quae est in porta
1CHR|11|18|tres ergo isti per media castra Philisthinorum perrexerunt et hauserunt aquam de cisterna Bethleem quae erat in porta et adtulerunt ad David ut biberet qui noluit sed magis libavit illam Domino
1CHR|11|19|dicens absit ut in conspectu Dei mei hoc faciam et sanguinem virorum istorum bibam quia in periculo animarum suarum adtulerunt mihi aquam et ob hanc causam noluit bibere haec fecerunt tres robustissimi
1CHR|11|20|Abisai quoque frater Ioab ipse erat princeps trium et ipse levavit hastam suam contra trecentos vulneratos et ipse erat inter tres nominatissimus
1CHR|11|21|inter tres secundos inclitus et princeps eorum verumtamen usque ad tres primos non pervenerat
1CHR|11|22|Banaia filius Ioiadae viri robustissimi qui multa opera perpetrarat de Capsehel ipse percussit duos Arihel Moab et ipse descendit et interfecit leonem in media cisterna tempore nivis
1CHR|11|23|et ipse percussit virum aegyptium cuius statura erat quinque cubitorum et habebat lanceam ut liciatorium texentium descendit ergo ad eum cum virga et rapuit hastam quam tenebat manu et interfecit eum hasta sua
1CHR|11|24|haec fecit Banaia filius Ioiada qui erat inter tres robustos nominatissimus
1CHR|11|25|inter triginta primus verumtamen ad tres usque non pervenerat posuit autem eum David ad auriculam suam
1CHR|11|26|porro fortissimi in exercitu Asahel frater Ioab et Eleanan filius patrui eius de Bethleem
1CHR|11|27|Semmoth Arorites Helles Phallonites
1CHR|11|28|Iras filius Acces Thecuites Abiezer Anathothites
1CHR|11|29|Sobbochai Asothites Ilai Ahoites
1CHR|11|30|Marai Netophathites Heled filius Baana Netophathites
1CHR|11|31|Ethai filius Ribai de Gabaath filiorum Beniamin Banaia Pharathonites
1CHR|11|32|Uri de torrente Gaas Abial Arabathites Azmoth Bauramites Eliaba Salabonites
1CHR|11|33|filii Asom Gezonites Ionathan filius Sega Ararites
1CHR|11|34|Ahiam filius Sachar Ararites
1CHR|11|35|Eliphal filius Ur
1CHR|11|36|Apher Mechurathites Ahia Phellonites
1CHR|11|37|Asrai Carmelites Noorai filius Azbi
1CHR|11|38|Iohel frater Nathan Mabar filius Agarai
1CHR|11|39|Sellec Ammonites Noorai Berothites armiger Ioab filii Sarviae
1CHR|11|40|Iras Iethreus Gareb Iethreus
1CHR|11|41|Urias Ettheus Zabad filius Ooli
1CHR|11|42|Adina filius Seza Rubenites princeps Rubenitarum et cum eo triginta
1CHR|11|43|Hanan filius Maacha et Iosaphat Mathanites
1CHR|11|44|Ozias Astharothites Semma et Iaihel filii Hotam Aroerites
1CHR|11|45|Iedihel filius Samri et Ioha frater eius Thosaites
1CHR|11|46|Elihel Maumites et Ieribai et Iosaia filii Elnaem et Iethma Moabites Elihel et Obed et Iasihel de Masobia
1CHR|12|1|hii quoque venerunt ad David in Siceleg cum adhuc fugeret Saul filium Cis qui erant fortissimi et egregii pugnatores
1CHR|12|2|tendentes arcum et utraque manu fundis saxa iacientes et dirigentes sagittas de fratribus Saul ex Beniamin
1CHR|12|3|princeps Ahiezer et Ioas filii Sammaa Gabathites et Iazihel et Phallet filii Azmoth et Baracha et Ieu Anathothites
1CHR|12|4|Samaias quoque Gabaonites fortissimus inter triginta et super triginta Hieremias et Iezihel et Iohanan et Iezbad Gaderothites
1CHR|12|5|Eluzai et Ierimuth et Baalia et Samaria et Saphatia Aruphites
1CHR|12|6|Helcana et Iesia et Azrahel et Ioezer et Iesbaam de Careim
1CHR|12|7|Ioeela quoque et Zabadia filii Ieroam de Gedor
1CHR|12|8|sed et de Gaddi transfugerunt ad David cum lateret in deserto viri robustissimi et pugnatores optimi tenentes clypeum et hastam facies eorum quasi facies leonis et veloces quasi capreae in montibus
1CHR|12|9|Ezer princeps Obdias secundus Eliab tertius
1CHR|12|10|Masmana quartus Hieremias quintus
1CHR|12|11|Hetthi sextus Helihel septimus
1CHR|12|12|Iohanan octavus Helzebad nonus
1CHR|12|13|Hieremias decimus Bachannai undecimus
1CHR|12|14|hii de filiis Gad principes exercitus novissimus centum militibus praeerat et maximus mille
1CHR|12|15|isti sunt qui transierunt Iordanem mense primo quando inundare consuevit super ripas suas et omnes fugaverunt qui morabantur in vallibus ad orientalem plagam et occidentalem
1CHR|12|16|venerunt autem et de Beniamin et de Iuda ad praesidium in quo morabatur David
1CHR|12|17|egressusque est David obviam eis et ait si pacifice venistis ad me ut auxiliemini mihi cor meum iungatur vobis si autem insidiamini mihi pro adversariis meis cum ego iniquitatem in manibus non habeam videat Deus patrum nostrorum et iudicet
1CHR|12|18|spiritus vero induit Amessai principem inter triginta et ait tui sumus o David et tecum fili Isai pax pax tibi et pax adiutoribus tuis te enim adiuvat Deus tuus suscepit ergo eos David et constituit principes turmae
1CHR|12|19|porro de Manasse transfugerunt ad David quando veniebat cum Philisthim adversum Saul ut pugnaret et non dimicavit cum eis quia inito consilio remiserunt eum principes Philisthinorum dicentes periculo capitis nostri revertetur ad dominum suum Saul
1CHR|12|20|quando igitur reversus est in Siceleg transfugerunt ad eum de Manasse Ednas et Iozabad et Iedihel et Michahel et Iozabad et Heliu et Salathi principes milium in Manasse
1CHR|12|21|hii praebuerunt auxilium David adversum latrunculos omnes enim erant viri fortissimi et facti sunt principes in exercitu
1CHR|12|22|sed et per singulos dies veniebant ad David ad auxiliandum ei usque dum fieret grandis numerus quasi exercitus Dei
1CHR|12|23|iste quoque est numerus principum exercitus qui venerunt ad David cum esset in Hebron ut transferrent regnum Saul ad eum iuxta verbum Domini
1CHR|12|24|filii Iuda portantes clypeum et hastam sex milia octingenti expediti ad proelium
1CHR|12|25|de filiis Symeon virorum fortissimorum ad pugnandum septem milia centum
1CHR|12|26|de filiis Levi quattuor milia sescenti
1CHR|12|27|Ioiada quoque princeps de stirpe Aaron et cum eo tria milia septingenti
1CHR|12|28|Sadoc etiam puer egregiae indolis et domus patris eius principes viginti duo
1CHR|12|29|de filiis autem Beniamin fratribus Saul tria milia magna enim pars eorum adhuc sequebatur domum Saul
1CHR|12|30|porro de filiis Ephraim viginti milia octingenti fortissimi robore viri nominati in cognationibus suis
1CHR|12|31|et ex dimidia parte tribus Manasse decem et octo milia singuli per nomina sua venerunt ut constituerent regem David
1CHR|12|32|de filiis quoque Isachar viri eruditi qui norant singula tempora ad praecipiendum quid facere deberet Israhel principes ducenti omnis autem reliqua tribus eorum consilium sequebatur
1CHR|12|33|porro de Zabulon qui egrediebantur ad proelium et stabant in acie instructi armis bellicis quinquaginta milia venerunt in auxilium non in corde duplici
1CHR|12|34|et de Nepthali principes mille et cum eis instructa clypeo et hasta triginta septem milia
1CHR|12|35|de Dan etiam praeparata ad proelium viginti octo milia sescentorum
1CHR|12|36|et de Aser egredientes ad pugnam et in acie provocantes quadraginta milia
1CHR|12|37|trans Iordanem autem de filiis Ruben et Gad et dimidia parte tribus Manasse instructa armis bellicis centum viginti milia
1CHR|12|38|omnes isti viri bellatores et expediti ad pugnandum corde perfecto venerunt in Hebron ut constituerent regem David super universum Israhel sed et omnes reliqui ex Israhel uno corde erant ut rex fieret David
1CHR|12|39|fueruntque ibi apud David tribus diebus comedentes et bibentes praeparaverunt enim eis fratres sui
1CHR|12|40|sed et qui iuxta eos erant usque ad Isachar et Zabulon et Nepthalim adferebant panes in asinis et camelis et mulis et bubus ad vescendum farinam palatas uvam passam vinum oleum boves arietes ad omnem copiam gaudium quippe erat in Israhel
1CHR|13|1|iniit autem consilium David cum tribunis et centurionibus et universis principibus
1CHR|13|2|et ait ad omnem coetum Israhel si placet vobis et a Domino Deo nostro egreditur sermo quem loquor mittamus ad fratres nostros reliquos in universas regiones Israhel et ad sacerdotes et Levitas qui habitant in suburbanis urbium ut congregentur ad nos
1CHR|13|3|et reducamus arcam Dei nostri ad nos non enim requisivimus eam in diebus Saul
1CHR|13|4|et respondit universa multitudo ut ita fieret placuerat enim sermo omni populo
1CHR|13|5|congregavit ergo David cunctum Israhel a Sior Aegypti usque dum ingrediaris Emath ut adduceret arcam Dei de Cariathiarim
1CHR|13|6|et ascendit David et omnis vir Israhel ad collem Cariathiarim quae est in Iuda ut adferrent inde arcam Dei Domini sedentis super cherubin ubi invocatum est nomen eius
1CHR|13|7|inposueruntque arcam Dei super plaustrum novum de domo Aminadab Oza autem et fratres eius minabant plaustrum
1CHR|13|8|porro David et universus Israhel ludebant coram Deo omni virtute in canticis et in citharis et psalteriis et tympanis et cymbalis et tubis
1CHR|13|9|cum autem pervenissent ad aream Chidon tetendit Oza manum suam ut sustentaret arcam bos quippe lasciviens paululum inclinaverat eam
1CHR|13|10|iratus est itaque Dominus contra Ozam et percussit eum eo quod contigisset arcam et mortuus est ibi coram Deo
1CHR|13|11|contristatusque David eo quod divisisset Dominus Ozam vocavit locum illum Divisio Oza usque in praesentem diem
1CHR|13|12|et timuit Deum tunc temporis dicens quomodo possum ad me introducere arcam Dei
1CHR|13|13|et ob hanc causam non eam adduxit ad se hoc est in civitatem David sed avertit in domum Obededom Getthei
1CHR|13|14|mansit ergo arca Dei in domo Obededom tribus mensibus et benedixit Dominus domui eius et omnibus quae habebat
1CHR|14|1|misit quoque Hiram rex Tyri nuntios ad David et ligna cedrina et artifices parietum lignorumque ut aedificarent ei domum
1CHR|14|2|cognovitque David eo quod confirmasset eum Dominus in regem super Israhel et sublevatum esset regnum suum super populum eius Israhel
1CHR|14|3|accepit quoque David alias uxores in Hierusalem genuitque filios et filias
1CHR|14|4|et haec nomina eorum qui nati sunt ei in Hierusalem Sammu et Sobab Nathan et Salomon
1CHR|14|5|Iebar et Helisu et Eliphaleth
1CHR|14|6|Noga quoque et Napheg et Iaphiae
1CHR|14|7|Elisama et Baliada et Eliphaleth
1CHR|14|8|audientes autem Philisthim eo quod unctus esset David in regem super universum Israhel ascenderunt omnes ut quaererent eum quod cum audisset David egressus est obviam eis
1CHR|14|9|porro Philisthim venientes diffusi sunt in valle Raphaim
1CHR|14|10|consuluitque David Deum dicens si ascendam ad Philistheos si trades eos in manu mea et dixit ei Dominus ascende et tradam eos in manu tua
1CHR|14|11|cumque illi ascendissent in Baalpharasim percussit eos ibi David et dixit divisit Deus inimicos meos per manum meam sicuti dividuntur aquae et idcirco vocatum est nomen loci illius Baalpharasim
1CHR|14|12|dereliqueruntque ibi deos suos quos David iussit exuri
1CHR|14|13|alia etiam vice Philisthim inruerunt et diffusi sunt in valle
1CHR|14|14|consuluitque rursum David Deum et dixit ei Deus non ascendas post eos recede ab eis et venies contra illos ex adverso pirorum
1CHR|14|15|cumque audieris sonitum gradientis in cacumine pirorum tunc egredieris ad bellum egressus est enim Deus ante te ut percutiat castra Philisthim
1CHR|14|16|fecit ergo David sicut praeceperat ei Deus et percussit castra Philisthinorum de Gabaon usque Gazera
1CHR|14|17|divulgatumque est nomen David in universis regionibus et Dominus dedit pavorem eius super omnes gentes
1CHR|15|1|fecit quoque sibi domos in civitate David et aedificavit locum arcae Dei tetenditque ei tabernaculum
1CHR|15|2|tunc dixit David inlicitum est ut a quocumque portetur arca Dei nisi a Levitis quos elegit Dominus ad portandum eam et ad ministrandum sibi usque in aeternum
1CHR|15|3|congregavitque universum Israhel in Hierusalem ut adferretur arca Dei in locum suum quem praeparaverat ei
1CHR|15|4|necnon et filios Aaron et Levitas
1CHR|15|5|de filiis Caath Urihel princeps fuit et fratres eius centum viginti
1CHR|15|6|de filiis Merari Asaia princeps et fratres eius ducenti viginti
1CHR|15|7|de filiis Gersom Iohel princeps et fratres eius centum triginta
1CHR|15|8|de filiis Elisaphan Semeias princeps et fratres eius ducenti
1CHR|15|9|de filiis Hebron Elihel princeps et fratres eius octoginta
1CHR|15|10|de filiis Ozihel Aminadab princeps et fratres eius centum duodecim
1CHR|15|11|vocavitque David Sadoc et Abiathar sacerdotes et Levitas Urihel Asaiam Iohel Semeiam Elihel et Aminadab
1CHR|15|12|et dixit ad eos vos qui estis principes familiarum leviticarum sanctificamini cum fratribus vestris et adferte arcam Domini Dei Israhel ad locum qui ei praeparatus est
1CHR|15|13|ne ut a principio quia non eratis praesentes percussit nos Dominus sic et nunc fiat inlicitum quid nobis agentibus
1CHR|15|14|sanctificati sunt ergo sacerdotes et Levitae ut portarent arcam Domini Dei Israhel
1CHR|15|15|et tulerunt filii Levi arcam Dei sicut praeceperat Moses iuxta verbum Domini umeris suis in vectibus
1CHR|15|16|dixit quoque David principibus Levitarum ut constituerent de fratribus suis cantores in organis musicorum nablis videlicet et lyris et cymbalis ut resonaret in excelsum sonitus laetitiae
1CHR|15|17|constitueruntque Levitas Heman filium Iohel et de fratribus eius Asaph filium Barachiae de filiis vero Merari fratribus eorum Ethan filium Casaiae
1CHR|15|18|et cum eis fratres eorum in secundo ordine Zacchariam et Ben et Iazihel et Semiramoth et Iahihel et Ani Eliab et Banaiam et Maasiam et Matthathiam et Eliphalu et Macheniam et Obededom et Ieihel ianitores
1CHR|15|19|porro cantores Heman Asaph et Ethan in cymbalis aeneis concrepantes
1CHR|15|20|Zaccharias autem et Ozihel et Semiramoth et Iahihel et Ani et Eliab et Maasias et Banaias in nablis arcana cantabant
1CHR|15|21|porro Matthathias et Eliphalu et Machenias et Obededom et Ieihel et Ozaziu in citharis pro octava canebant epinikion
1CHR|15|22|Chonenias autem princeps Levitarum prophetiae praeerat ad praecinendam melodiam erat quippe valde sapiens
1CHR|15|23|et Barachias et Helcana ianitores arcae
1CHR|15|24|porro Sebenias et Iosaphat et Nathanahel et Amasai et Zaccharias et Banaias et Eliezer sacerdotes clangebant tubis coram arca Dei et Obededom et Ahias erant ianitores arcae
1CHR|15|25|igitur David et maiores natu Israhel et tribuni ierunt ad deportandam arcam foederis Domini de domo Obededom cum laetitia
1CHR|15|26|cumque adiuvisset Deus Levitas qui portabant arcam foederis Domini immolabantur septem tauri et septem arietes
1CHR|15|27|porro David erat indutus stola byssina et universi Levitae qui portabant arcam cantoresque et Chonenias princeps prophetiae inter cantores David autem indutus erat etiam ephod lineo
1CHR|15|28|universusque Israhel deducebant arcam foederis Domini in iubilo et sonitu bucinae et tubis et cymbalis et nablis et citharis concrepantes
1CHR|15|29|cumque pervenisset arca foederis Domini usque ad civitatem David Michol filia Saul prospiciens per fenestram vidit regem David saltantem atque ludentem et despexit eum in corde suo
1CHR|16|1|adtulerunt igitur arcam Dei et constituerunt eam in medio tabernaculi quod tetenderat ei David et obtulerunt holocausta et pacifica coram Deo
1CHR|16|2|cumque conplesset David offerens holocausta et pacifica benedixit populo in nomine Domini
1CHR|16|3|et divisit universis per singulos a viro usque ad mulierem tortam panis et partem assae carnis bubulae et frixam oleo similam
1CHR|16|4|constituitque coram arca Domini de Levitis qui ministrarent et recordarentur operum eius et glorificarent atque laudarent Dominum Deum Israhel
1CHR|16|5|Asaph principem et secundum eius Zacchariam porro Iahihel et Semiramoth et Ieihel et Matthathiam et Eliab et Banaiam et Obededom et Ieihel super organa psalterii et lyras Asaph autem ut cymbalis personaret
1CHR|16|6|Banaiam vero et Azihel sacerdotes canere tuba iugiter coram arca foederis Domini
1CHR|16|7|in illo die fecit David principem ad confitendum Domino Asaph et fratres eius
1CHR|16|8|confitemini Domino invocate nomen eius notas facite in populis adinventiones illius
1CHR|16|9|canite ei et psallite et narrate omnia mirabilia eius
1CHR|16|10|laudate nomen sanctum eius laetetur cor quaerentium Dominum
1CHR|16|11|quaerite Dominum et virtutem eius quaerite faciem eius semper
1CHR|16|12|recordamini mirabilium eius quae fecit signorum illius et iudiciorum oris eius
1CHR|16|13|semen Israhel servi eius filii Iacob electi illius
1CHR|16|14|ipse Dominus Deus noster in universa terra iudicia eius
1CHR|16|15|recordamini in sempiternum pacti eius sermonis quem praecepit in mille generationes
1CHR|16|16|quem pepigit cum Abraham et iuramenti illius cum Isaac
1CHR|16|17|et constituit illud Iacob in praeceptum et Israhel in pactum sempiternum
1CHR|16|18|dicens tibi dabo terram Chanaan funiculum hereditatis vestrae
1CHR|16|19|cum essent pauci numero parvi et coloni eius
1CHR|16|20|et transierunt de gente in gentem et de regno ad populum alterum
1CHR|16|21|non dimisit quemquam calumniari eos sed increpuit pro eis reges
1CHR|16|22|nolite tangere christos meos et in prophetis meis nolite malignari
1CHR|16|23|canite Domino omnis terra adnuntiate ex die in diem salutare eius
1CHR|16|24|narrate in gentibus gloriam eius in cunctis populis mirabilia illius
1CHR|16|25|quia magnus Dominus et laudabilis nimis et horribilis super omnes deos
1CHR|16|26|omnes enim dii populorum idola Dominus autem caelos fecit
1CHR|16|27|confessio et magnificentia coram eo fortitudo et gaudium in loco eius
1CHR|16|28|adferte Domino familiae populorum adferte Domino gloriam et imperium
1CHR|16|29|date Domino gloriam nomini eius levate sacrificium et venite in conspectu eius et adorate Dominum in decore sancto
1CHR|16|30|commoveatur a facie illius omnis terra ipse enim fundavit orbem inmobilem
1CHR|16|31|laetentur caeli et exultet terra et dicant in nationibus Dominus regnavit
1CHR|16|32|tonet mare et plenitudo eius exultent agri et omnia quae in eis sunt
1CHR|16|33|tunc laudabunt ligna saltus coram Domino quia venit iudicare terram
1CHR|16|34|confitemini Domino quoniam bonus quoniam in aeternum misericordia eius
1CHR|16|35|et dicite salva nos Deus salvator noster et congrega nos et erue de gentibus ut confiteamur nomini sancto tuo et exultemus in carminibus tuis
1CHR|16|36|benedictus Dominus Deus Israhel ab aeterno usque in aeternum et dicat omnis populus amen et hymnus Domino
1CHR|16|37|dereliquit itaque ibi coram arca foederis Domini Asaph et fratres eius ut ministrarent in conspectu arcae iugiter per singulos dies et vices suas
1CHR|16|38|porro Obededom et fratres eius sexaginta octo et Obededom filium Idithun et Osa constituit ianitores
1CHR|16|39|Sadoc autem sacerdotem et fratres illius sacerdotes coram tabernaculo Domini in excelso quod erat in Gabaon
1CHR|16|40|ut offerrent holocausta Domino super altare holocaustomatis iugiter mane et vespere iuxta omnia quae scripta sunt in lege Domini quam praecepit Israheli
1CHR|16|41|et post eum Heman et Idithun et reliquos electos unumquemque vocabulo suo ad confitendum Domino quoniam in aeternum misericordia eius
1CHR|16|42|Heman quoque et Idithun canentes tuba et quatientes cymbala et omnia musicorum organa ad canendum Deo filios autem Idithun fecit esse portarios
1CHR|16|43|reversusque est omnis populus in domum suam et David ut benediceret etiam domui suae
1CHR|17|1|cum autem habitaret David in domo sua dixit ad Nathan prophetam ecce ego habito in domo cedrina arca autem foederis Domini sub pellibus est
1CHR|17|2|et ait Nathan ad David omnia quae in corde tuo sunt fac Deus enim tecum est
1CHR|17|3|igitur nocte illa factus est sermo Dei ad Nathan dicens
1CHR|17|4|vade et loquere David servo meo haec dicit Dominus non aedificabis tu mihi domum ad habitandum
1CHR|17|5|neque enim mansi in domo ex eo tempore quo eduxi Israhel usque ad hanc diem sed fui semper mutans loca tabernaculi et in tentorio
1CHR|17|6|manens cum omni Israhel numquid locutus sum saltim uni iudicum Israhel quibus praeceperam ut pascerent populum meum et dixi quare non aedificastis mihi domum cedrinam
1CHR|17|7|nunc itaque sic loqueris ad servum meum David haec dicit Dominus exercituum ego tuli te cum in pascuis sequereris gregem ut esses dux populi mei Israhel
1CHR|17|8|et fui tecum quocumque perrexisti et interfeci omnes inimicos tuos coram te fecique tibi nomen quasi unius magnorum qui celebrantur in terra
1CHR|17|9|et dedi locum populo meo Israhel plantabitur et habitabit in eo et ultra non commovebitur nec filii iniquitatis adterent eos sicut a principio
1CHR|17|10|ex diebus quibus dedi iudices populo meo Israhel et humiliavi universos inimicos tuos adnuntio ergo tibi quod aedificaturus sit domum tibi Dominus
1CHR|17|11|cumque impleveris dies tuos ut vadas ad patres tuos suscitabo semen tuum post te quod erit de filiis tuis et stabiliam regnum eius
1CHR|17|12|ipse aedificabit mihi domum et firmabo solium eius usque in aeternum
1CHR|17|13|ego ero ei in patrem et ipse erit mihi in filium et misericordiam meam non auferam ab eo sicut abstuli ab eo qui ante te fuit
1CHR|17|14|et statuam eum in domo mea et in regno meo usque in sempiternum et thronus eius erit firmissimus in perpetuum
1CHR|17|15|iuxta omnia verba haec et iuxta universam visionem istam sic locutus est Nathan ad David
1CHR|17|16|cumque venisset rex David et sedisset coram Domino dixit quis ego sum Domine Deus et quae domus mea ut praestares mihi talia
1CHR|17|17|sed et hoc parum visum est in conspectu tuo ideoque locutus es super domum servi tui etiam in futurum et fecisti me spectabilem super omnes homines Domine Deus meus
1CHR|17|18|quid ultra addere potest David cum ita glorificaveris servum tuum et cognoveris eum
1CHR|17|19|Domine propter famulum tuum iuxta cor tuum fecisti omnem magnificentiam hanc et nota esse voluisti universa magnalia
1CHR|17|20|Domine non est similis tui et non est alius deus absque te ex omnibus quos audivimus auribus nostris
1CHR|17|21|quis autem est alius ut populus tuus Israhel gens una in terra ad quam perrexit Deus ut liberaret et faceret populum sibi et magnitudine sua atque terroribus eiceret nationes a facie eius quem de Aegypto liberarat
1CHR|17|22|et posuisti populum tuum Israhel tibi in populum usque in aeternum et tu Domine factus es Deus eius
1CHR|17|23|nunc igitur Domine sermo quem locutus es famulo tuo et super domum eius confirmetur in perpetuum et fac sicut locutus es
1CHR|17|24|permaneatque et magnificetur nomen tuum usque in sempiternum et dicatur Dominus exercituum Deus Israhel et domus David servi eius permanens coram eo
1CHR|17|25|tu enim Domine Deus meus revelasti auriculam servi tui ut aedificares ei domum et idcirco invenit servus tuus fiduciam ut oret coram te
1CHR|17|26|nunc ergo Domine tu es Deus et locutus es ad servum tuum tanta beneficia
1CHR|17|27|et coepisti benedicere domui servi tui ut sit semper coram te te enim Domine benedicente benedicta erit in perpetuum
1CHR|18|1|factum est autem post haec ut percuteret David Philisthim et humiliaret eos et tolleret Geth et filias eius de manu Philisthim
1CHR|18|2|percuteretque Moab et fierent Moabitae servi David offerentes ei munera
1CHR|18|3|eo tempore percussit David etiam Adadezer regem Suba regionis Emath quando perrexit ut dilataret imperium suum usque ad flumen Eufraten
1CHR|18|4|cepit ergo David mille quadrigas eius et septem milia equites ac viginti milia virorum peditum subnervavitque omnes equos curruum exceptis centum quadrigis quas reservavit sibi
1CHR|18|5|supervenit autem et Syrus damascenus ut auxilium praeberet Adadezer regi Suba sed et huius percussit David viginti duo milia virorum
1CHR|18|6|et posuit milites in Damasco ut Syria quoque serviret sibi et offerret munera adiuvitque eum Dominus in cunctis ad quae perrexerat
1CHR|18|7|tulit quoque David faretras aureas quas habuerant servi Adadezer et adtulit eas in Hierusalem
1CHR|18|8|necnon de Thebath et Chun urbibus Adadezer aeris plurimum de quo fecit Salomon mare aeneum et columnas et vasa aenea
1CHR|18|9|quod cum audisset Thou rex Emath percussisse videlicet David omnem exercitum Adadezer regis Suba
1CHR|18|10|misit Aduram filium suum ad regem David ut postularet ab eo pacem et congratularetur ei eo quod expugnasset et percussisset Adadezer adversarius quippe Thou erat Adadezer
1CHR|18|11|sed et omnia vasa aurea et argentea et aenea consecravit rex David Domino cum argento et auro quod tulerat ex universis gentibus tam de Idumea et Moab et filiis Ammon quam de Philisthim et Amalech
1CHR|18|12|Abisai vero filius Sarviae percussit Edom in valle Salinarum decem et octo milia
1CHR|18|13|et constituit in Edom praesidium ut serviret Idumea David salvavitque Dominus David in cunctis ad quae perrexerat
1CHR|18|14|regnavit ergo David super universum Israhel et faciebat iudicium atque iustitiam cuncto populo suo
1CHR|18|15|porro Ioab filius Sarviae erat super exercitum et Iosaphat filius Ahilud a commentariis
1CHR|18|16|Sadoc autem filius Ahitob et Ahimelech filius Abiathar sacerdotes et Susa scriba
1CHR|18|17|Banaias vero filius Ioiada super legiones Cherethi et Felethi porro filii David primi ad manum regis
1CHR|19|1|accidit autem ut moreretur Naas rex filiorum Ammon et regnaret filius eius pro eo
1CHR|19|2|dixitque David faciam misericordiam cum Hanon filio Naas praestitit enim pater eius mihi gratiam misitque David nuntios ad consolandum eum super morte patris sui qui cum pervenissent in terram filiorum Ammon ut consolarentur Hanon
1CHR|19|3|dixerunt principes filiorum Ammon ad Hanon tu forsitan putas quod David honoris causa in patrem tuum miserit qui consolentur te nec animadvertis quod ut explorent et investigent et scrutentur terram tuam venerint ad te servi eius
1CHR|19|4|igitur Hanon pueros David decalvavit et rasit et praecidit tunicas eorum a natibus usque ad pedes et dimisit eos
1CHR|19|5|qui cum abissent et hoc mandassent David misit in occursum eorum grandem enim contumeliam sustinuerant et praecepit ut manerent in Hiericho donec cresceret barba eorum et tunc reverterentur
1CHR|19|6|videntes autem filii Ammon quod iniuriam fecissent David tam Hanon quam reliquus populus miserunt mille talenta argenti ut conducerent sibi de Mesopotamia et de Syria Macha et de Suba currus et equites
1CHR|19|7|conduxeruntque triginta duo milia curruum et regem Macha cum populo eius qui cum venissent castrametati sunt e regione Medaba filii quoque Ammon congregati de urbibus suis venerunt ad bellum
1CHR|19|8|quod cum audisset David misit Ioab et omnem exercitum virorum fortium
1CHR|19|9|egressique filii Ammon direxerunt aciem iuxta portam civitatis reges autem qui ad auxilium venerant separatim in agro steterunt
1CHR|19|10|igitur Ioab intellegens bellum et ex adverso et post tergum contra se fieri elegit viros fortissimos de universo Israhel et perrexit contra Syrum
1CHR|19|11|reliquam autem partem populi dedit sub manu Abisai fratris sui et perrexerunt contra filios Ammon
1CHR|19|12|dixitque si vicerit me Syrus auxilio eris mihi sin autem superaverint te filii Ammon ero tibi in praesidium
1CHR|19|13|confortare et agamus viriliter pro populo nostro et pro urbibus Dei nostri Dominus autem quod in conspectu suo bonum est faciet
1CHR|19|14|perrexit ergo Ioab et populus qui cum eo erat contra Syrum ad proelium et fugavit eos
1CHR|19|15|porro filii Ammon videntes quod fugisset Syrus ipsi quoque fugerunt Abisai fratrem eius et ingressi sunt civitatem reversusque est etiam Ioab in Hierusalem
1CHR|19|16|videns autem Syrus quod cecidisset coram Israhel misit nuntios et adduxit Syrum qui erat trans Fluvium Sophach autem princeps militiae Adadezer erat dux eorum
1CHR|19|17|quod cum nuntiatum esset David congregavit universum Israhel et transivit Iordanem inruitque in eos et direxit ex adverso aciem illis contra pugnantibus
1CHR|19|18|fugit autem Syrus Israhel et interfecit David de Syris septem milia curruum et quadraginta milia peditum et Sophach exercitus principem
1CHR|19|19|videntes autem servi Adadezer se ab Israhel esse superatos transfugerunt ad David et servierunt ei noluitque ultra Syria auxilium praebere filiis Ammon
1CHR|20|1|factum est autem post anni circulum eo tempore quo solent reges ad bella procedere congregavit Ioab exercitum et robur militiae et vastavit terram filiorum Ammon perrexitque et obsedit Rabba porro David manebat in Hierusalem quando Ioab percussit Rabba et destruxit eam
1CHR|20|2|tulit autem David coronam Melchom de capite eius et invenit in ea auri pondo talentum et pretiosissimas gemmas fecitque sibi inde diadema manubias quoque urbis plurimas tulit
1CHR|20|3|populum autem qui erat in ea eduxit et fecit super eos tribulas et trahas et ferrata carpenta transire ita ut dissicarentur et contererentur sic fecit David cunctis urbibus filiorum Ammon et reversus est cum omni populo suo in Hierusalem
1CHR|20|4|post haec initum est bellum in Gazer adversus Philistheos in quo percussit Sobbochai Usathites Saphai de genere Raphaim et humiliavit eos
1CHR|20|5|aliud quoque bellum gestum est adversum Philistheos in quo percussit Adeodatus filius Saltus Lehemites fratrem Goliath Getthei cuius hastae lignum erat quasi liciatorium texentium
1CHR|20|6|sed et aliud bellum accidit in Geth in quo fuit homo longissimus habens digitos senos id est simul viginti quattuor qui et ipse de Rapha fuerat stirpe generatus
1CHR|20|7|hic blasphemavit Israhel et percussit eum Ionathan filius Sammaa fratris David hii sunt filii Rapha in Geth qui ceciderunt in manu David et servorum eius
1CHR|21|1|consurrexit autem Satan contra Israhel et incitavit David ut numeraret Israhel
1CHR|21|2|dixitque David ad Ioab et ad principes populi ite et numerate Israhel a Bersabee usque Dan et adferte mihi numerum ut sciam
1CHR|21|3|responditque Ioab augeat Dominus populum suum centuplum quam sunt nonne domine mi rex omnes servi tui sunt quare hoc quaerit dominus meus quod in peccatum reputetur Israheli
1CHR|21|4|sed sermo regis magis praevaluit egressusque est Ioab et circuivit universum Israhel et reversus est Hierusalem
1CHR|21|5|deditque David numerum eorum quos circumierat et inventus est omnis Israhel numerus mille milia et centum milia virorum educentium gladium de Iuda autem trecenta septuaginta milia bellatorum
1CHR|21|6|nam Levi et Beniamin non numeravit eo quod invitus exsequeretur regis imperium
1CHR|21|7|displicuit autem Deo quod iussum erat et percussit Israhel
1CHR|21|8|dixitque David ad Deum peccavi nimis ut hoc facerem obsecro aufer iniquitatem servi tui quia insipienter egi
1CHR|21|9|et locutus est Dominus ad Gad videntem David dicens
1CHR|21|10|vade et loquere ad David et dic haec dicit Dominus trium tibi optionem do unum quod volueris elige et faciam tibi
1CHR|21|11|cumque venisset Gad ad David dixit ei haec dicit Dominus elige quod volueris
1CHR|21|12|aut tribus annis pestilentiam aut tribus mensibus fugere te hostes tuos et gladium eorum non posse evadere aut tribus diebus gladium Domini et mortem versari in terra et angelum Domini interficere in universis finibus Israhel nunc igitur vide quid respondeam ei qui misit me
1CHR|21|13|et dixit David ad Gad ex omni parte me angustiae premunt sed melius mihi est ut incidam in manus Domini quia multae sunt miserationes eius quam in manus hominum
1CHR|21|14|misit ergo Dominus pestilentiam in Israhel et ceciderunt de Israhel septuaginta milia virorum
1CHR|21|15|misit quoque angelum in Hierusalem ut percuteret eam cumque percuteretur vidit Dominus et misertus est super magnitudinem mali et imperavit angelo qui percutiebat sufficit iam cesset manus tua porro angelus Domini stabat iuxta aream Ornan Iebusei
1CHR|21|16|levansque David oculos suos vidit angelum Domini stantem inter terram et caelum et evaginatum gladium in manu eius et versum contra Hierusalem et ceciderunt tam ipse quam maiores natu vestiti ciliciis et proni in terram
1CHR|21|17|dixitque David ad Deum nonne ego sum qui iussi ut numeraretur populus ego qui peccavi ego qui malum feci iste grex quid commeruit Domine Deus meus vertatur obsecro manus tua in me et in domum patris mei populus autem tuus non percutiatur
1CHR|21|18|angelus autem Domini praecepit Gad ut diceret David et ascenderet extrueretque altare Domino Deo in area Ornan Iebusei
1CHR|21|19|ascendit ergo David iuxta sermonem Gad quem locutus fuerat ex nomine Domini
1CHR|21|20|porro Ornan cum suspexisset et vidisset angelum quattuorque filii eius cum eo absconderunt se nam eo tempore terebat in area triticum
1CHR|21|21|igitur cum venisset David ad Ornan conspexit eum Ornan et processit ei obviam de area et adoravit illum pronus in terram
1CHR|21|22|dixitque ei David da mihi locum areae tuae ut aedificem in ea altare Domini ita ut quantum valet argenti accipias et cesset plaga a populo
1CHR|21|23|dixit autem Ornan ad David tolle et faciat dominus meus rex quodcumque ei placet sed et boves do in holocaustum et tribulas in ligna et triticum in sacrificium omnia libens praebeo
1CHR|21|24|dixitque ei rex David nequaquam ita fiet sed argentum dabo quantum valet neque enim tibi auferre debeo et sic offerre Domino holocausta gratuita
1CHR|21|25|dedit ergo David Ornan pro loco siclos auri iustissimi ponderis sescentos
1CHR|21|26|et aedificavit ibi altare Domino obtulitque holocausta et pacifica et invocavit Dominum et exaudivit eum in igne de caelo super altare holocausti
1CHR|21|27|praecepitque Dominus angelo et convertit gladium suum in vaginam
1CHR|21|28|protinus ergo David videns quod exaudisset eum Dominus in area Ornan Iebusei immolavit ibi victimas
1CHR|21|29|tabernaculum autem Domini quod fecerat Moses in deserto et altare holocaustorum ea tempestate erat in excelso Gabaon
1CHR|21|30|et non praevaluit David ire ad altare ut ibi obsecraret Deum nimio enim fuerat timore perterritus videns gladium angeli Domini
1CHR|22|1|dixitque David haec est domus Dei et hoc altare in holocaustum Israhel
1CHR|22|2|et praecepit ut congregarentur omnes proselyti de terra Israhel et constituit ex eis latomos ad caedendos lapides et poliendos ut aedificaretur domus Dei
1CHR|22|3|ferrum quoque plurimum ad clavos ianuarum et ad commissuras atque iuncturas praeparavit David et aeris pondus innumerabile
1CHR|22|4|ligna quoque cedrina non poterant aestimari quae Sidonii et Tyrii deportaverant ad David
1CHR|22|5|et dixit David Salomon filius meus puer parvulus est et delicatus domus autem quam aedificari volo Domino talis esse debet ut in cunctis regionibus nominetur praeparabo ergo ei necessaria et ob hanc causam ante mortem suam omnes paravit inpensas
1CHR|22|6|vocavitque Salomonem filium suum et praecepit ei ut aedificaret domum Domino Deo Israhel
1CHR|22|7|dixitque David ad Salomonem fili mi voluntatis meae fuit ut aedificarem domum nomini Domini Dei mei
1CHR|22|8|sed factus est ad me sermo Domini dicens multum sanguinem effudisti et plurima bella bellasti non poteris aedificare domum nomini meo tanto effuso sanguine coram me
1CHR|22|9|filius qui nascetur tibi et erit vir quietissimus faciam enim eum requiescere ab omnibus inimicis suis per circuitum et ob hanc causam pacificus vocabitur et pacem et otium dabo in Israhel cunctis diebus eius
1CHR|22|10|ipse aedificabit domum nomini meo et ipse erit mihi in filium et ego ero ei in patrem firmaboque solium regni eius super Israhel in aeternum
1CHR|22|11|nunc ergo fili mi sit Dominus tecum et prosperare et aedifica domum Domino Deo tuo sicut locutus est de te
1CHR|22|12|det quoque tibi Dominus prudentiam et sensum ut regere possis Israhel et custodire legem Domini Dei tui
1CHR|22|13|tunc enim proficere poteris si custodieris mandata et iudicia quae praecepit Dominus Mosi ut doceret Israhel confortare viriliter age ne timeas neque paveas
1CHR|22|14|ecce ego in paupertatula mea praeparavi inpensas domus Domini auri talenta centum milia et argenti mille milia talentorum aeris vero et ferri non est pondus vincitur enim numerus magnitudine ligna et lapides praeparavi ad universa inpendia
1CHR|22|15|habes quoque plurimos artifices latomos et cementarios artificesque lignorum et omnium artium ad faciendum opus prudentissimos
1CHR|22|16|in auro et argento aere et ferro cuius non est numerus surge igitur et fac et erit Dominus tecum
1CHR|22|17|praecepit quoque David cunctis principibus Israhel ut adiuvarent Salomonem filium suum
1CHR|22|18|cernitis inquiens quod Dominus Deus vester vobiscum sit et dederit vobis requiem per circuitum et tradiderit omnes inimicos in manu vestra et subiecta sit terra coram Domino et coram populo eius
1CHR|22|19|praebete igitur corda vestra et animas vestras ut quaeratis Dominum Deum vestrum et consurgite et aedificate sanctuarium Domino Deo ut introducatur arca foederis Domini et vasa Domino consecrata in domum quae aedificatur nomini Domini
1CHR|23|1|igitur David senex et plenus dierum regem constituit Salomonem filium suum super Israhel
1CHR|23|2|et congregavit omnes principes Israhel et sacerdotes atque Levitas
1CHR|23|3|numeratique sunt Levitae a triginta annis et supra et inventa sunt triginta octo milia virorum
1CHR|23|4|ex his electi sunt et distributi in ministerium domus Domini viginti quattuor milia praepositorum autem et iudicum sex milia
1CHR|23|5|porro quattuor milia ianitores et totidem psaltae canentes Domino in organis quae fecerat ad canendum
1CHR|23|6|et distribuit eos David per vices filiorum Levi Gersom videlicet et Caath et Merari
1CHR|23|7|Gersom Leedan et Semei
1CHR|23|8|filii Leedan princeps Ieihel et Zetham et Iohel tres
1CHR|23|9|filii Semei Salomith et Ozihel et Aran tres isti principes familiarum Leedan
1CHR|23|10|porro filii Semei Ieeth et Ziza et Iaus et Baria isti filii Semei quattuor
1CHR|23|11|erat autem Ieeth prior Ziza secundus porro Iaus et Baria non habuerunt plurimos filios et idcirco in una familia unaque domo conputati sunt
1CHR|23|12|filii Caath Amram et Isaar Hebron et Ozihel quattuor
1CHR|23|13|filii Amram Aaron et Moses separatusque est Aaron ut ministraret in sancto sanctorum ipse et filii eius in sempiternum et adoleret incensum Domino secundum ritum suum ac benediceret nomini eius in perpetuum
1CHR|23|14|Mosi quoque hominis Dei filii adnumerati sunt in tribu Levi
1CHR|23|15|filii Mosi Gersom et Eliezer
1CHR|23|16|filii Gersom Subuhel primus
1CHR|23|17|fuerunt autem filii Eliezer Roobia primus et non erant Eliezer filii alii porro filii Roobia multiplicati sunt nimis
1CHR|23|18|filii Isaar Salumith primus
1CHR|23|19|filii Hebron Ieriau primus Amarias secundus Iazihel tertius Iecmaam quartus
1CHR|23|20|filii Ozihel Micha primus Iesia secundus
1CHR|23|21|filii Merari Mooli et Musi filii Mooli Eleazar et Cis
1CHR|23|22|mortuus est autem Eleazar et non habuit filios sed filias acceperuntque eas filii Cis fratres earum
1CHR|23|23|filii Musi Mooli et Eder et Ierimuth tres
1CHR|23|24|hii filii Levi in cognationibus et familiis suis principes per vices et numerum capitum singulorum qui faciebant opera ministerii domus Domini a viginti annis et supra
1CHR|23|25|dixit enim David requiem dedit Dominus Deus Israhel populo suo et habitationem Hierusalem usque in aeternum
1CHR|23|26|nec erit officii Levitarum ut ultra portent tabernaculum et omnia vasa eius ad ministrandum
1CHR|23|27|iuxta praecepta quoque David novissima supputabitur numerus filiorum Levi a viginti annis et supra
1CHR|23|28|et erunt sub manu filiorum Aaron in cultum domus Domini in vestibulis et in exedris et in loco purificationis et in sanctuario et in universis operibus ministerii templi Domini
1CHR|23|29|sacerdotes autem super panes propositionis et ad similae sacrificium et ad lagana et azyma et sartaginem et ad ferventem similam et super omne pondus atque mensuram
1CHR|23|30|Levitae vero ut stent mane ad confitendum et canendum Domino similiterque ad vesperam
1CHR|23|31|tam in oblatione holocaustorum Domini quam in sabbatis et kalendis et sollemnitatibus reliquis iuxta numerum et caerimonias uniuscuiusque rei iugiter coram Domino
1CHR|23|32|et custodiant observationes tabernaculi foederis et ritum sanctuarii et observationem filiorum Aaron fratrum suorum ut ministrent in domo Domini
1CHR|24|1|porro filiis Aaron hae partitiones erunt filii Aaron Nadab et Abiu et Eleazar et Ithamar
1CHR|24|2|mortui sunt autem Nadab et Abiu ante patrem suum absque liberis sacerdotioque functus est Eleazar et Ithamar
1CHR|24|3|et divisit eos David id est Sadoc de filiis Eleazar et Ahimelech de filiis Ithamar secundum vices suas et ministerium
1CHR|24|4|inventique sunt multo plures filii Eleazar in principibus viris quam filii Ithamar divisit autem eis hoc est filiis Eleazar principes per familias sedecim et filiis Ithamar per familias et domos suas octo
1CHR|24|5|porro divisit utrasque inter se familias sortibus erant enim principes sanctuarii et principes Dei tam de filiis Eleazar quam de filiis Ithamar
1CHR|24|6|descripsitque eos Semeias filius Nathanahel scriba Levites coram rege et principibus et Sadoc sacerdote et Ahimelech filio Abiathar principibus quoque familiarum sacerdotalium et leviticarum unam domum quae ceteris praeerat Eleazar et alteram domum quae sub se habebat ceteros Ithamar
1CHR|24|7|exivit autem sors prima Ioiarib secunda Iedeiae
1CHR|24|8|tertia Arim quarta Seorim
1CHR|24|9|quinta Melchia sexta Maiman
1CHR|24|10|septima Accos octava Abia
1CHR|24|11|nona Hiesu decima Sechenia
1CHR|24|12|undecima Eliasib duodecima Iacim
1CHR|24|13|tertiadecima Oppa quartadecima Isbaal
1CHR|24|14|quintadecima Belga sextadecima Emmer
1CHR|24|15|septimadecima Ezir octavadecima Hapses
1CHR|24|16|nonadecima Phetheia vicesima Iezecel
1CHR|24|17|vicesima prima Iachin vicesima secunda Gamul
1CHR|24|18|vicesima tertia Dalaiau vicesima quarta Mazziau
1CHR|24|19|hae vices eorum secundum ministeria sua ut ingrediantur domum Domini et iuxta ritum suum sub manu Aaron patris eorum sicut praecepit Dominus Deus Israhel
1CHR|24|20|porro filiorum Levi qui reliqui fuerant de filiis Amram erat Subahel et filiis Subahel Iedeia
1CHR|24|21|de filiis quoque Roobiae princeps Iesias
1CHR|24|22|Isaaris vero Salemoth filiusque Salemoth Iaath
1CHR|24|23|filiusque eius Ieriahu Amarias secundus Iazihel tertius Iecmaam quartus
1CHR|24|24|filius Ozihel Micha filius Micha Samir
1CHR|24|25|frater Micha Iesia filiusque Iesiae Zaccharias
1CHR|24|26|filii Merari Mooli et Musi filius Ioziau Benno
1CHR|24|27|filius quoque Merari Oziau et Soem et Zacchur et Hebri
1CHR|24|28|porro Mooli filius Eleazar qui non habebat liberos
1CHR|24|29|filius vero Cis Ierahemel
1CHR|24|30|filii Musi Mooli Eder et Ierimoth isti filii Levi secundum domos familiarum suarum
1CHR|24|31|miseruntque et ipsi sortes contra fratres suos filios Aaron coram David rege et Sadoc et Ahimelech et principibus familiarum sacerdotalium et leviticarum tam maiores quam minores omnes sors aequaliter dividebat
1CHR|25|1|igitur David et magistratus exercitus secreverunt in ministerium filios Asaph et Heman et Idithun qui prophetarent in citharis et psalteriis et cymbalis secundum numerum suum dedicato sibi officio servientes
1CHR|25|2|de filiis Asaph Zacchur et Ioseph et Nathania et Asarela filii Asaph sub manu Asaph prophetantis iuxta regem
1CHR|25|3|porro Idithun filii Idithun Godolias Sori Iesaias et Sabias et Matthathias sex sub manu patris sui Idithun qui in cithara prophetabat super confitentes et laudantes Dominum
1CHR|25|4|Heman quoque filii Heman Bocciau Matthaniau Ozihel Subuhel et Ierimoth Ananias Anani Elietha Geddelthi et Romemthiezer et Iesbacasa Mellothi Othir Mazioth
1CHR|25|5|omnes isti filii Heman videntis regis in sermonibus Dei ut exaltaret cornu deditque Deus Heman filios quattuordecim et filias tres
1CHR|25|6|universi sub manu patris sui ad cantandum in templo Domini distributi erant in cymbalis et psalteriis et citharis in ministeria domus Domini iuxta regem Asaph videlicet et Idithun et Heman
1CHR|25|7|fuit autem numerus eorum cum fratribus suis qui erudiebant canticum Domini cuncti doctores ducenti octoginta octo
1CHR|25|8|miseruntque sortes per vices suas ex aequo tam maior quam minor doctus pariter et indoctus
1CHR|25|9|egressaque est sors prima Ioseph qui erat de Asaph secunda Godoliae ipsi et filiis eius et fratribus duodecim
1CHR|25|10|tertia Zacchur filiis et fratribus eius duodecim
1CHR|25|11|quarta Isari filiis et fratribus eius duodecim
1CHR|25|12|quinta Nathaniae filiis et fratribus eius duodecim
1CHR|25|13|sexta Bocciau filiis et fratribus eius duodecim
1CHR|25|14|septima Israhela filiis et fratribus eius duodecim
1CHR|25|15|octava Isaiae filiis et fratribus eius duodecim
1CHR|25|16|nona Matthaniae filiis et fratribus eius duodecim
1CHR|25|17|decima Semeiae filiis et fratribus eius duodecim
1CHR|25|18|undecima Ezrahel filiis et fratribus eius duodecim
1CHR|25|19|duodecima Asabiae filiis et fratribus eius duodecim
1CHR|25|20|tertiadecima Subahel filiis et fratribus eius duodecim
1CHR|25|21|quartadecima Matthathiae filiis et fratribus eius duodecim
1CHR|25|22|quintadecima Ierimoth filiis et fratribus eius duodecim
1CHR|25|23|sextadecima Ananiae filiis et fratribus eius duodecim
1CHR|25|24|septimadecima Iesbocasae filiis et fratribus eius duodecim
1CHR|25|25|octavadecima Anani filiis et fratribus eius duodecim
1CHR|25|26|nonadecima Mellothi filiis et fratribus eius duodecim
1CHR|25|27|vicesima Eliatha filiis et fratribus eius duodecim
1CHR|25|28|vicesima prima Othir filiis et fratribus eius duodecim
1CHR|25|29|vicesima secunda Godollathi filiis et fratribus eius duodecim
1CHR|25|30|vicesima tertia Maziuth filiis et fratribus eius duodecim
1CHR|25|31|vicesima quarta Romamthiezer filiis et fratribus eius duodecim
1CHR|26|1|divisiones autem ianitorum de Coritis Mesellemia filius Core de filiis Asaph
1CHR|26|2|filii Mesellemiae Zaccharias primogenitus Iadihel secundus Zabadias tertius Iathanahel quartus
1CHR|26|3|Ahilam quintus Iohanan sextus Helioenai septimus
1CHR|26|4|filii autem Obededom Semeias primogenitus Iozabad secundus Iohaa tertius Sachar quartus Nathanahel quintus
1CHR|26|5|Amihel sextus Isachar septimus Phollathi octavus quia benedixit illi Dominus
1CHR|26|6|Semeiae autem filio eius nati sunt filii praefecti familiarum suarum erant enim viri fortissimi
1CHR|26|7|filii ergo Semeiae Othni et Raphahel et Obedihel Zabad fratres eius viri fortissimi Heliu quoque et Samachias
1CHR|26|8|omnes hii de filiis Obededom ipsi et filii et fratres eorum fortissimi ad ministrandum sexaginta duo de Obededom
1CHR|26|9|porro Mesellamiae filii et fratres robustissimi decem et octo
1CHR|26|10|de Hosa autem id est de filiis Merari Semri princeps non enim habuerat primogenitum et idcirco posuerat eum pater eius in principem
1CHR|26|11|Helchias secundus Tabelias tertius Zaccharias quartus omnes hii filii et fratres Hosa tredecim
1CHR|26|12|hii divisi sunt in ianitores ut semper principes custodiarum sicut et fratres eorum ministrarent in domo Domini
1CHR|26|13|missae sunt autem sortes ex aequo et parvis et magnis per familias suas in unamquamque portarum
1CHR|26|14|cecidit igitur sors orientalis Selemiae porro Zacchariae filio eius viro prudentissimo et erudito sortito obtigit plaga septentrionalis
1CHR|26|15|Obededom vero et filiis eius ad austrum in qua parte domus erat seniorum concilium
1CHR|26|16|Sepphima et Hosa ad occidentem iuxta portam quae ducit ad viam ascensionis custodia contra custodiam
1CHR|26|17|ad orientem vero Levitae sex et ad aquilonem quattuor per diem atque ad meridiem similiter in die quattuor et ubi erat concilium bini et bini
1CHR|26|18|in cellulis quoque ianitorum ad occidentem quattuor in via binique per cellulas
1CHR|26|19|hae sunt divisiones ianitorum filiorum Core et Merari
1CHR|26|20|porro Achias erat super thesauros domus Dei ac vasa sanctorum
1CHR|26|21|filii Ledan filii Gersonni de Ledan principes familiarum Ledan et Gersonni Ieiheli
1CHR|26|22|filii Ieiheli Zathan et Iohel frater eius super thesauros domus Domini
1CHR|26|23|Amramitis et Isaaritis et Hebronitis et Ozihelitibus
1CHR|26|24|Subahel autem filius Gersom filii Mosi praepositus thesauris
1CHR|26|25|fratres quoque eius Eliezer cuius filius Raabia et huius filius Isaias et huius filius Ioram huius quoque filius Zechri sed et huius filius Selemith
1CHR|26|26|ipse Selemith et fratres eius super thesauros sanctorum quae sanctificavit David rex et principes familiarum et tribuni et centuriones et duces exercitus
1CHR|26|27|de bellis et manubiis proeliorum quae consecraverant ad instaurationem et supellectilem templi Domini
1CHR|26|28|haec autem universa sanctificavit Samuhel videns et Saul filius Cis et Abner filius Ner et Ioab filius Sarviae omnes qui sanctificaverunt ea per manum Salemith et fratrum eius
1CHR|26|29|Saaritis vero praeerat Chonenias et filii eius ad opera forinsecus super Israhel ad docendum et ad iudicandum eos
1CHR|26|30|porro de Hebronitis Asabias et fratres eius viri fortissimi mille septingenti praeerant Israheli trans Iordanem contra occidentem in cunctis operibus Domini et in ministerium regis
1CHR|26|31|Hebronitarum autem princeps fuit Hieria secundum familias et cognationes eorum quadragesimo anno regni David recensiti sunt et inventi viri fortissimi in Iazer Galaad
1CHR|26|32|fratresque eius robustioris aetatis duo milia septingenti principes familiarum praeposuit autem eos David rex Rubenitis et Gadditis et dimidio tribus Manasse in omne ministerium Dei et regis
1CHR|27|1|filii autem Israhel secundum numerum suum principes familiarum tribuni et centuriones et praefecti qui ministrabant regi iuxta turmas suas ingredientes et egredientes per singulos menses in anno viginti quattuor milibus singuli praeerant
1CHR|27|2|primae turmae in primo mense Isboam praeerat filius Zabdihel et sub eo viginti quattuor milia
1CHR|27|3|de filiis Phares princeps cunctorum principum in exercitu mense primo
1CHR|27|4|secundi mensis habebat turmam Dudi Ahohites et post se alterum nomine Macelloth qui regebat partem exercitus viginti quattuor milium
1CHR|27|5|dux quoque turmae tertiae in mense tertio erat Banaias filius Ioiadae sacerdos et in divisione sua viginti quattuor milia
1CHR|27|6|ipse est Banaias fortissimus inter triginta et super triginta praeerat autem turmae ipsius Amizabad filius eius
1CHR|27|7|quartus mense quarto Asahel frater Ioab et Zabadias filius eius post eum et in turma eius viginti quattuor milia
1CHR|27|8|quintus mense quinto princeps Samaoth Iezarites et in turma eius viginti quattuor milia
1CHR|27|9|sextus mense sexto Hira filius Acces Thecuites et in turma eius viginti quattuor milia
1CHR|27|10|septimus mense septimo Helles Phallonites de filiis Ephraim et in turma eius viginti quattuor milia
1CHR|27|11|octavus mense octavo Sobochai Asothites de stirpe Zarai et in turma eius viginti quattuor milia
1CHR|27|12|nonus mense nono Abiezer Anathothites de filiis Iemini et in turma eius viginti quattuor milia
1CHR|27|13|decimus mense decimo Marai et ipse Netophathites de stirpe Zarai et in turma eius viginti quattuor milia
1CHR|27|14|undecimus mense undecimo Banaias Pharathonites de filiis Ephraim et in turma eius viginti quattuor milia
1CHR|27|15|duodecimus mense duodecimo Holdai Netophathites de stirpe Gothonihel et in turma eius viginti quattuor milia
1CHR|27|16|porro tribubus praeerant Israhel Rubenitis dux Eliezer filius Zechri Symeonitis dux Saphatias filius Macha
1CHR|27|17|Levitis Asabias filius Camuhel Aaronitis Sadoc
1CHR|27|18|Iuda Heliu frater David Isachar Amri filius Michahel
1CHR|27|19|Zabulonitis Iesmaias filius Abdiae Nepthalitibus Ierimoth filius Ozihel
1CHR|27|20|filiis Ephraim Osee filius Ozaziu dimidio tribus Manasse Iohel filius Phadiae
1CHR|27|21|et dimidio tribus Manasse in Galaad Iaddo filius Zacchariae Beniamin autem Iasihel filius Abner
1CHR|27|22|Dan vero Ezrihel filius Hieroam hii principes filiorum Israhel
1CHR|27|23|noluit autem David numerare eos a viginti annis inferius quia dixerat Dominus ut multiplicaret Israhel quasi stellas caeli
1CHR|27|24|Ioab filius Sarviae coeperat numerare nec conplevit quia super hoc ira inruerat in Israhel et idcirco numerus eorum qui fuerant recensiti non est relatus in fastos regis David
1CHR|27|25|super thesauros autem regis fuit Azmoth filius Adihel his autem thesauris qui erant in urbibus et in vicis et in turribus praesidebat Ionathan filius Oziae
1CHR|27|26|operi autem rustico et agricolis qui exercebant terram praeerat Ezri filius Chelub
1CHR|27|27|vinearumque cultoribus Semeias Ramathites cellis autem vinariis Zabdias Aphonites
1CHR|27|28|nam super oliveta et ficeta quae erant in campestribus Balanan Gaderites super apothecas autem olei Ioas
1CHR|27|29|porro armentis quae pascebantur in Sarona praepositus fuit Setrai Saronites et super boves in vallibus Saphat filius Adli
1CHR|27|30|super camelos vero Ubil Ismahelites et super asinos Iadias Meronathites
1CHR|27|31|super oves quoque Iaziz Agarenus omnes hii principes substantiae regis David
1CHR|27|32|Ionathan autem patruus David consiliarius vir prudens et litteratus ipse et Iaihel filius Achamoni erant cum filiis regis
1CHR|27|33|Ahitophel etiam consiliarius regis et Husi Arachites amicus regis
1CHR|27|34|post Ahitophel fuit Ioiada filius Banaiae et Abiathar princeps autem exercitus regis erat Ioab
1CHR|28|1|convocavit igitur David omnes principes Israhel duces tribuum et praepositos turmarum qui ministrabant regi tribunos quoque et centuriones et qui praeerant substantiae et possessionibus regis filiosque suos cum eunuchis et potentes et robustissimos quosque in exercitu Hierusalem
1CHR|28|2|cumque surrexisset rex et stetisset ait audite me fratres mei et populus meus cogitavi ut aedificarem domum in qua requiesceret arca foederis Domini et scabillum pedum Dei nostri et ad aedificandum omnia praeparavi
1CHR|28|3|Deus autem dixit mihi non aedificabis domum nomini meo eo quod sis vir bellator et sanguinem fuderis
1CHR|28|4|sed elegit Dominus Deus Israhel me de universa domo patris mei ut essem rex super Israhel in sempiternum de Iuda enim elegit principes porro de domo Iuda domum patris mei et de filiis patris mei placuit ei ut me eligeret regem super cunctum Israhel
1CHR|28|5|sed et de filiis meis filios enim multos dedit mihi Dominus elegit Salomonem filium meum ut sederet in throno regni Domini super Israhel
1CHR|28|6|dixitque mihi Salomon filius tuus aedificabit domum meam et atria mea ipsum enim elegi mihi in filium et ego ero ei in patrem
1CHR|28|7|et firmabo regnum eius usque in aeternum si perseveraverit facere praecepta mea et iudicia sicut et hodie
1CHR|28|8|nunc igitur coram universo coetu Israhel audiente Deo nostro custodite et perquirite cuncta mandata Domini Dei nostri ut possideatis terram bonam et relinquatis eam filiis vestris post vos usque in sempiternum
1CHR|28|9|tu autem Salomon fili mi scito Deum patris tui et servi ei corde perfecto et animo voluntario omnia enim corda scrutatur Dominus et universas mentium cogitationes intellegit si quaesieris eum invenies si autem dereliqueris illum proiciet te in aeternum
1CHR|28|10|nunc ergo quia elegit te Dominus ut aedificares domum sanctuarii confortare et perfice
1CHR|28|11|dedit autem David Salomoni filio suo descriptionem porticus et templi et cellariorum et cenaculi et cubiculorum in adytis et domus propitiationis
1CHR|28|12|necnon et omnium quae cogitaverat atriorum et exedrarum per circuitum in thesauros domus Domini et in thesauros sanctorum
1CHR|28|13|divisionumque sacerdotalium et leviticarum in omnia opera domus Domini et in universa vasa ministerii templi Domini
1CHR|28|14|aurum in pondere per singula vasa ministerii argenti quoque pondus pro vasorum ad opera diversitate
1CHR|28|15|sed et ad candelabra aurea et ad lucernas eorum aurum pro mensura uniuscuiusque candelabri et lucernarum similiter et in candelabris argenteis et in lucernis eorum pro diversitate mensurae pondus argenti tradidit
1CHR|28|16|aurum quoque dedit in mensas propositionis pro diversitate mensarum similiter et argentum in alias mensas argenteas
1CHR|28|17|ad fuscinulas quoque et fialas et turibula ex auro purissimo et leunculos aureos pro qualitate mensurae pondus distribuit in leunculum et leunculum similiter et in leones argenteos diversum argenti pondus separavit
1CHR|28|18|altari autem in quo adoletur incensum aurum purissimum dedit ut ex ipso fieret similitudo quadrigae cherubin extendentium alas et velantium arcam foederis Domini
1CHR|28|19|omnia inquit venerunt scripta manu Domini ad me ut intellegerem universa opera exemplaris
1CHR|28|20|dixit quoque David Salomoni filio suo viriliter age et confortare et fac ne timeas et ne paveas Dominus enim Deus meus tecum erit et non dimittet te nec derelinquet donec perficias omne opus ministerii domus Domini
1CHR|28|21|ecce divisiones sacerdotum et Levitarum in omne ministerium domus Domini adsistunt tibi et parati sunt et noverunt tam principes quam populus facere omnia praecepta tua
1CHR|29|1|locutusque est David rex ad omnem ecclesiam Salomonem filium meum unum elegit Deus adhuc puerum et tenellum opus autem grande est neque enim homini praeparatur habitatio sed Deo
1CHR|29|2|ego autem totis viribus meis praeparavi inpensas domus Dei mei aurum ad vasa aurea et argentum in argentea aes in aenea ferrum in ferrea lignum ad lignea lapides onychinos et quasi stibinos et diversorum colorum omnem pretiosum lapidem et marmor parium abundantissime
1CHR|29|3|et super haec quae obtuli in domum Dei mei de peculio meo aurum et argentum do in templum Dei mei exceptis his quae paravi in aedem sanctam
1CHR|29|4|tria milia talenta auri de auro Ophir et septem milia talentorum argenti probatissimi ad deaurandos parietes templi
1CHR|29|5|ut ubicumque opus est aurum de auro et ubicumque opus est argentum argenti opera fiant per manus artificum et si quis sponte offert impleat manum suam hodie et offerat quod voluerit Domino
1CHR|29|6|polliciti sunt itaque principes familiarum et proceres tribuum Israhel tribuni quoque et centuriones et principes possessionum regis
1CHR|29|7|dederuntque in opera domus Dei auri talenta quinque milia et solidos decem milia argenti talenta decem milia et aeris talenta decem et octo milia ferri quoque centum milia talentorum
1CHR|29|8|et apud quemcumque inventi sunt lapides dederunt in thesaurum domus Domini per manum Ieihel Gersonitis
1CHR|29|9|laetatusque est populus cum vota sponte promitterent quia corde toto offerebant ea Domino sed et David rex laetatus est gaudio magno
1CHR|29|10|et benedixit Domino coram universa multitudine et ait benedictus es Domine Deus Israhel patris nostri ab aeterno in aeternum
1CHR|29|11|tua est Domine magnificentia et potentia et gloria atque victoria et tibi laus cuncta enim quae in caelo sunt et in terra tua sunt tuum Domine regnum et tu es super omnes principes
1CHR|29|12|tuae divitiae et tua est gloria tu dominaris omnium in manu tua virtus et potentia in manu tua magnitudo et imperium omnium
1CHR|29|13|nunc igitur Deus noster confitemur tibi et laudamus nomen tuum inclitum
1CHR|29|14|quis ego et quis populus meus ut possimus haec tibi universa promittere tua sunt omnia et quae de manu tua accepimus dedimus tibi
1CHR|29|15|peregrini enim sumus coram te et advenae sicut omnes patres nostri dies nostri quasi umbra super terram et nulla est mora
1CHR|29|16|Domine Deus noster omnis haec copia quam paravimus ut aedificaretur domus nomini sancto tuo de manu tua est et tua sunt omnia
1CHR|29|17|scio Deus meus quod probes corda et simplicitatem diligas unde et ego in simplicitate cordis mei laetus obtuli universa haec et populum tuum qui hic reppertus est vidi cum ingenti gaudio tibi offerre donaria
1CHR|29|18|Domine Deus Abraham et Isaac et Israhel patrum nostrorum custodi in aeternum hanc voluntatem cordis eorum et semper in venerationem tui mens ista permaneat
1CHR|29|19|Salomoni quoque filio meo da cor perfectum ut custodiat mandata tua testimonia tua caerimonias tuas et faciat universa et aedificet aedem cuius inpensas paravi
1CHR|29|20|praecepit autem David universae ecclesiae benedicite Domino Deo nostro et benedixit omnis ecclesia Domino Deo patrum suorum et inclinaverunt se et adoraverunt Deum et deinde regem
1CHR|29|21|immolaveruntque victimas Domino et obtulerunt holocausta die sequenti tauros mille arietes mille agnos mille cum libaminibus suis et universo ritu abundantissime in omnem Israhel
1CHR|29|22|et comederunt et biberunt coram Domino in die illo cum grandi laetitia et unxerunt secundo Salomonem filium David unxerunt autem Domino in principem et Sadoc in pontificem
1CHR|29|23|seditque Salomon super solium Domini in regem pro David patre suo et cunctis placuit et paruit illi omnis Israhel
1CHR|29|24|sed et universi principes et potentes et cuncti filii regis David dederunt manum et subiecti fuerunt Salomoni regi
1CHR|29|25|magnificavit ergo Dominus Salomonem super omnem Israhel et dedit illi gloriam regni qualem nullus habuit ante eum rex Israhel
1CHR|29|26|igitur David filius Isai regnavit super universum Israhel
1CHR|29|27|et dies quibus regnavit super Israhel fuerunt quadraginta anni in Hebron regnavit septem annis et in Hierusalem triginta tribus
1CHR|29|28|et mortuus est in senectute bona plenus dierum et divitiis et gloria regnavitque Salomon filius eius pro eo
1CHR|29|29|gesta autem David regis priora et novissima scripta sunt in libro Samuhel videntis et in libro Nathan prophetae atque in volumine Gad videntis
1CHR|29|30|universique regni eius et fortitudinis et temporum quae transierunt sub eo sive in Israhel sive in cunctis regnis terrarum
2CHR|1|1|confortatus est ergo Salomon filius David in regno suo et Dominus erat cum eo et magnificavit eum in excelsum
2CHR|1|2|praecepitque Salomon universo Israheli tribunis et centurionibus et ducibus et iudicibus omnis Israhel et principibus familiarum
2CHR|1|3|et abiit cum universa multitudine in excelsum Gabaon ubi erat tabernaculum foederis Dei quod fecit Moses famulus Dei in solitudine
2CHR|1|4|arcam autem Dei adduxerat David de Cariathiarim in locum quem paraverat ei et ubi fixerat illi tabernaculum hoc est in Hierusalem
2CHR|1|5|altare quoque aeneum quod fabricatus fuerat Beselehel filius Uri filii Ur ibi erat coram tabernaculo Domini quod et requisivit Salomon et omnis ecclesia
2CHR|1|6|ascenditque Salomon ad altare aeneum coram tabernaculo foederis Domini et obtulit in eo mille hostias
2CHR|1|7|ecce autem in ipsa nocte apparuit ei Deus dicens postula quod vis ut dem tibi
2CHR|1|8|dixitque Salomon Deo tu fecisti cum David patre meo misericordiam magnam et constituisti me regem pro eo
2CHR|1|9|nunc igitur Domine Deus impleatur sermo tuus quem pollicitus es David patri meo tu enim fecisti me regem super populum tuum multum qui tam innumerabilis est quam pulvis terrae
2CHR|1|10|da mihi sapientiam et intellegentiam ut egrediar coram populo tuo et ingrediar quis enim potest hunc populum tuum digne qui tam grandis est iudicare
2CHR|1|11|dixit autem Deus ad Salomonem quia hoc magis placuit cordi tuo et non postulasti divitias et substantiam et gloriam neque animas eorum qui te oderunt sed nec dies vitae plurimos petisti autem sapientiam et scientiam ut iudicare possis populum meum super quem constitui te regem
2CHR|1|12|sapientia et scientia data sunt tibi divitias autem et substantiam et gloriam dabo tibi ita ut nullus in regibus nec ante te nec post te fuerit similis tui
2CHR|1|13|venit ergo Salomon ab excelso Gabaon in Hierusalem coram tabernaculo foederis et regnavit super Israhel
2CHR|1|14|congregavitque sibi currus et equites et facti sunt ei mille quadringenti currus et duodecim milia equitum et fecit eos esse in urbibus quadrigarum et cum rege in Hierusalem
2CHR|1|15|praebuitque rex argentum et aurum in Hierusalem quasi lapides et cedros quasi sycomoros quae nascuntur in campestribus multitudine magna
2CHR|1|16|adducebantur autem ei et equi de Aegypto et de Coa a negotiatoribus regis qui ibant et coemebant pretio
2CHR|1|17|quadrigam equorum sescentis argenteis et equum centum quinquaginta similiter de universis regnis Cettheorum et a regibus Syriae emptio celebrabatur
2CHR|2|1|decrevit autem Salomon aedificare domum nomini Domini et palatium sibi
2CHR|2|2|et numeravit septuaginta milia virorum portantium umeris et octoginta milia qui caederent lapides in montibus praepositosque eorum tria milia sescentos
2CHR|2|3|misit quoque ad Hiram regem Tyri dicens sicut egisti cum David patre meo et misisti ei ligna cedrina ut aedificaret sibi domum in qua et habitavit
2CHR|2|4|sic fac mecum ut aedificem domum nomini Domini Dei mei et consecrem eam ad adolendum incensum coram illo et fumiganda aromata et ad propositionem panum sempiternam et holocaustomata mane et vespere sabbatis quoque et neomeniis et sollemnitatibus Domini Dei nostri in sempiternum quae mandata sunt Israheli
2CHR|2|5|domus autem quam aedificare cupio magna est magnus est enim Deus noster super omnes deos
2CHR|2|6|quis ergo poterit praevalere ut aedificet ei dignam domum si caelum et caeli caelorum capere eum non queunt quantus ego sum ut possim ei aedificare domum sed ad hoc tantum ut adoleatur incensum coram illo
2CHR|2|7|mitte igitur mihi virum eruditum qui noverit operari in auro et argento aere ferro purpura coccino et hyacintho et qui sciat scalpere celata cum his artificibus quos mecum habeo in Iudaea et in Hierusalem quos praeparavit David pater meus
2CHR|2|8|sed et ligna cedrina mitte mihi et arceuthina et pinea de Libano scio enim quod servi tui noverint caedere ligna de Libano et erunt servi mei cum servis tuis
2CHR|2|9|ut parentur mihi ligna plurima domus enim quam cupio aedificare magna est nimis et inclita
2CHR|2|10|praeterea operariis qui caesuri sunt ligna servis tuis dabo in cibaria tritici choros viginti milia et hordei choros totidem olei quoque sata viginti milia
2CHR|2|11|dixit autem Hiram rex Tyri per litteras quas miserat Salomoni quia dilexit Dominus populum suum idcirco te regnare fecit super eum
2CHR|2|12|et addidit dicens benedictus Dominus Deus Israhel qui fecit caelum et terram qui dedit David regi filium sapientem et eruditum et sensatum atque prudentem ut aedificaret domum Domino et palatium sibi
2CHR|2|13|misi ergo tibi virum prudentem et scientissimum Hiram patrem meum
2CHR|2|14|filium mulieris de filiabus Dan cuius pater Tyrius fuit qui noverit operari in auro et argento et aere et ferro et marmore et lignis in purpura quoque et hyacintho et bysso et coccino et qui sciat celare omnem scalpturam et adinvenire prudenter quodcumque in opere necessarium est cum artificibus tuis et cum artificibus domini mei David patris tui
2CHR|2|15|triticum ergo et hordeum et oleum et vinum quae pollicitus es domine mi mitte servis tuis
2CHR|2|16|nos autem caedemus ligna de Libano quot necessaria habueris et adplicabimus ea ratibus per mare in Ioppe tuum erit transferre ea in Hierusalem
2CHR|2|17|numeravit igitur Salomon omnes viros proselytos qui erant in terra Israhel post dinumerationem quam dinumeravit David pater eius et inventi sunt centum quinquaginta milia et tria milia sescenti
2CHR|2|18|fecitque ex eis septuaginta milia qui umeris onera portarent et octoginta milia qui lapides in montibus caederent tria milia autem et sescentos praepositos operum populi
2CHR|3|1|et coepit Salomon aedificare domum Domini in Hierusalem in monte Moria qui demonstratus fuerat David patri eius in loco quem paraverat David in area Ornan Iebusei
2CHR|3|2|coepit autem aedificare mense secundo anno quarto regni sui
2CHR|3|3|et haec sunt fundamenta quae iecit Salomon ut aedificaret domum Dei longitudinis cubitos in mensura prima sexaginta latitudinis cubitos viginti
2CHR|3|4|porticum vero ante frontem quae tendebatur in longum iuxta mensuram latitudinis domus cubitorum viginti porro altitudo centum viginti cubitorum erat et deauravit eam intrinsecus auro mundissimo
2CHR|3|5|domum quoque maiorem texit tabulis ligneis abiegnis et lamminas auri obrizi adfixit per totum scalpsitque in ea palmas et quasi catenulas se invicem conplectentes
2CHR|3|6|stravit quoque pavimentum templi pretiosissimo marmore decore multo
2CHR|3|7|porro aurum erat probatissimum de cuius lamminis texit domum et trabes eius et postes et parietes et ostia et celavit cherubin in parietibus
2CHR|3|8|fecit quoque domum sancti sanctorum longitudinem iuxta latitudinem domus cubitorum viginti et latitudinem similiter viginti cubitorum et lamminis aureis texit eam quasi talentis sescentis
2CHR|3|9|sed et clavos fecit aureos ita ut singuli clavi siclos quinquagenos adpenderent cenacula quoque texit auro
2CHR|3|10|fecit etiam in domo sancti sanctorum cherubin duo opere statuario et texit eos auro
2CHR|3|11|alae cherubin viginti cubitis extendebantur ita ut una ala haberet cubitos quinque et tangeret parietem domus et altera quinque cubitos habens alam tangeret alterius cherub
2CHR|3|12|similiter cherub alterius ala quinque habebat cubitos et tangebat parietem et ala eius altera quinque cubitorum alam cherub alterius contingebat
2CHR|3|13|igitur alae utriusque cherubin expansae erant et extendebantur per cubitos viginti ipsi autem stabant erectis pedibus et facies eorum versae erant ad exteriorem domum
2CHR|3|14|fecit quoque velum ex hyacintho purpura coccino et bysso et intexuit ei cherubin
2CHR|3|15|ante fores etiam templi duas columnas quae triginta et quinque cubitos habebant altitudinis porro capita earum quinque cubitorum
2CHR|3|16|necnon et quasi catenulas in oraculo et superposuit eas capitibus columnarum malagranata etiam centum quae catenulis interposuit
2CHR|3|17|ipsas quoque columnas posuit in vestibulo templi unam a dextris et alteram a sinistris eam quae a dextris erat vocavit Iachin et quae ad levam Booz
2CHR|4|1|fecit quoque altare aeneum viginti cubitorum longitudinis et viginti cubitorum latitudinis et decem cubitorum altitudinis
2CHR|4|2|mare etiam fusile decem cubitis a labio usque ad labium rotundum per circuitum quinque cubitos habebat altitudinis et funiculus triginta cubitorum ambiebat gyrum eius
2CHR|4|3|similitudo quoque boum erat subter illud et decem cubitis quaedam extrinsecus celaturae quasi duobus versibus alvum maris circuibant boves autem erant fusiles
2CHR|4|4|et ipsum mare super duodecim boves inpositum erat quorum tres respiciebant aquilonem et alii tres occidentem porro tres alii meridiem et tres qui reliqui erant orientem mare habentes superpositum posteriora autem boum erant intrinsecus sub mari
2CHR|4|5|porro vastitas eius habebat mensuram palmi et labium illius erat quasi labium calicis vel repandi lilii capiebatque mensurae tria milia metretas
2CHR|4|6|fecit quoque concas decem et posuit quinque a dextris et quinque a sinistris ut lavarent in eis omnia quae in holocaustum oblaturi erant porro in mari sacerdotes lavabantur
2CHR|4|7|fecit autem et candelabra aurea decem secundum speciem qua iussa erant fieri et posuit ea in templo quinque a dextris et quinque a sinistris
2CHR|4|8|necnon et mensas decem posuitque eas in templo quinque a dextris et quinque a sinistris fialas quoque aureas centum
2CHR|4|9|fecit etiam atrium sacerdotum et basilicam grandem et ostia in basilica quae texit aere
2CHR|4|10|porro mare posuit in latere dextro contra orientem ad meridiem
2CHR|4|11|fecit autem Hiram lebetas quoque et creagras et fialas et conplevit omne opus regis in domo Dei
2CHR|4|12|hoc est columnas duas et epistylia et capita et quasi quaedam retiacula quae capita tegerent super epistylia
2CHR|4|13|malagranata quoque quadringenta et retiacula duo ita ut bini ordines malagranatorum singulis retiaculis iungerentur quae protegerent epistylia et capita columnarum
2CHR|4|14|bases etiam fecit et concas quas superposuit basibus
2CHR|4|15|mare unum bovesque duodecim sub mari
2CHR|4|16|et lebetas et creagras et fialas omnia vasa fecit Salomoni Hiram pater eius in domo Domini ex aere mundissimo
2CHR|4|17|in regione Iordanis fudit ea rex in argillosa terra inter Socchoth et Saredatha
2CHR|4|18|erat autem multitudo vasorum innumerabilis ita ut ignoraretur pondus aeris
2CHR|4|19|fecitque Salomon omnia vasa domus Dei et altare aureum et mensas et super eas panes propositionis
2CHR|4|20|candelabra quoque cum lucernis suis ut lucerent ante oraculum iuxta ritum ex auro purissimo
2CHR|4|21|et florentia quaedam et lucernas et forcipes aureos omnia de auro mundissimo facta sunt
2CHR|4|22|thymiamateria quoque et turibula et fialas et mortariola ex auro purissimo et ostia celavit templi interioris id est in sancto sanctorum et ostia templi forinsecus aurea sicque conpletum est omne opus quod fecit Salomon in domo Domini
2CHR|5|1|intulit igitur Salomon omnia quae voverat David pater suus argentum et aurum et universa vasa posuit in thesauris domus Dei
2CHR|5|2|post quae congregavit maiores natu Israhel et cunctos principes tribuum et capita familiarum de filiis Israhel in Hierusalem ut adducerent arcam foederis Domini de civitate David quae est Sion
2CHR|5|3|venerunt igitur ad regem omnes viri Israhel in die sollemni mensis septimi
2CHR|5|4|cumque venissent cuncti seniorum Israhel portaverunt Levitae arcam
2CHR|5|5|et intulerunt eam et omnem paraturam tabernaculi porro vasa sanctuarii quae erant in tabernaculo portaverunt sacerdotes cum Levitis
2CHR|5|6|rex autem Salomon et universus coetus Israhel et omnes qui fuerant congregati ante arcam immolabant arietes et boves absque ullo numero tanta enim erat multitudo victimarum
2CHR|5|7|et intulerunt sacerdotes arcam foederis Domini in locum suum id est ad oraculum templi in sancta sanctorum subter alas cherubin
2CHR|5|8|ita ut cherubin expanderent alas suas super locum in quo posita erat arca et ipsam arcam tegerent cum vectibus eius
2CHR|5|9|vectium autem quibus portabatur arca quia paululum longiores erant capita parebant ante oraculum si vero quis paululum fuisset extrinsecus eos videre non poterat fuit itaque arca ibi usque in praesentem diem
2CHR|5|10|nihilque erat aliud in arca nisi duae tabulae quas posuerat Moses in Horeb quando legem dedit Dominus filiis Israhel egredientibus ex Aegypto
2CHR|5|11|egressis autem sacerdotibus de sanctuario omnes enim sacerdotes qui ibi potuerant inveniri sanctificati sunt nec adhuc illo tempore vices et ministeriorum ordo inter eos divisus erat
2CHR|5|12|tam Levitae quam cantores id est et qui sub Asaph erant et qui sub Heman et qui sub Idithun filii et fratres eorum vestiti byssinis cymbalis et psalteriis et citharis concrepabant stantes ad orientalem plagam altaris cumque eis sacerdotes centum viginti canentes tubis
2CHR|5|13|igitur cunctis pariter et tubis et voce et cymbalis et organis et diversi generis musicorum concinentibus et vocem in sublime tollentibus longe sonitus audiebatur ita ut cum Dominum laudare coepissent et dicere confitemini Domino quoniam bonus quoniam in aeternum misericordia eius impleretur domus Domini nube
2CHR|5|14|nec possent sacerdotes stare et ministrare propter caliginem conpleverat enim gloria Domini domum Dei
2CHR|6|1|tunc Salomon ait Dominus pollicitus est ut habitaret in caligine
2CHR|6|2|ego autem aedificavi domum nomini eius ut habitaret ibi in perpetuum
2CHR|6|3|et convertit faciem suam et benedixit universae multitudini Israhel nam omnis turba stabat intenta et ait
2CHR|6|4|benedictus Dominus Deus Israhel qui quod locutus est David patri meo opere conplevit dicens
2CHR|6|5|a die qua eduxi populum meum de terra Aegypti non elegi civitatem de cunctis tribubus Israhel ut aedificaretur in ea domus nomini meo neque elegi quemquam alium virum ut esset dux in populo meo Israhel
2CHR|6|6|sed elegi Hierusalem ut sit nomen meum in ea et elegi David ut constituerem eum super populum meum Israhel
2CHR|6|7|cumque fuisset voluntatis David patris mei ut aedificaret domum nomini Domini Dei Israhel
2CHR|6|8|dixit Dominus ad eum quia haec fuit voluntas tua ut aedificares domum nomini meo bene quidem fecisti habere huiuscemodi voluntatem
2CHR|6|9|sed non tu aedificabis domum verum filius tuus qui egredietur de lumbis tuis ipse aedificabit domum nomini meo
2CHR|6|10|conplevit ergo Dominus sermonem suum quem locutus fuerat et ego surrexi pro David patre meo et sedi super thronum Israhel sicut locutus est Dominus et aedificavi domum nomini Domini Dei Israhel
2CHR|6|11|et posui in ea arcam in qua est pactum Domini quod pepigit cum filiis Israhel
2CHR|6|12|stetit ergo coram altare Domini ex adverso universae multitudinis Israhel et extendit manus suas
2CHR|6|13|siquidem fecerat Salomon basem aeneam et posuerat eam in medio basilicae habentem quinque cubitos longitudinis et quinque cubitos latitudinis et tres cubitos in altum stetitque super eam et deinceps flexis genibus contra universam multitudinem Israhel et palmis in caelum levatis
2CHR|6|14|ait Domine Deus Israhel non est similis tui Deus in caelo et in terra qui custodis pactum et misericordiam cum servis tuis qui ambulant coram te in toto corde suo
2CHR|6|15|qui praestitisti servo tuo David patri meo quaecumque locutus fueras ei et quae ore promiseras opere conplesti sicut et praesens tempus probat
2CHR|6|16|nunc ergo Domine Deus Israhel imple servo tuo patri meo David quaecumque locutus es dicens non deficiet ex te vir coram me qui sedeat super thronum Israhel ita tamen si custodierint filii tui vias suas et ambulaverint in lege mea sicut et tu ambulasti coram me
2CHR|6|17|et nunc Domine Deus Israhel firmetur sermo tuus quem locutus es servo tuo David
2CHR|6|18|ergone credibile est ut habitet Deus cum hominibus super terram si caelum et caeli caelorum non te capiunt quanto magis domus ista quam aedificavi
2CHR|6|19|sed ad hoc tantum facta est ut respicias orationem servi tui et obsecrationem eius Domine Deus meus audias et preces quas fundit famulus tuus coram te
2CHR|6|20|ut aperias oculos tuos super domum istam diebus et noctibus super locum in quo pollicitus es ut invocaretur nomen tuum
2CHR|6|21|et exaudires orationem quam servus tuus orat in eo exaudi preces famuli tui et populi tui Israhel quicumque oraverit in loco isto et exaudi de habitaculo tuo id est de caelis et propitiare
2CHR|6|22|si peccaverit quispiam in proximum suum et iurare contra eum paratus venerit seque maledicto constrinxerit coram altari in domo ista
2CHR|6|23|tu audies de caelo et facies iudicium servorum tuorum ita ut reddas iniquo viam suam in caput proprium et ulciscaris iustum retribuens ei secundum iustitiam suam
2CHR|6|24|si superatus fuerit populus tuus Israhel ab inimicis peccabunt enim tibi et conversi egerint paenitentiam et obsecraverint nomen tuum et fuerint deprecati in loco isto
2CHR|6|25|tu exaudi de caelo et propitiare peccato populi tui Israhel et reduc eos in terram quam dedisti eis et patribus eorum
2CHR|6|26|si clauso caelo pluvia non fluxerit propter peccata populi et deprecati te fuerint in loco isto et confessi nomini tuo et conversi a peccatis suis cum eos adflixeris
2CHR|6|27|exaudi de caelo Domine et dimitte peccata servis tuis et populi tui Israhel et doce eos viam bonam per quam ingrediantur et da pluviam terrae quam dedisti populo tuo ad possidendum
2CHR|6|28|fames si orta fuerit in terra et pestilentia erugo et aurugo et lucusta et brucus et hostes vastatis regionibus portas obsederint civitatis omnisque plaga et infirmitas presserit
2CHR|6|29|si quis de populo tuo Israhel fuerit deprecatus cognoscens plagam et infirmitatem suam et expanderit manus suas in domo hac
2CHR|6|30|tu exaudi de caelo de sublimi scilicet habitaculo tuo et propitiare et redde unicuique secundum vias suas quas nosti eum habere in corde suo tu enim solus nosti corda filiorum hominum
2CHR|6|31|ut timeant te et ambulent in viis tuis cunctis diebus quibus vivunt super faciem terrae quam dedisti patribus nostris
2CHR|6|32|externum quoque qui non est de populo tuo Israhel si venerit de terra longinqua propter nomen tuum magnum et propter manum tuam robustam et brachium tuum extentum et adoraverit in loco isto
2CHR|6|33|tu exaudies de caelo firmissimo habitaculo tuo et facies cuncta pro quibus invocaverit te ille peregrinus ut sciant omnes populi terrae nomen tuum et timeant te sicut populus tuus Israhel et cognoscant quia nomen tuum invocatum est super domum hanc quam aedificavi
2CHR|6|34|si egressus fuerit populus tuus ad bellum contra adversarios suos per viam in qua miseris eos adorabunt te contra viam in qua civitas haec est quam elegisti et domus quam aedificavi nomini tuo
2CHR|6|35|ut exaudias de caelo preces eorum et obsecrationem et ulciscaris
2CHR|6|36|si autem et peccaverint tibi neque enim est homo qui non peccet et iratus fueris eis et tradideris hostibus et captivos eos duxerint in terram longinquam vel certe quae iuxta est
2CHR|6|37|et conversi corde suo in terra ad quam captivi ducti fuerant egerint paenitentiam et deprecati te fuerint in terra captivitatis suae dicentes peccavimus inique fecimus iniuste egimus
2CHR|6|38|et reversi fuerint ad te in toto corde suo et in tota anima sua in terra captivitatis suae ad quam ducti sunt adorabunt te contra viam terrae suae quam dedisti patribus eorum et urbis quam elegisti et domus quam aedificavi nomini tuo
2CHR|6|39|ut exaudias de caelo hoc est de firmo habitaculo tuo preces eorum et facias iudicium et dimittas populo tuo quamvis peccatori
2CHR|6|40|tu es enim Deus meus aperiantur quaeso oculi tui et aures tuae intentae sint ad orationem quae fit in loco isto
2CHR|6|41|nunc igitur consurge Domine Deus in requiem tuam tu et arca fortitudinis tuae sacerdotes tui Domine Deus induantur salute et sancti tui laetentur in bonis
2CHR|6|42|Domine Deus ne averseris faciem christi tui memento misericordiarum David servi tui
2CHR|7|1|cumque conplesset Salomon fundens preces ignis descendit de caelo et devoravit holocausta et victimas et maiestas Domini implevit domum
2CHR|7|2|nec poterant sacerdotes ingredi templum Domini eo quod implesset maiestas Domini templum Domini
2CHR|7|3|sed et omnes filii Israhel videbant descendentem ignem et gloriam Domini super domum et corruentes proni in terram super pavimentum stratum lapide adoraverunt et laudaverunt Dominum quoniam bonus quoniam in aeternum misericordia eius
2CHR|7|4|rex autem et omnis populus immolabant victimas coram Domino
2CHR|7|5|mactavit igitur rex Salomon hostias boum viginti duo milia arietum centum viginti milia et dedicavit domum Dei rex et universus populus
2CHR|7|6|sacerdotes autem stabant in officiis suis et Levitae in organis carminum Domini quae fecit David rex ad laudandum Dominum quoniam in aeternum misericordia eius hymnos David canentes per manus suas porro sacerdotes canebant tubis ante eos cunctusque Israhel stabat
2CHR|7|7|sanctificavit quoque Salomon medium atrii ante templum Domini obtulerat enim ibi holocausta et adipes pacificorum quia altare aeneum quod fecerat non poterat sustinere holocausta et sacrificia et adipes
2CHR|7|8|fecit ergo Salomon sollemnitatem in tempore illo septem diebus et omnis Israhel cum eo ecclesia magna valde ab introitu Emath usque ad torrentem Aegypti
2CHR|7|9|fecitque die octavo collectam eo quod dedicasset altare septem diebus et sollemnitatem celebrasset diebus septem
2CHR|7|10|igitur in die vicesimo tertio mensis septimi dimisit populos ad tabernacula sua laetantes atque gaudentes super bono quod fecerat Dominus David et Salomoni et Israhel populo suo
2CHR|7|11|conplevitque Salomon domum Domini et domum regis et omnia quae disposuerat in corde suo ut faceret in domo Domini et in domo sua et prosperatus est
2CHR|7|12|apparuit autem ei Dominus nocte et ait audivi orationem tuam et elegi locum istum mihi in domum sacrificii
2CHR|7|13|si clausero caelum et pluvia non fluxerit et mandavero et praecepero lucustae ut devoret terram et misero pestilentiam in populum meum
2CHR|7|14|conversus autem populus meus super quos invocatum est nomen meum deprecatus me fuerit et exquisierit faciem meam et egerit paenitentiam a viis suis pessimis et ego exaudiam de caelo et propitius ero peccatis eorum et sanabo terram eorum
2CHR|7|15|oculi quoque mei erunt aperti et aures meae erectae ad orationem eius qui in loco isto oraverit
2CHR|7|16|elegi enim et sanctificavi locum istum ut sit nomen meum ibi in sempiternum et permaneant oculi mei et cor meum ibi cunctis diebus
2CHR|7|17|tu quoque si ambulaveris coram me sicut ambulavit David pater tuus et feceris iuxta omnia quae praecepi tibi et iustitias meas iudiciaque servaveris
2CHR|7|18|suscitabo thronum regni tui sicut pollicitus sum David patri tuo dicens non auferetur de stirpe tua vir qui sit princeps in Israhel
2CHR|7|19|si autem aversi fueritis et dereliqueritis iustitias meas et praecepta mea quae proposui vobis et abeuntes servieritis diis alienis et adoraveritis eos
2CHR|7|20|evellam vos de terra mea quam dedi vobis et domum hanc quam sanctificavi nomini meo proiciam a facie mea et tradam eam in parabolam et in exemplum cunctis populis
2CHR|7|21|et domus ista erit in proverbium universis transeuntibus et dicent stupentes quare fecit Dominus sic terrae huic et domui huic
2CHR|7|22|respondebuntque quia dereliquerunt Dominum Deum patrum suorum qui eduxit eos de terra Aegypti et adprehenderunt deos alienos et adoraverunt eos atque coluerunt idcirco venerunt super eos universa haec mala
2CHR|8|1|expletis autem viginti annis postquam aedificavit Salomon domum Domini et domum suam
2CHR|8|2|civitates quas dederat Hiram Salomoni aedificavit et habitare ibi fecit filios Israhel
2CHR|8|3|abiit quoque in Emath Suba et obtinuit eam
2CHR|8|4|et aedificavit Palmyram in deserto et alias civitates munitissimas aedificavit in Emath
2CHR|8|5|extruxitque Bethoron superiorem et Bethoron inferiorem civitates muratas habentes portas et vectes et seras
2CHR|8|6|Baalath etiam et omnes urbes firmissimas quae fuerunt Salomonis cunctasque urbes quadrigarum et urbes equitum omnia quae voluit Salomon atque disposuit aedificavit in Hierusalem et in Libano et in universa terra potestatis suae
2CHR|8|7|omnem populum qui derelictus fuerat de Hettheis et Amorreis et Ferezeis et Eveis et Iebuseis qui non erant de stirpe Israhel
2CHR|8|8|de filiis eorum et de posteris quos non interfecerant filii Israhel subiugavit Salomon in tributarios usque in diem hanc
2CHR|8|9|porro de filiis Israhel non posuit ut servirent operibus regis ipsi enim erant viri bellatores et duces primi et principes quadrigarum et equitum eius
2CHR|8|10|omnes autem principes exercitus regis Salomonis fuerunt ducenti quinquaginta qui erudiebant populum
2CHR|8|11|filiam vero Pharaonis transtulit de civitate David in domum quam aedificaverat ei dixit enim non habitabit uxor mea in domo David regis Israhel eo quod sanctificata sit quia ingressa est eam arca Domini
2CHR|8|12|tunc obtulit Salomon holocausta Domino super altare Domini quod extruxerat ante porticum
2CHR|8|13|ut per singulos dies offerretur in eo iuxta praeceptum Mosi in sabbatis et in kalendis et in festis diebus ter per annum id est in sollemnitate azymorum et in sollemnitate ebdomadarum et in sollemnitate tabernaculorum
2CHR|8|14|et constituit iuxta dispositionem David patris sui officia sacerdotum in ministeriis suis et Levitas in ordine suo ut laudarent et ministrarent coram sacerdotibus iuxta ritum uniuscuiusque diei et ianitores in divisionibus suis per portam et portam sic enim praeceperat David homo Dei
2CHR|8|15|nec praetergressi sunt de mandatis regis tam sacerdotes quam Levitae ex omnibus quae praeceperat et in custodiis thesaurorum
2CHR|8|16|omnes inpensas praeparatas habuit Salomon ex eo die quo fundavit domum Domini usque in diem quo perfecit eam
2CHR|8|17|tunc abiit Salomon in Hesiongaber et in Ahilath ad oram maris Rubri quae est in terra Edom
2CHR|8|18|misit autem ei Hiram per manum servorum suorum naves et nautas gnaros maris et abierunt cum servis Salomonis in Ophir tuleruntque inde quadringenta quinquaginta talenta auri et adtulerunt ad regem Salomonem
2CHR|9|1|regina quoque Saba cum audisset famam Salomonis venit ut temptaret eum enigmatibus in Hierusalem cum magnis opibus et camelis qui portabant aromata et auri plurimum gemmasque pretiosas cumque venisset ad Salomonem locuta est ei quaecumque erant in corde suo
2CHR|9|2|et exposuit ei Salomon omnia quae proposuerat nec quicquam fuit quod ei non perspicuum fecerit
2CHR|9|3|quod postquam vidit sapientiam scilicet Salomonis et domum quam aedificaverat
2CHR|9|4|necnon cibaria mensae eius et habitacula servorum et officia ministrorum eius et vestimenta eorum pincernas quoque et vestes eorum et victimas quas immolabat in domo Domini non erat prae stupore ultra in ea spiritus
2CHR|9|5|dixitque ad regem verus sermo quem audieram in terra mea de virtutibus et sapientia tua
2CHR|9|6|non credebam narrantibus donec ipsa venissem et vidissent oculi mei et probassem vix medietatem mihi sapientiae tuae fuisse narratam vicisti famam virtutibus tuis
2CHR|9|7|beati viri tui et beati servi tui hii qui adsistunt coram te in omni tempore et audiunt sapientiam tuam
2CHR|9|8|sit Dominus Deus tuus benedictus qui voluit te ordinare super thronum suum regem Domini Dei tui quia diligit Deus Israhel et vult servare eum in aeternum idcirco posuit te super eum regem ut facias iudicia atque iustitiam
2CHR|9|9|dedit autem regi centum viginti talenta auri et aromata multa nimis et gemmas pretiosissimas non fuerunt aromata talia ut haec quae dedit regina Saba regi Salomoni
2CHR|9|10|sed et servi Hiram cum servis Salomonis adtulerunt aurum de Ophir et ligna thyina et gemmas pretiosissimas
2CHR|9|11|de quibus fecit rex de lignis scilicet thyinis gradus in domo Domini et in domo regia citharas quoque et psalteria cantoribus numquam visa sunt in terra Iuda ligna talia
2CHR|9|12|rex autem Salomon dedit reginae Saba cuncta quae voluit et quae postulavit multo plura quam adtulerat ad eum quae reversa abiit in terram suam cum servis suis
2CHR|9|13|erat autem pondus auri quod adferebatur Salomoni per annos singulos sescenta sexaginta sex talenta auri
2CHR|9|14|excepta ea summa quam legati diversarum gentium et negotiatores adferre consueverant omnesque reges Arabiae et satrapae terrarum qui conportabant aurum et argentum Salomoni
2CHR|9|15|fecit igitur rex Salomon ducentas hastas aureas de summa sescentorum aureorum qui in hastis singulis expendebantur
2CHR|9|16|trecenta quoque scuta aurea trecentorum aureorum quibus tegebantur scuta singula posuitque ea rex in armamentario quod erat consitum nemore
2CHR|9|17|fecit quoque rex solium eburneum grande et vestivit illud auro mundissimo
2CHR|9|18|sexque gradus quibus ascendebatur ad solium et scabillum aureum et brachiola duo altrinsecus et duos leones stantes iuxta brachiola
2CHR|9|19|sed et alios duodecim leunculos stantes super sex gradus ex utraque parte non fuit tale solium in universis regnis
2CHR|9|20|omnia quoque vasa convivii regis erant aurea et vasa domus saltus Libani ex auro purissimo argentum enim in diebus illis pro nihilo reputabatur
2CHR|9|21|siquidem naves regis ibant in Tharsis cum servis Hiram semel in annis tribus et deferebant inde aurum et argentum et ebur et simias et pavos
2CHR|9|22|magnificatus est igitur Salomon super omnes reges terrae divitiis et gloria
2CHR|9|23|omnesque reges terrarum desiderabant faciem videre Salomonis ut audirent sapientiam quam dederat Deus in corde eius
2CHR|9|24|et deferebant ei munera vasa argentea et aurea et vestes et arma et aromata equos et mulos per singulos annos
2CHR|9|25|habuit quoque Salomon quadraginta milia equorum in stabulis et curruum equitumque duodecim milia constituitque eos in urbibus quadrigarum et ubi erat rex in Hierusalem
2CHR|9|26|exercuit etiam potestatem super cunctos reges a fluvio Eufraten usque ad terram Philisthinorum id est usque ad terminos Aegypti
2CHR|9|27|tantamque copiam praebuit argenti in Hierusalem quasi lapidum et cedrorum tantam multitudinem velut sycaminorum quae gignuntur in campestribus
2CHR|9|28|adducebantur autem ei equi de Aegypto cunctisque regionibus
2CHR|9|29|reliqua vero operum Salomonis priorum et novissimorum scripta sunt in verbis Nathan prophetae et in libris Ahiae Silonitis in visione quoque Iaddo videntis contra Hieroboam filium Nabath
2CHR|9|30|regnavit autem Salomon in Hierusalem super omnem Israhel quadraginta annis
2CHR|9|31|dormivitque cum patribus suis et sepelierunt eum in civitate David regnavitque pro eo Roboam filius eius
2CHR|10|1|profectus est autem Roboam in Sychem illuc enim cunctus Israhel convenerat ut constituerent eum regem
2CHR|10|2|quod cum audisset Hieroboam filius Nabath qui erat in Aegypto fugerat quippe illuc ante Salomonem statim reversus est
2CHR|10|3|vocaveruntque eum et venit cum universo Israhel et locuti sunt ad Roboam dicentes
2CHR|10|4|pater tuus durissimo iugo nos pressit tu leviora impera patre tuo qui nobis gravem inposuit servitutem et paululum de onere subleva ut serviamus tibi
2CHR|10|5|qui ait post tres dies revertimini ad me cumque abisset populus
2CHR|10|6|iniit consilium cum senibus qui steterant coram patre eius Salomone dum adviveret dicens quid datis consilii ut respondeam populo
2CHR|10|7|qui dixerunt ei si placueris populo huic et lenieris eos verbis clementibus servient tibi omni tempore
2CHR|10|8|at ille reliquit consilium senum et cum iuvenibus tractare coepit qui cum eo nutriti fuerant et erant in comitatu illius
2CHR|10|9|dixitque ad eos quid vobis videtur vel respondere quid debeo populo huic qui dixit mihi subleva iugum quod inposuit nobis pater tuus
2CHR|10|10|at illi responderunt ut iuvenes et nutriti cum eo in deliciis atque dixerunt sic loqueris populo qui dixit tibi pater tuus adgravavit iugum nostrum tu subleva et sic respondebis eis minimus digitus meus grossior est lumbis patris mei
2CHR|10|11|pater meus inposuit vobis iugum grave et ego maius pondus adponam pater meus cecidit vos flagellis ego vero caedam scorpionibus
2CHR|10|12|venit ergo Hieroboam et universus populus ad Roboam die tertio sicut praeceperat eis
2CHR|10|13|responditque rex dura derelicto consilio seniorum
2CHR|10|14|locutusque est iuxta iuvenum voluntatem pater meus grave vobis inposuit iugum quod ego gravius faciam pater meus cecidit vos flagellis ego vero caedam scorpionibus
2CHR|10|15|et non adquievit populi precibus erat enim voluntatis Dei ut conpleretur sermo eius quem locutus fuerat per manum Ahiae Silonitis ad Hieroboam filium Nabath
2CHR|10|16|populus autem universus rege duriora dicente sic locutus est ad eum non est nobis pars in David neque hereditas in filio Isai revertere in tabernacula tua Israhel tu autem pasce domum tuam David et abiit Israhel in tabernacula sua
2CHR|10|17|super filios autem Israhel qui habitabant in civitatibus Iuda regnavit Roboam
2CHR|10|18|misitque rex Roboam Aduram qui praeerat tributis et lapidaverunt eum filii Israhel et mortuus est porro rex Roboam currum festinavit ascendere et fugit in Hierusalem
2CHR|10|19|recessitque Israhel a domo David usque ad diem hanc
2CHR|11|1|venit autem Roboam in Hierusalem et convocavit universam domum Iuda et Beniamin in centum octoginta milibus electorum atque bellantium ut dimicaret contra Israhel et converteret ad se regnum suum
2CHR|11|2|factusque est sermo Domini ad Semeiam hominem Dei dicens
2CHR|11|3|loquere ad Roboam filium Salomonis regem Iuda et ad universum Israhel qui est in Iuda et Beniamin
2CHR|11|4|haec dicit Dominus non ascendetis neque pugnabitis contra fratres vestros revertatur unusquisque in domum suam quia mea hoc gestum est voluntate qui cum audissent sermonem Domini reversi sunt nec perrexerunt contra Hieroboam
2CHR|11|5|habitavit autem Roboam in Hierusalem et aedificavit civitates muratas in Iuda
2CHR|11|6|extruxitque Bethleem et Aetham et Thecue
2CHR|11|7|Bethsur quoque et Soccho et Odollam
2CHR|11|8|necnon Geth et Maresa et Ziph
2CHR|11|9|sed et Aduram et Lachis et Azecha
2CHR|11|10|Saraa quoque et Ahilon et Hebron quae erant in Iuda et Beniamin civitates munitissimas
2CHR|11|11|cumque clausisset eas muris posuit in eis principes ciborumque horrea hoc est olei et vini
2CHR|11|12|sed et in singulis urbibus fecit armamentaria scutorum et hastarum firmavitque eas multa diligentia et imperavit super Iudam et Beniamin
2CHR|11|13|sacerdotes autem et Levitae qui erant in universo Israhel venerunt ad eum de cunctis sedibus suis
2CHR|11|14|relinquentes suburbana et possessiones suas et transeuntes ad Iudam et Hierusalem eo quod abiecisset eos Hieroboam et posteri eius ne sacerdotio Domini fungerentur
2CHR|11|15|qui constituit sibi sacerdotes excelsorum et daemonum vitulorumque quos fecerat
2CHR|11|16|sed et de cunctis tribubus Israhel quicumque dederant cor suum ut quaererent Dominum Deum Israhel venerunt Hierusalem ad immolandas victimas Domino Deo patrum suorum
2CHR|11|17|et roboraverunt regnum Iuda et confirmaverunt Roboam filium Salomonis per tres annos ambulaverunt enim in viis David et Salomonis annis tantum tribus
2CHR|11|18|duxit autem Roboam uxorem Maalath filiam Hierimuth filii David Abiail quoque filiam Heliab filii Isai
2CHR|11|19|quae peperit ei filios Ieus et Somoriam et Zoom
2CHR|11|20|post hanc quoque accepit Maacha filiam Absalom quae peperit ei Abia et Ethai et Ziza et Salumith
2CHR|11|21|amavit autem Roboam Maacha filiam Absalom super omnes uxores suas et concubinas nam uxores decem et octo duxerat concubinasque sexaginta et genuit viginti octo filios et sexaginta filias
2CHR|11|22|constituit vero in capite Abiam filium Maacha ducem super fratres suos ipsum enim regem facere cogitabat
2CHR|11|23|qui sapientior fuit et potentior super omnes filios eius et in cunctis finibus Iuda et Beniamin et in universis civitatibus muratis praebuitque eis escas plurimas et multas petivit uxores
2CHR|12|1|cumque roboratum fuisset regnum Roboam et confortatum dereliquit legem Domini et omnis Israhel cum eo
2CHR|12|2|anno autem quinto regni Roboam ascendit Sesac rex Aegypti in Hierusalem quia peccaverunt Domino
2CHR|12|3|cum mille ducentis curribus et sexaginta milibus equitum nec erat numerus vulgi quod venerat cum eo ex Aegypto Lybies scilicet et Trogoditae et Aethiopes
2CHR|12|4|cepitque civitates munitissimas in Iuda et venit usque Hierusalem
2CHR|12|5|Semeias autem propheta ingressus est ad Roboam et principes Iuda qui congregati fuerant in Hierusalem fugientes Sesac dixitque ad eos haec dicit Dominus vos reliquistis me et ego reliqui vos in manu Sesac
2CHR|12|6|consternatique principes Israhel et rex dixerunt iustus est Dominus
2CHR|12|7|cumque vidisset Dominus quod humiliati essent factus est sermo Domini ad Semeiam dicens quia humiliati sunt non disperdam eos daboque eis pauxillum auxilii et non stillabit furor meus super Hierusalem per manum Sesac
2CHR|12|8|verumtamen servient ei ut sciant distantiam servitutis meae et servitutis regni terrarum
2CHR|12|9|recessit itaque Sesac rex Aegypti ab Hierusalem sublatis thesauris domus Domini et domus regis omniaque secum tulit et clypeos aureos quos fecerat Salomon
2CHR|12|10|pro quibus fecit rex aeneos et tradidit illos principibus scutariorum qui custodiebant vestibulum palatii
2CHR|12|11|cumque introiret rex domum Domini veniebant scutarii et tollebant eos iterumque referebant ad armamentarium suum
2CHR|12|12|verumtamen quia humiliati sunt aversa est ab eis ira Domini nec deleti sunt penitus siquidem et in Iuda inventa sunt opera bona
2CHR|12|13|confortatus est igitur rex Roboam in Hierusalem atque regnavit quadraginta autem et unius anni erat cum regnare coepisset et decem septemque annis regnavit in Hierusalem urbe quam elegit Dominus ut confirmaret nomen suum ibi de cunctis tribubus Israhel nomenque matris eius Naama Ammanitis
2CHR|12|14|fecit autem malum et non praeparavit cor suum ut quaereret Dominum
2CHR|12|15|opera vero Roboam prima et novissima scripta sunt in libris Semeiae prophetae et Addo videntis et diligenter exposita pugnaveruntque adversum se Roboam et Hieroboam cunctis diebus
2CHR|12|16|et dormivit Roboam cum patribus suis sepultusque est in civitate David et regnavit Abia filius eius pro eo
2CHR|13|1|anno octavodecimo regis Hieroboam regnavit Abia super Iudam
2CHR|13|2|tribus annis regnavit in Hierusalem nomenque matris eius Michaia filia Urihel de Gabaa et erat bellum inter Abia et Hieroboam
2CHR|13|3|cumque inisset Abia certamen et haberet bellicosissimos viros et electorum quadringenta milia Hieroboam instruxit e contra aciem octingenta milia virorum qui et ipsi electi erant et ad bella fortissimi
2CHR|13|4|stetit igitur Abia super montem Someron qui erat in Ephraim et ait audi Hieroboam et omnis Israhel
2CHR|13|5|num ignoratis quod Dominus Deus Israhel dederit regnum David super Israhel in sempiternum ipsi et filiis eius pactum salis
2CHR|13|6|et surrexit Hieroboam filius Nabath servus Salomonis filii David et rebellavit contra dominum suum
2CHR|13|7|congregatique sunt ad eum viri vanissimi et filii Belial et praevaluerunt contra Roboam filium Salomonis porro Roboam erat rudis et corde pavido nec potuit resistere eis
2CHR|13|8|nunc ergo vos dicitis quod resistere possitis regno Domini quod possidet per filios David habetisque grandem populi multitudinem atque vitulos aureos quos fecit vobis Hieroboam in deos
2CHR|13|9|et eiecistis sacerdotes Domini filios Aaron atque Levitas et fecistis vobis sacerdotes sicut omnes populi terrarum quicumque venerit et initiaverit manum suam in tauro in bubus et in arietibus septem fit sacerdos eorum qui non sunt dii
2CHR|13|10|noster autem Dominus Deus est quem non relinquimus sacerdotesque ministrant Domino de filiis Aaron et Levitae sunt in ordine suo
2CHR|13|11|holocausta quoque offerunt Domino per singulos dies mane et vespere et thymiama iuxta legis praecepta confectum et proponuntur panes in mensa mundissima estque apud nos candelabrum aureum et lucernae eius ut accendantur semper ad vesperam nos quippe custodimus praecepta Domini Dei nostri quem vos reliquistis
2CHR|13|12|ergo in exercitu nostro dux Deus est et sacerdotes eius qui clangunt tubis et resonant contra vos filii Israhel nolite pugnare contra Dominum Deum patrum vestrorum quia non vobis expedit
2CHR|13|13|haec illo loquente Hieroboam retro moliebatur insidias cumque ex adverso hostium staret ignorantem Iudam suo ambiebat exercitu
2CHR|13|14|respiciensque Iudas vidit instare bellum ex adverso et post tergum et clamavit ad Dominum ac sacerdotes tubis canere coeperunt
2CHR|13|15|omnesque viri Iuda vociferati sunt et ecce illis clamantibus perterruit Deus Hieroboam et omnem Israhel qui stabat ex adverso Abia et Iuda
2CHR|13|16|fugeruntque filii Israhel Iudam et tradidit eos Deus in manu eorum
2CHR|13|17|percussit ergo eos Abia et populus eius plaga magna et corruerunt vulnerati ex Israhel quingenta milia virorum fortium
2CHR|13|18|humiliatique sunt filii Israhel in tempore illo et vehementissime confortati filii Iuda eo quod sperassent in Domino Deo patrum suorum
2CHR|13|19|persecutus est autem Abia fugientem Hieroboam et cepit civitates eius Bethel et filias eius et Hiesena cum filiabus suis Ephron quoque et filias eius
2CHR|13|20|nec valuit ultra resistere Hieroboam in diebus Abia quem percussit Dominus et mortuus est
2CHR|13|21|igitur Abia confortato imperio suo accepit uxores quattuordecim procreavitque viginti duos filios et sedecim filias
2CHR|13|22|reliqua autem sermonum Abia viarumque et operum eius scripta sunt diligentissime in libro prophetae Addo
2CHR|14|1|dormivit autem Abia cum patribus suis et sepelierunt eum in civitate David regnavitque Asa filius eius pro eo in cuius diebus quievit terra annis decem
2CHR|14|2|fecit autem Asa quod bonum et placitum erat in conspectu Dei sui et subvertit altaria peregrini cultus et excelsa
2CHR|14|3|et confregit statuas lucosque succidit
2CHR|14|4|ac praecepit Iudae ut quaereret Dominum Deum patrum suorum et faceret legem et universa mandata
2CHR|14|5|et abstulit e cunctis urbibus Iuda aras et fana et regnavit in pace
2CHR|14|6|aedificavit quoque urbes munitas in Iuda quia quietus erat et nulla temporibus eius bella surrexerant pacem Domino largiente
2CHR|14|7|dixit autem Iudae aedificemus civitates istas et vallemus muris et roboremus turribus et portis et seris donec a bellis quieta sunt omnia eo quod quaesierimus Dominum Deum patrum nostrorum et dederit nobis pacem per gyrum aedificaverunt igitur et nullum in extruendo inpedimentum fuit
2CHR|14|8|habuit autem Asa in exercitu suo portantium scuta et hastas de Iuda trecenta milia de Beniamin vero scutariorum et sagittariorum ducenta octoginta milia omnes isti viri fortissimi
2CHR|14|9|egressus est autem contra eos Zara Aethiops cum exercitu decies centena milia et curribus trecentis et venit usque Maresa
2CHR|14|10|porro Asa perrexit obviam et instruxit aciem ad bellum in valle Sephata quae est iuxta Maresa
2CHR|14|11|et invocavit Dominum Deum et ait Domine non est apud te ulla distantia utrum in paucis auxilieris an in pluribus adiuva nos Domine Deus noster in te enim et in tuo nomine habentes fiduciam venimus contra hanc multitudinem Domine Deus noster tu es non praevaleat contra te homo
2CHR|14|12|exterruit itaque Dominus Aethiopas coram Asa et Iuda fugeruntque Aethiopes
2CHR|14|13|et persecutus est eos Asa et populus qui cum eo erat usque Gerar et ruerunt Aethiopes usque ad internicionem quia Domino caedente contriti sunt et exercitu illius proeliante tulerunt ergo spolia multa
2CHR|14|14|et percusserunt omnes civitates per circuitum Gerare grandis quippe cunctos terror invaserat et diripuerunt urbes et multam praedam asportaverunt
2CHR|14|15|sed et caulas ovium destruentes tulerunt pecorum infinitam multitudinem et camelorum reversique sunt Hierusalem
2CHR|15|1|Azarias autem filius Oded facto in se spiritu Dei
2CHR|15|2|egressus est in occursum Asa et dixit ei audite me Asa et omnis Iuda et Beniamin Dominus vobiscum quia fuistis cum eo si quaesieritis eum invenietis si autem dereliqueritis derelinquet vos
2CHR|15|3|transibunt autem multi dies in Israhel absque Deo vero et absque sacerdote doctore et absque lege
2CHR|15|4|cumque reversi fuerint in angustia sua ad Dominum Deum Israhel et quaesierint eum repperient
2CHR|15|5|in tempore illo non erit pax egredienti et ingredienti sed terrores undique in cunctis habitatoribus terrarum
2CHR|15|6|pugnabit enim gens contra gentem et civitas contra civitatem quia Dominus conturbabit eos in omni angustia
2CHR|15|7|vos ergo confortamini et non dissolvantur manus vestrae erit enim merces operi vestro
2CHR|15|8|quod cum audisset Asa verba scilicet et prophetiam Oded prophetae confortatus est et abstulit idola de omni terra Iuda et Beniamin et ex urbibus quas ceperat montis Ephraim et dedicavit altare Domini quod erat ante porticum Domini
2CHR|15|9|congregavitque universum Iuda et Beniamin et advenas cum eis de Ephraim et de Manasse et de Symeon plures enim ad eum confugerant ex Israhel videntes quod Dominus Deus illius esset cum eo
2CHR|15|10|cumque venissent Hierusalem mense tertio anno quintodecimo regni Asa
2CHR|15|11|immolaverunt Domino in die illa de manubiis et praeda quam adduxerant boves septingentos et arietes septem milia
2CHR|15|12|et intravit ex more ad corroborandum foedus ut quaererent Dominum Deum patrum suorum in toto corde et in tota anima sua
2CHR|15|13|si quis autem inquit non quaesierit Dominum Deum Israhel moriatur a minimo usque ad maximum a viro usque ad mulierem
2CHR|15|14|iuraveruntque Domino voce magna in iubilo et in clangore tubae et in sonitu bucinarum
2CHR|15|15|omnes qui erant in Iuda cum execratione in omni enim corde suo iuraverunt et in tota voluntate quaesierunt eum et invenerunt praestititque eis Dominus requiem per circuitum
2CHR|15|16|sed et Maacham matrem Asa regis ex augusto deposuit imperio eo quod fecisset in luco simulacrum Priapi quod omne contrivit et in frusta comminuens conbusit in torrente Cedron
2CHR|15|17|excelsa autem derelicta sunt in Israhel attamen cor Asa erat perfectum cunctis diebus eius
2CHR|15|18|ea quae voverat pater suus et ipse intulit in domum Domini argentum et aurum vasorumque diversam supellectilem
2CHR|15|19|bellum vero non fuit usque ad tricesimum quintum annum regni Asa
2CHR|16|1|anno autem tricesimo sexto regni eius ascendit Baasa rex Israhel in Iudam et muro circumdabat Rama ut nullus tute posset egredi et ingredi de regno Asa
2CHR|16|2|protulit ergo Asa argentum et aurum de thesauris domus Domini et de thesauris regis misitque ad Benadad regem Syriae qui habitabat in Damasco dicens
2CHR|16|3|foedus inter me et te est pater quoque meus et pater tuus habuere concordiam quam ob rem misi tibi argentum et aurum ut rupto foedere quod habes cum Baasa rege Israhel facias eum a me recedere
2CHR|16|4|quo conperto Benadad misit principes exercituum suorum ad urbes Israhel qui percusserunt Ahion et Dan et Abelmaim et universas urbes muratas Nepthalim
2CHR|16|5|quod cum audisset Baasa desivit aedificare Rama et intermisit opus suum
2CHR|16|6|porro Asa rex adsumpsit universum Iudam et tulerunt lapides Rama et ligna quae aedificationi praeparaverat Baasa aedificavitque ex eis Gabaa et Maspha
2CHR|16|7|in tempore illo venit Anani propheta ad Asam regem Iuda et dixit ei quia habuisti fiduciam in rege Syriae et non in Domino Deo tuo idcirco evasit Syriae regis exercitus de manu tua
2CHR|16|8|nonne Aethiopes et Lybies multo plures erant quadrigis et equitibus et multitudine nimia quos cum Domino credidisses tradidit in manu tua
2CHR|16|9|oculi enim eius contemplantur universam terram et praebent fortitudinem his qui corde perfecto credunt in eum stulte igitur egisti et propter hoc ex praesenti tempore contra te bella consurgent
2CHR|16|10|iratusque Asa adversus videntem iussit eum mitti in nervum valde quippe super hoc fuerat indignatus et interfecit de populo in tempore illo plurimos
2CHR|16|11|opera autem Asa prima et novissima scripta sunt in libro regum Iuda et Israhel
2CHR|16|12|aegrotavit etiam Asa anno tricesimo nono regni sui dolore pedum vehementissimo et nec in infirmitate sua quaesivit Dominum sed magis in medicorum arte confisus est
2CHR|16|13|dormivitque cum patribus suis et mortuus est anno quadragesimo primo regni sui
2CHR|16|14|et sepelierunt eum in sepulchro suo quod foderat sibi in civitate David posueruntque eum super lectulum suum plenum aromatibus et unguentis meretriciis quae erant pigmentariorum arte confecta et conbuserunt super eum ambitione nimia
2CHR|17|1|regnavit autem Iosaphat filius eius pro eo et invaluit contra Israhel
2CHR|17|2|constituitque militum numeros in cunctis urbibus Iudae quae erant vallatae muris praesidiaque disposuit in terra Iuda et in civitatibus Ephraim quas ceperat Asa pater eius
2CHR|17|3|et fuit Dominus cum Iosaphat quia ambulavit in viis David patris sui primis et non speravit in Baalim
2CHR|17|4|sed in Deo patris sui et perrexit in praeceptis illius et non iuxta peccata Israhel
2CHR|17|5|confirmavitque Dominus regnum in manu eius et dedit omnis Iuda munera Iosaphat factaeque sunt ei infinitae divitiae et multa gloria
2CHR|17|6|cumque sumpsisset cor eius audaciam propter vias Domini etiam excelsa et lucos de Iuda abstulit
2CHR|17|7|tertio autem anno regni sui misit de principibus suis Benail et Obdiam et Zacchariam et Nathanahel et Micheam ut docerent in civitatibus Iuda
2CHR|17|8|et cum eis Levitas Semeiam et Nathaniam et Zabadiam Asahel quoque et Semiramoth et Ionathan Adoniam et Tobiam et Tobadoniam Levitas et cum eis Elisama et Ioram sacerdotes
2CHR|17|9|docebantque in Iuda habentes librum legis Domini et circuibant cunctas urbes Iuda atque erudiebant populum
2CHR|17|10|itaque factus est pavor Domini super omnia regna terrarum quae erant per gyrum Iuda nec audebant bellare contra Iosaphat
2CHR|17|11|sed et Philisthei Iosaphat munera deferebant et vectigal argenti Arabes quoque adducebant pecora arietum septem milia septingentos et hircos totidem
2CHR|17|12|crevit ergo Iosaphat et magnificatus est usque in sublime atque aedificavit in Iuda domos ad instar turrium urbesque muratas
2CHR|17|13|et multa opera patravit in urbibus Iuda viri quoque bellatores et robusti erant in Hierusalem
2CHR|17|14|quorum iste numerus per domos atque familias singulorum in Iuda principes exercitus Ednas dux et cum eo robustissimorum trecenta milia
2CHR|17|15|post hunc Iohanan princeps et cum eo ducenta octoginta milia
2CHR|17|16|post istum quoque Amasias filius Zechri consecratus Domino et cum eo ducenta milia virorum fortium
2CHR|17|17|hunc sequebatur robustus ad proelia Heliada et cum eo tenentium arcum et clypeum ducenta milia
2CHR|17|18|post istum etiam Iozabath et cum eo centum octoginta milia expeditorum militum
2CHR|17|19|hii omnes erant ad manum regis exceptis aliis quos posuerat in urbibus muratis et in universo Iuda
2CHR|18|1|fuit ergo Iosaphat dives et inclitus multum et adfinitate coniunctus est Ahab
2CHR|18|2|descenditque post annos ad eum in Samariam ad cuius adventum mactavit Ahab arietes et boves plurimos et populo qui venerat cum eo persuasitque illi ut ascenderet in Ramoth Galaad
2CHR|18|3|dixitque Ahab rex Israhel ad Iosaphat regem Iuda veni mecum in Ramoth Galaad cui ille respondit ut ego et tu sicut populus tuus sic et populus meus tecumque erimus in bello
2CHR|18|4|dixitque Iosaphat ad regem Israhel consule obsecro inpraesentiarum sermonem Domini
2CHR|18|5|congregavitque rex Israhel prophetarum quadringentos viros et dixit ad eos in Ramoth Galaad ad bellandum ire debemus an quiescere at illi ascende inquiunt et tradet Deus in manu regis
2CHR|18|6|dixitque Iosaphat numquid non est hic prophetes Domini ut ab illo etiam requiramus
2CHR|18|7|et ait rex Israhel ad Iosaphat est vir unus a quo possumus quaerere Domini voluntatem sed ego odi eum quia non prophetat mihi bonum sed malum omni tempore est autem Micheas filius Iembla dixitque Iosaphat ne loquaris rex hoc modo
2CHR|18|8|vocavit ergo rex Israhel unum de eunuchis et dixit ei voca cito Micheam filium Iembla
2CHR|18|9|porro rex Israhel et Iosaphat rex Iuda uterque sedebant in solio suo vestiti cultu regio sedebant autem in area iuxta portam Samariae omnesque prophetae vaticinabantur coram eis
2CHR|18|10|Sedecias vero filius Chanana fecit sibi cornua ferrea et ait haec dicit Dominus his ventilabis Syriam donec conteras eam
2CHR|18|11|omnesque prophetae similiter prophetabant atque dicebant ascende in Ramoth Galaad et prosperaberis et tradet eos Dominus in manu regis
2CHR|18|12|nuntius autem qui ierat ad vocandum Micheam ait illi en verba omnium prophetarum uno ore bona regi adnuntiant quaeso ergo te ut et sermo tuus ab eis non dissentiat loquarisque prospera
2CHR|18|13|cui respondit Micheas vivit Dominus quia quodcumque dixerit Deus meus hoc loquar
2CHR|18|14|venit ergo ad regem cui rex ait Michea ire debemus in Ramoth Galaad ad bellandum an quiescere cui ille respondit ascendite cuncta enim prospera evenient et tradentur hostes in manus vestras
2CHR|18|15|dixitque rex iterum atque iterum te adiuro ut non mihi loquaris nisi quod verum est in nomine Domini
2CHR|18|16|at ille ait vidi universum Israhel dispersum in montibus sicut oves absque pastore et dixit Dominus non habent isti dominos revertatur unusquisque ad domum suam in pace
2CHR|18|17|et ait rex Israhel ad Iosaphat nonne dixi tibi quod non prophetaret iste mihi quicquam boni sed ea quae mala sunt
2CHR|18|18|at ille idcirco ait audite verbum Domini vidi Dominum sedentem in solio suo et omnem exercitum caeli adsistentem ei a dextris et sinistris
2CHR|18|19|et dixit Dominus quis decipiet Ahab regem Israhel ut ascendat et corruat in Ramoth Galaad cumque diceret unus hoc modo et alter alio
2CHR|18|20|processit spiritus et stetit coram Domino et ait ego decipiam eum cui Dominus in quo inquit decipies
2CHR|18|21|at ille respondit egrediar et ero spiritus mendax in ore omnium prophetarum eius dixitque Dominus decipies et praevalebis egredere et fac ita
2CHR|18|22|nunc igitur ecce dedit Dominus spiritum mendacii in ore omnium prophetarum tuorum et Dominus locutus est de te mala
2CHR|18|23|accessit autem Sedecias filius Chanana et percussit Micheae maxillam et ait per quam viam transivit spiritus Domini a me ut loqueretur tibi
2CHR|18|24|dixitque Micheas tu ipse videbis in die illo quando ingressus fueris cubiculum de cubiculo ut abscondaris
2CHR|18|25|praecepit autem rex Israhel dicens tollite Micheam et ducite eum ad Amon principem civitatis et ad Ioas filium Ammelech
2CHR|18|26|et dicetis haec dicit rex mittite hunc in carcerem et date ei panis modicum et aquae pauxillum donec revertar in pace
2CHR|18|27|dixitque Micheas si reversus fueris in pace non est locutus Dominus in me et ait audite populi omnes
2CHR|18|28|igitur ascenderunt rex Israhel et Iosaphat rex Iuda in Ramoth Galaad
2CHR|18|29|dixitque rex Israhel ad Iosaphat mutabo habitum et sic ad pugnandum vadam tu autem induere vestibus tuis mutatoque rex Israhel habitu venit ad bellum
2CHR|18|30|rex autem Syriae praeceperat ducibus equitatus sui dicens ne pugnetis contra minimum aut contra maximum nisi contra solum regem Israhel
2CHR|18|31|itaque cum vidissent principes equitatus Iosaphat dixerunt rex Israhel iste est et circumdederunt eum dimicantes at ille clamavit ad Dominum et auxiliatus est ei atque avertit eos ab illo
2CHR|18|32|cum enim vidissent duces equitatus quod non esset rex Israhel reliquerunt eum
2CHR|18|33|accidit autem ut unus e populo sagittam in incertum iaceret et percuteret regem Israhel inter cervicem et scapulas at ille aurigae suo ait converte manum tuam et educ me de acie quia vulneratus sum
2CHR|18|34|et finita est pugna in die illo porro rex Israhel stabat in curru suo contra Syros usque ad vesperam et mortuus est occidente sole
2CHR|19|1|reversus est autem Iosaphat rex Iuda domum suam pacifice in Hierusalem
2CHR|19|2|cui occurrit Hieu filius Anani videns et ait ad eum impio praebes auxilium et his qui oderunt Dominum amicitia iungeris et idcirco iram quidem Domini merebaris
2CHR|19|3|sed bona opera inventa sunt in te eo quod abstuleris lucos de terra Iuda et praeparaveris cor tuum ut requireres Dominum
2CHR|19|4|habitavit ergo Iosaphat in Hierusalem rursumque egressus est ad populum de Bersabee usque ad montem Ephraim et revocavit eos ad Dominum Deum patrum suorum
2CHR|19|5|constituitque iudices terrae in cunctis civitatibus Iuda munitis per singula loca
2CHR|19|6|et praecipiens iudicibus videte ait quid faciatis non enim hominis exercetis iudicium sed Domini et quodcumque iudicaveritis in vos redundabit
2CHR|19|7|sit timor Domini vobiscum et cum diligentia cuncta facite non est enim apud Dominum Deum nostrum iniquitas nec personarum acceptio nec cupido munerum
2CHR|19|8|in Hierusalem quoque constituit Iosaphat Levitas et sacerdotes et principes familiarum ex Israhel ut iudicium et causam Domini iudicarent habitatoribus eius
2CHR|19|9|praecepitque eis dicens sic agetis in timore Dei fideliter et corde perfecto
2CHR|19|10|omnem causam quae venerit ad vos fratrum vestrorum qui habitant in urbibus suis inter cognationem et cognationem ubicumque quaestio est de lege de mandato de caerimoniis de iustificationibus ostendite eis ut non peccent in Dominum et ne veniat ira super vos et super fratres vestros sic ergo agetis et non peccabitis
2CHR|19|11|Amarias autem sacerdos et pontifex vester in his quae ad Dominum pertinent praesidebit porro Zabadias filius Ismahel qui est dux in domo Iuda super ea opera erit quae ad regis officium pertinent habetisque magistros Levitas coram vobis confortamini et agite diligenter et erit Dominus cum bonis
2CHR|20|1|post haec congregati sunt filii Moab et filii Ammon et cum eis de Ammanitis ad Iosaphat ut pugnarent contra eum
2CHR|20|2|veneruntque nuntii et indicaverunt Iosaphat dicentes venit contra te multitudo magna de his locis quae trans mare sunt et de Syria et ecce consistunt in Asasonthamar quae est Engaddi
2CHR|20|3|Iosaphat autem timore perterritus totum se contulit ad rogandum Dominum et praedicavit ieiunium universo Iuda
2CHR|20|4|congregatusque Iudas ad precandum Dominum sed et omnes de urbibus suis venerunt ad obsecrandum eum
2CHR|20|5|cumque stetisset Iosaphat in medio coetu Iudae et Hierusalem in domo Domini ante atrium novum
2CHR|20|6|ait Domine Deus patrum nostrorum tu es Deus in caelo et dominaris cunctis regnis gentium in manu tua est fortitudo et potentia nec quisquam tibi potest resistere
2CHR|20|7|nonne tu Deus noster interfecisti omnes habitatores terrae huius coram populo tuo Israhel et dedisti eam semini Abraham amici tui in sempiternum
2CHR|20|8|habitaveruntque in ea et extruxerunt in illa sanctuarium nomini tuo dicentes
2CHR|20|9|si inruerint super nos mala gladius iudicii pestilentia et fames stabimus coram domo hac in conspectu tuo in qua invocatum est nomen tuum et clamabimus ad te in tribulationibus nostris et exaudies salvosque facies
2CHR|20|10|nunc igitur ecce filii Ammon et Moab et mons Seir per quos non concessisti Israheli ut transirent quando egrediebantur de Aegypto sed declinaverunt ab eis et non interfecerunt illos
2CHR|20|11|e contrario agunt et nituntur eicere nos de possessione quam tradidisti nobis
2CHR|20|12|Deus noster ergo non iudicabis eos in nobis quidem non tanta est fortitudo ut possimus huic multitudini resistere quae inruit super nos sed cum ignoremus quid agere debeamus hoc solum habemus residui ut oculos nostros dirigamus ad te
2CHR|20|13|omnis vero Iuda stabat coram Domino cum parvulis et uxoribus et liberis suis
2CHR|20|14|erat autem Hiazihel filius Zacchariae filii Banaiae filii Hiehihel filii Mathaniae Levites de filiis Asaph super quem factus est spiritus Domini in medio turbae
2CHR|20|15|et ait adtendite omnis Iuda et qui habitatis Hierusalem et tu rex Iosaphat haec dicit Dominus vobis nolite timere nec paveatis hanc multitudinem non est enim vestra pugna sed Dei
2CHR|20|16|cras descendetis contra eos ascensuri enim sunt per clivum nomine Sis et invenietis illos in summitate torrentis qui est contra solitudinem Hieruhel
2CHR|20|17|non eritis vos qui dimicabitis sed tantummodo confidenter state et videbitis auxilium Domini super vos o Iuda et Hierusalem nolite timere nec paveatis cras egredimini contra eos et Dominus erit vobiscum
2CHR|20|18|Iosaphat ergo et Iuda et omnes habitatores Hierusalem ceciderunt proni in terram coram Domino et adoraverunt eum
2CHR|20|19|porro Levitae de filiis Caath et de filiis Core laudabant Dominum Deum Israhel voce magna in excelsum
2CHR|20|20|cumque mane surrexissent egressi sunt per desertum Thecuae profectisque eis stans Iosaphat in medio eorum dixit audite me Iuda et omnes habitatores Hierusalem credite in Domino Deo vestro et securi eritis credite prophetis eius et cuncta evenient prospera
2CHR|20|21|deditque consilium populo et statuit cantores Domini ut laudarent eum in turmis suis et antecederent exercitum ac voce consona dicerent confitemini Domino quoniam in aeternum misericordia eius
2CHR|20|22|cumque coepissent laudes canere vertit Dominus insidias eorum in semet ipsos filiorum scilicet Ammon et Moab et montis Seir qui egressi fuerant ut pugnarent contra Iudam et percussi sunt
2CHR|20|23|namque filii Ammon et Moab consurrexerunt adversum habitatores montis Seir ut interficerent et delerent eos cumque hoc opere perpetrassent etiam in semet ipsos versi mutuis concidere vulneribus
2CHR|20|24|porro Iudas cum venisset ad speculam quae respicit solitudinem vidit procul omnem late regionem plenam cadaveribus nec superesse quemquam qui necem potuisset evadere
2CHR|20|25|venit ergo Iosaphat et omnis populus cum eo ad detrahenda spolia mortuorum inveneruntque inter cadavera variam supellectilem vestes quoque et vasa pretiosissima et diripuerunt ita ut omnia portare non possent nec per tres dies spolia auferre pro praedae magnitudine
2CHR|20|26|die autem quarto congregati sunt in valle Benedictionis etenim quoniam ibi benedixerant Domino vocaverunt locum illum vallis Benedictionis usque in praesentem diem
2CHR|20|27|reversusque est omnis vir Iuda et habitatores Hierusalem et Iosaphat ante eos in Hierusalem cum laetitia magna eo quod dedisset eis Dominus gaudium de inimicis suis
2CHR|20|28|ingressique sunt Hierusalem cum psalteriis et citharis et tubis in domum Domini
2CHR|20|29|inruit autem pavor Domini super universa regna terrarum cum audissent quod pugnasset Dominus contra inimicos Israhel
2CHR|20|30|quievitque regnum Iosaphat et praebuit ei Deus pacem per circuitum
2CHR|20|31|regnavit igitur Iosaphat super Iudam et erat triginta quinque annorum cum regnare coepisset viginti autem et quinque annis regnavit in Hierusalem nomen matris eius Azuba filia Selachi
2CHR|20|32|et ambulavit in via patris sui Asa nec declinavit ab ea faciens quae placita erant coram Domino
2CHR|20|33|verumtamen excelsa non abstulit et adhuc populus non direxerat cor suum ad Dominum Deum patrum suorum
2CHR|20|34|reliqua autem gestorum Iosaphat priorum et novissimorum scripta sunt in verbis Hieu filii Anani quae digessit in libro regum Israhel
2CHR|20|35|post haec iniit amicitias Iosaphat rex Iuda cum Ochozia rege Israhel cuius opera fuerunt impiissima
2CHR|20|36|et particeps fuit ut facerent naves quae irent in Tharsis feceruntque classem in Asiongaber
2CHR|20|37|prophetavit autem Eliezer filius Dodoau de Maresa ad Iosaphat dicens quia habuisti foedus cum Ochozia percussit Dominus opera tua contritaeque sunt naves nec potuerunt ire in Tharsis
2CHR|21|1|dormivit autem Iosaphat cum patribus suis et sepultus est cum eis in civitate David regnavitque Ioram filius eius pro eo
2CHR|21|2|qui habuit fratres filios Iosaphat Azariam et Hiahihel et Zacchariam et Azariam et Michahel et Saphatiam omnes hii filii Iosaphat regis Israhel
2CHR|21|3|deditque eis pater suus multa munera argenti et auri et pensitationes cum civitatibus munitissimis in Iuda regnum autem tradidit Ioram eo quod esset primogenitus
2CHR|21|4|surrexit ergo Ioram super regnum patris sui cumque se confirmasset occidit omnes fratres suos gladio et quosdam de principibus Israhel
2CHR|21|5|triginta duo annorum erat Ioram cum regnare coepisset et octo annis regnavit in Hierusalem
2CHR|21|6|ambulavitque in viis regum Israhel sicut egerat domus Ahab filia quippe Ahab erat uxor eius et fecit malum in conspectu Domini
2CHR|21|7|noluit autem Dominus disperdere domum David propter pactum quod inierat cum eo et quia promiserat ut daret illi lucernam et filiis eius omni tempore
2CHR|21|8|in diebus illis rebellavit Edom ne esset subditus Iudae et constituit sibi regem
2CHR|21|9|cumque transisset Ioram cum principibus suis et cuncto equitatu qui erat secum surrexit nocte et percussit Edom qui se circumdederat et omnes duces equitatus eius
2CHR|21|10|attamen rebellavit Edom ne esset sub dicione Iuda usque ad hanc diem eo tempore et Lobna recessit ne esset sub manu illius dereliquerat enim Dominum Deum patrum suorum
2CHR|21|11|insuper et excelsa fabricatus est in urbibus Iuda et fornicari fecit habitatores Hierusalem et praevaricari Iudam
2CHR|21|12|adlatae sunt autem ei litterae ab Helia propheta in quibus scriptum erat haec dicit Dominus Deus David patris tui quoniam non ambulasti in viis Iosaphat patris tui et in viis Asa regis Iuda
2CHR|21|13|sed incessisti per iter regum Israhel et fornicari fecisti Iudam et habitatores Hierusalem imitatus fornicationem domus Ahab insuper et fratres tuos domum patris tui meliores te occidisti
2CHR|21|14|ecce Dominus percutiet te plaga magna cum populo tuo et filiis et uxoribus tuis universaque substantia tua
2CHR|21|15|tu autem aegrotabis pessimo languore uteri donec egrediantur vitalia tua paulatim per dies singulos
2CHR|21|16|suscitavit ergo Dominus contra Ioram spiritum Philisthinorum et Arabum qui confines sunt Aethiopibus
2CHR|21|17|et ascenderunt in terram Iuda et vastaverunt eam diripueruntque cunctam substantiam quae inventa est in domo regis insuper et filios eius et uxores nec remansit ei filius nisi Ioachaz qui minimus natu erat
2CHR|21|18|et super haec omnia percussit eum Dominus alvi languore insanabili
2CHR|21|19|cumque diei succederet dies et temporum spatia volverentur duorum annorum expletus est circulus et sic longa consumptus tabe ita ut egereret etiam viscera sua languore pariter et vita caruit mortuusque est in infirmitate pessima et non fecit ei populus secundum morem conbustionis exequias sicut fecerat maioribus eius
2CHR|21|20|triginta duum annorum fuit cum regnare coepisset et octo annis regnavit in Hierusalem ambulavitque non recte et sepelierunt eum in civitate David verumtamen non in sepulchro regum
2CHR|22|1|constituerunt autem habitatores Hierusalem Ochoziam filium eius minimum regem pro eo omnes enim maiores natu qui ante eum fuerant interfecerant latrones Arabum qui inruerant in castra regnavitque Ochozias filius Ioram regis Iuda
2CHR|22|2|filius quadraginta duo annorum erat Ochozias cum regnare coepisset et uno anno regnavit in Hierusalem nomen matris eius Otholia filia Amri
2CHR|22|3|sed et ipse ingressus est per vias domus Ahab mater enim eius inpulit eum ut impie ageret
2CHR|22|4|fecit igitur malum in conspectu Domini sicut domus Ahab ipsi enim fuerunt ei consiliarii post mortem patris sui in interitum eius
2CHR|22|5|ambulavitque in consiliis eorum et perrexit cum Ioram filio Ahab rege Israhel in bellum contra Azahel regem Syriae in Ramoth Galaad vulneraveruntque Syri Ioram
2CHR|22|6|qui reversus est ut curaretur in Hiezrahel multas enim plagas acceperat in supradicto certamine igitur Azarias filius Ioram rex Iuda descendit ut inviseret Ioram filium Ahab in Hiezrahel aegrotantem
2CHR|22|7|voluntatis quippe fuit Dei adversum Ochoziam ut veniret ad Ioram et cum venisset egrederetur cum eo adversum Hieu filium Namsi quem unxit Dominus ut deleret domum Ahab
2CHR|22|8|cum ergo subverteret Hieu domum Ahab invenit principes Iuda et filios fratrum Ochoziae qui ministrabant ei et interfecit illos
2CHR|22|9|ipsumque perquirens Ochoziam conprehendit latentem in Samaria adductumque ad se occidit et sepelierunt eum eo quod esset filius Iosaphat qui quaesierat Dominum in toto corde suo nec erat ultra spes aliqua ut de stirpe regnaret Ochoziae
2CHR|22|10|siquidem Otholia mater eius videns quod mortuus esset filius suus surrexit et interfecit omnem stirpem regiam domus Ioram
2CHR|22|11|porro Iosabeth filia regis tulit Ioas filium Ochoziae et furata est eum de medio filiorum regis cum interficerentur absconditque cum nutrice sua in cubiculo lectulorum Iosabeth autem quae absconderat eum erat filia regis Ioram uxor Ioiadae pontificis soror Ochoziae et idcirco Otholia non interfecit eum
2CHR|22|12|fuit ergo cum eis in domo Dei absconditus sex annis quibus regnavit Otholia super terram
2CHR|23|1|anno autem septimo confortatus Ioiadae adsumpsit centuriones Azariam videlicet filium Hieroam et Ismahel filium Iohanan Azariam quoque filium Oded et Maasiam filium Adaiae et Elisaphat filium Zechri et iniit cum eis foedus
2CHR|23|2|qui circumeuntes Iudam congregaverunt Levitas de cunctis urbibus Iuda et principes familiarum Israhel veneruntque in Hierusalem
2CHR|23|3|iniit igitur omnis multitudo pactum in domo Domini cum rege dixitque ad eos Ioiadae ecce filius regis regnabit sicut locutus est Dominus super filios David
2CHR|23|4|iste est ergo sermo quem facietis
2CHR|23|5|tertia pars vestrum qui veniunt ad sabbatum sacerdotum et Levitarum et ianitorum erit in portis tertia vero pars ad domum regis et tertia in porta quae appellatur Fundamenti omne vero reliquum vulgus sit in atriis domus Domini
2CHR|23|6|nec quisquam alius ingrediatur domum Domini nisi sacerdotes et qui ministrant de Levitis ipsi tantummodo ingrediantur quia sanctificati sunt et omne reliquum vulgus observet custodias Domini
2CHR|23|7|Levitae autem circumdent regem habentes singuli arma sua et si quis alius ingressus fuerit templum interficiatur sintque cum rege et intrante et egrediente
2CHR|23|8|fecerunt igitur Levitae et universus Iuda iuxta omnia quae praeceperat Ioiadae pontifex et adsumpserunt singuli viros qui sub se erant et veniebant per ordinem sabbati cum his qui iam impleverant sabbatum et egressuri erant siquidem Ioiadae pontifex non dimiserat abire turmas quae sibi per singulas ebdomadas succedere consueverant
2CHR|23|9|deditque Ioiadae sacerdos centurionibus lanceas clypeosque et peltas regis David quas consecraverat in domo Domini
2CHR|23|10|constituitque omnem populum tenentium pugiones a parte templi dextra usque ad partem templi sinistram coram altari et templo per circuitum regis
2CHR|23|11|et eduxerunt filium regis et inposuerunt ei diadema dederuntque in manu eius tenendam legem et constituerunt eum regem unxit quoque illum Ioiadae pontifex et filii eius inprecatique sunt atque dixerunt vivat rex
2CHR|23|12|quod cum audisset Otholia vocem scilicet currentium atque laudantium regem ingressa est ad populum in templum Domini
2CHR|23|13|cumque vidisset regem stantem super gradum in introitu et principes turmasque circa eum omnem quoque populum terrae gaudentem atque clangentem tubis et diversi generis organis concinentem vocemque laudantium scidit vestimenta sua et ait insidiae insidiae
2CHR|23|14|egressus autem Ioiadae pontifex ad centuriones et principes exercitus dixit eis educite illam extra septa templi et interficiatur foris gladio praecepitque sacerdos ne occideretur in domo Domini
2CHR|23|15|et inposuerunt cervicibus eius manus cumque intrasset portam Equorum domus regis interfecerunt eam ibi
2CHR|23|16|pepigit autem Ioiadae foedus inter se universumque populum et regem ut esset populus Domini
2CHR|23|17|itaque ingressus est omnis populus domum Baal et destruxerunt eam et altaria ac simulacra illius confregerunt Matthan quoque sacerdotem Baal interfecerunt ante aras
2CHR|23|18|constituit autem Ioiadae praepositos in domo Domini et sub manibus sacerdotum ac Levitarum quos distribuit David in domo Domini ut offerrent holocausta Domino sicut scriptum est in lege Mosi in gaudio et canticis iuxta dispositionem David
2CHR|23|19|constituit quoque ianitores in portis domus Domini ut non ingrederetur eam inmundus in omni re
2CHR|23|20|adsumpsitque centuriones et fortissimos viros ac principes populi et omne vulgus terrae et fecerunt descendere regem de domo Domini et introire per medium portae superioris in domum regis et conlocaverunt eum in solio regali
2CHR|23|21|laetatusque est omnis populus terrae et urbs quievit porro Otholia interfecta est gladio
2CHR|24|1|septem annorum erat Ioas cum regnare coepisset et quadraginta annis regnavit in Hierusalem nomen matris eius Sebia de Bersabee
2CHR|24|2|fecitque quod bonum est coram Domino cunctis diebus Ioiadae sacerdotis
2CHR|24|3|accepit autem ei Ioiadae uxores duas e quibus genuit filios et filias
2CHR|24|4|post quae placuit Ioas ut instauraret domum Domini
2CHR|24|5|congregavitque sacerdotes et Levitas et dixit eis egredimini ad civitates Iuda et colligite de universo Israhel pecuniam ad sarta tecta templi Dei vestri per singulos annos festinatoque hoc facite porro Levitae egere neglegentius
2CHR|24|6|vocavitque rex Ioiadae principem et dixit ei quare non tibi fuit curae ut cogeres Levitas inferre de Iuda et de Hierusalem pecuniam quae constituta est a Mose servo Domini ut inferret eam omnis multitudo Israhel in tabernaculum testimonii
2CHR|24|7|Otholia enim impiissima et filii eius destruxerunt domum Domini et de universis quae sanctificata fuerant templo Domini ornaverunt fanum Baalim
2CHR|24|8|praecepit ergo rex et fecerunt arcam posueruntque eam iuxta portam domus Domini forinsecus
2CHR|24|9|et praedicatum est in Iuda et Hierusalem ut deferrent singuli pretium Domino quod constituit Moses servus Dei super omnem Israhel in deserto
2CHR|24|10|laetatique sunt cuncti principes et omnis populus et ingressi contulerunt in arcam Domini atque miserunt ita ut impleretur
2CHR|24|11|cumque tempus esset ut deferrent arcam coram rege per manus Levitarum videbant enim multam pecuniam ingrediebatur scriba regis et quem primus sacerdos constituerat effundebantque pecuniam quae erat in arca porro arcam reportabant ad locum suum sicque faciebant per singulos dies et congregata est infinita pecunia
2CHR|24|12|quam dederunt rex et Ioiada his qui praeerant operibus domus Domini at illi conducebant ex ea caesores lapidum et artifices operum singulorum ut instaurarent domum Domini fabros quoque ferri et aeris ut quod cadere coeperat fulciretur
2CHR|24|13|egeruntque hii qui operabantur industrie et obducebatur parietum cicatrix per manus eorum ac suscitaverunt domum Domini in statum pristinum et firme eam stare fecerunt
2CHR|24|14|cumque conplessent omnia opera detulerunt coram rege et Ioiadae reliquam partem pecuniae de qua facta sunt vasa templi in ministerium et ad holocausta fialae quoque et cetera vasa aurea et argentea et offerebantur holocausta in domo Domini iugiter cunctis diebus Ioiadae
2CHR|24|15|senuit autem Ioiadae plenus dierum et mortuus est cum centum triginta esset annorum
2CHR|24|16|sepelieruntque eum in civitate David cum regibus eo quod fecisset bonum cum Israhel et cum domo eius
2CHR|24|17|postquam autem obiit Ioiada ingressi sunt principes Iuda et adoraverunt regem qui delinitus obsequiis eorum adquievit eis
2CHR|24|18|et dereliquerunt templum Domini Dei patrum suorum servieruntque lucis et sculptilibus et facta est ira contra Iudam et Hierusalem propter hoc peccatum
2CHR|24|19|mittebatque eis prophetas ut reverterentur ad Dominum quos protestantes illi audire nolebant
2CHR|24|20|spiritus itaque Dei induit Zacchariam filium Ioiadae sacerdotem et stetit in conspectu populi et dixit eis haec dicit Dominus quare transgredimini praeceptum Domini quod vobis non proderit et dereliquistis Dominum ut derelinqueret vos
2CHR|24|21|qui congregati adversus eum miserunt lapides iuxta regis imperium in atrio domus Domini
2CHR|24|22|et non est recordatus Ioas rex misericordiae quam fecerat Ioiadae pater illius secum sed interfecit filium eius qui cum moreretur ait videat Dominus et requirat
2CHR|24|23|cumque evolutus esset annus ascendit contra eum exercitus Syriae venitque in Iudam et Hierusalem et interfecit cunctos principes populi atque universam praedam miserunt regi Damascum
2CHR|24|24|et certe cum permodicus venisset numerus Syrorum tradidit Dominus manibus eorum infinitam multitudinem eo quod reliquissent Dominum Deum patrum suorum in Ioas quoque ignominiosa exercuere iudicia
2CHR|24|25|et abeuntes dimiserunt eum in languoribus magnis surrexerunt autem contra eum servi sui in ultionem sanguinis filii Ioiadae sacerdotis et occiderunt eum in lectulo suo et mortuus est sepelieruntque eum in civitate David sed non in sepulchris regum
2CHR|24|26|insidiati vero sunt ei Zabath filius Semath Ammanitidis et Iozabath filius Semarith Moabitidis
2CHR|24|27|porro filii eius ac summa pecuniae quae adunata fuerat sub eo et instauratio domus Dei scripta sunt diligentius in libro regum regnavitque Amasias filius eius pro eo
2CHR|25|1|viginti quinque annorum erat Amasias cum regnare coepisset et viginti novem annis regnavit in Hierusalem nomen matris eius Ioaden de Hierusalem
2CHR|25|2|fecitque bonum in conspectu Domini verumtamen non in corde perfecto
2CHR|25|3|cumque roboratum sibi videret imperium iugulavit servos qui occiderant regem patrem suum
2CHR|25|4|sed filios eorum non interfecit sicut scriptum est in libro legis Mosi ubi praecepit Dominus dicens non occidentur patres pro filiis neque filii pro patribus suis sed unusquisque in suo peccato morietur
2CHR|25|5|congregavit igitur Amasias Iudam et constituit eos per familias tribunosque et centuriones in universo Iuda et Beniamin et recensuit a viginti annis sursum invenitque triginta milia iuvenum qui egrederentur ad pugnam et tenerent hastam et clypeum
2CHR|25|6|mercede quoque conduxit de Israhel centum milia robustorum centum talentis argenti
2CHR|25|7|venit autem homo Dei ad illum et ait o rex ne egrediatur tecum exercitus Israhel non est enim Dominus cum Israhel et cunctis filiis Ephraim
2CHR|25|8|quod si putas in robore exercitus bella consistere superari te faciet Deus ab hostibus Dei quippe est et adiuvare et in fugam vertere
2CHR|25|9|dixitque Amasias ad hominem Dei quid ergo fiet de centum talentis quae dedi militibus Israhel et respondit ei homo Dei habet Dominus unde tibi dare possit multo his plura
2CHR|25|10|separavit itaque Amasias exercitum qui venerat ad eum ex Ephraim ut reverteretur in locum suum at illi contra Iudam vehementer irati reversi sunt in regionem suam
2CHR|25|11|porro Amasias confidenter eduxit populum suum et abiit in vallem Salinarum percussitque filios Seir decem milia
2CHR|25|12|et alia decem milia virorum ceperunt filii Iuda et adduxerunt ad praeruptum cuiusdam petrae praecipitaveruntque eos de summo in praeceps qui universi crepuerunt
2CHR|25|13|at ille exercitus quem remiserat Amasias ne secum iret ad proelium diffusus est in civitatibus Iuda a Samaria usque Bethoron et interfectis tribus milibus diripuit praedam magnam
2CHR|25|14|Amasias vero post caedem Idumeorum et adlatos deos filiorum Seir statuit illos in deos sibi et adorabat eos et illis adolebat incensum
2CHR|25|15|quam ob rem iratus Dominus contra Amasiam misit ad illum prophetam qui diceret ei cur adorasti deos qui non liberaverunt populum suum de manu tua
2CHR|25|16|cumque haec ille loqueretur respondit ei num consiliarius regis es quiesce ne interficiam te discedensque propheta scio inquit quod cogitaverit Dominus occidere te qui et fecisti hoc malum et insuper non adquievisti consilio meo
2CHR|25|17|igitur Amasias rex Iuda inito pessimo consilio misit ad Ioas filium Ioachaz filii Hieu regem Israhel dicens veni videamus nos mutuo
2CHR|25|18|at ille remisit nuntium dicens carduus qui est in Libano misit ad cedrum Libani dicens da filiam tuam filio meo uxorem et ecce bestiae quae erant in silva Libani transierunt et conculcaverunt carduum
2CHR|25|19|dixisti percussi Edom et idcirco erigitur cor tuum in superbiam sede in domo tua cur malum adversum te provocas ut cadas et tu et Iudas tecum
2CHR|25|20|noluit audire Amasias eo quod Domini esset voluntas ut traderetur in manibus hostium propter deos Edom
2CHR|25|21|ascendit igitur Ioas rex Israhel et mutuos sibi praebuere conspectus Amasias autem rex Iuda erat in Bethsames Iudae
2CHR|25|22|corruitque Iudas coram Israhel et fugit in tabernacula sua
2CHR|25|23|porro Amasiam regem Iuda filium Ioas filii Ioachaz cepit Ioas rex Israhel in Bethsames et adduxit in Hierusalem destruxitque murum eius a porta Ephraim usque ad portam Anguli quadringentis cubitis
2CHR|25|24|omne quoque aurum et argentum et universa vasa quae reppererat in domo Dei et apud Obededom in thesauris etiam domus regiae necnon et filios obsidum reduxit Samariam
2CHR|25|25|vixit autem Amasias filius Ioas rex Iuda postquam mortuus est Ioas filius Ioachaz rex Israhel quindecim annis
2CHR|25|26|reliqua vero sermonum Amasiae priorum et novissimorum scripta sunt in libro regum Iuda et Israhel
2CHR|25|27|qui postquam recessit a Domino tetenderunt ei insidias in Hierusalem cumque fugisset Lachis miserunt et interfecerunt eum ibi
2CHR|25|28|reportantesque super equos sepelierunt eum cum patribus suis in civitate David
2CHR|26|1|omnis autem populus Iuda filium eius Oziam annorum sedecim constituit regem pro patre suo Amasia
2CHR|26|2|ipse aedificavit Ahilath et restituit eam dicioni Iudae postquam dormivit rex cum patribus suis
2CHR|26|3|sedecim annorum erat Ozias cum regnare coepisset et quinquaginta duobus annis regnavit in Hierusalem nomen matris eius Hiechelia de Hierusalem
2CHR|26|4|fecitque quod erat rectum in oculis Domini iuxta omnia quae fecerat Amasias pater eius
2CHR|26|5|et exquisivit Deum in diebus Zacchariae intellegentis et videntis Deum cumque requireret Dominum direxit eum in omnibus
2CHR|26|6|denique egressus est et pugnavit contra Philisthim et destruxit murum Geth et murum Iabniae murumque Azoti aedificavit quoque oppida in Azoto et in Philisthim
2CHR|26|7|et adiuvit eum Deus contra Philisthim et contra Arabas qui habitabant in Gurbaal et contra Ammanitas
2CHR|26|8|pendebantque Ammanitae munera Oziae et divulgatum est nomen eius usque ad introitum Aegypti propter crebras victorias
2CHR|26|9|aedificavitque Ozias turres in Hierusalem super portam Anguli et super portam Vallis et reliquas in eodem muri latere firmavitque eas
2CHR|26|10|extruxit etiam turres in solitudine et fodit cisternas plurimas eo quod haberet multa pecora tam in campestribus quam in heremi vastitate vineas quoque habuit et vinitores in montibus et in Carmelo erat quippe homo agriculturae deditus
2CHR|26|11|fuit autem exercitus bellatorum eius qui procedebant ad proelia sub manu Hiehihel scribae Maasiaeque doctoris et sub manu Ananiae qui erat de ducibus regis
2CHR|26|12|omnisque numerus principum per familias virorum fortium duum milium sescentorum
2CHR|26|13|et sub eis universus exercitus trecentorum et septem milium quingentorum qui erant apti ad bella et pro rege contra adversarios dimicabant
2CHR|26|14|praeparavit quoque eis Ozias id est cuncto exercitui clypeos et hastas et galeas et loricas arcusque et fundas ad iaciendos lapides
2CHR|26|15|et fecit in Hierusalem diversi generis machinas quas in turribus conlocavit et in angulis murorum ut mitterent sagittas et saxa grandia egressumque est nomen eius procul eo quod auxiliaretur ei Dominus et corroborasset illum
2CHR|26|16|sed cum roboratus esset elevatum est cor eius in interitum suum et neglexit Dominum Deum suum ingressusque templum Domini adolere voluit incensum super altare thymiamatis
2CHR|26|17|statimque ingressus post eum Azarias sacerdos et cum eo sacerdotes Domini octoginta viri fortissimi
2CHR|26|18|restiterunt regi atque dixerunt non est tui officii Ozia ut adoleas incensum Domino sed sacerdotum hoc est filiorum Aaron qui consecrati sunt ad huiuscemodi ministerium egredere de sanctuario ne contempseris quia non reputabitur tibi in gloriam hoc a Domino Deo
2CHR|26|19|iratusque est Ozias et tenens in manu turibulum ut adoleret incensum minabatur sacerdotibus statimque orta est lepra in fronte eius coram sacerdotibus in domo Domini super altare thymiamatis
2CHR|26|20|cumque respexisset eum Azarias pontifex et omnes reliqui sacerdotes viderunt lepram in fronte eius et festinato expulerunt eum sed et ipse perterritus adceleravit egredi eo quod sensisset ilico plagam Domini
2CHR|26|21|fuit igitur Ozias rex leprosus usque ad diem mortis suae et habitavit in domo separata plenus lepra ob quam et eiectus fuerat de domo Domini porro Ioatham filius eius rexit domum regis et iudicabat populum terrae
2CHR|26|22|reliqua autem sermonum Oziae priorum et novissimorum scripsit Esaias filius Amos propheta
2CHR|26|23|dormivitque Ozias cum patribus suis et sepelierunt eum in agro regalium sepulchrorum eo quod esset leprosus regnavitque Ioatham filius eius pro eo
2CHR|27|1|viginti quinque annorum erat Ioatham cum regnare coepisset et sedecim annis regnavit in Hierusalem nomen matris eius Hierusa filia Sadoc
2CHR|27|2|fecitque quod rectum erat coram Domino iuxta omnia quae fecerat Ozias pater suus excepto quod non est ingressus templum Domini et adhuc populus delinquebat
2CHR|27|3|ipse aedificavit portam domus Domini Excelsam et in muro Ophel multa construxit
2CHR|27|4|urbes quoque aedificavit in montibus Iuda et in saltibus castella et turres
2CHR|27|5|ipse pugnavit contra regem filiorum Ammon et vicit eos dederuntque ei filii Ammon in tempore illo centum talenta argenti et decem milia choros tritici ac totidem choros hordei haec ei praebuerunt filii Ammon in anno secundo et tertio
2CHR|27|6|corroboratusque est Ioatham eo quod direxisset vias suas coram Domino Deo suo
2CHR|27|7|reliqua autem sermonum Ioatham et omnes pugnae eius et opera scripta sunt in libro regum Israhel et Iuda
2CHR|27|8|viginti quinque annorum erat cum regnare coepisset et sedecim annis regnavit in Hierusalem
2CHR|27|9|dormivitque Ioatham cum patribus suis et sepelierunt eum in civitate David et regnavit Achaz filius eius pro eo
2CHR|28|1|viginti annorum erat Achaz cum regnare coepisset et sedecim annis regnavit in Hierusalem non fecit rectum in conspectu Domini sicut David pater eius
2CHR|28|2|sed ambulavit in viis regum Israhel insuper et statuas fudit Baalim
2CHR|28|3|ipse est qui adolevit incensum in valle Benennon et lustravit filios suos in igne iuxta ritum gentium quas interfecit Dominus in adventu filiorum Israhel
2CHR|28|4|sacrificabat quoque et thymiama succendebat in excelsis et in collibus et sub omni ligno frondoso
2CHR|28|5|tradiditque eum Dominus Deus eius in manu regis Syriae qui percussit eum magnamque praedam de eius cepit imperio et adduxit in Damascum manibus quoque regis Israhel traditus est et percussus plaga grandi
2CHR|28|6|occiditque Phacee filius Romeliae de Iuda centum viginti milia in die uno omnes viros bellatores eo quod reliquissent Dominum Deum patrum suorum
2CHR|28|7|eodem tempore occidit Zechri vir potens ex Ephraim Masiam filium regis et Ezricam ducem domus eius Helcanam quoque secundum a rege
2CHR|28|8|ceperuntque filii Israhel de fratribus suis ducenta milia mulierum puerorum et puellarum et infinitam praedam pertuleruntque eam in Samariam
2CHR|28|9|ea tempestate erat ibi propheta Domini nomine Oded qui egressus obviam exercitui venientium in Samariam dixit eis ecce iratus Dominus Deus patrum vestrorum contra Iudam tradidit eos manibus vestris et occidistis illos atrociter ita ut caelum pertingeret vestra crudelitas
2CHR|28|10|insuper filios Iuda et Hierusalem vultis vobis subicere in servos et ancillas quod nequaquam facto opus est peccatis enim super hoc Domino Deo vestro
2CHR|28|11|sed audite consilium meum et reducite captivos quos adduxistis de fratribus vestris quia magnus furor Domini inminet vobis
2CHR|28|12|steterunt itaque viri de principibus filiorum Ephraim Azarias filius Iohanan Barachias filius Mosollamoth Hiezechias filius Sellum et Amasa filius Adali contra eos qui veniebant de proelio
2CHR|28|13|et dixerunt eis non introducetis huc captivos ne peccemus Domino quare vultis adicere super peccata nostra et vetera cumulare delicta grande quippe peccatum est et ira furoris Domini inminet super Israhel
2CHR|28|14|dimiseruntque viri bellatores praedam et universa quae ceperant coram principibus et omni multitudine
2CHR|28|15|steteruntque viri quos supra memoravimus et adprehendentes captivos omnesque qui nudi erant vestierunt de spoliis cumque vestissent eos et calciassent et refecissent cibo ac potu unxissent quoque propter laborem et adhibuissent eis curam quicumque ambulare non poterant et erant inbecillo corpore inposuerunt eos iumentis et adduxerunt Hierichum civitatem Palmarum ad fratres eorum ipsique reversi sunt Samariam
2CHR|28|16|tempore illo misit rex Achaz ad regem Assyriorum auxilium postulans
2CHR|28|17|veneruntque Idumei et percusserunt multos ex Iuda et ceperunt praedam magnam
2CHR|28|18|Philisthim quoque diffusi sunt per urbes campestres et ad meridiem Iuda ceperuntque Bethsames et Ahilon et Gaderoth Soccho quoque et Thamnam et Gamzo cum viculis suis et habitaverunt in eis
2CHR|28|19|humiliaverat enim Dominus Iudam propter Achaz regem Iuda eo quod nudasset eum auxilio et contemptui habuisset Dominum
2CHR|28|20|adduxitque contra eum Thaglathphalnasar regem Assyriorum qui et adflixit eum et nullo resistente vastavit
2CHR|28|21|igitur Achaz spoliata domo Domini et domo regum et principum dedit regi Assyriorum munera et tamen nihil ei profuit
2CHR|28|22|insuper et in tempore angustiae suae auxit contemptum in Dominum ipse per se rex Achaz
2CHR|28|23|immolavit diis Damasci victimas percussoribus suis et dixit dii regum Syriae auxiliantur eis quos ego placabo hostiis et aderunt mihi cum e contrario ipsi fuerint ruina eius et universo Israhel
2CHR|28|24|direptis itaque Achaz omnibus vasis domus Dei atque confractis clusit ianuas templi Dei et fecit sibi altaria in universis angulis Hierusalem
2CHR|28|25|in omnibus quoque urbibus Iuda extruxit aras ad cremandum tus atque ad iracundiam provocavit Dominum Deum patrum suorum
2CHR|28|26|reliqua autem sermonum eius et omnium operum priorum et novissimorum scripta sunt in libro regum Iuda et Israhel
2CHR|28|27|dormivitque Achaz cum patribus suis et sepelierunt eum in civitate Hierusalem neque enim receperunt eum in sepulchra regum Israhel regnavitque Ezechias filius eius pro eo
2CHR|29|1|igitur Ezechias regnare coepit cum viginti quinque esset annorum et viginti novem annis regnavit in Hierusalem nomen matris eius Abia filia Zacchariae
2CHR|29|2|fecitque quod erat placitum in conspectu Domini iuxta omnia quae fecerat David pater eius
2CHR|29|3|ipse anno et mense primo regni sui aperuit valvas domus Domini et instauravit eas
2CHR|29|4|adduxitque sacerdotes atque Levitas et congregavit eos in plateam orientalem
2CHR|29|5|dixitque ad eos audite me Levitae et sanctificamini mundate domum Domini Dei patrum vestrorum auferte omnem inmunditiam de sanctuario
2CHR|29|6|peccaverunt patres nostri et fecerunt malum in conspectu Domini Dei nostri derelinquentes eum averterunt facies suas a tabernaculo Domini et praebuerunt dorsum
2CHR|29|7|cluserunt ostia quae erant in porticu et extinxerunt lucernas incensumque non adoleverunt et holocausta non obtulerunt in sanctuario Deo Israhel
2CHR|29|8|concitatus est itaque furor Domini super Iudam et Hierusalem tradiditque eos in commotionem et in interitum et in sibilum sicut ipsi cernitis oculis vestris
2CHR|29|9|en corruerunt patres nostri gladiis filii nostri et filiae nostrae et coniuges captivae ductae sunt propter hoc scelus
2CHR|29|10|nunc igitur placet mihi ut ineamus foedus cum Domino Deo Israhel et avertat a nobis furorem irae suae
2CHR|29|11|filii mi nolite neglegere vos elegit Dominus ut stetis coram eo et ministretis illi colatis eum et cremetis incensum
2CHR|29|12|surrexerunt ergo Levitae Maath filius Amasiae et Iohel filius Azariae de filiis Caath porro de filiis Merari Cis filius Abdai et Azarias filius Iallelel de filiis autem Gersom Ioha filius Zemma et Eden filius Ioaha
2CHR|29|13|at vero de filiis Elisaphan Samri et Iahihel de filiis quoque Asaph Zaccharias et Mathanias
2CHR|29|14|necnon de filiis Heman Iahihel et Semei sed et de filiis Idithun Semeias et Ozihel
2CHR|29|15|congregaveruntque fratres suos et sanctificati sunt et ingressi iuxta mandatum regis et imperium Domini ut expiarent domum Dei
2CHR|29|16|sacerdotes quoque ingressi templum Domini ut sanctificarent illud extulerunt omnem inmunditiam quam intro reppererant in vestibulum domus Domini quam tulerunt Levitae et asportaverunt ad torrentem Cedron foras
2CHR|29|17|coeperunt autem prima die mensis primi mundare et in die octava eiusdem mensis ingressi sunt porticum templi Domini expiaveruntque templum diebus octo et in die sextadecima mensis eiusdem quod coeperant impleverunt
2CHR|29|18|ingressi quoque sunt ad Ezechiam regem et dixerunt ei sanctificavimus omnem domum Domini et altare holocaustoseos vasaque eius necnon et mensam propositionis cum omnibus vasis suis
2CHR|29|19|cunctamque templi supellectilem quam polluerat rex Achaz in regno suo postquam praevaricatus est et ecce exposita sunt omnia coram altari Domini
2CHR|29|20|consurgensque diluculo Ezechias rex adunavit omnes principes civitatis et ascendit domum Domini
2CHR|29|21|obtuleruntque simul tauros septem arietes septem agnos septem et hircos septem pro peccato pro regno pro sanctuario pro Iuda dixit quoque sacerdotibus filiis Aaron ut offerrent super altare Domini
2CHR|29|22|mactaverunt igitur tauros et susceperunt sacerdotes sanguinem et fuderunt illud super altare mactaverunt etiam arietes et illorum sanguinem super altare fuderunt immolaverunt agnos et fuderunt super altare sanguinem
2CHR|29|23|adplicaverunt hircos pro peccato coram rege et universa multitudine inposueruntque manus suas super eos
2CHR|29|24|et immolaverunt illos sacerdotes et asperserunt sanguinem eorum altari pro piaculo universi Israhelis pro omni quippe Israhel praeceperat rex ut holocaustum fieret et pro peccato
2CHR|29|25|constituit quoque Levitas in domo Domini cum cymbalis et psalteriis et citharis secundum dispositionem David et Gad videntis regis et Nathan prophetae siquidem Domini praeceptum fuit per manum prophetarum eius
2CHR|29|26|steteruntque Levitae tenentes organa David et sacerdotes tubas
2CHR|29|27|et iussit Ezechias ut offerrent holocaustum super altare cumque offerrentur holocausta coeperunt laudes canere Domino et clangere tubis atque in diversis organis quae David rex Israhel reppererat concrepare
2CHR|29|28|omni autem turba adorante cantores et hii qui tenebant tubas erant in officio suo donec conpleretur holocaustum
2CHR|29|29|cumque finita esset oblatio incurvatus est rex et omnes qui erant cum eo et adoraverunt
2CHR|29|30|praecepitque Ezechias et principes Levitis ut laudarent Dominum sermonibus David et Asaph videntis qui laudaverunt eum magna laetitia et curvato genu adoraverunt
2CHR|29|31|Ezechias autem etiam haec addidit implestis manus vestras Domino accedite et offerte victimas et laudes in domo Domini obtulit ergo universa multitudo hostias et laudes et holocausta mente devota
2CHR|29|32|porro numerus holocaustorum quae obtulit multitudo hic fuit tauros septuaginta arietes centum agnos ducentos
2CHR|29|33|sanctificaveruntque Domino boves sescentos et oves tria milia
2CHR|29|34|sacerdotes vero pauci erant nec poterant sufficere ut pelles holocaustorum detraherent unde et Levitae fratres eorum adiuverunt eos donec impleretur opus et sanctificarentur antistites Levitae quippe faciliori ritu sanctificantur quam sacerdotes
2CHR|29|35|fuerunt igitur holocausta plurima adipes pacificorum et libamina holocaustorum et conpletus est cultus domus Domini
2CHR|29|36|laetatusque est Ezechias et omnis populus eo quod ministerium Domini esset expletum de repente quippe hoc fieri placuerat
2CHR|30|1|misit quoque Ezechias ad omnem Israhel et Iudam scripsitque epistulas ad Ephraim et Manassem ut venirent ad domum Domini in Hierusalem et facerent phase Domino Deo Israhel
2CHR|30|2|inito ergo consilio regis et principum et universi coetus Hierusalem decreverunt ut facerent phase mense secundo
2CHR|30|3|non enim occurrerant facere in tempore suo quia sacerdotes qui possent sufficere sanctificati non fuerant et populus necdum congregatus erat in Hierusalem
2CHR|30|4|placuitque sermo regi et omni multitudini
2CHR|30|5|et decreverunt ut mitterent nuntios in universum Israhel de Bersabee usque Dan ut venirent et facerent phase Domino Deo Israhel in Hierusalem multi enim non fecerant sicut lege praescriptum est
2CHR|30|6|perrexeruntque cursores cum epistulis ex regis imperio et principum eius in universum Israhel et Iudam iuxta quod rex iusserat praedicantes filii Israhel revertimini ad Dominum Deum Abraham et Isaac et Israhel et revertetur ad reliquias quae effugerunt manum regis Assyriorum
2CHR|30|7|nolite fieri sicut patres vestri et fratres qui recesserunt a Domino Deo patrum suorum et tradidit eos in interitum ut ipsi cernitis
2CHR|30|8|nolite indurare cervices vestras sicut patres vestri tradite manus Domino et venite ad sanctuarium eius quod sanctificavit in aeternum servite Domino Deo patrum vestrorum et avertetur a vobis ira furoris eius
2CHR|30|9|si enim vos reversi fueritis ad Dominum fratres vestri et filii habebunt misericordiam coram dominis suis qui illos duxere captivos et revertentur in terram hanc pius enim et clemens est Dominus Deus vester et non avertet faciem suam a vobis si reversi fueritis ad eum
2CHR|30|10|igitur cursores pergebant velociter de civitate in civitatem per terram Ephraim et Manasse usque Zabulon illis inridentibus et subsannantibus eos
2CHR|30|11|attamen quidam viri ex Aser et Manasse et Zabulon adquiescentes consilio venerunt Hierusalem
2CHR|30|12|in Iuda vero facta est manus Domini ut daret eis cor unum et facerent iuxta praeceptum regis et principum verbum Domini
2CHR|30|13|congregatique sunt in Hierusalem populi multi ut facerent sollemnitatem azymorum in mense secundo
2CHR|30|14|et surgentes destruxerunt altaria quae erant in Hierusalem atque universa in quibus idolis adolebatur incensum subvertentes proiecerunt in torrentem Cedron
2CHR|30|15|immolaverunt autem phase quartadecima die mensis secundi sacerdotes quoque atque Levitae tandem sanctificati obtulerunt holocausta in domo Domini
2CHR|30|16|steteruntque in ordine suo iuxta dispositionem et legem Mosi hominis Dei sacerdotes vero suscipiebant effundendum sanguinem de manibus Levitarum
2CHR|30|17|eo quod multa turba sanctificata non esset et idcirco Levitae immolarent phase his qui non occurrerant sanctificari Domino
2CHR|30|18|magna etiam pars populi de Ephraim et Manasse et Isachar et Zabulon quae sanctificata non fuerat comedit phase non iuxta quod scriptum est et oravit pro eis Ezechias dicens Dominus bonus propitiabitur
2CHR|30|19|cunctis qui in toto corde requirunt Dominum Deum patrum suorum et non inputabit eis quod minus sanctificati sunt
2CHR|30|20|quem exaudivit Dominus et placatus est populo
2CHR|30|21|feceruntque filii Israhel qui inventi sunt in Hierusalem sollemnitatem azymorum septem diebus in laetitia magna laudantes Dominum per singulos dies Levitae quoque et sacerdotes per organa quae suo officio congruebant
2CHR|30|22|et locutus est Ezechias ad cor omnium Levitarum qui habebant intellegentiam bonam super Domino et comederunt septem diebus sollemnitatis immolantes victimas pacificorum et laudantes Dominum Deum patrum suorum
2CHR|30|23|placuitque universae multitudini ut celebrarent etiam alios dies septem quod et fecerunt cum ingenti gaudio
2CHR|30|24|Ezechias enim rex Iuda praebuerat multitudini mille tauros et septem milia ovium principes vero dederant populo tauros mille et oves decem milia sanctificata ergo est sacerdotum plurima multitudo
2CHR|30|25|et hilaritate perfusa omnis turba Iuda tam sacerdotum et Levitarum quam universae frequentiae quae venerat ex Israhel proselytorum quoque de terra Israhel et habitantium in Iuda
2CHR|30|26|factaque est grandis celebritas in Hierusalem qualis a diebus Salomonis filii David regis Israhel in ea urbe non fuerat
2CHR|30|27|surrexerunt autem sacerdotes atque Levitae benedicentes populo et exaudita est vox eorum pervenitque oratio in habitaculum sanctum caeli
2CHR|31|1|cumque haec fuissent rite celebrata egressus est omnis Israhel qui inventus fuerat in urbibus Iuda et fregerunt simulacra succideruntque lucos demoliti sunt excelsa et altaria destruxerunt non solum de universo Iuda et Beniamin sed de Ephraim quoque et Manasse donec penitus everterent reversique sunt omnes filii Israhel in possessiones et civitates suas
2CHR|31|2|Ezechias vero constituit turmas sacerdotales et leviticas per divisiones suas unumquemque in officio proprio tam sacerdotum videlicet quam Levitarum ad holocausta et pacifica ut ministrarent et confiterentur canerentque in portis castrorum Domini
2CHR|31|3|pars autem regis erat ut de propria eius substantia offerretur holocaustum mane semper et vespere sabbatis quoque et kalendis et sollemnitatibus ceteris sicut scriptum est in lege Mosi
2CHR|31|4|praecepit etiam populo habitantium Hierusalem ut darent partes sacerdotibus et Levitis et possent vacare legi Domini
2CHR|31|5|quod cum percrebruisset in auribus multitudinis plurimas obtulere primitias filii Israhel frumenti vini et olei mellis quoque et omnium quae gignit humus decimas obtulerunt
2CHR|31|6|sed et filii Israhel et Iuda qui habitabant in urbibus Iuda obtulerunt decimas boum et ovium decimasque sanctorum quae voverant Domino Deo suo atque universa portantes fecerunt acervos plurimos
2CHR|31|7|mense tertio coeperunt acervorum iacere fundamenta et mense septimo conpleverunt eos
2CHR|31|8|cumque ingressi fuissent Ezechias et principes eius viderunt acervos et benedixerunt Domino ac populo Israhel
2CHR|31|9|interrogavitque Ezechias sacerdotes et Levitas cur ita iacerent acervi
2CHR|31|10|respondit illi Azarias sacerdos primus de stirpe Sadoc dicens ex quo coeperunt offerri primitiae in domo Domini comedimus et saturati sumus remanseruntque plurima eo quod benedixerit Dominus populo suo reliquiarum autem copia est ista quam cernis
2CHR|31|11|praecepit igitur Ezechias ut praepararent horrea in domo Domini quod cum fecissent
2CHR|31|12|intulerunt tam primitias quam decimas et quaecumque voverant fideliter fuit autem praefectus eorum Chonenias Levita et Semei frater eius secundus
2CHR|31|13|post quem Ieihel et Azazias et Naath et Asahel et Ierimoth Iozabath quoque et Helihel et Iesmachias et Maath et Banaias praepositi sub manibus Choneniae et Semei fratris eius ex imperio Ezechiae regis et Azariae pontificis domus Domini ad quos omnia pertinebant
2CHR|31|14|Core vero filius Iemna Levites et ianitor orientalis portae praepositus erat his quae sponte offerebantur Domino primitiisque et consecratis in sancta sanctorum
2CHR|31|15|et sub cura eius Eden et Meniamin Hiesue et Sameias Amarias quoque et Sechenias in civitatibus sacerdotum ut fideliter distribuerent fratribus suis partes minoribus atque maioribus
2CHR|31|16|exceptis maribus ab annis tribus et supra cunctis qui ingrediebantur templum Domini et quicquid per dies singulos conducebat in ministerio atque observationibus iuxta divisiones suas
2CHR|31|17|sacerdotibus per familias et Levitis a vicesimo anno et supra per ordines et turmas suas
2CHR|31|18|universaeque multitudini tam uxoribus quam liberis eorum utriusque sexus fideliter cibi de his quae sanctificata fuerant praebebantur
2CHR|31|19|sed et filiorum Aaron per agros et suburbana urbium singularum dispositi erant viri qui partes distribuerent universo sexui masculino de sacerdotibus et Levitis
2CHR|31|20|fecit ergo Ezechias universa quae diximus in omni Iuda operatusque est bonum et rectum et verum coram Domino Deo suo
2CHR|31|21|in universa cultura ministerii domus Domini iuxta legem et caerimonias volens requirere Deum suum in toto corde suo fecitque et prosperatus est
2CHR|32|1|post quae et huiuscemodi veritatem venit Sennacherib rex Assyriorum et ingressus Iudam obsedit civitates munitas volens eas capere
2CHR|32|2|quod cum vidisset Ezechias venisse scilicet Sennacherib et totum belli impetum verti contra Hierusalem
2CHR|32|3|inito cum principibus consilio virisque fortissimis ut obturarent capita fontium quae erant extra urbem et hoc omnium decernente sententia
2CHR|32|4|congregavit plurimam multitudinem et obturaverunt cunctos fontes et rivum qui fluebat in medio terrae dicentes ne veniant reges Assyriorum et inveniant aquarum abundantiam
2CHR|32|5|aedificavit quoque agens industrie omnem murum qui fuerat dissipatus et extruxit turres desuper et forinsecus alterum murum instauravitque Mello in civitate David et fecit universi generis armaturam et clypeos
2CHR|32|6|constituitque principes bellatorum in exercitu et convocavit universos in platea portae civitatis ac locutus est ad cor eorum dicens
2CHR|32|7|viriliter agite et confortamini nolite timere nec paveatis regem Assyriorum et universam multitudinem quae est cum eo multo enim plures nobiscum sunt quam cum illo
2CHR|32|8|cum illo est brachium carneum nobiscum Dominus Deus noster qui auxiliator est noster pugnatque pro nobis confortatusque est populus huiuscemodi verbis Ezechiae regis Iuda
2CHR|32|9|quae postquam gesta sunt misit Sennacherib rex Assyriorum servos suos Hierusalem ipse enim cum universo exercitu obsidebat Lachis ad Ezechiam regem Iuda et ad omnem populum qui erat in urbe dicens
2CHR|32|10|haec dicit Sennacherib rex Assyriorum in quo habentes fiduciam sedetis obsessi in Hierusalem
2CHR|32|11|num Ezechias decipit vos ut tradat morti in fame et siti adfirmans quod Dominus Deus vester liberet vos de manu regis Assyriorum
2CHR|32|12|numquid non iste est Ezechias qui destruxit excelsa illius et altaria et praecepit Iudae et Hierusalem dicens coram altari uno adorabitis et in ipso conburetis incensum
2CHR|32|13|an ignoratis quae ego fecerim et patres mei cunctis terrarum populis numquid praevaluerunt dii gentium omniumque terrarum liberare regionem suam de manu mea
2CHR|32|14|quis est de universis diis gentium quas vastaverunt patres mei qui potuerit eruere populum suum de manu mea ut possit etiam Deus vester eruere vos de hac manu
2CHR|32|15|non vos ergo decipiat Ezechias nec vana persuasione deludat neque credatis ei si enim nullus potuit deus cunctarum gentium atque regnorum liberare populum suum de manu mea et de manu patrum meorum consequenter nec Deus vester poterit eruere vos de hac manu
2CHR|32|16|sed et alia multa locuti sunt servi eius contra Dominum Deum et contra Ezechiam servum eius
2CHR|32|17|epistulas quoque scripsit plenas blasphemiae in Dominum Deum Israhel et locutus est adversus eum sicut dii gentium ceterarum non potuerunt liberare populos suos de manu mea sic et Deus Ezechiae eruere non poterit populum suum de manu ista
2CHR|32|18|insuper et clamore magno lingua iudaica contra populum qui sedebat in muris Hierusalem personabat ut terreret eos et caperet civitatem
2CHR|32|19|locutusque est contra Deum Hierusalem sicut adversum deos populorum terrae opera manuum hominum
2CHR|32|20|oraverunt igitur Ezechias rex et Esaias filius Amos prophetes adversum hanc blasphemiam ac vociferati sunt usque in caelum
2CHR|32|21|et misit Dominus angelum qui percussit omnem virum robustum et bellatorem et principem exercitus regis Assyriorum reversusque est cum ignominia in terram suam cumque ingressus esset domum dei sui filii qui egressi fuerant de utero eius interfecerunt eum gladio
2CHR|32|22|salvavitque Dominus Ezechiam et habitatores Hierusalem de manu Sennacherib regis Assyriorum et de manu omnium et praestitit ei quietem per circuitum
2CHR|32|23|multi etiam deferebant hostias et sacrificia Domino Hierusalem et munera Ezechiae regi Iuda qui exaltatus est post haec coram cunctis gentibus
2CHR|32|24|in diebus illis aegrotavit Ezechias usque ad mortem et oravit Dominum exaudivitque eum et dedit ei signum
2CHR|32|25|sed non iuxta beneficia quae acceperat retribuit quia elevatum est cor eius et facta est contra eum ira et contra Iudam ac Hierusalem
2CHR|32|26|humiliatusque est postea eo quod exaltatum fuisset cor eius tam ipse quam habitatores Hierusalem et idcirco non venit super eos ira Domini in diebus Ezechiae
2CHR|32|27|fuit autem Ezechias dives et inclitus valde et thesauros sibi plurimos congregavit argenti auri et lapidis pretiosi aromatum et armorum universi generis et vasorum magni pretii
2CHR|32|28|apothecas quoque frumenti vini et olei et praesepia omnium iumentorum caulasque pecoribus
2CHR|32|29|et urbes exaedificavit habebat quippe greges ovium et armentorum innumerabiles eo quod dedisset ei Dominus substantiam multam nimis
2CHR|32|30|ipse est Ezechias qui obturavit superiorem fontem aquarum Gion et avertit eas subter ad occidentem urbis David in omnibus operibus suis fecit prospere quae voluit
2CHR|32|31|attamen in legatione principum Babylonis qui missi fuerant ad eum ut interrogarent de portento quod acciderat super terram dereliquit eum Deus ut temptaretur et nota fierent omnia quae erant in corde eius
2CHR|32|32|reliqua autem sermonum Ezechiae et misericordiarum eius scripta sunt in visione Esaiae filii Amos prophetae et in libro regum Iuda et Israhel
2CHR|32|33|dormivitque Ezechias cum patribus suis et sepelierunt eum supra sepulchra filiorum David et celebravit eius exequias universus Iuda et omnes habitatores Hierusalem regnavitque Manasses filius eius pro eo
2CHR|33|1|duodecim annorum erat Manasses cum regnare coepisset et quinquaginta quinque annis regnavit in Hierusalem
2CHR|33|2|fecit autem malum coram Domino iuxta abominationes gentium quas subvertit Dominus coram filiis Israhel
2CHR|33|3|et conversus instauravit excelsa quae demolitus fuerat Ezechias pater eius construxitque aras Baalim et fecit lucos et adoravit omnem militiam caeli et coluit eam
2CHR|33|4|aedificavit quoque altaria in domo Domini de qua dixerat Dominus in Hierusalem erit nomen meum in aeternum
2CHR|33|5|aedificavit autem ea cuncto exercitui caeli in duobus atriis domus Domini
2CHR|33|6|transireque fecit filios suos per ignem in valle Benennon observabat somnia sectabatur auguria maleficis artibus inserviebat habebat secum magos et incantatores multaque mala operatus est coram Domino ut inritaret eum
2CHR|33|7|sculptile quoque et conflatile signum posuit in domo Domini de qua locutus est Dominus ad David et ad Salomonem filium eius dicens in domo hac et in Hierusalem quam elegi de cunctis tribubus Israhel ponam nomen meum in sempiternum
2CHR|33|8|et movere non faciam pedem Israhel de terra quam tradidi patribus eorum ita dumtaxat si custodierint facere quae praecepi eis cunctamque legem et caerimonias atque iudicia per manum Mosi
2CHR|33|9|igitur Manasses seduxit Iudam et habitatores Hierusalem ut facerent malum super omnes gentes quas subverterat Dominus a facie filiorum Israhel
2CHR|33|10|locutusque est Dominus ad eum et ad populum illius et adtendere noluerunt
2CHR|33|11|idcirco superinduxit eis principes exercitus regis Assyriorum ceperuntque Manassen et vinctum catenis atque conpedibus duxerunt Babylonem
2CHR|33|12|qui postquam coangustatus est oravit Dominum Deum suum et egit paenitentiam valde coram Deo patrum suorum
2CHR|33|13|deprecatusque est eum et obsecravit intente et exaudivit orationem eius reduxitque eum Hierusalem in regnum suum et cognovit Manasses quod Dominus ipse esset Deus
2CHR|33|14|post haec aedificavit murum extra civitatem David ad occidentem Gion in convalle ab introitu portae Piscium per circuitum usque ad Ophel et exaltavit illum vehementer constituitque principes exercitus in cunctis civitatibus Iuda munitis
2CHR|33|15|et abstulit deos alienos et simulacrum de domo Domini aras quoque quas fecerat in monte domus Domini et in Hierusalem et proiecit omnia extra urbem
2CHR|33|16|porro instauravit altare Domini et immolavit super illud victimas et pacifica et laudem praecepitque Iudae ut serviret Domino Deo Israhel
2CHR|33|17|attamen adhuc populus immolabat in excelsis Domino Deo suo
2CHR|33|18|reliqua autem gestorum Manasse et obsecratio eius ad Deum suum verba quoque videntium qui loquebantur ad eum in nomine Domini Dei Israhel continentur in sermonibus regum Israhel
2CHR|33|19|oratio quoque eius et exauditio et cuncta peccata atque contemptus loca etiam in quibus aedificavit excelsa et fecit lucos et statuas antequam ageret paenitentiam scripta sunt in sermonibus Ozai
2CHR|33|20|dormivit ergo Manasses cum patribus suis et sepelierunt eum in domo sua regnavitque pro eo filius eius Amon
2CHR|33|21|viginti duo annorum erat Amon cum regnare coepisset et duobus annis regnavit in Hierusalem
2CHR|33|22|fecitque malum in conspectu Domini sicut fecerat Manasses pater eius et cunctis idolis quae Manasses fuerat fabricatus immolavit atque servivit
2CHR|33|23|et non est reveritus faciem Domini sicut reveritus est Manasses pater eius et multo maiora deliquit
2CHR|33|24|cumque coniurassent adversus eum servi sui interfecerunt eum in domo sua
2CHR|33|25|porro reliqua populi multitudo caesis his qui Amon percusserant constituit regem Iosiam filium eius pro eo
2CHR|34|1|octo annorum erat Iosias cum regnare coepisset et triginta et uno annis regnavit in Hierusalem
2CHR|34|2|fecitque quod erat rectum in conspectu Domini et ambulavit in viis David patris sui non declinavit neque ad dexteram neque ad sinistram
2CHR|34|3|octavo autem anno regni sui cum adhuc esset puer coepit quaerere Deum patris sui David et duodecimo anno postquam coeperat mundavit Iudam et Hierusalem ab excelsis et lucis simulacrisque et sculptilibus
2CHR|34|4|destruxeruntque coram eo aras Baalim et simulacra quae superposita fuerant demoliti sunt lucos etiam et sculptilia succidit atque comminuit et super tumulos eorum qui eis immolare consueverant fragmenta dispersit
2CHR|34|5|ossa praeterea sacerdotum conbusit in altaribus idolorum mundavitque Iudam et Hierusalem
2CHR|34|6|sed et in urbibus Manasse et Ephraim et Symeon usque Nepthalim cuncta subvertit
2CHR|34|7|cumque altaria dissipasset et lucos et sculptilia contrivisset in frusta cunctaque delubra demolitus esset de universa terra Israhel reversus est Hierusalem
2CHR|34|8|igitur anno octavodecimo regni sui mundata iam terra et templo Domini misit Saphan filium Eseliae et Maasiam principem civitatis et Ioha filium Ioachaz a commentariis ut instaurarent domum Domini Dei sui
2CHR|34|9|qui venerunt ad Helciam sacerdotem magnum acceptamque ab eo pecuniam quae inlata fuerat in domum Domini et quam congregaverant Levitae ianitores de Manasse et Ephraim et universis reliquiis Israhel ab omni quoque Iuda et Beniamin et habitatoribus Hierusalem
2CHR|34|10|tradiderunt in manibus eorum qui praeerant operariis in domo Domini ut instaurarent templum et infirma quaeque sarcirent
2CHR|34|11|at illi dederunt eam artificibus et cementariis ut emerent lapides de lapidicinis et ligna ad commissuras aedificii et ad contignationem domorum quas destruxerant reges Iuda
2CHR|34|12|qui fideliter cuncta faciebant erant autem praepositi operantium Iaath et Abdias de filiis Merari Zaccharias et Mosollam de filiis Caath qui urguebant opus omnes Levitae scientes organis canere
2CHR|34|13|super eos vero qui ad varios usus onera portabant erant scribae et magistri de Levitis ianitores
2CHR|34|14|cumque efferrent pecuniam quae inlata fuerat in templum Domini repperit Helcias sacerdos librum legis Domini per manum Mosi
2CHR|34|15|et ait ad Saphan scribam librum legis inveni in domo Domini et tradidit ei
2CHR|34|16|at ille intulit volumen ad regem et nuntiavit ei dicens omnia quae dedisti in manu servorum tuorum ecce conplentur
2CHR|34|17|argentum quod reppertum est in domo Domini conflaverunt datumque est praefectis artificum et diversa opera fabricantium
2CHR|34|18|praeterea tradidit mihi Helcias sacerdos hunc librum quem cum rege praesente recitasset
2CHR|34|19|audissetque ille verba legis scidit vestimenta sua
2CHR|34|20|et praecepit Helciae et Ahicam filio Saphan et Abdon filio Micha Saphan quoque scribae et Asaiae servo regis dicens
2CHR|34|21|ite et orate Dominum pro me et pro reliquiis Israhel et Iuda super universis sermonibus libri istius qui reppertus est magnus enim furor Domini stillavit super nos eo quod non custodierint patres nostri verba Domini ut facerent omnia quae scripta sunt in isto volumine
2CHR|34|22|abiit igitur Helcias et hii qui simul a rege missi fuerant ad Holdan propheten uxorem Sellum filii Thecuath filii Hasra custodis vestium quae habitabat Hierusalem in secunda et locuti sunt ei verba quae supra narravimus
2CHR|34|23|at illa respondit eis haec dicit Dominus Deus Israhel dicite viro qui misit vos ad me
2CHR|34|24|haec dicit Dominus ecce ego inducam mala super locum istum et super habitatores eius cunctaque maledicta quae scripta sunt in libro hoc quem legerunt coram rege Iuda
2CHR|34|25|quia dereliquerunt me et sacrificaverunt diis alienis ut me ad iracundiam provocarent in cunctis operibus manuum suarum idcirco stillavit furor meus super locum istum et non extinguetur
2CHR|34|26|ad regem autem Iuda qui misit vos pro Domino deprecando sic loquimini haec dicit Dominus Deus Israhel quoniam audisti verba voluminis
2CHR|34|27|atque emollitum est cor tuum et humiliatus es in conspectu Dei super his quae dicta sunt contra locum hunc et habitatores Hierusalem reveritusque faciem meam scidisti vestimenta tua et flevisti coram me ego quoque exaudivi te dicit Dominus
2CHR|34|28|iam enim colligam te ad patres tuos et infereris in sepulchrum tuum in pace nec videbunt oculi tui omne malum quod ego inducturus sum super locum istum et super habitatores eius rettulerunt itaque regi cuncta quae dixerat
2CHR|34|29|at ille convocatis universis maioribus natu Iuda et Hierusalem
2CHR|34|30|ascendit domum Domini unaque omnes viri Iuda et habitatores Hierusalem sacerdotes et Levitae et cunctus populus a minimo usque ad maximum quibus audientibus in domo Domini legit rex omnia verba voluminis
2CHR|34|31|et stans in tribunali suo percussit foedus coram Domino ut ambularet post eum et custodiret praecepta et testimonia et iustificationes eius in toto corde suo et in tota anima sua faceretque quae scripta sunt in volumine illo quem legerat
2CHR|34|32|adiuravit quoque super hoc omnes qui repperti fuerant in Hierusalem et Beniamin et fecerunt habitatores Hierusalem iuxta pactum Domini Dei patrum suorum
2CHR|34|33|abstulit ergo Iosias cunctas abominationes de universis regionibus filiorum Israhel et fecit omnes qui residui erant in Israhel servire Domino Deo suo cunctis diebus eius non recesserunt a Domino Deo patrum suorum
2CHR|35|1|fecit autem Iosias in Hierusalem phase Domino quod immolatum est quartadecima die mensis primi
2CHR|35|2|et constituit sacerdotes in officiis suis hortatusque est eos ut ministrarent in domo Domini
2CHR|35|3|Levitis quoque ad quorum eruditionem omnis Israhel sanctificabatur Domino locutus est ponite arcam in sanctuario templi quod aedificavit Salomon filius David rex Israhel nequaquam enim eam ultra portabitis nunc autem ministrate Domino Deo vestro et populo eius Israhel
2CHR|35|4|et praeparate vos per domos et cognationes vestras in divisionibus singulorum sicut praecepit David rex Israhel et descripsit Salomon filius eius
2CHR|35|5|ministrate in sanctuario per familias turmasque leviticas
2CHR|35|6|et sanctificati immolate phase fratres etiam vestros ut possint iuxta verba quae locutus est Dominus in manu Mosi facere praeparate
2CHR|35|7|dedit praeterea Iosias omni populo qui ibi fuerat inventus in sollemnitatem phase agnos et hedos de gregibus et reliqui pecoris triginta milia boumque tria milia haec de regis universa substantia
2CHR|35|8|duces quoque eius sponte quod voluerant obtulerunt tam populo quam sacerdotibus et Levitis porro Helcias et Zaccharias et Iehihel principes domus Domini dederunt sacerdotibus ad faciendum phase pecora commixtim duo milia sescenta et boves trecentos
2CHR|35|9|Chonenias autem Semeias etiam et Nathanahel fratres eius necnon Asabias et Iahihel et Iozabath principes Levitarum dederunt ceteris Levitis ad celebrandum phase quinque milia pecorum et boves quingentos
2CHR|35|10|praeparatumque est ministerium et steterunt sacerdotes in officio suo Levitae quoque in turmis iuxta regis imperium
2CHR|35|11|et immolatum est phase asperseruntque sacerdotes manu sua sanguinem et Levitae detraxerunt pelles holocaustorum
2CHR|35|12|et separaverunt ea ut darent per domos et familias singulorum et offerrentur Domino sicut scriptum est in libro Mosi de bubus quoque fecere similiter
2CHR|35|13|et assaverunt phase super ignem iuxta quod lege praeceptum est pacificas vero hostias coxerunt in lebetis et caccabis et ollis et festinato distribuerunt universae plebi
2CHR|35|14|sibi autem et sacerdotibus postea paraverunt nam in oblatione holocaustorum et adipum usque ad noctem sacerdotes fuerant occupati unde Levitae et sibi et sacerdotibus filiis Aaron paraverunt novissimis
2CHR|35|15|porro cantores filii Asaph stabant in ordine suo iuxta praeceptum David et Asaph et Heman et Idithun prophetarum regis ianitores vero per portas singulas observabant ita ut ne puncto quidem discederent a ministerio quam ob rem et fratres eorum Levitae paraverunt eis cibos
2CHR|35|16|omnis igitur cultura Domini rite conpleta est in die illa ut facerent phase et offerrent holocausta super altare Domini iuxta praeceptum regis Iosiae
2CHR|35|17|feceruntque filii Israhel qui repperti fuerant ibi phase in tempore illo et sollemnitatem azymorum septem diebus
2CHR|35|18|non fuit phase simile huic in Israhel a diebus Samuhelis prophetae sed nec quisquam de cunctis regibus Israhel fecit phase sicut Iosias sacerdotibus et Levitis et omni Iuda et Israhel qui reppertus fuerat et habitantibus in Hierusalem
2CHR|35|19|octavodecimo anno regni Iosiae hoc phase celebratum est
2CHR|35|20|postquam instauraverat Iosias templum ascendit Nechao rex Aegypti ad pugnandum in Charchamis iuxta Eufraten et processit in occursum eius Iosias
2CHR|35|21|at ille missis ad eum nuntiis ait quid mihi et tibi est rex Iuda non adversum te hodie venio sed contra aliam pugno domum ad quam me Deus festinato ire praecepit desine adversum Deum facere qui mecum est ne interficiat te
2CHR|35|22|noluit Iosias reverti sed praeparavit contra eum bellum nec adquievit sermonibus Nechao ex ore Dei verum perrexit ut dimicaret in campo Mageddo
2CHR|35|23|ibique vulneratus a sagittariis dixit pueris suis educite me de proelio quia oppido vulneratus sum
2CHR|35|24|qui transtulerunt eum de curru in alterum currum qui sequebatur eum more regio et asportaverunt in Hierusalem mortuusque est et sepultus in mausoleo patrum suorum et universus Iuda et Hierusalem luxerunt eum
2CHR|35|25|Hieremias maxime cuius omnes cantores atque cantrices usque in praesentem diem lamentationes super Iosia replicant et quasi lex obtinuit in Israhel ecce scriptum fertur in Lamentationibus
2CHR|35|26|reliqua autem sermonum Iosiae et misericordiarum eius quae lege praecepta sunt Domini
2CHR|35|27|opera quoque illius prima et novissima scripta sunt in libro regum Israhel et Iuda
2CHR|36|1|tulit ergo populus terrae Ioachaz filium Iosiae et constituit regem pro patre suo in Hierusalem
2CHR|36|2|viginti trium annorum erat Ioachaz cum regnare coepisset et tribus mensibus regnavit in Hierusalem
2CHR|36|3|amovit autem eum rex Aegypti cum venisset Hierusalem et condemnavit terram centum talentis argenti et talento auri
2CHR|36|4|constituitque regem pro eo Eliacim fratrem eius super Iudam et Hierusalem et vertit nomen eius Ioacim ipsum vero Ioachaz tulit secum et adduxit in Aegyptum
2CHR|36|5|viginti quinque annorum erat Ioacim cum regnare coepisset et undecim annis regnavit in Hierusalem fecitque malum coram Domino Deo suo
2CHR|36|6|contra hunc ascendit Nabuchodonosor rex Chaldeorum et vinctum catenis duxit in Babylonem
2CHR|36|7|ad quam et vasa Domini transtulit et posuit ea in templo suo
2CHR|36|8|reliqua autem verborum Ioacim et abominationum eius quas operatus est et quae inventa sunt in eo continentur in libro regum Israhel et Iuda regnavitque Ioachin filius eius pro eo
2CHR|36|9|octo annorum erat Ioachin cum regnare coepisset et tribus mensibus ac decem diebus regnavit in Hierusalem fecitque malum in conspectu Domini
2CHR|36|10|cumque anni circulus volveretur misit Nabuchodonosor rex qui et adduxerunt eum in Babylonem asportatis simul pretiosissimis vasis domus Domini regem vero constituit Sedeciam fratrem eius super Iudam et Hierusalem
2CHR|36|11|viginti et unius anni erat Sedecias cum regnare coepisset et undecim annis regnavit in Hierusalem
2CHR|36|12|fecitque malum in oculis Domini Dei sui nec erubuit faciem Hieremiae prophetae loquentis ad se ex ore Domini
2CHR|36|13|a rege quoque Nabuchodonosor recessit qui adiuraverat eum per Deum et induravit cervicem suam et cor ut non reverteretur ad Dominum Deum Israhel
2CHR|36|14|sed et universi principes sacerdotum et populus praevaricati sunt inique iuxta universas abominationes gentium et polluerunt domum Domini quam sanctificaverat sibi in Hierusalem
2CHR|36|15|mittebat autem Dominus Deus patrum suorum ad illos per manum nuntiorum suorum de nocte consurgens et cotidie commonens eo quod parceret populo et habitaculo suo
2CHR|36|16|at illi subsannabant nuntios Dei et parvipendebant sermones eius inludebantque prophetis donec ascenderet furor Domini in populum eius et esset nulla curatio
2CHR|36|17|adduxit enim super eos regem Chaldeorum et interfecit iuvenes eorum gladio in domo sanctuarii sui non est misertus adulescentis et virginis et senis nec decrepiti quidem sed omnes tradidit manibus eius
2CHR|36|18|universaque vasa domus Domini tam maiora quam minora et thesauros templi et regis et principum transtulit in Babylonem
2CHR|36|19|incenderunt hostes domum Dei destruxerunt murum Hierusalem universas turres conbuserunt et quicquid pretiosum fuerat demoliti sunt
2CHR|36|20|si quis evaserat gladium ductus in Babylonem servivit regi et filiis eius donec imperaret rex Persarum
2CHR|36|21|et conpleretur sermo Domini ex ore Hieremiae et celebraret terra sabbata sua cunctis enim diebus desolationis egit sabbatum usque dum conplerentur septuaginta anni
2CHR|36|22|anno autem primo Cyri regis Persarum ad explendum sermonem Domini quem locutus fuerat per os Hieremiae suscitavit Dominus spiritum Cyri regis Persarum qui iussit praedicari in universo regno suo etiam per scripturam dicens
2CHR|36|23|haec dicit Cyrus rex Persarum omnia regna terrae dedit mihi Dominus Deus caeli et ipse praecepit mihi ut aedificarem ei domum in Hierusalem quae est in Iudaea quis ex vobis est in omni populo eius sit Dominus Deus suus cum eo et ascendat
EZRA|1|1|in anno primo Cyri regis Persarum ut conpleretur verbum Domini ex ore Hieremiae suscitavit Dominus spiritum Cyri regis Persarum et transduxit vocem in universo regno suo etiam per scripturam dicens
EZRA|1|2|haec dicit Cyrus rex Persarum omnia regna terrae dedit mihi Dominus Deus caeli et ipse praecepit mihi ut aedificarem ei domum in Hierusalem quae est in Iudaea
EZRA|1|3|quis est in vobis de universo populo eius sit Deus illius cum ipso ascendat Hierusalem quae est in Iudaea et aedificet domum Domini Dei Israhel ipse est Deus qui est in Hierusalem
EZRA|1|4|et omnes reliqui in cunctis locis ubicumque habitant adiuvent eum viri de loco suo argento et auro et substantia et pecoribus excepto quod voluntarie offerunt templo Dei quod est in Hierusalem
EZRA|1|5|et surrexerunt principes patrum de Iuda et Beniamin et sacerdotes et Levitae omnis cuius suscitavit Deus spiritum ut ascenderent ad aedificandum templum Domini quod erat in Hierusalem
EZRA|1|6|universique qui erant in circuitu adiuverunt manus eorum in vasis argenteis et aureis in substantia in iumentis in supellectili exceptis his quae sponte obtulerunt
EZRA|1|7|rex quoque Cyrus protulit vasa templi Domini quae tulerat Nabuchodonosor de Hierusalem et posuerat ea in templo dei sui
EZRA|1|8|protulit autem ea Cyrus rex Persarum per manum Mitridatis filii Gazabar et adnumeravit ea Sasabassar principi Iudae
EZRA|1|9|et hic est numerus eorum fialae aureae triginta fialae argenteae mille cultri viginti novem scyphi aurei triginta
EZRA|1|10|scyphi argentei secundi quadringenti decem vasa alia mille
EZRA|1|11|omnia vasa aurea et argentea quinque milia quadringenta universa tulit Sasabassar cum his qui ascendebant de transmigratione Babylonis in Hierusalem
EZRA|2|1|hii sunt autem filii provinciae qui ascenderunt de captivitate quam transtulerat Nabuchodonosor rex Babylonis in Babylonem et reversi sunt in Hierusalem et Iudam unusquisque in civitatem suam
EZRA|2|2|qui venerunt cum Zorobabel Hiesua Neemia Saraia Rahelaia Mardochai Belsan Mesphar Beguai Reum Baana numerus virorum populi Israhel
EZRA|2|3|filii Pharos duo milia centum septuaginta duo
EZRA|2|4|filii Sephetia trecenti septuaginta duo
EZRA|2|5|filii Area septingenti septuaginta quinque
EZRA|2|6|filii Phaethmoab filiorum Iosue Ioab duo milia octingenti duodecim
EZRA|2|7|filii Helam mille ducenti quinquaginta quattuor
EZRA|2|8|filii Zeththua nongenti quadraginta quinque
EZRA|2|9|filii Zacchai septingenti sexaginta
EZRA|2|10|filii Bani sescenti quadraginta duo
EZRA|2|11|filii Bebai sescenti viginti tres
EZRA|2|12|filii Azgad mille ducenti viginti duo
EZRA|2|13|filii Adonicam sescenti sexaginta sex
EZRA|2|14|filii Beguai duo milia quinquaginta sex
EZRA|2|15|filii Adin quadringenti quinquaginta quattuor
EZRA|2|16|filii Ater qui erant ex Hiezechia nonaginta octo
EZRA|2|17|filii Besai trecenti viginti tres
EZRA|2|18|filii Iora centum duodecim
EZRA|2|19|filii Asom ducenti viginti tres
EZRA|2|20|filii Gebbar nonaginta quinque
EZRA|2|21|filii Bethleem centum viginti tres
EZRA|2|22|viri Netupha quinquaginta sex
EZRA|2|23|viri Anathoth centum viginti octo
EZRA|2|24|filii Azmaveth quadraginta duo
EZRA|2|25|filii Cariathiarim Caephira et Beroth septingenti quadraginta tres
EZRA|2|26|filii Arama et Gaba sescenti viginti unus
EZRA|2|27|viri Machmas centum viginti duo
EZRA|2|28|viri Bethel et Gai ducenti viginti tres
EZRA|2|29|filii Nebo quinquaginta duo
EZRA|2|30|filii Megbis centum quinquaginta sex
EZRA|2|31|filii Helam alterius mille ducenti quinquaginta quattuor
EZRA|2|32|filii Arim trecenti viginti
EZRA|2|33|filii Lod Adid et Ono septingenti viginti quinque
EZRA|2|34|filii Hiericho trecenti quadraginta quinque
EZRA|2|35|filii Sennaa tria milia sescenti triginta
EZRA|2|36|sacerdotes filii Idaia in domo Hiesue nongenti septuaginta tres
EZRA|2|37|filii Emmer mille quinquaginta duo
EZRA|2|38|filii Phessur mille ducenti quadraginta septem
EZRA|2|39|filii Arim mille decem et septem
EZRA|2|40|Levitae filii Hiesue et Cedmihel filiorum Odevia septuaginta quattuor
EZRA|2|41|cantores filii Asaph centum viginti octo
EZRA|2|42|filii ianitorum filii Sellum filii Ater filii Telmon filii Accub filii Atita filii Sobai universi centum triginta novem
EZRA|2|43|Nathinnei filii Sia filii Asupha filii Tebbaoth
EZRA|2|44|filii Ceros filii Siaa filii Phadon
EZRA|2|45|filii Levana filii Agaba filii Accub
EZRA|2|46|filii Agab filii Selmai filii Anan
EZRA|2|47|filii Gaddel filii Gaer filii Rahaia
EZRA|2|48|filii Rasin filii Nechoda filii Gazem
EZRA|2|49|filii Aza filii Phasea filii Besee
EZRA|2|50|filii Asenaa filii Munim filii Nephusim
EZRA|2|51|filii Becbuc filii Acupha filii Arur
EZRA|2|52|filii Besluth filii Maida filii Arsa
EZRA|2|53|filii Bercos filii Sisara filii Thema
EZRA|2|54|filii Nasia filii Atupha
EZRA|2|55|filii servorum Salomonis filii Sotei filii Suphereth filii Pharuda
EZRA|2|56|filii Iala filii Dercon filii Gedel
EZRA|2|57|filii Saphatia filii Athil filii Phocereth qui erant de Asebaim filii Ammi
EZRA|2|58|omnes Nathinnei et filii servorum Salomonis trecenti nonaginta duo
EZRA|2|59|et hii qui ascenderunt de Thelmela Thelarsa Cherub et Don et Mer et non potuerunt indicare domum patrum suorum et semen suum utrum ex Israhel essent
EZRA|2|60|filii Delaia filii Tobia filii Necoda sescenti quinquaginta duo
EZRA|2|61|et de filiis sacerdotum filii Obia filii Accos filii Berzellai qui accepit de filiabus Berzellai Galaditis uxorem et vocatus est nomine eorum
EZRA|2|62|hii quaesierunt scripturam genealogiae suae et non invenerunt et eiecti sunt de sacerdotio
EZRA|2|63|et dixit Athersatha eis ut non comederent de sancto sanctorum donec surgeret sacerdos doctus atque perfectus
EZRA|2|64|omnis multitudo quasi unus quadraginta duo milia trecenti sexaginta
EZRA|2|65|exceptis servis eorum et ancillis qui erant septem milia trecenti triginta septem et in ipsis cantores atque cantrices ducentae
EZRA|2|66|equi eorum septingenti triginta sex muli eorum ducenti quadraginta quinque
EZRA|2|67|cameli eorum quadringenti triginta quinque asini eorum sex milia septingenti viginti
EZRA|2|68|et de principibus patrum cum ingrederentur templum Domini quod est in Hierusalem sponte obtulerunt in domum Dei ad extruendam eam in loco suo
EZRA|2|69|secundum vires suas dederunt in inpensas operis auri solidos sexaginta milia et mille argenti minas quinque milia et vestes sacerdotales centum
EZRA|2|70|habitaverunt ergo sacerdotes et Levitae et de populo et cantores et ianitores et Nathinnei in urbibus suis universusque Israhel in civitatibus suis
EZRA|3|1|iamque venerat mensis septimus et erant filii Israhel in civitatibus suis congregatus est ergo populus quasi vir unus in Hierusalem
EZRA|3|2|et surrexit Iosue filius Iosedech et fratres eius sacerdotes et Zorobabel filius Salathihel et fratres eius et aedificaverunt altare Dei Israhel ut offerrent in eo holocaustomata sicut scriptum est in lege Mosi viri Dei
EZRA|3|3|conlocaverunt autem altare super bases suas deterrentibus eos per circuitum populis terrarum et obtulerunt super illud holocaustum Domino mane et vespere
EZRA|3|4|feceruntque sollemnitatem tabernaculorum sicut scriptum est et holocaustum diebus singulis per ordinem secundum praeceptum opus diei in die suo
EZRA|3|5|et post haec holocaustum iuge tam in kalendis quam in universis sollemnitatibus Domini quae erant consecratae et in omnibus in quibus ultro offerebatur munus Deo
EZRA|3|6|a primo die mensis septimi coeperunt offerre holocaustum Domino porro templum Dei fundatum necdum erat
EZRA|3|7|dederunt autem pecunias latomis et cementariis cibum quoque et potum et oleum Sidoniis Tyriisque ut deferrent ligna cedrina de Libano ad mare Ioppes iuxta quod praeceperat Cyrus rex Persarum eis
EZRA|3|8|anno autem secundo adventus eorum ad templum Dei in Hierusalem mense secundo coeperunt Zorobabel filius Salathihel et Iosue filius Iosedech et reliqui de fratribus eorum sacerdotes et Levitae et omnes qui venerant de captivitate in Hierusalem et constituerunt Levitas a viginti annis et supra ut urguerent opus Domini
EZRA|3|9|stetitque Iosue filii eius et fratres eius Cedmihel et filii eius et filii Iuda quasi unus ut instarent super eos qui faciebant opus in templo Dei filii Enadad filii eorum et fratres eorum Levitae
EZRA|3|10|fundato igitur a cementariis templo Domini steterunt sacerdotes in ornatu suo cum tubis et Levitae filii Asaph in cymbalis ut laudarent Deum per manus David regis Israhel
EZRA|3|11|et concinebant in hymnis et confessione Domino quoniam bonus quoniam in aeternum misericordia eius super Israhel omnis quoque populus vociferabatur clamore magno in laudando Dominum eo quod fundatum esset templum Domini
EZRA|3|12|plurimi etiam de sacerdotibus et Levitis et principes patrum seniores qui viderant templum prius cum fundatum esset et hoc templum in oculis eorum flebant voce magna et multi vociferantes in laetitia elevabant vocem
EZRA|3|13|nec poterat quisquam agnoscere vocem clamoris laetantium et vocem fletus populi commixtim enim populus vociferabatur clamore magno et vox audiebatur procul
EZRA|4|1|audierunt autem hostes Iudae et Beniamin quia filii captivitatis aedificarent templum Domino Deo Israhel
EZRA|4|2|et accedentes ad Zorobabel et ad principes patrum dixerunt eis aedificemus vobiscum quia ita ut vos quaerimus Deum vestrum ecce nos immolamus victimas ex diebus Asoraddan regis Assur qui adduxit nos huc
EZRA|4|3|et dixit eis Zorobabel et Iosue et reliqui principes patrum Israhel non est vobis et nobis ut aedificemus domum Deo nostro sed nos ipsi soli aedificabimus Domino Deo nostro sicut praecepit nobis rex Cyrus rex Persarum
EZRA|4|4|factum est igitur ut populus terrae inpediret manus populi Iudae et turbaret eos in aedificando
EZRA|4|5|conduxerunt quoque adversum eos consiliatores ut destruerent consilium eorum omnibus diebus Cyri regis Persarum et usque ad regnum Darii regis Persarum
EZRA|4|6|in regno autem Asueri principio regni eius scripserunt accusationem adversum habitatores Iudae et Hierusalem
EZRA|4|7|et in diebus Artarxersis scripsit Beselam Mitridatis et Tabel et reliqui qui erant in consilio eorum ad Artarxersen regem Persarum epistula autem accusationis scripta erat syriace et legebatur sermone syro
EZRA|4|8|Reum Beelteem et Samsai scriba scripserunt epistulam unam de Hierusalem Artarxersi regi huiuscemodi
EZRA|4|9|Reum Beelteem et Samsai scriba et reliqui consiliatores eorum Dinei et Apharsathei Terphalei Apharsei Erchuei Babylonii Susannechei Deaei Aelamitae
EZRA|4|10|et ceteri de gentibus quas transtulit Asennaphar magnus et gloriosus et habitare eas fecit in civitatibus Samariae et in reliquis regionibus trans Flumen in pace
EZRA|4|11|hoc est exemplar epistulae quam miserunt ad eum Artarxersi regi servi tui viri qui sunt trans Fluvium salutem dicunt
EZRA|4|12|notum sit regi quia Iudaei qui ascenderunt a te ad nos venerunt in Hierusalem civitatem rebellem et pessimam quam aedificant extruentes muros eius et parietes conponentes
EZRA|4|13|nunc igitur notum sit regi quia si civitas illa aedificata fuerit et muri eius instaurati tributum et vectigal et annuos reditus non dabunt et usque ad reges haec noxa perveniet
EZRA|4|14|nos ergo memores salis quod in palatio comedimus et quia laesiones regis videre nefas ducimus idcirco misimus et nuntiavimus regi
EZRA|4|15|ut recenseas in libris historiarum patrum tuorum et invenies scriptum in commentariis et scies quoniam urbs illa urbs rebellis est et nocens regibus et provinciis et bella concitant in ea ex diebus antiquis quam ob rem et civitas ipsa destructa est
EZRA|4|16|nuntiamus nos regi quoniam si civitas illa aedificata fuerit et muri ipsius instaurati possessionem trans Fluvium non habebis
EZRA|4|17|verbum misit rex ad Reum Beelteem et Samsai scribam et ad reliquos qui erant in consilio eorum habitatores Samariae et ceteris trans Fluvium salutem dicens et pacem
EZRA|4|18|accusationem quam misistis ad nos manifeste lecta est coram me
EZRA|4|19|et a me praeceptum est et recensuerunt inveneruntque quoniam civitas illa a diebus antiquis adversum reges rebellat et seditiones et proelia concitantur in ea
EZRA|4|20|nam et reges fortissimi fuerunt in Hierusalem qui et dominati sunt omni regioni quae trans Fluvium est tributum quoque et vectigal et reditus accipiebant
EZRA|4|21|nunc ergo audite sententiam ut prohibeatis viros illos et urbs illa non aedificetur donec si forte a me iussum fuerit
EZRA|4|22|videte ne neglegenter hoc impleatis et paulatim crescat malum contra reges
EZRA|4|23|itaque exemplum edicti Artarxersis regis lectum est coram Reum et Samsai scriba et consiliariis eorum et abierunt festini in Hierusalem ad Iudaeos et prohibuerunt eos in brachio et robore
EZRA|4|24|tunc intermissum est opus domus Dei in Hierusalem et non fiebat usque ad annum secundum regni Darii regis Persarum
EZRA|5|1|prophetaverunt autem Aggeus propheta et Zaccharias filius Addo prophetantes ad Iudaeos qui erant in Iudaea et Hierusalem in nomine Dei Israhel
EZRA|5|2|tunc surrexerunt Zorobabel filius Salathihel et Iosue filius Iosedech et coeperunt aedificare templum Dei in Hierusalem et cum eis prophetae Dei adiuvantes eos
EZRA|5|3|in ipso tempore venit ad eos Tatannai qui erat dux trans Flumen et Starbuzannai et consiliarii eorum sicque dixerunt eis quis dedit vobis consilium ut domum hanc aedificaretis et muros hos instauraretis
EZRA|5|4|ad quod respondimus eis quae essent nomina hominum auctorum illius aedificationis
EZRA|5|5|oculus autem Dei eorum factus est super senes Iudaeorum et non potuerunt inhibere eos placuitque ut res ad Darium referretur et tunc satisfacerent adversus accusationem illam
EZRA|5|6|exemplar epistulae quam misit Tatannai dux regionis trans Flumen et Starbuzannai et consiliatores eius Apharsacei qui erant trans Flumen ad Darium regem
EZRA|5|7|sermo quem miserant ei sic scriptus erat Dario regi pax omnis
EZRA|5|8|notum sit regi isse nos ad Iudaeam provinciam ad domum Dei magni quae aedificatur lapide inpolito et ligna ponuntur in parietibus opusque illud diligenter extruitur et crescit in manibus eorum
EZRA|5|9|interrogavimus ergo senes illos et ita diximus eis quis dedit vobis potestatem ut domum hanc aedificaretis et muros instauraretis
EZRA|5|10|sed et nomina eorum quaesivimus ab eis ut nuntiaremus tibi quae scripsimus nomina virorum qui sunt principes in eis
EZRA|5|11|huiuscemodi autem sermonem responderunt nobis dicentes nos sumus servi Dei caeli et terrae et aedificamus templum quod erat extructum ante hos annos multos quodque rex Israhel magnus aedificaverat et extruxerat
EZRA|5|12|postquam autem ad iracundiam provocaverunt patres nostri Deum caeli et tradidit eos in manu Nabuchodonosor regis Babylonis Chaldei domum quoque hanc destruxit et populum eius transtulit in Babylonem
EZRA|5|13|anno autem primo Cyri regis Babylonis Cyrus rex proposuit edictum ut domus Dei aedificaretur
EZRA|5|14|nam et vasa templi Dei aurea et argentea quae Nabuchodonosor tulerat de templo quod erat in Hierusalem et asportaverat ea in templum Babylonis protulit Cyrus rex de templo Babylonis et data sunt Sasabassar vocabulo quem et principem constituit
EZRA|5|15|dixitque ei haec vasa tolle et vade et pone ea in templo quod est in Hierusalem et domus Dei aedificetur in loco suo
EZRA|5|16|tunc itaque Sasabassar ille venit et posuit fundamenta templi Dei in Hierusalem et ex eo tempore usque nunc aedificatur et necdum conpletum est
EZRA|5|17|nunc ergo si videtur regi bonum recenseat in bibliotheca regis quae est in Babylone utrumnam a Cyro rege iussum sit ut aedificaretur domus Dei in Hierusalem et voluntatem regis super hac re mittat ad nos
EZRA|6|1|tunc Darius rex praecepit et recensuerunt in bibliotheca librorum qui erant repositi in Babylone
EZRA|6|2|et inventum est in Ecbathanis quod est castrum in Madena provincia volumen unum talisque scriptus erat in eo commentarius
EZRA|6|3|anno primo Cyri regis Cyrus rex decrevit ut domus Dei quae est in Hierusalem aedificaretur in loco ubi immolent hostias et ut ponant fundamenta subportantia altitudinem cubitorum sexaginta et latitudinem cubitorum sexaginta
EZRA|6|4|ordines de lapidibus inpolitis tres et sic ordines de lignis novis sumptus autem de domo regis dabuntur
EZRA|6|5|sed et vasa templi Dei aurea et argentea quae Nabuchodonosor tulerat de templo Hierusalem et adtulerat ea in Babylonem reddantur et referantur in templo Hierusalem in locum suum quae et posita sunt in templo Dei
EZRA|6|6|nunc ergo Tatannai dux regionis quae est trans Flumen Starbuzannai et consiliarii vestri Apharsacei qui estis trans Flumen procul recedite ab illis
EZRA|6|7|et dimittite fieri templum Dei illud a duce Iudaeorum et a senioribus eorum domum Dei illam aedificent in loco suo
EZRA|6|8|sed et a me praeceptum est quid oporteat fieri a presbyteris Iudaeorum illis ut aedificetur domus Dei scilicet ut de arca regis id est de tributis quae dantur de regione trans Flumen studiose sumptus dentur viris illis ne inpediatur opus
EZRA|6|9|quod si necesse fuerit et vitulos et agnos et hedos in holocaustum Deo caeli frumentum sal vinum et oleum secundum ritum sacerdotum qui sunt in Hierusalem detur eis per dies singulos ne sit in aliquo querimonia
EZRA|6|10|et offerant oblationes Deo caeli orentque pro vita regis et filiorum eius
EZRA|6|11|a me ergo positum est decretum ut omnis homo qui hanc mutaverit iussionem tollatur lignum de domo ipsius et erigatur et configatur in eo domus autem eius publicetur
EZRA|6|12|Deus autem qui habitare fecit nomen suum ibi dissipet omnia regna et populum qui extenderit manum suam ut repugnet et dissipet domum Dei illam quae est in Hierusalem ego Darius statui decretum quod studiose impleri volo
EZRA|6|13|igitur Tatannai dux regionis trans Flumen et Starbuzannai et consiliarii eius secundum quod praeceperat Darius rex sic diligenter exsecuti sunt
EZRA|6|14|seniores autem Iudaeorum aedificabant et prosperabantur iuxta prophetiam Aggei prophetae et Zacchariae filii Addo et aedificaverunt et construxerunt iubente Deo Israhel et iubente Cyro et Dario et Artarxerse regibus Persarum
EZRA|6|15|et conpleverunt domum Dei istam usque ad diem tertium mensis adar qui est annus sextus regni Darii regis
EZRA|6|16|fecerunt autem filii Israhel sacerdotes et Levitae et reliqui filiorum transmigrationis dedicationem domus Dei in gaudio
EZRA|6|17|et obtulerunt in dedicationem domus Dei vitulos centum arietes ducentos agnos quadringentos hircos caprarum pro peccato totius Israhel duodecim iuxta numerum tribuum Israhel
EZRA|6|18|et statuerunt sacerdotes in ordinibus suis et Levitas in vicibus suis super opera Dei in Hierusalem sicut scriptum est in libro Mosi
EZRA|6|19|fecerunt autem filii transmigrationis pascha quartadecima die mensis primi
EZRA|6|20|purificati enim fuerant sacerdotes et Levitae quasi unus omnes mundi ad immolandum pascha universis filiis transmigrationis et fratribus suis sacerdotibus et sibi
EZRA|6|21|et comederunt filii Israhel qui reversi fuerant de transmigratione et omnis qui se separaverat a coinquinatione gentium terrae ad eos ut quaererent Dominum Deum Israhel
EZRA|6|22|et fecerunt sollemnitatem azymorum septem diebus in laetitia quoniam laetificaverat eos Dominus et converterat cor regis Assur ad eos ut adiuvaret manus eorum in opere domus Domini Dei Israhel
EZRA|7|1|post haec autem verba in regno Artarxersis regis Persarum Ezras filius Saraiae filii Azariae filii Helciae
EZRA|7|2|filii Sellum filii Sadoc filii Achitob
EZRA|7|3|filii Amariae filii Azariae filii Maraioth
EZRA|7|4|filii Zaraiae filii Ozi filii Bocci
EZRA|7|5|filii Abisue filii Finees filii Eleazar filii Aaron sacerdotis ab initio
EZRA|7|6|ipse Ezras ascendit de Babylone et ipse scriba velox in lege Mosi quam dedit Dominus Deus Israhel et dedit ei rex secundum manum Domini Dei eius super eum omnem petitionem eius
EZRA|7|7|et ascenderunt de filiis Israhel et de filiis sacerdotum et de filiis Levitarum et de cantoribus et de ianitoribus et de Nathinneis in Hierusalem anno septimo Artarxersis regis
EZRA|7|8|et venerunt in Hierusalem mense quinto ipse est annus septimus regis
EZRA|7|9|quia in primo die mensis primi coepit ascendere de Babylone et in primo mensis quinti venit in Hierusalem iuxta manum Dei sui bonam super se
EZRA|7|10|Ezras enim paravit cor suum ut investigaret legem Domini et faceret et doceret in Israhel praeceptum et iudicium
EZRA|7|11|hoc est autem exemplar epistulae edicti quod dedit rex Artarxersis Ezrae sacerdoti scribae erudito in sermonibus et praeceptis Domini et caerimoniis eius in Israhel
EZRA|7|12|Artarxersis rex regum Ezrae sacerdoti scribae legis Dei caeli doctissimo salutem
EZRA|7|13|a me decretum est ut cuicumque placuerit in regno meo de populo Israhel et de sacerdotibus eius et de Levitis ire in Hierusalem tecum vadat
EZRA|7|14|a facie enim regis et septem consiliatorum eius missus es ut visites Iudaeam et Hierusalem in lege Dei tui quae est in manu tua
EZRA|7|15|et ut feras argentum et aurum quod rex et consiliatores eius sponte obtulerunt Deo Israhel cuius in Hierusalem tabernaculum est
EZRA|7|16|et omne argentum et aurum quodcumque inveneris in universa provincia Babylonis et populus offerre voluerit et de sacerdotibus qui sponte obtulerint domui Dei sui quae est in Hierusalem
EZRA|7|17|libere accipe et studiose eme de hac pecunia vitulos arietes agnos et sacrificia et libamina eorum et offer ea super altare templi Dei vestri quod est in Hierusalem
EZRA|7|18|sed et si quid tibi et fratribus tuis placuerit de reliquo argento et auro ut faciatis iuxta voluntatem Dei vestri facite
EZRA|7|19|vasa quoque quae dantur tibi in ministerium domus Dei tui trade in conspectu Dei Hierusalem
EZRA|7|20|sed et cetera quibus opus fuerit in domo Dei tui quantumcumque necesse est ut expendas dabis de thesauro et de fisco regis
EZRA|7|21|et a me ego Artarxersis rex statui atque decrevi omnibus custodibus arcae publicae qui sunt trans Flumen ut quodcumque petierit a vobis Ezras sacerdos scriba legis Dei caeli absque mora detis
EZRA|7|22|usque ad argenti talenta centum et usque ad frumenti choros centum et usque ad vini batos centum et usque ad batos olei centum sal vero absque mensura
EZRA|7|23|omne quod ad ritum Dei caeli pertinet tribuatur diligenter in domo Dei caeli ne forte irascatur contra regnum regis et filiorum eius
EZRA|7|24|vobisque notum facimus de universis sacerdotibus et Levitis cantoribus ianitoribus Nathinneis et ministris domus Dei huius ut vectigal et tributum et annonas non habeatis potestatem inponendi super eos
EZRA|7|25|tu autem Ezras secundum sapientiam Dei tui quae est in manu tua constitue iudices et praesides ut iudicent omni populo qui est trans Flumen his videlicet qui noverunt legem Dei tui sed et inperitos docete libere
EZRA|7|26|et omnis qui non fecerit legem Dei tui et legem regis diligenter iudicium erit de eo sive in mortem sive in exilium sive in condemnationem substantiae eius vel certe in carcerem
EZRA|7|27|benedictus Dominus Deus patrum nostrorum qui dedit hoc in corde regis ut glorificaret domum Domini quae est in Hierusalem
EZRA|7|28|et in me inclinavit misericordiam coram rege et consiliatoribus eius et universis principibus regis potentibus et ego confortatus manu Domini Dei mei quae erat in me congregavi de Israhel principes qui ascenderent mecum
EZRA|8|1|hii sunt ergo principes familiarum et genealogia eorum qui ascenderunt mecum in regno Artarxersis regis de Babylone
EZRA|8|2|de filiis Finees Gersom de filiis Ithamar Danihel de filiis David Attus
EZRA|8|3|de filiis Secheniae et de filiis Pharos Zaccharias et cum eo numerati sunt viri centum quinquaginta
EZRA|8|4|de filiis Phaethmoab Helioenai filius Zareae et cum eo ducenti viri
EZRA|8|5|de filiis Secheniae filius Hiezihel et cum eo trecenti viri
EZRA|8|6|de filiis Adden Abeth filius Ionathan et cum eo quinquaginta viri
EZRA|8|7|de filiis Helam Isaias filius Athaliae et cum eo septuaginta viri
EZRA|8|8|de filiis Saphatiae Zebedia filius Michahel et cum eo octoginta viri
EZRA|8|9|de filiis Ioab Obedia filius Iehihel et cum eo ducenti decem et octo viri
EZRA|8|10|de filiis Selomith filius Iosphiae et cum eo centum sexaginta viri
EZRA|8|11|de filiis Bebai Zaccharias filius Bebai et cum eo viginti octo viri
EZRA|8|12|de filiis Ezgad Iohanan filius Eccetan et cum eo centum decem viri
EZRA|8|13|de filiis Adonicam qui erant novissimi et haec nomina eorum Helifeleth et Heihel et Samaias et cum eis sexaginta viri
EZRA|8|14|de filiis Beggui Uthai et Zacchur et cum eo septuaginta viri
EZRA|8|15|congregavi autem eos ad fluvium qui decurrit ad Ahavva et mansimus ibi diebus tribus quaesivique in populo et in sacerdotibus de filiis Levi et non inveni ibi
EZRA|8|16|itaque misi Heliezer et Arihel et Semeam et Helnathan et Iarib et alterum Helnathan et Nathan et Zacchariam et Mesolam principes et Ioarib et Helnathan sapientes
EZRA|8|17|et misi eos ad Heddo qui est primus in Casphiae loco et posui in ore eorum verba quae loquerentur ad Addom et ad fratres eius Nathinneos in loco Casphiae ut adducerent nobis ministros domus Dei nostri
EZRA|8|18|et adduxerunt nobis per manum Dei nostri bonam super nos virum doctissimum de filiis Moolli filii Levi filii Israhel et Sarabiam et filios eius et fratres eius decem et octo
EZRA|8|19|et Asabiam et cum eo Isaiam de filiis Merari fratres eius et filios eius viginti
EZRA|8|20|et de Nathinneis quos dederat David et principes ad ministeria Levitarum Nathinneos ducentos viginti omnes hii suis nominibus vocabantur
EZRA|8|21|et praedicavi ibi ieiunium iuxta fluvium Ahavva ut adfligeremur coram Domino Deo nostro et peteremus ab eo viam rectam nobis et filiis nostris universaeque substantiae nostrae
EZRA|8|22|erubui enim petere regem auxilium et equites qui defenderent nos ab inimico in via quia dixeramus regi manus Dei nostri est super omnes qui quaerunt eum in bonitate et imperium eius et fortitudo eius et furor super omnes qui derelinquunt eum
EZRA|8|23|ieiunavimus autem et rogavimus Deum nostrum pro hoc et evenit nobis prospere
EZRA|8|24|et separavi de principibus sacerdotum duodecim Sarabian Asabian et cum eis de fratribus eorum decem
EZRA|8|25|adpendique eis argentum et aurum et vasa consecrata domus Dei nostri quae obtulerat rex et consiliatores eius et principes eius universusque Israhel eorum qui inventi fuerant
EZRA|8|26|et adpendi in manibus eorum argenti talenta sescenta quinquaginta et vasa argentea centum auri centum talenta
EZRA|8|27|et crateras aureos viginti qui habebant solidos millenos et vasa aeris fulgentis optimi duo pulchra ut aurum
EZRA|8|28|et dixi eis vos sancti Domini et vasa sancta et argentum et aurum quod sponte oblatum est Domino Deo patrum vestrorum
EZRA|8|29|vigilate et custodite donec adpendatis coram principibus sacerdotum et Levitarum et ducibus familiarum Israhel in Hierusalem et thesaurum domus Domini
EZRA|8|30|susceperunt autem sacerdotes et Levitae pondus argenti et auri et vasorum ut deferrent in Hierusalem in domum Dei nostri
EZRA|8|31|promovimus ergo a flumine Ahavva duodecimo die mensis primi ut pergeremus Hierusalem et manus Dei nostri fuit super nos et liberavit nos de manu inimici et insidiatoris in via
EZRA|8|32|et venimus Hierusalem et mansimus ibi diebus tribus
EZRA|8|33|die autem quarta adpensum est argentum et aurum et vasa in domo Dei nostri per manum Meremoth filii Uriae sacerdotis et cum eo Eleazar filius Finees cumque eis Iozaded filius Iosue et Noadaia filius Bennoi Levitae
EZRA|8|34|iuxta numerum et pondus omnium descriptumque est omne pondus in tempore illo
EZRA|8|35|sed et qui venerant de captivitate filii transmigrationis obtulerunt holocaustomata Deo Israhel vitulos duodecim pro omni Israhel arietes nonaginta sex agnos septuaginta septem hircos pro peccato duodecim omnia in holocaustum Domino
EZRA|8|36|dederunt autem edicta regis satrapis qui erant de conspectu regis et ducibus trans Flumen et elevaverunt populum et domum Dei
EZRA|9|1|postquam autem haec conpleta sunt accesserunt ad me principes dicentes non est separatus populus Israhel et sacerdotes et Levitae a populis terrarum et de abominationibus eorum Chananei videlicet et Hetthei et Ferezei et Iebusei et Ammanitarum et Moabitarum et Aegyptiorum et Amorreorum
EZRA|9|2|tulerunt enim de filiabus eorum sibi et filiis suis et commiscuerunt semen sanctum cum populis terrarum manus etiam principum et magistratuum fuit in transgressione hac prima
EZRA|9|3|cumque audissem sermonem istum scidi pallium meum et tunicam et evelli capillos capitis mei et barbae et sedi maerens
EZRA|9|4|convenerunt autem ad me omnes qui timebant verbum Dei Israhel pro transgressione eorum qui de captivitate venerant et ego sedebam tristis usque ad sacrificium vespertinum
EZRA|9|5|et in sacrificio vespertino surrexi de adflictione mea et scisso pallio et tunica curvavi genua mea et expandi manus meas ad Dominum Deum meum
EZRA|9|6|et dixi Deus meus confundor et erubesco levare Deus meus faciem meam ad te quoniam iniquitates nostrae multiplicatae sunt super caput et delicta nostra creverunt usque in caelum
EZRA|9|7|a diebus patrum nostrorum sed et nos ipsi peccavimus granditer usque ad diem hanc et in iniquitatibus nostris traditi sumus ipsi et reges nostri et sacerdotes nostri in manum regum terrarum in gladium in captivitatem in rapinam et in confusionem vultus sicut et die hac
EZRA|9|8|et nunc quasi parum et ad momentum facta est deprecatio nostra apud Dominum Deum nostrum ut dimitterentur nobis reliquiae et daretur paxillus in loco sancto eius et inluminaret oculos nostros Deus noster et daret nobis vitam modicam in servitute nostra
EZRA|9|9|quia servi sumus et in servitute nostra non dereliquit nos Deus noster et inclinavit super nos misericordiam coram rege Persarum ut daret nobis vitam et sublimaret domum Dei nostri et extrueret solitudines eius et daret nobis sepem in Iuda et in Hierusalem
EZRA|9|10|et nunc quid dicemus Deus noster post haec quia dereliquimus mandata tua
EZRA|9|11|quae praecepisti in manu servorum tuorum prophetarum dicens terram ad quam vos ingredimini ut possideatis eam terra inmunda est iuxta inmunditiam populorum ceterarumque terrarum abominationibus eorum qui repleverunt eam ab ore usque ad os in coinquinatione sua
EZRA|9|12|nunc ergo filias vestras ne detis filiis eorum et filias eorum non accipiatis filiis vestris et non quaeratis pacem eorum et prosperitatem eorum usque in aeternum ut confortemini et comedatis quae bona sunt terrae et heredes habeatis filios vestros usque in saeculum
EZRA|9|13|et post omnia quae venerunt super nos in operibus nostris pessimis et in delicto nostro magno quia tu Deus noster liberasti nos de iniquitate nostra et dedisti nobis salutem sicut est hodie
EZRA|9|14|ut non converteremur et irrita faceremus mandata tua neque matrimonia iungeremus cum populis abominationum istarum numquid iratus es nobis usque ad consummationem ne dimitteres nobis reliquias et salutem
EZRA|9|15|Domine Deus Israhel iustus tu quoniam derelicti sumus qui salvaremur sicut die hac ecce coram te sumus in delicto nostro non enim stari potest coram te super hoc
EZRA|10|1|sic ergo orante Ezra et inplorante eo et flente et iacente ante templum Dei collectus est ad eum de Israhel coetus grandis nimis virorum et mulierum puerorumque et flevit populus multo fletu
EZRA|10|2|et respondit Sechenia filius Iehihel de filiis Helam et dixit Ezrae nos praevaricati sumus in Deum nostrum et duximus uxores alienigenas de populis terrae et nunc si est paenitentia Israhel super hoc
EZRA|10|3|percutiamus foedus cum Deo nostro ut proiciamus universas uxores et eos qui de his nati sunt iuxta voluntatem Domini et eorum qui timent praeceptum Dei nostri secundum legem fiat
EZRA|10|4|surge tuum est decernere nosque erimus tecum confortare et fac
EZRA|10|5|surrexit ergo Ezras et adiuravit principes sacerdotum Levitarum et omnem Israhel ut facerent secundum verbum hoc et iuraverunt
EZRA|10|6|et surrexit Ezras ante domum Dei et abiit ad cubiculum Iohanan filii Eliasib et ingressus est illuc panem non comedit et aquam non bibit lugebat enim in transgressione eorum qui de captivitate venerant
EZRA|10|7|et missa est vox in Iuda et in Hierusalem omnibus filiis transmigrationis ut congregarentur in Hierusalem
EZRA|10|8|et omnis qui non venerit in tribus diebus iuxta consilium principum et seniorum auferetur universa substantia eius et ipse abicietur de coetu transmigrationis
EZRA|10|9|convenerunt igitur omnes viri Iuda et Beniamin in Hierusalem tribus diebus ipse est mensis nonus vicesimo die mensis et sedit omnis populus in platea domus Dei trementes pro peccato et pluviis
EZRA|10|10|et surrexit Ezras sacerdos et dixit ad eos vos transgressi estis et duxistis uxores alienigenas ut adderetis super delictum Israhel
EZRA|10|11|et nunc date confessionem Domino Deo patrum vestrorum et facite placitum eius et separamini a populis terrae et ab uxoribus alienigenis
EZRA|10|12|et respondit universa multitudo dixitque voce magna iuxta verbum tuum ad nos sic fiat
EZRA|10|13|verumtamen quia populus multus est et tempus pluviae et non sustinemus stare foris et opus non est diei unius vel duorum vehementer quippe peccavimus in sermone isto
EZRA|10|14|constituantur principes in universa multitudine et omnes in civitatibus nostris qui duxerunt uxores alienigenas veniant in temporibus statutis et cum his seniores per civitatem et civitatem et iudices eius donec avertatur ira Dei nostri a nobis super peccato hoc
EZRA|10|15|igitur Ionathan filius Asahel et Iaazia filius Thecuae steterunt super hoc et Mesollam et Sebethai Levites adiuverunt eos
EZRA|10|16|feceruntque sic filii transmigrationis et abierunt Ezras sacerdos et viri principes familiarum in domum patrum suorum et omnes per nomina sua et sederunt in die primo mensis decimi ut quaererent rem
EZRA|10|17|et consummati sunt omnes viri qui duxerant uxores alienigenas usque ad diem primam mensis primi
EZRA|10|18|et inventi sunt de filiis sacerdotum qui duxerant uxores alienigenas de filiis Iosue filii Iosedech et fratres eius Maasia et Eliezer et Iarib et Godolia
EZRA|10|19|et dederunt manus suas ut eicerent uxores suas et pro delicto suo arietem de ovibus offerrent
EZRA|10|20|et de filiis Emmer Anani et Zebedia
EZRA|10|21|et de filiis Erim Masia et Helia et Semeia et Hiehihel et Ozias
EZRA|10|22|et de filiis Phessur Helioenai Maasia Ismahel Nathanahel Iozabeth et Elasa
EZRA|10|23|et de filiis Levitarum Iozabeth et Semei et Celaia ipse est Calita Phataia Iuda et Eliezer
EZRA|10|24|et de cantoribus Eliasub et de ianitoribus Sellum et Telem et Uri
EZRA|10|25|et ex Israhel de filiis Pharos Remia et Ezia et Melchia et Miamin et Eliezer et Melchia et Banea
EZRA|10|26|et de filiis Helam Mathania Zaccharias et Hiehil et Abdi et Irimoth et Helia
EZRA|10|27|et de filiis Zethua Helioenai Eliasib Mathania et Ierimuth et Zabeth et Aziza
EZRA|10|28|et de filiis Bebai Iohanan Anania Zabbai Athalai
EZRA|10|29|et de filiis Bani Mosollam et Melluch et Adaia Iasub et Saal et Ramoth
EZRA|10|30|et de filiis Phaethmoab Edna et Chalal Banaias Maasias Mathanias Beselehel et Bennui et Manasse
EZRA|10|31|et de filiis Erem Eliezer Iesue Melchias Semeias Symeon
EZRA|10|32|Beniamin Maloch Samarias
EZRA|10|33|de filiis Asom Matthanai Matthetha Zabed Elipheleth Iermai Manasse Semei
EZRA|10|34|de filiis Bani Maaddi Amram et Huhel
EZRA|10|35|Baneas et Badaias Cheiliau
EZRA|10|36|Vannia Marimuth et Eliasib
EZRA|10|37|Matthanias Mathanai et Iasi
EZRA|10|38|et Bani et Bennui Semei
EZRA|10|39|et Salmias et Nathan et Adaias
EZRA|10|40|Mechnedabai Sisai Sarai
EZRA|10|41|Ezrel et Selemau Semeria
EZRA|10|42|Sellum Amaria Ioseph
EZRA|10|43|de filiis Nebu Iaihel Matthathias Zabed Zabina Ieddu et Iohel Banaia
EZRA|10|44|omnes hii acceperunt uxores alienigenas et fuerunt ex eis mulieres quae pepererant filios
NEH|1|1|verba Neemiae filii Echliae et factum est in mense casleu anno vicesimo et ego eram in Susis castro
NEH|1|2|et venit Anani unus de fratribus meis ipse et viri ex Iuda et interrogavi eos de Iudaeis qui remanserant et supererant de captivitate et de Hierusalem
NEH|1|3|et dixerunt mihi qui remanserunt et derelicti sunt de captivitate ibi in provincia in adflictione magna sunt et in obprobrio et murus Hierusalem dissipatus est et portae eius conbustae sunt igni
NEH|1|4|cumque audissem verba huiuscemodi sedi et flevi et luxi diebus et ieiunabam et orabam ante faciem Dei caeli
NEH|1|5|et dixi quaeso Domine Deus caeli fortis magne atque terribilis qui custodis pactum et misericordiam cum his qui te diligunt et custodiunt mandata tua
NEH|1|6|fiat auris tua auscultans et oculi tui aperti ut audias orationem servi tui quam ego oro coram te hodie nocte et die pro filiis Israhel servis tuis et confiteor pro peccatis filiorum Israhel quibus peccaverunt tibi et ego et domus patris mei peccavimus
NEH|1|7|vanitate seducti sumus et non custodivimus mandatum et caerimonias et iudicia quae praecepisti Mosi servo tuo
NEH|1|8|memento verbi quod mandasti Mosi famulo tuo dicens cum transgressi fueritis ego dispergam vos in populos
NEH|1|9|et si revertamini ad me et custodiatis mandata mea et faciatis ea etiam si abducti fueritis ad extrema caeli inde congregabo vos et inducam in locum quem elegi ut habitaret nomen meum ibi
NEH|1|10|et ipsi servi tui et populus tuus quos redemisti in fortitudine tua magna et in manu tua valida
NEH|1|11|obsecro Domine sit auris tua adtendens ad orationem servi tui et ad orationem servorum tuorum qui volunt timere nomen tuum et dirige servum tuum hodie et da ei misericordiam ante virum hunc ego enim eram pincerna regis
NEH|2|1|factum est autem in mense nisan anno vicesimo Artarxersis regis et vinum erat ante eum et levavi vinum et dedi regi et non eram quasi languidus ante faciem eius
NEH|2|2|dixitque mihi rex quare vultus tuus tristis cum te aegrotum non videam non est hoc frustra sed malum nescio quid in corde tuo est et timui valde ac nimis
NEH|2|3|et dixi regi rex in aeternum vive quare non maereat vultus meus quia civitas domus sepulchrorum patris mei deserta est et portae eius conbustae sunt igni
NEH|2|4|et ait mihi rex pro qua re postulas et oravi Deum caeli
NEH|2|5|et dixi ad regem si videtur regi bonum et si placet servus tuus ante faciem tuam ut mittas me in Iudaeam ad civitatem sepulchri patris mei et aedificabo eam
NEH|2|6|dixitque mihi rex et regina quae sedebat iuxta eum usque ad quod tempus erit iter tuum et quando reverteris et placuit ante vultum regis et misit me et constitui ei tempus
NEH|2|7|et dixi regi si regi videtur bonum epistulas det mihi ad duces regionis trans Flumen ut transducant me donec veniam in Iudaeam
NEH|2|8|et epistulam ad Asaph custodem saltus regis ut det mihi ligna et tegere possim portas turris domus et muri civitatis et domum quam ingressus fuero et dedit mihi rex iuxta manum Dei mei bonam mecum
NEH|2|9|et veni ad duces regionis trans Flumen dedique eis epistulas regis miserat autem mecum rex principes militum et equites
NEH|2|10|et audierunt Sanaballat Horonites et Tobias servus ammanites et contristati sunt adflictione magna quod venisset homo qui quaereret prosperitatem filiorum Israhel
NEH|2|11|et veni Hierusalem et eram ibi diebus tribus
NEH|2|12|et surrexi nocte ego et viri pauci mecum et non indicavi cuiquam quid Deus dedisset in corde meo ut facerem in Hierusalem et iumentum non erat mecum nisi animal cui sedebam
NEH|2|13|et egressus sum per portam Vallis nocte et ante fontem Draconis et ad portam Stercoris et considerabam murum Hierusalem dissipatum et portas eius consumptas igni
NEH|2|14|et transivi ad portam Fontis et ad aquaeductum Regis et non erat locus iumento cui sedebam ut transiret
NEH|2|15|et ascendi per torrentem nocte et considerabam murum et reversus veni ad portam Vallis et redii
NEH|2|16|magistratus autem nesciebant quo abissem aut quid ego facerem sed et Iudaeis et sacerdotibus et optimatibus et magistratibus et reliquis qui faciebant opus usque ad id locorum nihil indicaveram
NEH|2|17|et dixi eis vos nostis adflictionem in qua sumus quia Hierusalem deserta est et portae eius consumptae sunt igni venite et aedificemus muros Hierusalem et non simus ultra obprobrium
NEH|2|18|et indicavi eis manum Dei mei quod esset bona mecum et verba regis quae locutus est mihi et aio surgamus et aedificemus et confortatae sunt manus eorum in bono
NEH|2|19|audierunt autem Sanaballat Horonites et Tobias servus ammanites et Gosem Arabs et subsannaverunt nos et despexerunt dixeruntque quae est haec res quam facitis numquid contra regem vos rebellatis
NEH|2|20|et reddidi eis sermonem dixique ad eos Deus caeli ipse nos iuvat et nos servi eius sumus surgamus et aedificemus vobis autem non est pars et iustitia et memoria in Hierusalem
NEH|3|1|et surrexit Eliasib sacerdos magnus et fratres eius sacerdotes et aedificaverunt portam Gregis ipsi sanctificaverunt eam et statuerunt valvas eius et usque ad turrem centum cubitorum sanctificaverunt eam usque ad turrem Ananehel
NEH|3|2|et iuxta eum aedificaverunt viri Hiericho et iuxta eum aedificavit Zecchur filius Amri
NEH|3|3|portam autem Piscium aedificaverunt filii Asanaa ipsi texerunt eam et statuerunt valvas eius et seras et vectes et iuxta eos aedificavit Marimuth filius Uriae filii Accus
NEH|3|4|et iuxta eos aedificavit Mosollam filius Barachiae filii Mesezebel et iuxta eos aedificavit Sadoc filius Baana
NEH|3|5|et iuxta eos aedificaverunt Thecueni optimates autem eorum non subposuerunt colla sua in opere Domini sui
NEH|3|6|et portam Veterem aedificaverunt Ioiada filius Fasea et Mosollam filius Besodia ipsi texerunt eam et statuerunt valvas eius et seras et vectes
NEH|3|7|et iuxta eos aedificavit Meletias Gabaonites et Iadon Meronathites viri de Gabaon et Maspha pro duce qui erat in regione trans Flumen
NEH|3|8|et iuxta eum aedificavit Ezihel filius Araia aurifex et iuxta eum aedificavit Anania filius pigmentarii et dimiserunt Hierusalem usque ad murum plateae latioris
NEH|3|9|et iuxta eum aedificavit Rafaia filius Ahur princeps vici Hierusalem
NEH|3|10|et iuxta eos aedificavit Ieiada filius Aromath contra domum suam et iuxta eum aedificavit Attus filius Asebeniae
NEH|3|11|mediam partem vici aedificavit Melchias filius Erem et Asub filius Phaethmoab et turrem Furnorum
NEH|3|12|iuxta eum aedificavit Sellum filius Alloes princeps mediae partis vici Hierusalem ipse et filiae eius
NEH|3|13|et portam Vallis aedificavit Anun et habitatores Zanoe ipsi aedificaverunt eam et statuerunt valvas eius et seras et vectes et mille cubitos in muro usque ad portam Sterquilinii
NEH|3|14|et portam Sterquilinii aedificavit Melchias filius Rechab princeps vici Bethaccharem ipse aedificavit eam et statuit valvas eius et seras et vectes
NEH|3|15|et portam Fontis aedificavit Sellum filius Choloozai princeps pagi Maspha ipse aedificavit eam et texit et statuit valvas eius et seras et vectes et muros piscinae Siloae in hortum regis et usque ad gradus qui descendunt de civitate David
NEH|3|16|post eum aedificavit Neemias filius Azboc princeps dimidiae partis vici Bethsur usque contra sepulchra David et usque ad piscinam quae grandi opere constructa est et usque ad domum Fortium
NEH|3|17|post eum aedificaverunt Levitae Reum filius Benni post eum aedificavit Asebias princeps dimidiae partis vici Ceilae in vico suo
NEH|3|18|post eum aedificaverunt fratres eorum Behui filius Enadad princeps dimidiae partis Ceila
NEH|3|19|et aedificavit iuxta eum Azer filius Iosue princeps Maspha mensuram secundam contra ascensum firmissimi anguli
NEH|3|20|post eum in monte aedificavit Baruch filius Zacchai mensuram secundam ab angulo usque ad portam domus Eliasib sacerdotis magni
NEH|3|21|post eum aedificavit Meremuth filius Uriae filii Accus mensuram secundam a porta domus Eliasib donec extenderetur domus Eliasib
NEH|3|22|et post eum aedificaverunt sacerdotes viri de campestribus Iordanis
NEH|3|23|post eum aedificavit Beniamin et Asub contra domum suam et post eum aedificavit Azarias filius Maasiae filii Ananiae contra domum suam
NEH|3|24|post eum aedificavit Bennui filius Enadda mensuram secundam a domo Azariae usque ad flexuram et usque ad angulum
NEH|3|25|Falel filius Ozi contra flexuram et turrem quae eminet de domo regis excelsa id est in atrio carceris post eum Phadaia filius Pheros
NEH|3|26|Nathinnei autem habitabant in Ofel usque contra portam Aquarum ad orientem et turrem quae prominebat
NEH|3|27|post eum aedificaverunt Thecueni mensuram secundam e regione a turre magna et eminenti usque ad murum templi
NEH|3|28|sursum autem a porta Equorum aedificaverunt sacerdotes unusquisque contra domum suam
NEH|3|29|post eos aedificavit Seddo filius Emmer contra domum suam et post eum aedificavit Semeia filius Secheniae custos portae orientalis
NEH|3|30|post eum aedificavit Anania filius Selemiae et Anon filius Selo sextus mensuram secundam post eum aedificavit Mosollam filius Barachiae contra gazofilacium suum post eum aedificavit Melchias filius aurificis usque ad domum Nathinneorum et scruta vendentium contra portam Iudicialem et usque ad cenaculum Anguli
NEH|3|31|et inter cenaculum Anguli in porta Gregis aedificaverunt artifices et negotiatores
NEH|4|1|factum est autem cum audisset Sanaballat quod aedificaremus murum iratus est valde et motus nimis subsannavit Iudaeos
NEH|4|2|et dixit coram fratribus suis et frequentia Samaritanorum quid Iudaei inbecilli faciunt num dimittent eos gentes num sacrificabunt et conplebunt in una die numquid aedificare poterunt lapides de acervis pulveris qui conbusti sunt
NEH|4|3|sed et Tobias Ammanites proximus eius ait aedificent si ascenderit vulpis transiliet murum eorum lapideum
NEH|4|4|audi Deus noster quia facti sumus despectio converte obprobrium super caput eorum et da eos in despectionem in terra captivitatis
NEH|4|5|ne operias iniquitatem eorum et peccatum eorum coram facie tua non deleatur quia inriserunt aedificantes
NEH|4|6|itaque aedificavimus murum et coniunximus totum usque ad partem dimidiam et provocatum est cor populi ad operandum
NEH|4|7|factum est autem cum audisset Sanaballat et Tobias et Arabes et Ammanitae et Azotii quod obducta esset cicatrix muri Hierusalem et quod coepissent interrupta concludi irati sunt nimis
NEH|4|8|et congregati omnes pariter ut venirent et pugnarent contra Hierusalem et molirentur insidias
NEH|4|9|et oravimus Deum nostrum et posuimus custodes super murum die et nocte contra eos
NEH|4|10|dixit autem Iudas debilitata est fortitudo portantis et humus nimia est et nos non poterimus aedificare murum
NEH|4|11|et dixerunt hostes nostri nesciant et ignorent donec veniamus in medio eorum et interficiamus eos et cessare faciamus opus
NEH|4|12|factum est autem venientibus Iudaeis qui habitabant iuxta eos et dicentibus nobis per decem vices ex omnibus locis quibus venerant ad nos
NEH|4|13|statui in loco post murum per circuitum populum in ordine cum gladiis suis et lanceis et arcis
NEH|4|14|perspexi atque surrexi et aio ad optimates et ad magistratus et ad reliquam partem vulgi nolite timere a facie eorum Domini magni et terribilis mementote et pugnate pro fratribus vestris filiis vestris et filiabus vestris uxoribus vestris et domibus
NEH|4|15|factum est autem cum audissent inimici nostri nuntiatum esse nobis dissipavit Deus consilium eorum et reversi sumus omnes ad muros unusquisque ad opus suum
NEH|4|16|et factum est a die illa media pars iuvenum eorum faciebant opus et media parata erat ad bellum et lanceae et scuta et arcus et loricae et principes post eos in omni domo Iuda
NEH|4|17|aedificantium in muro et portantium onera et inponentium una manu sua faciebat opus et altera tenebat gladium
NEH|4|18|aedificantium enim unusquisque gladio erat accinctus renes et aedificabant et clangebant bucina iuxta me
NEH|4|19|et dixi ad optimates et ad magistratus et ad reliquam partem vulgi opus grande est et latum et nos separati sumus in muro procul alter ab altero
NEH|4|20|in loco quocumque audieritis clangorem tubae illuc concurrite ad nos Deus noster pugnabit pro nobis
NEH|4|21|et nos ipsi faciamus opus et media pars nostrum teneat lanceas ab ascensu aurorae donec egrediantur astra
NEH|4|22|in tempore quoque illo dixi populo unusquisque cum puero suo maneat in medio Hierusalem et sint vobis vices per noctem et diem ad operandum
NEH|4|23|ego autem et fratres mei et pueri mei et custodes qui erant post me non deponebamus vestimenta nostra unusquisque tantum nudabatur ad baptismum
NEH|5|1|et factus est clamor populi et uxorum eius magnus adversus fratres suos iudaeos
NEH|5|2|et erant qui dicerent filii nostri et filiae nostrae multae sunt nimis accipiamus pro pretio eorum frumentum et comedamus et vivamus
NEH|5|3|et erant qui dicerent agros nostros et vineas et domos nostras opponamus et accipiamus frumentum in fame
NEH|5|4|et alii dicebant mutuo sumamus pecunias in tributa regis demusque agros nostros et vineas
NEH|5|5|et nunc sicut carnes fratrum nostrorum sic carnes nostrae sunt sicut filii eorum ita filii nostri ecce nos subiugamus filios nostros et filias nostras in servitutem et de filiabus nostris sunt famulae nec habemus unde possint redimi et agros nostros et vineas alii possident
NEH|5|6|et iratus sum nimis cum audissem clamorem eorum secundum verba haec
NEH|5|7|cogitavitque cor meum mecum et increpui optimates et magistratus et dixi eis usurasne singuli a fratribus vestris exigatis et congregavi adversus eos contionem magnam
NEH|5|8|et dixi eis nos ut scitis redemimus fratres nostros iudaeos qui venditi fuerant gentibus secundum possibilitatem nostram et vos igitur vendite fratres vestros et emimus eos et siluerunt nec invenerunt quid responderent
NEH|5|9|dixique ad eos non est bona res quam facitis quare non in timore Dei nostri ambulatis ne exprobretur nobis a gentibus inimicis nostris
NEH|5|10|et ego et fratres mei et pueri mei commodavimus plurimis pecuniam et frumentum non repetamus in commune istud aes alienum concedamus quod debetur nobis
NEH|5|11|reddite eis hodie agros suos vineas suas oliveta sua et domos suas quin potius et centesimam pecuniae frumenti vini et olei quam exigere soletis ab eis date pro illis
NEH|5|12|et dixerunt reddimus et ab eis nihil quaerimus sicque faciemus ut loqueris et vocavi sacerdotes et adiuravi eos ut facerent iuxta quod dixeram
NEH|5|13|insuper et sinum meum excussi et dixi sic excutiat Deus omnem virum qui non conpleverit verbum istud de domo sua et de laboribus suis sic excutiatur et vacuus fiat et dixit universa multitudo amen et laudaverunt Deum fecit ergo populus sicut dictum erat
NEH|5|14|a die autem illa qua praeceperat mihi ut essem dux in terra Iuda ab anno vicesimo usque ad annum tricesimum secundum Artarxersis regis per annos duodecim ego et fratres mei annonas quae ducibus debebantur non comedimus
NEH|5|15|duces autem primi qui fuerant ante me gravaverunt populum et acceperunt ab eis in pane vino et pecunia cotidie siclos quadraginta sed et ministri eorum depresserant populum ego autem non feci ita propter timorem Dei
NEH|5|16|quin potius in opere muri aedificavi et agrum non emi et omnes pueri mei congregati ad opus erant
NEH|5|17|Iudaei quoque et magistratus centum quinquaginta viri et qui veniebant ad nos de gentibus quae in circuitu nostro sunt in mensa mea erant
NEH|5|18|parabatur autem mihi per dies singulos bos unus arietes sex electi exceptis volatilibus et inter dies decem vina diversa et alia multa tribuebam insuper et annonas ducatus mei non quaesivi valde enim erat adtenuatus populus
NEH|5|19|memento mei Deus meus in bonum secundum omnia quae feci populo huic
NEH|6|1|factum est autem cum audisset Sanaballat et Tobia et Gosem Arabs et ceteri inimici nostri quod aedificassem ego murum et non esset in ipso residua interruptio usque ad tempus autem illud valvas non posueram in portis
NEH|6|2|miserunt Sanaballat et Gosem ad me dicentes veni et percutiamus foedus pariter in viculis in campo Ono ipsi autem cogitabant ut facerent mihi malum
NEH|6|3|misi ergo ad eos nuntios dicens opus grande ego facio et non possum descendere ne forte neglegatur cum venero et descendero ad vos
NEH|6|4|miserunt autem ad me secundum verbum hoc per quattuor vices et respondi eis iuxta sermonem priorem
NEH|6|5|et misit ad me Sanaballat iuxta verbum prius quinta vice puerum suum et epistulam habebat in manu scriptam hoc modo
NEH|6|6|in gentibus auditum est et Gosem dixit quod tu et Iudaei cogitetis rebellare et propterea aedifices murum et levare te velis super eos regem propter quam causam
NEH|6|7|et prophetas posueris qui praedicent de te in Hierusalem dicentes rex in Iudaea est auditurus est rex verba haec idcirco nunc veni ut ineamus consilium pariter
NEH|6|8|et misi ad eos dicens non est factum secundum verba haec quae tu loqueris de corde enim tuo tu conponis haec
NEH|6|9|omnes autem hii terrebant nos cogitantes quod cessarent manus nostrae ab opere et quiesceremus quam ob causam magis confortavi manus meas
NEH|6|10|et ingressus sum domum Samaiae filii Dalaiae filii Metabehel secreto qui ait tractemus nobiscum in domo Dei in medio templi et claudamus portas aedis quia venturi sunt ut interficiant te et nocte venturi sunt ad occidendum te
NEH|6|11|et dixi num quisquam similis mei fugit et quis ut ego ingredietur templum et vivet non ingrediar
NEH|6|12|et intellexi quod Deus non misisset eum sed quasi vaticinans locutus esset ad me et Tobia et Sanaballat conduxissent eum
NEH|6|13|acceperat enim pretium ut territus facerem et peccarem et haberent malum quod exprobrarent mihi
NEH|6|14|memento Domine mei pro Tobia et Sanaballat iuxta opera eorum talia sed et Noadiae prophetae et ceterorum prophetarum qui terrebant me
NEH|6|15|conpletus est autem murus vicesimo quinto die mensis elul quinquaginta duobus diebus
NEH|6|16|factum est ergo cum audissent omnes inimici nostri ut timerent universae gentes quae erant in circuitu nostro et conciderent intra semet ipsos et scirent quod a Deo factum esset opus hoc
NEH|6|17|sed et in diebus illis multae optimatium Iudaeorum epistulae mittebantur ad Tobiam et a Tobia veniebant ad eos
NEH|6|18|multi enim erant in Iudaea habentes iuramentum eius quia gener erat Secheniae filii Orei et Iohanan filius eius acceperat filiam Mosollam filii Barachiae
NEH|6|19|sed et laudabant eum coram me et verba mea nuntiabant ei et Tobias mittebat epistulas ut terreret me
NEH|7|1|postquam autem aedificatus est murus et posui valvas et recensui ianitores et cantores et Levitas
NEH|7|2|praecepi Aneni fratri meo et Ananiae principi domus de Hierusalem ipse enim quasi vir verax et timens Deum plus ceteris videbatur
NEH|7|3|et dixi eis non aperiantur portae Hierusalem usque ad calorem solis cumque adhuc adsisterent clausae portae sunt et oppilatae et posui custodes de habitatoribus Hierusalem singulos per vices suas et unumquemque contra domum suam
NEH|7|4|civitas autem erat lata nimis et grandis et populus parvus in medio eius et non erant domus aedificatae
NEH|7|5|dedit autem Deus in corde meo et congregavi optimates et magistratus et vulgum ut recenserem eos et inveni librum census eorum qui ascenderant primum et inventum est scriptum in eo
NEH|7|6|isti filii provinciae qui ascenderunt de captivitate migrantium quos transtulerat Nabuchodonosor rex Babylonis et reversi sunt in Hierusalem et in Iudaeam unusquisque in civitatem suam
NEH|7|7|qui venerunt cum Zorobabel Hiesuae Neemias Azarias Raamias Naamni Mardocheus Belsar Mespharath Beggoai Naum Baana numerus virorum populi Israhel
NEH|7|8|filii Pharos duo milia centum septuaginta duo
NEH|7|9|filii Saphatiae trecenti septuaginta duo
NEH|7|10|filii Area sescenti quinquaginta duo
NEH|7|11|filii Phaethmoab filiorum Hiesuae et Ioab duo milia octingenti decem et octo
NEH|7|12|filii Helam mille octingenti quinquaginta quattuor
NEH|7|13|filii Zethua octingenti quadraginta quinque
NEH|7|14|filii Zacchai septingenti sexaginta
NEH|7|15|filii Bennui sescenti quadraginta octo
NEH|7|16|filii Bebai sescenti viginti octo
NEH|7|17|filii Azgad duo milia trecenti viginti duo
NEH|7|18|filii Adonicam sescenti sexaginta septem
NEH|7|19|filii Baggoaim duo milia sexaginta septem
NEH|7|20|filii Adin sescenti quinquaginta quinque
NEH|7|21|filii Ater filii Ezechiae nonaginta octo
NEH|7|22|filii Asem trecenti viginti octo
NEH|7|23|filii Besai trecenti viginti quattuor
NEH|7|24|filii Areph centum duodecim
NEH|7|25|filii Gabaon nonaginta quinque
NEH|7|26|viri Bethleem et Netupha centum octoginta octo
NEH|7|27|viri Anathoth centum viginti octo
NEH|7|28|viri Bethamoth quadraginta duo
NEH|7|29|viri Cariathiarim Cephira et Beroth septingenti quadraginta tres
NEH|7|30|viri Rama et Geba sescenti viginti unus
NEH|7|31|viri Machmas centum viginti duo
NEH|7|32|viri Bethel et Hai centum viginti tres
NEH|7|33|viri Nebo alterius quinquaginta duo
NEH|7|34|viri Helam alterius mille ducenti quinquaginta quattuor
NEH|7|35|filii Arem trecenti viginti
NEH|7|36|filii Hiericho trecenti quadraginta quinque
NEH|7|37|filii Lod Adid et Ono septingenti viginti unus
NEH|7|38|filii Senaa tria milia nongenti triginta
NEH|7|39|sacerdotes filii Idaia in domo Iosua nongenti septuaginta tres
NEH|7|40|filii Emmer mille quinquaginta duo
NEH|7|41|filii Phassur mille ducenti quadraginta septem
NEH|7|42|filii Arem mille decem et septem Levitae
NEH|7|43|filii Iosue et Cadmihel filiorum
NEH|7|44|Oduia septuaginta quattuor cantores
NEH|7|45|filii Asaph centum quadraginta octo
NEH|7|46|ianitores filii Sellum filii Ater filii Telmon filii Accub filii Atita filii Sobai centum triginta octo
NEH|7|47|Nathinnei filii Soa filii Asfa filii Tebaoth
NEH|7|48|filii Ceros filii Siaa filii Fado filii Lebana filii Agaba filii Selmon
NEH|7|49|filii Anan filii Geddel filii Gaer
NEH|7|50|filii Raaia filii Rasim filii Necoda
NEH|7|51|filii Gezem filii Aza filii Fasea
NEH|7|52|filii Besai filii Munim filii Nephusim
NEH|7|53|filii Becbuc filii Acupha filii Arur
NEH|7|54|filii Besloth filii Meida filii Arsa
NEH|7|55|filii Bercos filii Sisara filii Thema
NEH|7|56|filii Nesia filii Atipha
NEH|7|57|filii servorum Salomonis filii Sotai filii Sophereth filii Pherida
NEH|7|58|filii Iahala filii Dercon filii Geddel
NEH|7|59|filii Saphatia filii Athil filii Phocereth qui erat ortus ex Sabaim filio Amon
NEH|7|60|omnes Nathinnei et filii servorum Salomonis trecenti nonaginta duo
NEH|7|61|hii sunt autem qui ascenderunt de Thelmella Thelarsa Cherub Addon et Emmer et non potuerunt indicare domum patrum suorum et semen suum utrum ex Israhel essent
NEH|7|62|filii Dalaia filii Tobia filii Necoda sescenti quadraginta duo
NEH|7|63|et de sacerdotibus filii Abia filii Accos filii Berzellai qui accepit de filiabus Berzellai Galaditis uxorem et vocatus est nomine eorum
NEH|7|64|hii quaesierunt scripturam suam in censu et non invenerunt et eiecti sunt de sacerdotio
NEH|7|65|dixitque Athersatha eis ut non manducarent de sanctis sanctorum donec staret sacerdos doctus et eruditus
NEH|7|66|omnis multitudo quasi unus quadraginta duo milia sescenti sexaginta
NEH|7|67|absque servis et ancillis eorum qui erant septem milia trecenti triginta et septem et inter eos cantores et cantrices ducentae quadraginta quinque
NEH|7|68|
NEH|7|69|cameli quadringenti triginta quinque asini sex milia septingenti viginti
NEH|7|70|nonnulli autem de principibus familiarum dederunt in opus Athersatha dedit in thesaurum auri dragmas mille fialas quinquaginta tunicas sacerdotales quingentas triginta
NEH|7|71|et de principibus familiarum dederunt in thesaurum operis auri dragmas viginti milia et argenti minas duo milia ducentas
NEH|7|72|et quod dedit reliquus populus auri dragmas viginti milia et argenti minas duo milia et tunicas sacerdotales sexaginta septem
NEH|7|73|habitaverunt autem sacerdotes et Levitae et ianitores et cantores et reliquum vulgus et Nathinnei et omnis Israhel in civitatibus suis
NEH|8|1|et venerat mensis septimus filii autem Israhel erant in civitatibus suis congregatusque est omnis populus quasi vir unus ad plateam quae est ante portam Aquarum et dixerunt Ezrae scribae ut adferret librum legis Mosi quam praecepit Dominus Israheli
NEH|8|2|adtulit ergo Ezras sacerdos legem coram multitudine virorum et mulierum cunctisque qui poterant intellegere in die prima mensis septimi
NEH|8|3|et legit in eo aperte in platea quae erat ante portam Aquarum de mane usque ad mediam diem in conspectu virorum et mulierum et sapientium et aures omnis populi erant erectae ad librum
NEH|8|4|stetit autem Ezras scriba super gradum ligneum quem fecerat ad loquendum et steterunt iuxta eum Matthathia et Sema et Ania et Uria et Helcia et Maasia ad dextram eius et ad sinistram Phadaia Misahel et Melchia et Asum et Asephdana Zaccharia et Mosollam
NEH|8|5|et aperuit Ezras librum coram omni populo super universum quippe populum eminebat et cum aperuisset eum stetit omnis populus
NEH|8|6|et benedixit Ezras Domino Deo magno et respondit omnis populus amen amen elevans manus suas et incurvati sunt et adoraverunt Deum proni in terram
NEH|8|7|porro Hiesue et Baani et Serebia Iamin Accub Septhai Odia Maasia Celita Azarias Iozabed Anam Phalaia Levitae silentium faciebant in populo ad audiendam legem populus autem stabat in gradu suo
NEH|8|8|et legerunt in libro legis Dei distincte et adposite ad intellegendum et intellexerunt cum legeretur
NEH|8|9|dixit autem Neemias ipse est Athersatha et Ezras sacerdos scriba et Levitae interpretantes universo populo dies sanctificatus est Domino Deo nostro nolite lugere et nolite flere flebat enim omnis populus cum audiret verba legis
NEH|8|10|et dixit eis ite comedite pinguia et bibite mulsum et mittite partes ei qui non praeparavit sibi quia sanctus dies Domini est et nolite contristari gaudium enim Domini est fortitudo nostra
NEH|8|11|Levitae autem silentium faciebant in omni populo dicentes tacete quia dies sanctus est et nolite dolere
NEH|8|12|abiit itaque omnis populus ut comederet et biberet et mitteret partes et faceret laetitiam magnam quia intellexerant verba quae docuerat eos
NEH|8|13|et in die secundo congregati sunt principes familiarum universi populi sacerdotes et Levitae ad Ezram scribam ut interpretaretur eis verba legis
NEH|8|14|et invenerunt scriptum in lege praecepisse Dominum in manu Mosi ut habitent filii Israhel in tabernaculis in die sollemni mense septimo
NEH|8|15|et ut praedicent et divulgent vocem in universis urbibus suis et in Hierusalem dicentes egredimini in montem et adferte frondes olivae et frondes ligni pulcherrimi frondes myrti et ramos palmarum et frondes ligni nemorosi ut fiant tabernacula sicut scriptum est
NEH|8|16|et egressus est populus et adtulerunt feceruntque sibi tabernacula unusquisque in domate suo et in atriis suis et in atriis domus Dei et in platea portae Aquarum et in platea portae Ephraim
NEH|8|17|fecit ergo universa ecclesia eorum qui redierant de captivitate tabernacula et habitaverunt in tabernaculis non enim fecerant a diebus Iosue filii Nun taliter filii Israhel usque ad diem illum et fuit laetitia magna nimis
NEH|8|18|legit autem in libro legis Dei per dies singulos a die primo usque ad diem novissimum et fecerunt sollemnitatem septem diebus et in die octavo collectum iuxta ritum
NEH|9|1|in die autem vicesimo quarto mensis huius convenerunt filii Israhel in ieiunio et in saccis et humus super eos
NEH|9|2|et separatum est semen filiorum Israhel ab omni filio alienigena et steterunt et confitebantur peccata sua et iniquitates patrum suorum
NEH|9|3|et consurrexerunt ad standum et legerunt in volumine legis Domini Dei sui quater in die et quater confitebantur et adorabant Dominum Deum suum
NEH|9|4|surrexit autem super gradum Levitarum Iosue et Bani Cedmihel Sebnia Bani Sarebias Bani Chanani et inclamaverunt voce magna Dominum Deum suum
NEH|9|5|et dixerunt Levitae Iosue et Cedmihel Bonni Asebia Serebia Odoia Sebna Fataia surgite benedicite Domino Deo vestro ab aeterno usque in aeternum et benedicant nomini gloriae tuae excelso in omni benedictione et laude
NEH|9|6|tu ipse Domine solus tu fecisti caelum caelum caelorum et omnem exercitum eorum terram et universa quae in ea sunt maria et omnia quae in eis sunt et tu vivificas omnia haec et exercitus caeli te adorat
NEH|9|7|tu ipse Domine Deus qui elegisti Abram et eduxisti eum de igne Chaldeorum et posuisti nomen eius Abraham
NEH|9|8|et invenisti cor eius fidele coram te et percussisti cum eo foedus ut dares ei terram Chananei Chetthei Amorrei et Ferezei et Iebusei et Gergesei ut dares semini eius et implesti verba tua quoniam iustus es
NEH|9|9|et vidisti adflictionem patrum nostrorum in Aegypto clamoremque eorum audisti super mare Rubrum
NEH|9|10|et dedisti signa et portenta in Pharao et in universis servis eius et in omni populo terrae illius cognovisti enim quia superbe egerant contra eos et fecisti tibi nomen sicut et in hac die
NEH|9|11|et mare divisisti ante eos et transierunt per medium maris in sicca persecutores autem eorum proiecisti in profundum quasi lapidem in aquas validas
NEH|9|12|et in columna nubis ductor eorum fuisti per diem et in columna ignis per noctem ut appareret eis via per quam ingrediebantur
NEH|9|13|ad montem quoque Sinai descendisti et locutus es cum eis de caelo et dedisti eis iudicia recta et legem veritatis caerimonias et praecepta bona
NEH|9|14|et sabbatum sanctificatum tuum ostendisti eis et mandata et caerimonias et legem praecepisti eis in manu Mosi servi tui
NEH|9|15|panem quoque de caelo dedisti eis in fame eorum et aquam de petra eduxisti eis sitientibus et dixisti eis ut ingrederentur et possiderent terram super quam levasti manum tuam ut traderes eis
NEH|9|16|ipsi vero et patres nostri superbe egerunt et induraverunt cervices suas et non audierunt mandata tua
NEH|9|17|et noluerunt audire et non sunt recordati mirabilium tuorum quae feceras eis et induraverunt cervices suas et dederunt caput ut converterentur ad servitutem suam quasi per contentionem tu autem Deus propitius clemens et misericors longanimis et multae miserationis non dereliquisti eos
NEH|9|18|et quidem cum fecissent sibi vitulum conflatilem et dixissent iste est Deus tuus qui eduxit te de Aegypto feceruntque blasphemias magnas
NEH|9|19|tu autem in misericordiis tuis multis non dimisisti eos in deserto columna nubis non recessit ab eis per diem ut duceret eos in via et columna ignis in nocte ut ostenderet eis iter per quod ingrederentur
NEH|9|20|et spiritum tuum bonum dedisti qui doceret eos et manna tuum non prohibuisti ab ore eorum et aquam dedisti eis in siti
NEH|9|21|quadraginta annis pavisti eos in deserto nihilque eis defuit vestimenta eorum non inveteraverunt et pedes eorum non sunt adtriti
NEH|9|22|et dedisti eis regna et populos et partitus es eis sortes et possederunt terram Seon et terram regis Esebon et terram Og regis Basan
NEH|9|23|et filios eorum multiplicasti sicut stellas caeli et adduxisti eos ad terram de qua dixeras patribus eorum ut ingrederentur et possiderent
NEH|9|24|et venerunt filii et possederunt terram et humiliasti coram eis habitatores terrae Chananeos et dedisti eos in manu eorum et reges eorum et populos terrae ut facerent eis sicut placebat illis
NEH|9|25|ceperunt itaque urbes munitas et humum pinguem et possederunt domos plenas cunctis bonis cisternas ab aliis fabricatas vineas et oliveta et ligna pomifera multa et comederunt et saturati sunt et inpinguati sunt et abundavere deliciis in bonitate tua magna
NEH|9|26|provocaverunt autem te ad iracundiam et recesserunt a te et proiecerunt legem tuam post terga sua et prophetas tuos occiderunt qui contestabantur eos ut reverterentur ad te feceruntque blasphemias grandes
NEH|9|27|et dedisti eos in manu hostium suorum et adflixerunt eos et in tempore tribulationis suae clamaverunt ad te et tu de caelo audisti et secundum miserationes tuas multas dedisti eis salvatores qui salvaverunt eos de manu hostium suorum
NEH|9|28|cumque requievissent reversi sunt ut facerent malum in conspectu tuo et dereliquisti eos in manu inimicorum suorum et possederunt eos conversique sunt et clamaverunt ad te tu autem de caelo audisti et liberasti eos in misericordiis tuis multis temporibus
NEH|9|29|et contestatus es eos ut reverterentur ad legem tuam ipsi vero superbe egerunt et non audierunt mandata tua et in iudiciis tuis peccaverunt quae faciet homo et vivet in eis et dederunt umerum recedentem et cervicem suam induraverunt nec audierunt
NEH|9|30|et protraxisti super eos annos multos et contestatus es eos in spiritu tuo per manum prophetarum tuorum et non audierunt et tradidisti eos in manu populorum terrarum
NEH|9|31|in misericordiis autem tuis plurimis non fecisti eos in consumptione nec dereliquisti eos quoniam Deus miserationum et clemens tu es
NEH|9|32|nunc itaque Deus noster Deus magne fortis et terribilis custodiens pactum et misericordiam ne avertas a facie tua omnem laborem qui invenit nos reges nostros principes nostros et sacerdotes nostros prophetas nostros et patres nostros et omnem populum tuum a diebus regis Assur usque in diem hanc
NEH|9|33|et tu iustus in omnibus quae venerunt super nos quia veritatem fecisti nos autem impie egimus
NEH|9|34|reges nostri principes nostri sacerdotes nostri et patres nostri non fecerunt legem tuam et non adtenderunt mandata tua et testimonia tua quae testificatus es in eis
NEH|9|35|et ipsi in regnis suis bonis et in bonitate tua multa quam dederas eis et in terra latissima et pingui quam tradideras in conspectu eorum non servierunt tibi nec reversi sunt ab studiis suis pessimis
NEH|9|36|ecce nos ipsi hodie servi sumus et terram quam dedisti patribus nostris ut comederent panem eius et quae bona sunt eius et nos ipsi servi sumus in ea
NEH|9|37|et fruges eius multiplicantur regibus quos posuisti super nos propter peccata nostra et in corporibus nostris dominantur et in iumentis nostris secundum voluntatem suam et in tribulatione magna sumus
NEH|9|38|super omnibus ergo his nos ipsi percutimus foedus et scribimus et signant principes nostri Levitae nostri et sacerdotes nostri
NEH|10|1|signatores autem fuerunt Neemias Athersatha filius Achelai et Sedecias
NEH|10|2|Saraias Azarias Hieremias
NEH|10|3|Phessur Amaria Melchia
NEH|10|4|Attus Sebenia Melluc
NEH|10|5|Arem Mermuth Obdias
NEH|10|6|Danihel Genton Baruch
NEH|10|7|Mosollam Abia Miamin
NEH|10|8|Mazia Belga Semaia hii sacerdotes
NEH|10|9|porro Levitae Iosue filius Azaniae Bennui de filiis Enadad Cedmihel
NEH|10|10|et fratres eorum Sechenia Odevia Celita Phalaia Anan
NEH|10|11|Micha Roob Asebia
NEH|10|12|Zacchur Serebia Sabania
NEH|10|13|Odia Bani Baninu
NEH|10|14|capita populi Pheros Phaethmoab Helam Zethu Bani
NEH|10|15|Bonni Azgad Bebai
NEH|10|16|Adonia Beggoai Adin
NEH|10|17|Ater Ezechia Azur
NEH|10|18|Odevia Asum Besai
NEH|10|19|Ares Anathoth Nebai
NEH|10|20|Mecphia Mosollam Azir
NEH|10|21|Mesizabel Sadoc Ieddua
NEH|10|22|Felthia Anan Ania
NEH|10|23|Osee Anania Asub
NEH|10|24|Aloes Phaleam Sobec
NEH|10|25|Reum Asebna Madsia
NEH|10|26|et Haia Hanam Anan
NEH|10|27|Melluc Arem Baana
NEH|10|28|et reliqui de populo sacerdotes Levitae ianitores et cantores Nathinnei et omnes qui se separaverunt de populis terrarum ad legem Dei uxores eorum filii eorum et filiae eorum
NEH|10|29|omnis qui poterat sapere spondentes pro fratribus suis optimates eorum et qui veniebant ad pollicendum et iurandum ut ambularent in lege Dei quam dederat in manu Mosi servi Dei ut facerent et custodirent universa mandata Domini Dei nostri et iudicia eius et caerimonias eius
NEH|10|30|et ut non daremus filias nostras populo terrae et filias eorum non acciperemus filiis nostris
NEH|10|31|populi quoque terrae qui inportant venalia et omnia ad usum per diem sabbati ut vendant non accipiemus ab eis in sabbato et in die sanctificata et dimittemus annum septimum et exactionem universae manus
NEH|10|32|et statuemus super nos praecepta ut demus tertiam partem sicli per annum ad opus domus Dei nostri
NEH|10|33|ad panes propositionis et ad sacrificium sempiternum et in holocaustum sempiternum in sabbatis in kalendis in sollemnitatibus et in sanctificatis et pro peccato ut exoretur pro Israhel et in omnem usum domus Dei nostri
NEH|10|34|sortes ergo misimus super oblatione lignorum inter sacerdotes et Levitas et populos ut inferrentur in domum Dei nostri per domos patrum nostrorum per tempora a temporibus anni usque ad annum ut arderent super altare Domini Dei nostri sicut scriptum est in lege Mosi
NEH|10|35|et ut adferremus primogenita terrae nostrae et primitiva universi fructus omnis ligni ab anno in annum in domo Domini
NEH|10|36|et primitiva filiorum nostrorum et pecorum nostrorum sicut scriptum est in lege et primitiva boum nostrorum et ovium nostrarum ut offerrentur in domo Dei nostri sacerdotibus qui ministrant in domo Dei nostri
NEH|10|37|et primitias ciborum nostrorum et libaminum nostrorum et poma omnis ligni vindemiae quoque et olei adferemus sacerdotibus ad gazofilacium Dei nostri et decimam partem terrae nostrae Levitis ipsi Levitae decimas accipient ex omnibus civitatibus operum nostrorum
NEH|10|38|erit autem sacerdos filius Aaron cum Levitis in decimis Levitarum et Levitae offerent decimam partem decimae suae in domum Dei nostri ad gazofilacium in domo thesauri
NEH|10|39|ad gazofilacium enim deportabunt filii Israhel et filii Levi primitias frumenti vini et olei et ibi erunt vasa sanctificata et sacerdotes et cantores et ianitores et ministri et non dimittemus domum Dei nostri
NEH|11|1|habitaverunt autem principes populi in Hierusalem reliqua vero plebs misit sortem ut tollerent unam partem de decem qui habitaturi essent in Hierusalem in civitate sancta novem vero partes in civitatibus
NEH|11|2|benedixit autem populus omnibus viris qui se sponte obtulerunt ut habitarent in Hierusalem
NEH|11|3|hii sunt itaque principes provinciae qui habitaverunt in Hierusalem et in civitatibus Iuda habitavit unusquisque in possessione sua in urbibus suis Israhel sacerdotes Levitae Nathinnei et filii servorum Salomonis
NEH|11|4|et in Hierusalem habitaverunt de filiis Iuda et de filiis Beniamin de filiis Iuda Athaias filius Aziam filii Zacchariae filii Amariae filii Saphatia filii Malelehel de filiis Phares
NEH|11|5|Imaasia filius Baruch filius Coloza filius Azia filius Adaia filius Ioiarib filius Zacchariae filius Silonites
NEH|11|6|omnes filii Phares qui habitaverunt in Hierusalem quadringenti sexaginta octo viri fortes
NEH|11|7|hii sunt autem filii Beniamin Sellum filius Mosollam filius Ioed filius Phadaia filius Colaia filius Masia filius Ethehel filius Isaia
NEH|11|8|et post eum Gabbai Sellai nongenti viginti octo
NEH|11|9|et Iohel filius Zechri praepositus eorum et Iuda filius Sennua super civitatem secundus
NEH|11|10|et de sacerdotibus Idaia filius Ioarib Iachin
NEH|11|11|Saraia filius Elcia filius Mesollam filius Sadoc filius Meraioth filius Ahitub princeps domus Dei
NEH|11|12|et fratres eorum facientes opera templi octingenti viginti duo et Adaia filius Ieroam filius Felelia filius Amsi filius Zacchariae filius Phessur filius Melchiae
NEH|11|13|et fratres eius principes patrum ducenti quadraginta duo et Amassai filius Azrihel filius Aazi filius Mosollamoth filius Emmer
NEH|11|14|et fratres eorum potentes nimis centum viginti octo et praepositus eorum Zabdihel filius potentium
NEH|11|15|et de Levitis Sebenia filius Asob filius Azaricam filius Asabia filius Boni
NEH|11|16|et Sabathai et Iozabed super opera quae erant forinsecus in domo Dei a principibus Levitarum
NEH|11|17|et Mathania filius Micha filius Zebdaei filius Asaph princeps ad laudandum et confitendum in oratione et Becbecia secundus de fratribus eius et Abda filius Sammua filius Galal filius Idithun
NEH|11|18|omnes Levitae in civitate sancta ducenti octoginta quattuor
NEH|11|19|et ianitores Accob Telmon et fratres eorum qui custodiebant ostia centum septuaginta duo
NEH|11|20|et reliqui ex Israhel sacerdotes et Levitae in universis civitatibus Iuda unusquisque in possessione sua
NEH|11|21|et Nathinnei qui habitabant in Ofel et Siaha et Gaspha de Nathinneis
NEH|11|22|et episcopus Levitarum in Hierusalem Azzi filius Bani filius Asabiae filius Matthaniae filius Michae de filiis Asaph cantores in ministerio domus Dei
NEH|11|23|praeceptum quippe regis super eos erat et ordo in cantoribus per dies singulos
NEH|11|24|et Fataia filius Mesezebel de filiis Zera filii Iuda in manu regis iuxta omne verbum populi
NEH|11|25|et in domibus per omnes regiones eorum de filiis Iuda habitaverunt in Cariatharbe et in filiabus eius et in Dibon et in filiabus eius et in Capsel et in viculis eius
NEH|11|26|et in Iesue et in Molada et in Bethfaleth
NEH|11|27|et in Asersual et in Bersabee et in filiabus eius
NEH|11|28|et in Siceleg et in Mochona et in filiabus eius
NEH|11|29|et in Ainremmon et in Sara et in Irimuth
NEH|11|30|Zanoa Odollam et villis earum Lachis et regionibus eius Azeca et filiabus eius et manserunt in Bersabee usque ad vallem Ennom
NEH|11|31|filii autem Beniamin a Geba Mechmas et Aia et Bethel et filiabus eius
NEH|11|32|Anathoth Nob Anania
NEH|11|33|Asor Rama Getthaim
NEH|11|34|Adid Seboim Neballa Loth
NEH|11|35|et Ono valle Artificum
NEH|11|36|et de Levitis partitiones Iuda et Beniamin
NEH|12|1|hii autem sacerdotes et Levitae qui ascenderunt cum Zorobabel filio Salathihel et Iosue Saraia Hieremias Ezra
NEH|12|2|Amaria Melluch Attus
NEH|12|3|Sechenia Reum Meremuth
NEH|12|4|Addo Genthon Abia
NEH|12|5|Miamin Madia Belga
NEH|12|6|Semaia et Ioarib Idaia Sellum Amoc Elceia
NEH|12|7|Idaia isti principes sacerdotum et fratres eorum in diebus Iosue
NEH|12|8|porro Levitae Iesua Bennui Cedmihel Sarabia Iuda Mathanias super hymnos ipsi et fratres eorum
NEH|12|9|et Becbecia atque et Hanni fratres eorum unusquisque in officio suo
NEH|12|10|Hiesue autem genuit Ioachim et Ioachim genuit Eliasib et Eliasib genuit Ioiada
NEH|12|11|et Ioiada genuit Ionathan et Ionathan genuit Ieddoa
NEH|12|12|in diebus autem Ioachim erant sacerdotes principes familiarum Saraiae Amaria Hieremiae Anania
NEH|12|13|Ezrae Mosollam Amariae Iohanan
NEH|12|14|Milico Ionathan Sebeniae Ioseph
NEH|12|15|Arem Edna Maraioth Elci
NEH|12|16|Addaiae Zaccharia Genthon Mosollam
NEH|12|17|Abiae Zecheri Miamin et Moadiae Felti
NEH|12|18|Belgae Sammua Semaiae Ionathan
NEH|12|19|Ioiarib Matthanai Iadaiae Azzi
NEH|12|20|Sellaiae Celai Amoc Eber
NEH|12|21|Elciae Asebia Idaiae Nathanahel
NEH|12|22|Levitae in diebus Eliasib et Ioiada et Ionan et Ieddoa scripti principes familiarum et sacerdotes in regno Darii Persae
NEH|12|23|filii Levi principes familiarum scripti in libro verborum dierum et usque ad dies Ionathan filii Eliasib
NEH|12|24|et principes Levitarum Asebia Serebia et Iesue filius Cedmihel et fratres eorum per vices suas ut laudarent et confiterentur iuxta praeceptum David viri Dei et observarent aeque per ordinem
NEH|12|25|Matthania et Becbecia Obedia Mosollam Thelmon Accub custodes portarum et vestibulorum ante portas
NEH|12|26|hii in diebus Ioachim filii Iesue filii Iosedech et in diebus Neemiae ducis et Ezrae sacerdotis scribaeque
NEH|12|27|in dedicatione autem muri Hierusalem requisierunt Levitas de omnibus locis suis ut adducerent eos in Hierusalem et facerent dedicationem et laetitiam in actione gratiarum et in cantico in cymbalis psalteriis et citharis
NEH|12|28|congregati sunt ergo filii cantorum et de campestribus circa Hierusalem et de villis Netuphati
NEH|12|29|et de domo Galgal et de regionibus Geba et Azmaveth quoniam villas aedificaverunt sibi cantores in circuitu Hierusalem
NEH|12|30|et mundati sunt sacerdotes et Levitae et mundaverunt populum et portas et murum
NEH|12|31|ascendere autem feci principes Iuda super murum et statui duos choros laudantium magnos et ierunt ad dexteram super murum ad portam Sterquilinii
NEH|12|32|et ivit post eos Osaias et media pars principum Iuda
NEH|12|33|et Azarias Ezras et Mosollam Iuda et Beniamin et Semeia et Hieremia
NEH|12|34|et de filiis sacerdotum in tubis Zaccharias filius Ionathan filius Semeiae filius Mathaniae filius Michaiae filius Zecchur filius Asaph
NEH|12|35|et fratres eius Semeia et Azarel Malalai Galalai Maai Nathanel et Iuda et Anani in vasis cantici David viri Dei et Ezras scriba ante eos in porta Fontis
NEH|12|36|et contra eos ascenderunt in gradibus civitatis David in ascensu muri super domum David et usque ad portam Aquarum ad orientem
NEH|12|37|et chorus secundus gratias referentium ibat ex adverso et ego post eum et media pars populi super murum et super turrem Furnorum et usque ad murum latissimum
NEH|12|38|et super portam Ephraim et super portam Antiquam et super portam Piscium et turrem Ananehel et turrem Ema et usque ad portam Gregis et steterunt in porta Custodiae
NEH|12|39|steteruntque duo chori laudantium in domo Dei et ego et dimidia pars magistratuum mecum
NEH|12|40|et sacerdotes Eliachim Maasia Miniamin Michea Elioenai Zaccharia Anania in tubis
NEH|12|41|et Maasia et Semea et Eleazar et Azi et Iohanan et Melchia et Elam et Ezer et clare cecinerunt cantores et Iezraia praepositus
NEH|12|42|et immolaverunt in die illa victimas magnas et laetati sunt Deus enim laetificaverat eos laetitia magna sed et uxores eorum et liberi gavisi sunt et audita est laetitia Hierusalem procul
NEH|12|43|recensuerunt quoque in die illa viros super gazofilacia thesauri ad libamina et ad primitias et ad decimas ut introferrent per eos principes civitatis in decore gratiarum actionis sacerdotes et Levitas quia laetatus est Iuda in sacerdotibus et Levitis adstantibus
NEH|12|44|et custodierunt observationem Dei sui et observationem expiationis et cantores et ianitores iuxta praeceptum David et Salomonis filii eius
NEH|12|45|quia in diebus David et Asaph ab exordio erant principes constituti cantorum in carmine laudantium et confitentium Deo
NEH|12|46|et omnis Israhel in diebus Zorobabel et in diebus Neemiae dabat partes cantoribus et ianitoribus per dies singulos et sanctificabant Levitas et Levitae sanctificabant filios Aaron
NEH|13|1|in die autem illo lectum est in volumine Mosi audiente populo et inventum est scriptum in eo quod non debeat introire Ammanites et Moabites in ecclesiam Dei usque in aeternum
NEH|13|2|eo quod non occurrerint filiis Israhel cum pane et aqua et conduxerint adversum eum Balaam ad maledicendum ei et convertit Deus noster maledictionem in benedictionem
NEH|13|3|factum est autem cum audissent legem separaverunt omnem alienigenam ab Israhel
NEH|13|4|et super hoc erat Eliasib sacerdos qui fuerat positus in gazofilacio domus Dei nostri et proximus Tobiae
NEH|13|5|fecit ergo sibi gazofilacium grande et ibi erant ante eum reponentes munera et tus et vasa et decimam frumenti et vini et olei partes Levitarum et cantorum et ianitorum et primitias sacerdotales
NEH|13|6|in omnibus autem his non fui in Hierusalem quia in anno tricesimo secundo Artarxersis regis Babylonis veni ad regem et in fine dierum rogavi regem
NEH|13|7|et veni in Hierusalem et intellexi malum quod fecerat Eliasib Tobiae ut faceret ei thesaurum in vestibulis domus Dei
NEH|13|8|et malum mihi visum est valde et proieci vasa domus Tobiae foras de gazofilacio
NEH|13|9|praecepique et mundaverunt gazofilacia et rettuli ibi vasa domus Dei sacrificium et tus
NEH|13|10|et cognovi quoniam partes Levitarum non fuissent datae et fugisset unusquisque in regionem suam de Levitis et de cantoribus et de his qui ministrabant
NEH|13|11|et egi causam adversus magistratus et dixi quare dereliquimus domum Dei et congregavi eos et feci stare in stationibus suis
NEH|13|12|et omnis Iuda adportabat decimam frumenti et vini et olei in horrea
NEH|13|13|et constituimus super horrea Selemiam sacerdotem et Sadoc scribam et Phadaiam de Levitis et iuxta eos Anan filium Zacchur filium Matthaniae quoniam fideles conprobati sunt et ipsis creditae sunt partes fratrum suorum
NEH|13|14|memento mei Deus meus pro hoc et ne deleas miserationes meas quas feci in domo Dei mei et in caerimoniis eius
NEH|13|15|in diebus illis vidi in Iuda calcabant torcularia in sabbato portantes acervos et onerantes super asinos vinum et uvas et ficus et omne onus et inferentes Hierusalem in die sabbati et contestatus sum ut in die qua vendere liceret venderent
NEH|13|16|et Tyrii habitaverunt in ea inferentes pisces et omnia venalia et vendebant in sabbatis filiis Iuda et in Hierusalem
NEH|13|17|et obiurgavi optimates Iuda et dixi eis quae est res haec mala quam vos facitis et profanatis diem sabbati
NEH|13|18|numquid non haec fecerunt patres nostri et adduxit Deus noster super nos omne malum hoc et super civitatem hanc et vos additis iracundiam super Israhel violando sabbatum
NEH|13|19|factum est itaque cum quievissent portae Hierusalem die sabbati dixi et cluserunt ianuas et praecepi ut non aperirent eas usque post sabbatum et de pueris meis constitui super portas ut nullus inferret onus in die sabbati
NEH|13|20|et manserunt negotiatores et vendentes universa venalia foris Hierusalem semel et bis
NEH|13|21|et contestatus sum eos et dixi eis quare manetis ex adverso muri si secundo hoc feceritis manum mittam in vos itaque ex tempore illo non venerunt in sabbato
NEH|13|22|dixi quoque Levitis ut mundarentur et venirent ad custodiendas portas et sanctificandum diem sabbati et pro hoc ergo memento mei Deus meus et parce mihi secundum multitudinem miserationum tuarum
NEH|13|23|sed et in diebus illis vidi Iudaeos ducentes uxores azotias ammanitidas et moabitidas
NEH|13|24|et filii eorum ex media parte loquebantur azotice et nesciebant loqui iudaice et loquebantur iuxta linguam populi et populi
NEH|13|25|et obiurgavi eos et maledixi et cecidi ex ipsis viros et decalvavi eos et adiuravi in Deo ut non darent filias suas filiis eorum et non acciperent de filiabus eorum filiis suis et sibimet ipsis dicens
NEH|13|26|numquid non in huiuscemodi re peccavit Salomon rex Israhel et certe in gentibus multis non erat rex similis ei et dilectus Deo suo erat et posuit eum Deus regem super omnem Israhel et ipsum ergo ad peccatum duxerunt mulieres alienigenae
NEH|13|27|numquid et nos inoboedientes faciemus omne malum grande hoc ut praevaricemur in Deo nostro et ducamus uxores peregrinas
NEH|13|28|de filiis autem Ioiada filii Eliasib sacerdotis magni gener erat Sanaballat Horonitis quem fugavi a me
NEH|13|29|recordare Domine Deus meus adversum eos qui polluunt sacerdotium iusque sacerdotale et leviticum
NEH|13|30|igitur mundavi eos ab omnibus alienigenis et constitui ordines sacerdotum et Levitarum unumquemque in ministerio suo
NEH|13|31|et in oblatione lignorum in temporibus constitutis et in primitiis memento mei Deus meus in bonum
ESTH|1|1|in diebus Asueri qui regnavit ab India usque Aethiopiam super centum viginti septem provincias
ESTH|1|2|quando sedit in solio regni sui Susa civitas regni eius exordium fuit
ESTH|1|3|tertio igitur anno imperii sui fecit grande convivium cunctis principibus et pueris suis fortissimis Persarum et Medorum inclitis et praefectis provinciarum coram se
ESTH|1|4|ut ostenderet divitias gloriae regni sui ac magnitudinem atque iactantiam potentiae suae multo tempore centum videlicet et octoginta diebus
ESTH|1|5|cumque implerentur dies convivii invitavit omnem populum qui inventus est Susis a maximo usque ad minimum et septem diebus iussit convivium praeparari in vestibulo horti et nemoris quod regio cultu et manu consitum erat
ESTH|1|6|et pendebant ex omni parte tentoria aerii coloris et carpasini et hyacinthini sustentata funibus byssinis atque purpureis qui eburneis circulis inserti erant et columnis marmoreis fulciebantur lectuli quoque aurei et argentei super pavimentum zmaragdino et pario stratum lapide dispositi erant quod mira varietate pictura decorabat
ESTH|1|7|bibebant autem qui invitati erant aureis poculis et aliis atque aliis vasis cibi inferebantur vinum quoque ut magnificentia regia dignum erat abundans et praecipuum ponebatur
ESTH|1|8|nec erat qui nolentes cogeret ad bibendum sed sic rex statuerat praeponens mensis singulos de principibus suis ut sumeret unusquisque quod vellet
ESTH|1|9|Vasthi quoque regina fecit convivium feminarum in palatio ubi rex Asuerus manere consueverat
ESTH|1|10|itaque die septimo cum rex esset hilarior et post nimiam potionem incaluisset mero praecepit Mauman et Bazatha et Arbona et Bagatha et Abgatha et Zarath et Charchas septem eunuchis qui in conspectu eius ministrabant
ESTH|1|11|ut introducerent reginam Vasthi coram rege posito super caput eius diademate et ostenderet cunctis populis et principibus illius pulchritudinem erat enim pulchra valde
ESTH|1|12|quae rennuit et ad regis imperium quod per eunuchos mandaverat venire contempsit unde iratus rex et nimio furore succensus
ESTH|1|13|interrogavit sapientes qui ex more regio semper ei aderant et illorum faciebat cuncta consilio scientium leges ac iura maiorum
ESTH|1|14|erant autem primi et proximi Charsena et Sethar et Admatha et Tharsis et Mares et Marsana et Mamucha septem duces Persarum atque Medorum qui videbant faciem regis et primi post eum residere soliti erant
ESTH|1|15|cui sententiae Vasthi regina subiaceret quae Asueri regis imperium quod per eunuchos mandaverat facere noluisset
ESTH|1|16|responditque Mamuchan audiente rege atque principibus non solum regem laesit regina Vasthi sed omnes principes et populos qui sunt in cunctis provinciis regis Asueri
ESTH|1|17|egredietur enim sermo reginae ad omnes mulieres ut contemnant viros suos et dicant rex Asuerus iussit ut regina Vasthi intraret ad eum et illa noluit
ESTH|1|18|atque hoc exemplo omnes principum coniuges Persarum atque Medorum parvipendent imperia maritorum unde regis iusta est indignatio
ESTH|1|19|et si tibi placet egrediatur edictum a facie tua et scribatur iuxta legem Persarum atque Medorum quam praeteriri inlicitum est ut nequaquam ultra Vasthi ingrediatur ad regem sed regnum illius altera quae melior illa est accipiat
ESTH|1|20|et hoc in omne quod latissimum est provinciarum tuarum divulgetur imperium et cunctae uxores tam maiorum quam minorum deferant maritis suis
ESTH|1|21|placuit consilium eius regi et principibus fecitque rex iuxta consultum Mamuchan
ESTH|1|22|et misit epistulas ad universas provincias regni sui ut quaeque gens audire et legere poterat diversis linguis et litteris esse viros principes ac maiores in domibus suis et hoc per cunctos populos divulgari
ESTH|2|1|his itaque gestis postquam regis Asueri deferbuerat indignatio recordatus est Vasthi et quae fecisset vel quae passa esset
ESTH|2|2|dixeruntque pueri regis ac ministri eius quaerantur regi puellae virgines ac speciosae
ESTH|2|3|et mittantur qui considerent per universas provincias puellas speciosas et virgines et adducant eas ad civitatem Susan et tradant in domum feminarum sub manu Aegaei eunuchi qui est praepositus et custos mulierum regiarum et accipiant mundum muliebrem et cetera ad usus necessaria
ESTH|2|4|et quaecumque inter omnes oculis regis placuerit ipsa regnet pro Vasthi placuit sermo regi et ita ut suggesserant iussit fieri
ESTH|2|5|erat vir iudaeus in Susis civitate vocabulo Mardocheus filius Iair filii Semei filii Cis de stirpe Iemini
ESTH|2|6|qui translatus fuerat de Hierusalem eo tempore quo Iechoniam regem Iuda Nabuchodonosor rex Babylonis transtulerat
ESTH|2|7|qui fuit nutricius filiae fratris sui Edessae quae altero nomine Hester vocabatur et utrumque parentem amiserat pulchra nimis et decora facie mortuisque patre eius ac matre Mardocheus sibi eam adoptavit in filiam
ESTH|2|8|cumque percrebuisset regis imperium et iuxta mandata illius multae virgines pulchrae adducerentur Susan et Aegaeo traderentur eunucho Hester quoque inter ceteras puellas ei tradita est ut servaretur in numero feminarum
ESTH|2|9|quae placuit ei et invenit gratiam in conspectu illius ut adceleraret mundum muliebrem et traderet ei partes suas et septem puellas speciosissimas de domo regis et tam ipsam quam pedisequas eius ornaret atque excoleret
ESTH|2|10|quae noluit indicare ei populum et patriam suam Mardocheus enim praeceperat ut de hac re omnino reticeret
ESTH|2|11|qui deambulabat cotidie ante vestibulum domus in qua electae virgines servabantur curam agens salutis Hester et scire volens quid ei accideret
ESTH|2|12|cum autem venisset tempus singularum per ordinem puellarum ut intrarent ad regem expletis omnibus quae ad cultum muliebrem pertinebant mensis duodecimus vertebatur ita dumtaxat ut sex menses oleo unguerentur myrtino et aliis sex quibusdam pigmentis et aromatibus uterentur
ESTH|2|13|ingredientesque ad regem quicquid postulassent ad ornatum pertinens accipiebant et ut eis placuerat conpositae de triclinio feminarum ad regis cubiculum transiebant
ESTH|2|14|et quae intraverat vespere egrediebatur mane atque inde in secundas aedes deducebatur quae sub manu Sasagazi eunuchi erant qui concubinis regis praesidebat nec habebat potestatem ad regem ultra redeundi nisi voluisset rex et eam venire iussisset ex nomine
ESTH|2|15|evoluto autem tempore per ordinem instabat dies quo Hester filia Abiahil fratris Mardochei quam sibi adoptaverat in filiam intrare deberet ad regem quae non quaesivit muliebrem cultum sed quaecumque voluit Aegaeus eunuchus custos virginum haec ei ad ornatum dedit erat enim formonsa valde et incredibili pulchritudine omnium oculis gratiosa et amabilis videbatur
ESTH|2|16|ducta est itaque ad cubiculum regis Asueri mense decimo qui vocatur tebeth septimo anno regni eius
ESTH|2|17|et amavit eam rex plus quam omnes mulieres habuitque gratiam et misericordiam coram eo super omnes mulieres et posuit diadema regni in capite eius fecitque eam regnare in loco Vasthi
ESTH|2|18|et iussit convivium praeparari permagnificum cunctis principibus et servis suis pro coniunctione et nuptiis Hester et dedit requiem in universis provinciis ac dona largitus est iuxta magnificentiam principalem
ESTH|2|19|cumque et secundo quaererentur virgines et congregarentur Mardocheus manebat ad regis ianuam
ESTH|2|20|necdumque prodiderat Hester patriam et populum suum iuxta mandatum eius quicquid enim ille praecipiebat observabat Hester et ita cuncta faciebat ut eo tempore solita erat quo eam parvulam nutriebat
ESTH|2|21|eo igitur tempore quo Mardocheus ad regis ianuam morabatur irati sunt Bagathan et Thares duo eunuchi regis qui ianitores erant et in primo palatii limine praesidebant volueruntque insurgere in regem et occidere eum
ESTH|2|22|quod Mardocheum non latuit statimque nuntiavit reginae Hester et illa regi ex nomine Mardochei qui ad se rem detulerat
ESTH|2|23|quaesitum est et inventum et adpensus uterque eorum in patibulo mandatumque historiis et annalibus traditum coram rege
ESTH|3|1|post haec rex Asuerus exaltavit Aman filium Amadathi qui erat de stirpe Agag et posuit solium eius super omnes principes quos habebat
ESTH|3|2|cunctique servi regis qui in foribus palatii versabantur flectebant genu et adorabant Aman sic enim eis praeceperat imperator solus Mardocheus non flectebat genu neque adorabat eum
ESTH|3|3|cui dixerunt regis pueri qui ad fores palatii praesidebant cur praeter ceteros non observas mandata regis
ESTH|3|4|cumque hoc crebrius dicerent et ille nollet audire nuntiaverunt Aman scire cupientes utrum perseveraret in sententia dixerat enim eis se esse Iudaeum
ESTH|3|5|quod cum audisset Aman et experimento probasset quod Mardocheus non sibi flecteret genu nec se adoraret iratus est valde
ESTH|3|6|et pro nihilo duxit in unum Mardocheum mittere manus suas audierat enim quod esset gentis iudaeae magisque voluit omnem Iudaeorum qui erant in regno Asueri perdere nationem
ESTH|3|7|mense primo cuius vocabulum est nisan anno duodecimo regni Asueri missa est sors in urnam quae hebraice dicitur phur coram Aman quo die et quo mense gens Iudaeorum deberet interfici et exivit mensis duodecimus qui vocatur adar
ESTH|3|8|dixitque Aman regi Asuero est populus per omnes provincias regni tui dispersus et a se mutuo separatus novis utens legibus et caerimoniis insuper et regis scita contemnens et optime nosti quod non expediat regno tuo ut insolescat per licentiam
ESTH|3|9|si tibi placet decerne ut pereat et decem milia talentorum adpendam arcariis gazae tuae
ESTH|3|10|tulit ergo rex anulum quo utebatur de manu sua et dedit eum Aman filio Amadathi de progenie Agag hosti Iudaeorum
ESTH|3|11|dixitque ad eum argentum quod polliceris tuum sit de populo age quod tibi placet
ESTH|3|12|vocatique sunt scribae regis mense primo nisan tertiadecima die eius et scriptum est ut iusserat Aman ad omnes satrapas regis et iudices provinciarum diversarumque gentium ut quaeque gens legere poterat et audire pro varietate linguarum ex nomine regis Asueri et litterae ipsius signatae anulo
ESTH|3|13|missae sunt per cursores regis ad universas provincias ut occiderent atque delerent omnes Iudaeos a puero usque ad senem parvulos et mulieres uno die hoc est tertiodecimo mensis duodecimi qui vocatur adar et bona eorum diriperent
ESTH|3|14|summa autem epistularum haec fuit ut omnes provinciae scirent et pararent se ad praedictam diem
ESTH|3|15|festinabant cursores qui missi erant explere regis imperium statimque in Susis pependit edictum rege et Aman celebrante convivium et cunctis qui in urbe erant flentibus
ESTH|4|1|quae cum audisset Mardocheus scidit vestimenta sua et indutus est sacco spargens cinerem capiti et in platea mediae civitatis voce magna clamabat ostendens amaritudinem animi sui
ESTH|4|2|et hoc heiulatu usque ad fores palatii gradiens non enim erat licitum indutum sacco aulam regis intrare
ESTH|4|3|in omnibus quoque provinciis oppidis ac locis ad quae crudele regis dogma pervenerat planctus ingens erat apud Iudaeos ieiunium ululatus et fletus sacco et cinere multis pro strato utentibus
ESTH|4|4|ingressae sunt autem puellae Hester et eunuchi nuntiaveruntque ei quod audiens consternata est et misit vestem ut ablato sacco induerent eum quam accipere noluit
ESTH|4|5|accitoque Athac eunucho quem rex ministrum ei dederat praecepit ut iret ad Mardocheum et disceret ab eo cur hoc faceret
ESTH|4|6|egressusque Athac ivit ad Mardocheum stantem in platea civitatis ante ostium palatii
ESTH|4|7|qui indicavit ei omnia quae acciderant quomodo Aman promisisset ut in thesauros regis pro Iudaeorum nece inferret argentum
ESTH|4|8|exemplarque edicti quod pendebat in Susis dedit ei ut reginae ostenderet et moneret eam ut intraret ad regem et deprecaretur eum pro populo suo
ESTH|4|9|regressus Athac nuntiavit Hester omnia quae Mardocheus dixerat
ESTH|4|10|quae respondit ei et iussit ut diceret Mardocheo
ESTH|4|11|omnes servi regis et cunctae quae sub dicione eius sunt norunt provinciae quod sive vir sive mulier invocatus interius atrium regis intraverit absque ulla cunctatione statim interficiatur nisi forte rex auream virgam ad eum tetenderit pro signo clementiae atque ita possit vivere ego igitur quomodo ad regem intrare potero quae triginta iam diebus non sum vocata ad eum
ESTH|4|12|quod cum audisset Mardocheus
ESTH|4|13|rursum mandavit Hester dicens ne putes quod animam tuam tantum liberes quia in domo regis es prae cunctis Iudaeis
ESTH|4|14|si enim nunc silueris per aliam occasionem liberabuntur Iudaei et tu et domus patris tui peribitis et quis novit utrum idcirco ad regnum veneris ut in tali tempore parareris
ESTH|4|15|rursumque Hester haec Mardocheo verba mandavit
ESTH|4|16|vade et congrega omnes Iudaeos quos in Susis reppereris et orate pro me non comedatis et non bibatis tribus diebus ac noctibus et ego cum ancillulis meis similiter ieiunabo et tunc ingrediar ad regem contra legem faciens invocata tradensque me morti et periculo
ESTH|4|17|ivit itaque Mardocheus et fecit omnia quae ei Hester praeceperat
ESTH|5|1|die autem tertio induta est Hester regalibus vestimentis et stetit in atrio domus regiae quod erat interius contra basilicam regis at ille sedebat super solium in consistorio palatii contra ostium domus
ESTH|5|2|cumque vidisset Hester reginam stantem placuit oculis eius et extendit contra eam virgam auream quam tenebat manu quae accedens osculata est summitatem virgae eius
ESTH|5|3|dixitque ad eam rex quid vis Hester regina quae est petitio tua etiam si dimidiam regni partem petieris dabitur tibi
ESTH|5|4|at illa respondit si regi placet obsecro ut venias ad me hodie et Aman tecum ad convivium quod paravi
ESTH|5|5|statimque rex vocate inquit cito Aman ut Hester oboediat voluntati venerunt itaque rex et Aman ad convivium quod eis regina paraverat
ESTH|5|6|dixitque ei rex postquam vinum biberat abundanter quid petis ut detur tibi et pro qua re postulas etiam si dimidiam partem regni mei petieris inpetrabis
ESTH|5|7|cui respondit Hester petitio mea et preces istae sunt
ESTH|5|8|si inveni gratiam in conspectu regis et si regi placet ut det mihi quod postulo et meam impleat petitionem veniat rex et Aman ad convivium quod paravi eis et cras regi aperiam voluntatem meam
ESTH|5|9|egressus est itaque illo die Aman laetus et alacer cumque vidisset Mardocheum sedentem ante fores palatii et non solum non adsurrexisse sibi sed nec motum quidem de loco sessionis suae indignatus est valde
ESTH|5|10|et dissimulata ira reversus in domum suam convocavit ad se amicos et Zares uxorem suam
ESTH|5|11|et exposuit illis magnitudinem divitiarum suarum filiorumque turbam et quanta eum gloria super omnes principes et servos suos rex elevasset
ESTH|5|12|et post haec ait regina quoque Hester nullum alium vocavit cum rege ad convivium praeter me apud quam etiam cras cum rege pransurus sum
ESTH|5|13|et cum haec omnia habeam nihil me habere puto quamdiu videro Mardocheum Iudaeum sedentem ante fores regias
ESTH|5|14|responderuntque ei Zares uxor eius et ceteri amici iube parari excelsam trabem habentem altitudinem quinquaginta cubitos et dic mane regi ut adpendatur super eam Mardocheus et sic ibis cum rege laetus ad convivium placuit ei consilium et iussit excelsam parari crucem
ESTH|6|1|noctem illam rex duxit insomnem iussitque adferri sibi historias et annales priorum temporum qui cum illo praesente legerentur
ESTH|6|2|ventum est ad eum locum ubi scriptum erat quomodo nuntiasset Mardocheus insidias Bagathan et Thares eunuchorum regem Asuerum iugulare cupientium
ESTH|6|3|quod cum rex audisset ait quid pro hac fide honoris ac praemii Mardocheus consecutus est dixeruntque ei servi illius ac ministri nihil omnino mercedis accepit
ESTH|6|4|statimque rex quis est inquit in atrio Aman quippe interius atrium domus regiae intraverat ut suggereret regi et iuberet Mardocheum adfigi patibulo quod ei fuerat praeparatum
ESTH|6|5|responderunt pueri Aman stat in atrio dixitque rex ingrediatur
ESTH|6|6|cumque esset ingressus ait illi quid debet fieri viro quem rex honorare desiderat cogitans Aman in corde suo et reputans quod nullum alium rex nisi se vellet honorare
ESTH|6|7|respondit homo quem rex honorare cupit
ESTH|6|8|debet indui vestibus regiis et inponi super equum qui de sella regis est et accipere regium diadema super caput suum
ESTH|6|9|et primus de regis principibus ac tyrannis teneat equum eius et per plateam civitatis incedens clamet ac dicat sic honorabitur quemcumque rex voluerit honorare
ESTH|6|10|dixitque ei rex festina et sumpta stola et equo fac ita ut locutus es Mardocheo Iudaeo qui sedet ante fores palatii cave ne quicquam de his quae locutus es praetermittas
ESTH|6|11|tulit itaque Aman stolam et equum indutumque Mardocheum in platea civitatis et inpositum equo praecedebat atque clamabat hoc honore condignus est quemcumque rex voluerit honorare
ESTH|6|12|reversus est Mardocheus ad ianuam palatii et Aman festinavit ire in domum suam lugens et operto capite
ESTH|6|13|narravitque Zares uxori suae et amicis omnia quae evenissent sibi cui responderunt sapientes quos habebat in consilio et uxor eius si de semine Iudaeorum est Mardocheus ante quem cadere coepisti non poteris ei resistere sed cades in conspectu eius
ESTH|6|14|adhuc illis loquentibus venerunt eunuchi regis et cito eum ad convivium quod regina paraverat pergere conpulerunt
ESTH|7|1|intravit itaque rex et Aman ut biberent cum regina
ESTH|7|2|dixitque ei rex etiam in secundo die postquam vino incaluerat quae est petitio tua Hester ut detur tibi et quid vis fieri etiam si dimidiam regni mei partem petieris inpetrabis
ESTH|7|3|ad quem illa respondit si inveni gratiam in oculis tuis o rex et si tibi placet dona mihi animam meam pro qua rogo et populum meum pro quo obsecro
ESTH|7|4|traditi enim sumus ego et populus meus ut conteramur iugulemur et pereamus atque utinam in servos et famulas venderemur esset tolerabile malum et gemens tacerem nunc autem hostis noster est cuius crudelitas redundat in regem
ESTH|7|5|respondensque rex Asuerus ait quis est iste et cuius potentiae ut haec audeat facere
ESTH|7|6|dixit Hester hostis et inimicus noster pessimus iste est Aman quod ille audiens ilico obstipuit vultum regis ac reginae ferre non sustinens
ESTH|7|7|rex autem surrexit iratus et de loco convivii intravit in hortum arboribus consitum Aman quoque surrexit ut rogaret Hester reginam pro anima sua intellexit enim a rege sibi paratum malum
ESTH|7|8|qui cum reversus esset de horto nemoribus consito et intrasset convivii locum repperit Aman super lectulum corruisse in quo iacebat Hester et ait etiam reginam vult opprimere me praesente in domo mea necdum verbum de ore regis exierat et statim operuerunt faciem eius
ESTH|7|9|dixitque Arbona unus de eunuchis qui stabant in ministerio regis en lignum quod paraverat Mardocheo qui locutus est pro rege stat in domo Aman habens altitudinis quinquaginta cubitos cui dixit rex adpendite eum in eo
ESTH|7|10|suspensus est itaque Aman in patibulo quod paraverat Mardocheo et regis ira quievit
ESTH|8|1|die illo dedit rex Asuerus Hester reginae domum Aman adversarii Iudaeorum et Mardocheus ingressus est ante faciem regis confessa est enim ei Hester quod esset patruus suus
ESTH|8|2|tulitque rex anulum quem ab Aman recipi iusserat et tradidit Mardocheo Hester autem constituit Mardocheum super domum suam
ESTH|8|3|nec his contenta procidit ad pedes regis flevitque et locuta ad eum oravit ut malitiam Aman Agagitae et machinationes eius pessimas quas excogitaverat contra Iudaeos iuberet irritas fieri
ESTH|8|4|at ille ex more sceptrum aureum protendit manu quo signum clementiae monstrabatur illaque consurgens stetit ante eum
ESTH|8|5|et ait si placet regi et inveni gratiam coram oculis eius et deprecatio mea non ei videtur esse contraria obsecro ut novis epistulis veteres Aman litterae insidiatoris et hostis Iudaeorum quibus eos in cunctis regis provinciis perire praeceperat corrigantur
ESTH|8|6|quomodo enim potero sustinere necem et interfectionem populi mei
ESTH|8|7|responditque rex Asuerus Hester reginae et Mardocheo Iudaeo domum Aman concessi Hester et ipsum iussi adfigi cruci qui ausus est manum in Iudaeos mittere
ESTH|8|8|scribite ergo Iudaeis sicut vobis placet ex regis nomine signantes litteras anulo meo haec enim consuetudo erat ut epistulis quae ex regis nomine mittebantur et illius anulo signatae erant nemo auderet contradicere
ESTH|8|9|accitisque scribis et librariis regis erat autem tempus tertii mensis qui appellatur siban vicesima et tertia illius die scriptae sunt epistulae ut Mardocheus voluerat ad Iudaeos et ad principes procuratoresque et iudices qui centum viginti septem provinciis ab India usque Aethiopiam praesidebant provinciae atque provinciae populo et populo iuxta linguas et litteras suas et Iudaeis ut legere poterant et audire
ESTH|8|10|ipsaeque epistulae quae ex regis nomine mittebantur anulo illius obsignatae sunt et missae per veredarios qui per omnes provincias discurrentes veteres litteras novis nuntiis praevenirent
ESTH|8|11|quibus imperavit rex ut convenirent Iudaeos per singulas civitates et in unum praeciperent congregari ut starent pro animabus suis et omnes inimicos suos cum coniugibus ac liberis et universis domibus interficerent atque delerent
ESTH|8|12|et constituta est per omnes provincias una ultionis dies id est tertiadecima mensis duodecimi adar
ESTH|8|13|summaque epistulae fuit ut in omnibus terris ac populis qui regis Asueri imperio subiacebant notum fieret paratos esse Iudaeos ad capiendam vindictam de hostibus suis
ESTH|8|14|egressique sunt veredarii celeres nuntios perferentes et edictum regis pependit in Susis
ESTH|8|15|Mardocheus autem de palatio et de conspectu regis egrediens fulgebat vestibus regiis hyacinthinis videlicet et aerinis coronam auream portans capite et amictus pallio serico atque purpureo omnisque civitas exultavit atque laetata est
ESTH|8|16|Iudaeis autem nova lux oriri visa est gaudium honor et tripudium
ESTH|8|17|apud omnes populos urbes atque provincias quocumque regis iussa veniebant mira exultatio epulae atque convivia et festus dies in tantum ut plures alterius gentis et sectae eorum religioni et caerimoniis iungerentur grandis enim cunctos iudaici nominis terror invaserat
ESTH|9|1|igitur duodecimi mensis quem adar vocari ante iam diximus tertiadecima die quando cunctis Iudaeis interfectio parabatur et hostes eorum inhiabant sanguini versa vice Iudaei superiores esse coeperunt et se de adversariis vindicare
ESTH|9|2|congregatique sunt per singulas civitates oppida et loca ut extenderent manum contra inimicos et persecutores suos nullusque ausus est resistere eo quod omnes populos magnitudinis eorum formido penetrarat
ESTH|9|3|nam et provinciarum iudices duces et procuratores omnisque dignitas quae singulis locis et operibus praeerat extollebant Iudaeos timore Mardochei
ESTH|9|4|quem principem esse palatii et plurimum posse cognoverant fama quoque nominis eius crescebat cotidie et per cunctorum ora volitabat
ESTH|9|5|itaque percusserunt Iudaei inimicos suos plaga magna et occiderunt eos reddentes eis quod sibi paraverant facere
ESTH|9|6|in tantum ut etiam in Susis quingentos viros interficerent et decem extra filios Aman Agagitae hostis Iudaeorum quorum ista sunt nomina
ESTH|9|7|Pharsandatha et Delphon et Esphata
ESTH|9|8|et Phorata et Adalia et Aridatha
ESTH|9|9|et Ephermesta et Arisai et Aridai et Vaizatha
ESTH|9|10|quos cum occidissent praedas de substantiis eorum agere noluerunt
ESTH|9|11|statimque numerus eorum qui occisi erant in Susis ad regem relatus est
ESTH|9|12|qui dixit reginae in urbe Susis interfecere Iudaei quingentos viros et alios decem filios Aman quantam putas eos exercere caedem in universis provinciis quid ultra postulas et quid vis ut fieri iubeam
ESTH|9|13|cui illa respondit si regi placet detur potestas Iudaeis ut sicut hodie fecerunt in Susis sic et cras faciant et decem filii Aman in patibulis suspendantur
ESTH|9|14|praecepitque rex ut ita fieret statimque in Susis pependit edictum et decem Aman filii suspensi sunt
ESTH|9|15|congregatis Iudaeis quartadecima adar mensis die interfecti sunt in Susis trecenti viri nec eorum ab illis direpta substantia est
ESTH|9|16|sed et per omnes provincias quae dicioni regis subiacebant pro animabus suis stetere Iudaei interfectis hostibus ac persecutoribus suis in tantum ut septuaginta quinque milia occisorum implerentur et nullus de substantiis eorum quicquam contingeret
ESTH|9|17|dies autem tertiusdecimus mensis adar unus apud omnes interfectionis fuit et quartodecimo die caedere desierunt quem constituerunt esse sollemnem ut in eo omni deinceps tempore vacarent epulis gaudio atque conviviis
ESTH|9|18|at hii qui in urbe Susis caedem exercuerant tertiodecimo et quartodecimo eiusdem mensis die in caede versati sunt quintodecimo autem die percutere desierunt et idcirco eandem diem constituere sollemnem epularum atque laetitiae
ESTH|9|19|hii vero Iudaei qui in oppidis non muratis ac villis morabantur quartumdecimum diem mensis adar conviviorum et gaudii decreverunt ita ut exultent in eo et mittant sibi mutuo partes epularum et ciborum
ESTH|9|20|scripsit itaque Mardocheus omnia haec et litteris conprehensa misit ad Iudaeos qui in omnibus regis provinciis morabantur tam in vicino positis quam procul
ESTH|9|21|ut quartamdecimam et quintamdecimam diem mensis adar pro festis susciperent et revertente semper anno sollemni honore celebrarent
ESTH|9|22|quia in ipsis diebus se ulti sunt Iudaei de inimicis suis et luctus atque tristitia in hilaritatem gaudiumque conversa sint essentque istae dies epularum atque laetitiae et mitterent sibi invicem ciborum partes et pauperibus munuscula largirentur
ESTH|9|23|susceperuntque Iudaei in sollemnem ritum cuncta quae eo tempore facere coeperant et quae Mardocheus litteris facienda mandaverat
ESTH|9|24|Aman enim filius Amadathi stirpis Agag hostis et adversarius Iudaeorum cogitavit contra eos malum ut occideret illos atque deleret et misit phur quod nostra lingua vertitur in sortem
ESTH|9|25|et postea ingressa est Hester ad regem obsecrans ut conatus eius litteris regis irriti fierent et malum quod contra Iudaeos cogitaverat reverteretur in caput eius denique et ipsum et filios eius adfixerunt cruci
ESTH|9|26|atque ex illo tempore dies isti appellati sunt Phurim id est Sortium eo quod phur id est sors in urnam missa fuerit et cuncta quae gesta sunt epistulae id est libri huius volumine continentur
ESTH|9|27|quaeque sustinuerint et quae deinceps inmutata sint suscepere Iudaei super se et semen suum et super cunctos qui religioni eorum voluerint copulari ut nulli liceat duos hos dies absque sollemnitate transigere quam scriptura testatur et certa expetunt tempora annis sibi iugiter succedentibus
ESTH|9|28|isti sunt dies quos nulla umquam delebit oblivio et per singulas generationes cunctae in toto orbe provinciae celebrabunt nec est ulla civitas in qua dies Phurim id est Sortium non observentur a Iudaeis et ab eorum progenie quae his caerimoniis obligata est
ESTH|9|29|scripseruntque Hester regina filia Abiahil et Mardocheus Iudaeus etiam secundam epistulam ut omni studio dies ista sollemnis sanciretur in posterum
ESTH|9|30|et miserunt ad omnes Iudaeos qui in centum viginti septem regis Asueri provinciis versabantur ut haberent pacem et susciperent veritatem
ESTH|9|31|observantes dies Sortium et suo tempore cum gaudio celebrarent sicut constituerat Mardocheus et Hester et illi observanda susceperant a se et a semine suo ieiunia atque clamores et Sortium dies
ESTH|9|32|et omnia quae libri huius qui vocatur Hester historia continentur
ESTH|10|1|rex vero Asuerus omnem terram et cunctas maris insulas fecit tributarias
ESTH|10|2|cuius fortitudo et imperium et dignitas atque sublimitas qua exaltavit Mardocheum scripta sunt in libris Medorum atque Persarum
ESTH|10|3|et quomodo Mardocheus iudaici generis secundus a rege Asuero fuerit et magnus inter Iudaeos et acceptabilis plebi fratrum suorum quaerens bona populo suo et loquens ea quae ad pacem sui seminis pertinerent
JOB|1|1|vir erat in terra Hus nomine Iob et erat vir ille simplex et rectus ac timens Deum et recedens a malo
JOB|1|2|natique sunt ei septem filii et tres filiae
JOB|1|3|et fuit possessio eius septem milia ovium et tria milia camelorum quingenta quoque iuga boum et quingentae asinae ac familia multa nimis eratque vir ille magnus inter omnes Orientales
JOB|1|4|et ibant filii eius et faciebant convivium per domos unusquisque in die suo et mittentes vocabant tres sorores suas ut comederent et biberent cum eis
JOB|1|5|cumque in orbem transissent dies convivii mittebat ad eos Iob et sanctificabat illos consurgensque diluculo offerebat holocausta per singulos dicebat enim ne forte peccaverint filii mei et benedixerint Deo in cordibus suis sic faciebat Iob cunctis diebus
JOB|1|6|quadam autem die cum venissent filii Dei ut adsisterent coram Domino adfuit inter eos etiam Satan
JOB|1|7|cui dixit Dominus unde venis qui respondens ait circuivi terram et perambulavi eam
JOB|1|8|dixitque Dominus ad eum numquid considerasti servum meum Iob quod non sit ei similis in terra homo simplex et rectus et timens Deum ac recedens a malo
JOB|1|9|cui respondens Satan ait numquid frustra timet Iob Deum
JOB|1|10|nonne tu vallasti eum ac domum eius universamque substantiam per circuitum operibus manuum eius benedixisti et possessio illius crevit in terra
JOB|1|11|sed extende paululum manum tuam et tange cuncta quae possidet nisi in facie tua benedixerit tibi
JOB|1|12|dixit ergo Dominus ad Satan ecce universa quae habet in manu tua sunt tantum in eum ne extendas manum tuam egressusque est Satan a facie Domini
JOB|1|13|cum autem quadam die filii et filiae eius comederent et biberent vinum in domo fratris sui primogeniti
JOB|1|14|nuntius venit ad Iob qui diceret boves arabant et asinae pascebantur iuxta eos
JOB|1|15|et inruerunt Sabei tuleruntque omnia et pueros percusserunt gladio et evasi ego solus ut nuntiarem tibi
JOB|1|16|cumque adhuc ille loqueretur venit alter et dixit ignis Dei cecidit e caelo et tactas oves puerosque consumpsit et effugi ego solus ut nuntiarem tibi
JOB|1|17|sed et illo adhuc loquente venit alius et dixit Chaldei fecerunt tres turmas et invaserunt camelos et tulerunt eos necnon et pueros percusserunt gladio et ego fugi solus ut nuntiarem tibi
JOB|1|18|loquebatur ille et ecce alius intravit et dixit filiis tuis et filiabus vescentibus et bibentibus vinum in domo fratris sui primogeniti
JOB|1|19|repente ventus vehemens inruit a regione deserti et concussit quattuor angulos domus quae corruens oppressit liberos tuos et mortui sunt et effugi ego solus ut nuntiarem tibi
JOB|1|20|tunc surrexit Iob et scidit tunicam suam et tonso capite corruens in terram adoravit
JOB|1|21|et dixit nudus egressus sum de utero matris meae et nudus revertar illuc Dominus dedit Dominus abstulit sit nomen Domini benedictum
JOB|1|22|in omnibus his non peccavit Iob neque stultum quid contra Deum locutus est
JOB|2|1|factum est autem cum quadam die venissent filii Dei et starent coram Domino venisset quoque Satan inter eos et staret in conspectu eius
JOB|2|2|ut diceret Dominus ad Satan unde venis qui respondens ait circuivi terram et perambulavi eam
JOB|2|3|et dixit Dominus ad Satan numquid considerasti servum meum Iob quod non sit ei similis in terra vir simplex et rectus timens Deum ac recedens a malo et adhuc retinens innocentiam tu autem commovisti me adversus eum ut adfligerem illum frustra
JOB|2|4|cui respondens Satan ait pellem pro pelle et cuncta quae habet homo dabit pro anima sua
JOB|2|5|alioquin mitte manum tuam et tange os eius et carnem et tunc videbis quod in facie benedicat tibi
JOB|2|6|dixit ergo Dominus ad Satan ecce in manu tua est verumtamen animam illius serva
JOB|2|7|egressus igitur Satan a facie Domini percussit Iob ulcere pessimo a planta pedis usque ad verticem eius
JOB|2|8|qui testa saniem deradebat sedens in sterquilinio
JOB|2|9|dixit autem illi uxor sua adhuc tu permanes in simplicitate tua benedic Deo et morere
JOB|2|10|qui ait ad illam quasi una de stultis locuta es si bona suscepimus de manu Domini quare mala non suscipiamus in omnibus his non peccavit Iob labiis suis
JOB|2|11|igitur audientes tres amici Iob omne malum quod accidisset ei venerunt singuli de loco suo Eliphaz Themanites et Baldad Suites et Sophar Naamathites condixerant enim ut pariter venientes visitarent eum et consolarentur
JOB|2|12|cumque levassent procul oculos suos non cognoverunt eum et exclamantes ploraverunt scissisque vestibus sparserunt pulverem super caput suum in caelum
JOB|2|13|et sederunt cum eo in terram septem diebus et septem noctibus et nemo loquebatur ei verbum videbant enim dolorem esse vehementem
JOB|3|1|post haec aperuit Iob os suum et maledixit diei suo
JOB|3|2|et locutus est
JOB|3|3|pereat dies in qua natus sum et nox in qua dictum est conceptus est homo
JOB|3|4|dies ille vertatur in tenebras non requirat eum Deus desuper et non inlustret lumine
JOB|3|5|obscurent eum tenebrae et umbra mortis occupet eum caligo et involvatur amaritudine
JOB|3|6|noctem illam tenebrosus turbo possideat non conputetur in diebus anni nec numeretur in mensibus
JOB|3|7|sit nox illa solitaria nec laude digna
JOB|3|8|maledicant ei qui maledicunt diei qui parati sunt suscitare Leviathan
JOB|3|9|obtenebrentur stellae caligine eius expectet lucem et non videat nec ortum surgentis aurorae
JOB|3|10|quia non conclusit ostia ventris qui portavit me nec abstulit mala ab oculis meis
JOB|3|11|quare non in vulva mortuus sum egressus ex utero non statim perii
JOB|3|12|quare exceptus genibus cur lactatus uberibus
JOB|3|13|nunc enim dormiens silerem et somno meo requiescerem
JOB|3|14|cum regibus et consulibus terrae qui aedificant sibi solitudines
JOB|3|15|aut cum principibus qui possident aurum et replent domos suas argento
JOB|3|16|aut sicut abortivum absconditum non subsisterem vel qui concepti non viderunt lucem
JOB|3|17|ibi impii cessaverunt a tumultu et ibi requieverunt fessi robore
JOB|3|18|et quondam vincti pariter sine molestia non audierunt vocem exactoris
JOB|3|19|parvus et magnus ibi sunt et servus liber a domino suo
JOB|3|20|quare data est misero lux et vita his qui in amaritudine animae sunt
JOB|3|21|qui expectant mortem et non venit quasi effodientes thesaurum
JOB|3|22|gaudentque vehementer cum invenerint sepulchrum
JOB|3|23|viro cuius abscondita est via et circumdedit eum Deus tenebris
JOB|3|24|antequam comedam suspiro et quasi inundantes aquae sic rugitus meus
JOB|3|25|quia timor quem timebam evenit mihi et quod verebar accidit
JOB|3|26|nonne dissimulavi nonne silui nonne quievi et venit super me indignatio
JOB|4|1|respondens autem Eliphaz Themanites dixit
JOB|4|2|si coeperimus loqui tibi forsitan moleste accipias sed conceptum sermonem tenere quis possit
JOB|4|3|ecce docuisti multos et manus lassas roborasti
JOB|4|4|vacillantes confirmaverunt sermones tui et genua trementia confortasti
JOB|4|5|nunc autem venit super te plaga et defecisti tetigit te et conturbatus es
JOB|4|6|timor tuus fortitudo tua patientia tua et perfectio viarum tuarum
JOB|4|7|recordare obsecro te quis umquam innocens perierit aut quando recti deleti sint
JOB|4|8|quin potius vidi eos qui operantur iniquitatem et seminant dolores et metunt eos
JOB|4|9|flante Deo perisse et spiritu irae eius esse consumptos
JOB|4|10|rugitus leonis et vox leaenae et dentes catulorum leonum contriti sunt
JOB|4|11|tigris periit eo quod non haberet praedam et catuli leonis dissipati sunt
JOB|4|12|porro ad me dictum est verbum absconditum et quasi furtive suscepit auris mea venas susurri eius
JOB|4|13|in horrore visionis nocturnae quando solet sopor occupare homines
JOB|4|14|pavor tenuit me et tremor et omnia ossa mea perterrita sunt
JOB|4|15|et cum spiritus me praesente transiret inhorruerunt pili carnis meae
JOB|4|16|stetit quidam cuius non agnoscebam vultum imago coram oculis meis et vocem quasi aurae lenis audivi
JOB|4|17|numquid homo Dei conparatione iustificabitur aut factore suo purior erit vir
JOB|4|18|ecce qui serviunt ei non sunt stabiles et in angelis suis repperit pravitatem
JOB|4|19|quanto magis hii qui habitant domos luteas qui terrenum habent fundamentum consumentur velut a tinea
JOB|4|20|de mane usque ad vesperum succidentur et quia nullus intellegit in aeternum peribunt
JOB|4|21|qui autem reliqui fuerint auferentur ex eis morientur et non in sapientia
JOB|5|1|voca ergo si est qui tibi respondeat et ad aliquem sanctorum convertere
JOB|5|2|vere stultum interficit iracundia et parvulum occidit invidia
JOB|5|3|ego vidi stultum firma radice et maledixi pulchritudini eius statim
JOB|5|4|longe fient filii eius a salute et conterentur in porta et non erit qui eruat
JOB|5|5|cuius messem famelicus comedet et ipsum rapiet armatus et ebibent sitientes divitias eius
JOB|5|6|nihil in terra sine causa fit et de humo non orietur dolor
JOB|5|7|homo ad laborem nascitur et avis ad volatum
JOB|5|8|quam ob rem ego deprecabor Dominum et ad Deum ponam eloquium meum
JOB|5|9|qui facit magna et inscrutabilia et mirabilia absque numero
JOB|5|10|qui dat pluviam super faciem terrae et inrigat aquis universa
JOB|5|11|qui ponit humiles in sublimi et maerentes erigit sospitate
JOB|5|12|qui dissipat cogitationes malignorum ne possint implere manus eorum quod coeperant
JOB|5|13|qui adprehendit sapientes in astutia eorum et consilium pravorum dissipat
JOB|5|14|per diem incurrent tenebras et quasi in nocte sic palpabunt in meridie
JOB|5|15|porro salvum faciet a gladio oris eorum et de manu violenti pauperem
JOB|5|16|et erit egeno spes iniquitas autem contrahet os suum
JOB|5|17|beatus homo qui corripitur a Domino increpationem ergo Domini ne reprobes
JOB|5|18|quia ipse vulnerat et medetur percutit et manus eius sanabunt
JOB|5|19|in sex tribulationibus liberabit te et in septima non tanget te malum
JOB|5|20|in fame eruet te de morte et in bello de manu gladii
JOB|5|21|a flagello linguae absconderis et non timebis calamitatem cum venerit
JOB|5|22|in vastitate et fame ridebis et bestiam terrae non formidabis
JOB|5|23|sed cum lapidibus regionum pactum tuum et bestiae terrae pacificae erunt tibi
JOB|5|24|et scies quod pacem habeat tabernaculum tuum et visitans speciem tuam non peccabis
JOB|5|25|scies quoque quoniam multiplex erit semen tuum et progenies tua quasi herba terrae
JOB|5|26|ingredieris in abundantia sepulchrum sicut infertur acervus in tempore suo
JOB|5|27|ecce hoc ut investigavimus ita est quod auditum mente pertracta
JOB|6|1|respondens autem Iob dixit
JOB|6|2|utinam adpenderentur peccata mea quibus iram merui et calamitas quam patior in statera
JOB|6|3|quasi harena maris haec gravior appareret unde et verba mea dolore sunt plena
JOB|6|4|quia sagittae Domini in me sunt quarum indignatio ebibit spiritum meum et terrores Domini militant contra me
JOB|6|5|numquid rugiet onager cum habuerit herbam aut mugiet bos cum ante praesepe plenum steterit
JOB|6|6|aut poterit comedi insulsum quod non est sale conditum aut potest aliquis gustare quod gustatum adfert mortem
JOB|6|7|quae prius tangere nolebat anima mea nunc prae angustia cibi mei sunt
JOB|6|8|quis det ut veniat petitio mea et quod expecto tribuat mihi Deus
JOB|6|9|et qui coepit ipse me conterat solvat manum suam et succidat me
JOB|6|10|et haec mihi sit consolatio ut adfligens me dolore non parcat nec contradicam sermonibus Sancti
JOB|6|11|quae est enim fortitudo mea ut sustineam aut quis finis meus ut patienter agam
JOB|6|12|nec fortitudo lapidum fortitudo mea nec caro mea aerea est
JOB|6|13|ecce non est auxilium mihi in me et necessarii quoque mei recesserunt a me
JOB|6|14|qui tollit ab amico suo misericordiam timorem Domini derelinquit
JOB|6|15|fratres mei praeterierunt me sicut torrens qui raptim transit in convallibus
JOB|6|16|qui timent pruinam inruet super eos nix
JOB|6|17|tempore quo fuerint dissipati peribunt et ut incaluerit solventur de loco suo
JOB|6|18|involutae sunt semitae gressuum eorum ambulabunt in vacuum et peribunt
JOB|6|19|considerate semitas Theman itinera Saba et expectate paulisper
JOB|6|20|confusi sunt quia speravi venerunt quoque usque ad me et pudore cooperti sunt
JOB|6|21|nunc venistis et modo videntes plagam meam timetis
JOB|6|22|numquid dixi adferte mihi et de substantia vestra donate mihi
JOB|6|23|vel liberate me de manu hostis et de manu robustorum eruite me
JOB|6|24|docete me et ego tacebo et si quid forte ignoravi instruite me
JOB|6|25|quare detraxistis sermonibus veritatis cum e vobis nullus sit qui possit arguere
JOB|6|26|ad increpandum tantum eloquia concinnatis et in ventum verba profertis
JOB|6|27|super pupillum inruitis et subvertere nitimini amicum vestrum
JOB|6|28|verumtamen quod coepistis explete praebete aurem et videte an mentiar
JOB|6|29|respondete obsecro absque contentione et loquentes id quod iustum est iudicate
JOB|6|30|et non invenietis in lingua mea iniquitatem nec in faucibus meis stultitia personabit
JOB|7|1|militia est vita hominis super terram et sicut dies mercennarii dies eius
JOB|7|2|sicut servus desiderat umbram et sicut mercennarius praestolatur finem operis sui
JOB|7|3|sic et ego habui menses vacuos et noctes laboriosas enumeravi mihi
JOB|7|4|si dormiero dico quando consurgam et rursum expectabo vesperam et replebor doloribus usque ad tenebras
JOB|7|5|induta est caro mea putredine et sordibus pulveris cutis mea aruit et contracta est
JOB|7|6|dies mei velocius transierunt quam a texente tela succiditur et consumpti sunt absque ulla spe
JOB|7|7|memento quia ventus est vita mea et non revertetur oculus meus ut videat bona
JOB|7|8|nec aspiciet me visus hominis oculi tui in me et non subsistam
JOB|7|9|sicut consumitur nubes et pertransit sic qui descenderit ad inferos non ascendet
JOB|7|10|nec revertetur ultra in domum suam neque cognoscet eum amplius locus eius
JOB|7|11|quapropter et ego non parcam ori meo loquar in tribulatione spiritus mei confabulabor cum amaritudine animae meae
JOB|7|12|numquid mare sum ego aut cetus quia circumdedisti me carcere
JOB|7|13|si dixero consolabitur me lectulus meus et relevabor loquens mecum in strato meo
JOB|7|14|terrebis me per somnia et per visiones horrore concuties
JOB|7|15|quam ob rem elegit suspendium anima mea et mortem ossa mea
JOB|7|16|desperavi nequaquam ultra iam vivam parce mihi nihil enim sunt dies mei
JOB|7|17|quid est homo quia magnificas eum aut quia ponis erga eum cor tuum
JOB|7|18|visitas eum diluculo et subito probas illum
JOB|7|19|usquequo non parces mihi nec dimittis me ut gluttiam salivam meam
JOB|7|20|peccavi quid faciam tibi o custos hominum quare posuisti me contrarium tibi et factus sum mihimet ipsi gravis
JOB|7|21|cur non tolles peccatum meum et quare non auferes iniquitatem meam ecce nunc in pulvere dormiam et si mane me quaesieris non subsistam
JOB|8|1|respondens autem Baldad Suites dixit
JOB|8|2|usquequo loqueris talia et spiritus multiplex sermones oris tui
JOB|8|3|numquid Deus subplantat iudicium et Omnipotens subvertit quod iustum est
JOB|8|4|etiam si filii tui peccaverunt ei et dimisit eos in manu iniquitatis suae
JOB|8|5|tu tamen si diluculo consurrexeris ad Deum et Omnipotentem fueris deprecatus
JOB|8|6|si mundus et rectus incesseris statim evigilabit ad te et pacatum reddet habitaculum iustitiae tuae
JOB|8|7|in tantum ut priora tua fuerint parva et novissima tua multiplicentur nimis
JOB|8|8|interroga enim generationem pristinam et diligenter investiga patrum memoriam
JOB|8|9|hesterni quippe sumus et ignoramus quoniam sicut umbra dies nostri sunt super terram
JOB|8|10|et ipsi docebunt te loquentur tibi et de corde suo proferent eloquia
JOB|8|11|numquid vivere potest scirpus absque humore aut crescet carectum sine aqua
JOB|8|12|cum adhuc sit in flore nec carpatur manu ante omnes herbas arescit
JOB|8|13|sic viae omnium qui obliviscuntur Deum et spes hypocritae peribit
JOB|8|14|non ei placebit vecordia sua et sicut tela aranearum fiducia eius
JOB|8|15|innitetur super domum suam et non stabit fulciet eam et non consurget
JOB|8|16|humectus videtur antequam veniat sol et in horto suo germen eius egreditur
JOB|8|17|super acervum petrarum radices eius densabuntur et inter lapides commorabitur
JOB|8|18|si absorbuerit eum de loco suo negabit eum et dicet non novi te
JOB|8|19|haec est enim laetitia viae eius ut rursum de terra alii germinentur
JOB|8|20|Deus non proiciet simplicem nec porriget manum malignis
JOB|8|21|donec impleatur risu os tuum et labia tua iubilo
JOB|8|22|qui oderunt te induentur confusione et tabernaculum impiorum non subsistet
JOB|9|1|et respondens Iob ait
JOB|9|2|vere scio quod ita sit et quod non iustificetur homo conpositus Deo
JOB|9|3|si voluerit contendere cum eo non poterit ei respondere unum pro mille
JOB|9|4|sapiens corde est et fortis robore quis restitit ei et pacem habuit
JOB|9|5|qui transtulit montes et nescierunt hii quos subvertit in furore suo
JOB|9|6|qui commovet terram de loco suo et columnae eius concutiuntur
JOB|9|7|qui praecipit soli et non oritur et stellas claudit quasi sub signaculo
JOB|9|8|qui extendit caelos solus et graditur super fluctus maris
JOB|9|9|qui facit Arcturum et Oriona et Hyadas et interiora austri
JOB|9|10|qui facit magna et inconprehensibilia et mirabilia quorum non est numerus
JOB|9|11|si venerit ad me non videbo si abierit non intellegam eum
JOB|9|12|si repente interroget quis respondebit ei vel quis dicere potest cur facis
JOB|9|13|Deus cuius resistere irae nemo potest et sub quo curvantur qui portant orbem
JOB|9|14|quantus ergo sum ego qui respondeam ei et loquar verbis meis cum eo
JOB|9|15|qui etiam si habuero quippiam iustum non respondebo sed meum iudicem deprecabor
JOB|9|16|et cum invocantem exaudierit me non credo quod audierit vocem meam
JOB|9|17|in turbine enim conteret me et multiplicabit vulnera mea etiam sine causa
JOB|9|18|non concedit requiescere spiritum meum et implet me amaritudinibus
JOB|9|19|si fortitudo quaeritur robustissimus est si aequitas iudicii nemo pro me audet testimonium dicere
JOB|9|20|si iustificare me voluero os meum condemnabit me si innocentem ostendere pravum me conprobabit
JOB|9|21|etiam si simplex fuero hoc ipsum ignorabit anima mea et taedebit me vitae meae
JOB|9|22|unum est quod locutus sum et innocentem et impium ipse consumit
JOB|9|23|si flagellat occidat semel et non de poenis innocentum rideat
JOB|9|24|terra data est in manu impii vultum iudicum eius operit quod si non ille est quis ergo est
JOB|9|25|dies mei velociores fuerunt cursore fugerunt et non viderunt bonum
JOB|9|26|pertransierunt quasi naves poma portantes sicut aquila volans ad escam
JOB|9|27|cum dixero nequaquam ita loquar commuto faciem meam et dolore torqueor
JOB|9|28|verebar omnia opera mea sciens quod non parceres delinquenti
JOB|9|29|si autem et sic impius sum quare frustra laboravi
JOB|9|30|si lotus fuero quasi aquis nivis et fulserint velut mundissimae manus meae
JOB|9|31|tamen sordibus intingues me et abominabuntur me vestimenta mea
JOB|9|32|neque enim viro qui similis mei est respondebo nec qui mecum in iudicio ex aequo possit audiri
JOB|9|33|non est qui utrumque valeat arguere et ponere manum suam in ambobus
JOB|9|34|auferat a me virgam suam et pavor eius non me terreat
JOB|9|35|loquar et non timebo eum neque enim possum metuens respondere
JOB|10|1|taedet animam meam vitae meae dimittam adversum me eloquium meum loquar in amaritudine animae meae
JOB|10|2|dicam Deo noli me condemnare indica mihi cur me ita iudices
JOB|10|3|numquid bonum tibi videtur si calumnieris et opprimas me opus manuum tuarum et consilium impiorum adiuves
JOB|10|4|numquid oculi carnei tibi sunt aut sicut videt homo et tu videbis
JOB|10|5|numquid sicut dies hominis dies tui et anni tui sicut humana sunt tempora
JOB|10|6|ut quaeras iniquitatem meam et peccatum meum scruteris
JOB|10|7|et scias quia nihil impium fecerim cum sit nemo qui de manu tua possit eruere
JOB|10|8|manus tuae plasmaverunt me et fecerunt me totum in circuitu et sic repente praecipitas me
JOB|10|9|memento quaeso quod sicut lutum feceris me et in pulverem reduces me
JOB|10|10|nonne sicut lac mulsisti me et sicut caseum me coagulasti
JOB|10|11|pelle et carnibus vestisti me et ossibus et nervis conpegisti me
JOB|10|12|vitam et misericordiam tribuisti mihi et visitatio tua custodivit spiritum meum
JOB|10|13|licet haec celes in corde tuo tamen scio quia universorum memineris
JOB|10|14|si peccavi et ad horam pepercisti mihi cur ab iniquitate mea mundum me esse non pateris
JOB|10|15|et si impius fuero vae mihi est et si iustus non levabo caput saturatus adflictione et miseria
JOB|10|16|et propter superbiam quasi leaenam capies me reversusque mirabiliter me crucias
JOB|10|17|instauras testes tuos contra me et multiplicas iram tuam adversum me et poenae militant in me
JOB|10|18|quare de vulva eduxisti me qui utinam consumptus essem ne oculus me videret
JOB|10|19|fuissem quasi qui non essem de utero translatus ad tumulum
JOB|10|20|numquid non paucitas dierum meorum finietur brevi dimitte ergo me ut plangam paululum dolorem meum
JOB|10|21|antequam vadam et non revertar ad terram tenebrosam et opertam mortis caligine
JOB|10|22|terram miseriae et tenebrarum ubi umbra mortis et nullus ordo et sempiternus horror inhabitans
JOB|11|1|respondens autem Sophar Naamathites dixit
JOB|11|2|numquid qui multa loquitur non et audiet aut vir verbosus iustificabitur
JOB|11|3|tibi soli tacebunt homines et cum ceteros inriseris a nullo confutaberis
JOB|11|4|dixisti enim purus est sermo meus et mundus sum in conspectu tuo
JOB|11|5|atque utinam Deus loqueretur tecum et aperiret labia sua tibi
JOB|11|6|ut ostenderet tibi secreta sapientiae et quod multiplex esset lex eius et intellegeres quod multo minora exigaris a Deo quam meretur iniquitas tua
JOB|11|7|forsitan vestigia Dei conprehendes et usque ad perfectum Omnipotentem repperies
JOB|11|8|excelsior caelo est et quid facies profundior inferno et unde cognosces
JOB|11|9|longior terrae mensura eius et latior mari
JOB|11|10|si subverterit omnia vel in unum coartaverit quis contradicet ei
JOB|11|11|ipse enim novit hominum vanitatem et videns iniquitatem nonne considerat
JOB|11|12|vir vanus in superbiam erigitur et tamquam pullum onagri se liberum natum putat
JOB|11|13|tu autem firmasti cor tuum et expandisti ad eum manus tuas
JOB|11|14|si iniquitatem quod est in manu tua abstuleris a te et non manserit in tabernaculo tuo iniustitia
JOB|11|15|tum levare poteris faciem tuam absque macula et eris stabilis et non timebis
JOB|11|16|miseriae quoque oblivisceris et quasi aquarum quae praeterierint recordaberis
JOB|11|17|et quasi meridianus fulgor consurget tibi ad vesperam et cum te consumptum putaveris orieris ut lucifer
JOB|11|18|et habebis fiduciam proposita tibi spe et defossus securus dormies
JOB|11|19|requiesces et non erit qui te exterreat et deprecabuntur faciem tuam plurimi
JOB|11|20|oculi autem impiorum deficient et effugium peribit ab eis et spes eorum abominatio animae
JOB|12|1|respondens autem Iob dixit
JOB|12|2|ergo vos estis soli homines et vobiscum morietur sapientia
JOB|12|3|et mihi est cor sicut et vobis nec inferior vestri sum quis enim haec quae nostis ignorat
JOB|12|4|qui deridetur ab amico suo sicut ego invocabit Deum et exaudiet eum deridetur enim iusti simplicitas
JOB|12|5|lampas contempta apud cogitationes divitum parata ad tempus statutum
JOB|12|6|abundant tabernacula praedonum et audacter provocant Deum cum ipse dederit omnia in manibus eorum
JOB|12|7|nimirum interroga iumenta et docebunt te et volatilia caeli et indicabunt tibi
JOB|12|8|loquere terrae et respondebit tibi et narrabunt pisces maris
JOB|12|9|quis ignorat quod omnia haec manus Domini fecerit
JOB|12|10|in cuius manu anima omnis viventis et spiritus universae carnis hominis
JOB|12|11|nonne auris verba diiudicat et fauces comedentis saporem
JOB|12|12|in antiquis est sapientia et in multo tempore prudentia
JOB|12|13|apud ipsum est sapientia et fortitudo ipse habet consilium et intellegentiam
JOB|12|14|si destruxerit nemo est qui aedificet et si incluserit hominem nullus est qui aperiat
JOB|12|15|si continuerit aquas omnia siccabuntur et si emiserit eas subvertent terram
JOB|12|16|apud ipsum est fortitudo et sapientia ipse novit et decipientem et eum qui decipitur
JOB|12|17|adducit consiliarios in stultum finem et iudices in stuporem
JOB|12|18|balteum regum dissolvit et praecingit fune renes eorum
JOB|12|19|ducit sacerdotes inglorios et optimates subplantat
JOB|12|20|commutans labium veracium et doctrinam senum auferens
JOB|12|21|effundit despectionem super principes et eos qui oppressi fuerant relevans
JOB|12|22|qui revelat profunda de tenebris et producit in lucem umbram mortis
JOB|12|23|qui multiplicat gentes et perdet eas et subversas in integrum restituet
JOB|12|24|qui inmutat cor principum populi terrae et decipit eos ut frustra incedant per invium
JOB|12|25|palpabunt quasi in tenebris et non in luce et errare eos faciet quasi ebrios
JOB|13|1|ecce omnia et vidit oculus meus et audivit auris mea et intellexi singula
JOB|13|2|secundum scientiam vestram et ego novi nec inferior vestri sum
JOB|13|3|sed tamen ad Omnipotentem loquar et disputare cum Deo cupio
JOB|13|4|prius vos ostendens fabricatores mendacii et cultores perversorum dogmatum
JOB|13|5|atque utinam taceretis ut putaremini esse sapientes
JOB|13|6|audite ergo correptiones meas et iudicium labiorum meorum adtendite
JOB|13|7|numquid Deus indiget vestro mendacio ut pro illo loquamini dolos
JOB|13|8|numquid faciem eius accipitis et pro Deo iudicare nitimini
JOB|13|9|aut placebit ei quem celare nihil potest aut decipietur ut homo vestris fraudulentiis
JOB|13|10|ipse vos arguet quoniam in abscondito faciem eius accipitis
JOB|13|11|statim ut se commoverit turbabit vos et terror eius inruet super vos
JOB|13|12|memoria vestra conparabitur cineri et redigentur in lutum cervices vestrae
JOB|13|13|tacete paulisper ut loquar quodcumque mihi mens suggesserit
JOB|13|14|quare lacero carnes meas dentibus meis et animam meam porto in manibus meis
JOB|13|15|etiam si occiderit me in ipso sperabo verumtamen vias meas in conspectu eius arguam
JOB|13|16|et ipse erit salvator meus non enim veniet in conspectu eius omnis hypocrita
JOB|13|17|audite sermonem meum et enigmata percipite auribus vestris
JOB|13|18|si fuero iudicatus scio quod iustus inveniar
JOB|13|19|quis est qui iudicetur mecum veniat quare tacens consumor
JOB|13|20|duo tantum ne facias mihi et tunc a facie tua non abscondar
JOB|13|21|manum tuam longe fac a me et formido tua non me terreat
JOB|13|22|et voca me et respondebo tibi aut certe loquar et tu responde mihi
JOB|13|23|quantas habeo iniquitates et peccata scelera mea et delicta ostende mihi
JOB|13|24|cur faciem tuam abscondis et arbitraris me inimicum tuum
JOB|13|25|contra folium quod vento rapitur ostendis potentiam tuam et stipulam siccam persequeris
JOB|13|26|scribis enim contra me amaritudines et consumere me vis peccatis adulescentiae meae
JOB|13|27|posuisti in nervo pedem meum et observasti omnes semitas meas et vestigia pedum meorum considerasti
JOB|13|28|qui quasi putredo consumendus sum et quasi vestimentum quod comeditur a tinea
JOB|14|1|homo natus de muliere brevi vivens tempore repletus multis miseriis
JOB|14|2|quasi flos egreditur et conteritur et fugit velut umbra et numquam in eodem statu permanet
JOB|14|3|et dignum ducis super huiuscemodi aperire oculos tuos et adducere eum tecum in iudicium
JOB|14|4|quis potest facere mundum de inmundo conceptum semine nonne tu qui solus es
JOB|14|5|breves dies hominis sunt numerus mensuum eius apud te est constituisti terminos eius qui praeterire non poterunt
JOB|14|6|recede paululum ab eo ut quiescat donec optata veniat sicut mercennarii dies eius
JOB|14|7|lignum habet spem si praecisum fuerit rursum virescit et rami eius pullulant
JOB|14|8|si senuerit in terra radix eius et in pulvere emortuus fuerit truncus illius
JOB|14|9|ad odorem aquae germinabit et faciet comam quasi cum primum plantatum est
JOB|14|10|homo vero cum mortuus fuerit et nudatus atque consumptus ubi quaeso est
JOB|14|11|quomodo si recedant aquae de mari et fluvius vacuefactus arescat
JOB|14|12|sic homo cum dormierit non resurget donec adteratur caelum non evigilabit nec consurget de somno suo
JOB|14|13|quis mihi hoc tribuat ut in inferno protegas me ut abscondas me donec pertranseat furor tuus et constituas mihi tempus in quo recorderis mei
JOB|14|14|putasne mortuus homo rursum vivet cunctis diebus quibus nunc milito expecto donec veniat inmutatio mea
JOB|14|15|vocabis et ego respondebo tibi operi manuum tuarum porriges dexteram
JOB|14|16|tu quidem gressus meos dinumerasti sed parces peccatis meis
JOB|14|17|signasti quasi in sacculo delicta mea sed curasti iniquitatem meam
JOB|14|18|mons cadens defluet et saxum transfertur de loco suo
JOB|14|19|lapides excavant aquae et adluvione paulatim terra consumitur et homines ergo similiter perdes
JOB|14|20|roborasti eum paululum ut in perpetuum pertransiret inmutabis faciem eius et emittes eum
JOB|14|21|sive nobiles fuerint filii eius sive ignobiles non intelleget
JOB|14|22|attamen caro eius dum vivet dolebit et anima illius super semet ipso lugebit
JOB|15|1|respondens autem Eliphaz Themanites dixit
JOB|15|2|numquid sapiens respondebit quasi in ventum loquens et implebit ardore stomachum suum
JOB|15|3|arguis verbis eum qui non est aequalis tui et loqueris quod tibi non expedit
JOB|15|4|quantum in te est evacuasti timorem et tulisti preces coram Deo
JOB|15|5|docuit enim iniquitas tua os tuum et imitaris linguam blasphemantium
JOB|15|6|condemnabit te os tuum et non ego et labia tua respondebunt tibi
JOB|15|7|numquid primus homo tu natus es et ante colles formatus
JOB|15|8|numquid consilium Dei audisti et inferior te erit eius sapientia
JOB|15|9|quid nosti quod ignoremus quid intellegis quod nesciamus
JOB|15|10|et senes et antiqui sunt in nobis multo vetustiores quam patres tui
JOB|15|11|numquid grande est ut consoletur te Deus sed verba tua prava hoc prohibent
JOB|15|12|quid te elevat cor tuum et quasi magna cogitans adtonitos habes oculos
JOB|15|13|quid tumet contra Deum spiritus tuus ut proferas de ore huiuscemodi sermones
JOB|15|14|quid est homo ut inmaculatus sit et ut iustus appareat natus de muliere
JOB|15|15|ecce inter sanctos eius nemo inmutabilis et caeli non sunt mundi in conspectu eius
JOB|15|16|quanto magis abominabilis et inutilis homo qui bibit quasi aquas iniquitatem
JOB|15|17|ostendam tibi audi me quod vidi narrabo tibi
JOB|15|18|sapientes confitentur et non abscondunt patres suos
JOB|15|19|quibus solis data est terra et non transibit alienus per eos
JOB|15|20|cunctis diebus suis impius superbit et numerus annorum incertus est tyrannidis eius
JOB|15|21|sonitus terroris semper in auribus illius et cum pax sit ille insidias suspicatur
JOB|15|22|non credit quod reverti possit de tenebris circumspectans undique gladium
JOB|15|23|cum se moverit ad quaerendum panem novit quod paratus sit in manu eius tenebrarum dies
JOB|15|24|terrebit eum tribulatio et angustia vallabit eum sicut regem qui praeparatur ad proelium
JOB|15|25|tetendit enim adversus Deum manum suam et contra Omnipotentem roboratus est
JOB|15|26|cucurrit adversus eum erecto collo et pingui cervice armatus est
JOB|15|27|operuit faciem eius crassitudo et de lateribus eius arvina dependet
JOB|15|28|habitavit in civitatibus desolatis et in domibus desertis quae in tumulos sunt redactae
JOB|15|29|non ditabitur nec perseverabit substantia eius nec mittet in terra radicem suam
JOB|15|30|non recedet de tenebris ramos eius arefaciet flamma et auferetur spiritu oris sui
JOB|15|31|non credat frustra errore deceptus quod aliquo pretio redimendus sit
JOB|15|32|antequam dies eius impleantur peribit et manus eius arescet
JOB|15|33|laedetur quasi vinea in primo flore botrus eius et quasi oliva proiciens florem suum
JOB|15|34|congregatio enim hypocritae sterilis et ignis devorabit tabernacula eorum qui munera libenter accipiunt
JOB|15|35|concepit dolorem et peperit iniquitatem et uterus eius praeparat dolos
JOB|16|1|respondens autem Iob dixit
JOB|16|2|audivi frequenter talia consolatores onerosi omnes vos estis
JOB|16|3|numquid habebunt finem verba ventosa aut aliquid tibi molestum est si loquaris
JOB|16|4|poteram et ego similia vestri loqui atque utinam esset anima vestra pro anima mea
JOB|16|5|consolarer et ego vos sermonibus et moverem caput meum super vos
JOB|16|6|roborarem vos ore meo et moverem labia quasi parcens vobis
JOB|16|7|sed quid agam si locutus fuero non quiescet dolor meus et si tacuero non recedet a me
JOB|16|8|nunc autem oppressit me dolor meus et in nihili redacti sunt omnes artus mei
JOB|16|9|rugae meae testimonium dicunt contra me et suscitatur falsiloquus adversus faciem meam contradicens mihi
JOB|16|10|collegit furorem suum in me et comminans mihi infremuit contra me dentibus suis hostis meus terribilibus oculis me intuitus est
JOB|16|11|aperuerunt super me ora sua exprobrantes percusserunt maxillam meam satiati sunt poenis meis
JOB|16|12|conclusit me Deus apud iniquum et manibus impiorum me tradidit
JOB|16|13|ego ille quondam opulentus repente contritus sum tenuit cervicem meam confregit me et posuit sibi quasi in signum
JOB|16|14|circumdedit me lanceis suis convulneravit lumbos meos non pepercit et effudit in terra viscera mea
JOB|16|15|concidit me vulnere super vulnus inruit in me quasi gigans
JOB|16|16|saccum consui super cutem meam et operui cinere cornu meum
JOB|16|17|facies mea intumuit a fletu et palpebrae meae caligaverunt
JOB|16|18|haec passus sum absque iniquitate manus meae cum haberem mundas ad Deum preces
JOB|16|19|terra ne operias sanguinem meum neque inveniat locum in te latendi clamor meus
JOB|16|20|ecce enim in caelo testis meus et conscius meus in excelsis
JOB|16|21|verbosi mei amici mei ad Deum stillat oculus meus
JOB|16|22|atque utinam sic iudicaretur vir cum Deo quomodo iudicatur filius hominis cum collega suo
JOB|16|23|ecce enim breves anni transeunt et semitam per quam non revertar ambulo
JOB|17|1|spiritus meus adtenuabitur dies mei breviabuntur et solum mihi superest sepulchrum
JOB|17|2|non peccavi et in amaritudinibus moratur oculus meus
JOB|17|3|libera me et pone iuxta te et cuiusvis manus pugnet contra me
JOB|17|4|cor eorum longe fecisti a disciplina et propterea non exaltabuntur
JOB|17|5|praedam pollicetur sociis et oculi filiorum eius deficient
JOB|17|6|posuit me quasi in proverbium vulgi et exemplum sum coram eis
JOB|17|7|caligavit ab indignatione oculus meus et membra mea quasi in nihili redacta sunt
JOB|17|8|stupebunt iusti super hoc et innocens contra hypocritam suscitabitur
JOB|17|9|et tenebit iustus viam suam et mundis manibus addet fortitudinem
JOB|17|10|igitur vos omnes convertimini et venite et non inveniam in vobis ullum sapientem
JOB|17|11|dies mei transierunt cogitationes meae dissipatae sunt torquentes cor meum
JOB|17|12|noctem verterunt in diem et rursum post tenebras spero lucem
JOB|17|13|si sustinuero infernus domus mea est in tenebris stravi lectulum meum
JOB|17|14|putredini dixi pater meus es mater mea et soror mea vermibus
JOB|17|15|ubi est ergo nunc praestolatio mea et patientiam meam quis considerat
JOB|17|16|in profundissimum infernum descendent omnia mea putasne saltim ibi erit requies mihi
JOB|18|1|respondens autem Baldad Suites dixit
JOB|18|2|usque ad quem finem verba iactabitis intellegite prius et sic loquamur
JOB|18|3|quare reputati sumus ut iumenta et sorduimus coram vobis
JOB|18|4|qui perdis animam tuam in furore tuo numquid propter te derelinquetur terra et transferentur rupes de loco suo
JOB|18|5|nonne lux impii extinguetur nec splendebit flamma ignis eius
JOB|18|6|lux obtenebrescet in tabernaculo illius et lucerna quae super eum est extinguetur
JOB|18|7|artabuntur gressus virtutis eius et praecipitabit eum consilium suum
JOB|18|8|inmisit enim in rete pedes suos et in maculis eius ambulat
JOB|18|9|tenebitur planta illius laqueo et exardescet contra eum sitis
JOB|18|10|abscondita est in terra pedica eius et decipula illius super semitam
JOB|18|11|undique terrebunt eum formidines et involvent pedes eius
JOB|18|12|adtenuetur fame robur eius et inedia invadat costas illius
JOB|18|13|devoret pulchritudinem cutis eius consumat brachia illius primogenita mors
JOB|18|14|avellatur de tabernaculo suo fiducia eius et calcet super eum quasi rex interitus
JOB|18|15|habitent in tabernaculo illius socii eius qui non est aspergatur in tabernaculo eius sulphur
JOB|18|16|deorsum radices eius siccentur sursum autem adteratur messis eius
JOB|18|17|memoria illius pereat de terra et non celebretur nomen eius in plateis
JOB|18|18|expellet eum de luce in tenebras et de orbe transferet eum
JOB|18|19|non erit semen eius neque progenies in populo suo nec ullae reliquiae in regionibus eius
JOB|18|20|in die eius stupebunt novissimi et primos invadet horror
JOB|18|21|haec sunt ergo tabernacula iniqui et iste locus eius qui ignorat Deum
JOB|19|1|respondens autem Iob dixit
JOB|19|2|usquequo adfligitis animam meam et adteritis me sermonibus
JOB|19|3|en decies confunditis me et non erubescitis opprimentes me
JOB|19|4|nempe et si ignoravi mecum erit ignorantia mea
JOB|19|5|at vos contra me erigimini et arguitis me obprobriis meis
JOB|19|6|saltim nunc intellegite quia Deus non aequo iudicio adflixerit me et flagellis suis me cinxerit
JOB|19|7|ecce clamabo vim patiens et nemo audiet vociferabor et non est qui iudicet
JOB|19|8|semitam meam circumsepsit et transire non possum et in calle meo tenebras posuit
JOB|19|9|spoliavit me gloria mea et abstulit coronam de capite meo
JOB|19|10|destruxit me undique et pereo et quasi evulsae arbori abstulit spem meam
JOB|19|11|iratus est contra me furor eius et sic me habuit quasi hostem suum
JOB|19|12|simul venerunt latrones eius et fecerunt sibi viam per me et obsederunt in gyro tabernaculum meum
JOB|19|13|fratres meos longe fecit a me et noti mei quasi alieni recesserunt a me
JOB|19|14|dereliquerunt me propinqui mei et qui me noverant obliti sunt mei
JOB|19|15|inquilini domus meae et ancillae meae sicut alienum habuerunt me et quasi peregrinus fui in oculis eorum
JOB|19|16|servum meum vocavi et non respondit ore proprio deprecabar illum
JOB|19|17|halitum meum exhorruit uxor mea et orabam filios uteri mei
JOB|19|18|stulti quoque despiciebant me et cum ab eis recessissem detrahebant mihi
JOB|19|19|abominati sunt me quondam consiliarii mei et quem maxime diligebam aversatus est me
JOB|19|20|pelli meae consumptis carnibus adhesit os meum et derelicta sunt tantummodo labia circa dentes meos
JOB|19|21|miseremini mei miseremini mei saltim vos amici mei quia manus Domini tetigit me
JOB|19|22|quare persequimini me sicut Deus et carnibus meis saturamini
JOB|19|23|quis mihi tribuat ut scribantur sermones mei quis mihi det ut exarentur in libro
JOB|19|24|stilo ferreo et plumbi lammina vel certe sculpantur in silice
JOB|19|25|scio enim quod redemptor meus vivat et in novissimo de terra surrecturus sim
JOB|19|26|et rursum circumdabor pelle mea et in carne mea videbo Deum
JOB|19|27|quem visurus sum ego ipse et oculi mei conspecturi sunt et non alius reposita est haec spes mea in sinu meo
JOB|19|28|quare ergo nunc dicitis persequamur eum et radicem verbi inveniamus contra eum
JOB|19|29|fugite ergo a facie gladii quoniam ultor iniquitatum gladius est et scitote esse iudicium
JOB|20|1|respondens autem Sophar Naamathites dixit
JOB|20|2|idcirco cogitationes meae variae succedunt sibi et mens in diversa rapitur
JOB|20|3|doctrinam qua me arguis audiam et spiritus intellegentiae meae respondebit mihi
JOB|20|4|hoc scio a principio ex quo positus est homo super terram
JOB|20|5|quod laus impiorum brevis sit et gaudium hypocritae ad instar puncti
JOB|20|6|si ascenderit usque ad caelum superbia eius et caput eius nubes tetigerit
JOB|20|7|quasi sterquilinium in fine perdetur et qui eum viderant dicent ubi est
JOB|20|8|velut somnium avolans non invenietur transiet sicut visio nocturna
JOB|20|9|oculus qui eum viderat non videbit neque ultra intuebitur eum locus suus
JOB|20|10|filii eius adterentur egestate et manus illius reddent ei dolorem suum
JOB|20|11|ossa eius implebuntur vitiis adulescentiae eius et cum eo in pulverem dormient
JOB|20|12|cum enim dulce fuerit in ore eius malum abscondet illud sub lingua sua
JOB|20|13|parcet illi et non derelinquet illud et celabit in gutture suo
JOB|20|14|panis eius in utero illius vertetur in fel aspidum intrinsecus
JOB|20|15|divitias quas devoravit evomet et de ventre illius extrahet eas Deus
JOB|20|16|caput aspidum suget occidet eum lingua viperae
JOB|20|17|non videat rivulos fluminis torrentes mellis et butyri
JOB|20|18|luet quae fecit omnia nec tamen consumetur iuxta multitudinem adinventionum suarum sic et sustinebit
JOB|20|19|quoniam confringens nudavit pauperes domum rapuit et non aedificavit eam
JOB|20|20|nec est satiatus venter eius et cum habuerit quae cupierat possidere non poterit
JOB|20|21|non remansit de cibo eius et propterea nihil permanebit de bonis eius
JOB|20|22|cum satiatus fuerit artabitur aestuabit et omnis dolor inruet in eum
JOB|20|23|utinam impleatur venter eius ut emittat in eum iram furoris sui et pluat super illum bellum suum
JOB|20|24|fugiet arma ferrea et inruet in arcum aereum
JOB|20|25|eductus et egrediens de vagina sua et fulgurans in amaritudine sua vadent et venient super eum horribiles
JOB|20|26|omnes tenebrae absconditae sunt in occultis eius devorabit eum ignis qui non succenditur adfligetur relictus in tabernaculo suo
JOB|20|27|revelabunt caeli iniquitatem eius et terra consurget adversus eum
JOB|20|28|apertum erit germen domus illius detrahetur in die furoris Dei
JOB|20|29|haec est pars hominis impii a Deo et hereditas verborum eius a Domino
JOB|21|1|respondens autem Iob dixit
JOB|21|2|audite quaeso sermones meos et agetis paenitentiam
JOB|21|3|sustinete me ut et ego loquar et post mea si videbitur verba ridete
JOB|21|4|numquid contra hominem disputatio mea est ut merito non debeam contristari
JOB|21|5|adtendite me et obstupescite et superponite digitum ori vestro
JOB|21|6|et ego quando recordatus fuero pertimesco et concutit carnem meam tremor
JOB|21|7|quare ergo impii vivunt sublevati sunt confortatique divitiis
JOB|21|8|semen eorum permanet coram eis propinquorum turba et nepotum in conspectu eorum
JOB|21|9|domus eorum securae sunt et pacatae et non est virga Dei super illos
JOB|21|10|bos eorum concepit et non abortit vacca peperit et non est privata fetu suo
JOB|21|11|egrediuntur quasi greges parvuli eorum et infantes eorum exultant lusibus
JOB|21|12|tenent tympanum et citharam et gaudent ad sonitum organi
JOB|21|13|ducunt in bonis dies suos et in puncto ad inferna descendunt
JOB|21|14|qui dixerunt Deo recede a nobis et scientiam viarum tuarum nolumus
JOB|21|15|quid est Omnipotens ut serviamus ei et quid nobis prodest si oraverimus illum
JOB|21|16|verumtamen quia non sunt in manu eorum bona sua consilium impiorum longe sit a me
JOB|21|17|quotiens lucerna impiorum extinguetur et superveniet eis inundatio et dolores dividet furoris sui
JOB|21|18|erunt sicut paleae ante faciem venti et sicut favilla quam turbo dispergit
JOB|21|19|Deus servabit filiis illius dolorem patris et cum reddiderit tunc sciet
JOB|21|20|videbunt oculi eius interfectionem suam et de furore Omnipotentis bibet
JOB|21|21|quid enim ad eum pertinet de domo sua post se et si numerus mensuum eius dimidietur
JOB|21|22|numquid Deum quispiam docebit scientiam qui excelsos iudicat
JOB|21|23|iste moritur robustus et sanus dives et felix
JOB|21|24|viscera eius plena sunt adipe et medullis ossa illius inrigantur
JOB|21|25|alius vero moritur in amaritudine animae absque ullis opibus
JOB|21|26|et tamen simul in pulverem dormient et vermes operient eos
JOB|21|27|certe novi cogitationes vestras et sententias contra me iniquas
JOB|21|28|dicitis enim ubi est domus principis et ubi tabernacula impiorum
JOB|21|29|interrogate quemlibet de viatoribus et haec eadem eum intellegere cognoscetis
JOB|21|30|quia in diem perditionis servabitur malus et ad diem furoris ducitur
JOB|21|31|quis arguet coram eo viam eius et quae fecit quis reddet illi
JOB|21|32|ipse ad sepulchra ducetur et in congerie mortuorum vigilabit
JOB|21|33|dulcis fuit glareis Cocyti et post se omnem hominem trahet et ante se innumerabiles
JOB|21|34|quomodo igitur consolamini me frustra cum responsio vestra repugnare ostensa sit veritati
JOB|22|1|respondens autem Eliphaz Themanites dixit
JOB|22|2|numquid Deo conparari potest homo etiam cum perfectae fuerit scientiae
JOB|22|3|quid prodest Deo si iustus fueris aut quid ei confers si inmaculata fuerit via tua
JOB|22|4|numquid timens arguet te et veniet tecum in iudicium
JOB|22|5|et non propter malitiam tuam plurimam et infinitas iniquitates tuas
JOB|22|6|abstulisti enim pignus fratrum tuorum sine causa et nudos spoliasti vestibus
JOB|22|7|aquam lasso non dedisti et esurienti subtraxisti panem
JOB|22|8|in fortitudine brachii tui possidebas terram et potentissimus obtinebas eam
JOB|22|9|viduas dimisisti vacuas et lacertos pupillorum comminuisti
JOB|22|10|propterea circumdatus es laqueis et conturbat te formido subita
JOB|22|11|et putabas te tenebras non visurum et impetu aquarum inundantium non oppressurum
JOB|22|12|an cogitas quod Deus excelsior caelo et super stellarum vertices sublimetur
JOB|22|13|et dicis quid enim novit Deus et quasi per caliginem iudicat
JOB|22|14|nubes latibulum eius nec nostra considerat et circa cardines caeli perambulat
JOB|22|15|numquid semitam saeculorum custodire cupis quam calcaverunt viri iniqui
JOB|22|16|qui sublati sunt ante tempus suum et fluvius subvertit fundamentum eorum
JOB|22|17|qui dicebant Deo recede a nobis et quasi nihil possit facere Omnipotens aestimabant eum
JOB|22|18|cum ille implesset domos eorum bonis quorum sententia procul sit a me
JOB|22|19|videbunt iusti et laetabuntur et innocens subsannabit eos
JOB|22|20|nonne succisa est erectio eorum et reliquias eorum devoravit ignis
JOB|22|21|adquiesce igitur ei et habeto pacem et per haec habebis fructus optimos
JOB|22|22|suscipe ex ore illius legem et pone sermones eius in corde tuo
JOB|22|23|si reversus fueris ad Omnipotentem aedificaberis et longe facies iniquitatem a tabernaculo tuo
JOB|22|24|dabit pro terra silicem et pro silice torrentes aureos
JOB|22|25|eritque Omnipotens contra hostes tuos et argentum coacervabitur tibi
JOB|22|26|tunc super Omnipotentem deliciis afflues et elevabis ad Deum faciem tuam
JOB|22|27|rogabis eum et exaudiet te et vota tua reddes
JOB|22|28|decernes rem et veniet tibi et in viis tuis splendebit lumen
JOB|22|29|qui enim humiliatus fuerit erit in gloria et qui inclinaverit oculos suos ipse salvabitur
JOB|22|30|salvabitur innocens salvabitur autem munditia manuum suarum
JOB|23|1|respondens autem Iob dixit
JOB|23|2|nunc quoque in amaritudine est sermo meus et manus plagae meae adgravata est super gemitum meum
JOB|23|3|quis mihi tribuat ut cognoscam et inveniam illum et veniam usque ad solium eius
JOB|23|4|ponam coram eo iudicium et os meum replebo increpationibus
JOB|23|5|ut sciam verba quae mihi respondeat et intellegam quid loquatur mihi
JOB|23|6|nolo multa fortitudine contendat mecum nec magnitudinis suae mole me premat
JOB|23|7|proponat aequitatem contra me et perveniat ad victoriam iudicium meum
JOB|23|8|si ad orientem iero non apparet si ad occidentem non intellegam eum
JOB|23|9|si ad sinistram quid agat non adprehendam eum si me vertam ad dextram non videbo illum
JOB|23|10|ipse vero scit viam meam et probavit me quasi aurum quod per ignem transit
JOB|23|11|vestigia eius secutus est pes meus viam eius custodivi et non declinavi ex ea
JOB|23|12|a mandatis labiorum eius non recessi et in sinu meo abscondi verba oris eius
JOB|23|13|ipse enim solus est et nemo avertere potest cogitationem eius et anima eius quodcumque voluerit hoc facit
JOB|23|14|cum expleverit in me voluntatem suam et alia multa similia praesto sunt ei
JOB|23|15|et idcirco a facie eius turbatus sum et considerans eum timore sollicitor
JOB|23|16|Deus mollivit cor meum et Omnipotens conturbavit me
JOB|23|17|non enim perii propter inminentes tenebras nec faciem meam operuit caligo
JOB|24|1|ab Omnipotente non sunt abscondita tempora qui autem noverunt eum ignorant dies illius
JOB|24|2|alii terminos transtulerunt diripuerunt greges et paverunt eos
JOB|24|3|asinum pupillorum abigerunt et abstulerunt pro pignore bovem viduae
JOB|24|4|subverterunt pauperum viam et oppresserunt pariter mansuetos terrae
JOB|24|5|alii quasi onagri in deserto egrediuntur ad opus suum vigilantesque ad praedam praeparant panem liberis
JOB|24|6|agrum non suum demetunt et vineam eius quem vi oppresserunt vindemiant
JOB|24|7|nudos dimittunt homines indumenta tollentes quibus non est operimentum in frigore
JOB|24|8|quos imbres montium rigant et non habentes velamen amplexantur lapides
JOB|24|9|vim fecerunt depraedantes pupillos et vulgum pauperem spoliaverunt
JOB|24|10|nudis et incedentibus absque vestitu et esurientibus tulerunt spicas
JOB|24|11|inter acervos eorum meridiati sunt qui calcatis torcularibus sitiunt
JOB|24|12|de civitatibus fecerunt viros gemere et anima vulneratorum clamavit et Deus inultum abire non patitur
JOB|24|13|ipsi fuerunt rebelles luminis nescierunt vias eius nec reversi sunt per semitas illius
JOB|24|14|mane primo consurgit homicida interficit egenum et pauperem per noctem vero erit quasi fur
JOB|24|15|oculus adulteri observat caliginem dicens non me videbit oculus et operiet vultum suum
JOB|24|16|perfodit in tenebris domos sicut in die condixerant sibi et ignoraverunt lucem
JOB|24|17|si subito apparuerit aurora arbitrantur umbram mortis et sic in tenebris quasi in luce ambulant
JOB|24|18|levis est super faciem aquae maledicta sit pars eius in terra nec ambulet per viam vinearum
JOB|24|19|ad nimium calorem transeat ab aquis nivium et usque ad inferos peccatum illius
JOB|24|20|obliviscatur eius misericordia dulcedo illius vermes non sit in recordatione sed conteratur quasi lignum infructuosum
JOB|24|21|pavit enim sterilem et quae non parit et viduae bene non fecit
JOB|24|22|detraxit fortes in fortitudine sua et cum steterit non credet vitae suae
JOB|24|23|dedit ei Deus locum paenitentiae et ille abutitur eo in superbiam oculi autem eius sunt in viis illius
JOB|24|24|elevati sunt ad modicum et non subsistent et humiliabuntur sicut omnia et auferentur et sicut summitates spicarum conterentur
JOB|24|25|quod si non est ita quis me potest arguere esse mentitum et ponere ante Deum verba mea
JOB|25|1|respondens autem Baldad Suites dixit
JOB|25|2|potestas et terror apud eum est qui facit concordiam in sublimibus suis
JOB|25|3|numquid est numerus militum eius et super quem non surget lumen illius
JOB|25|4|numquid iustificari potest homo conparatus Deo aut apparere mundus natus de muliere
JOB|25|5|ecce etiam luna non splendet et stellae non sunt mundae in conspectu eius
JOB|25|6|quanto magis homo putredo et filius hominis vermis
JOB|26|1|respondens autem Iob dixit
JOB|26|2|cuius adiutor es numquid inbecilli et sustentas brachium eius qui non est fortis
JOB|26|3|cui dedisti consilium forsitan illi qui non habet sapientiam et prudentiam tuam ostendisti plurimam
JOB|26|4|quem docere voluisti nonne eum qui fecit spiramen tuum
JOB|26|5|ecce gigantes gemunt sub aquis et qui habitant cum eis
JOB|26|6|nudus est inferus coram illo et nullum est operimentum perditioni
JOB|26|7|qui extendit aquilonem super vacuum et adpendit terram super nihili
JOB|26|8|qui ligat aquas in nubibus suis ut non erumpant pariter deorsum
JOB|26|9|qui tenet vultum solii sui et expandit super illud nebulam suam
JOB|26|10|terminum circumdedit aquis usque dum finiantur lux et tenebrae
JOB|26|11|columnae caeli contremescunt et pavent ad nutum eius
JOB|26|12|in fortitudine illius repente maria congregata sunt et prudentia eius percussit superbum
JOB|26|13|spiritus eius ornavit caelos et obsetricante manu eius eductus est coluber tortuosus
JOB|26|14|ecce haec ex parte dicta sunt viarum eius et cum vix parvam stillam sermonis eius audierimus quis poterit tonitruum magnitudinis illius intueri
JOB|27|1|addidit quoque Iob adsumens parabolam suam et dixit
JOB|27|2|vivit Deus qui abstulit iudicium meum et Omnipotens qui ad amaritudinem adduxit animam meam
JOB|27|3|quia donec superest halitus in me et spiritus Dei in naribus meis
JOB|27|4|non loquentur labia mea iniquitatem nec lingua mea meditabitur mendacium
JOB|27|5|absit a me ut iustos vos esse iudicem donec deficiam non recedam ab innocentia mea
JOB|27|6|iustificationem meam quam coepi tenere non deseram nec enim reprehendit me cor meum in omni vita mea
JOB|27|7|sit ut impius inimicus meus et adversarius meus quasi iniquus
JOB|27|8|quae enim spes est hypocritae si avare rapiat et non liberet Deus animam eius
JOB|27|9|numquid clamorem eius Deus audiet cum venerit super illum angustia
JOB|27|10|aut poterit in Omnipotente delectari et invocare Deum in omni tempore
JOB|27|11|docebo vos per manum Dei quae Omnipotens habeat nec abscondam
JOB|27|12|ecce vos omnes nostis et quid sine causa vana loquimini
JOB|27|13|haec est pars hominis impii apud Deum et hereditas violentorum quam ab Omnipotente suscipient
JOB|27|14|si multiplicati fuerint filii eius in gladio erunt et nepotes eius non saturabuntur pane
JOB|27|15|qui reliqui fuerint ex eo sepelientur in interitu et viduae illius non plorabunt
JOB|27|16|si conportaverit quasi terram argentum et sicut lutum praeparaverit vestimenta
JOB|27|17|praeparabit quidem sed iustus vestietur illis et argentum innocens dividet
JOB|27|18|aedificavit sicut tinea domum suam et sicut custos fecit umbraculum
JOB|27|19|dives cum dormierit nihil secum auferet aperit oculos suos et nihil inveniet
JOB|27|20|adprehendit eum quasi aqua inopia nocte opprimet eum tempestas
JOB|27|21|tollet eum ventus urens et auferet et velut turbo rapiet eum de loco suo
JOB|27|22|et mittet super eum et non parcet de manu eius fugiens fugiet
JOB|27|23|stringet super eum manus suas et sibilabit super illum intuens locum eius
JOB|28|1|habet argentum venarum suarum principia et auro locus est in quo conflatur
JOB|28|2|ferrum de terra tollitur et lapis solutus calore in aes vertitur
JOB|28|3|tempus posuit tenebris et universorum finem ipse considerat lapidem quoque caliginis et umbram mortis
JOB|28|4|dividit torrens a populo peregrinante eos quos oblitus est pes egentis hominum et invios
JOB|28|5|terra de qua oriebatur panis in loco suo igne subversa est
JOB|28|6|locus sapphyri lapides eius et glebae illius aurum
JOB|28|7|semitam ignoravit avis nec intuitus est oculus vulturis
JOB|28|8|non calcaverunt eam filii institorum nec pertransivit per eam leaena
JOB|28|9|ad silicem extendit manum suam subvertit a radicibus montes
JOB|28|10|in petris rivos excidit et omne pretiosum vidit oculus eius
JOB|28|11|profunda quoque fluviorum scrutatus est et abscondita produxit in lucem
JOB|28|12|sapientia vero ubi invenitur et quis est locus intellegentiae
JOB|28|13|nescit homo pretium eius nec invenitur in terra suaviter viventium
JOB|28|14|abyssus dicit non est in me et mare loquitur non est mecum
JOB|28|15|non dabitur aurum obrizum pro ea nec adpendetur argentum in commutatione eius
JOB|28|16|non conferetur tinctis Indiae coloribus nec lapidi sardonico pretiosissimo vel sapphyro
JOB|28|17|non adaequabitur ei aurum vel vitrum nec commutabuntur pro ea vasa auri
JOB|28|18|excelsa et eminentia non memorabuntur conparatione eius trahitur autem sapientia de occultis
JOB|28|19|non adaequabitur ei topazium de Aethiopia nec tincturae mundissimae conponetur
JOB|28|20|unde ergo sapientia veniet et quis est locus intellegentiae
JOB|28|21|abscondita est ab oculis omnium viventium volucres quoque caeli latet
JOB|28|22|perditio et mors dixerunt auribus nostris audivimus famam eius
JOB|28|23|Deus intellegit viam eius et ipse novit locum illius
JOB|28|24|ipse enim fines mundi intuetur et omnia quae sub caelo sunt respicit
JOB|28|25|qui fecit ventis pondus et aquas adpendit mensura
JOB|28|26|quando ponebat pluviis legem et viam procellis sonantibus
JOB|28|27|tunc vidit illam et enarravit et praeparavit et investigavit
JOB|28|28|et dixit homini ecce timor Domini ipsa est sapientia et recedere a malo intellegentia
JOB|29|1|addidit quoque Iob adsumens parabolam suam et dixit
JOB|29|2|quis mihi tribuat ut sim iuxta menses pristinos secundum dies quibus Deus custodiebat me
JOB|29|3|quando splendebat lucerna eius super caput meum et ad lumen eius ambulabam in tenebris
JOB|29|4|sicut fui in diebus adulescentiae meae quando secreto Deus erat in tabernaculo meo
JOB|29|5|quando erat Omnipotens mecum et in circuitu meo pueri mei
JOB|29|6|quando lavabam pedes meos butyro et petra fundebat mihi rivos olei
JOB|29|7|quando procedebam ad portam civitatis et in platea parabant cathedram mihi
JOB|29|8|videbant me iuvenes et abscondebantur et senes adsurgentes stabant
JOB|29|9|principes cessabant loqui et digitum superponebant ori suo
JOB|29|10|vocem suam cohibebant duces et lingua eorum gutturi suo adherebat
JOB|29|11|auris audiens beatificabat me et oculus videns testimonium reddebat mihi
JOB|29|12|quod liberassem pauperem vociferantem et pupillum cui non esset adiutor
JOB|29|13|benedictio perituri super me veniebat et cor viduae consolatus sum
JOB|29|14|iustitia indutus sum et vestivit me sicut vestimento et diademate iudicio meo
JOB|29|15|oculus fui caeco et pes claudo
JOB|29|16|pater eram pauperum et causam quam nesciebam diligentissime investigabam
JOB|29|17|conterebam molas iniqui et de dentibus illius auferebam praedam
JOB|29|18|dicebamque in nidulo meo moriar et sicut palma multiplicabo dies
JOB|29|19|radix mea aperta est secus aquas et ros morabitur in messione mea
JOB|29|20|gloria mea semper innovabitur et arcus meus in manu mea instaurabitur
JOB|29|21|qui me audiebant expectabant sententiam et intenti tacebant ad consilium meum
JOB|29|22|verbis meis addere nihil audebant et super illos stillabat eloquium meum
JOB|29|23|expectabant me sicut pluviam et os suum aperiebant quasi ad imbrem serotinum
JOB|29|24|si quando ridebam ad eos non credebant et lux vultus mei non cadebat in terram
JOB|29|25|si voluissem ire ad eos sedebam primus cumque sederem quasi rex circumstante exercitu eram tamen maerentium consolator
JOB|30|1|nunc autem derident me iuniores tempore quorum non dignabar patres ponere cum canibus gregis mei
JOB|30|2|quorum virtus manuum erat mihi pro nihilo et vita ipsa putabantur indigni
JOB|30|3|egestate et fame steriles qui rodebant in solitudine squalentes calamitate et miseria
JOB|30|4|et mandebant herbas et arborum cortices et radix iuniperorum erat cibus eorum
JOB|30|5|qui de convallibus ista rapientes cum singula repperissent ad ea cum clamore currebant
JOB|30|6|in desertis habitabant torrentium et in cavernis terrae vel super glaream
JOB|30|7|qui inter huiuscemodi laetabantur et esse sub sentibus delicias conputabant
JOB|30|8|filii stultorum et ignobilium et in terra penitus non parentes
JOB|30|9|nunc in eorum canticum versus sum et factus sum eis proverbium
JOB|30|10|abominantur me et longe fugiunt a me et faciem meam conspuere non verentur
JOB|30|11|faretram enim suam aperuit et adflixit me et frenum posuit in os meum
JOB|30|12|ad dexteram orientis calamitatis meae ilico surrexerunt pedes meos subverterunt et oppresserunt quasi fluctibus semitis suis
JOB|30|13|dissipaverunt itinera mea insidiati sunt mihi et praevaluerunt et non fuit qui ferret auxilium
JOB|30|14|quasi rupto muro et aperta ianua inruerunt super me et ad meas miserias devoluti sunt
JOB|30|15|redactus sum in nihili abstulisti quasi ventus desiderium meum et velut nubes pertransiit salus mea
JOB|30|16|nunc autem in memet ipso marcescit anima mea et possident me dies adflictionis
JOB|30|17|nocte os meum perforatur doloribus et qui me comedunt non dormiunt
JOB|30|18|in multitudine eorum consumitur vestimentum meum et quasi capitio tunicae sic cinxerunt me
JOB|30|19|conparatus sum luto et adsimilatus favillae et cineri
JOB|30|20|clamo ad te et non exaudis me sto et non respicis me
JOB|30|21|mutatus es mihi in crudelem et in duritia manus tuae adversaris mihi
JOB|30|22|elevasti me et quasi super ventum ponens elisisti me valide
JOB|30|23|scio quia morti tradas me ubi constituta domus est omni viventi
JOB|30|24|verumtamen non ad consumptionem eorum emittis manum tuam et si corruerint ipse salvabis
JOB|30|25|flebam quondam super eum qui adflictus erat et conpatiebatur anima mea pauperi
JOB|30|26|expectabam bona et venerunt mihi mala praestolabar lucem et eruperunt tenebrae
JOB|30|27|interiora mea efferbuerunt absque ulla requie praevenerunt me dies adflictionis
JOB|30|28|maerens incedebam sine furore consurgens in turba clamavi
JOB|30|29|frater fui draconum et socius strutionum
JOB|30|30|cutis mea denigrata est super me et ossa mea aruerunt prae caumate
JOB|30|31|versa est in luctum cithara mea et organum meum in vocem flentium
JOB|31|1|pepigi foedus cum oculis meis ut ne cogitarem quidem de virgine
JOB|31|2|quam enim partem haberet Deus in me desuper et hereditatem Omnipotens de excelsis
JOB|31|3|numquid non perditio est iniquo et alienatio operantibus iniustitiam
JOB|31|4|nonne ipse considerat vias meas et cunctos gressus meos dinumerat
JOB|31|5|si ambulavi in vanitate et festinavit in dolo pes meus
JOB|31|6|adpendat me in statera iusta et sciat Deus simplicitatem meam
JOB|31|7|si declinavit gressus meus de via et si secutum est oculos meos cor meum et in manibus meis adhesit macula
JOB|31|8|seram et alius comedat et progenies mea eradicetur
JOB|31|9|si deceptum est cor meum super mulierem et si ad ostium amici mei insidiatus sum
JOB|31|10|scortum sit alteri uxor mea et super illam incurventur alii
JOB|31|11|hoc enim nefas est et iniquitas maxima
JOB|31|12|ignis est usque ad perditionem devorans et omnia eradicans genimina
JOB|31|13|si contempsi subire iudicium cum servo meo et ancillae meae cum disceptarent adversum me
JOB|31|14|quid enim faciam cum surrexerit ad iudicandum Deus et cum quaesierit quid respondebo illi
JOB|31|15|numquid non in utero fecit me qui et illum operatus est et formavit in vulva unus
JOB|31|16|si negavi quod volebant pauperibus et oculos viduae expectare feci
JOB|31|17|si comedi buccellam meam solus et non comedit pupillus ex ea
JOB|31|18|quia ab infantia mea crevit mecum miseratio et de utero matris meae egressa est mecum
JOB|31|19|si despexi pereuntem eo quod non habuerit indumentum et absque operimento pauperem
JOB|31|20|si non benedixerunt mihi latera eius et de velleribus ovium mearum calefactus est
JOB|31|21|si levavi super pupillum manum meam etiam cum viderem me in porta superiorem
JOB|31|22|umerus meus a iunctura sua cadat et brachium meum cum suis ossibus confringatur
JOB|31|23|semper enim quasi tumentes super me fluctus timui Deum et pondus eius ferre non potui
JOB|31|24|si putavi aurum robur meum et obrizae dixi fiducia mea
JOB|31|25|si laetatus sum super multis divitiis meis et quia plurima repperit manus mea
JOB|31|26|si vidi solem cum fulgeret et lunam incedentem clare
JOB|31|27|et lactatum est in abscondito cor meum et osculatus sum manum meam ore meo
JOB|31|28|quae est iniquitas maxima et negatio contra Deum altissimum
JOB|31|29|si gavisus sum ad ruinam eius qui me oderat et exultavi quod invenisset eum malum
JOB|31|30|non enim dedi ad peccandum guttur meum ut expeterem maledicens animam eius
JOB|31|31|si non dixerunt viri tabernaculi mei quis det de carnibus eius ut saturemur
JOB|31|32|foris non mansit peregrinus ostium meum viatori patuit
JOB|31|33|si abscondi quasi homo peccatum meum et celavi in sinu meo iniquitatem meam
JOB|31|34|si expavi ad multitudinem nimiam et despectio propinquorum terruit me et non magis tacui nec egressus sum ostium
JOB|31|35|quis mihi tribuat auditorem ut desiderium meum Omnipotens audiat et librum scribat ipse qui iudicat
JOB|31|36|ut in umero meo portem illum et circumdem illum quasi coronam mihi
JOB|31|37|per singulos gradus meos pronuntiabo illum et quasi principi offeram eum
JOB|31|38|si adversum me terra mea clamat et cum ipsa sulci eius deflent
JOB|31|39|si fructus eius comedi absque pecunia et animam agricolarum eius adflixi
JOB|31|40|pro frumento oriatur mihi tribulus et pro hordeo spina finita sunt verba Iob
JOB|32|1|omiserunt autem tres viri isti respondere Iob eo quod iustus sibi videretur
JOB|32|2|et iratus indignatusque Heliu filius Barachel Buzites de cognatione Ram iratus est autem adversus Iob eo quod iustum se esse diceret coram Deo
JOB|32|3|porro adversum amicos eius indignatus est eo quod non invenissent responsionem rationabilem sed tantummodo condemnassent Iob
JOB|32|4|igitur Heliu expectavit Iob loquentem eo quod seniores se essent qui loquebantur
JOB|32|5|cum autem vidisset quod tres respondere non potuissent iratus est vehementer
JOB|32|6|respondensque Heliu filius Barachel Buzites dixit iunior sum tempore vos autem antiquiores idcirco dimisso capite veritus sum indicare vobis meam sententiam
JOB|32|7|sperabam enim quod aetas prolixior loqueretur et annorum multitudo doceret sapientiam
JOB|32|8|sed ut video spiritus est in hominibus et inspiratio Omnipotentis dat intellegentiam
JOB|32|9|non sunt longevi sapientes nec senes intellegunt iudicium
JOB|32|10|ideo dicam audite me ostendam vobis etiam ego meam scientiam
JOB|32|11|expectavi enim sermones vestros audivi prudentiam vestram donec disceptaremini sermonibus
JOB|32|12|et donec putabam vos aliquid dicere considerabam sed ut video non est qui arguere possit Iob et respondere ex vobis sermonibus eius
JOB|32|13|ne forte dicatis invenimus sapientiam Deus proiecit eum non homo
JOB|32|14|nihil locutus est mihi et ego non secundum vestros sermones respondebo illi
JOB|32|15|extimuerunt non responderunt ultra abstuleruntque a se eloquia
JOB|32|16|quoniam igitur expectavi et non sunt locuti steterunt nec responderunt ultra
JOB|32|17|respondebo et ego partem meam et ostendam scientiam meam
JOB|32|18|plenus sum enim sermonibus et coartat me spiritus uteri mei
JOB|32|19|en venter meus quasi mustum absque spiraculo quod lagunculas novas disrumpit
JOB|32|20|loquar et respirabo paululum aperiam labia mea et respondebo
JOB|32|21|non accipiam personam viri et Deum homini non aequabo
JOB|32|22|nescio enim quamdiu subsistam et si post modicum tollat me factor meus
JOB|33|1|audi igitur Iob eloquia mea et omnes sermones meos ausculta
JOB|33|2|ecce aperui os meum loquatur lingua mea in faucibus meis
JOB|33|3|simplici corde meo sermones mei et sententiam labia mea puram loquentur
JOB|33|4|spiritus Dei fecit me et spiraculum Omnipotentis vivificavit me
JOB|33|5|si potes responde mihi et adversus faciem meam consiste
JOB|33|6|ecce et me sicut et te fecit Deus et de eodem luto ego quoque formatus sum
JOB|33|7|verumtamen miraculum meum non te terreat et eloquentia mea non sit tibi gravis
JOB|33|8|dixisti ergo in auribus meis et vocem verborum audivi
JOB|33|9|mundus sum ego absque delicto inmaculatus et non est iniquitas in me
JOB|33|10|quia querellas in me repperit ideo arbitratus est me inimicum sibi
JOB|33|11|posuit in nervo pedes meos custodivit omnes semitas meas
JOB|33|12|hoc est ergo in quo non es iustificatus respondebo tibi quia maior sit Deus homine
JOB|33|13|adversum eum contendis quod non ad omnia verba responderit tibi
JOB|33|14|semel loquitur Deus et secundo id ipsum non repetit
JOB|33|15|per somnium in visione nocturna quando inruit sopor super homines et dormiunt in lectulo
JOB|33|16|tunc aperit aures virorum et erudiens eos instruit disciplinam
JOB|33|17|ut avertat hominem ab his quae facit et liberet eum de superbia
JOB|33|18|eruens animam eius a corruptione et vitam illius ut non transeat in gladium
JOB|33|19|increpat quoque per dolorem in lectulo et omnia ossa eius marcescere facit
JOB|33|20|abominabilis ei fit in vita sua panis et animae illius cibus ante desiderabilis
JOB|33|21|tabescet caro eius et ossa quae tecta fuerant nudabuntur
JOB|33|22|adpropinquabit corruptioni anima eius et vita illius mortiferis
JOB|33|23|si fuerit pro eo angelus loquens unum de milibus ut adnuntiet hominis aequitatem
JOB|33|24|miserebitur eius et dicet libera eum et non descendat in corruptionem inveni in quo ei propitier
JOB|33|25|consumpta est caro eius a suppliciis revertatur ad dies adulescentiae suae
JOB|33|26|deprecabitur Deum et placabilis ei erit et videbit faciem eius in iubilo et reddet homini iustitiam suam
JOB|33|27|respiciet homines et dicet peccavi et vere deliqui et ut eram dignus non recepi
JOB|33|28|liberavit animam suam ne pergeret in interitum sed vivens lucem videret
JOB|33|29|ecce haec omnia operatur Deus tribus vicibus per singulos
JOB|33|30|ut revocet animas eorum a corruptione et inluminet luce viventium
JOB|33|31|adtende Iob et audi me et tace dum ego loquar
JOB|33|32|si autem habes quod loquaris responde mihi loquere volo enim te apparere iustum
JOB|33|33|quod si non habes audi me tace et docebo te sapientiam
JOB|34|1|pronuntians itaque Heliu etiam haec locutus est
JOB|34|2|audite sapientes verba mea et eruditi auscultate me
JOB|34|3|auris enim verba probat et guttur escas gustu diiudicat
JOB|34|4|iudicium eligamus nobis et inter nos videamus quid sit melius
JOB|34|5|quia dixit Iob iustus sum et Deus subvertit iudicium meum
JOB|34|6|in iudicando enim me mendacium est violenta sagitta mea absque ullo peccato
JOB|34|7|quis est vir ut est Iob qui bibit subsannationem quasi aquam
JOB|34|8|qui graditur cum operantibus iniquitatem et ambulat cum viris impiis
JOB|34|9|dixit enim non placebit vir Deo etiam si cucurrerit cum eo
JOB|34|10|ideo viri cordati audite me absit a Deo impietas et ab Omnipotente iniquitas
JOB|34|11|opus enim hominis reddet ei et iuxta vias singulorum restituet
JOB|34|12|vere enim Deus non condemnabit frustra nec Omnipotens subvertet iudicium
JOB|34|13|quem constituit alium super terram aut quem posuit super orbem quem fabricatus est
JOB|34|14|si direxerit ad eum cor suum spiritum illius et flatum ad se trahet
JOB|34|15|deficiet omnis caro simul et homo in cinerem revertetur
JOB|34|16|si habes ergo intellectum audi quod dicitur et ausculta vocem eloquii mei
JOB|34|17|numquid qui non amat iudicium sanare potest et quomodo tu eum qui iustus est in tantum condemnas
JOB|34|18|qui dicit regi apostata qui vocat duces impios
JOB|34|19|qui non accipit personas principum nec cognovit tyrannum cum disceptaret contra pauperem opus enim manuum eius sunt universi
JOB|34|20|subito morientur et in media nocte turbabuntur populi et pertransibunt et auferent violentum absque manu
JOB|34|21|oculi enim eius super vias hominum et omnes gressus eorum considerat
JOB|34|22|non sunt tenebrae et non est umbra mortis ut abscondantur ibi qui operantur iniquitatem
JOB|34|23|neque enim ultra in hominis potestate est ut veniat ad Deum in iudicium
JOB|34|24|conteret multos innumerabiles et stare faciet alios pro eis
JOB|34|25|novit enim opera eorum et idcirco inducet noctem et conterentur
JOB|34|26|quasi impios percussit eos in loco videntium
JOB|34|27|qui quasi de industria recesserunt ab eo et omnes vias eius intellegere noluerunt
JOB|34|28|ut pervenire facerent ad eum clamorem egeni et audiret vocem pauperum
JOB|34|29|ipso enim concedente pacem quis est qui condemnet ex quo absconderit vultum quis est qui contempletur eum et super gentem et super omnes homines
JOB|34|30|qui regnare facit hominem hypocritam propter peccata populi
JOB|34|31|quia ergo ego locutus sum ad Deum te quoque non prohibeo
JOB|34|32|si erravi tu doce me si iniquitatem locutus sum ultra non addam
JOB|34|33|numquid a te Deus expetit eam quia displicuit tibi tu enim coepisti loqui et non ego quod si quid nosti melius loquere
JOB|34|34|viri intellegentes loquantur mihi et vir sapiens audiat me
JOB|34|35|Iob autem stulte locutus est et verba illius non sonant disciplinam
JOB|34|36|pater mi probetur Iob usque ad finem ne desinas in hominibus iniquitatis
JOB|34|37|quia addit super peccata sua blasphemiam inter nos interim constringatur et tunc ad iudicium provocet sermonibus suis Deum
JOB|35|1|igitur Heliu haec rursum locutus est
JOB|35|2|numquid aequa tibi videtur tua cogitatio ut diceres iustior Deo sum
JOB|35|3|dixisti enim non tibi placet quod rectum est vel quid tibi proderit si ego peccavero
JOB|35|4|itaque ego respondebo sermonibus tuis et amicis tuis tecum
JOB|35|5|suspice caelum et intuere et contemplare aethera quod altior te sit
JOB|35|6|si peccaveris quid ei nocebis et si multiplicatae fuerint iniquitates tuae quid facies contra eum
JOB|35|7|porro si iuste egeris quid donabis ei aut quid de manu tua accipiet
JOB|35|8|homini qui similis tui est nocebit impietas tua et filium hominis adiuvabit iustitia tua
JOB|35|9|propter multitudinem calumniatorum clamabunt et heiulabunt propter vim brachii tyrannorum
JOB|35|10|et non dixit ubi est Deus qui fecit me qui dedit carmina in nocte
JOB|35|11|qui docet nos super iumenta terrae et super volucres caeli erudit nos
JOB|35|12|ibi clamabunt et non exaudiet propter superbiam malorum
JOB|35|13|non ergo frustra audiet Deus et Omnipotens singulorum causas intuebitur
JOB|35|14|etiam cum dixeris non considerat iudicare coram eo et expecta eum
JOB|35|15|nunc enim non infert furorem suum nec ulciscitur scelus valde
JOB|35|16|ergo Iob frustra aperit os suum et absque scientia verba multiplicat
JOB|36|1|addens quoque Heliu haec locutus est
JOB|36|2|sustine me paululum et indicabo tibi adhuc enim habeo quod pro Deo loquar
JOB|36|3|repetam scientiam meam a principio et operatorem meum probabo iustum
JOB|36|4|vere enim absque mendacio sermones mei et perfecta scientia probabitur tibi
JOB|36|5|Deus potentes non abicit cum et ipse sit potens
JOB|36|6|sed non salvat impios et iudicium pauperibus tribuit
JOB|36|7|non aufert a iusto oculos suos et reges in solio conlocat in perpetuum et illi eriguntur
JOB|36|8|et si fuerint in catenis et vinciantur funibus paupertatis
JOB|36|9|indicabit eis opera eorum et scelera eorum quia violenti fuerint
JOB|36|10|revelabit quoque aurem eorum ut corripiat et loquetur ut revertantur ab iniquitate
JOB|36|11|si audierint et observaverint conplebunt dies suos in bono et annos suos in gloria
JOB|36|12|si autem non audierint transibunt per gladium et consumentur in stultitia
JOB|36|13|simulatores et callidi provocant iram Dei neque clamabunt cum vincti fuerint
JOB|36|14|morietur in tempestate anima eorum et vita eorum inter effeminatos
JOB|36|15|eripiet pauperem de angustia sua et revelabit in tribulatione aurem eius
JOB|36|16|igitur salvabit te de ore angusto latissime et non habentis fundamentum subter se requies autem mensae tuae erit plena pinguedine
JOB|36|17|causa tua quasi impii iudicata est causam iudiciumque recipies
JOB|36|18|non te ergo superet ira ut aliquem opprimas nec multitudo donorum inclinet te
JOB|36|19|depone magnitudinem tuam absque tribulatione et omnes robustos fortitudine
JOB|36|20|ne protrahas noctem ut ascendant populi pro eis
JOB|36|21|cave ne declines ad iniquitatem hanc enim coepisti sequi post miseriam
JOB|36|22|ecce Deus excelsus in fortitudine sua et nullus ei similis in legislatoribus
JOB|36|23|quis poterit scrutari vias eius aut quis ei dicere operatus es iniquitatem
JOB|36|24|memento quod ignores opus eius de quo cecinerunt viri
JOB|36|25|omnes homines vident eum unusquisque intuetur procul
JOB|36|26|ecce Deus magnus vincens scientiam nostram numerus annorum eius inaestimabilis
JOB|36|27|qui aufert stillas pluviae et effundit imbres ad instar gurgitum
JOB|36|28|qui de nubibus fluunt quae praetexunt cuncta desuper
JOB|36|29|si voluerit extendere nubes quasi tentorium suum
JOB|36|30|et fulgurare lumine suo desuper cardines quoque maris operiet
JOB|36|31|per haec enim iudicat populos et dat escas multis mortalibus
JOB|36|32|in manibus abscondit lucem et praecipit ei ut rursus adveniat
JOB|36|33|adnuntiat de ea amico suo quod possessio eius sit et ad eam possit ascendere
JOB|37|1|super hoc expavit cor meum et emotum est de loco suo
JOB|37|2|audite auditionem in terrore vocis eius et sonum de ore illius procedentem
JOB|37|3|subter omnes caelos ipse considerat et lumen illius super terminos terrae
JOB|37|4|post eum rugiet sonitus tonabit voce magnitudinis suae et non investigabitur cum audita fuerit vox eius
JOB|37|5|tonabit Deus in voce sua mirabiliter qui facit magna et inscrutabilia
JOB|37|6|qui praecipit nivi ut descendat in terram et hiemis pluviis et imbri fortitudinis suae
JOB|37|7|qui in manu omnium hominum signat ut noverint singuli opera sua
JOB|37|8|ingredietur bestia latibulum et in antro suo morabitur
JOB|37|9|ab interioribus egreditur tempestas et ab Arcturo frigus
JOB|37|10|flante Deo concrescit gelu et rursum latissimae funduntur aquae
JOB|37|11|frumentum desiderat nubes et nubes spargunt lumen suum
JOB|37|12|quae lustrant per circuitum quocumque eas voluntas gubernantis duxerit ad omne quod praeceperit illis super faciem orbis terrarum
JOB|37|13|sive in una tribu sive in terra sua sive in quocumque loco misericordiae suae eas iusserit inveniri
JOB|37|14|ausculta haec Iob sta et considera miracula Dei
JOB|37|15|numquid scis quando praeceperit Deus pluviis ut ostenderent lucem nubium eius
JOB|37|16|numquid nosti semitas nubium magnas et perfectas scientias
JOB|37|17|nonne vestimenta tua calida sunt cum perflata fuerit terra austro
JOB|37|18|tu forsitan cum eo fabricatus es caelos qui solidissimi quasi aere fusi sunt
JOB|37|19|ostende nobis quid dicamus illi nos quippe involvimur tenebris
JOB|37|20|quis narrabit ei quae loquor etiam si locutus fuerit homo devorabitur
JOB|37|21|at nunc non vident lucem subito aer cogitur in nubes et ventus transiens fugabit eas
JOB|37|22|ab aquilone aurum venit et ad Deum formidolosa laudatio
JOB|37|23|digne eum invenire non possumus magnus fortitudine et iudicio et iustitia et enarrari non potest
JOB|37|24|ideo timebunt eum viri et non audebunt contemplari omnes qui sibi videntur esse sapientes
JOB|38|1|respondens autem Dominus Iob de turbine dixit
JOB|38|2|quis est iste involvens sententias sermonibus inperitis
JOB|38|3|accinge sicut vir lumbos tuos interrogabo te et responde mihi
JOB|38|4|ubi eras quando ponebam fundamenta terrae indica mihi si habes intellegentiam
JOB|38|5|quis posuit mensuras eius si nosti vel quis tetendit super eam lineam
JOB|38|6|super quo bases illius solidatae sunt aut quis dimisit lapidem angularem eius
JOB|38|7|cum me laudarent simul astra matutina et iubilarent omnes filii Dei
JOB|38|8|quis conclusit ostiis mare quando erumpebat quasi de vulva procedens
JOB|38|9|cum ponerem nubem vestimentum eius et caligine illud quasi pannis infantiae obvolverem
JOB|38|10|circumdedi illud terminis meis et posui vectem et ostia
JOB|38|11|et dixi usque huc venies et non procedes amplius et hic confringes tumentes fluctus tuos
JOB|38|12|numquid post ortum tuum praecepisti diluculo et ostendisti aurorae locum suum
JOB|38|13|et tenuisti concutiens extrema terrae et excussisti impios ex ea
JOB|38|14|restituetur ut lutum signaculum et stabit sicut vestimentum
JOB|38|15|auferetur ab impiis lux sua et brachium excelsum confringetur
JOB|38|16|numquid ingressus es profunda maris et in novissimis abyssis deambulasti
JOB|38|17|numquid apertae tibi sunt portae mortis et ostia tenebrosa vidisti
JOB|38|18|numquid considerasti latitudines terrae indica mihi si nosti omnia
JOB|38|19|in qua via habitet lux et tenebrarum quis locus sit
JOB|38|20|ut ducas unumquodque ad terminos suos et intellegas semitas domus eius
JOB|38|21|sciebas tunc quod nasciturus esses et numerum dierum tuorum noveras
JOB|38|22|numquid ingressus es thesauros nivis aut thesauros grandinis aspexisti
JOB|38|23|quae praeparavi in tempus hostis in diem pugnae et belli
JOB|38|24|per quam viam spargitur lux dividitur aestus super terram
JOB|38|25|quis dedit vehementissimo imbri cursum et viam sonantis tonitrui
JOB|38|26|ut plueret super terram absque homine in deserto ubi nullus mortalium commoratur
JOB|38|27|ut impleret inviam et desolatam et produceret herbas virentes
JOB|38|28|quis est pluviae pater vel quis genuit stillas roris
JOB|38|29|de cuius utero egressa est glacies et gelu de caelo quis genuit
JOB|38|30|in similitudinem lapidis aquae durantur et superficies abyssi constringitur
JOB|38|31|numquid coniungere valebis micantes stellas Pliadis aut gyrum Arcturi poteris dissipare
JOB|38|32|numquid producis luciferum in tempore suo et vesperum super filios terrae consurgere facis
JOB|38|33|numquid nosti ordinem caeli et pones rationem eius in terra
JOB|38|34|numquid elevabis in nebula vocem tuam et impetus aquarum operiet te
JOB|38|35|numquid mittes fulgura et ibunt et revertentia dicent tibi adsumus
JOB|38|36|quis posuit in visceribus hominis sapientiam vel quis dedit gallo intellegentiam
JOB|38|37|quis enarravit caelorum rationem et concentum caeli quis dormire faciet
JOB|38|38|quando fundebatur pulvis in terram et glebae conpingebantur
JOB|38|39|numquid capies leaenae praedam et animam catulorum eius implebis
JOB|38|40|quando cubant in antris et in specubus insidiantur
JOB|38|41|quis praeparat corvo escam suam quando pulli eius ad Deum clamant vagantes eo quod non habeant cibos
JOB|39|1|numquid nosti tempus partus hibicum in petris vel parturientes cervas observasti
JOB|39|2|dinumerasti menses conceptus earum et scisti tempus partus earum
JOB|39|3|incurvantur ad fetum et pariunt et rugitus emittunt
JOB|39|4|separantur filii earum pergunt ad pastum egrediuntur et non revertuntur ad eas
JOB|39|5|quis dimisit onagrum liberum et vincula eius quis solvit
JOB|39|6|cui dedi in solitudine domum et tabernacula eius in terra salsuginis
JOB|39|7|contemnit multitudinem civitatis clamorem exactoris non audit
JOB|39|8|circumspicit montes pascuae suae et virentia quaeque perquirit
JOB|39|9|numquid volet rinoceros servire tibi aut morabitur ad praesepe tuum
JOB|39|10|numquid alligabis rinocerota ad arandum loro tuo aut confringet glebas vallium post te
JOB|39|11|numquid fiduciam habebis in magna fortitudine eius et derelinques ei labores tuos
JOB|39|12|numquid credes ei quoniam reddat sementem tibi et aream tuam congreget
JOB|39|13|pinna strutionum similis est pinnis herodii et accipitris
JOB|39|14|quando derelinquit in terra ova sua tu forsitan in pulvere calefacis ea
JOB|39|15|obliviscitur quod pes conculcet ea aut bestiae agri conterant
JOB|39|16|duratur ad filios suos quasi non sint sui frustra laboravit nullo timore cogente
JOB|39|17|privavit enim eam Deus sapientia nec dedit illi intellegentiam
JOB|39|18|cum tempus fuerit in altum alas erigit deridet equitem et ascensorem eius
JOB|39|19|numquid praebebis equo fortitudinem aut circumdabis collo eius hinnitum
JOB|39|20|numquid suscitabis eum quasi lucustas gloria narium eius terror
JOB|39|21|terram ungula fodit exultat audacter in occursum pergit armatis
JOB|39|22|contemnit pavorem nec cedit gladio
JOB|39|23|super ipsum sonabit faretra vibrabit hasta et clypeus
JOB|39|24|fervens et fremens sorbet terram nec reputat tubae sonare clangorem
JOB|39|25|ubi audierit bucinam dicet va procul odoratur bellum exhortationem ducum et ululatum exercitus
JOB|39|26|numquid per sapientiam tuam plumescit accipiter expandens alas suas ad austrum
JOB|39|27|aut ad praeceptum tuum elevabitur aquila et in arduis ponet nidum suum
JOB|39|28|in petris manet et in praeruptis silicibus commoratur atque inaccessis rupibus
JOB|39|29|inde contemplatur escam et de longe oculi eius prospiciunt
JOB|39|30|pulli eius lambent sanguinem et ubicumque cadaver fuerit statim adest
JOB|39|31|et adiecit Dominus et locutus est ad Iob
JOB|39|32|numquid qui contendit cum Deo tam facile conquiescit utique qui arguit Deum debet respondere ei
JOB|39|33|respondens autem Iob Domino dixit
JOB|39|34|qui leviter locutus sum respondere quid possum manum meam ponam super os meum
JOB|39|35|unum locutus sum quod utinam non dixissem et alterum quibus ultra non addam
JOB|40|1|respondens autem Dominus Iob de turbine ait
JOB|40|2|accinge sicut vir lumbos tuos interrogabo te et indica mihi
JOB|40|3|numquid irritum facies iudicium meum et condemnabis me ut tu iustificeris
JOB|40|4|et si habes brachium sicut Deus et si voce simili tonas
JOB|40|5|circumda tibi decorem et in sublime erigere et esto gloriosus et speciosis induere vestibus
JOB|40|6|disperge superbos furore tuo et respiciens omnem arrogantem humilia
JOB|40|7|respice cunctos superbos et confunde eos et contere impios in loco suo
JOB|40|8|absconde eos in pulvere simul et facies eorum demerge in foveam
JOB|40|9|et ego confitebor quod salvare te possit dextera tua
JOB|40|10|ecce Behemoth quem feci tecum faenum quasi bos comedet
JOB|40|11|fortitudo eius in lumbis eius et virtus illius in umbilicis ventris eius
JOB|40|12|constringit caudam suam quasi cedrum nervi testiculorum eius perplexi sunt
JOB|40|13|ossa eius velut fistulae aeris cartilago illius quasi lamminae ferreae
JOB|40|14|ipse principium est viarum Dei qui fecit eum adplicabit gladium eius
JOB|40|15|huic montes herbas ferunt omnes bestiae agri ludent ibi
JOB|40|16|sub umbra dormit in secreto calami et locis humentibus
JOB|40|17|protegunt umbrae umbram eius circumdabunt eum salices torrentis
JOB|40|18|ecce absorbebit fluvium et non mirabitur habet fiduciam quod influat Iordanis in os eius
JOB|40|19|in oculis eius quasi hamo capiet eum et in sudibus perforabit nares eius
JOB|40|20|an extrahere poteris Leviathan hamo et fune ligabis linguam eius
JOB|40|21|numquid pones circulum in naribus eius et armilla perforabis maxillam eius
JOB|40|22|numquid multiplicabit ad te preces aut loquetur tibi mollia
JOB|40|23|numquid feriet tecum pactum et accipies eum servum sempiternum
JOB|40|24|numquid inludes ei quasi avi aut ligabis illum ancillis tuis
JOB|40|25|concident eum amici divident illum negotiatores
JOB|40|26|numquid implebis sagenas pelle eius et gurgustium piscium capite illius
JOB|40|27|pone super eum manum tuam memento belli nec ultra addas loqui
JOB|40|28|ecce spes eius frustrabitur eum et videntibus cunctis praecipitabitur
JOB|41|1|non quasi crudelis suscitabo eum quis enim resistere potest vultui meo
JOB|41|2|quis ante dedit mihi ut reddam ei omnia quae sub caelo sunt mea sunt
JOB|41|3|non parcam ei et verbis potentibus et ad deprecandum conpositis
JOB|41|4|quis revelavit faciem indumenti eius et in medium oris eius quis intrabit
JOB|41|5|portas vultus eius quis aperiet per gyrum dentium eius formido
JOB|41|6|corpus illius quasi scuta fusilia et conpactum squamis se prementibus
JOB|41|7|una uni coniungitur et ne spiraculum quidem incedit per eas
JOB|41|8|una alteri adherebunt et tenentes se nequaquam separabuntur
JOB|41|9|sternutatio eius splendor ignis et oculi eius ut palpebrae diluculi
JOB|41|10|de ore eius lampades procedunt sicut taedae ignis accensae
JOB|41|11|de naribus eius procedit fumus sicut ollae succensae atque ferventis
JOB|41|12|halitus eius prunas ardere facit et flamma de ore eius egreditur
JOB|41|13|in collo eius morabitur fortitudo et faciem eius praecedet egestas
JOB|41|14|membra carnium eius coherentia sibi mittet contra eum fulmina et ad locum alium non ferentur
JOB|41|15|cor eius indurabitur quasi lapis et stringetur quasi malleatoris incus
JOB|41|16|cum sublatus fuerit timebunt angeli et territi purgabuntur
JOB|41|17|cum adprehenderit eum gladius subsistere non poterit neque hasta neque torax
JOB|41|18|reputabit enim quasi paleas ferrum et quasi lignum putridum aes
JOB|41|19|non fugabit eum vir sagittarius in stipulam versi sunt ei lapides fundae
JOB|41|20|quasi stipulam aestimabit malleum et deridebit vibrantem hastam
JOB|41|21|sub ipso erunt radii solis sternet sibi aurum quasi lutum
JOB|41|22|fervescere faciet quasi ollam profundum mare ponet quasi cum unguenta bulliunt
JOB|41|23|post eum lucebit semita aestimabit abyssum quasi senescentem
JOB|41|24|non est super terram potestas quae conparetur ei qui factus est ut nullum timeret
JOB|41|25|omne sublime videt ipse est rex super universos filios superbiae
JOB|42|1|respondens autem Iob Domino dixit
JOB|42|2|scio quia omnia potes et nulla te latet cogitatio
JOB|42|3|quis est iste qui celat consilium absque scientia ideo insipienter locutus sum et quae ultra modum excederent scientiam meam
JOB|42|4|audi et ego loquar interrogabo et ostende mihi
JOB|42|5|auditu auris audivi te nunc autem oculus meus videt te
JOB|42|6|idcirco ipse me reprehendo et ago paenitentiam in favilla et cinere
JOB|42|7|postquam autem locutus est Dominus verba haec ad Iob dixit ad Eliphaz Themaniten iratus est furor meus in te et in duos amicos tuos quoniam non estis locuti coram me rectum sicut servus meus Iob
JOB|42|8|sumite igitur vobis septem tauros et septem arietes et ite ad servum meum Iob et offerte holocaustum pro vobis Iob autem servus meus orabit pro vobis faciem eius suscipiam ut non vobis inputetur stultitia neque enim locuti estis ad me recta sicut servus meus Iob
JOB|42|9|abierunt ergo Eliphaz Themanites et Baldad Suites et Sophar Naamathites et fecerunt sicut locutus fuerat ad eos Dominus et suscepit Dominus faciem Iob
JOB|42|10|Dominus quoque conversus est ad paenitentiam Iob cum oraret ille pro amicis suis et addidit Dominus omnia quaecumque fuerant Iob duplicia
JOB|42|11|venerunt autem ad eum omnes fratres sui et universae sorores suae et cuncti qui noverant eum prius et comederunt cum eo panem in domo eius et moverunt super eum caput et consolati sunt eum super omni malo quod intulerat Dominus super eum et dederunt ei unusquisque ovem unam et inaurem auream unam
JOB|42|12|Dominus autem benedixit novissimis Iob magis quam principio eius et facta sunt ei quattuordecim milia ovium et sex milia camelorum et mille iuga boum et mille asinae
JOB|42|13|et fuerunt ei septem filii et filiae tres
JOB|42|14|et vocavit nomen unius Diem et nomen secundae Cassia et nomen tertiae Cornu stibii
JOB|42|15|non sunt autem inventae mulieres speciosae sicut filiae Iob in universa terra deditque eis pater suus hereditatem inter fratres earum
JOB|42|16|vixit autem Iob post haec centum quadraginta annis et vidit filios suos et filios filiorum suorum usque ad quartam generationem et mortuus est senex et plenus dierum
PS|1|1|beatus vir qui non abiit in consilio impiorum et in via peccatorum non stetit et in cathedra pestilentiae non sedit
PS|1|2|sed in lege Domini voluntas eius et in lege eius meditabitur die ac nocte
PS|1|3|et erit tamquam lignum quod plantatum est secus decursus aquarum quod fructum suum dabit in tempore suo et folium eius non defluet et omnia quaecumque faciet prosperabuntur
PS|1|4|non sic impii non sic; sed tamquam pulvis quem proicit ventus a facie terrae;
PS|1|5|ideo non resurgent impii in iudicio neque peccatores in consilio iustorum
PS|1|6|quoniam novit Dominus viam iustorum et iter impiorum peribit
PS|2|1|psalmus David quare fremuerunt gentes et populi meditati sunt inania
PS|2|2|adstiterunt reges terrae et principes convenerunt in unum adversus Dominum et adversus christum eius diapsalma
PS|2|3|disrumpamus vincula eorum et proiciamus a nobis iugum ipsorum
PS|2|4|qui habitat in caelis inridebit eos et Dominus subsannabit eos
PS|2|5|tunc loquetur ad eos in ira sua et in furore suo conturbabit eos
PS|2|6|ego autem constitutus sum rex ab eo super Sion montem sanctum eius praedicans praeceptum eius
PS|2|7|Dominus dixit ad me filius meus es tu ego hodie genui te
PS|2|8|postula a me et dabo tibi gentes hereditatem tuam et possessionem tuam terminos terrae
PS|2|9|reges eos in virga ferrea tamquam vas figuli confringes eos
PS|2|10|et nunc reges intellegite erudimini qui iudicatis terram
PS|2|11|servite Domino in timore et exultate ei in tremore
PS|2|12|adprehendite disciplinam nequando irascatur Dominus et pereatis de via iusta
PS|2|13|cum exarserit in brevi ira eius beati omnes qui confidunt in eo
PS|3|1|psalmus David cum fugeret a facie Abessalon filii sui
PS|3|2|Domine quid multiplicati sunt qui tribulant me multi insurgunt adversum me
PS|3|3|multi dicunt animae meae non est salus ipsi in Deo eius; diapsalma
PS|3|4|tu autem Domine susceptor meus es gloria mea et exaltans caput meum
PS|3|5|voce mea ad Dominum clamavi et exaudivit me de monte sancto suo diapsalma
PS|3|6|ego dormivi et soporatus sum exsurrexi quia Dominus suscipiet me
PS|3|7|non timebo milia populi circumdantis me exsurge Domine salvum me fac Deus meus
PS|3|8|quoniam tu percussisti omnes adversantes mihi sine causa dentes peccatorum contrivisti
PS|3|9|Domini est salus et super populum tuum benedictio tua
PS|4|1|in finem in carminibus psalmus David
PS|4|2|cum invocarem exaudivit me Deus iustitiae meae in tribulatione dilatasti mihi miserere mei et exaudi orationem meam
PS|4|3|filii hominum usquequo gravi corde ut quid diligitis vanitatem et quaeritis mendacium diapsalma
PS|4|4|et scitote quoniam mirificavit Dominus sanctum suum Dominus exaudiet me cum clamavero ad eum
PS|4|5|irascimini et nolite peccare quae dicitis in cordibus vestris in cubilibus vestris conpungimini diapsalma
PS|4|6|sacrificate sacrificium iustitiae et sperate in Domino multi dicunt quis ostendet nobis bona
PS|4|7|signatum est super nos lumen vultus tui Domine dedisti laetitiam in corde meo
PS|4|8|a fructu frumenti et vini et olei sui multiplicati sunt
PS|4|9|in pace in id ipsum dormiam et requiescam
PS|4|10|quoniam tu Domine singulariter in spe constituisti me
PS|5|1|in finem pro ea quae hereditatem consequitur psalmus David
PS|5|2|verba mea auribus percipe Domine intellege clamorem meum
PS|5|3|intende voci orationis meae rex meus et Deus meus
PS|5|4|quoniam ad te orabo Domine mane exaudies vocem meam
PS|5|5|mane adstabo tibi et videbo quoniam non deus volens iniquitatem tu es
PS|5|6|neque habitabit iuxta te malignus neque permanebunt iniusti ante oculos tuos
PS|5|7|odisti omnes qui operantur iniquitatem perdes %omnes; qui loquuntur mendacium virum sanguinum et dolosum abominabitur Dominus
PS|5|8|ego autem in multitudine misericordiae tuae introibo in domum tuam adorabo ad templum sanctum tuum in timore tuo
PS|5|9|Domine deduc me in iustitia tua propter inimicos meos dirige in conspectu meo viam tuam
PS|5|10|quoniam non est in ore eorum veritas cor eorum vanum est
PS|5|11|sepulchrum patens est guttur eorum linguis suis dolose agebant iudica illos Deus decidant a cogitationibus suis secundum multitudinem impietatum eorum expelle eos quoniam inritaverunt te Domine
PS|5|12|et laetentur omnes qui sperant in te in aeternum exultabunt et habitabis in eis et gloriabuntur in te omnes qui diligunt nomen tuum
PS|5|13|quoniam tu benedices iusto Domine ut scuto bonae voluntatis coronasti nos
PS|6|1|in finem in carminibus pro octava psalmus David
PS|6|2|Domine ne in furore tuo arguas me neque in ira tua corripias me
PS|6|3|miserere mei Domine quoniam infirmus sum sana me Domine quoniam conturbata sunt ossa mea
PS|6|4|et anima mea turbata est valde et tu Domine usquequo
PS|6|5|convertere Domine eripe animam meam salvum me fac propter misericordiam tuam
PS|6|6|quoniam non est in morte qui memor sit tui in inferno autem quis confitebitur tibi
PS|6|7|laboravi in gemitu meo lavabo per singulas noctes lectum meum in lacrimis meis stratum meum rigabo
PS|6|8|turbatus est a furore oculus meus inveteravi inter omnes inimicos meos
PS|6|9|discedite a me omnes qui operamini iniquitatem quoniam exaudivit Dominus vocem fletus mei
PS|6|10|exaudivit Dominus deprecationem meam Dominus orationem meam suscepit
PS|6|11|erubescant et conturbentur vehementer omnes inimici mei convertantur et erubescant valde velociter
PS|7|1|psalmus David quem cantavit Domino pro verbis Chusi filii Iemini
PS|7|2|Domine Deus meus in te speravi salvum me fac ex omnibus persequentibus me et libera me
PS|7|3|nequando rapiat ut leo animam meam dum non est qui redimat neque qui salvum faciat
PS|7|4|Domine Deus meus si feci istud si est iniquitas in manibus meis
PS|7|5|si reddidi retribuentibus mihi mala decidam merito ab inimicis meis inanis
PS|7|6|persequatur inimicus animam meam et conprehendat et conculcet in terra vitam meam et gloriam meam in pulverem deducat diapsalma
PS|7|7|exsurge Domine in ira tua exaltare in finibus inimicorum meorum et exsurge Domine Deus meus in praecepto quod mandasti
PS|7|8|et synagoga populorum circumdabit te et propter hanc in altum regredere
PS|7|9|Dominus iudicat populos iudica me Domine secundum iustitiam meam et secundum innocentiam meam super me
PS|7|10|consummetur nequitia peccatorum et diriges iustum et scrutans corda et renes Deus
PS|7|11|iustum adiutorium meum a Deo qui salvos facit rectos corde
PS|7|12|Deus iudex iustus et fortis et patiens numquid irascitur per singulos dies
PS|7|13|nisi conversi fueritis gladium suum vibrabit arcum suum tetendit et paravit illum
PS|7|14|et in eo paravit vasa mortis sagittas suas ardentibus effecit
PS|7|15|ecce parturiit iniustitiam et; concepit dolorem et peperit iniquitatem
PS|7|16|lacum aperuit et effodit eum et incidet in foveam quam fecit
PS|7|17|convertetur dolor eius in caput eius et in verticem ipsius iniquitas eius descendet
PS|7|18|confitebor Domino secundum iustitiam eius et psallam nomini Domini altissimi
PS|8|1|in finem pro torcularibus psalmus David
PS|8|2|Domine Dominus noster quam admirabile est nomen tuum in universa terra quoniam elevata est magnificentia tua super caelos
PS|8|3|ex ore infantium et lactantium perfecisti laudem propter inimicos tuos ut destruas inimicum et ultorem
PS|8|4|quoniam videbo caelos tuos; opera digitorum tuorum lunam et stellas quae tu fundasti
PS|8|5|quid est homo quod memor es eius aut filius hominis quoniam visitas eum
PS|8|6|minuisti eum paulo minus ab angelis gloria et honore coronasti eum
PS|8|7|et constituisti eum super opera manuum tuarum
PS|8|8|omnia subiecisti sub pedibus eius oves et boves universas insuper et pecora campi
PS|8|9|volucres caeli et pisces maris qui perambulant semitas maris
PS|8|10|Domine Dominus noster quam admirabile est nomen tuum in universa terra
PS|9|1|in finem pro occultis filii psalmus David
PS|9|2|confitebor tibi Domine in toto corde meo narrabo omnia mirabilia tua
PS|9|3|laetabor et exultabo in te psallam nomini tuo Altissime
PS|9|4|in convertendo inimicum meum retrorsum infirmabuntur et peribunt a facie tua
PS|9|5|quoniam fecisti iudicium meum et causam meam sedisti super thronum qui iudicas iustitiam
PS|9|6|increpasti gentes %et; periit impius nomen eorum delisti in aeternum et in saeculum %saeculi;
PS|9|7|inimici defecerunt frameae in finem et civitates destruxisti periit memoria eorum cum sonitu
PS|9|8|et Dominus in aeternum permanet paravit in iudicio thronum suum
PS|9|9|et ipse iudicabit orbem terrae in aequitate iudicabit populos in iustitia
PS|9|10|et factus est Dominus refugium pauperi adiutor in oportunitatibus in tribulatione
PS|9|11|et sperent in te qui noverunt nomen tuum quoniam non dereliquisti quaerentes te Domine
PS|9|12|psallite Domino qui habitat in Sion adnuntiate inter gentes studia eius
PS|9|13|quoniam requirens sanguinem eorum recordatus est non est oblitus clamorem pauperum
PS|9|14|miserere mei Domine vide humilitatem meam de inimicis meis
PS|9|15|qui exaltas me de portis mortis ut adnuntiem omnes laudationes tuas in portis filiae Sion
PS|9|16|exultabo in salutari tuo infixae sunt gentes in interitu quem fecerunt in laqueo isto quem absconderunt conprehensus est pes eorum
PS|9|17|cognoscitur Dominus iudicia faciens in operibus manuum suarum conprehensus est peccator canticum diapsalmatis
PS|9|18|convertantur peccatores in infernum omnes gentes quae obliviscuntur Deum
PS|9|19|quoniam non in finem oblivio erit pauperis patientia pauperum non peribit in finem
PS|9|20|exsurge Domine non confortetur homo iudicentur gentes in conspectu tuo
PS|9|21|constitue Domine legislatorem super eos sciant gentes quoniam homines sunt diapsalma
PS|9|22|ut quid Domine recessisti longe dispicis in oportunitatibus in tribulatione
PS|9|23|dum superbit impius incenditur pauper conprehenduntur in consiliis quibus cogitant
PS|9|24|quoniam laudatur peccator in desideriis animae suae et iniquus benedicitur
PS|9|25|exacerbavit Dominum peccator secundum multitudinem irae suae non quaeret
PS|9|26|non est Deus in conspectu eius inquinatae sunt viae illius in omni tempore auferuntur iudicia tua a facie eius omnium inimicorum suorum dominabitur
PS|9|27|dixit enim in corde suo non movebor a generatione in generationem sine malo
PS|9|28|cuius maledictione os plenum est et amaritudine et dolo sub lingua eius labor et dolor
PS|9|29|sedet in insidiis cum divitibus in occultis ut interficiat innocentem
PS|9|30|oculi eius in pauperem respiciunt insidiatur in abscondito quasi leo in spelunca sua insidiatur ut rapiat pauperem rapere pauperem dum adtrahit eum
PS|9|31|in laqueo suo humiliabit eum inclinabit se et cadet cum dominatus fuerit pauperum
PS|9|32|dixit enim in corde suo oblitus est Deus avertit faciem suam ne videat in finem
PS|9|33|exsurge Domine Deus exaltetur manus tua ne obliviscaris pauperum
PS|9|34|propter quid inritavit impius Deum dixit enim in corde suo non requiret
PS|9|35|vides quoniam tu laborem et dolorem consideras ut tradas eos in manus tuas tibi derelictus est pauper orfano tu eras adiutor
PS|9|36|contere brachium peccatoris et maligni quaeretur peccatum illius et non invenietur
PS|9|37|Dominus regnabit in aeternum et in saeculum %saeculi; peribitis gentes de terra illius
PS|9|38|desiderium pauperum exaudivit Dominus praeparationem cordis eorum audivit auris tua
PS|9|39|iudicare pupillo et humili ut non adponat ultra magnificare se homo super terram
PS|10|1|in finem psalmus David
PS|10|2|in Domino confido quomodo dicitis animae meae transmigra in montes sicut passer
PS|10|3|quoniam ecce peccatores intenderunt arcum paraverunt sagittas suas in faretra ut sagittent in obscuro rectos corde
PS|10|4|quoniam quae perfecisti destruxerunt iustus %autem; quid fecit
PS|10|5|Dominus in templo sancto suo Dominus in caelo sedis eius oculi eius %in pauperem; respiciunt palpebrae eius interrogant filios hominum
PS|10|6|Dominus interrogat iustum et impium qui autem diligit iniquitatem odit animam suam
PS|10|7|pluet super peccatores laqueos ignis et sulphur et spiritus procellarum pars calicis eorum
PS|10|8|quoniam iustus Dominus %et; iustitias dilexit aequitatem vidit vultus eius
PS|11|1|in finem pro octava psalmus David
PS|11|2|salvum me fac Domine quoniam defecit sanctus quoniam deminutae sunt veritates a filiis hominum
PS|11|3|vana locuti sunt unusquisque ad proximum suum labia dolosa in corde et corde locuti sunt
PS|11|4|disperdat Dominus universa labia dolosa linguam magniloquam
PS|11|5|qui dixerunt linguam nostram magnificabimus labia nostra a nobis sunt quis noster dominus est
PS|11|6|propter miseriam inopum et gemitum pauperum nunc exsurgam dicit Dominus ponam in salutari fiducialiter agam in eo
PS|11|7|eloquia Domini eloquia casta argentum igne examinatum probatum terrae purgatum septuplum
PS|11|8|tu Domine servabis nos et custodies nos a generatione hac et in aeternum
PS|11|9|in circuitu impii ambulant secundum altitudinem tuam multiplicasti filios hominum
PS|12|1|in finem psalmus David usquequo Domine oblivisceris me in finem usquequo avertis faciem tuam a me
PS|12|2|quamdiu ponam consilia in anima mea dolorem in corde meo per diem
PS|12|3|usquequo exaltabitur inimicus meus super me
PS|12|4|respice exaudi me Domine Deus meus inlumina oculos meos ne umquam obdormiam in mortem
PS|12|5|nequando dicat inimicus meus praevalui adversus eum qui tribulant me exultabunt si motus fuero
PS|12|6|ego autem in misericordia tua speravi exultabit cor meum in salutari tuo cantabo Domino qui bona tribuit mihi et psallam nomini Domini altissimi
PS|13|1|in finem psalmus David dixit insipiens in corde suo non est Deus corrupti sunt et abominabiles facti sunt in studiis %suis; non est qui faciat bonum %non est usque ad unum;
PS|13|2|Dominus de caelo prospexit super filios hominum ut videat si est intellegens %aut; requirens Deum
PS|13|3|omnes declinaverunt simul inutiles facti sunt non est qui faciat bonum non est usque ad unum = sepulchrum patens est guttur eorum = linguis suis dolose agebant = venenum aspidum sub labiis eorum = quorum os maledictione et amaritudine plenum est = veloces pedes eorum ad effundendum sanguinem = contritio et infelicitas in viis eorum = et viam pacis non cognoverunt % non est timor Dei ante oculos eorum;
PS|13|4|nonne cognoscent omnes qui operantur iniquitatem qui devorant plebem meam sicut escam panis
PS|13|5|Dominum non invocaverunt illic trepidaverunt timore %ubi non erat timor;
PS|13|6|quoniam Deus in generatione iusta consilium inopis confudistis quoniam Dominus spes eius est
PS|13|7|quis dabit ex Sion salutare Israhel cum averterit Dominus captivitatem plebis suae exultabit Iacob et laetabitur Israhel
PS|14|1|psalmus David Domine quis habitabit in tabernaculo tuo aut quis requiescet in monte sancto tuo
PS|14|2|qui ingreditur sine macula et operatur iustitiam
PS|14|3|qui loquitur veritatem in corde suo qui non egit dolum in lingua sua nec fecit proximo suo malum et obprobrium non accepit adversus proximos suos
PS|14|4|ad nihilum deductus est in conspectu eius malignus timentes autem Dominum glorificat qui iurat proximo suo et non decipit
PS|14|5|qui pecuniam suam non dedit ad usuram et munera super innocentes non accepit qui facit haec non movebitur in aeternum
PS|15|1|tituli inscriptio ipsi David conserva me Domine quoniam in te speravi
PS|15|2|dixi Domino Dominus meus es tu quoniam bonorum meorum non eges
PS|15|3|sanctis qui sunt in terra eius mirificavit mihi; omnes voluntates meas in eis
PS|15|4|multiplicatae sunt infirmitates eorum postea adceleraverunt non congregabo conventicula eorum de sanguinibus nec memor ero nominum eorum per labia mea
PS|15|5|Dominus pars hereditatis meae et calicis mei tu es qui restitues hereditatem meam mihi
PS|15|6|funes ceciderunt mihi in praeclaris etenim hereditas mea praeclara est mihi
PS|15|7|benedicam Domino qui tribuit mihi intellectum insuper et usque ad noctem increpaverunt me renes mei
PS|15|8|providebam Dominum in conspectu meo semper quoniam a dextris est mihi ne commovear
PS|15|9|propter hoc laetatum est cor meum et exultavit lingua mea insuper et caro mea requiescet in spe
PS|15|10|quoniam non derelinques animam meam in inferno non dabis sanctum tuum videre corruptionem notas mihi fecisti vias vitae adimplebis me laetitia cum vultu tuo delectatio in dextera tua usque in finem
PS|16|1|oratio David exaudi Domine iustitiam meam intende deprecationem meam auribus percipe orationem meam non in labiis dolosis
PS|16|2|de vultu tuo iudicium meum prodeat oculi tui videant aequitates
PS|16|3|probasti cor meum visitasti nocte igne me examinasti et non est inventa in me iniquitas
PS|16|4|ut non loquatur os meum opera hominum propter verba labiorum tuorum ego custodivi vias duras
PS|16|5|perfice gressus meos in semitis tuis ut non moveantur vestigia mea
PS|16|6|ego clamavi quoniam exaudisti me Deus inclina aurem tuam mihi et exaudi verba mea
PS|16|7|mirifica misericordias tuas qui salvos facis sperantes in te
PS|16|8|a resistentibus dexterae tuae custodi me ut pupillam oculi sub umbra alarum tuarum proteges me
PS|16|9|a facie impiorum qui me adflixerunt inimici mei animam meam circumdederunt super me;
PS|16|10|adipem suum concluserunt os eorum locutum est superbia
PS|16|11|proicientes me nunc circumdederunt me oculos suos statuerunt declinare in terram
PS|16|12|susceperunt me sicut leo paratus ad praedam et sicut catulus leonis habitans in abditis
PS|16|13|exsurge Domine praeveni eum et subplanta eum eripe animam meam ab impio frameam tuam
PS|16|14|ab inimicis manus tuae Domine a paucis de terra divide eos in vita eorum de absconditis tuis adimpletus est venter eorum saturati sunt filiis et dimiserunt reliquias suas parvulis suis
PS|16|15|ego autem in iustitia apparebo conspectui tuo satiabor cum apparuerit gloria tua
PS|17|1|in finem puero Domini David quae locutus est Domino verba cantici huius in die qua eripuit eum Dominus de manu omnium inimicorum eius et de manu Saul et dixit
PS|17|2|diligam te Domine fortitudo mea
PS|17|3|Dominus firmamentum meum et refugium meum et liberator meus Deus meus adiutor meus et sperabo in eum protector meus et cornu salutis meae et susceptor meus
PS|17|4|laudans invocabo Dominum et ab inimicis meis salvus ero
PS|17|5|circumdederunt me dolores mortis et torrentes iniquitatis conturbaverunt me
PS|17|6|dolores inferni circumdederunt me praeoccupaverunt me laquei mortis
PS|17|7|cum tribularer invocavi Dominum et ad Deum meum clamavi exaudivit de templo %sancto; suo vocem meam et clamor meus in conspectu eius introibit in aures eius
PS|17|8|et commota est et contremuit terra et fundamenta montium conturbata sunt et commota sunt quoniam iratus est eis
PS|17|9|ascendit fumus in ira eius et ignis a facie eius exarsit carbones succensi sunt ab eo
PS|17|10|inclinavit caelos et descendit et caligo sub pedibus eius
PS|17|11|et ascendit super cherubin et volavit volavit super pinnas ventorum
PS|17|12|et posuit tenebras latibulum suum in circuitu eius tabernaculum eius tenebrosa aqua in nubibus aeris
PS|17|13|prae fulgore in conspectu eius nubes eius; transierunt grando et carbones ignis
PS|17|14|et intonuit de caelo Dominus et Altissimus dedit vocem suam grando et carbones ignis;
PS|17|15|et misit sagittas et dissipavit eos et fulgora multiplicavit et conturbavit eos
PS|17|16|et apparuerunt fontes aquarum et revelata sunt fundamenta orbis terrarum ab increpatione tua Domine ab inspiratione spiritus irae tuae
PS|17|17|misit de summo et accepit me adsumpsit me de aquis multis
PS|17|18|eripiet me de inimicis meis fortissimis et ab his qui oderunt me quoniam confirmati sunt super me
PS|17|19|praevenerunt me in die adflictionis meae et factus est Dominus protector meus
PS|17|20|et eduxit me in latitudinem salvum me faciet quoniam voluit me
PS|17|21|%et; retribuet mihi Dominus secundum iustitiam meam %et; secundum puritatem manuum mearum retribuet mihi
PS|17|22|quia custodivi vias Domini nec impie gessi a Deo meo
PS|17|23|quoniam omnia iudicia eius in conspectu meo sunt et iustitias eius non reppuli a me
PS|17|24|et ero inmaculatus cum eo et observabo ab iniquitate mea
PS|17|25|et retribuet mihi Dominus secundum iustitiam meam et secundum puritatem manuum mearum in conspectu oculorum eius
PS|17|26|cum sancto sanctus eris et cum viro innocente innocens eris
PS|17|27|et cum electo electus eris et cum perverso perverteris
PS|17|28|quoniam tu populum humilem salvum facies et oculos superborum humiliabis
PS|17|29|quoniam tu inluminas lucernam meam Domine Deus meus inluminas tenebras meas
PS|17|30|quoniam in te eripiar a temptatione et in Deo meo transgrediar murum
PS|17|31|Deus meus inpolluta via eius eloquia Domini igne examinata protector est omnium sperantium in eum
PS|17|32|quoniam quis deus praeter Dominum et quis deus praeter Deum nostrum
PS|17|33|Deus qui praecingit me virtute et posuit inmaculatam viam meam
PS|17|34|qui perfecit pedes meos tamquam cervorum et super excelsa statuens me
PS|17|35|qui doces manus meas in proelium et posuisti arcum aereum brachia mea
PS|17|36|et dedisti mihi protectionem salutis tuae et dextera tua suscepit me et disciplina tua correxit me in finem et disciplina tua ipsa me docebit
PS|17|37|dilatasti gressus meos subtus me et non sunt infirmata vestigia mea
PS|17|38|persequar inimicos meos et conprehendam illos et non convertar donec deficiant
PS|17|39|confringam illos nec poterunt stare cadent subtus pedes meos
PS|17|40|et praecinxisti me virtute ad bellum subplantasti insurgentes in me subtus me
PS|17|41|et inimicos meos dedisti mihi dorsum et odientes me disperdisti
PS|17|42|clamaverunt nec erat qui salvos faceret ad Dominum nec exaudivit eos
PS|17|43|et comminuam illos ut pulverem ante faciem venti ut lutum platearum delebo eos
PS|17|44|eripe me de contradictionibus populi constitues me in caput gentium
PS|17|45|populus quem non cognovi servivit mihi in auditu auris oboedivit mihi
PS|17|46|filii alieni mentiti sunt mihi filii alieni inveterati sunt et claudicaverunt a semitis suis
PS|17|47|vivit Dominus et benedictus Deus meus et exaltetur Deus salutis meae
PS|17|48|Deus qui dat vindictas mihi et subdidit populos sub me liberator meus de gentibus iracundis
PS|17|49|et ab insurgentibus in me exaltabis me a viro iniquo eripies me
PS|17|50|propterea confitebor tibi in nationibus Domine et psalmum dicam nomini tuo
PS|17|51|magnificans salutes regis eius et faciens misericordiam christo suo David et semini eius usque in saeculum
PS|18|1|in finem psalmus David
PS|18|2|caeli enarrant gloriam Dei et opera manuum eius adnuntiat firmamentum
PS|18|3|dies diei eructat verbum et nox nocti indicat scientiam
PS|18|4|non sunt loquellae neque sermones quorum non audiantur voces eorum
PS|18|5|in omnem terram exivit sonus eorum et in fines orbis terrae verba eorum
PS|18|6|in sole posuit tabernaculum suum et ipse tamquam sponsus procedens de thalamo suo exultavit ut gigans ad currendam viam %suam;
PS|18|7|a summo caeli egressio eius et occursus eius usque ad summum eius nec est qui se abscondat a calore eius
PS|18|8|lex Domini inmaculata convertens animas testimonium Domini fidele sapientiam praestans parvulis
PS|18|9|iustitiae Domini rectae laetificantes corda praeceptum Domini lucidum inluminans oculos
PS|18|10|timor Domini sanctus permanens in saeculum saeculi iudicia Domini vera iustificata in semet ipsa
PS|18|11|desiderabilia super aurum et lapidem pretiosum multum et dulciora super mel et favum
PS|18|12|etenim servus tuus custodit ea in custodiendis illis retributio multa
PS|18|13|delicta quis intellegit ab occultis meis munda me
PS|18|14|et ab alienis parce servo tuo si mei non fuerint dominati tunc inmaculatus ero et emundabor a delicto maximo
PS|18|15|et erunt ut conplaceant eloquia oris mei et meditatio cordis mei in conspectu tuo semper Domine adiutor meus et redemptor meus
PS|19|1|in finem psalmus David
PS|19|2|exaudiat te Dominus in die tribulationis protegat te nomen Dei Iacob
PS|19|3|mittat tibi auxilium de sancto et de Sion tueatur te
PS|19|4|memor sit omnis sacrificii tui et holocaustum tuum pingue fiat diapsalma
PS|19|5|tribuat tibi secundum cor tuum et omne consilium tuum confirmet
PS|19|6|laetabimur in salutari tuo et in nomine Dei nostri magnificabimur
PS|19|7|impleat Dominus omnes petitiones tuas nunc cognovi quoniam salvum fecit Dominus christum suum exaudiet illum de caelo sancto suo in potentatibus salus dexterae eius
PS|19|8|hii in curribus et hii in equis nos autem in nomine Domini Dei nostri invocabimus
PS|19|9|ipsi obligati sunt et ceciderunt nos vero surreximus et erecti sumus
PS|19|10|Domine salvum fac regem et exaudi nos in die qua invocaverimus te
PS|20|1|in finem psalmus David
PS|20|2|Domine in virtute tua laetabitur rex et super salutare tuum exultabit vehementer
PS|20|3|desiderium animae eius tribuisti ei et voluntate labiorum eius non fraudasti eum diapsalma
PS|20|4|quoniam praevenisti eum in benedictionibus dulcedinis posuisti in capite eius coronam de lapide pretioso
PS|20|5|vitam petiit a te et tribuisti ei longitudinem dierum in saeculum et in saeculum saeculi
PS|20|6|magna gloria eius in salutari tuo gloriam et magnum decorem inpones super eum
PS|20|7|quoniam dabis eum benedictionem in saeculum saeculi laetificabis eum in gaudio cum vultu tuo
PS|20|8|quoniam rex sperat in Domino et in misericordia Altissimi non commovebitur
PS|20|9|inveniatur manus tua omnibus inimicis tuis dextera tua inveniat %omnes; qui te oderunt
PS|20|10|pones eos ut clibanum ignis in tempore vultus tui Dominus in ira sua conturbabit eos et devorabit eos ignis
PS|20|11|fructum eorum de terra perdes et semen eorum a filiis hominum
PS|20|12|quoniam declinaverunt in te mala cogitaverunt consilia quae non potuerunt %stabilire;
PS|20|13|quoniam pones eos dorsum in reliquis tuis praeparabis vultum eorum
PS|20|14|exaltare Domine in virtute tua cantabimus et psallemus virtutes tuas
PS|21|1|in finem pro adsumptione matutina psalmus David
PS|21|2|Deus Deus meus respice me; quare me dereliquisti longe a salute mea verba delictorum meorum
PS|21|3|Deus meus clamabo per diem et non exaudies et nocte et non ad insipientiam mihi
PS|21|4|tu autem in sancto habitas Laus Israhel
PS|21|5|in te speraverunt patres nostri speraverunt et liberasti eos
PS|21|6|ad te clamaverunt et salvi facti sunt in te speraverunt et non sunt confusi
PS|21|7|ego autem sum vermis et non homo obprobrium hominum et abiectio plebis
PS|21|8|omnes videntes me deriserunt me locuti sunt labiis moverunt caput
PS|21|9|speravit in Domino eripiat eum salvum faciat eum quoniam vult eum
PS|21|10|quoniam tu es qui extraxisti me de ventre spes mea ab uberibus matris meae
PS|21|11|in te proiectus sum ex utero de ventre matris meae Deus meus es tu
PS|21|12|ne discesseris a me quoniam tribulatio proxima est quoniam non est qui adiuvet
PS|21|13|circumdederunt me vituli multi tauri pingues obsederunt me
PS|21|14|aperuerunt super me os suum sicut leo rapiens et rugiens
PS|21|15|sicut aqua effusus sum et dispersa sunt universa ossa mea factum est cor meum tamquam cera liquescens in medio ventris mei
PS|21|16|aruit tamquam testa virtus mea et lingua mea adhesit faucibus meis et in limum mortis deduxisti me
PS|21|17|quoniam circumdederunt me canes multi concilium malignantium obsedit me foderunt manus meas et pedes meos
PS|21|18|dinumeraverunt omnia ossa mea ipsi vero consideraverunt et inspexerunt me
PS|21|19|diviserunt sibi vestimenta mea et super vestem meam miserunt sortem
PS|21|20|tu autem Domine ne elongaveris auxilium tuum ad defensionem meam conspice
PS|21|21|erue a framea animam meam et de manu canis unicam meam
PS|21|22|salva me ex ore leonis et a cornibus unicornium humilitatem meam
PS|21|23|narrabo nomen tuum fratribus meis in media ecclesia laudabo te
PS|21|24|qui timetis Dominum laudate eum universum semen Iacob magnificate eum
PS|21|25|timeat eum omne semen Israhel quoniam non sprevit neque dispexit deprecationem pauperis nec avertit faciem suam a me et cum clamarem ad eum exaudivit %me;
PS|21|26|apud te laus mea in ecclesia magna vota mea reddam in conspectu timentium eum
PS|21|27|edent pauperes et saturabuntur et laudabunt Dominum qui requirunt eum vivent corda eorum in saeculum saeculi
PS|21|28|reminiscentur et convertentur ad Dominum universi fines terrae et adorabunt in conspectu eius universae familiae gentium
PS|21|29|quoniam Dei est regnum et %ipse; dominabitur gentium
PS|21|30|manducaverunt et adoraverunt omnes pingues terrae in conspectu eius cadent omnes qui descendunt in terram
PS|21|31|et anima mea illi vivet et semen meum serviet ipsi
PS|21|32|adnuntiabitur Domino generatio ventura et adnuntiabunt iustitiam eius populo qui nascetur quem fecit %Dominus;
PS|22|1|psalmus David Dominus reget me et nihil mihi deerit
PS|22|2|in loco pascuae %ibi; me conlocavit super aquam refectionis educavit me
PS|22|3|animam meam convertit deduxit me super semitas iustitiae propter nomen suum
PS|22|4|nam et si ambulavero in medio umbrae mortis non timebo mala quoniam tu mecum es virga tua et baculus tuus ipsa me consolata sunt
PS|22|5|parasti in conspectu meo mensam adversus eos qui tribulant me inpinguasti in oleo caput meum et calix meus inebrians quam praeclarus est
PS|22|6|et misericordia tua subsequitur me omnibus diebus vitae meae et ut inhabitem in domo Domini in longitudinem dierum
PS|23|1|psalmus David prima sabbati Domini est terra et plenitudo eius orbis terrarum et %universi; qui habitant in eo
PS|23|2|quia; ipse super maria fundavit eum et super flumina praeparavit eum
PS|23|3|quis ascendit in montem Domini aut quis stabit in loco sancto eius
PS|23|4|innocens manibus et mundo corde qui non accepit in vano animam suam nec iuravit in dolo proximo suo
PS|23|5|hic accipiet benedictionem a Domino et misericordiam a Deo salvatore suo
PS|23|6|haec est generatio quaerentium eum quaerentium faciem Dei Iacob diapsalma
PS|23|7|adtollite portas principes vestras et elevamini portae aeternales et introibit rex gloriae
PS|23|8|quis est iste rex gloriae Dominus fortis et potens Dominus potens in proelio
PS|23|9|adtollite portas principes vestras et elevamini portae aeternales et introibit rex gloriae
PS|23|10|quis est iste rex gloriae Dominus virtutum ipse est rex gloriae diapsalma
PS|24|1|psalmus David ad te Domine levavi animam meam
PS|24|2|Deus meus in te confido non erubescam
PS|24|3|neque inrideant me inimici mei etenim universi qui sustinent te non confundentur
PS|24|4|confundantur %omnes; iniqua agentes supervacue vias tuas Domine demonstra mihi %et; semitas tuas doce me
PS|24|5|dirige me in veritatem tuam et doce me quoniam tu es Deus salvator meus et te sustinui tota die
PS|24|6|reminiscere miserationum tuarum Domine et misericordiarum tuarum quia a saeculo sunt
PS|24|7|delicta iuventutis meae et ignorantias meas ne memineris secundum misericordiam tuam memento mei tu; propter bonitatem tuam Domine
PS|24|8|dulcis et rectus Dominus propter hoc legem dabit delinquentibus in via
PS|24|9|diriget mansuetos in iudicio docebit mites vias suas
PS|24|10|universae viae Domini misericordia et veritas requirentibus testamentum eius et testimonia eius
PS|24|11|propter nomen tuum Domine et propitiaberis peccato meo multum est enim
PS|24|12|quis est homo qui timet Dominum legem statuet ei in via quam elegit
PS|24|13|anima eius in bonis demorabitur et semen ipsius hereditabit terram
PS|24|14|firmamentum est Dominus timentibus eum et testamentum ipsius ut manifestetur illis
PS|24|15|oculi mei semper ad Dominum quoniam ipse evellet de laqueo pedes meos
PS|24|16|respice in me et miserere mei quia unicus et pauper sum ego
PS|24|17|tribulationes cordis mei multiplicatae sunt de necessitatibus meis erue me
PS|24|18|vide humilitatem meam et laborem meum et dimitte universa delicta mea
PS|24|19|respice inimicos meos quoniam multiplicati sunt et odio iniquo oderunt me
PS|24|20|custodi animam meam et erue me non erubescam quoniam speravi in te
PS|24|21|innocentes et recti adheserunt mihi quia sustinui te
PS|24|22|libera Deus Israhel ex omnibus tribulationibus suis
PS|25|1|psalmus David iudica me Domine quoniam ego in innocentia mea ingressus sum et in Domino sperans non infirmabor
PS|25|2|proba me Domine et tempta me ure renes meos et cor meum
PS|25|3|quoniam misericordia tua ante oculos meos est et conplacui in veritate tua
PS|25|4|non sedi cum concilio vanitatis et cum iniqua gerentibus non introibo
PS|25|5|odivi ecclesiam malignantium et cum impiis non sedebo
PS|25|6|lavabo inter innocentes manus meas et circumdabo altare tuum Domine
PS|25|7|ut audiam vocem laudis et enarrem universa mirabilia tua
PS|25|8|Domine dilexi decorem domus tuae et locum habitationis gloriae tuae
PS|25|9|ne perdas cum impiis animam meam et cum viris sanguinum vitam meam
PS|25|10|in quorum manibus iniquitates sunt dextera eorum repleta est muneribus
PS|25|11|ego autem in innocentia mea ingressus sum redime me et miserere mei
PS|25|12|pes meus stetit in directo in ecclesiis benedicam %te; Domine
PS|26|1|David priusquam liniretur Dominus inluminatio mea et salus mea quem timebo Dominus protector vitae meae a quo trepidabo
PS|26|2|dum adpropiant super me nocentes ut edant carnes meas qui tribulant me et inimici mei ipsi infirmati sunt et ceciderunt
PS|26|3|si consistant adversus me castra non timebit cor meum si exsurgat adversus me proelium in hoc ego sperabo
PS|26|4|unam petii a Domino hanc requiram ut inhabitem in domo Domini omnes dies vitae meae ut videam voluntatem Domini et visitem templum eius
PS|26|5|quoniam abscondit me in tabernaculo in die malorum protexit me in abscondito tabernaculi sui
PS|26|6|in petra exaltavit me et nunc exaltavit caput meum super inimicos meos circuivi et immolavi in tabernaculo eius hostiam vociferationis cantabo et psalmum dicam Domino
PS|26|7|exaudi Domine vocem meam qua clamavi miserere mei et exaudi me
PS|26|8|tibi dixit cor meum exquisivit facies mea faciem tuam Domine requiram
PS|26|9|ne avertas faciem tuam a me ne declines in ira a servo tuo adiutor meus esto ne derelinquas me neque dispicias me Deus salvator meus
PS|26|10|quoniam pater meus et mater mea dereliquerunt me Dominus autem adsumpsit me
PS|26|11|legem pone mihi Domine in via tua et dirige me in semita recta propter inimicos meos
PS|26|12|ne tradideris me in animas tribulantium me quoniam insurrexerunt in me testes iniqui et mentita est iniquitas sibi
PS|26|13|credo videre bona Domini in terra viventium
PS|26|14|expecta Dominum viriliter age et confortetur cor tuum et sustine Dominum
PS|27|1|huic David ad te Domine clamabo Deus meus ne sileas a me nequando taceas a me et adsimilabor descendentibus in lacum
PS|27|2|exaudi vocem deprecationis meae dum oro ad te dum extollo manus meas ad templum sanctum tuum
PS|27|3|ne simul tradas me cum peccatoribus et cum operantibus iniquitatem %ne perdideris me; qui loquuntur pacem cum proximo suo mala autem sunt in cordibus eorum
PS|27|4|da illis secundum opera ipsorum et secundum nequitiam adinventionum ipsorum secundum opera manuum eorum tribue illis redde retributionem eorum ipsis
PS|27|5|quoniam non intellexerunt opera Domini et in opera manuum eius destrues illos et non aedificabis eos
PS|27|6|benedictus Dominus quoniam exaudivit vocem deprecationis meae
PS|27|7|Dominus adiutor meus et protector meus in ipso speravit cor meum et adiutus sum et refloruit caro mea et ex voluntate mea confitebor ei
PS|27|8|Dominus fortitudo plebis suae et protector salvationum christi sui est
PS|27|9|salvam fac plebem tuam et benedic hereditati tuae et rege eos et extolle eos usque in aeternum
PS|28|1|psalmus David in consummatione tabernaculi adferte Domino filii Dei adferte Domino filios arietum
PS|28|2|adferte Domino gloriam et honorem adferte Domino gloriam nomini eius adorate Dominum in atrio sancto eius
PS|28|3|vox Domini super aquas Deus maiestatis intonuit Dominus super aquas multas
PS|28|4|vox Domini in virtute vox Domini in magnificentia
PS|28|5|vox Domini confringentis cedros et confringet Dominus cedros Libani
PS|28|6|et comminuet eas tamquam vitulum Libani et dilectus quemadmodum filius unicornium
PS|28|7|vox Domini intercidentis flammam ignis
PS|28|8|vox Domini concutientis desertum et commovebit Dominus desertum Cades
PS|28|9|vox Domini praeparantis cervos et revelabit condensa et in templo eius omnis dicet gloriam
PS|28|10|Dominus diluvium inhabitare facit et sedebit Dominus rex in aeternum
PS|28|11|Dominus virtutem populo suo dabit Dominus benedicet populo suo in pace
PS|29|1|psalmus cantici in dedicatione domus David
PS|29|2|exaltabo te Domine quoniam suscepisti me nec delectasti inimicos meos super me
PS|29|3|Domine Deus meus clamavi ad te et sanasti me
PS|29|4|Domine eduxisti ab inferno animam meam salvasti me a descendentibus in lacum
PS|29|5|psallite Domino sancti eius et confitemini memoriae sanctitatis eius
PS|29|6|quoniam ira in indignatione eius et vita in voluntate eius ad vesperum demorabitur fletus et ad matutinum laetitia
PS|29|7|ego autem dixi in abundantia mea non movebor in aeternum
PS|29|8|Domine in voluntate tua praestitisti decori meo virtutem avertisti faciem tuam et factus sum conturbatus
PS|29|9|ad te Domine clamabo et ad Deum meum deprecabor
PS|29|10|quae utilitas in sanguine meo dum descendo in corruptionem numquid confitebitur tibi pulvis aut adnuntiabit veritatem tuam
PS|29|11|audivit Dominus et misertus est mei Dominus factus est adiutor meus
PS|29|12|convertisti planctum meum in gaudium mihi conscidisti saccum meum et circumdedisti me laetitia
PS|29|13|ut cantet tibi gloria mea et non conpungar Domine Deus meus in aeternum confitebor tibi
PS|30|1|in finem psalmus David
PS|30|2|in te Domine speravi non confundar in aeternum in iustitia tua libera me
PS|30|3|inclina ad me aurem tuam adcelera ut eruas me esto mihi in Deum protectorem et in domum refugii ut salvum me facias
PS|30|4|quoniam fortitudo mea et refugium meum es tu et propter nomen tuum deduces me et enutries me
PS|30|5|educes me de laqueo hoc quem absconderunt mihi quoniam tu es protector meus
PS|30|6|in manus tuas commendabo spiritum meum redemisti me Domine Deus veritatis
PS|30|7|odisti observantes vanitates supervacue ego autem in Domino speravi
PS|30|8|exultabo et laetabor in misericordia tua quoniam respexisti humilitatem meam salvasti de necessitatibus animam meam
PS|30|9|nec conclusisti me in manibus inimici statuisti in loco spatioso pedes meos
PS|30|10|miserere mei Domine quoniam tribulor conturbatus est in ira oculus meus anima mea et venter meus
PS|30|11|quoniam defecit in dolore vita mea et anni mei in gemitibus infirmata est in paupertate virtus mea et ossa mea conturbata sunt
PS|30|12|super omnes inimicos meos factus sum obprobrium et vicinis meis valde et timor notis meis qui videbant me foras fugerunt a me
PS|30|13|oblivioni datus sum tamquam mortuus a corde factus sum tamquam vas perditum
PS|30|14|quoniam audivi vituperationem multorum commorantium in circuitu in eo dum convenirent simul adversus me accipere animam meam consiliati sunt
PS|30|15|ego autem in te speravi Domine dixi Deus meus es tu
PS|30|16|in manibus tuis sortes meae eripe me de manu inimicorum meorum et a persequentibus me
PS|30|17|inlustra faciem tuam super servum tuum salvum me fac in misericordia tua
PS|30|18|Domine ne confundar quoniam invocavi te erubescant impii et deducantur in infernum
PS|30|19|muta fiant labia dolosa quae loquuntur adversus iustum iniquitatem in superbia et in abusione
PS|30|20|quam magna multitudo dulcedinis tuae %Domine; quam abscondisti timentibus te perfecisti eis qui sperant in te in conspectu filiorum hominum
PS|30|21|abscondes eos in abdito faciei tuae a conturbatione hominum proteges eos in tabernaculo a contradictione linguarum
PS|30|22|benedictus Dominus quoniam mirificavit misericordiam suam mihi in civitate munita
PS|30|23|ego autem dixi in excessu mentis meae proiectus sum a facie oculorum tuorum ideo exaudisti vocem orationis meae dum clamarem ad te
PS|30|24|diligite Dominum omnes sancti eius %quoniam; veritates requirit Dominus et retribuit abundanter facientibus superbiam
PS|30|25|viriliter agite et confortetur cor vestrum omnes qui speratis in Domino
PS|31|1|huic David intellectus beati quorum remissae sunt iniquitates et quorum tecta sunt peccata
PS|31|2|beatus vir cui non inputabit Dominus peccatum nec est in spiritu eius dolus
PS|31|3|quoniam tacui inveteraverunt ossa mea dum clamarem tota die
PS|31|4|quoniam die ac nocte gravata est super me manus tua conversus sum in aerumna mea; dum configitur %mihi; spina diapsalma
PS|31|5|delictum meum cognitum tibi; feci et iniustitiam meam non abscondi dixi confitebor adversus me iniustitiam meam Domino et tu remisisti impietatem peccati mei diapsalma
PS|31|6|pro hac orabit ad te omnis sanctus in tempore oportuno verumtamen in diluvio aquarum multarum ad eum non adproximabunt
PS|31|7|tu es refugium meum a tribulatione quae circumdedit me exultatio mea erue me a circumdantibus me diapsalma
PS|31|8|intellectum tibi dabo et instruam te in via hac qua gradieris firmabo super te oculos meos
PS|31|9|nolite fieri sicut equus et mulus quibus non est intellectus in camo et freno maxillas eorum constringe qui non adproximant ad te
PS|31|10|multa flagella peccatoris sperantem autem in Domino misericordia circumdabit
PS|31|11|laetamini in Domino et exultate iusti et gloriamini omnes recti corde
PS|32|1|psalmus David exultate iusti in Domino rectos decet laudatio
PS|32|2|confitemini Domino in cithara in psalterio decem cordarum psallite illi
PS|32|3|cantate ei canticum novum bene psallite in vociferatione
PS|32|4|quia rectum est verbum Domini et omnia opera eius in fide
PS|32|5|diligit misericordiam et iudicium misericordia Domini plena est terra
PS|32|6|verbo Domini caeli firmati sunt et spiritu oris eius omnis virtus eorum
PS|32|7|congregans sicut in utre aquas maris ponens in thesauris abyssos
PS|32|8|timeat Dominum omnis terra ab eo autem commoveantur omnes inhabitantes orbem
PS|32|9|quoniam ipse dixit et facta sunt ipse mandavit et creata sunt
PS|32|10|Dominus dissipat consilia gentium reprobat autem cogitationes populorum %et reprobat consilia principum;
PS|32|11|consilium autem Domini in aeternum manet cogitationes cordis eius in generatione et generationem
PS|32|12|beata gens cuius est Dominus Deus eius populus quem elegit in hereditatem sibi
PS|32|13|de caelo respexit Dominus vidit omnes filios hominum
PS|32|14|de praeparato habitaculo suo respexit super omnes qui habitant terram
PS|32|15|qui finxit singillatim corda eorum qui intellegit omnia opera illorum
PS|32|16|non salvatur rex per multam virtutem et gigans non salvabitur in multitudine virtutis suae
PS|32|17|fallax equus ad salutem in abundantia autem virtutis suae non salvabitur
PS|32|18|ecce oculi Domini super metuentes eum qui sperant super misericordia eius
PS|32|19|ut eruat a morte animas eorum et alat eos in fame
PS|32|20|anima nostra sustinet Dominum quoniam adiutor et protector noster est
PS|32|21|quia in eo laetabitur cor nostrum et in nomine sancto eius speravimus
PS|32|22|fiat misericordia tua Domine super nos quemadmodum speravimus in te
PS|33|1|David cum inmutavit vultum suum coram Abimelech et dimisit eum et abiit
PS|33|2|benedicam Dominum in omni tempore semper laus eius in ore meo
PS|33|3|in Domino laudabitur anima mea audiant mansueti et laetentur
PS|33|4|magnificate Dominum mecum et exaltemus nomen eius in id ipsum
PS|33|5|exquisivi Dominum et exaudivit me et ex omnibus tribulationibus meis eripuit me
PS|33|6|accedite ad eum et inluminamini et facies vestrae non confundentur
PS|33|7|iste pauper clamavit et Dominus exaudivit %eum; et de omnibus tribulationibus eius salvavit eum
PS|33|8|vallabit angelus Domini in circuitu timentium eum et eripiet eos
PS|33|9|gustate et videte quoniam suavis est Dominus beatus vir qui sperat in eo
PS|33|10|timete Dominum %omnes; sancti eius quoniam non est inopia timentibus eum
PS|33|11|divites eguerunt et esurierunt inquirentes autem Dominum non minuentur omni bono diapsalma
PS|33|12|venite filii audite me timorem Domini docebo vos
PS|33|13|quis est homo qui vult vitam cupit videre dies bonos
PS|33|14|prohibe linguam tuam a malo et labia tua ne loquantur dolum
PS|33|15|deverte a malo et fac bonum inquire pacem et persequere eam
PS|33|16|oculi Domini super iustos et aures eius in precem eorum
PS|33|17|facies Domini super facientes mala ut perdat de terra memoriam eorum
PS|33|18|clamaverunt iusti et Dominus exaudivit et ex omnibus tribulationibus eorum liberavit eos
PS|33|19|iuxta est Dominus his qui tribulato sunt corde et humiles spiritu salvabit
PS|33|20|multae tribulationes iustorum et de omnibus his liberavit eos
PS|33|21|Dominus custodit omnia ossa eorum unum ex his non conteretur
PS|33|22|mors peccatorum pessima et qui oderunt iustum delinquent
PS|33|23|redimet Dominus animas servorum suorum et non delinquent omnes qui sperant in eum
PS|34|1|huic David iudica Domine nocentes me expugna expugnantes me
PS|34|2|adprehende arma et scutum et exsurge in adiutorium mihi
PS|34|3|effunde frameam et conclude adversus eos qui persequuntur me dic animae meae salus tua ego sum
PS|34|4|confundantur et revereantur quaerentes animam meam avertantur retrorsum et confundantur cogitantes mihi mala
PS|34|5|fiant tamquam pulvis ante faciem venti et angelus Domini coartans eos
PS|34|6|fiat via illorum tenebrae et lubricum et angelus Domini persequens eos
PS|34|7|quoniam gratis absconderunt mihi interitum laquei sui supervacue exprobraverunt animam meam
PS|34|8|veniat illi laqueus quem ignorat et captio quam abscondit conprehendat eum et in laqueo cadat in ipso
PS|34|9|anima autem mea exultabit in Domino delectabitur super salutari suo
PS|34|10|omnia ossa mea dicent Domine quis similis tui eripiens inopem de manu fortiorum eius egenum et pauperem a diripientibus eum
PS|34|11|surgentes testes iniqui quae ignorabam interrogabant me
PS|34|12|retribuebant mihi mala pro bonis sterilitatem animae meae
PS|34|13|ego autem cum mihi molesti essent induebar cilicio humiliabam in ieiunio animam meam et oratio mea in sinum meum convertetur
PS|34|14|quasi proximum quasi fratrem nostrum sic conplacebam quasi lugens et contristatus sic humiliabar
PS|34|15|et adversum me laetati sunt et convenerunt congregata sunt super me flagella et ignoravi
PS|34|16|dissipati sunt nec conpuncti temptaverunt me subsannaverunt me subsannatione frenduerunt super me dentibus suis
PS|34|17|Domine quando respicies restitue animam meam a malignitate eorum a leonibus unicam meam
PS|34|18|confitebor tibi in ecclesia magna in populo gravi laudabo te
PS|34|19|non supergaudeant mihi qui adversantur mihi inique qui oderunt me gratis et annuunt oculis
PS|34|20|quoniam mihi quidem pacifice loquebantur et in iracundia terrae loquentes; dolos cogitabant
PS|34|21|et dilataverunt super me os suum dixerunt euge euge viderunt oculi nostri
PS|34|22|vidisti Domine ne sileas Domine ne discedas a me
PS|34|23|exsurge et intende iudicio meo Deus meus et Dominus meus in causam meam
PS|34|24|iudica me secundum iustitiam tuam Domine Deus meus et non supergaudeant mihi
PS|34|25|non dicant in cordibus suis euge euge animae nostrae nec dicant devoravimus eum
PS|34|26|erubescant et revereantur simul qui gratulantur malis meis induantur confusione et reverentia qui magna loquuntur super me
PS|34|27|exultent et laetentur qui volunt iustitiam meam et dicant semper magnificetur Dominus qui volunt pacem servi eius
PS|34|28|et lingua mea meditabitur iustitiam tuam tota die laudem tuam
PS|35|1|in finem servo Domini David
PS|35|2|dixit iniustus ut delinquat in semet ipso non est timor Dei ante oculos eius
PS|35|3|quoniam dolose egit in conspectu eius ut inveniatur iniquitas eius ad odium
PS|35|4|verba oris eius iniquitas et dolus noluit intellegere ut bene ageret
PS|35|5|iniquitatem meditatus est in cubili suo adstetit omni viae non bonae malitiam autem non odivit
PS|35|6|Domine in caelo misericordia tua et veritas tua usque ad nubes
PS|35|7|iustitia tua sicut montes Dei iudicia tua abyssus multa homines et iumenta salvabis Domine
PS|35|8|quemadmodum multiplicasti misericordiam tuam Deus filii autem hominum in tegmine alarum tuarum sperabunt
PS|35|9|inebriabuntur ab ubertate domus tuae et torrente voluntatis tuae potabis eos
PS|35|10|quoniam apud te fons vitae in lumine tuo videbimus lumen
PS|35|11|praetende misericordiam tuam scientibus te et iustitiam tuam his qui recto sunt corde
PS|35|12|non veniat mihi pes superbiae et manus peccatoris non moveat me
PS|35|13|ibi ceciderunt qui operantur iniquitatem expulsi sunt nec potuerunt stare
PS|36|1|ipsi David noli aemulari in malignantibus neque zelaveris facientes iniquitatem
PS|36|2|quoniam tamquam faenum velociter arescent et quemadmodum holera herbarum cito decident
PS|36|3|spera in Domino et fac bonitatem et inhabita terram et pasceris in divitiis eius
PS|36|4|delectare in Domino et dabit tibi petitiones cordis tui
PS|36|5|revela Domino viam tuam et spera in eum et ipse faciet
PS|36|6|et educet quasi lumen iustitiam tuam et iudicium tuum tamquam meridiem
PS|36|7|subditus esto Domino et ora eum noli aemulari in eo qui prosperatur in via sua in homine faciente iniustitias
PS|36|8|desine ab ira et derelinque furorem noli aemulari ut maligneris
PS|36|9|quoniam qui malignantur exterminabuntur sustinentes autem Dominum ipsi hereditabunt terram
PS|36|10|et adhuc pusillum et non erit peccator et quaeres locum eius et non invenies
PS|36|11|mansueti autem hereditabunt terram et delectabuntur in multitudine pacis
PS|36|12|observabit peccator iustum et stridebit super eum dentibus suis
PS|36|13|Dominus autem inridebit eum quia prospicit quoniam veniet dies eius
PS|36|14|gladium evaginaverunt peccatores intenderunt arcum suum ut decipiant pauperem et inopem ut trucident rectos corde
PS|36|15|gladius eorum intret in corda ipsorum et arcus ipsorum confringatur
PS|36|16|melius est modicum iusto super divitias peccatorum multas
PS|36|17|quoniam brachia peccatorum conterentur confirmat autem iustos Dominus
PS|36|18|novit Dominus dies inmaculatorum et hereditas eorum in aeternum erit
PS|36|19|non confundentur in tempore malo et in diebus famis saturabuntur
PS|36|20|quia peccatores peribunt inimici vero Domini mox honorificati fuerint et exaltati deficientes quemadmodum fumus defecerunt
PS|36|21|mutuabitur peccator et non solvet iustus autem miseretur et tribuet
PS|36|22|quia benedicentes ei hereditabunt terram maledicentes autem ei disperibunt
PS|36|23|apud Dominum gressus hominis dirigentur et viam eius volet
PS|36|24|cum ceciderit non conlidetur quia Dominus subponit manum suam
PS|36|25|iunior fui et senui et non vidi iustum derelictum nec semen eius quaerens panes
PS|36|26|tota die miseretur et commodat et semen illius in benedictione erit
PS|36|27|declina a malo et fac bonum et inhabita in saeculum saeculi
PS|36|28|quia Dominus amat iudicium et non derelinquet sanctos suos in aeternum conservabuntur iniusti punientur et semen impiorum peribit
PS|36|29|iusti autem hereditabunt terram et inhabitabunt in saeculum %saeculi; super eam
PS|36|30|os iusti meditabitur sapientiam et lingua eius loquetur iudicium
PS|36|31|lex Dei eius in corde ipsius et non subplantabuntur gressus eius
PS|36|32|considerat peccator iustum et quaerit mortificare eum
PS|36|33|Dominus autem non derelinquet eum in manus eius nec damnabit eum cum iudicabitur illi
PS|36|34|expecta Dominum et custodi viam eius et exaltabit te ut hereditate capias terram cum perierint peccatores videbis
PS|36|35|vidi impium superexaltatum et elevatum sicut cedros Libani
PS|36|36|et transivi et ecce non erat et quaesivi eum et non est inventus locus eius
PS|36|37|custodi innocentiam et vide aequitatem quoniam sunt reliquiae homini pacifico
PS|36|38|iniusti autem disperibunt simul reliquiae impiorum peribunt
PS|36|39|salus autem iustorum a Domino et protector eorum in tempore tribulationis
PS|36|40|et adiuvabit eos Dominus et liberabit eos et eruet eos a peccatoribus et salvabit eos quia speraverunt in eo
PS|37|1|psalmus David in rememorationem de sabbato
PS|37|2|Domine ne in furore tuo arguas me neque in ira tua corripias me
PS|37|3|quoniam sagittae tuae infixae sunt mihi et confirmasti super me manum tuam
PS|37|4|non est sanitas carni meae a facie irae tuae non est pax ossibus meis a facie peccatorum meorum
PS|37|5|quoniam iniquitates meae supergressae sunt caput meum sicut onus grave gravatae sunt super me
PS|37|6|putruerunt et corruptae sunt cicatrices meae a facie insipientiae meae
PS|37|7|miser factus sum et curvatus sum usque ad finem tota die contristatus ingrediebar
PS|37|8|quoniam lumbi mei impleti sunt inlusionibus et non est sanitas in carne mea
PS|37|9|adflictus sum et humiliatus sum nimis rugiebam a gemitu cordis mei
PS|37|10|Domine ante te omne desiderium meum et gemitus meus a te non est absconditus
PS|37|11|cor meum conturbatum est dereliquit me virtus mea et lumen oculorum meorum et ipsum non est mecum
PS|37|12|amici mei et proximi mei adversus me adpropinquaverunt et steterunt et qui iuxta me erant de longe steterunt
PS|37|13|et vim faciebant qui quaerebant animam meam et qui inquirebant mala mihi locuti sunt vanitates et dolos tota die meditabantur
PS|37|14|ego autem tamquam surdus non audiebam et sicut mutus non aperiens os suum
PS|37|15|et factus sum sicut homo non audiens et non habens in ore suo redargutiones
PS|37|16|quoniam in te Domine speravi tu exaudies Domine Deus meus
PS|37|17|quia dixi nequando supergaudeant mihi inimici mei et dum commoventur pedes mei super me magna locuti sunt
PS|37|18|quoniam ego in flagella paratus et dolor meus in conspectu meo semper
PS|37|19|quoniam iniquitatem meam adnuntiabo %et; cogitabo pro peccato meo
PS|37|20|inimici autem mei vivent et firmati sunt super me et multiplicati sunt qui oderunt me inique
PS|37|21|qui retribuunt mala pro bonis detrahebant mihi quoniam sequebar bonitatem
PS|37|22|non derelinquas me Domine Deus meus ne discesseris a me
PS|37|23|intende in adiutorium meum Domine salutis meae
PS|38|1|in finem Idithun canticum David
PS|38|2|dixi custodiam vias meas ut non delinquam in lingua mea posui ori meo custodiam cum consisteret peccator adversum me
PS|38|3|obmutui et humiliatus sum et silui a bonis et dolor meus renovatus est
PS|38|4|concaluit cor meum intra me et in meditatione mea exardescet ignis
PS|38|5|locutus sum in lingua mea notum fac mihi Domine finem meum et numerum dierum meorum quis est ut sciam quid desit mihi
PS|38|6|ecce mensurabiles posuisti dies meos et substantia mea tamquam nihilum ante te verumtamen universa vanitas omnis homo vivens diapsalma
PS|38|7|verumtamen in imagine pertransit homo sed et frustra conturbatur thesaurizat et ignorat cui congregabit ea
PS|38|8|et nunc quae est expectatio mea nonne Dominus et substantia mea apud te est
PS|38|9|ab omnibus iniquitatibus meis erue me obprobrium insipienti dedisti me
PS|38|10|obmutui %et; non aperui os meum quoniam tu fecisti
PS|38|11|amove a me plagas tuas
PS|38|12|a fortitudine manus tuae ego defeci in increpationibus propter iniquitatem corripuisti hominem et tabescere fecisti sicut araneam animam eius verumtamen vane %conturbatur; omnis homo diapsalma
PS|38|13|exaudi orationem meam Domine et deprecationem meam auribus percipe lacrimas meas ne sileas quoniam advena sum apud te et peregrinus sicut omnes patres mei
PS|38|14|remitte mihi ut refrigerer priusquam abeam et amplius non ero
PS|39|1|in finem David psalmus
PS|39|2|expectans expectavi Dominum et intendit mihi
PS|39|3|et exaudivit preces meas et eduxit me de lacu miseriae et de luto fecis et statuit super petram pedes meos et direxit gressus meos
PS|39|4|et inmisit in os meum canticum novum carmen Deo nostro videbunt multi et timebunt et sperabunt in Domino
PS|39|5|beatus vir cuius est nomen Domini spes ipsius et non respexit in vanitates et insanias falsas
PS|39|6|multa fecisti tu Domine Deus meus mirabilia tua et cogitationibus tuis non est qui similis sit tibi adnuntiavi et locutus sum multiplicati sunt super numerum
PS|39|7|sacrificium et oblationem noluisti aures autem perfecisti mihi holocaustum et pro peccato non postulasti
PS|39|8|tunc dixi ecce venio in capite libri scriptum est de me
PS|39|9|ut facerem voluntatem tuam Deus meus volui et legem tuam in medio cordis mei
PS|39|10|adnuntiavi iustitiam in ecclesia magna ecce labia mea non prohibebo Domine tu scisti
PS|39|11|iustitiam tuam non abscondi in corde meo veritatem tuam et salutare tuum dixi non abscondi misericordiam tuam et veritatem tuam a concilio multo
PS|39|12|tu autem Domine ne longe facias miserationes tuas a me misericordia tua et veritas tua semper susceperunt me
PS|39|13|quoniam circumdederunt me mala quorum non est numerus conprehenderunt me iniquitates meae et non potui ut viderem multiplicatae sunt super capillos capitis mei et cor meum dereliquit me
PS|39|14|conplaceat tibi Domine ut eruas me Domine ad adiuvandum me respice
PS|39|15|confundantur et revereantur simul qui quaerunt animam meam ut auferant eam convertantur retrorsum et revereantur qui volunt mihi mala
PS|39|16|ferant confestim confusionem suam qui dicunt mihi euge euge
PS|39|17|exultent et laetentur super te omnes quaerentes te et dicant semper magnificetur Dominus qui diligunt salutare tuum
PS|39|18|ego autem mendicus sum et pauper Dominus sollicitus est mei adiutor meus et protector meus tu es Deus meus ne tardaveris
PS|40|1|in finem psalmus David
PS|40|2|beatus qui intellegit super egenum et pauperem in die mala liberabit eum Dominus
PS|40|3|Dominus conservet eum et vivificet eum et beatum faciat eum in terra et non tradat eum in animam inimicorum eius
PS|40|4|Dominus opem ferat illi super lectum doloris eius universum stratum eius versasti in infirmitate eius
PS|40|5|ego dixi Domine miserere mei sana animam meam quoniam peccavi tibi
PS|40|6|inimici mei dixerunt mala mihi quando morietur et peribit nomen eius
PS|40|7|et si ingrediebatur ut videret vane loquebatur cor eius congregavit iniquitatem sibi egrediebatur foras et loquebatur
PS|40|8|in id ipsum adversum me susurrabant omnes inimici mei adversus me cogitabant mala mihi
PS|40|9|verbum iniquum constituerunt adversus me numquid qui dormit non adiciet ut resurgat
PS|40|10|etenim homo pacis meae in quo speravi qui edebat panes meos magnificavit super me subplantationem
PS|40|11|tu autem Domine miserere mei et resuscita me et retribuam eis
PS|40|12|in hoc cognovi quoniam voluisti me quoniam non gaudebit inimicus meus super me
PS|40|13|me autem propter innocentiam suscepisti et confirmasti me in conspectu tuo in aeternum
PS|40|14|benedictus Dominus Deus Israhel a saeculo et in saeculum fiat fiat
PS|41|1|in finem in intellectum filiis Core
PS|41|2|quemadmodum desiderat cervus ad fontes aquarum ita desiderat anima mea ad te Deus
PS|41|3|sitivit anima mea ad Deum fortem; vivum quando veniam et parebo ante faciem Dei
PS|41|4|fuerunt mihi lacrimae meae panis die ac nocte dum dicitur mihi cotidie ubi est Deus tuus
PS|41|5|haec recordatus sum et effudi in me animam meam quoniam transibo in loco tabernaculi admirabilis usque ad domum Dei in voce exultationis et confessionis sonus epulantis
PS|41|6|quare tristis es anima mea et quare conturbas me spera in Deo quoniam confitebor illi salutare vultus mei
PS|41|7|Deus meus ad me ipsum anima mea conturbata est propterea memor ero tui de terra Iordanis et Hermoniim a monte modico
PS|41|8|abyssus ad; abyssum invocat in voce cataractarum tuarum omnia excelsa tua et fluctus tui super me transierunt
PS|41|9|in die mandavit Dominus misericordiam suam et nocte canticum eius apud me oratio Deo vitae meae
PS|41|10|dicam Deo susceptor meus es quare oblitus es mei quare contristatus incedo dum adfligit me inimicus
PS|41|11|dum confringuntur ossa mea exprobraverunt mihi qui tribulant me dum dicunt mihi per singulos dies ubi est Deus tuus
PS|41|12|quare tristis es anima mea et quare conturbas me spera in Deum quoniam adhuc; confitebor illi salutare vultus mei et; Deus meus
PS|42|1|psalmus David iudica me Deus et discerne causam meam de gente non sancta ab homine iniquo et doloso erue me
PS|42|2|quia tu es Deus fortitudo mea quare me reppulisti quare tristis incedo dum adfligit me inimicus
PS|42|3|emitte lucem tuam et veritatem tuam ipsa me deduxerunt et adduxerunt in montem sanctum tuum et in tabernacula tua
PS|42|4|et introibo ad altare Dei ad Deum qui laetificat iuventutem meam confitebor tibi in cithara Deus Deus meus
PS|42|5|quare tristis es anima mea et quare conturbas me spera in Deum quoniam adhuc; confitebor illi salutare vultus mei et; Deus meus
PS|43|1|in finem filiis Core ad intellectum
PS|43|2|Deus auribus nostris audivimus patres nostri adnuntiaverunt nobis opus quod operatus es in diebus eorum in diebus antiquis
PS|43|3|manus tua gentes disperdit et plantasti eos adflixisti populos et expulisti eos
PS|43|4|nec enim in gladio suo possederunt terram et brachium eorum non salvavit eos sed dextera tua et brachium tuum et inluminatio faciei tuae quoniam conplacuisti in eis
PS|43|5|tu es ipse rex meus et Deus meus qui mandas salutes Iacob
PS|43|6|in te inimicos nostros ventilabimus cornu et in nomine tuo spernemus insurgentes in nobis
PS|43|7|non enim in arcu meo sperabo et gladius meus non salvabit me
PS|43|8|salvasti enim nos de adfligentibus nos et odientes nos confudisti
PS|43|9|in Deo laudabimur tota die et in nomine tuo confitebimur in saeculum diapsalma
PS|43|10|nunc autem reppulisti et confudisti nos et non egredieris in virtutibus nostris
PS|43|11|avertisti nos retrorsum post inimicos nostros et qui oderunt nos diripiebant sibi
PS|43|12|dedisti nos tamquam oves escarum et in gentibus dispersisti nos
PS|43|13|vendidisti populum tuum sine pretio et non fuit multitudo in commutationibus nostris
PS|43|14|posuisti nos obprobrium vicinis nostris subsannationem et derisum his qui in circuitu nostro
PS|43|15|posuisti nos in similitudinem gentibus commotionem capitis in populis
PS|43|16|tota die verecundia mea contra me est et confusio faciei meae cooperuit me
PS|43|17|a voce exprobrantis et obloquentis a facie inimici et persequentis
PS|43|18|haec omnia venerunt super nos nec obliti sumus te et inique non egimus in testamento tuo
PS|43|19|et non recessit retrorsum cor nostrum et declinasti semitas nostras a via tua
PS|43|20|quoniam humiliasti nos in loco adflictionis et cooperuit nos umbra mortis
PS|43|21|si obliti sumus nomen Dei nostri et %si; expandimus manus nostras ad deum alienum
PS|43|22|nonne Deus requiret ista ipse enim novit abscondita cordis quoniam propter te mortificamur omni die aestimati sumus sicut oves occisionis
PS|43|23|exsurge quare dormis Domine exsurge %et; ne repellas in finem
PS|43|24|quare faciem tuam avertis oblivisceris inopiae nostrae et tribulationis nostrae
PS|43|25|quoniam humiliata est in pulvere anima nostra conglutinatus est in terra venter noster
PS|43|26|exsurge adiuva nos et redime nos propter nomen tuum
PS|44|1|in finem pro his qui commutabuntur filiis Core ad intellectum canticum pro dilecto
PS|44|2|eructavit cor meum verbum bonum dico ego opera mea regi lingua mea calamus scribae velociter scribentis
PS|44|3|speciosus forma prae filiis hominum diffusa est gratia in labiis tuis propterea benedixit te Deus in aeternum
PS|44|4|accingere gladio tuo super femur tuum potentissime
PS|44|5|specie tua et pulchritudine tua et intende prospere procede et regna propter veritatem et mansuetudinem et iustitiam et deducet te mirabiliter dextera tua
PS|44|6|sagittae tuae acutae populi sub te cadent in corde inimicorum regis
PS|44|7|sedis tua Deus in saeculum saeculi virga directionis virga regni tui
PS|44|8|dilexisti iustitiam et odisti iniquitatem propterea unxit te Deus Deus tuus oleo laetitiae prae consortibus tuis
PS|44|9|murra et gutta et cassia a vestimentis tuis a domibus eburneis ex quibus delectaverunt te
PS|44|10|filiae regum in honore tuo adstetit regina a dextris tuis in vestitu deaurato circumdata varietate
PS|44|11|audi filia et vide et inclina aurem tuam et obliviscere populum tuum et domum patris tui
PS|44|12|et concupiscet rex decorem tuum quoniam ipse est dominus tuus et adorabunt eum
PS|44|13|et; filiae Tyri in muneribus vultum tuum deprecabuntur divites plebis
PS|44|14|omnis gloria eius filiae regis ab intus in fimbriis aureis
PS|44|15|circumamicta varietatibus adducentur regi virgines post eam proximae eius adferentur tibi
PS|44|16|adferentur in laetitia et exultatione adducentur in templum regis
PS|44|17|pro patribus tuis nati sunt tibi filii constitues eos principes super omnem terram
PS|44|18|memor ero nominis tui in omni generatione et generatione propterea populi confitebuntur tibi in aeternum et in saeculum saeculi
PS|45|1|in finem pro filiis Core pro arcanis psalmus
PS|45|2|Deus noster refugium et virtus adiutor in tribulationibus quae invenerunt nos nimis
PS|45|3|propterea non timebimus dum turbabitur terra et transferentur montes in cor maris
PS|45|4|sonaverunt et turbatae sunt aquae eorum conturbati sunt montes in fortitudine eius diapsalma
PS|45|5|fluminis impetus laetificat civitatem Dei sanctificavit tabernaculum suum Altissimus
PS|45|6|Deus in medio eius non commovebitur adiuvabit eam Deus mane diluculo
PS|45|7|conturbatae sunt gentes inclinata sunt regna dedit vocem suam mota est terra
PS|45|8|Dominus virtutum nobiscum susceptor noster Deus Iacob diapsalma
PS|45|9|venite et videte opera Domini quae posuit prodigia super terram
PS|45|10|auferens bella usque ad finem terrae arcum conteret et confringet arma et scuta conburet in igne
PS|45|11|vacate et videte quoniam ego sum Deus exaltabor in gentibus exaltabor in terra
PS|45|12|Dominus virtutum nobiscum susceptor noster Deus Iacob
PS|46|1|in finem pro filiis Core psalmus
PS|46|2|omnes gentes plaudite manibus iubilate Deo in voce exultationis
PS|46|3|quoniam Dominus excelsus terribilis rex magnus super omnem terram
PS|46|4|subiecit populos nobis et gentes sub pedibus nostris
PS|46|5|elegit nobis hereditatem suam speciem Iacob quam dilexit diapsalma
PS|46|6|ascendit Deus in iubilo Dominus in voce tubae
PS|46|7|psallite Deo nostro psallite psallite regi nostro psallite
PS|46|8|quoniam rex omnis terrae Deus psallite sapienter
PS|46|9|regnavit Deus super gentes Deus sedit super sedem sanctam suam
PS|46|10|principes populorum congregati sunt cum Deo Abraham quoniam Dei fortes terrae vehementer elevati sunt
PS|47|1|canticum psalmi filiis Core secunda sabbati
PS|47|2|magnus Dominus et laudabilis nimis in civitate Dei nostri in monte sancto eius
PS|47|3|fundatur exultatione universae terrae montes Sion latera aquilonis civitas regis magni
PS|47|4|Deus in domibus eius cognoscitur cum suscipiet eam
PS|47|5|quoniam ecce reges congregati sunt convenerunt in unum
PS|47|6|ipsi videntes sic admirati sunt conturbati sunt commoti sunt
PS|47|7|tremor adprehendit eos ibi dolores ut parturientis
PS|47|8|in spiritu vehementi conteres naves Tharsis
PS|47|9|sicut audivimus sic vidimus in civitate Domini virtutum in civitate Dei nostri Deus fundavit eam in aeternum diapsalma
PS|47|10|suscepimus Deus misericordiam tuam in medio templi tui
PS|47|11|secundum nomen tuum Deus sic et laus tua in fines terrae iustitia plena est dextera tua
PS|47|12|laetetur mons Sion exultent filiae Iudaeae propter iudicia tua %Domine;
PS|47|13|circumdate Sion et conplectimini eam narrate in turribus eius
PS|47|14|ponite corda vestra in virtute eius et distribuite domus eius ut enarretis in progeniem alteram
PS|47|15|quoniam hic est Deus Deus noster in aeternum et in saeculum saeculi ipse reget nos in saecula
PS|48|1|in finem filiis Core psalmus
PS|48|2|audite haec omnes gentes auribus percipite omnes qui habitatis orbem
PS|48|3|quique terriginae et filii hominum in unum dives et pauper
PS|48|4|os meum loquetur sapientiam et meditatio cordis mei prudentiam
PS|48|5|inclinabo in parabolam aurem meam aperiam in psalterio propositionem meam
PS|48|6|cur timebo in die malo iniquitas calcanei mei circumdabit me
PS|48|7|qui confidunt in virtute sua et in multitudine divitiarum suarum gloriantur
PS|48|8|frater non redimit redimet homo non dabit Deo placationem suam
PS|48|9|et pretium redemptionis animae suae et laboravit in aeternum
PS|48|10|et vivet adhuc; in finem
PS|48|11|non videbit interitum cum viderit sapientes morientes simul insipiens et stultus peribunt et relinquent alienis divitias suas
PS|48|12|%et; sepulchra eorum domus illorum in aeternum tabernacula eorum in progeniem et progeniem vocaverunt nomina sua in terris suis
PS|48|13|et homo cum in honore esset non intellexit conparatus est iumentis insipientibus et similis factus est illis
PS|48|14|haec via illorum scandalum ipsis et postea in ore suo conplacebunt diapsalma
PS|48|15|sicut oves in inferno positi sunt mors depascet eos et dominabuntur eorum iusti in matutino et auxilium eorum veterescet in inferno a gloria eorum
PS|48|16|verumtamen Deus redimet animam meam de manu inferi cum acceperit me diapsalma
PS|48|17|ne timueris cum dives factus fuerit homo et cum multiplicata fuerit gloria domus eius
PS|48|18|quoniam cum interierit non sumet omnia neque descendet cum eo pone; gloria eius
PS|48|19|quia anima eius in vita ipsius benedicetur confitebitur tibi cum benefeceris ei
PS|48|20|introibit usque in progenies patrum suorum usque in aeternum non videbit lumen
PS|48|21|homo in honore cum esset non intellexit conparatus est iumentis %insipientibus; et similis factus est illis
PS|49|1|psalmus Asaph Deus deorum Dominus locutus est et vocavit terram a solis ortu usque ad occasum
PS|49|2|ex Sion species decoris eius
PS|49|3|Deus manifeste veniet Deus noster et non silebit ignis in conspectu eius exardescet et in circuitu eius tempestas valida
PS|49|4|advocabit caelum desursum et terram discernere populum suum
PS|49|5|congregate illi sanctos eius qui ordinant testamentum eius super sacrificia
PS|49|6|et adnuntiabunt caeli iustitiam eius quoniam Deus iudex est diapsalma
PS|49|7|audi populus meus et loquar tibi Israhel et testificabor tibi Deus Deus tuus ego sum
PS|49|8|non in sacrificiis tuis arguam te holocausta autem tua in conspectu meo sunt semper
PS|49|9|non accipiam de domo tua vitulos neque de gregibus tuis hircos
PS|49|10|quoniam meae sunt omnes ferae silvarum iumenta in montibus et boves
PS|49|11|cognovi omnia volatilia caeli et pulchritudo agri mecum est
PS|49|12|si esuriero non dicam tibi meus est enim orbis terrae et plenitudo eius
PS|49|13|numquid manducabo carnes taurorum aut sanguinem hircorum potabo
PS|49|14|immola Deo sacrificium laudis et redde Altissimo vota tua
PS|49|15|et invoca me in die tribulationis et eruam te et honorificabis me diapsalma
PS|49|16|peccatori autem dixit Deus quare tu enarras iustitias meas et adsumis testamentum meum per os tuum
PS|49|17|tu vero odisti disciplinam et proiecisti sermones meos retrorsum
PS|49|18|si videbas furem currebas cum eo et cum adulteris portionem tuam ponebas
PS|49|19|os tuum abundavit malitia et lingua tua concinnabat dolos
PS|49|20|sedens adversus fratrem tuum loquebaris et adversus filium matris tuae ponebas scandalum
PS|49|21|haec fecisti et tacui existimasti inique quod ero tui similis arguam te et statuam contra faciem tuam
PS|49|22|intellegite nunc haec qui obliviscimini Deum nequando rapiat et non sit qui eripiat
PS|49|23|sacrificium laudis honorificabit me et illic iter quod ostendam illi salutare Dei
PS|50|1|in finem psalmus David
PS|50|2|cum venit ad eum Nathan propheta quando intravit ad Bethsabee
PS|50|3|miserere mei Deus secundum %magnam; misericordiam tuam %et; secundum multitudinem miserationum tuarum dele iniquitatem meam
PS|50|4|amplius lava me ab iniquitate mea et a peccato meo munda me
PS|50|5|quoniam iniquitatem meam ego cognosco et peccatum meum contra me est semper
PS|50|6|tibi soli peccavi et malum coram te feci ut iustificeris in sermonibus tuis et vincas cum iudicaris
PS|50|7|ecce enim in iniquitatibus conceptus sum et in peccatis concepit me mater mea
PS|50|8|ecce enim veritatem dilexisti incerta et occulta sapientiae tuae manifestasti mihi
PS|50|9|asparges me hysopo et mundabor lavabis me et super nivem dealbabor
PS|50|10|auditui meo dabis gaudium et laetitiam exultabunt ossa humiliata
PS|50|11|averte faciem tuam a peccatis meis et omnes iniquitates meas dele
PS|50|12|cor mundum crea in me Deus et spiritum rectum innova in visceribus meis
PS|50|13|ne proicias me a facie tua et spiritum sanctum tuum ne auferas a me
PS|50|14|redde mihi laetitiam salutaris tui et spiritu principali confirma me
PS|50|15|docebo iniquos vias tuas et impii ad te convertentur
PS|50|16|libera me de sanguinibus Deus Deus salutis meae exultabit lingua mea iustitiam tuam
PS|50|17|Domine labia mea aperies et os meum adnuntiabit laudem tuam
PS|50|18|quoniam si voluisses sacrificium dedissem utique holocaustis non delectaberis
PS|50|19|sacrificium Deo spiritus contribulatus cor contritum et humiliatum Deus non spernet
PS|50|20|benigne fac Domine in bona voluntate tua Sion et aedificentur muri Hierusalem
PS|50|21|tunc acceptabis sacrificium iustitiae oblationes et holocausta tunc inponent super altare tuum vitulos
PS|51|1|in finem intellectus David
PS|51|2|cum venit Doec Idumeus et adnuntiavit Saul et dixit venit David in domo Achimelech
PS|51|3|quid gloriatur in malitia qui potens est iniquitate
PS|51|4|tota die iniustitiam cogitavit lingua tua sicut novacula acuta fecisti dolum
PS|51|5|dilexisti malitiam super benignitatem iniquitatem magis quam loqui aequitatem diapsalma
PS|51|6|dilexisti omnia verba praecipitationis linguam dolosam
PS|51|7|propterea Deus destruet te in finem evellet te et emigrabit te de tabernaculo et radicem tuam de terra viventium diapsalma
PS|51|8|videbunt iusti et timebunt et super eum ridebunt et dicent
PS|51|9|ecce homo qui non posuit Deum adiutorem suum sed speravit in multitudine divitiarum suarum et praevaluit in vanitate sua
PS|51|10|ego autem sicut oliva fructifera in domo Dei speravi in misericordia Dei in aeternum et in saeculum saeculi
PS|51|11|confitebor tibi in saeculum quia fecisti et expectabo nomen tuum quoniam bonum in conspectu sanctorum tuorum
PS|52|1|in finem pro Melech intellegentiae David dixit insipiens in corde suo non est Deus
PS|52|2|corrupti sunt et abominabiles facti sunt in iniquitatibus non est qui faciat bonum
PS|52|3|Deus de caelo prospexit in filios hominum ut videat si est intellegens %aut; requirens Deum
PS|52|4|omnes declinaverunt simul inutiles facti sunt non est qui faciat bonum non est usque ad unum
PS|52|5|nonne scient %omnes; qui operantur iniquitatem qui devorant plebem meam ut cibum panis
PS|52|6|Deum non invocaverunt illic trepidabunt timore ubi non fuit timor quoniam Deus dissipavit ossa eorum qui hominibus placent confusi sunt quoniam Deus sprevit eos
PS|52|7|quis dabit ex Sion salutare Israhel dum convertit Deus captivitatem plebis suae exultabit Iacob et laetabitur Israhel
PS|53|1|in finem in carminibus intellectus David
PS|53|2|cum venissent Ziphei et dixissent ad Saul nonne David absconditus est apud nos
PS|53|3|Deus in nomine tuo salvum me fac et in virtute tua iudica me
PS|53|4|Deus exaudi orationem meam auribus percipe verba oris mei
PS|53|5|quoniam alieni insurrexerunt adversum me et fortes quaesierunt animam meam non proposuerunt Deum ante conspectum suum diapsalma
PS|53|6|ecce enim Deus adiuvat me Dominus susceptor animae meae
PS|53|7|avertet mala inimicis meis in veritate tua disperde illos
PS|53|8|voluntarie sacrificabo tibi confitebor nomini tuo Domine quoniam bonum
PS|53|9|quoniam ex omni tribulatione eripuisti me et super inimicos meos despexit oculus meus
PS|54|1|in finem in carminibus intellectus David
PS|54|2|exaudi Deus orationem meam et ne despexeris deprecationem meam
PS|54|3|intende mihi et exaudi me contristatus sum in exercitatione mea et conturbatus sum
PS|54|4|a voce inimici et a tribulatione peccatoris quoniam declinaverunt in me iniquitatem et in ira molesti erant mihi
PS|54|5|cor meum conturbatum est in me et formido mortis cecidit super me
PS|54|6|timor et tremor venit super me et contexit me tenebra
PS|54|7|et dixi quis dabit mihi pinnas sicut columbae et volabo et requiescam
PS|54|8|ecce elongavi fugiens et mansi in solitudine diapsalma
PS|54|9|expectabam eum qui salvum me fecit a pusillanimitate spiritus et a tempestate
PS|54|10|praecipita Domine divide linguas eorum quoniam vidi iniquitatem et contradictionem in civitate
PS|54|11|die et nocte circumdabit eam super muros eius et iniquitas et labor in medio eius
PS|54|12|et iniustitia et non defecit de plateis eius usura et dolus
PS|54|13|quoniam si inimicus maledixisset mihi sustinuissem utique et si is qui oderat me super me magna locutus fuisset abscondissem me forsitan ab eo
PS|54|14|tu vero homo unianimis dux meus et notus meus
PS|54|15|qui simul mecum dulces capiebas cibos in domo Dei ambulavimus cum consensu
PS|54|16|veniat mors super illos et descendant in infernum viventes quoniam nequitiae in habitaculis eorum in medio eorum
PS|54|17|ego %autem; ad Deum clamavi et Dominus salvabit me
PS|54|18|vespere et mane et meridie narrabo et adnuntiabo et exaudiet vocem meam
PS|54|19|redimet in pace animam meam ab his qui adpropinquant mihi quoniam inter multos erant mecum
PS|54|20|exaudiet Deus et humiliabit illos qui est ante saecula diapsalma non enim est illis commutatio et non timuerunt Deum
PS|54|21|extendit manum suam in retribuendo contaminaverunt testamentum eius
PS|54|22|divisi sunt ab ira vultus eius et adpropinquavit cor illius molliti sunt sermones eius super oleum et ipsi sunt iacula
PS|54|23|iacta super Dominum curam tuam et ipse te enutriet non dabit in aeternum fluctuationem iusto
PS|54|24|tu vero Deus deduces eos in puteum interitus viri sanguinum et doli non dimidiabunt dies suos ego autem sperabo in te Domine
PS|55|1|in finem pro populo qui a sanctis longe factus est David in tituli inscriptione cum tenuerunt eum Allophili in Geth
PS|55|2|miserere mei Deus quoniam conculcavit me homo tota die inpugnans tribulavit me
PS|55|3|conculcaverunt me inimici mei tota die quoniam multi bellantes adversum me
PS|55|4|ab altitudine diei timebo ego vero in te sperabo
PS|55|5|in Deo laudabo sermones meos in Deo speravi non timebo quid faciat mihi caro
PS|55|6|tota die verba mea execrabantur adversum me omnia consilia eorum in malum
PS|55|7|inhabitabunt et abscondent ipsi calcaneum meum observabunt sicut sustinuerunt animam meam
PS|55|8|pro nihilo salvos facies illos in ira populos confringes Deus
PS|55|9|vitam meam adnuntiavi tibi posuisti lacrimas meas in conspectu tuo sicut et in promissione tua
PS|55|10|tunc convertentur inimici mei retrorsum in quacumque die invocavero te ecce cognovi quoniam Deus meus es
PS|55|11|in Deo laudabo verbum in Domino laudabo sermonem in Deo speravi non timebo quid faciat mihi homo
PS|55|12|in me sunt Deus vota tua; % quae; reddam laudationes tibi
PS|55|13|quoniam eripuisti animam meam de morte et pedes meos de lapsu ut placeam coram Deo in lumine viventium
PS|56|1|in finem ne disperdas David in tituli inscriptione cum fugeret a facie Saul in spelunca
PS|56|2|miserere mei Deus miserere mei quoniam in te confidit anima mea et in umbra alarum tuarum sperabo donec transeat iniquitas
PS|56|3|clamabo ad Deum altissimum Deum qui benefecit mihi
PS|56|4|misit de caelo et liberavit me dedit in obprobrium conculcantes me diapsalma misit Deus misericordiam suam et veritatem suam
PS|56|5|et eripuit animam meam de medio catulorum leonum dormivi conturbatus filii hominum dentes eorum arma et sagittae et lingua eorum gladius acutus
PS|56|6|exaltare super caelos Deus et in omnem terram gloria tua
PS|56|7|laqueum paraverunt pedibus meis et incurvaverunt animam meam foderunt ante faciem meam foveam et inciderunt in eam diapsalma
PS|56|8|paratum cor meum Deus paratum cor meum cantabo et psalmum dicam
PS|56|9|exsurge gloria mea exsurge psalterium et cithara exsurgam diluculo
PS|56|10|confitebor tibi in populis Domine psalmum dicam tibi in gentibus
PS|56|11|quoniam magnificata est usque ad caelos misericordia tua et usque ad nubes veritas tua
PS|56|12|exaltare super caelos Deus et super omnem terram gloria tua
PS|57|1|in finem ne disperdas David in tituli inscriptione
PS|57|2|si vere utique iustitiam loquimini recta iudicate filii hominum
PS|57|3|etenim in corde iniquitates operamini in terra iniustitiam manus vestrae concinnant
PS|57|4|alienati sunt peccatores a vulva erraverunt ab utero locuti sunt falsa
PS|57|5|furor illis secundum similitudinem serpentis sicut aspidis surdae et obturantis aures suas
PS|57|6|quae non exaudiet vocem incantantium et venefici incantantis sapienter
PS|57|7|Deus conteret dentes eorum in ore ipsorum molas leonum confringet Dominus
PS|57|8|ad nihilum devenient tamquam aqua decurrens intendit arcum suum donec infirmentur
PS|57|9|sicut cera quae fluit auferentur supercecidit ignis et non viderunt solem
PS|57|10|priusquam intellegerent spinae vestrae ramnum sicut viventes sicut in ira absorbet vos
PS|57|11|laetabitur iustus cum viderit vindictam manus suas lavabit in sanguine peccatoris
PS|57|12|et dicet homo si utique est fructus iusto utique est Deus iudicans eos in terra
PS|58|1|in finem ne disperdas David in tituli inscriptione quando misit Saul et custodivit domum eius ut interficeret eum
PS|58|2|eripe me de inimicis meis Deus et ab insurgentibus in me libera me
PS|58|3|eripe me de operantibus iniquitatem et de viris sanguinum salva me
PS|58|4|quia ecce ceperunt animam meam inruerunt in me fortes
PS|58|5|neque iniquitas mea neque peccatum meum Domine sine iniquitate cucurri et direxi
PS|58|6|exsurge in occursum meum et vide et tu Domine Deus virtutum Deus Israhel intende ad visitandas omnes gentes non miserearis omnibus qui operantur iniquitatem diapsalma
PS|58|7|convertentur ad vesperam et famem patientur ut canes et circuibunt civitatem
PS|58|8|ecce loquentur in ore suo et gladius in labiis eorum quoniam quis audivit
PS|58|9|et tu Domine deridebis eos ad nihilum deduces omnes gentes
PS|58|10|fortitudinem meam ad te custodiam quia Deus susceptor meus
PS|58|11|Deus meus voluntas eius praeveniet me
PS|58|12|Deus ostendet mihi super inimicos meos ne occidas eos nequando obliviscantur populi mei disperge illos in virtute tua et depone eos protector meus Domine
PS|58|13|delictum oris eorum sermonem labiorum ipsorum et conprehendantur in superbia sua et de execratione et mendacio adnuntiabuntur
PS|58|14|in consummatione in ira consummationis et non erunt et scient quia Deus dominatur Iacob finium terrae diapsalma
PS|58|15|convertentur ad vesperam et famem patientur ut canes et circuibunt civitatem
PS|58|16|ipsi dispergentur ad manducandum si vero non fuerint saturati et murmurabunt
PS|58|17|ego autem cantabo fortitudinem tuam et exultabo mane misericordiam tuam quia factus es susceptor meus et refugium meum in die tribulationis meae
PS|58|18|adiutor meus tibi psallam quia Deus susceptor meus es Deus meus misericordia mea
PS|59|1|in finem his qui inmutabuntur in tituli inscriptione David in doctrina
PS|59|2|cum succendit Syriam Mesopotamiam et Syriam Soba et convertit Ioab et percussit vallem Salinarum duodecim milia
PS|59|3|Deus reppulisti nos et destruxisti nos iratus es et misertus es nobis
PS|59|4|commovisti terram et turbasti eam sana contritiones eius quia commota est
PS|59|5|ostendisti populo tuo dura potasti nos vino conpunctionis
PS|59|6|dedisti metuentibus te significationem ut fugiant a facie arcus diapsalma ut liberentur dilecti tui
PS|59|7|salvum fac dextera tua et exaudi me
PS|59|8|Deus locutus est in sancto suo laetabor et partibor Sicima et convallem tabernaculorum metibor
PS|59|9|meus est Galaad et meus %est; Manasses et Effraim fortitudo capitis mei Iuda rex meus
PS|59|10|Moab olla spei meae in Idumeam extendam calciamentum meum mihi alienigenae subditi sunt
PS|59|11|quis deducet me in civitatem munitam quis deducet me usque in Idumeam
PS|59|12|nonne tu Deus qui reppulisti nos et non egredieris Deus in virtutibus nostris
PS|59|13|da nobis auxilium de tribulatione et vana salus hominis
PS|59|14|in Deo faciemus virtutem et ipse ad nihilum deducet tribulantes nos
PS|60|1|in finem in hymnis David
PS|60|2|exaudi Deus deprecationem meam intende orationi meae
PS|60|3|a finibus terrae ad te clamavi dum anxiaretur cor meum in petra exaltasti me deduxisti me
PS|60|4|quia factus es spes mea turris fortitudinis a facie inimici
PS|60|5|inhabitabo in tabernaculo tuo in saecula protegar in velamento alarum tuarum diapsalma
PS|60|6|quoniam tu Deus meus exaudisti orationem meam dedisti hereditatem timentibus nomen tuum
PS|60|7|dies super dies regis adicies annos eius usque in diem generationis et generationis
PS|60|8|permanet in aeternum in conspectu Dei misericordiam et veritatem quis requiret eius
PS|60|9|sic psalmum dicam nomini tuo in saeculum saeculi ut reddam vota mea de die in diem
PS|61|1|in finem pro Idithun psalmus David
PS|61|2|nonne Deo subiecta erit anima mea ab ipso enim salutare meum
PS|61|3|nam et ipse Deus meus et salutaris meus susceptor meus non movebor amplius
PS|61|4|quousque inruitis in hominem interficitis universi vos tamquam parieti inclinato et maceriae depulsae
PS|61|5|verumtamen pretium meum cogitaverunt repellere cucurri in siti ore suo benedicebant et corde suo maledicebant diapsalma
PS|61|6|verumtamen Deo subiecta esto anima mea quoniam ab ipso patientia mea
PS|61|7|quia ipse Deus meus et salvator meus adiutor meus non emigrabo
PS|61|8|in Deo salutare meum et gloria mea Deus auxilii mei et spes mea in Deo est
PS|61|9|sperate in eo omnis congregatio populi effundite coram illo corda vestra Deus adiutor noster in aeternum
PS|61|10|verumtamen vani filii hominum mendaces filii hominum in stateris ut decipiant ipsi de vanitate in id ipsum
PS|61|11|nolite sperare in iniquitate et rapinas nolite concupiscere divitiae si affluant nolite cor adponere
PS|61|12|semel locutus est Deus duo haec audivi quia potestas Dei
PS|61|13|et tibi Domine misericordia quia tu reddes unicuique iuxta opera sua
PS|62|1|psalmus David cum esset in deserto Iudaeae
PS|62|2|Deus Deus meus ad te de luce vigilo sitivit in te anima mea quam multipliciter tibi caro mea
PS|62|3|in terra deserta et invia et inaquosa sic in sancto apparui tibi ut viderem virtutem tuam et gloriam tuam
PS|62|4|quoniam melior est misericordia tua super vitas labia mea laudabunt te
PS|62|5|sic benedicam te in vita mea in nomine tuo levabo manus meas
PS|62|6|sicut adipe et pinguidine repleatur anima mea et labia exultationis laudabit os meum
PS|62|7|si memor fui tui super stratum meum in matutinis meditabar in te
PS|62|8|quia fuisti adiutor meus et in velamento alarum tuarum exultabo
PS|62|9|adhesit anima mea post te me suscepit dextera tua
PS|62|10|ipsi vero in vanum quaesierunt animam meam introibunt in inferiora terrae
PS|62|11|tradentur in manus gladii partes vulpium erunt
PS|62|12|rex vero laetabitur in Deo laudabitur omnis qui iurat in eo quia obstructum est os loquentium iniqua
PS|63|1|in finem psalmus David
PS|63|2|exaudi Deus orationem meam cum deprecor a timore inimici eripe animam meam
PS|63|3|protexisti me a conventu malignantium a multitudine operantium iniquitatem
PS|63|4|quia exacuerunt ut gladium linguas suas intenderunt arcum rem amaram
PS|63|5|ut sagittent in occultis inmaculatum
PS|63|6|subito sagittabunt eum et non timebunt firmaverunt sibi sermonem nequam narraverunt ut absconderent laqueos dixerunt quis videbit eos
PS|63|7|scrutati sunt iniquitates defecerunt scrutantes scrutinio accedet homo et cor altum
PS|63|8|et exaltabitur Deus sagittae parvulorum factae sunt plagae eorum
PS|63|9|et infirmatae sunt contra eos linguae eorum conturbati sunt omnes qui videbant eos
PS|63|10|et timuit omnis homo et adnuntiaverunt opera Dei et facta eius intellexerunt
PS|63|11|laetabitur iustus in Domino et sperabit in eo et laudabuntur omnes recti corde
PS|64|1|in finem psalmus David canticum; Hieremiae et Aggei de verbo peregrinationis quando incipiebant proficisci
PS|64|2|te decet hymnus Deus in Sion et tibi reddetur votum in Hierusalem
PS|64|3|exaudi orationem ad te omnis caro veniet
PS|64|4|verba iniquorum praevaluerunt super nos et impietatibus nostris tu propitiaberis
PS|64|5|beatus quem elegisti et adsumpsisti inhabitabit in atriis tuis replebimur in bonis domus tuae sanctum est templum tuum
PS|64|6|mirabile in aequitate exaudi nos Deus salutaris noster spes omnium finium terrae et in mari longe
PS|64|7|praeparans montes in virtute tua accinctus potentia
PS|64|8|qui conturbas profundum maris sonum fluctuum eius turbabuntur gentes
PS|64|9|et timebunt qui inhabitant terminos a signis tuis exitus matutini et vespere delectabis
PS|64|10|visitasti terram et inebriasti eam multiplicasti locupletare eam flumen Dei repletum est aquis parasti cibum illorum quoniam ita est praeparatio eius
PS|64|11|rivos eius inebria multiplica genimina eius in stillicidiis eius laetabitur germinans
PS|64|12|benedices coronae anni benignitatis tuae et campi tui replebuntur ubertate
PS|64|13|pinguescent speciosa deserti et exultatione colles accingentur
PS|64|14|induti sunt arietes ovium et valles abundabunt frumento clamabunt etenim hymnum dicent
PS|65|1|in finem canticum psalmi resurrectionis iubilate Deo omnis terra
PS|65|2|psalmum dicite nomini eius date gloriam laudi eius
PS|65|3|dicite Deo quam terribilia sunt opera tua Domine in multitudine virtutis tuae mentientur tibi inimici tui
PS|65|4|omnis terra adorent te et psallant tibi psalmum dicant nomini tuo diapsalma
PS|65|5|venite et videte opera Dei terribilis in consiliis super filios hominum
PS|65|6|qui convertit mare in aridam in flumine pertransibunt pede ibi laetabimur in ipso
PS|65|7|qui dominatur in virtute sua in aeternum oculi eius super gentes respiciunt qui exasperant non exaltentur in semet ipsis diapsalma
PS|65|8|benedicite gentes Deum nostrum et auditam facite vocem laudis eius
PS|65|9|qui posuit animam meam ad vitam et non dedit in commotionem pedes meos
PS|65|10|quoniam probasti nos Deus igne nos examinasti sicut examinatur argentum
PS|65|11|induxisti nos in laqueum posuisti tribulationes in dorso nostro
PS|65|12|inposuisti homines super capita nostra transivimus per ignem et aquam et eduxisti nos in refrigerium
PS|65|13|introibo in domum tuam in holocaustis reddam tibi vota mea
PS|65|14|quae distinxerunt labia mea et locutum est os meum in tribulatione mea
PS|65|15|holocausta medullata offeram tibi cum incensu arietum offeram tibi boves cum hircis diapsalma
PS|65|16|venite audite et narrabo omnes qui timetis Deum quanta fecit animae meae
PS|65|17|ad ipsum ore meo clamavi et exaltavi sub lingua mea
PS|65|18|iniquitatem si aspexi in corde meo non exaudiat Dominus
PS|65|19|propterea exaudivit Deus adtendit voci deprecationis meae
PS|65|20|benedictus Deus qui non amovit orationem meam et misericordiam suam a me
PS|66|1|in finem in hymnis psalmus cantici
PS|66|2|Deus misereatur nostri et benedicat nobis inluminet vultum suum super nos et misereatur nostri diapsalma
PS|66|3|ut cognoscamus in terra viam tuam in omnibus gentibus salutare tuum
PS|66|4|confiteantur tibi populi Deus confiteantur tibi populi omnes
PS|66|5|laetentur et exultent gentes quoniam iudicas populos in aequitate et gentes in terra diriges diapsalma
PS|66|6|confiteantur tibi populi Deus confiteantur tibi populi omnes
PS|66|7|terra dedit fructum suum benedicat nos Deus Deus noster
PS|66|8|benedicat nos Deus et metuant eum omnes fines terrae
PS|67|1|in finem David psalmus cantici
PS|67|2|exsurgat Deus et dissipentur inimici eius et fugiant qui oderunt eum a facie eius
PS|67|3|sicut deficit fumus deficiant sicut fluit cera a facie ignis sic pereant peccatores a facie Dei
PS|67|4|et iusti epulentur exultent in conspectu Dei delectentur in laetitia
PS|67|5|cantate Deo psalmum dicite nomini eius iter facite ei qui ascendit super occasum Dominus nomen illi et exultate in conspectu eius turbabuntur a facie eius
PS|67|6|patris orfanorum et iudicis viduarum Deus in loco sancto suo
PS|67|7|Deus inhabitare facit unius moris in domo qui educit vinctos in fortitudine similiter eos qui exasperant qui habitant in sepulchris
PS|67|8|Deus cum egredereris in conspectu populi tui cum pertransieris in deserto diapsalma
PS|67|9|terra mota est etenim caeli distillaverunt a facie Dei Sinai a facie Dei Israhel
PS|67|10|pluviam voluntariam segregabis Deus hereditati tuae et infirmata est tu vero perfecisti eam
PS|67|11|animalia tua habitant in ea parasti in dulcedine tua pauperi Deus
PS|67|12|Dominus dabit verbum evangelizantibus virtute multa
PS|67|13|rex virtutum dilecti dilecti; et speciei domus dividere spolia
PS|67|14|si dormiatis inter medios cleros pinnae columbae deargentatae et posteriora dorsi eius in pallore auri
PS|67|15|dum discernit Caelestis reges super eam nive dealbabuntur in Selmon
PS|67|16|mons Dei mons pinguis mons coagulatus mons pinguis
PS|67|17|ut quid suspicamini montes coagulatos mons in quo beneplacitum est Deo habitare in eo etenim Dominus habitabit in finem
PS|67|18|currus Dei decem milibus multiplex milia laetantium Dominus in eis in Sina in sancto
PS|67|19|ascendisti in altum cepisti captivitatem accepisti dona in hominibus etenim non credentes inhabitare Dominum Deus
PS|67|20|benedictus Dominus die cotidie prosperum iter faciet nobis Deus salutarium nostrorum diapsalma
PS|67|21|Deus noster Deus salvos faciendi et Domini Domini exitus mortis
PS|67|22|verumtamen Deus confringet capita inimicorum suorum verticem capilli perambulantium in delictis suis
PS|67|23|dixit Dominus ex Basan convertam convertam in profundis maris
PS|67|24|ut intinguatur pes tuus in sanguine lingua canum tuorum ex inimicis ab ipso
PS|67|25|viderunt ingressus tui Deus ingressus Dei mei regis mei qui est in sancto
PS|67|26|praevenerunt principes coniuncti psallentibus in medio iuvencularum tympanistriarum
PS|67|27|in ecclesiis benedicite Deum Dominum de fontibus Israhel
PS|67|28|ibi Beniamin adulescentulus in mentis excessu principes Iuda duces eorum principes Zabulon principes Nepthali
PS|67|29|manda Deus virtutem tuam confirma Deus hoc quod operatus es nobis
PS|67|30|a templo tuo in Hierusalem tibi adferent reges munera
PS|67|31|increpa feras harundinis congregatio taurorum in vaccis populorum ut excludant eos qui probati sunt argento dissipa gentes quae bella volunt
PS|67|32|venient legati ex Aegypto Aethiopia praeveniet manus eius Deo
PS|67|33|regna terrae cantate Deo psallite Domino diapsalma %psallite Deo;
PS|67|34|qui ascendit super caelum caeli ad orientem ecce dabit voci suae vocem virtutis
PS|67|35|date gloriam Deo super Israhel magnificentia eius et virtus eius in nubibus
PS|67|36|mirabilis Deus in sanctis suis Deus Israhel ipse dabit virtutem et fortitudinem plebi suae benedictus Deus
PS|68|1|in finem pro his qui commutabuntur David
PS|68|2|salvum me fac Deus quoniam intraverunt aquae usque ad animam meam
PS|68|3|infixus sum in limum profundi et non est substantia veni in altitudines maris et tempestas demersit me
PS|68|4|laboravi clamans raucae factae sunt fauces meae defecerunt oculi mei dum spero in Deum meum
PS|68|5|multiplicati sunt super capillos capitis mei qui oderunt me gratis confortati sunt qui persecuti sunt me inimici mei iniuste quae non rapui tunc exsolvebam
PS|68|6|Deus tu scis insipientiam meam et delicta mea a te non sunt abscondita
PS|68|7|non erubescant in me qui expectant te Domine Domine virtutum non confundantur super me qui quaerunt te Deus Israhel
PS|68|8|quoniam propter te sustinui obprobrium operuit confusio faciem meam
PS|68|9|extraneus factus sum fratribus meis et peregrinus filiis matris meae
PS|68|10|quoniam zelus domus tuae comedit me et obprobria exprobrantium tibi ceciderunt super me
PS|68|11|et operui in ieiunio animam meam et factum est in obprobrium mihi
PS|68|12|et posui vestimentum meum cilicium et factus sum illis in parabolam
PS|68|13|adversum me exercebantur qui sedebant in porta et in me psallebant qui bibebant vinum
PS|68|14|ego vero orationem meam ad te Domine tempus beneplaciti Deus in multitudine misericordiae tuae exaudi me in veritate salutis tuae
PS|68|15|eripe me de luto ut non infigar liberer ab his qui oderunt me et de profundis aquarum
PS|68|16|non me demergat tempestas aquae neque absorbeat me profundum neque urgeat super me puteus os suum
PS|68|17|exaudi me Domine quoniam benigna est misericordia tua secundum multitudinem miserationum tuarum respice me
PS|68|18|et ne avertas faciem tuam a puero tuo quoniam tribulor velociter exaudi me
PS|68|19|intende animae meae et libera eam propter inimicos meos eripe me
PS|68|20|tu scis inproperium meum et confusionem et reverentiam meam
PS|68|21|in conspectu tuo sunt omnes qui tribulant me inproperium expectavit cor meum et miseriam et sustinui qui simul contristaretur et non fuit et qui consolaretur et non inveni
PS|68|22|et dederunt in escam meam fel et in siti mea potaverunt me aceto
PS|68|23|fiat mensa eorum coram ipsis in laqueum et in retributiones et in scandalum
PS|68|24|obscurentur oculi eorum ne videant et dorsum eorum semper incurva
PS|68|25|effunde super eos iram tuam et furor irae tuae conprehendat eos
PS|68|26|fiat habitatio eorum deserta et in tabernaculis eorum non sit qui inhabitet
PS|68|27|quoniam quem tu percussisti persecuti sunt et super dolorem vulnerum meorum addiderunt
PS|68|28|adpone iniquitatem super iniquitatem eorum et non intrent in iustitia tua
PS|68|29|deleantur de libro viventium et cum iustis non scribantur
PS|68|30|ego sum pauper et dolens salus tua Deus suscepit me
PS|68|31|laudabo nomen Dei cum cantico magnificabo eum in laude
PS|68|32|et placebit Deo super vitulum novellum cornua producentem et ungulas
PS|68|33|videant pauperes et laetentur quaerite Deum et vivet anima vestra
PS|68|34|quoniam exaudivit pauperes Dominus et vinctos suos non despexit
PS|68|35|laudent illum caeli et terra mare et omnia reptilia in eis
PS|68|36|quoniam Deus salvam faciet Sion et aedificabuntur civitates Iudaeae et inhabitabunt ibi et hereditate adquirent eam
PS|68|37|et semen servorum eius possidebunt eam et qui diligunt nomen eius habitabunt in ea
PS|69|1|in finem David in rememoratione eo quod salvum me fecit Dominus
PS|69|2|Deus in adiutorium meum intende Domine ad adiuvandum me festina;
PS|69|3|confundantur et revereantur qui quaerunt animam meam
PS|69|4|avertantur retrorsum et erubescant qui volunt mihi mala avertantur statim erubescentes qui dicunt %mihi; euge euge
PS|69|5|exultent et laetentur in te omnes qui quaerunt te et dicant semper magnificetur Deus qui diligunt salutare tuum
PS|69|6|ego vero egenus et pauper Deus adiuva me adiutor meus et liberator meus es tu Domine ne moreris
PS|69|7|
PS|69|8|
PS|69|9|
PS|70|1|David psalmus filiorum Ionadab et priorum captivorum in te Domine speravi non confundar in aeternum
PS|70|2|in iustitia tua libera me et eripe me inclina ad me aurem tuam et salva me
PS|70|3|esto mihi in Deum protectorem et in locum munitum ut salvum me facias quoniam firmamentum meum et refugium meum es tu
PS|70|4|Deus meus eripe me de manu peccatoris de manu contra legem agentis et iniqui
PS|70|5|quoniam tu es patientia mea Domine Domine spes mea a iuventute mea
PS|70|6|in te confirmatus sum ex utero de ventre matris meae tu es protector meus in te cantatio mea semper
PS|70|7|tamquam prodigium factus sum multis et tu adiutor fortis
PS|70|8|repleatur os meum laude ut cantem gloriam tuam tota die magnitudinem tuam
PS|70|9|non proicias me in tempore senectutis cum deficiet virtus mea ne derelinquas me
PS|70|10|quia dixerunt inimici mei mihi et qui custodiebant animam meam consilium fecerunt in unum
PS|70|11|dicentes Deus dereliquit eum persequimini et conprehendite eum quia non est qui eripiat
PS|70|12|Deus ne elongeris a me Deus meus in adiutorium meum respice
PS|70|13|confundantur et deficiant detrahentes animae meae operiantur confusione et pudore qui quaerunt mala mihi
PS|70|14|ego autem semper sperabo et adiciam super omnem laudem tuam
PS|70|15|os meum adnuntiabit iustitiam tuam tota die salutem tuam quoniam non cognovi litteraturam
PS|70|16|introibo in potentiam Domini Domine memorabor iustitiae tuae solius
PS|70|17|Deus docuisti me ex iuventute mea et usque nunc pronuntiabo mirabilia tua
PS|70|18|et usque in senectam et senium Deus ne derelinquas me donec adnuntiem brachium tuum generationi omni quae ventura est potentiam tuam
PS|70|19|et iustitiam tuam Deus usque in altissima quae fecisti magnalia Deus quis similis tibi
PS|70|20|quantas ostendisti mihi tribulationes multas et malas et conversus vivificasti me et de abyssis terrae iterum reduxisti me
PS|70|21|multiplicasti magnificentiam tuam et conversus consolatus es me
PS|70|22|nam et ego confitebor tibi in vasis psalmi veritatem tuam Deus psallam tibi in cithara Sanctus Israhel
PS|70|23|exultabunt labia mea cum cantavero tibi et anima mea quam redemisti
PS|70|24|sed et lingua mea tota die meditabitur iustitiam tuam cum confusi et reveriti fuerint qui quaerunt mala mihi
PS|71|1|in Salomonem
PS|71|2|Deus iudicium tuum regi da et iustitiam tuam filio regis iudicare populum tuum in iustitia et pauperes tuos in iudicio
PS|71|3|suscipiant montes pacem populo et colles iustitiam
PS|71|4|iudicabit pauperes populi et salvos faciet filios pauperum et humiliabit calumniatorem
PS|71|5|et permanebit cum sole et ante lunam generationes generationum
PS|71|6|descendet sicut pluvia in vellus et sicut stillicidia stillantia super terram
PS|71|7|orietur in diebus eius iustitia et abundantia pacis donec auferatur luna
PS|71|8|et dominabitur a mari usque ad mare et a flumine usque ad terminos orbis terrarum
PS|71|9|coram illo procident Aethiopes et inimici eius terram lingent
PS|71|10|reges Tharsis et insulae munera offerent reges Arabum et Saba dona adducent
PS|71|11|et adorabunt eum omnes reges omnes gentes servient ei
PS|71|12|quia liberavit pauperem a potente et pauperem cui non erat adiutor
PS|71|13|parcet pauperi et inopi et animas pauperum salvas faciet
PS|71|14|ex usuris et iniquitate redimet animas eorum et honorabile nomen eorum coram illo
PS|71|15|et vivet et dabitur ei de auro Arabiae et orabunt de ipso semper tota die benedicent ei
PS|71|16|erit firmamentum in terra in summis montium superextolletur super Libanum fructus eius et florebunt de civitate sicut faenum terrae
PS|71|17|sit nomen eius benedictum in saecula ante solem permanet nomen eius et benedicentur in ipso omnes tribus terrae omnes gentes beatificabunt eum
PS|71|18|benedictus Dominus Deus Deus Israhel qui facit mirabilia solus
PS|71|19|et benedictum nomen maiestatis eius in aeternum et replebitur maiestate eius omnis terra fiat fiat
PS|71|20|defecerunt laudes David filii Iesse
PS|72|1|psalmus Asaph quam bonus Israhel Deus his qui recto sunt corde
PS|72|2|mei autem paene moti sunt pedes paene effusi sunt gressus mei
PS|72|3|quia zelavi super iniquis pacem peccatorum videns
PS|72|4|quia non est respectus morti eorum et firmamentum in plaga eorum
PS|72|5|in labore hominum non sunt et cum hominibus non flagellabuntur
PS|72|6|ideo tenuit eos superbia operti sunt iniquitate et impietate sua
PS|72|7|prodiet quasi ex adipe iniquitas eorum transierunt in affectum cordis
PS|72|8|cogitaverunt et locuti sunt in nequitia iniquitatem in excelso locuti sunt
PS|72|9|posuerunt in caelum os suum et lingua eorum transivit in terra
PS|72|10|ideo convertetur populus meus hic et dies pleni invenientur in eis
PS|72|11|et dixerunt quomodo scit Deus et si est scientia in Excelso
PS|72|12|ecce ipsi peccatores et abundantes in saeculo obtinuerunt divitias
PS|72|13|%et dixi; ergo sine causa iustificavi cor meum et lavi inter innocentes manus meas
PS|72|14|et fui flagellatus tota die et castigatio mea in matutino
PS|72|15|si dicebam narrabo sic ecce nationem filiorum tuorum reprobavi
PS|72|16|et existimabam cognoscere hoc labor est ante me
PS|72|17|donec intrem in sanctuarium Dei intellegam in novissimis eorum
PS|72|18|verumtamen propter dolos posuisti eis deiecisti eos dum adlevarentur
PS|72|19|quomodo facti sunt in desolationem subito defecerunt perierunt propter iniquitatem suam
PS|72|20|velut somnium surgentium Domine in civitate tua imaginem ipsorum ad nihilum rediges
PS|72|21|quia inflammatum est cor meum et renes mei commutati sunt
PS|72|22|et ego ad nihilum redactus sum et nescivi
PS|72|23|ut iumentum factus sum apud te et ego semper tecum
PS|72|24|tenuisti manum dexteram meam et in voluntate tua deduxisti me et cum gloria suscepisti me
PS|72|25|quid enim mihi est in caelo et a te quid volui super terram
PS|72|26|defecit caro mea et cor meum Deus cordis mei et pars mea Deus in aeternum
PS|72|27|quia ecce qui elongant se a te peribunt perdidisti omnem qui fornicatur abs te
PS|72|28|mihi autem adherere Deo bonum est ponere in Domino Deo spem meam ut adnuntiem omnes praedicationes tuas % in portis filiae Sion;
PS|73|1|intellectus Asaph ut quid Deus reppulisti in finem iratus est furor tuus super oves pascuae tuae
PS|73|2|memor esto congregationis tuae quam possedisti ab initio redemisti virgam hereditatis tuae mons Sion in quo habitasti in eo
PS|73|3|leva manus tuas in superbias eorum in finem quanta malignatus est inimicus in sancto
PS|73|4|et gloriati sunt qui oderunt te in medio sollemnitatis tuae posuerunt signa sua signa
PS|73|5|et non cognoverunt sicut in exitu super summum quasi in silva lignorum securibus
PS|73|6|exciderunt ianuas eius in id ipsum in securi et ascia deiecerunt %eam;
PS|73|7|incenderunt igni sanctuarium tuum in terra polluerunt tabernaculum nominis tui
PS|73|8|dixerunt in corde suo cognatio eorum simul quiescere faciamus omnes dies festos Dei a terra
PS|73|9|signa nostra non vidimus iam non est propheta et nos non cognoscet amplius
PS|73|10|usquequo Deus inproperabit inimicus inritat adversarius nomen tuum in finem
PS|73|11|ut quid avertis manum tuam et dexteram tuam de medio sinu tuo in finem
PS|73|12|Deus autem rex noster ante saeculum operatus est salutes in medio terrae
PS|73|13|tu confirmasti in virtute tua mare contribulasti capita draconum in aquis
PS|73|14|tu confregisti capita draconis dedisti eum escam populis Aethiopum
PS|73|15|tu disrupisti fontem et torrentes tu siccasti fluvios Aetham;
PS|73|16|tuus est dies et tua est nox tu fabricatus es auroram et solem
PS|73|17|tu fecisti omnes terminos terrae aestatem et ver tu plasmasti ea
PS|73|18|memor esto huius inimicus inproperavit Dominum et populus insipiens incitavit nomen tuum
PS|73|19|ne tradas bestiis animam confitentem tibi animas pauperum tuorum ne obliviscaris in finem
PS|73|20|respice in testamentum tuum quia repleti sunt qui obscurati sunt terrae domibus iniquitatum
PS|73|21|ne avertatur humilis factus confusus pauper et inops laudabunt nomen tuum
PS|73|22|exsurge Deus iudica causam tuam memor esto inproperiorum tuorum eorum qui ab insipiente sunt tota die
PS|73|23|ne obliviscaris voces inimicorum tuorum superbia eorum qui te oderunt ascendit semper
PS|74|1|in finem ne corrumpas psalmus Asaph cantici
PS|74|2|confitebimur tibi Deus confitebimur et invocabimus nomen tuum narrabimus mirabilia tua
PS|74|3|cum accepero tempus ego iustitias iudicabo
PS|74|4|liquefacta est terra et omnes qui habitant in ea ego confirmavi columnas eius diapsalma
PS|74|5|dixi iniquis nolite inique facere et delinquentibus nolite exaltare cornu
PS|74|6|nolite extollere in altum cornu vestrum nolite loqui adversus Deum iniquitatem
PS|74|7|quia neque ab oriente neque ab occidente neque a desertis montibus
PS|74|8|quoniam Deus iudex est hunc humiliat et hunc exaltat
PS|74|9|quia calix in manu Domini vini meri plenus mixto et inclinavit ex hoc in hoc verum fex eius non est exinanita bibent omnes peccatores terrae
PS|74|10|ego autem adnuntiabo in saeculum cantabo Deo Iacob
PS|74|11|et omnia cornua peccatorum confringam et exaltabuntur cornua iusti
PS|75|1|in finem in laudibus psalmus Asaph canticum ad Assyrium
PS|75|2|notus in Iudaea Deus in Israhel magnum nomen eius
PS|75|3|et factus est in pace locus eius et habitatio eius in Sion
PS|75|4|ibi confregit potentias arcuum scutum et gladium et bellum diapsalma
PS|75|5|inluminas tu mirabiliter de montibus aeternis
PS|75|6|turbati sunt omnes insipientes corde dormierunt somnum suum et nihil invenerunt omnes viri divitiarum manibus suis
PS|75|7|ab increpatione tua Deus Iacob dormitaverunt qui ascenderunt equos
PS|75|8|tu terribilis es et quis resistet tibi ex tunc ira tua
PS|75|9|de caelo auditum fecisti iudicium terra timuit et quievit
PS|75|10|cum exsurgeret in iudicium Deus ut salvos faceret omnes mansuetos terrae diapsalma
PS|75|11|quoniam cogitatio hominis confitebitur tibi et reliquiae cogitationis diem festum agent tibi
PS|75|12|vovete et reddite Domino Deo vestro omnes qui in circuitu eius adferent munera terribili
PS|75|13|et ei qui aufert spiritus principum terribili apud reges terrae
PS|76|1|in finem pro Idithun psalmus Asaph
PS|76|2|voce mea ad Dominum clamavi voce mea ad Deum et intendit me
PS|76|3|in die tribulationis meae Deum exquisivi manibus meis nocte contra eum et non sum deceptus rennuit consolari anima mea
PS|76|4|memor fui Dei et delectatus sum exercitatus sum et defecit spiritus meus diapsalma
PS|76|5|anticipaverunt vigilias oculi mei turbatus sum et non sum locutus
PS|76|6|cogitavi dies antiquos et annos aeternos in mente habui
PS|76|7|et meditatus sum nocte cum corde meo exercitabar et scobebam spiritum meum
PS|76|8|numquid in aeternum proiciet Deus et non adponet ut conplacitior sit adhuc
PS|76|9|aut in finem misericordiam suam abscidet a generatione in generationem
PS|76|10|aut obliviscetur misereri Deus aut continebit in ira sua misericordias suas diapsalma
PS|76|11|et dixi nunc coepi haec mutatio dexterae Excelsi
PS|76|12|memor fui operum Domini quia memor ero ab initio mirabilium tuorum
PS|76|13|et meditabor in omnibus operibus tuis et in adinventionibus tuis exercebor
PS|76|14|Deus in sancto via tua quis deus magnus sicut Deus noster
PS|76|15|tu es Deus qui facis mirabilia notam fecisti in populis virtutem tuam
PS|76|16|redemisti in brachio tuo populum tuum filios Iacob et Ioseph diapsalma
PS|76|17|viderunt te aquae Deus viderunt te aquae et timuerunt et turbatae sunt abyssi
PS|76|18|multitudo sonitus aquarum vocem dederunt nubes etenim sagittae tuae transeunt
PS|76|19|vox tonitrui tui in rota inluxerunt coruscationes tuae orbi terrae commota est et contremuit terra
PS|76|20|in mari via tua et semitae tuae in aquis multis et vestigia tua non cognoscentur
PS|76|21|deduxisti sicut oves populum tuum in manu Mosi et Aaron
PS|77|1|intellectus Asaph adtendite populus meus legem meam inclinate aurem vestram in verba oris mei
PS|77|2|aperiam in parabola os meum eloquar propositiones ab initio
PS|77|3|quanta audivimus et cognovimus ea et patres nostri narraverunt nobis
PS|77|4|non sunt occultata a filiis eorum in generationem alteram narrantes laudes Domini et virtutes eius et mirabilia eius quae fecit
PS|77|5|et suscitavit testimonium in Iacob et legem posuit in Israhel quanta mandavit patribus nostris nota facere ea filiis suis
PS|77|6|ut cognoscat generatio altera filii qui nascentur et exsurgent et narrabunt filiis suis
PS|77|7|ut ponant in Deo spem suam et non obliviscantur opera Dei et mandata eius exquirant
PS|77|8|ne fiant sicut patres eorum generatio prava et exasperans generatio quae non direxit cor suum et non est creditus cum Deo spiritus eius
PS|77|9|filii Effrem intendentes et mittentes arcus conversi sunt in die belli
PS|77|10|non custodierunt testamentum Dei et in lege eius noluerunt ambulare
PS|77|11|et obliti sunt benefactorum eius et mirabilium eius quae ostendit eis
PS|77|12|coram patribus eorum quae fecit mirabilia in terra Aegypti in campo Taneos
PS|77|13|interrupit mare et perduxit eos statuit aquas quasi utrem
PS|77|14|et deduxit eos in nube diei et tota nocte in inluminatione ignis
PS|77|15|interrupit petram in heremo et adaquavit eos velut in abysso multa
PS|77|16|et eduxit aquam de petra et deduxit tamquam flumina aquas
PS|77|17|et adposuerunt adhuc peccare ei in ira excitaverunt Excelsum in inaquoso
PS|77|18|et temptaverunt Deum in cordibus suis ut peterent escas animabus suis
PS|77|19|et male locuti sunt de Deo dixerunt numquid poterit Deus parare mensam in deserto
PS|77|20|quoniam percussit petram et fluxerunt aquae et torrentes inundaverunt numquid et panem potest dare aut parare mensam populo suo
PS|77|21|ideo audivit Dominus et distulit et ignis accensus est in Iacob et ira ascendit in Israhel
PS|77|22|quia non crediderunt in Deo nec speraverunt in salutare eius
PS|77|23|et mandavit nubibus desuper et ianuas caeli aperuit
PS|77|24|et pluit illis manna ad manducandum et panem caeli dedit eis
PS|77|25|panem angelorum manducavit homo cibaria misit eis in abundantiam
PS|77|26|transtulit austrum de caelo et induxit in virtute sua africum
PS|77|27|et pluit super eos sicut pulverem carnes et sicut harenam maris volatilia pinnata
PS|77|28|et ceciderunt in medio castrorum eorum circa tabernacula eorum
PS|77|29|et manducaverunt et saturati sunt nimis et desiderium eorum adtulit eis
PS|77|30|non sunt fraudati a desiderio suo adhuc escae eorum erant in ore ipsorum
PS|77|31|et ira Dei ascendit in eos et occidit pingues eorum et electos Israhel inpedivit
PS|77|32|in omnibus his peccaverunt adhuc et non crediderunt mirabilibus eius
PS|77|33|et defecerunt in vanitate dies eorum et anni eorum cum festinatione
PS|77|34|cum occideret eos quaerebant eum et revertebantur et diluculo veniebant ad Deum
PS|77|35|et rememorati sunt quia Deus adiutor est eorum et Deus excelsus redemptor eorum est
PS|77|36|et dilexerunt eum in ore suo et lingua sua mentiti sunt ei
PS|77|37|cor autem ipsorum non erat rectum cum eo nec fideles habiti sunt in testamento eius
PS|77|38|ipse autem est misericors et propitius fiet peccatis eorum et non perdet eos et abundabit ut avertat iram suam et non accendet omnem iram suam
PS|77|39|et recordatus est quia caro sunt spiritus vadens et non rediens
PS|77|40|quotiens exacerbaverunt eum in deserto in ira concitaverunt eum in inaquoso
PS|77|41|et conversi sunt et temptaverunt Deum et Sanctum Israhel exacerbaverunt
PS|77|42|non sunt recordati manus eius die qua redemit eos de manu tribulantis
PS|77|43|sicut posuit in Aegypto signa sua et prodigia sua in campo Taneos
PS|77|44|et convertit in sanguine flumina eorum et imbres eorum ne biberent
PS|77|45|misit in eos cynomiam et comedit eos et ranam et disperdit eos
PS|77|46|et dedit erugini fructus eorum et labores eorum lucustae
PS|77|47|et occidit in grandine vineam eorum et moros eorum in pruina
PS|77|48|et tradidit grandini iumenta eorum et possessionem eorum igni
PS|77|49|misit in eos iram indignationis suae indignationem et iram et tribulationem inmissionem per angelos malos
PS|77|50|viam fecit semitae irae suae non pepercit a morte animarum eorum et iumenta eorum in morte conclusit
PS|77|51|et percussit omne primitivum in terra Aegypti primitias laborum eorum in tabernaculis Cham
PS|77|52|et abstulit sicut oves populum suum et perduxit eos tamquam gregem in deserto
PS|77|53|et deduxit eos in spe et non timuerunt et inimicos eorum operuit mare
PS|77|54|et induxit eos in montem sanctificationis suae montem quem adquisivit dextera eius et eiecit a facie eorum gentes et sorte divisit eis terram in funiculo distributionis
PS|77|55|et habitare fecit in tabernaculis eorum tribus Israhel
PS|77|56|et temptaverunt et exacerbaverunt Deum excelsum et testimonia eius non custodierunt
PS|77|57|et averterunt se et non servaverunt pactum quemadmodum patres eorum conversi sunt in arcum pravum
PS|77|58|et in ira concitaverunt eum in collibus suis et in sculptilibus suis ad aemulationem eum provocaverunt
PS|77|59|audivit Deus et sprevit et ad nihilum redegit valde Israhel
PS|77|60|et reppulit tabernaculum Selo tabernaculum suum ubi habitavit in hominibus
PS|77|61|et tradidit in captivitatem virtutem eorum et pulchritudinem eorum in manus inimici
PS|77|62|et conclusit in gladio populum suum et hereditatem suam sprevit
PS|77|63|iuvenes eorum comedit ignis et virgines eorum non sunt lamentatae
PS|77|64|sacerdotes eorum in gladio ceciderunt et viduae eorum non plorabuntur
PS|77|65|et excitatus est tamquam dormiens Dominus tamquam potens crapulatus a vino
PS|77|66|et percussit inimicos suos in posteriora obprobrium sempiternum dedit illis
PS|77|67|et reppulit tabernaculum Ioseph et tribum Effrem non elegit
PS|77|68|et elegit tribum Iuda montem Sion quem dilexit
PS|77|69|et aedificavit sicut unicornium sanctificium suum in terra quam fundavit in saecula
PS|77|70|et elegit David servum suum et sustulit eum de gregibus ovium de post fetantes accepit eum
PS|77|71|pascere Iacob servum suum et Israhel hereditatem suam
PS|77|72|et pavit eos in innocentia cordis sui et in intellectibus manuum suarum deduxit eos
PS|78|1|psalmus Asaph Deus venerunt gentes in hereditatem tuam polluerunt templum sanctum tuum posuerunt Hierusalem in pomorum custodiam
PS|78|2|posuerunt morticina servorum tuorum escas volatilibus caeli carnes sanctorum tuorum bestiis terrae
PS|78|3|effuderunt sanguinem ipsorum tamquam aquam in circuitu Hierusalem et non erat qui sepeliret
PS|78|4|facti sumus obprobrium vicinis nostris subsannatio et inlusio his qui circum nos sunt
PS|78|5|usquequo Domine irasceris in finem accendetur velut ignis zelus tuus
PS|78|6|effunde iram tuam in gentes quae te non noverunt et in regna quae nomen tuum non invocaverunt
PS|78|7|quia comederunt Iacob et locum eius desolaverunt
PS|78|8|ne memineris iniquitatum nostrarum antiquarum cito anticipent nos misericordiae tuae quia pauperes facti sumus nimis
PS|78|9|adiuva nos Deus salutaris noster propter gloriam nominis tui Domine libera nos et propitius esto peccatis nostris propter nomen tuum
PS|78|10|ne forte dicant in gentibus ubi est Deus eorum et innotescat in nationibus coram oculis nostris ultio sanguinis servorum tuorum qui effusus est
PS|78|11|introeat in conspectu tuo gemitus conpeditorum secundum magnitudinem brachii tui posside filios mortificatorum
PS|78|12|et redde vicinis nostris septuplum in sinu eorum inproperium ipsorum quod exprobraverunt tibi Domine
PS|78|13|nos autem populus tuus et oves pascuae tuae confitebimur tibi in saeculum in generationem et generationem adnuntiabimus laudem tuam
PS|79|1|in finem pro his qui commutabuntur testimonium Asaph psalmus
PS|79|2|qui regis Israhel intende qui deducis tamquam oves Ioseph qui sedes super cherubin manifestare
PS|79|3|coram Effraim et Beniamin et Manasse excita potentiam tuam et veni ut salvos facias nos
PS|79|4|Deus converte nos et ostende faciem tuam et salvi erimus
PS|79|5|Domine Deus virtutum quousque irasceris super orationem servi tui
PS|79|6|cibabis nos pane lacrimarum et potum dabis nobis in lacrimis in mensura
PS|79|7|posuisti nos in contradictionem vicinis nostris et inimici nostri subsannaverunt nos
PS|79|8|Deus virtutum converte nos et ostende faciem tuam et salvi erimus
PS|79|9|vineam de Aegypto transtulisti eiecisti gentes et plantasti eam
PS|79|10|dux itineris fuisti in conspectu eius et plantasti radices eius et implevit terram
PS|79|11|operuit montes umbra eius et arbusta eius cedros Dei
PS|79|12|extendit palmites suos usque ad mare et usque ad Flumen propagines eius
PS|79|13|ut quid destruxisti maceriam eius et vindemiant eam omnes qui praetergrediuntur viam
PS|79|14|exterminavit eam aper de silva et singularis ferus depastus est eam
PS|79|15|Deus virtutum convertere respice de caelo et vide et visita vineam istam
PS|79|16|et perfice eam quam plantavit dextera tua et super filium quem confirmasti tibi
PS|79|17|incensa igni et suffossa ab increpatione vultus tui peribunt
PS|79|18|fiat manus tua super virum dexterae tuae et super filium hominis quem confirmasti tibi
PS|79|19|et non discedimus a te vivificabis nos et nomen tuum invocabimus
PS|79|20|Domine Deus virtutum converte nos et ostende faciem tuam et salvi erimus
PS|80|1|in finem pro torcularibus Asaph
PS|80|2|exultate Deo adiutori nostro iubilate Deo Iacob
PS|80|3|sumite psalmum et date tympanum psalterium iucundum cum cithara
PS|80|4|bucinate in neomenia tuba in insigni die sollemnitatis nostrae
PS|80|5|quia praeceptum Israhel est et iudicium Dei Iacob
PS|80|6|testimonium in Ioseph posuit illud cum exiret de terra Aegypti linguam quam non noverat audivit
PS|80|7|devertit ab oneribus dorsum eius manus eius in cofino servierunt
PS|80|8|in tribulatione invocasti me et liberavi te exaudivi te in abscondito tempestatis probavi te apud aquam Contradictionis diapsalma
PS|80|9|audi populus meus et contestabor te Israhel si audias me
PS|80|10|non erit in te deus recens nec adorabis deum alienum
PS|80|11|ego enim sum Dominus Deus tuus qui eduxi te de terra Aegypti dilata os tuum et implebo illud
PS|80|12|et non audivit populus meus vocem meam et Israhel non intendit mihi
PS|80|13|et dimisi illos secundum desideria cordis eorum ibunt in adinventionibus suis
PS|80|14|si populus meus audisset me Israhel si in viis meis ambulasset
PS|80|15|pro nihilo forsitan inimicos eorum humiliassem et super tribulantes eos misissem manum meam
PS|80|16|inimici Domini mentiti sunt ei et erit tempus eorum in saeculo
PS|80|17|et cibavit illos ex adipe frumenti et de petra melle saturavit illos
PS|81|1|psalmus Asaph Deus stetit in synagoga deorum in medio autem Deus deiudicat
PS|81|2|usquequo iudicatis iniquitatem et facies peccatorum sumitis diapsalma
PS|81|3|iudicate egenum et pupillum humilem et pauperem iustificate
PS|81|4|eripite pauperem et egenum de manu peccatoris liberate
PS|81|5|nescierunt neque intellexerunt in tenebris ambulant movebuntur omnia fundamenta terrae
PS|81|6|ego dixi dii estis et filii Excelsi omnes
PS|81|7|vos autem sicut homines moriemini et sicut unus de principibus cadetis
PS|81|8|surge Deus iudica terram quoniam tu hereditabis in omnibus gentibus
PS|82|1|canticum psalmi Asaph
PS|82|2|Deus quis similis erit tibi ne taceas neque conpescaris Deus
PS|82|3|quoniam ecce inimici tui sonaverunt et qui oderunt te extulerunt caput
PS|82|4|super populum tuum malignaverunt consilium et cogitaverunt adversus sanctos tuos
PS|82|5|dixerunt venite et disperdamus eos de gente et non memoretur nomen Israhel ultra
PS|82|6|quoniam cogitaverunt unianimiter simul adversum te testamentum disposuerunt
PS|82|7|tabernacula Idumeorum et Ismahelitae Moab et Aggareni
PS|82|8|Gebal et Ammon et Amalech alienigenae cum habitantibus Tyrum
PS|82|9|etenim Assur venit cum illis facti sunt in adiutorium filiis Loth diapsalma
PS|82|10|fac illis sicut Madiam et Sisarae sicut Iabin in torrente Cison
PS|82|11|disperierunt in Endor facti sunt ut stercus terrae
PS|82|12|pone principes eorum sicut Oreb et Zeb et Zebee et Salmana omnes principes eorum
PS|82|13|qui dixerunt hereditate possideamus sanctuarium Dei
PS|82|14|Deus meus pone illos ut rotam sicut stipulam ante faciem venti
PS|82|15|sicut ignis qui conburit silvam sicut flamma conburens montes
PS|82|16|ita persequeris illos in tempestate tua et in ira tua turbabis eos
PS|82|17|imple facies illorum ignominia et quaerent nomen tuum Domine
PS|82|18|erubescant et conturbentur in saeculum saeculi et confundantur et pereant
PS|82|19|et cognoscant quia nomen tibi Dominus tu solus Altissimus in omni terra
PS|83|1|in finem pro torcularibus filiis Core psalmus
PS|83|2|quam dilecta tabernacula tua Domine virtutum
PS|83|3|concupiscit et defecit anima mea in atria Domini cor meum et caro mea exultavit in Deum vivum
PS|83|4|etenim passer invenit %sibi; domum et turtur nidum sibi ubi ponat pullos suos altaria tua Domine virtutum rex meus et Deus meus
PS|83|5|beati qui habitant in domo tua in saecula saeculorum laudabunt te diapsalma
PS|83|6|beatus vir cui est auxilium abs te ascensiones in corde suo disposuit
PS|83|7|in valle lacrimarum in loco quem posuit
PS|83|8|etenim benedictiones dabit legis dator ibunt de virtute in virtutem videbitur Deus deorum in Sion
PS|83|9|Domine Deus virtutum exaudi orationem meam auribus percipe Deus Iacob diapsalma
PS|83|10|protector noster aspice Deus et respice in faciem christi tui
PS|83|11|quia melior est dies una in atriis tuis super milia elegi abiectus esse in domo Dei mei magis quam habitare in tabernaculis peccatorum
PS|83|12|quia misericordiam et veritatem %diligit; Deus gratiam et gloriam dabit Dominus
PS|83|13|non privabit bonis eos qui ambulant in innocentia Domine virtutum beatus vir qui sperat in te
PS|84|1|in finem filiis Core psalmus
PS|84|2|benedixisti Domine terram tuam avertisti captivitatem Iacob
PS|84|3|remisisti iniquitates plebis tuae operuisti omnia peccata eorum diapsalma
PS|84|4|mitigasti omnem iram tuam avertisti ab ira indignationis tuae
PS|84|5|converte nos Deus salutum nostrarum et averte iram tuam a nobis
PS|84|6|numquid in aeternum irasceris nobis aut extendes iram tuam a generatione in generationem
PS|84|7|Deus tu conversus vivificabis nos et plebs tua laetabitur in te
PS|84|8|ostende nobis Domine misericordiam tuam et salutare tuum da nobis
PS|84|9|audiam quid loquatur % in me; Dominus Deus quoniam loquetur pacem in plebem suam et super sanctos suos et in eos qui convertuntur ad cor
PS|84|10|verumtamen prope timentes eum salutare ipsius ut inhabitet gloria in terra nostra
PS|84|11|misericordia et veritas obviaverunt % sibi; iustitia et pax osculatae sunt
PS|84|12|veritas de terra orta est et iustitia de caelo prospexit
PS|84|13|etenim Dominus dabit benignitatem et terra nostra dabit fructum suum
PS|84|14|iustitia ante eum ambulabit et ponet in via gressus suos
PS|85|1|oratio ipsi David inclina Domine aurem tuam %et; exaudi me quoniam inops et pauper sum ego
PS|85|2|custodi animam meam quoniam sanctus sum salvum fac servum tuum Deus meus sperantem in te
PS|85|3|miserere mei Domine quoniam ad te clamabo tota die
PS|85|4|laetifica animam servi tui quoniam ad te Domine animam meam levavi
PS|85|5|quoniam tu Domine suavis et mitis et multae misericordiae omnibus invocantibus te
PS|85|6|auribus percipe Domine orationem meam et intende voci orationis meae
PS|85|7|in die tribulationis meae clamavi ad te quia exaudisti me
PS|85|8|non est similis tui in diis Domine et non est secundum opera tua
PS|85|9|omnes gentes quascumque fecisti venient et adorabunt coram te Domine et glorificabunt nomen tuum
PS|85|10|quoniam magnus es tu et faciens mirabilia tu es Deus solus
PS|85|11|deduc me Domine in via tua et ingrediar in veritate tua laetetur cor meum ut timeat nomen tuum
PS|85|12|confitebor tibi Domine Deus meus in toto corde meo et glorificabo nomen tuum in aeternum
PS|85|13|quia misericordia tua magna est super me et eruisti animam meam ex inferno inferiori
PS|85|14|Deus iniqui insurrexerunt super me et synagoga potentium quaesierunt animam meam et non proposuerunt te in conspectu suo
PS|85|15|et tu Domine Deus miserator et misericors patiens et multae misericordiae et verax
PS|85|16|respice in me et miserere mei da imperium tuum puero tuo et salvum fac filium ancillae tuae
PS|85|17|fac mecum signum in bono et videant qui oderunt me et confundantur quoniam tu Domine adiuvasti me et consolatus es me
PS|86|1|filiis Core psalmus cantici fundamenta eius in montibus sanctis
PS|86|2|diligit Dominus portas Sion super omnia tabernacula Iacob
PS|86|3|gloriosa dicta sunt de te civitas Dei diapsalma
PS|86|4|memor ero Raab et Babylonis scientibus me ecce alienigenae et Tyrus et populus Aethiopum hii fuerunt illic
PS|86|5|numquid Sion dicet homo et homo natus est in ea et ipse fundavit eam Altissimus
PS|86|6|Dominus narrabit in scriptura populorum et principum horum qui fuerunt in ea diapsalma
PS|86|7|sicut laetantium omnium habitatio in te
PS|87|1|canticum psalmi filiis Core in finem pro Maeleth ad respondendum intellectus Eman Ezraitae
PS|87|2|Domine Deus salutis meae die clamavi et nocte coram te
PS|87|3|intret in conspectu tuo oratio mea inclina aurem tuam ad precem meam
PS|87|4|quia repleta est malis anima mea et vita mea in inferno adpropinquavit
PS|87|5|aestimatus sum cum descendentibus in lacum factus sum sicut homo sine adiutorio
PS|87|6|inter mortuos liber sicut vulnerati dormientes in sepulchris quorum non es memor amplius et ipsi de manu tua repulsi sunt
PS|87|7|posuerunt me in lacu inferiori in tenebrosis et in umbra mortis
PS|87|8|super me confirmatus est furor tuus et omnes fluctus tuos induxisti super me diapsalma
PS|87|9|longe fecisti notos meos a me posuerunt me abominationem sibi traditus sum et non egrediebar
PS|87|10|oculi mei languerunt prae inopia clamavi ad te Domine tota die expandi ad te manus meas
PS|87|11|numquid mortuis facies mirabilia aut medici suscitabunt et confitebuntur tibi diapsalma
PS|87|12|numquid narrabit aliquis in sepulchro misericordiam tuam et veritatem tuam in perditione
PS|87|13|numquid cognoscentur in tenebris mirabilia tua et iustitia tua in terra oblivionis
PS|87|14|et ego ad te Domine clamavi et mane oratio mea praeveniet te
PS|87|15|ut quid Domine repellis orationem meam avertis faciem tuam a me
PS|87|16|pauper sum ego et in laboribus a iuventute mea exaltatus autem humiliatus sum et conturbatus
PS|87|17|in me transierunt irae tuae et terrores tui conturbaverunt me
PS|87|18|circuierunt me sicut aqua tota die circumdederunt me simul
PS|87|19|elongasti a me amicum et proximum et notos meos a miseria
PS|88|1|intellectus Aethan Ezraitae
PS|88|2|misericordias Domini in aeternum cantabo in generationem et generationem adnuntiabo veritatem tuam in ore meo
PS|88|3|quoniam dixisti in aeternum misericordia aedificabitur in caelis praeparabitur veritas tua in eis;
PS|88|4|disposui testamentum electis meis iuravi David servo meo
PS|88|5|usque in aeternum praeparabo semen tuum et aedificabo in generationem et generationem sedem tuam diapsalma
PS|88|6|confitebuntur caeli mirabilia tua Domine etenim veritatem tuam in ecclesia sanctorum
PS|88|7|quoniam quis in nubibus aequabitur Domino similis erit Domino in filiis Dei
PS|88|8|Deus qui glorificatur in consilio sanctorum magnus et horrendus super omnes qui in circuitu eius sunt
PS|88|9|Domine Deus virtutum quis similis tibi potens es Domine et veritas tua in circuitu tuo
PS|88|10|tu dominaris potestatis maris motum autem fluctuum eius tu mitigas
PS|88|11|tu humiliasti sicut vulneratum superbum in brachio virtutis tuae dispersisti inimicos tuos
PS|88|12|tui sunt caeli et tua est terra orbem terrae et plenitudinem eius tu fundasti
PS|88|13|aquilonem et mare tu creasti Thabor et Hermon in nomine tuo exultabunt
PS|88|14|tuum brachium cum potentia firmetur manus tua et exaltetur dextera tua
PS|88|15|iustitia et iudicium praeparatio sedis tuae misericordia et veritas praecedent faciem tuam
PS|88|16|beatus populus qui scit iubilationem Domine in lumine vultus tui ambulabunt
PS|88|17|et in nomine tuo exultabunt tota die et in iustitia tua exaltabuntur
PS|88|18|quoniam gloria virtutis eorum tu es et in beneplacito tuo exaltabitur cornu nostrum
PS|88|19|quia Domini est adsumptio nostra; et Sancti Israhel regis nostri
PS|88|20|tunc locutus es in visione sanctis tuis et dixisti posui adiutorium in potentem exaltavi electum de plebe mea
PS|88|21|inveni David servum meum in oleo sancto meo linui eum
PS|88|22|manus enim mea auxiliabitur ei et brachium meum confirmabit eum
PS|88|23|nihil proficiet inimicus in eo et filius iniquitatis non adponet nocere eum
PS|88|24|et concidam a facie ipsius inimicos eius et odientes eum in fugam convertam
PS|88|25|et veritas mea et misericordia mea cum ipso et in nomine meo exaltabitur cornu eius
PS|88|26|et ponam in mari manum eius et in fluminibus dexteram eius
PS|88|27|ipse invocabit me pater meus es tu Deus meus et susceptor salutis meae
PS|88|28|et ego primogenitum ponam illum excelsum prae regibus terrae
PS|88|29|in aeternum servabo illi misericordiam meam et testamentum meum fidele ipsi
PS|88|30|et ponam in saeculum saeculi semen eius et thronum eius sicut dies caeli
PS|88|31|si dereliquerint filii eius legem meam et in iudiciis meis non ambulaverint
PS|88|32|si iustitias meas profanaverint et mandata mea non custodierint
PS|88|33|visitabo in virga iniquitates eorum et in verberibus peccata eorum
PS|88|34|misericordiam autem meam non dispergam ab eo neque nocebo in veritate mea
PS|88|35|neque profanabo testamentum meum et quae procedunt de labiis meis non faciam irrita
PS|88|36|semel iuravi in sancto meo si David mentiar
PS|88|37|semen eius in aeternum manebit
PS|88|38|et thronus eius sicut sol in conspectu meo et sicut luna perfecta in aeternum et testis in caelo fidelis diapsalma
PS|88|39|tu vero reppulisti et despexisti distulisti christum tuum
PS|88|40|evertisti testamentum servi tui profanasti in terram sanctuarium eius
PS|88|41|destruxisti omnes sepes eius posuisti firmamenta eius formidinem
PS|88|42|diripuerunt eum omnes transeuntes viam factus est obprobrium vicinis suis
PS|88|43|exaltasti dexteram deprimentium eum laetificasti omnes inimicos eius
PS|88|44|avertisti adiutorium gladii eius et non es auxiliatus ei in bello
PS|88|45|destruxisti eum a mundatione sedem eius in terram conlisisti
PS|88|46|minorasti dies temporis eius perfudisti eum confusione diapsalma
PS|88|47|usquequo Domine avertis in finem exardescet sicut ignis ira tua
PS|88|48|memorare quae mea substantia numquid enim vane constituisti omnes filios hominum
PS|88|49|quis est homo qui vivet et non videbit mortem eruet animam suam de manu inferi diapsalma
PS|88|50|ubi sunt misericordiae tuae antiquae Domine sicut iurasti David in veritate tua
PS|88|51|memor esto Domine obprobrii servorum tuorum quod continui in sinu meo multarum gentium
PS|88|52|quod exprobraverunt inimici tui Domine quod exprobraverunt commutationem christi tui
PS|88|53|benedictus Dominus in aeternum fiat fiat
PS|89|1|oratio Mosi hominis Dei Domine refugium tu factus es nobis in generatione et generatione
PS|89|2|priusquam montes fierent et formaretur terra et orbis a saeculo usque in saeculum tu es Deus
PS|89|3|ne avertas hominem in humilitatem et dixisti convertimini filii hominum
PS|89|4|quoniam mille anni ante oculos tuos tamquam dies hesterna quae praeteriit et custodia in nocte
PS|89|5|quae pro nihilo habentur eorum anni erunt
PS|89|6|mane sicut herba transeat mane floreat et transeat vespere decidat induret et arescat
PS|89|7|quia defecimus in ira tua et in furore tuo turbati sumus
PS|89|8|posuisti iniquitates nostras in conspectu tuo saeculum nostrum in inluminatione vultus tui
PS|89|9|quoniam omnes dies nostri defecerunt in ira tua defecimus anni nostri sicut aranea meditabantur
PS|89|10|dies annorum nostrorum in ipsis septuaginta anni si autem in potentatibus octoginta anni et amplius eorum labor et dolor quoniam supervenit mansuetudo et corripiemur
PS|89|11|quis novit potestatem irae tuae et prae timore tuo iram tuam
PS|89|12|dinumerare dexteram tuam sic notam fac et conpeditos corde in sapientia
PS|89|13|convertere Domine usquequo et deprecabilis esto super servos tuos
PS|89|14|repleti sumus mane misericordia tua et exultavimus et delectati sumus in omnibus diebus nostris
PS|89|15|laetati sumus pro diebus quibus nos humiliasti annis quibus vidimus mala
PS|89|16|et respice in servos tuos et in opera tua et dirige filios eorum
PS|89|17|et sit splendor Domini Dei nostri super nos et opera manuum nostrarum dirige super nos et opus manuum nostrarum dirige;
PS|90|1|laus cantici David qui habitat in adiutorio Altissimi in protectione Dei caeli commorabitur
PS|90|2|dicet Domino susceptor meus es tu et refugium meum Deus meus sperabo in eum
PS|90|3|quoniam ipse liberabit me de laqueo venantium et a verbo aspero
PS|90|4|in scapulis suis obumbrabit te et sub pinnis eius sperabis
PS|90|5|scuto circumdabit te veritas eius non timebis a timore nocturno
PS|90|6|a sagitta volante in die a negotio perambulante in tenebris ab incursu et daemonio meridiano
PS|90|7|cadent a latere tuo mille et decem milia a dextris tuis ad te autem non adpropinquabit
PS|90|8|verumtamen oculis tuis considerabis et retributionem peccatorum videbis
PS|90|9|quoniam tu Domine spes mea Altissimum posuisti refugium tuum
PS|90|10|non accedent ad te mala et flagellum non adpropinquabit tabernaculo tuo
PS|90|11|quoniam angelis suis mandabit de te ut custodiant te in omnibus viis tuis
PS|90|12|in manibus portabunt te ne forte offendas ad lapidem pedem tuum
PS|90|13|super aspidem et basiliscum ambulabis %et; conculcabis leonem et draconem
PS|90|14|quoniam in me speravit et liberabo eum protegam eum quia cognovit nomen meum
PS|90|15|clamabit ad me et exaudiam eum cum ipso sum in tribulatione eripiam eum et clarificabo eum
PS|90|16|longitudine dierum replebo eum et ostendam illi salutare meum
PS|91|1|psalmus cantici in die sabbati
PS|91|2|bonum est confiteri Domino et psallere nomini tuo Altissime
PS|91|3|ad adnuntiandum mane misericordiam tuam et veritatem tuam per noctem
PS|91|4|in decacordo psalterio cum cantico in cithara
PS|91|5|quia delectasti me Domine in factura tua et in operibus manuum tuarum exultabo
PS|91|6|quam magnificata sunt opera tua Domine nimis profundae factae sunt cogitationes tuae
PS|91|7|vir insipiens non cognoscet et stultus non intelleget haec
PS|91|8|cum exorti fuerint peccatores sicut faenum et apparuerint omnes qui operantur iniquitatem ut intereant in saeculum %saeculi;
PS|91|9|tu autem Altissimus in aeternum Domine
PS|91|10|quoniam ecce inimici tui Domine; quoniam ecce inimici tui peribunt et dispergentur omnes qui operantur iniquitatem
PS|91|11|et exaltabitur sicut unicornis cornu meum et senectus mea in misericordia uberi
PS|91|12|et despexit oculus meus inimicis meis et insurgentibus in me malignantibus audiet auris mea
PS|91|13|iustus ut palma florebit ut cedrus Libani multiplicabitur
PS|91|14|plantati in domo Domini in atriis Dei nostri florebunt
PS|91|15|adhuc multiplicabuntur in senecta uberi et bene patientes erunt
PS|91|16|ut adnuntient quoniam rectus Dominus Deus noster et non est iniquitas in eo
PS|92|1|laus cantici David in die ante sabbatum quando inhabitata est terra Dominus regnavit decore indutus est indutus est Dominus fortitudine et praecinxit se etenim firmavit orbem terrae qui non commovebitur
PS|92|2|parata sedis tua ex tunc a saeculo tu es
PS|92|3|elevaverunt flumina Domine elevaverunt flumina vocem suam elevabunt flumina fluctus suos;
PS|92|4|a vocibus aquarum multarum mirabiles elationes maris mirabilis in altis Dominus
PS|92|5|testimonia tua credibilia facta sunt nimis domum tuam decet sanctitudo Domine in longitudine dierum
PS|93|1|psalmus David quarta sabbati Deus ultionum Dominus Deus ultionum libere egit
PS|93|2|exaltare qui iudicas terram redde retributionem superbis
PS|93|3|usquequo peccatores Domine usquequo peccatores gloriabuntur
PS|93|4|effabuntur et loquentur iniquitatem loquentur omnes qui operantur iniustitiam
PS|93|5|populum tuum Domine humiliaverunt et hereditatem tuam vexaverunt
PS|93|6|viduam et advenam interfecerunt et pupillos occiderunt
PS|93|7|et dixerunt non videbit Dominus nec intelleget Deus Iacob
PS|93|8|intellegite qui insipientes estis in populo et stulti aliquando sapite
PS|93|9|qui plantavit aurem non audiet aut qui finxit oculum non considerat
PS|93|10|qui corripit gentes non arguet qui docet hominem scientiam
PS|93|11|Dominus scit cogitationes hominum quoniam vanae sunt
PS|93|12|beatus homo quem tu erudieris Domine et de lege tua docueris eum
PS|93|13|ut mitiges ei a diebus malis donec fodiatur peccatori fovea
PS|93|14|quia non repellet Dominus plebem suam et hereditatem suam non derelinquet
PS|93|15|quoadusque iustitia convertatur in iudicium et qui iuxta illam omnes qui recto sunt corde diapsalma
PS|93|16|quis consurget mihi adversus malignantes aut quis stabit mecum adversus operantes iniquitatem
PS|93|17|nisi quia Dominus adiuvit me paulo minus habitavit in inferno anima mea
PS|93|18|si dicebam motus est pes meus misericordia tua Domine adiuvabat me
PS|93|19|secundum multitudinem dolorum meorum in corde meo consolationes tuae laetificaverunt animam meam
PS|93|20|numquid aderit tibi sedis iniquitatis qui fingis dolorem in praecepto
PS|93|21|captabunt in animam iusti et sanguinem innocentem condemnabunt
PS|93|22|et factus est Dominus mihi in refugium et Deus meus in adiutorem spei meae
PS|93|23|et reddet illis iniquitatem ipsorum et in malitia eorum disperdet eos disperdet illos Dominus Deus noster
PS|94|1|laus cantici David venite exultemus Domino iubilemus Deo salutari nostro
PS|94|2|praeoccupemus faciem eius in confessione et in psalmis iubilemus ei
PS|94|3|quoniam Deus magnus Dominus et rex magnus super omnes deos
PS|94|4|quia in manu eius fines terrae et altitudines montium ipsius sunt
PS|94|5|quoniam ipsius est mare et ipse fecit illud et siccam manus eius formaverunt
PS|94|6|venite adoremus et procidamus et ploremus ante Dominum qui fecit nos
PS|94|7|quia ipse est Deus noster et nos populus pascuae eius et oves manus eius
PS|94|8|hodie si vocem eius audieritis nolite obdurare corda vestra
PS|94|9|sicut in inritatione secundum diem temptationis in deserto ubi temptaverunt me patres vestri probaverunt me; et viderunt opera mea
PS|94|10|quadraginta annis offensus fui generationi illi et dixi semper errant corde
PS|94|11|et isti non cognoverunt vias meas ut iuravi in ira mea si intrabunt in requiem meam
PS|95|1|quando domus aedificabatur post captivitatem canticum huic David cantate Domino canticum novum cantate Domino omnis terra
PS|95|2|cantate Domino benedicite nomini eius adnuntiate diem de die salutare eius
PS|95|3|adnuntiate inter gentes gloriam eius in omnibus populis mirabilia eius
PS|95|4|quoniam magnus Dominus et laudabilis valde terribilis est super omnes deos
PS|95|5|quoniam omnes dii gentium daemonia at vero Dominus caelos fecit
PS|95|6|confessio et pulchritudo in conspectu eius sanctimonia et magnificentia in sanctificatione eius
PS|95|7|adferte Domino patriae gentium adferte Domino gloriam et honorem
PS|95|8|adferte Domino gloriam nomini eius tollite hostias et introite in atria eius
PS|95|9|adorate Dominum in atrio sancto eius commoveatur a facie eius universa terra
PS|95|10|dicite in gentibus quia Dominus regnavit etenim correxit orbem qui non movebitur iudicabit populos in aequitate
PS|95|11|laetentur caeli et exultet terra commoveatur mare et plenitudo eius
PS|95|12|gaudebunt campi et omnia quae in eis sunt tunc exultabunt omnia ligna silvarum
PS|95|13|a facie Domini quia venit quoniam venit iudicare terram iudicabit orbem terrae in aequitate et populos in veritate sua
PS|96|1|huic David quando terra eius restituta est Dominus regnavit exultet terra laetentur insulae multae
PS|96|2|nubes et caligo in circuitu eius iustitia et iudicium correctio sedis eius
PS|96|3|ignis ante ipsum praecedet et inflammabit in circuitu inimicos eius
PS|96|4|adluxerunt fulgora eius orbi terrae vidit et commota est terra
PS|96|5|montes sicut cera fluxerunt a facie Domini; a facie Domini omnis terrae
PS|96|6|adnuntiaverunt caeli iustitiam eius et viderunt omnes populi gloriam eius
PS|96|7|confundantur omnes qui adorant sculptilia qui gloriantur in simulacris suis adorate eum omnes angeli eius
PS|96|8|audivit et laetata est Sion et exultaverunt filiae Iudaeae propter iudicia tua Domine
PS|96|9|quoniam tu Dominus Altissimus super omnem terram nimis superexaltatus es super omnes deos
PS|96|10|qui diligitis Dominum odite malum custodit animas sanctorum suorum de manu peccatoris liberabit eos
PS|96|11|lux orta est iusto et rectis corde laetitia
PS|96|12|laetamini iusti in Domino et confitemini memoriae sanctificationis eius
PS|97|1|psalmus David cantate Domino canticum novum quoniam mirabilia fecit salvavit sibi dextera eius et brachium sanctum eius
PS|97|2|notum fecit Dominus salutare suum in conspectu gentium revelavit iustitiam suam
PS|97|3|recordatus est misericordiae suae et veritatem suam domui Israhel viderunt omnes termini terrae salutare Dei nostri
PS|97|4|iubilate Domino omnis terra cantate et exultate et psallite
PS|97|5|psallite Domino in cithara in cithara et voce psalmi
PS|97|6|in tubis ductilibus et voce tubae corneae iubilate in conspectu regis Domini
PS|97|7|moveatur mare et plenitudo eius orbis terrarum et qui habitant in eo
PS|97|8|flumina plaudent manu simul montes exultabunt
PS|97|9|a conspectu Domini quoniam venit iudicare terram iudicabit orbem terrarum in iustitia et populos in aequitate
PS|98|1|psalmus David Dominus regnavit irascantur populi qui sedet super cherubin moveatur terra
PS|98|2|Dominus in Sion magnus et excelsus est super omnes populos
PS|98|3|confiteantur nomini tuo magno quoniam terribile et sanctum est
PS|98|4|et honor regis iudicium diligit tu parasti directiones iudicium et iustitiam in Iacob tu fecisti
PS|98|5|exaltate Dominum Deum nostrum et adorate scabillum pedum eius quoniam sanctum est
PS|98|6|Moses et Aaron in sacerdotibus eius et Samuhel inter eos qui invocant nomen eius invocabant Dominum et ipse exaudiebat illos
PS|98|7|in columna nubis loquebatur ad eos custodiebant testimonia eius et praeceptum quod dedit illis
PS|98|8|Domine Deus noster tu exaudiebas illos Deus tu propitius fuisti eis et ulciscens in omnes adinventiones eorum
PS|98|9|exaltate Dominum Deum nostrum et adorate in monte sancto eius quoniam sanctus Dominus Deus noster
PS|99|1|psalmus in confessione
PS|99|2|iubilate Domino omnis terra servite Domino in laetitia introite in conspectu eius in exultatione
PS|99|3|scitote quoniam Dominus ipse est Deus ipse fecit nos et non ipsi nos populus eius et oves pascuae eius
PS|99|4|introite portas eius in confessione atria eius in hymnis confitemini illi laudate nomen eius
PS|99|5|quoniam suavis Dominus in aeternum misericordia eius et usque in generationem et generationem veritas eius
PS|100|1|David psalmus misericordiam et iudicium cantabo tibi Domine psallam
PS|100|2|et intellegam in via inmaculata quando venies ad me perambulabam in innocentia cordis mei in medio domus meae
PS|100|3|non proponebam ante oculos meos rem iniustam facientes praevaricationes odivi non adhesit mihi
PS|100|4|cor pravum declinante a me maligno non cognoscebam
PS|100|5|detrahentem secreto proximo suo hunc persequebar superbo oculo et insatiabili corde cum hoc non edebam
PS|100|6|oculi mei ad fideles terrae ut sederent mecum ambulans in via inmaculata hic mihi ministrabat
PS|100|7|non habitabat in medio domus meae qui facit superbiam qui loquitur iniqua non direxit in conspectu oculorum meorum
PS|100|8|in matutino interficiebam omnes peccatores terrae ut disperderem de civitate Domini omnes operantes iniquitatem
PS|101|1|oratio pauperis cum anxius fuerit et coram Domino effuderit precem suam
PS|101|2|Domine exaudi orationem meam et clamor meus ad te veniat
PS|101|3|non avertas faciem tuam a me in quacumque die tribulor inclina ad me aurem tuam in quacumque die invocavero te velociter exaudi me
PS|101|4|quia defecerunt sicut fumus dies mei et ossa mea sicut gremium aruerunt
PS|101|5|percussum est ut faenum et aruit cor meum quia oblitus sum comedere panem meum
PS|101|6|a voce gemitus mei adhesit os meum carni meae
PS|101|7|similis factus sum pelicano solitudinis factus sum sicut nycticorax in domicilio
PS|101|8|vigilavi et factus sum sicut passer solitarius in tecto
PS|101|9|tota die exprobrabant mihi inimici mei et qui laudabant me adversus me iurabant
PS|101|10|quia cinerem tamquam panem manducavi et poculum meum cum fletu miscebam
PS|101|11|a facie irae et indignationis tuae quia elevans adlisisti me
PS|101|12|dies mei sicut umbra declinaverunt et ego sicut faenum arui
PS|101|13|tu autem Domine in aeternum permanes et memoriale tuum in generationem et generationem
PS|101|14|tu exsurgens misereberis Sion quia tempus miserendi eius quia venit tempus
PS|101|15|quoniam placuerunt servis tuis lapides eius et terrae eius miserebuntur
PS|101|16|et timebunt gentes nomen Domini et omnes reges terrae gloriam tuam
PS|101|17|quia aedificabit Dominus Sion et videbitur in gloria sua
PS|101|18|respexit in orationem humilium et non sprevit precem eorum
PS|101|19|scribantur haec in generationem alteram et populus qui creabitur laudabit Dominum
PS|101|20|quia prospexit de excelso sancto suo Dominus de caelo in terram aspexit
PS|101|21|ut audiret gemitum conpeditorum ut solvat filios interemptorum
PS|101|22|ut adnuntiet in Sion nomen Domini et laudem suam in Hierusalem
PS|101|23|in conveniendo populos in unum et reges ut serviant Domino
PS|101|24|respondit ei in via virtutis suae paucitatem dierum meorum nuntia mihi
PS|101|25|ne revoces me in dimidio dierum meorum in generationem et generationem anni tui
PS|101|26|initio tu Domine terram fundasti et opera manuum tuarum sunt caeli
PS|101|27|ipsi peribunt tu autem permanes et omnes sicut vestimentum veterescent et sicut opertorium mutabis eos et mutabuntur
PS|101|28|tu autem idem ipse es et anni tui non deficient
PS|101|29|filii servorum tuorum habitabunt et semen eorum in saeculum dirigetur
PS|102|1|ipsi David benedic anima mea Domino et omnia quae intra me sunt nomini sancto eius
PS|102|2|benedic anima mea Domino et noli oblivisci omnes retributiones eius
PS|102|3|qui propitiatur omnibus iniquitatibus tuis qui sanat omnes infirmitates tuas
PS|102|4|qui redimit de interitu vitam tuam qui coronat te in misericordia et miserationibus
PS|102|5|qui replet in bonis desiderium tuum renovabitur ut aquilae iuventus tua
PS|102|6|faciens misericordias Dominus et iudicium omnibus iniuriam patientibus
PS|102|7|notas fecit vias suas Mosi filiis Israhel voluntates suas
PS|102|8|miserator et misericors Dominus longanimis et multum misericors
PS|102|9|non in perpetuum irascetur neque in aeternum comminabitur
PS|102|10|non secundum peccata nostra fecit nobis nec secundum iniustitias nostras retribuit nobis
PS|102|11|quoniam secundum altitudinem caeli a terra corroboravit misericordiam suam super timentes se
PS|102|12|quantum distat ortus ab occidente longe fecit a nobis iniquitates nostras
PS|102|13|quomodo miseretur pater filiorum misertus est Dominus timentibus se
PS|102|14|quoniam ipse cognovit figmentum nostrum recordatus est quoniam pulvis sumus
PS|102|15|homo sicut faenum dies eius tamquam flos agri sic efflorebit
PS|102|16|quoniam spiritus pertransivit in illo et non subsistet et non cognoscet amplius locum suum
PS|102|17|misericordia autem Domini ab aeterno et usque in aeternum super timentes eum et iustitia illius in filios filiorum
PS|102|18|his qui servant testamentum eius et memores sunt mandatorum ipsius ad faciendum ea
PS|102|19|Dominus in caelo paravit sedem suam et regnum ipsius omnibus dominabitur
PS|102|20|benedicite Domino angeli eius potentes virtute facientes verbum illius ad audiendam vocem sermonum eius
PS|102|21|benedicite Domino omnes virtutes eius ministri eius qui facitis voluntatem eius
PS|102|22|benedicite Domino omnia opera eius in omni loco dominationis ipsius benedic anima mea Domino
PS|103|1|ipsi David benedic anima mea Domino Domine Deus meus magnificatus es vehementer confessionem et decorem induisti
PS|103|2|amictus lumine sicut vestimento extendens caelum sicut pellem
PS|103|3|qui tegis in aquis superiora eius qui ponis nubem ascensum tuum qui ambulas super pinnas ventorum
PS|103|4|qui facis angelos tuos spiritus et ministros tuos ignem urentem
PS|103|5|qui fundasti terram super stabilitatem suam non inclinabitur in saeculum saeculi
PS|103|6|abyssus sicut vestimentum amictus eius super montes stabunt aquae
PS|103|7|ab increpatione tua fugient a voce tonitrui tui formidabunt
PS|103|8|ascendunt montes et descendunt campi in locum quem fundasti eis
PS|103|9|terminum posuisti quem non transgredientur neque convertentur operire terram
PS|103|10|qui emittis fontes in convallibus inter medium montium pertransibunt aquae
PS|103|11|potabunt omnes bestiae agri expectabunt onagri in siti sua
PS|103|12|super ea volucres caeli habitabunt de medio petrarum dabunt vocem
PS|103|13|rigans montes de superioribus suis de fructu operum tuorum satiabitur terra
PS|103|14|producens faenum iumentis et herbam servituti hominum ut educas panem de terra
PS|103|15|et vinum laetificat cor hominis ut exhilaret faciem in oleo et panis cor hominis confirmat
PS|103|16|saturabuntur ligna campi et cedri Libani quas plantavit
PS|103|17|illic passeres nidificabunt erodii domus dux est eorum
PS|103|18|montes excelsi cervis petra refugium erinaciis
PS|103|19|fecit lunam in tempora sol cognovit occasum suum
PS|103|20|posuisti tenebras et facta est nox in ipsa pertransibunt omnes bestiae silvae
PS|103|21|catuli leonum rugientes ut rapiant et quaerant a Deo escam sibi
PS|103|22|ortus est sol et congregati sunt et in cubilibus suis conlocabuntur
PS|103|23|exibit homo ad opus suum et ad operationem suam usque ad vesperum
PS|103|24|quam magnificata sunt opera tua Domine omnia in sapientia fecisti impleta est terra possessione tua
PS|103|25|hoc mare magnum et spatiosum manibus; illic reptilia quorum non est numerus animalia pusilla cum magnis
PS|103|26|illic naves pertransibunt draco iste quem formasti ad inludendum ei
PS|103|27|omnia a te expectant ut des illis escam in tempore
PS|103|28|dante te illis colligent aperiente te manum tuam omnia implebuntur bonitate
PS|103|29|avertente autem te faciem turbabuntur auferes spiritum eorum et deficient et in pulverem suum revertentur
PS|103|30|emittes spiritum tuum et creabuntur et renovabis faciem terrae
PS|103|31|sit gloria Domini in saeculum laetabitur Dominus in operibus suis
PS|103|32|qui respicit terram et facit eam tremere qui tangit montes et fumigant
PS|103|33|cantabo Domino in vita mea psallam Deo meo quamdiu sum
PS|103|34|iucundum sit ei eloquium meum ego vero delectabor in Domino
PS|103|35|deficiant peccatores a terra et iniqui ita ut non sint benedic anima mea Domino
PS|104|1|alleluia confitemini Domino et invocate nomen eius adnuntiate inter gentes opera eius
PS|104|2|cantate ei et psallite ei narrate omnia mirabilia eius
PS|104|3|laudamini in nomine sancto eius laetetur cor quaerentium Dominum
PS|104|4|quaerite Dominum et confirmamini quaerite faciem eius semper
PS|104|5|mementote mirabilium eius quae fecit prodigia eius et iudicia oris eius
PS|104|6|semen Abraham servi eius filii Iacob electi eius
PS|104|7|ipse Dominus Deus noster in universa terra iudicia eius
PS|104|8|memor fuit in saeculum testamenti sui verbi quod mandavit in mille generationes
PS|104|9|quod disposuit ad Abraham et iuramenti sui ad Isaac
PS|104|10|et statuit illud Iacob in praeceptum et Israhel in testamentum aeternum
PS|104|11|dicens tibi dabo terram Chanaan funiculum hereditatis vestrae
PS|104|12|cum essent numero breves paucissimos et incolas eius
PS|104|13|et pertransierunt de gente in gentem et de regno ad populum alterum
PS|104|14|non reliquit hominem nocere eis et corripuit pro eis reges
PS|104|15|nolite tangere christos meos et in prophetis meis nolite malignari
PS|104|16|et vocavit famem super terram omne firmamentum panis contrivit
PS|104|17|misit ante eos virum in servum venundatus est Ioseph
PS|104|18|humiliaverunt in conpedibus pedes eius ferrum pertransiit anima eius
PS|104|19|donec veniret verbum eius eloquium Domini inflammavit eum
PS|104|20|misit rex et solvit eum princeps populorum et dimisit eum
PS|104|21|constituit eum dominum domus suae et principem omnis possessionis suae
PS|104|22|ut erudiret principes eius sicut semet ipsum et senes eius prudentiam doceret
PS|104|23|et intravit Israhel in Aegyptum et Iacob accola fuit in terra Cham
PS|104|24|et auxit populum eius vehementer et firmavit eum super inimicos eius
PS|104|25|convertit cor eorum ut odirent populum eius ut dolum facerent in servos eius
PS|104|26|misit Mosen servum suum Aaron quem elegit ipsum
PS|104|27|posuit in eis verba signorum suorum et prodigiorum in terra Cham
PS|104|28|misit tenebras et obscuravit et non exacerbavit sermones suos
PS|104|29|convertit aquas eorum in sanguinem et occidit pisces eorum
PS|104|30|dedit terra eorum ranas in penetrabilibus regum ipsorum
PS|104|31|dixit et venit cynomia et scinifes in omnibus finibus eorum
PS|104|32|posuit pluvias eorum grandinem ignem conburentem in terra ipsorum
PS|104|33|et percussit vineas eorum et ficulneas eorum et contrivit lignum finium eorum
PS|104|34|dixit et venit lucusta et bruchus cuius non erat numerus
PS|104|35|et comedit omne faenum in terra eorum et comedit omnem fructum terrae eorum
PS|104|36|et percussit omne primogenitum in terra eorum primitias omnis laboris eorum
PS|104|37|et eduxit eos in argento et auro et non erat in tribubus eorum infirmus
PS|104|38|laetata est Aegyptus in profectione eorum quia incubuit timor eorum super eos
PS|104|39|expandit nubem in protectionem eorum et ignem ut luceret eis per noctem
PS|104|40|petierunt et venit coturnix et panem caeli saturavit eos
PS|104|41|disrupit petram et fluxerunt aquae abierunt in sicco flumina
PS|104|42|quoniam memor fuit verbi sancti sui quod habuit ad Abraham puerum suum
PS|104|43|et eduxit populum suum in exultatione %et; electos suos in laetitia
PS|104|44|et dedit illis regiones gentium et labores populorum possederunt
PS|104|45|ut custodiant iustificationes eius et legem eius requirant
PS|105|1|alleluia confitemini Domino quoniam bonus quoniam in saeculum misericordia eius
PS|105|2|quis loquetur potentias Domini auditas faciet omnes laudes eius
PS|105|3|beati qui custodiunt iudicium et faciunt iustitiam in omni tempore
PS|105|4|memento nostri Domine in beneplacito populi tui visita nos in salutari tuo
PS|105|5|ad videndum in bonitate electorum tuorum ad laetandum in laetitia gentis tuae et lauderis cum hereditate tua
PS|105|6|peccavimus cum patribus nostris iniuste egimus iniquitatem fecimus
PS|105|7|patres nostri in Aegypto non intellexerunt mirabilia tua non fuerunt memores multitudinis misericordiae tuae et inritaverunt ascendentes in mare mare; Rubrum
PS|105|8|et salvavit eos propter nomen suum ut notam faceret potentiam suam
PS|105|9|et increpuit mare Rubrum et exsiccatum est et deduxit eos in abyssis sicut in deserto
PS|105|10|et salvavit eos de manu odientium et redemit eos de manu inimici
PS|105|11|et operuit aqua tribulantes eos unus ex eis non remansit
PS|105|12|et crediderunt in verbis eius et laudaverunt laudem eius
PS|105|13|cito fecerunt obliti sunt operum eius non sustinuerunt consilium eius
PS|105|14|et concupierunt concupiscentiam in deserto et temptaverunt Deum in inaquoso
PS|105|15|et dedit eis petitionem ipsorum et misit saturitatem in anima eorum
PS|105|16|et inritaverunt Mosen in castris Aaron sanctum Domini
PS|105|17|aperta est terra et degluttivit Dathan et operuit super congregationem Abiron
PS|105|18|et exarsit ignis in synagoga eorum flamma conbusit peccatores
PS|105|19|et fecerunt vitulum in Choreb et adoraverunt sculptile
PS|105|20|et mutaverunt gloriam suam in similitudine vituli comedentis faenum
PS|105|21|obliti sunt Deum qui salvavit eos qui fecit magnalia in Aegypto
PS|105|22|mirabilia in terra Cham terribilia in mari Rubro
PS|105|23|et dixit ut disperderet eos si non Moses electus eius stetisset in confractione in conspectu eius ut averteret iram eius ne disperderet eos
PS|105|24|et pro nihilo habuerunt terram desiderabilem non crediderunt verbo eius
PS|105|25|et murmurabant in tabernaculis suis non exaudierunt vocem Domini
PS|105|26|et elevavit manum suam super eos ut prosterneret eos in deserto
PS|105|27|et ut deiceret semen eorum in nationibus et dispergeret eos in regionibus
PS|105|28|et initiati sunt Beelphegor et comederunt sacrificia mortuorum
PS|105|29|et inritaverunt eum in adinventionibus suis et multiplicata est in eis ruina
PS|105|30|et stetit Finees et placavit et cessavit quassatio
PS|105|31|et reputatum est ei in iustitiam in generatione et generationem usque in sempiternum
PS|105|32|et inritaverunt ad aquam Contradictionis et vexatus est Moses propter eos
PS|105|33|quia exacerbaverunt spiritum eius et distinxit in labiis suis
PS|105|34|non disperdiderunt gentes quas dixit Dominus illis
PS|105|35|et commixti sunt inter gentes et didicerunt opera eorum
PS|105|36|et servierunt sculptilibus eorum et factum est illis in scandalum
PS|105|37|et immolaverunt filios suos et filias suas daemoniis
PS|105|38|et effuderunt sanguinem innocentem sanguinem filiorum suorum et filiarum suarum; quas sacrificaverunt sculptilibus Chanaan et interfecta est terra in sanguinibus
PS|105|39|et contaminata est in operibus eorum et fornicati sunt in adinventionibus suis
PS|105|40|et iratus est furore Dominus in populo suo et abominatus est hereditatem suam
PS|105|41|et tradidit eos in manus gentium et dominati sunt eorum qui oderant eos
PS|105|42|et tribulaverunt eos inimici eorum et humiliati sunt sub manibus eorum
PS|105|43|saepe liberavit eos ipsi autem exacerbaverunt eum in consilio suo et humiliati sunt in iniquitatibus suis
PS|105|44|et vidit cum tribularentur et audiret orationem eorum
PS|105|45|et memor fuit testamenti sui et paenituit eum secundum multitudinem misericordiae suae
PS|105|46|et dedit eos in misericordias in conspectu omnium qui ceperant eos
PS|105|47|salvos fac nos Domine Deus noster et congrega nos de nationibus ut confiteamur nomini tuo sancto et gloriemur in laude tua
PS|105|48|benedictus Dominus Deus Israhel a saeculo et usque in saeculum et dicet omnis populus fiat fiat
PS|106|1|alleluia confitemini Domino quoniam bonus quoniam in saeculum misericordia eius
PS|106|2|dicant qui redempti sunt a Domino quos redemit de manu inimici de regionibus congregavit eos
PS|106|3|a solis ortu et occasu et ab aquilone et mari
PS|106|4|erraverunt in solitudine in inaquoso viam civitatis habitaculi non invenerunt
PS|106|5|esurientes et sitientes anima eorum in ipsis defecit
PS|106|6|et clamaverunt ad Dominum cum tribularentur et de necessitatibus eorum eripuit eos
PS|106|7|et deduxit eos in viam rectam ut irent in civitatem habitationis
PS|106|8|confiteantur Domino misericordiae eius et mirabilia eius filiis hominum
PS|106|9|quia satiavit animam inanem et animam esurientem satiavit bonis
PS|106|10|sedentes in tenebris et umbra mortis vinctos in mendicitate et ferro
PS|106|11|quia exacerbaverunt eloquia Dei et consilium Altissimi inritaverunt
PS|106|12|et humiliatum est in laboribus cor eorum infirmati sunt nec fuit qui adiuvaret
PS|106|13|et clamaverunt ad Dominum cum tribularentur et de necessitatibus eorum liberavit eos
PS|106|14|et eduxit eos de tenebris et umbra mortis et vincula eorum disrupit
PS|106|15|confiteantur Domino misericordiae eius et mirabilia eius filiis hominum
PS|106|16|quia contrivit portas aereas et vectes ferreos confregit
PS|106|17|suscepit eos de via iniquitatis eorum propter iniustitias enim suas humiliati sunt
PS|106|18|omnem escam abominata est anima eorum et adpropinquaverunt usque ad portas mortis
PS|106|19|et clamaverunt ad Dominum cum tribularentur et de necessitatibus eorum liberavit eos
PS|106|20|misit verbum suum et sanavit eos et eripuit eos de interitionibus eorum
PS|106|21|confiteantur Domino misericordiae eius et mirabilia eius filiis hominum
PS|106|22|et sacrificent sacrificium laudis et adnuntient opera eius in exultatione
PS|106|23|qui descendunt mare in navibus facientes operationem in aquis multis
PS|106|24|ipsi viderunt opera Domini et mirabilia eius in profundo
PS|106|25|dixit et stetit spiritus procellae et exaltati sunt fluctus eius
PS|106|26|ascendunt usque ad caelos et descendunt usque ad abyssos anima eorum in malis tabescebat
PS|106|27|turbati sunt et moti sunt sicut ebrius et omnis sapientia eorum devorata est
PS|106|28|et clamaverunt ad Dominum cum tribularentur et de necessitatibus eorum eduxit eos
PS|106|29|et statuit procellam %eius; in auram et siluerunt fluctus eius
PS|106|30|et laetati sunt quia siluerunt et deduxit eos in portum voluntatis eorum
PS|106|31|confiteantur Domino misericordiae eius et mirabilia eius filiis hominum
PS|106|32|exaltent eum in ecclesia plebis et in cathedra seniorum laudent eum
PS|106|33|posuit flumina in desertum et exitus aquarum in sitim
PS|106|34|terram fructiferam in salsuginem a malitia inhabitantium in ea
PS|106|35|posuit desertum in stagna aquarum et terram sine aqua in exitus aquarum
PS|106|36|et conlocavit illic esurientes et constituerunt civitatem habitationis
PS|106|37|et seminaverunt agros et plantaverunt vineas et fecerunt fructum nativitatis
PS|106|38|et benedixit eis et multiplicati sunt nimis et iumenta eorum non minoravit
PS|106|39|et pauci facti sunt et vexati sunt a tribulatione malorum et dolore
PS|106|40|effusa est contemptio super principes et errare fecit eos in invio et non in via
PS|106|41|et adiuvit pauperem de inopia et posuit sicut oves familias
PS|106|42|videbunt recti et laetabuntur et omnis iniquitas oppilabit os suum
PS|106|43|quis sapiens et custodiet haec et intellegent misericordias Domini
PS|107|1|canticum psalmi David
PS|107|2|paratum cor meum Deus paratum cor meum cantabo et psallam in gloria mea
PS|107|3|exsurge psalterium et cithara exsurgam diluculo
PS|107|4|confitebor tibi in populis Domine et psallam tibi in nationibus
PS|107|5|quia magna super caelos misericordia tua et usque ad nubes veritas tua
PS|107|6|exaltare super caelos Deus et super omnem terram gloria tua
PS|107|7|ut liberentur dilecti tui salvum fac dextera tua et exaudi me
PS|107|8|Deus locutus est in sancto suo exaltabor et dividam Sicima et convallem tabernaculorum dimetiar
PS|107|9|meus est Galaad et meus est Manasse et Effraim susceptio capitis mei Iuda rex meus
PS|107|10|Moab lebes spei meae in Idumeam extendam calciamentum meum mihi alienigenae amici facti sunt
PS|107|11|quis deducet me in civitatem munitam quis deducet me usque in Idumeam
PS|107|12|nonne tu Deus qui reppulisti nos et non exibis Deus in virtutibus nostris
PS|107|13|da nobis auxilium de tribulatione quia vana salus hominis
PS|107|14|in Deo faciemus virtutem et ipse ad nihilum deducet inimicos nostros
PS|108|1|in finem David psalmus
PS|108|2|Deus laudem meam ne tacueris quia os peccatoris et os dolosi super me apertum est
PS|108|3|locuti sunt adversum me lingua dolosa et sermonibus odii circuierunt me et expugnaverunt me gratis
PS|108|4|pro eo ut me diligerent detrahebant mihi ego autem orabam
PS|108|5|et posuerunt adversus me mala pro bonis et odium pro dilectione mea
PS|108|6|constitue super eum peccatorem et diabulus stet a dextris eius
PS|108|7|cum iudicatur exeat condemnatus et oratio eius fiat in peccatum
PS|108|8|fiant dies eius pauci et episcopatum eius accipiat alter
PS|108|9|fiant filii eius orfani et uxor eius vidua
PS|108|10|nutantes transferantur filii eius et mendicent eiciantur de habitationibus suis
PS|108|11|scrutetur fenerator omnem substantiam eius et diripiant alieni labores eius
PS|108|12|non sit illi adiutor nec sit qui misereatur pupillis eius
PS|108|13|fiant nati eius in interitum in generatione una deleatur nomen eius
PS|108|14|in memoriam redeat iniquitas patrum eius in conspectu Domini et peccatum matris eius non deleatur
PS|108|15|fiant contra Dominum semper et dispereat de terra memoria eorum
PS|108|16|pro eo quod non est recordatus facere misericordiam
PS|108|17|et persecutus est hominem inopem et mendicum et conpunctum corde mortificare
PS|108|18|et dilexit maledictionem et veniet ei et noluit benedictionem et elongabitur ab eo et induit maledictionem sicut vestimentum et intravit sicut aqua in interiora eius et sicut oleum in ossibus eius
PS|108|19|fiat ei sicut vestimentum quo operitur et sicut zona qua semper praecingitur
PS|108|20|hoc opus eorum qui detrahunt mihi apud Dominum et qui loquuntur mala adversus animam meam
PS|108|21|et tu Domine Domine fac mecum propter nomen tuum quia suavis misericordia tua libera me
PS|108|22|quia egenus et pauper ego sum et cor meum turbatum est intra me
PS|108|23|sicut umbra cum declinat ablatus sum excussus sum sicut lucustae
PS|108|24|genua mea infirmata sunt a ieiunio et caro mea inmutata est propter oleum
PS|108|25|et ego factus sum obprobrium illis viderunt me moverunt capita sua
PS|108|26|adiuva me Domine Deus meus salvum fac me secundum misericordiam tuam
PS|108|27|et sciant quia manus tua haec tu Domine fecisti eam
PS|108|28|maledicent illi et tu benedices qui insurgunt in me confundantur servus autem tuus laetabitur
PS|108|29|induantur qui detrahunt mihi pudore et operiantur sicut deploide confusione sua
PS|108|30|confitebor Domino nimis in ore meo et in medio multorum laudabo eum
PS|108|31|quia adstetit a dextris pauperis ut salvam faceret a persequentibus animam meam
PS|109|1|David psalmus dixit Dominus Domino meo sede a dextris meis donec ponam inimicos tuos scabillum pedum tuorum
PS|109|2|virgam virtutis tuae emittet Dominus ex Sion dominare in medio inimicorum tuorum
PS|109|3|tecum principium in die virtutis tuae in splendoribus sanctorum ex utero ante luciferum genui te
PS|109|4|iuravit Dominus et non paenitebit eum tu es sacerdos in aeternum secundum ordinem Melchisedech
PS|109|5|Dominus a dextris tuis confregit in die irae suae reges
PS|109|6|iudicabit in nationibus implebit cadavera conquassabit capita in terra multorum
PS|109|7|de torrente in via bibet propterea exaltabit caput
PS|110|1|alleluia reversionis Aggei et Zacchariae confitebor tibi Domine in toto corde meo in consilio iustorum et congregatione
PS|110|2|magna opera Domini exquisita in omnes voluntates eius
PS|110|3|confessio et magnificentia opus eius et iustitia eius manet in saeculum saeculi
PS|110|4|memoriam fecit mirabilium suorum misericors et miserator Dominus
PS|110|5|escam dedit timentibus se memor erit in saeculum testamenti sui
PS|110|6|virtutem operum suorum adnuntiabit populo suo
PS|110|7|ut det illis hereditatem gentium opera manuum eius veritas et iudicium
PS|110|8|fidelia omnia mandata eius confirmata in saeculum saeculi facta in veritate et aequitate
PS|110|9|redemptionem misit populo suo mandavit in aeternum testamentum suum sanctum et terribile nomen eius
PS|110|10|initium sapientiae timor Domini intellectus bonus omnibus facientibus eum laudatio eius manet in saeculum %saeculi;
PS|111|1|alleluia reversionis Aggei et Zacchariae beatus vir qui timet Dominum in mandatis eius volet nimis
PS|111|2|potens in terra erit semen eius generatio rectorum benedicetur
PS|111|3|gloria et divitiae in domo eius et iustitia eius manet in saeculum saeculi
PS|111|4|exortum est in tenebris lumen rectis misericors et miserator et iustus
PS|111|5|iucundus homo qui miseretur et commodat disponet sermones suos in iudicio
PS|111|6|quia in aeternum non commovebitur
PS|111|7|in memoria aeterna erit iustus ab auditione mala non timebit paratum cor eius sperare in Domino
PS|111|8|confirmatum est cor eius non commovebitur donec dispiciat inimicos suos
PS|111|9|dispersit dedit pauperibus iustitia eius manet in saeculum saeculi cornu eius exaltabitur in gloria
PS|111|10|peccator videbit et irascetur dentibus suis fremet et tabescet desiderium peccatorum peribit
PS|112|1|alleluia laudate pueri Dominum laudate nomen Domini
PS|112|2|sit nomen Domini benedictum ex hoc nunc et usque in saeculum
PS|112|3|a solis ortu usque ad occasum laudabile nomen Domini
PS|112|4|excelsus super omnes gentes Dominus super caelos gloria eius
PS|112|5|quis sicut Dominus Deus noster qui in altis habitat
PS|112|6|et humilia respicit in caelo et in terra
PS|112|7|suscitans a terra inopem et de stercore erigens pauperem
PS|112|8|ut conlocet eum cum principibus cum principibus populi sui
PS|112|9|qui habitare facit sterilem in domo matrem filiorum laetantem
PS|113|1|alleluia in exitu Israhel de Aegypto domus Iacob de populo barbaro
PS|113|2|facta est Iudaea sanctificatio eius Israhel potestas eius
PS|113|3|mare vidit et fugit Iordanis conversus est retrorsum
PS|113|4|montes exultaverunt ut arietes colles sicut agni ovium
PS|113|5|quid est tibi mare quod fugisti et tu Iordanis quia conversus es retrorsum
PS|113|6|montes exultastis sicut arietes et colles sicut agni ovium
PS|113|7|a facie Domini mota est terra a facie Dei Iacob
PS|113|8|qui convertit petram in stagna aquarum et rupem in fontes aquarum
PS|113|9|non nobis Domine non nobis sed nomini tuo da gloriam
PS|113|10|super misericordia tua et veritate tua nequando dicant gentes ubi est Deus eorum
PS|113|11|Deus autem noster in caelo omnia quaecumque voluit fecit
PS|113|12|simulacra gentium argentum et aurum opera manuum hominum
PS|113|13|os habent et non loquentur oculos habent et non videbunt
PS|113|14|aures habent et non audient nares habent et non odorabuntur
PS|113|15|manus habent et non palpabunt pedes habent et non ambulabunt non clamabunt in gutture suo
PS|113|16|similes illis fiant qui faciunt ea et omnes qui confidunt in eis
PS|113|17|domus Israhel speravit in Domino adiutor eorum et protector eorum est
PS|113|18|domus Aaron speravit in Domino adiutor eorum et protector eorum est
PS|113|19|qui timent Dominum speraverunt in Domino adiutor eorum et protector eorum est
PS|113|20|Dominus memor fuit nostri et benedixit nobis benedixit domui Israhel benedixit domui Aaron
PS|113|21|benedixit omnibus qui timent Dominum pusillis cum maioribus
PS|113|22|adiciat Dominus super vos super vos et super filios vestros
PS|113|23|benedicti vos Domino qui fecit caelum et terram
PS|113|24|caelum caeli Domino terram autem dedit filiis hominum
PS|113|25|non mortui laudabunt te Domine neque omnes qui descendunt in infernum
PS|113|26|sed nos qui vivimus benedicimus Domino ex hoc nunc et usque in saeculum
PS|114|1|alleluia dilexi quoniam exaudiet Dominus vocem orationis meae
PS|114|2|quia inclinavit aurem suam mihi et in diebus meis invocabo te
PS|114|3|circumdederunt me dolores mortis pericula inferni invenerunt me tribulationem et dolorem inveni
PS|114|4|et nomen Domini invocavi o Domine libera animam meam
PS|114|5|misericors Dominus et iustus et Deus noster miseretur
PS|114|6|custodiens parvulos Dominus humiliatus sum et liberavit me
PS|114|7|convertere anima mea in requiem tuam quia Dominus benefecit tibi
PS|114|8|quia eripuit animam meam de morte oculos meos a lacrimis pedes meos a lapsu
PS|114|9|placebo Domino in regione vivorum
PS|115|1|alleluia credidi propter quod locutus sum ego autem humiliatus sum nimis
PS|115|2|ego dixi in excessu meo omnis homo mendax
PS|115|3|quid retribuam Domino pro omnibus quae retribuit mihi
PS|115|4|calicem salutaris accipiam et nomen Domini invocabo
PS|115|5|vota mea Domino reddam coram omni populo eius
PS|115|6|pretiosa in conspectu Domini mors sanctorum eius
PS|115|7|o Domine quia ego servus tuus ego servus tuus et filius ancillae tuae disrupisti vincula mea
PS|115|8|tibi sacrificabo hostiam laudis et in nomine Domini invocabo
PS|115|9|vota mea Domino reddam in conspectu omnis populi eius
PS|115|10|in atriis domus Domini in medio tui Hierusalem
PS|116|1|alleluia laudate Dominum omnes gentes laudate eum omnes populi
PS|116|2|quoniam confirmata est super nos misericordia eius et veritas Domini manet in saeculum
PS|117|1|alleluia confitemini Domino quoniam bonus quoniam in saeculum misericordia eius
PS|117|2|dicat nunc Israhel quoniam bonus quoniam in saeculum misericordia eius
PS|117|3|dicat nunc domus Aaron quoniam in saeculum misericordia eius
PS|117|4|dicant nunc qui timent Dominum quoniam in saeculum misericordia eius
PS|117|5|de tribulatione invocavi Dominum et exaudivit me in latitudinem Dominus
PS|117|6|Dominus mihi adiutor non timebo quid faciat mihi homo
PS|117|7|Dominus mihi adiutor et ego despiciam inimicos meos
PS|117|8|bonum est confidere in Domino quam confidere in homine
PS|117|9|bonum est sperare in Domino quam sperare in principibus
PS|117|10|omnes gentes circumierunt me et in nomine Domini quia; ultus sum in eos
PS|117|11|circumdantes circumdederunt me in nomine autem Domini quia; ultus sum in eos
PS|117|12|circumdederunt me sicut apes et exarserunt sicut ignis in spinis et in nomine Domini quia; ultus sum in eos
PS|117|13|inpulsus eversus sum ut caderem et Dominus suscepit me
PS|117|14|fortitudo mea et laudatio mea Dominus et factus est mihi in salutem
PS|117|15|vox exultationis et salutis in tabernaculis iustorum
PS|117|16|dextera Domini fecit virtutem dextera Domini exaltavit me dextera Domini fecit virtutem
PS|117|17|non moriar sed vivam et narrabo opera Domini
PS|117|18|castigans castigavit me Dominus et morti non tradidit me
PS|117|19|aperite mihi portas iustitiae ingressus in eas confitebor Domino
PS|117|20|haec porta Domini iusti intrabunt in eam
PS|117|21|confitebor tibi quoniam exaudisti me et factus es mihi in salutem
PS|117|22|lapidem quem reprobaverunt aedificantes hic factus est in caput anguli
PS|117|23|a Domino factum est istud hoc est mirabile in oculis nostris
PS|117|24|haec est dies quam fecit Dominus exultemus et laetemur in ea
PS|117|25|o Domine salvum fac o Domine prosperare
PS|117|26|benedictus qui venturus est in nomine Domini benediximus vobis de domo Domini
PS|117|27|Deus Dominus et inluxit nobis constituite diem sollemnem in condensis usque ad cornua altaris
PS|117|28|Deus meus es tu et confitebor tibi Deus meus % es tu; et exaltabo te confitebor tibi quoniam exaudisti me et factus es mihi in salutem
PS|117|29|confitemini Domino quoniam bonus quoniam in saeculum misericordia eius
PS|118|1|alleluia aleph beati inmaculati in via qui ambulant in lege Domini
PS|118|2|beati qui scrutantur testimonia eius in toto corde exquirent eum
PS|118|3|non enim qui operantur iniquitatem in viis eius ambulaverunt
PS|118|4|tu mandasti mandata tua custodire nimis
PS|118|5|utinam dirigantur viae meae ad custodiendas iustificationes tuas
PS|118|6|tunc non confundar cum perspexero in omnibus mandatis tuis
PS|118|7|confitebor tibi in directione cordis in eo quod didici iudicia iustitiae tuae
PS|118|8|iustificationes tuas custodiam non me derelinquas usquequaque
PS|118|9|beth in quo corriget adulescentior viam suam in custodiendo sermones tuos
PS|118|10|in toto corde meo exquisivi te non repellas me a mandatis tuis
PS|118|11|in corde meo abscondi eloquia tua ut non peccem tibi
PS|118|12|benedictus es Domine doce me iustificationes tuas
PS|118|13|in labiis meis pronuntiavi omnia iudicia oris tui
PS|118|14|in via testimoniorum tuorum delectatus sum sicut in omnibus divitiis
PS|118|15|in mandatis tuis exercebor et considerabo vias tuas
PS|118|16|in iustificationibus tuis meditabor non obliviscar sermones tuos
PS|118|17|gimel retribue servo tuo vivifica me et custodiam sermones tuos
PS|118|18|revela oculos meos et considerabo mirabilia de lege tua
PS|118|19|incola ego sum in terra non abscondas a me mandata tua
PS|118|20|concupivit anima mea desiderare iustificationes tuas in omni tempore
PS|118|21|increpasti superbos maledicti qui declinant a mandatis tuis
PS|118|22|aufer a me obprobrium et contemptum quia testimonia tua exquisivi
PS|118|23|etenim sederunt principes et adversum me loquebantur servus autem tuus exercebatur in iustificationibus tuis
PS|118|24|nam et testimonia tua meditatio mea et consilium meum iustificationes tuae
PS|118|25|deleth adhesit pavimento anima mea vivifica me secundum verbum tuum
PS|118|26|vias meas enuntiavi et exaudisti me doce me iustificationes tuas
PS|118|27|viam iustificationum tuarum instrue me et exercebor in mirabilibus tuis
PS|118|28|dormitavit anima mea prae taedio confirma me in verbis tuis
PS|118|29|viam iniquitatis amove a me et lege tua miserere mei
PS|118|30|viam veritatis elegi iudicia tua non sum oblitus
PS|118|31|adhesi testimoniis tuis Domine noli me confundere
PS|118|32|viam mandatorum tuorum cucurri cum dilatasti cor meum
PS|118|33|he legem pone mihi Domine viam iustificationum tuarum et exquiram eam semper
PS|118|34|da mihi intellectum et scrutabor legem tuam et custodiam illam in toto corde meo
PS|118|35|deduc me in semita mandatorum tuorum quia ipsam volui
PS|118|36|inclina cor meum in testimonia tua et non in avaritiam
PS|118|37|averte oculos meos ne videant vanitatem in via tua vivifica me
PS|118|38|statue servo tuo eloquium tuum in timore tuo
PS|118|39|amputa obprobrium meum quod suspicatus sum quia iudicia tua iucunda
PS|118|40|ecce concupivi mandata tua in aequitate tua vivifica me
PS|118|41|vav et veniat super me misericordia tua Domine salutare tuum secundum eloquium tuum
PS|118|42|et respondebo exprobrantibus mihi verbum quia speravi in sermonibus tuis
PS|118|43|et ne auferas de ore meo verbum veritatis usquequaque quia in iudiciis tuis supersperavi
PS|118|44|et custodiam legem tuam semper in saeculum et in saeculum saeculi
PS|118|45|et ambulabam in latitudine quia mandata tua exquisivi
PS|118|46|et loquebar in testimoniis tuis in conspectu regum et non confundebar
PS|118|47|et meditabar in mandatis tuis quae dilexi
PS|118|48|et levavi manus meas ad mandata quae dilexi et exercebar in iustificationibus tuis
PS|118|49|zai memor esto verbi tui servo tuo in quo mihi spem dedisti
PS|118|50|haec me consolata est in humilitate mea quia eloquium tuum vivificavit me
PS|118|51|superbi inique agebant usquequaque a lege autem tua non declinavi
PS|118|52|memor fui iudiciorum tuorum a saeculo Domine et consolatus sum
PS|118|53|defectio tenuit me prae peccatoribus derelinquentibus legem tuam
PS|118|54|cantabiles mihi erant iustificationes tuae in loco peregrinationis meae
PS|118|55|memor fui in nocte nominis tui Domine et custodivi legem tuam
PS|118|56|haec facta est mihi quia iustificationes tuas exquisivi
PS|118|57|heth portio mea Dominus dixi custodire legem tuam
PS|118|58|deprecatus sum faciem tuam in toto corde meo miserere mei secundum eloquium tuum
PS|118|59|cogitavi vias meas et avertisti pedes meos in testimonia tua
PS|118|60|paratus sum et non sum turbatus ut custodiam mandata tua
PS|118|61|funes peccatorum circumplexi sunt me et legem tuam non sum oblitus
PS|118|62|media nocte surgebam ad confitendum tibi super iudicia iustificationis tuae
PS|118|63|particeps ego sum omnium timentium te et custodientium mandata tua
PS|118|64|misericordia Domini plena est terra iustificationes tuas doce me
PS|118|65|teth bonitatem fecisti cum servo tuo Domine secundum verbum tuum
PS|118|66|bonitatem et disciplinam et scientiam doce me quia mandatis tuis credidi
PS|118|67|priusquam humiliarer ego deliqui propterea eloquium tuum custodivi
PS|118|68|bonus es tu et in bonitate tua doce me iustificationes tuas
PS|118|69|multiplicata est super me iniquitas superborum ego autem in toto corde scrutabor mandata tua
PS|118|70|coagulatum est sicut lac cor eorum ego vero legem tuam meditatus sum
PS|118|71|bonum mihi quia humiliasti me ut discam iustificationes tuas
PS|118|72|bonum mihi lex oris tui super milia auri et argenti
PS|118|73|ioth manus tuae fecerunt me et plasmaverunt me da mihi intellectum et discam mandata tua
PS|118|74|qui timent te videbunt me et laetabuntur quia in verba tua supersperavi
PS|118|75|cognovi Domine quia aequitas iudicia tua et veritate humiliasti me
PS|118|76|fiat misericordia tua ut consoletur me secundum eloquium tuum servo tuo
PS|118|77|veniant mihi miserationes tuae et vivam quia lex tua meditatio mea est
PS|118|78|confundantur superbi quia iniuste iniquitatem fecerunt in me ego autem exercebor in mandatis tuis
PS|118|79|convertantur mihi timentes te et qui noverunt testimonia tua
PS|118|80|fiat cor meum inmaculatum in iustificationibus tuis ut non confundar
PS|118|81|caf defecit in salutare tuum anima mea in verbum tuum supersperavi
PS|118|82|defecerunt oculi mei in eloquium tuum dicentes quando consolaberis me
PS|118|83|quia factus sum sicut uter in pruina iustificationes tuas non sum oblitus
PS|118|84|quot sunt dies servo tuo quando facies de persequentibus me iudicium
PS|118|85|narraverunt mihi iniqui fabulationes sed non ut lex tua
PS|118|86|omnia mandata tua veritas inique persecuti sunt me adiuva me
PS|118|87|paulo minus consummaverunt me in terra ego autem non dereliqui mandata tua
PS|118|88|secundum misericordiam tuam vivifica me et custodiam testimonia oris tui
PS|118|89|lamed in aeternum Domine verbum tuum permanet in caelo
PS|118|90|in generationem et generationem veritas tua fundasti terram et permanet
PS|118|91|ordinatione tua perseverat dies quoniam omnia serviunt tibi
PS|118|92|nisi quod lex tua meditatio mea est tunc forte perissem in humilitate mea
PS|118|93|in aeternum non obliviscar iustificationes tuas quia in ipsis vivificasti me
PS|118|94|tuus sum ego salvum me fac quoniam iustificationes tuas exquisivi
PS|118|95|me expectaverunt peccatores ut perderent me testimonia tua intellexi
PS|118|96|omni consummationi vidi finem latum mandatum tuum nimis
PS|118|97|mem quomodo dilexi legem tuam tota die meditatio mea est
PS|118|98|super inimicos meos prudentem me fecisti mandato tuo quia in aeternum mihi est
PS|118|99|super omnes docentes me intellexi quia testimonia tua meditatio mea est
PS|118|100|super senes intellexi quia mandata tua quaesivi
PS|118|101|ab omni via mala prohibui pedes meos ut custodiam verba tua
PS|118|102|a iudiciis tuis non declinavi quia tu legem posuisti mihi
PS|118|103|quam dulcia faucibus meis eloquia tua super mel ori meo
PS|118|104|a mandatis tuis intellexi propterea odivi omnem viam iniquitatis
PS|118|105|nun lucerna pedibus meis verbum tuum et lumen semitis meis
PS|118|106|iuravi et statui custodire iudicia iustitiae tuae
PS|118|107|humiliatus sum usquequaque Domine vivifica me secundum verbum tuum
PS|118|108|voluntaria oris mei beneplacita fac Domine et iudicia tua doce me
PS|118|109|anima mea in manibus meis semper et legem tuam non sum oblitus
PS|118|110|posuerunt peccatores laqueum mihi et de mandatis tuis non erravi
PS|118|111|hereditate adquisivi testimonia tua in aeternum quia exultatio cordis mei sunt
PS|118|112|inclinavi cor meum ad faciendas iustificationes tuas in aeternum propter retributionem
PS|118|113|samech iniquos odio habui et legem tuam dilexi
PS|118|114|adiutor meus et susceptor meus es tu in verbum tuum supersperavi
PS|118|115|declinate a me maligni et scrutabor mandata Dei mei
PS|118|116|suscipe me secundum eloquium tuum et vivam et non confundas me ab expectatione mea
PS|118|117|adiuva me et salvus ero et meditabor in iustificationibus tuis semper
PS|118|118|sprevisti omnes discedentes a iustitiis tuis quia iniusta cogitatio eorum
PS|118|119|praevaricantes reputavi omnes peccatores terrae ideo dilexi testimonia tua
PS|118|120|confige timore tuo carnes meas a iudiciis %enim; tuis timui
PS|118|121|ain feci iudicium et iustitiam non tradas me calumniantibus me
PS|118|122|suscipe servum tuum in bonum non calumnientur me superbi
PS|118|123|oculi mei defecerunt in salutare tuum et in eloquium iustitiae tuae
PS|118|124|fac cum servo tuo secundum misericordiam tuam et iustificationes tuas doce me
PS|118|125|servus tuus sum ego da mihi intellectum et sciam testimonia tua
PS|118|126|tempus faciendi Domino dissipaverunt legem tuam
PS|118|127|ideo dilexi mandata tua super aurum et topazion
PS|118|128|propterea ad omnia mandata tua dirigebar omnem viam iniquam odio habui
PS|118|129|fe mirabilia testimonia tua ideo scrutata est ea anima mea
PS|118|130|declaratio sermonum tuorum inluminat et intellectum dat parvulis
PS|118|131|os meum aperui et adtraxi spiritum quia mandata tua desiderabam
PS|118|132|aspice in me et miserere mei secundum iudicium diligentium nomen tuum
PS|118|133|gressus meos dirige secundum eloquium tuum et non dominetur mei omnis iniustitia
PS|118|134|redime me a calumniis hominum et custodiam mandata tua
PS|118|135|faciem tuam inlumina super servum tuum et doce me iustificationes tuas
PS|118|136|exitus aquarum deduxerunt oculi mei quia non custodierunt legem tuam
PS|118|137|sade iustus es Domine et rectum iudicium tuum
PS|118|138|mandasti iustitiam testimonia tua et veritatem tuam nimis
PS|118|139|tabescere me fecit zelus meus quia obliti sunt verba tua inimici mei
PS|118|140|ignitum eloquium tuum vehementer et servus tuus dilexit illud
PS|118|141|adulescentulus sum ego et contemptus iustificationes tuas non sum oblitus
PS|118|142|iustitia tua iustitia in aeternum et lex tua veritas
PS|118|143|tribulatio et angustia invenerunt me mandata tua meditatio mea
PS|118|144|aequitas testimonia tua in aeternum intellectum da mihi et vivam
PS|118|145|cof clamavi in toto corde exaudi me Domine iustificationes tuas requiram
PS|118|146|clamavi te salvum me fac et custodiam mandata tua
PS|118|147|praeveni in maturitate et clamavi in verba tua supersperavi
PS|118|148|praevenerunt oculi mei ad diluculum ut meditarer eloquia tua
PS|118|149|vocem meam audi secundum misericordiam tuam Domine secundum iudicium tuum vivifica me
PS|118|150|adpropinquaverunt persequentes me iniquitate a lege autem tua longe facti sunt
PS|118|151|prope es tu Domine et omnes viae tuae veritas
PS|118|152|initio cognovi de testimoniis tuis quia in aeternum fundasti ea
PS|118|153|res vide humilitatem meam et eripe me quia legem tuam non sum oblitus
PS|118|154|iudica iudicium meum et redime me propter eloquium tuum vivifica me
PS|118|155|longe a peccatoribus salus quia iustificationes tuas non exquisierunt
PS|118|156|misericordiae tuae multae Domine secundum iudicia tua vivifica me
PS|118|157|multi qui persequuntur me et tribulant me a testimoniis tuis non declinavi
PS|118|158|vidi praevaricantes et tabescebam quia eloquia tua non custodierunt
PS|118|159|vide quoniam mandata tua dilexi Domine in misericordia tua vivifica me
PS|118|160|principium verborum tuorum veritas et in aeternum omnia iudicia iustitiae tuae
PS|118|161|sen principes persecuti sunt me gratis et a verbis tuis formidavit cor meum
PS|118|162|laetabor ego super eloquia tua sicut qui invenit spolia multa
PS|118|163|iniquitatem odio habui et abominatus sum legem autem tuam dilexi
PS|118|164|septies in die laudem dixi tibi super iudicia iustitiae tuae
PS|118|165|pax multa diligentibus legem tuam et non est illis scandalum
PS|118|166|expectabam salutare tuum Domine et mandata tua dilexi
PS|118|167|custodivit anima mea testimonia tua et dilexi ea vehementer
PS|118|168|servavi mandata tua et testimonia tua quia omnes viae meae in conspectu tuo
PS|118|169|thau adpropinquet deprecatio mea in conspectu tuo Domine iuxta eloquium tuum da mihi intellectum
PS|118|170|intret postulatio mea in conspectu tuo secundum eloquium tuum eripe me
PS|118|171|eructabunt labia mea hymnum cum docueris me iustificationes tuas
PS|118|172|pronuntiabit lingua mea eloquium tuum quia omnia mandata tua aequitas
PS|118|173|fiat manus tua ut salvet me quoniam mandata tua elegi
PS|118|174|concupivi salutare tuum Domine et lex tua meditatio mea
PS|118|175|vivet anima mea et laudabit te et iudicia tua adiuvabunt me
PS|118|176|erravi sicut ovis quae periit quaere servum tuum quia mandata tua non sum oblitus
PS|119|1|canticum graduum ad Dominum cum tribularer clamavi et exaudivit me
PS|119|2|Domine libera animam meam a labiis iniquis a lingua dolosa
PS|119|3|quid detur tibi et quid adponatur tibi ad linguam dolosam
PS|119|4|sagittae potentis acutae cum carbonibus desolatoriis
PS|119|5|heu mihi quia incolatus meus prolongatus est habitavi cum habitationibus Cedar
PS|119|6|multum incola fuit anima mea
PS|119|7|cum his qui oderant pacem eram pacificus cum loquebar illis inpugnabant me gratis
PS|120|1|canticum graduum levavi oculos meos in montes unde veniet auxilium mihi
PS|120|2|auxilium meum a Domino qui fecit caelum et terram
PS|120|3|non det in commotionem pedem tuum neque dormitet qui custodit te
PS|120|4|ecce non dormitabit neque dormiet qui custodit Israhel
PS|120|5|Dominus custodit te Dominus protectio tua super manum dexteram tuam
PS|120|6|per diem sol non uret te neque luna per noctem
PS|120|7|Dominus custodit te ab omni malo custodiat animam tuam Dominus
PS|120|8|Dominus custodiat introitum tuum et exitum tuum ex hoc nunc et usque in saeculum
PS|121|1|canticum graduum huic David laetatus sum in his quae dicta sunt mihi in domum Domini ibimus
PS|121|2|stantes erant pedes nostri in atriis tuis Hierusalem
PS|121|3|Hierusalem quae aedificatur ut civitas cuius participatio eius in id ipsum
PS|121|4|illic enim ascenderunt tribus tribus Domini testimonium Israhel ad confitendum nomini Domini
PS|121|5|quia illic sederunt sedes in iudicium sedes super domum David
PS|121|6|rogate quae ad pacem sunt Hierusalem et abundantia diligentibus te
PS|121|7|fiat pax in virtute tua et abundantia in turribus tuis
PS|121|8|propter fratres meos et proximos meos loquebar pacem de te
PS|121|9|propter domum Domini Dei nostri quaesivi bona tibi
PS|122|1|canticum graduum ad te levavi oculos meos qui habitas in caelo
PS|122|2|ecce sicut oculi servorum in manibus dominorum suorum sicut oculi ancillae in manibus dominae eius ita oculi nostri ad Dominum Deum nostrum donec misereatur nostri
PS|122|3|miserere nostri Domine miserere nostri quia multum repleti sumus despectione
PS|122|4|quia multum repleta est anima nostra obprobrium abundantibus et despectio superbis
PS|123|1|canticum graduum huic David nisi quia Dominus erat in nobis dicat nunc Israhel
PS|123|2|nisi quia Dominus erat in nobis cum exsurgerent in nos homines
PS|123|3|forte vivos degluttissent nos cum irasceretur furor eorum in nos
PS|123|4|forsitan aqua absorbuisset nos
PS|123|5|torrentem pertransivit anima nostra forsitan pertransisset anima nostra aquam intolerabilem
PS|123|6|benedictus Dominus qui non dedit nos in captionem dentibus eorum
PS|123|7|anima nostra sicut passer erepta est de laqueo venantium laqueus contritus est et nos liberati sumus
PS|123|8|adiutorium nostrum in nomine Domini qui fecit caelum et terram
PS|124|1|canticum graduum qui confidunt in Domino sicut mons Sion non commovebitur in aeternum qui habitat
PS|124|2|in Hierusalem montes in circuitu eius et Dominus in circuitu populi sui ex hoc nunc et usque in saeculum
PS|124|3|quia non relinquet virgam peccatorum super sortem iustorum ut non extendant iusti ad iniquitatem manus suas
PS|124|4|benefac Domine bonis et rectis corde
PS|124|5|declinantes autem in obligationes adducet Dominus cum operantibus iniquitatem pax super Israhel
PS|125|1|canticum graduum in convertendo Dominum captivitatem Sion facti sumus sicut consolati
PS|125|2|tunc repletum est gaudio os nostrum et lingua nostra exultatione tunc dicent inter gentes magnificavit Dominus facere cum eis
PS|125|3|magnificavit Dominus facere nobiscum facti sumus laetantes
PS|125|4|converte Domine captivitatem nostram sicut torrens in austro
PS|125|5|qui seminant in lacrimis in exultatione metent
PS|125|6|euntes ibant et flebant portantes semina sua venientes autem venient in exultatione portantes manipulos suos
PS|126|1|canticum graduum Salomonis nisi Dominus aedificaverit domum in vanum laboraverunt qui aedificant eam nisi Dominus custodierit civitatem frustra vigilavit qui custodit
PS|126|2|vanum est vobis ante lucem surgere surgere postquam sederitis qui manducatis panem doloris cum dederit dilectis suis somnum
PS|126|3|ecce hereditas Domini filii mercis fructus ventris
PS|126|4|sicut sagittae in manu potentis ita filii excussorum
PS|126|5|beatus vir qui implebit desiderium suum ex ipsis non confundentur cum loquentur inimicis suis in porta
PS|127|1|canticum graduum beati omnes qui timent Dominum qui ambulant in viis eius
PS|127|2|labores manuum tuarum quia; manducabis beatus es et bene tibi erit
PS|127|3|uxor tua sicut vitis abundans in lateribus domus tuae filii tui sicut novella olivarum in circuitu mensae tuae
PS|127|4|ecce sic benedicetur homo qui timet Dominum
PS|127|5|benedicat te Dominus ex Sion et videas bona Hierusalem omnibus diebus vitae tuae
PS|127|6|et videas filios filiorum tuorum pax super Israhel
PS|128|1|canticum graduum saepe expugnaverunt me a iuventute mea dicat nunc Israhel
PS|128|2|saepe expugnaverunt me a iuventute mea etenim non potuerunt mihi
PS|128|3|supra dorsum meum fabricabantur peccatores prolongaverunt iniquitatem suam
PS|128|4|Dominus iustus concidet cervices peccatorum
PS|128|5|confundantur et convertantur retrorsum omnes qui oderunt Sion
PS|128|6|fiant sicut faenum tectorum quod priusquam evellatur exaruit
PS|128|7|de quo non implevit manum suam qui metit et sinum suum qui manipulos colligit
PS|128|8|et non dixerunt qui praeteribant benedictio Domini super vos benediximus vobis in nomine Domini
PS|129|1|canticum graduum de profundis clamavi ad te Domine
PS|129|2|Domine exaudi vocem meam fiant aures tuae intendentes in vocem deprecationis meae
PS|129|3|si iniquitates observabis Domine Domine quis sustinebit
PS|129|4|quia apud te propitiatio est propter legem tuam sustinui te Domine sustinuit anima mea in verbum eius
PS|129|5|speravit anima mea in Domino
PS|129|6|a custodia matutina usque ad noctem speret Israhel in Domino
PS|129|7|quia apud Dominum misericordia et copiosa apud eum redemptio
PS|129|8|et ipse redimet Israhel ex omnibus iniquitatibus eius
PS|130|1|canticum graduum David Domine non est exaltatum cor meum neque elati sunt oculi mei neque ambulavi in magnis neque in mirabilibus super me
PS|130|2|si non humiliter sentiebam sed exaltavi animam meam sicut ablactatum super matrem suam ita retributio in anima mea
PS|130|3|speret Israhel in Domino ex hoc nunc et usque in saeculum
PS|131|1|canticum graduum memento Domine David et omnis mansuetudinis eius
PS|131|2|sicut iuravit Domino votum vovit Deo Iacob
PS|131|3|si introiero in tabernaculum domus meae si ascendero in lectum strati mei
PS|131|4|si dedero somnum oculis meis et palpebris meis dormitationem
PS|131|5|et requiem temporibus meis donec inveniam locum Domino tabernaculum Deo Iacob
PS|131|6|ecce audivimus eam in Efrata invenimus eam in campis silvae
PS|131|7|introibimus in tabernacula eius adorabimus in loco ubi steterunt pedes eius
PS|131|8|surge Domine in requiem tuam tu et arca sanctificationis tuae
PS|131|9|sacerdotes tui induentur iustitia et sancti tui exultabunt
PS|131|10|propter David servum tuum non avertas faciem christi tui
PS|131|11|iuravit Dominus David veritatem et non frustrabit eum de fructu ventris tui ponam super sedem tuam
PS|131|12|si custodierint filii tui testamentum meum et testimonia mea haec quae docebo eos et filii eorum usque in saeculum sedebunt super sedem tuam
PS|131|13|quoniam elegit Dominus Sion elegit eam in habitationem sibi
PS|131|14|haec requies mea in saeculum saeculi hic habitabo quoniam elegi eam
PS|131|15|viduam eius benedicens benedicam pauperes eius saturabo panibus
PS|131|16|sacerdotes eius induam salutari et sancti eius exultatione exultabunt
PS|131|17|illic producam cornu David paravi lucernam christo meo
PS|131|18|inimicos eius induam confusione super ipsum autem efflorebit sanctificatio mea
PS|132|1|canticum graduum David ecce quam bonum et quam iucundum habitare fratres in unum
PS|132|2|sicut unguentum in capite quod descendit in barbam barbam Aaron quod descendit in ora vestimenti eius
PS|132|3|sicut ros Hermon qui descendit in montes Sion quoniam illic mandavit Dominus benedictionem et vitam usque in saeculum
PS|133|1|canticum graduum ecce nunc benedicite Dominum omnes servi Domini qui statis in domo Domini %in atriis domus Dei nostri;
PS|133|2|in noctibus extollite manus vestras in sancta et benedicite Domino
PS|133|3|benedicat te Dominus ex Sion qui fecit caelum et terram
PS|134|1|alleluia laudate nomen Domini laudate servi Dominum
PS|134|2|qui statis in domo Domini in atriis domus Dei nostri
PS|134|3|laudate Dominum quia bonus Dominus psallite nomini eius quoniam suave
PS|134|4|quoniam Iacob elegit sibi Dominus Israhel in possessionem sibi
PS|134|5|quia ego cognovi quod magnus est Dominus et Deus noster prae omnibus diis
PS|134|6|omnia quae voluit Dominus fecit in caelo et in terra in mare et in omnibus abyssis
PS|134|7|educens nubes ab extremo terrae fulgora in pluviam fecit qui producit ventos de thesauris suis
PS|134|8|qui percussit primogenita Aegypti ab homine usque ad pecus
PS|134|9|emisit signa et prodigia in medio tui Aegypte in Pharaonem et in omnes servos eius
PS|134|10|qui percussit gentes multas et occidit reges fortes
PS|134|11|Seon regem Amorreorum et Og regem Basan et omnia regna Chanaan
PS|134|12|et dedit terram eorum hereditatem hereditatem Israhel populo suo
PS|134|13|Domine nomen tuum in aeternum Domine memoriale tuum in generationem et generationem
PS|134|14|quia iudicabit Dominus populum suum et in servis suis deprecabitur
PS|134|15|simulacra gentium argentum et aurum opera manuum hominum
PS|134|16|os habent et non loquentur oculos habent et non videbunt
PS|134|17|aures habent et non audient neque enim est spiritus in ore eorum
PS|134|18|similes illis fiant qui faciunt ea et omnes qui sperant in eis
PS|134|19|domus Israhel benedicite Domino domus Aaron benedicite Domino
PS|134|20|domus Levi benedicite Domino qui timetis Dominum benedicite Domino
PS|134|21|benedictus Dominus ex Sion qui habitat in Hierusalem
PS|135|1|alleluia confitemini Domino quoniam bonus quoniam in aeternum misericordia eius
PS|135|2|confitemini Deo deorum quoniam in aeternum misericordia eius
PS|135|3|confitemini Domino dominorum quoniam in aeternum misericordia eius
PS|135|4|qui facit mirabilia magna solus quoniam in aeternum misericordia eius
PS|135|5|qui fecit caelos in intellectu quoniam in aeternum misericordia eius
PS|135|6|qui firmavit terram super aquas quoniam in aeternum misericordia eius
PS|135|7|qui fecit luminaria magna quoniam in aeternum misericordia eius
PS|135|8|solem in potestatem diei quoniam in aeternum misericordia eius
PS|135|9|lunam et stellas in potestatem noctis quoniam in aeternum misericordia eius
PS|135|10|qui percussit Aegyptum cum primogenitis eorum quoniam in aeternum misericordia eius
PS|135|11|qui eduxit Israhel de medio eorum quoniam in aeternum misericordia eius
PS|135|12|in manu potenti et brachio excelso quoniam in aeternum misericordia eius
PS|135|13|qui divisit Rubrum mare in divisiones quoniam in aeternum misericordia eius
PS|135|14|et duxit Israhel per medium eius quoniam in aeternum misericordia eius
PS|135|15|et excussit Pharaonem et virtutem eius in mari Rubro quoniam in aeternum misericordia eius
PS|135|16|qui transduxit populum suum in deserto quoniam in aeternum misericordia eius
PS|135|17|qui percussit reges magnos quoniam in aeternum misericordia eius
PS|135|18|et occidit reges fortes quoniam in aeternum misericordia eius
PS|135|19|Seon regem Amorreorum quoniam in aeternum misericordia eius
PS|135|20|et Og regem Basan quoniam in aeternum misericordia eius
PS|135|21|et dedit terram eorum hereditatem quoniam in aeternum misericordia eius
PS|135|22|hereditatem Israhel servo suo quoniam in aeternum misericordia eius
PS|135|23|quia in humilitate nostra memor fuit nostri quoniam in aeternum misericordia eius
PS|135|24|et redemit nos ab inimicis nostris quoniam in aeternum misericordia eius
PS|135|25|qui dat escam omni carni quoniam in aeternum misericordia eius
PS|135|26|confitemini Deo caeli quoniam in aeternum misericordia eius confitemini Domino dominorum quoniam in aeternum misericordia eius
PS|136|1|David Hieremiae super flumina Babylonis illic sedimus et flevimus cum recordaremur Sion
PS|136|2|in salicibus in medio eius suspendimus organa nostra
PS|136|3|quia illic interrogaverunt nos qui captivos duxerunt nos verba cantionum et qui abduxerunt nos hymnum cantate nobis de canticis Sion
PS|136|4|quomodo cantabimus canticum Domini in terra aliena
PS|136|5|si oblitus fuero tui Hierusalem oblivioni detur dextera mea
PS|136|6|adhereat lingua mea faucibus meis si non meminero tui si non praeposuero Hierusalem in principio laetitiae meae
PS|136|7|memor esto Domine filiorum Edom diem Hierusalem qui dicunt exinanite exinanite usque ad fundamentum in ea
PS|136|8|filia Babylonis misera beatus qui retribuet tibi retributionem tuam quam retribuisti nobis
PS|136|9|beatus qui tenebit et adlidet parvulos tuos ad petram
PS|137|1|ipsi David confitebor tibi Domine in toto corde meo quoniam audisti verba oris mei in conspectu angelorum psallam tibi
PS|137|2|adorabo ad templum sanctum tuum et confitebor nomini tuo super misericordia tua et veritate tua quoniam magnificasti super omne nomen sanctum tuum
PS|137|3|in quacumque die invocavero te exaudi me multiplicabis me in anima mea virtute
PS|137|4|confiteantur tibi Domine omnes reges terrae quia audierunt omnia verba oris tui
PS|137|5|et cantent in viis Domini quoniam magna gloria Domini
PS|137|6|quoniam excelsus Dominus et humilia respicit et alta a longe cognoscit
PS|137|7|si ambulavero in medio tribulationis vivificabis me super iram inimicorum meorum extendisti manum tuam et salvum me fecit dextera tua
PS|137|8|Dominus retribuet propter me Domine misericordia tua in saeculum opera manuum tuarum ne dispicias
PS|138|1|in finem David psalmus
PS|138|2|Domine probasti me et cognovisti me tu cognovisti sessionem meam et surrectionem meam
PS|138|3|intellexisti cogitationes meas de longe semitam meam et funiculum meum investigasti
PS|138|4|et omnes vias meas praevidisti quia non est sermo in lingua mea
PS|138|5|ecce Domine tu cognovisti omnia novissima et antiqua tu formasti me et posuisti super me manum tuam
PS|138|6|mirabilis facta est scientia tua ex me confortata est non potero ad eam
PS|138|7|quo ibo ab spiritu tuo et quo a facie tua fugiam
PS|138|8|si ascendero in caelum tu illic es si descendero ad infernum ades
PS|138|9|si sumpsero pinnas meas diluculo et habitavero in extremis maris
PS|138|10|etenim illuc manus tua deducet me et tenebit me dextera tua
PS|138|11|et dixi forsitan tenebrae conculcabunt me et nox inluminatio in deliciis meis
PS|138|12|quia tenebrae non obscurabuntur a te et nox sicut dies inluminabitur sicut tenebrae eius ita et lumen eius
PS|138|13|quia tu possedisti renes meos suscepisti me de utero matris meae
PS|138|14|confitebor tibi quia terribiliter magnificatus es mirabilia opera tua et anima mea cognoscit nimis
PS|138|15|non est occultatum os meum a te quod fecisti in occulto et substantia mea in inferioribus terrae
PS|138|16|inperfectum meum viderunt oculi tui et in libro tuo omnes scribentur die formabuntur et nemo in eis
PS|138|17|mihi autem nimis honorificati sunt amici tui Deus nimis confirmati sunt principatus eorum
PS|138|18|dinumerabo eos et super harenam multiplicabuntur exsurrexi et adhuc sum tecum
PS|138|19|si occideris Deus peccatores et viri sanguinum declinate a me
PS|138|20|quia dices in cogitatione accipient in vanitate civitates tuas
PS|138|21|nonne qui oderunt te Domine oderam et super inimicos tuos tabescebam
PS|138|22|perfecto odio oderam illos inimici facti sunt mihi
PS|138|23|proba me Deus et scito cor meum interroga me et cognosce semitas meas
PS|138|24|et vide si via iniquitatis in me est et deduc me in via aeterna
PS|139|1|in finem psalmus David
PS|139|2|eripe me Domine ab homine malo a viro iniquo eripe me
PS|139|3|qui cogitaverunt iniquitates in corde tota die constituebant proelia
PS|139|4|acuerunt linguam suam sicut serpentis venenum aspidum sub labiis eorum diapsalma
PS|139|5|custodi me Domine de manu peccatoris ab hominibus iniquis eripe me qui cogitaverunt subplantare gressus meos
PS|139|6|absconderunt superbi laqueum mihi et funes extenderunt in laqueum iuxta iter scandalum posuerunt mihi diapsalma
PS|139|7|dixi Domino Deus meus es tu exaudi Domine vocem deprecationis meae
PS|139|8|Domine Domine virtus salutis meae obumbrasti super caput meum in die belli
PS|139|9|non tradas Domine desiderio meo peccatori cogitaverunt contra me ne derelinquas me ne forte exaltentur diapsalma
PS|139|10|caput circuitus eorum labor labiorum ipsorum operiet eos
PS|139|11|cadent super eos carbones in igne deicies eos in miseriis non subsistent
PS|139|12|vir linguosus non dirigetur in terra virum iniustum mala capient in interitu
PS|139|13|cognovi quia faciet Dominus iudicium inopis et vindictam pauperum
PS|139|14|verumtamen iusti confitebuntur nomini tuo habitabunt recti cum vultu tuo
PS|140|1|psalmus David Domine clamavi ad te exaudi me intende voci meae cum clamavero ad te
PS|140|2|dirigatur oratio mea sicut incensum in conspectu tuo elevatio manuum mearum sacrificium vespertinum
PS|140|3|pone Domine custodiam ori meo et ostium circumstantiae labiis meis
PS|140|4|non declines cor meum in verba malitiae ad excusandas excusationes in peccatis cum hominibus operantibus iniquitatem et non communicabo cum electis eorum
PS|140|5|corripiet me iustus in misericordia et increpabit me oleum %autem; peccatoris non inpinguet caput meum quoniam adhuc et oratio mea in beneplacitis eorum
PS|140|6|absorti sunt iuncti petrae iudices eorum audient verba mea quoniam potuerunt
PS|140|7|sicut crassitudo terrae erupta est super terram dissipata sunt ossa nostra secus infernum
PS|140|8|quia ad te Domine Domine oculi mei in te speravi non auferas animam meam
PS|140|9|custodi me a laqueo quem statuerunt mihi et ab scandalis operantium iniquitatem
PS|140|10|cadent in retiaculo eius peccatores singulariter sum ego donec transeam
PS|141|1|intellectus David cum esset in spelunca oratio
PS|141|2|voce mea ad Dominum clamavi voce mea ad Dominum deprecatus sum
PS|141|3|effundo in conspectu eius deprecationem meam tribulationem meam ante ipsum pronuntio
PS|141|4|in deficiendo ex me spiritum meum et tu cognovisti semitas meas in via hac qua ambulabam absconderunt laqueum mihi
PS|141|5|considerabam ad dexteram et videbam et non erat qui cognosceret me periit fuga a me et non est qui requirit animam meam
PS|141|6|clamavi ad te Domine dixi tu es spes mea portio mea in terra viventium
PS|141|7|intende ad deprecationem meam quia humiliatus sum nimis libera me a persequentibus me quia confortati sunt super me
PS|141|8|educ de custodia animam meam ad confitendum nomini tuo me expectant iusti donec retribuas mihi
PS|142|1|psalmus David quando filius eum persequebatur Domine exaudi orationem meam auribus percipe obsecrationem meam in veritate tua exaudi me in tua iustitia
PS|142|2|et non intres in iudicio cum servo tuo quia non iustificabitur in conspectu tuo omnis vivens
PS|142|3|quia persecutus est inimicus animam meam humiliavit in terra vitam meam conlocavit me in obscuris sicut mortuos saeculi
PS|142|4|et anxiatus est super me spiritus meus in me turbatum est cor meum
PS|142|5|memor fui dierum antiquorum meditatus sum in omnibus operibus tuis in factis manuum tuarum meditabar
PS|142|6|expandi manus meas ad te anima mea sicut terra sine aqua tibi diapsalma
PS|142|7|velociter exaudi me Domine defecit spiritus meus non avertas faciem tuam a me et similis ero descendentibus in lacum
PS|142|8|auditam mihi fac mane misericordiam tuam quia in te speravi notam fac mihi viam in qua ambulem quia ad te levavi animam meam
PS|142|9|eripe me de inimicis meis Domine ad te confugi
PS|142|10|doce me facere voluntatem tuam quia Deus meus es tu spiritus tuus bonus deducet me in terra recta
PS|142|11|propter nomen tuum Domine vivificabis me in aequitate tua educes de tribulatione animam meam
PS|142|12|et in misericordia tua disperdes inimicos meos et perdes omnes qui tribulant animam meam quoniam ego servus tuus sum
PS|143|1|David adversus Goliad benedictus Dominus Deus meus qui docet manus meas ad proelium digitos meos ad bellum
PS|143|2|misericordia mea et refugium meum susceptor meus et liberator meus protector meus et in eo speravi qui subdis populum meum sub me
PS|143|3|Domine quid est homo quia innotuisti ei aut filius hominis quia reputas eum
PS|143|4|homo vanitati similis factus est dies eius sicut umbra praetereunt
PS|143|5|Domine inclina caelos tuos et descende tange montes et fumigabunt
PS|143|6|fulgora coruscationem et dissipabis eos emitte sagittas tuas et conturbabis eos
PS|143|7|emitte manum tuam de alto eripe me et libera me de aquis multis de manu filiorum alienorum
PS|143|8|quorum os locutum est vanitatem et dextera eorum dextera iniquitatis
PS|143|9|Deus canticum novum cantabo tibi in psalterio decacordo psallam tibi
PS|143|10|qui das salutem regibus qui redimit David servum suum de gladio maligno
PS|143|11|eripe me et eripe me de manu filiorum alienigenarum quorum os locutum est vanitatem et dextera eorum dextera iniquitatis
PS|143|12|quorum filii sicut novella plantationis in iuventute sua filiae eorum conpositae circumornatae ut similitudo templi
PS|143|13|promptuaria eorum plena eructantia ex hoc in illud oves eorum fetosae abundantes in egressibus suis
PS|143|14|boves eorum crassi non est ruina maceriae neque transitus neque clamor in plateis eorum
PS|143|15|beatum dixerunt populum cui haec sunt beatus populus cuius Dominus Deus eius
PS|144|1|laudatio David exaltabo te Deus meus rex et benedicam nomini tuo in saeculum et in saeculum saeculi
PS|144|2|per singulos dies benedicam tibi et laudabo nomen tuum in saeculum et in saeculum saeculi
PS|144|3|magnus Dominus et laudabilis nimis et magnitudinis eius non est finis
PS|144|4|generatio et generatio laudabit opera tua et potentiam tuam pronuntiabunt
PS|144|5|magnificentiam gloriae sanctitatis tuae loquentur et mirabilia tua narrabunt
PS|144|6|et virtutem terribilium tuorum dicent et magnitudinem tuam narrabunt
PS|144|7|memoriam abundantiae suavitatis tuae eructabunt et iustitia tua exultabunt
PS|144|8|miserator et misericors Dominus patiens et multum misericors
PS|144|9|suavis Dominus universis et miserationes eius super omnia opera eius
PS|144|10|confiteantur tibi Domine omnia opera tua et sancti tui confiteantur tibi
PS|144|11|gloriam regni tui dicent et potentiam tuam loquentur
PS|144|12|ut notam faciant filiis hominum potentiam tuam et gloriam magnificentiae regni tui
PS|144|13|regnum tuum regnum omnium saeculorum et dominatio tua in omni generatione et progenie fidelis Dominus in omnibus verbis suis et sanctus in omnibus operibus suis
PS|144|14|adlevat Dominus omnes qui corruunt et erigit omnes elisos
PS|144|15|oculi omnium in te sperant et tu das escam illorum in tempore oportuno
PS|144|16|aperis tu manum tuam et imples omne animal benedictione
PS|144|17|iustus Dominus in omnibus viis suis et sanctus in omnibus operibus suis
PS|144|18|prope est Dominus omnibus invocantibus eum omnibus invocantibus eum in veritate
PS|144|19|voluntatem timentium se faciet et deprecationem eorum exaudiet et salvos faciet eos
PS|144|20|custodit Dominus omnes diligentes se et omnes peccatores disperdet
PS|144|21|laudationem Domini loquetur os meum et benedicat omnis caro nomini sancto eius in saeculum et in saeculum saeculi
PS|145|1|alleluia Aggei et Zacchariae
PS|145|2|lauda anima mea Dominum laudabo Dominum in vita mea psallam Deo meo quamdiu fuero nolite confidere in principibus
PS|145|3|in filiis hominum quibus non est salus
PS|145|4|exibit spiritus eius et revertetur in terram suam in illa die peribunt omnes cogitationes eorum
PS|145|5|beatus cuius Deus Iacob adiutor eius spes eius in Domino Deo ipsius
PS|145|6|qui fecit caelum et terram mare et omnia quae in eis
PS|145|7|qui custodit veritatem in saeculum facit iudicium iniuriam patientibus dat escam esurientibus Dominus solvit conpeditos
PS|145|8|Dominus inluminat caecos Dominus erigit adlisos Dominus diligit iustos
PS|145|9|Dominus custodit advenas pupillum et viduam suscipiet et viam peccatorum disperdet
PS|145|10|regnabit Dominus in saecula Deus tuus Sion in generationem et generationem
PS|146|1|alleluia Aggei et Zacchariae laudate Dominum quoniam bonum psalmus Deo nostro sit iucunda decoraque; laudatio
PS|146|2|aedificans Hierusalem Dominus dispersiones Israhel congregabit
PS|146|3|qui sanat contritos corde et alligat contritiones illorum
PS|146|4|qui numerat multitudinem stellarum et omnibus eis nomina vocans
PS|146|5|magnus Dominus noster et magna virtus eius et sapientiae eius non est numerus
PS|146|6|suscipiens mansuetos Dominus humilians autem peccatores usque ad terram
PS|146|7|praecinite Domino in confessione psallite Deo nostro in cithara
PS|146|8|qui operit caelum nubibus et parat terrae pluviam qui producit in montibus faenum et herbam servituti hominum
PS|146|9|et dat iumentis escam ipsorum et pullis corvorum invocantibus eum
PS|146|10|non in fortitudine equi voluntatem habebit nec in tibiis viri beneplacitum erit ei
PS|146|11|beneplacitum est Domino super timentes eum et in eis qui sperant super misericordia eius
PS|147|1|alleluia lauda Hierusalem Dominum lauda Deum tuum Sion
PS|147|2|quoniam confortavit seras portarum tuarum benedixit filiis tuis in te
PS|147|3|qui posuit fines tuos pacem et adipe frumenti satiat te
PS|147|4|qui emittit eloquium suum terrae velociter currit sermo eius
PS|147|5|qui dat nivem sicut lanam nebulam sicut cinerem spargit
PS|147|6|mittit cristallum suum sicut buccellas ante faciem frigoris eius quis sustinebit
PS|147|7|emittet verbum suum et liquefaciet ea flabit spiritus eius et fluent aquae
PS|147|8|qui adnuntiat verbum suum Iacob iustitias et iudicia sua Israhel
PS|147|9|non fecit taliter omni nationi et iudicia sua non manifestavit eis
PS|148|1|alleluia laudate Dominum de caelis laudate eum in excelsis
PS|148|2|laudate eum omnes angeli eius laudate eum omnes virtutes eius
PS|148|3|laudate eum sol et luna laudate eum omnes stellae et lumen
PS|148|4|laudate eum caeli caelorum et aqua quae super caelum est
PS|148|5|laudent nomen Domini quia ipse dixit et facta sunt ipse mandavit et creata sunt
PS|148|6|statuit ea in saeculum et in saeculum saeculi praeceptum posuit et non praeteribit
PS|148|7|laudate Dominum de terra dracones et omnes abyssi
PS|148|8|ignis grando nix glacies spiritus procellarum quae faciunt verbum eius
PS|148|9|montes et omnes colles ligna fructifera et omnes cedri
PS|148|10|bestiae et universa pecora serpentes et volucres pinnatae
PS|148|11|reges terrae et omnes populi principes et omnes iudices terrae
PS|148|12|iuvenes et virgines senes cum iunioribus laudent nomen Domini
PS|148|13|quia exaltatum est nomen eius solius
PS|148|14|confessio eius super caelum et terram et exaltabit cornu populi sui hymnus omnibus sanctis eius filiis Israhel populo adpropinquanti sibi
PS|149|1|alleluia cantate Domino canticum novum laus eius in ecclesia sanctorum
PS|149|2|laetetur Israhel in eo qui fecit eum et filii Sion exultent in rege suo
PS|149|3|laudent nomen eius in choro in tympano et psalterio psallant ei
PS|149|4|quia beneplacitum est Domino in populo suo et exaltabit mansuetos in salute
PS|149|5|exultabunt sancti in gloria laetabuntur in cubilibus suis
PS|149|6|exaltationes Dei in gutture eorum et gladii ancipites in manibus eorum
PS|149|7|ad faciendam vindictam in nationibus increpationes in populis
PS|149|8|ad alligandos reges eorum in conpedibus et nobiles eorum in manicis ferreis
PS|149|9|ut faciant in eis iudicium conscriptum gloria haec est omnibus sanctis eius
PS|150|1|alleluia laudate Dominum in sanctis eius laudate eum in firmamento virtutis eius
PS|150|2|laudate eum in virtutibus eius laudate eum secundum multitudinem magnitudinis eius
PS|150|3|laudate eum in sono tubae laudate eum in psalterio et cithara
PS|150|4|laudate eum in tympano et choro laudate eum in cordis et organo
PS|150|5|laudate eum in cymbalis bene sonantibus laudate eum in cymbalis iubilationis
PS|150|6|omnis spiritus laudet Dominum
PROV|1|1|parabolae Salomonis filii David regis Israhel
PROV|1|2|ad sciendam sapientiam et disciplinam
PROV|1|3|ad intellegenda verba prudentiae et suscipiendam eruditionem doctrinae iustitiam et iudicium et aequitatem
PROV|1|4|ut detur parvulis astutia adulescenti scientia et intellectus
PROV|1|5|audiens sapiens sapientior erit et intellegens gubernacula possidebit
PROV|1|6|animadvertet parabolam et interpretationem verba sapientium et enigmata eorum
PROV|1|7|timor Domini principium scientiae sapientiam atque doctrinam stulti despiciunt
PROV|1|8|audi fili mi disciplinam patris tui et ne dimittas legem matris tuae
PROV|1|9|ut addatur gratia capiti tuo et torques collo tuo
PROV|1|10|fili mi si te lactaverint peccatores ne adquiescas
PROV|1|11|si dixerint veni nobiscum insidiemur sanguini abscondamus tendiculas contra insontem frustra
PROV|1|12|degluttiamus eum sicut infernus viventem et integrum quasi descendentem in lacum
PROV|1|13|omnem pretiosam substantiam repperiemus implebimus domos nostras spoliis
PROV|1|14|sortem mitte nobiscum marsuppium unum sit omnium nostrum
PROV|1|15|fili mi ne ambules cum eis prohibe pedem tuum a semitis eorum
PROV|1|16|pedes enim illorum ad malum currunt et festinant ut effundant sanguinem
PROV|1|17|frustra autem iacitur rete ante oculos pinnatorum
PROV|1|18|ipsique contra sanguinem suum insidiantur et moliuntur fraudes contra animas suas
PROV|1|19|sic semitae omnis avari animas possidentium rapiunt
PROV|1|20|sapientia foris praedicat in plateis dat vocem suam
PROV|1|21|in capite turbarum clamitat in foribus portarum urbis profert verba sua dicens
PROV|1|22|usquequo parvuli diligitis infantiam et stulti ea quae sibi sunt noxia cupiunt et inprudentes odibunt scientiam
PROV|1|23|convertimini ad correptionem meam en proferam vobis spiritum meum et ostendam verba mea
PROV|1|24|quia vocavi et rennuistis extendi manum meam et non fuit qui aspiceret
PROV|1|25|despexistis omne consilium meum et increpationes meas neglexistis
PROV|1|26|ego quoque in interitu vestro ridebo et subsannabo cum vobis quod timebatis advenerit
PROV|1|27|cum inruerit repentina calamitas et interitus quasi tempestas ingruerit quando venerit super vos tribulatio et angustia
PROV|1|28|tunc invocabunt me et non exaudiam mane consurgent et non invenient me
PROV|1|29|eo quod exosam habuerint disciplinam et timorem Domini non susceperint
PROV|1|30|nec adquieverint consilio meo et detraxerint universae correptioni meae
PROV|1|31|comedent igitur fructus viae suae suisque consiliis saturabuntur
PROV|1|32|aversio parvulorum interficiet eos et prosperitas stultorum perdet illos
PROV|1|33|qui autem me audierit absque terrore requiescet et abundantia perfruetur malorum timore sublato
PROV|2|1|fili mi si susceperis sermones meos et mandata mea absconderis penes te
PROV|2|2|ut audiat sapientiam auris tua inclina cor tuum ad noscendam prudentiam
PROV|2|3|si enim sapientiam invocaveris et inclinaveris cor tuum prudentiae
PROV|2|4|si quaesieris eam quasi pecuniam et sicut thesauros effoderis illam
PROV|2|5|tunc intelleges timorem Domini et scientiam Dei invenies
PROV|2|6|quia Dominus dat sapientiam et ex ore eius scientia et prudentia
PROV|2|7|custodiet rectorum salutem et proteget gradientes simpliciter
PROV|2|8|servans semitas iustitiae et vias sanctorum custodiens
PROV|2|9|tunc intelleges iustitiam et iudicium et aequitatem et omnem semitam bonam
PROV|2|10|si intraverit sapientia cor tuum et scientia animae tuae placuerit
PROV|2|11|consilium custodiet te prudentia servabit te
PROV|2|12|ut eruaris de via mala ab homine qui perversa loquitur
PROV|2|13|qui relinquunt iter rectum et ambulant per vias tenebrosas
PROV|2|14|qui laetantur cum malefecerint et exultant in rebus pessimis
PROV|2|15|quorum viae perversae et infames gressus eorum
PROV|2|16|ut eruaris a muliere aliena et ab extranea quae mollit sermones suos
PROV|2|17|et relinquit ducem pubertatis suae
PROV|2|18|et pacti Dei sui oblita est inclinata est enim ad mortem domus eius et ad impios semitae ipsius
PROV|2|19|omnes qui ingrediuntur ad eam non revertentur nec adprehendent semitas vitae
PROV|2|20|ut ambules in via bona et calles iustorum custodias
PROV|2|21|qui enim recti sunt habitabunt in terra et simplices permanebunt in ea
PROV|2|22|impii vero de terra perdentur et qui inique agunt auferentur ex ea
PROV|3|1|fili mi ne obliviscaris legis meae et praecepta mea custodiat cor tuum
PROV|3|2|longitudinem enim dierum et annos vitae et pacem adponent tibi
PROV|3|3|misericordia et veritas non te deserant circumda eas gutturi tuo et describe in tabulis cordis tui
PROV|3|4|et invenies gratiam et disciplinam bonam coram Deo et hominibus
PROV|3|5|habe fiduciam in Domino ex toto corde tuo et ne innitaris prudentiae tuae
PROV|3|6|in omnibus viis tuis cogita illum et ipse diriget gressus tuos
PROV|3|7|ne sis sapiens apud temet ipsum time Dominum et recede a malo
PROV|3|8|sanitas quippe erit umbilico tuo et inrigatio ossuum tuorum
PROV|3|9|honora Dominum de tua substantia et de primitiis omnium frugum tuarum
PROV|3|10|et implebuntur horrea tua saturitate et vino torcularia redundabunt
PROV|3|11|disciplinam Domini fili mi ne abicias nec deficias cum ab eo corriperis
PROV|3|12|quem enim diligit Dominus corripit et quasi pater in filio conplacet sibi
PROV|3|13|beatus homo qui invenit sapientiam et qui affluit prudentia
PROV|3|14|melior est adquisitio eius negotiatione argenti et auro primo fructus eius
PROV|3|15|pretiosior est cunctis opibus et omnia quae desiderantur huic non valent conparari
PROV|3|16|longitudo dierum in dextera eius in sinistra illius divitiae et gloria
PROV|3|17|viae eius viae pulchrae et omnes semitae illius pacificae
PROV|3|18|lignum vitae est his qui adprehenderint eam et qui tenuerit eam beatus
PROV|3|19|Dominus sapientia fundavit terram stabilivit caelos prudentia
PROV|3|20|sapientia illius eruperunt abyssi et nubes rore concrescunt
PROV|3|21|fili mi ne effluant haec ab oculis tuis custodi legem atque consilium
PROV|3|22|et erit vita animae tuae et gratia faucibus tuis
PROV|3|23|tunc ambulabis fiducialiter in via tua et pes tuus non inpinget
PROV|3|24|si dormieris non timebis quiesces et suavis erit somnus tuus
PROV|3|25|ne paveas repentino terrore et inruentes tibi potentias impiorum
PROV|3|26|Dominus enim erit in latere tuo et custodiet pedem tuum ne capiaris
PROV|3|27|noli prohibere benefacere eum qui potest si vales et ipse benefac
PROV|3|28|ne dicas amico tuo vade et revertere et cras dabo tibi cum statim possis dare
PROV|3|29|ne moliaris amico tuo malum cum ille in te habeat fiduciam
PROV|3|30|ne contendas adversus hominem frustra cum ipse tibi nihil mali fecerit
PROV|3|31|ne aemuleris hominem iniustum nec imiteris vias eius
PROV|3|32|quia abominatio Domini est omnis inlusor et cum simplicibus sermocinatio eius
PROV|3|33|egestas a Domino in domo impii habitacula autem iustorum benedicentur
PROV|3|34|inlusores ipse deludet et mansuetis dabit gratiam
PROV|3|35|gloriam sapientes possidebunt stultorum exaltatio ignominia
PROV|4|1|audite filii disciplinam patris et adtendite ut sciatis prudentiam
PROV|4|2|donum bonum tribuam vobis legem meam ne derelinquatis
PROV|4|3|nam et ego filius fui patris mei tenellus et unigenitus coram matre mea
PROV|4|4|et docebat me atque dicebat suscipiat verba mea cor tuum custodi praecepta mea et vives
PROV|4|5|posside sapientiam posside prudentiam ne obliviscaris neque declines a verbis oris mei
PROV|4|6|ne dimittas eam et custodiet te dilige eam et servabit te
PROV|4|7|principium sapientiae posside sapientiam et in omni possessione tua adquire prudentiam
PROV|4|8|arripe illam et exaltabit te glorificaberis ab ea cum eam fueris amplexatus
PROV|4|9|dabit capiti tuo augmenta gratiarum et corona inclita proteget te
PROV|4|10|audi fili mi et suscipe verba mea ut multiplicentur tibi anni vitae
PROV|4|11|viam sapientiae monstravi tibi duxi te per semitas aequitatis
PROV|4|12|quas cum ingressus fueris non artabuntur gressus tui et currens non habebis offendiculum
PROV|4|13|tene disciplinam ne dimittas eam custodi illam quia ipsa est vita tua
PROV|4|14|ne delecteris semitis impiorum nec tibi placeat malorum via
PROV|4|15|fuge ab ea ne transeas per illam declina et desere eam
PROV|4|16|non enim dormiunt nisi malefecerint et rapitur somnus ab eis nisi subplantaverint
PROV|4|17|comedunt panem impietatis et vinum iniquitatis bibunt
PROV|4|18|iustorum autem semita quasi lux splendens procedit et crescit usque ad perfectam diem
PROV|4|19|via impiorum tenebrosa nesciunt ubi corruant
PROV|4|20|fili mi ausculta sermones meos et ad eloquia mea inclina aurem tuam
PROV|4|21|ne recedant ab oculis tuis custodi ea in medio cordis tui
PROV|4|22|vita enim sunt invenientibus ea et universae carni sanitas
PROV|4|23|omni custodia serva cor tuum quia ex ipso vita procedit
PROV|4|24|remove a te os pravum et detrahentia labia sint procul a te
PROV|4|25|oculi tui recta videant et palpebrae tuae praecedant gressus tuos
PROV|4|26|dirige semitam pedibus tuis et omnes viae tuae stabilientur
PROV|4|27|ne declines ad dexteram et ad sinistram averte pedem tuum a malo
PROV|5|1|fili mi adtende sapientiam meam et prudentiae meae inclina aurem tuam
PROV|5|2|ut custodias cogitationes et disciplinam labia tua conservent
PROV|5|3|favus enim stillans labia meretricis et nitidius oleo guttur eius
PROV|5|4|novissima autem illius amara quasi absinthium et acuta quasi gladius biceps
PROV|5|5|pedes eius descendunt in mortem et ad inferos gressus illius penetrant
PROV|5|6|per semitam vitae non ambulat vagi sunt gressus eius et investigabiles
PROV|5|7|nunc ergo fili audi me et ne recedas a verbis oris mei
PROV|5|8|longe fac ab ea viam tuam et ne adpropinques foribus domus eius
PROV|5|9|ne des alienis honorem tuum et annos tuos crudeli
PROV|5|10|ne forte impleantur extranei viribus tuis et labores tui sint in domo aliena
PROV|5|11|et gemas in novissimis quando consumpseris carnes et corpus tuum et dicas
PROV|5|12|cur detestatus sum disciplinam et increpationibus non adquievit cor meum
PROV|5|13|nec audivi vocem docentium me et magistris non inclinavi aurem meam
PROV|5|14|paene fui in omni malo in medio ecclesiae et synagogae
PROV|5|15|bibe aquam de cisterna tua et fluenta putei tui
PROV|5|16|deriventur fontes tui foras et in plateis aquas tuas divide
PROV|5|17|habeto eas solus nec sint alieni participes tui
PROV|5|18|sit vena tua benedicta et laetare cum muliere adulescentiae tuae
PROV|5|19|cerva carissima et gratissimus hinulus ubera eius inebrient te omni tempore in amore illius delectare iugiter
PROV|5|20|quare seduceris fili mi ab aliena et foveris sinu alterius
PROV|5|21|respicit Dominus vias hominis et omnes gressus illius considerat
PROV|5|22|iniquitates suae capiunt impium et funibus peccatorum suorum constringitur
PROV|5|23|ipse morietur quia non habuit disciplinam et multitudine stultitiae suae decipietur
PROV|6|1|fili mi si spoponderis pro amico tuo defixisti apud extraneum manum tuam
PROV|6|2|inlaqueatus es verbis oris tui et captus propriis sermonibus
PROV|6|3|fac ergo quod dico fili mi et temet ipsum libera quia incidisti in manu proximi tui discurre festina suscita amicum tuum
PROV|6|4|ne dederis somnum oculis tuis nec dormitent palpebrae tuae
PROV|6|5|eruere quasi dammula de manu et quasi avis de insidiis aucupis
PROV|6|6|vade ad formicam o piger et considera vias eius et disce sapientiam
PROV|6|7|quae cum non habeat ducem nec praeceptorem nec principem
PROV|6|8|parat aestate cibum sibi et congregat in messe quod comedat
PROV|6|9|usquequo piger dormis quando consurges ex somno tuo
PROV|6|10|paululum dormies paululum dormitabis paululum conseres manus ut dormias
PROV|6|11|et veniet tibi quasi viator egestas et pauperies quasi vir armatus
PROV|6|12|homo apostata vir inutilis graditur ore perverso
PROV|6|13|annuit oculis terit pede digito loquitur
PROV|6|14|pravo corde machinatur malum et in omni tempore iurgia seminat
PROV|6|15|huic extemplo veniet perditio sua et subito conteretur nec habebit ultra medicinam
PROV|6|16|sex sunt quae odit Dominus et septimum detestatur anima eius
PROV|6|17|oculos sublimes linguam mendacem manus effundentes innoxium sanguinem
PROV|6|18|cor machinans cogitationes pessimas pedes veloces ad currendum in malum
PROV|6|19|proferentem mendacia testem fallacem et eum qui seminat inter fratres discordias
PROV|6|20|conserva fili mi praecepta patris tui et ne dimittas legem matris tuae
PROV|6|21|liga ea in corde tuo iugiter et circumda gutturi tuo
PROV|6|22|cum ambulaveris gradiantur tecum cum dormieris custodiant te et evigilans loquere cum eis
PROV|6|23|quia mandatum lucerna est et lex lux et via vitae increpatio disciplinae
PROV|6|24|ut custodiant te a muliere mala et a blanda lingua extraneae
PROV|6|25|non concupiscat pulchritudinem eius cor tuum nec capiaris nutibus illius
PROV|6|26|pretium enim scorti vix unius est panis mulier autem viri pretiosam animam capit
PROV|6|27|numquid abscondere potest homo ignem in sinu suo ut vestimenta illius non ardeant
PROV|6|28|aut ambulare super prunas et non conburentur plantae eius
PROV|6|29|sic qui ingreditur ad mulierem proximi sui non erit mundus cum tetigerit eam
PROV|6|30|non grandis est culpae cum quis furatus fuerit furatur enim ut esurientem impleat animam
PROV|6|31|deprehensus quoque reddet septuplum et omnem substantiam domus suae tradet
PROV|6|32|qui autem adulter est propter cordis inopiam perdet animam suam
PROV|6|33|turpitudinem et ignominiam congregat sibi et obprobrium illius non delebitur
PROV|6|34|quia zelus et furor viri non parcet in die vindictae
PROV|6|35|nec adquiescet cuiusquam precibus nec suscipiet pro redemptione dona plurima
PROV|7|1|fili mi custodi sermones meos et praecepta mea reconde tibi
PROV|7|2|serva mandata mea et vives et legem meam quasi pupillam oculi tui
PROV|7|3|liga eam in digitis tuis scribe illam in tabulis cordis tui
PROV|7|4|dic sapientiae soror mea es et prudentiam voca amicam tuam
PROV|7|5|ut custodiat te a muliere extranea et ab aliena quae verba sua dulcia facit
PROV|7|6|de fenestra enim domus meae per cancellos prospexi
PROV|7|7|et video parvulos considero vecordem iuvenem
PROV|7|8|qui transit in platea iuxta angulum et propter viam domus illius graditur
PROV|7|9|in obscuro advesperascente die in noctis tenebris et caligine
PROV|7|10|et ecce mulier occurrit illi ornatu meretricio praeparata ad capiendas animas garrula et vaga
PROV|7|11|quietis inpatiens nec valens in domo consistere pedibus suis
PROV|7|12|nunc foris nunc in plateis nunc iuxta angulos insidians
PROV|7|13|adprehensumque deosculatur iuvenem et procaci vultu blanditur dicens
PROV|7|14|victimas pro salute debui hodie reddidi vota mea
PROV|7|15|idcirco egressa sum in occursum tuum desiderans te videre et repperi
PROV|7|16|intexui funibus lectum meum stravi tapetibus pictis ex Aegypto
PROV|7|17|aspersi cubile meum murra et aloe et cinnamomo
PROV|7|18|veni inebriemur uberibus donec inlucescat dies et fruamur cupitis amplexibus
PROV|7|19|non est enim vir in domo sua abiit via longissima
PROV|7|20|sacculum pecuniae secum tulit in die plenae lunae reversurus est domum suam
PROV|7|21|inretivit eum multis sermonibus et blanditiis labiorum protraxit illum
PROV|7|22|statim eam sequitur quasi bos ductus ad victimam et quasi agnus lasciviens et ignorans quod ad vincula stultus trahatur
PROV|7|23|donec transfigat sagitta iecur eius velut si avis festinet ad laqueum et nescit quia de periculo animae illius agitur
PROV|7|24|nunc ergo fili audi me et adtende verba oris mei
PROV|7|25|ne abstrahatur in viis illius mens tua neque decipiaris semitis eius
PROV|7|26|multos enim vulneratos deiecit et fortissimi quique interfecti sunt ab ea
PROV|7|27|viae inferi domus eius penetrantes interiora mortis
PROV|8|1|numquid non sapientia clamitat et prudentia dat vocem suam
PROV|8|2|in summis excelsisque verticibus super viam in mediis semitis stans
PROV|8|3|iuxta portas civitatis in ipsis foribus loquitur dicens
PROV|8|4|o viri ad vos clamito et vox mea ad filios hominum
PROV|8|5|intellegite parvuli astutiam et insipientes animadvertite
PROV|8|6|audite quoniam de rebus magnis locutura sum et aperientur labia mea ut recta praedicent
PROV|8|7|veritatem meditabitur guttur meum et labia mea detestabuntur impium
PROV|8|8|iusti sunt omnes sermones mei non est in eis pravum quid neque perversum
PROV|8|9|recti sunt intellegentibus et aequi invenientibus scientiam
PROV|8|10|accipite disciplinam meam et non pecuniam doctrinam magis quam aurum eligite
PROV|8|11|melior est enim sapientia cunctis pretiosissimis et omne desiderabile ei non potest conparari
PROV|8|12|ego sapientia habito in consilio et eruditis intersum cogitationibus
PROV|8|13|timor Domini odit malum arrogantiam et superbiam et viam pravam et os bilingue detestor
PROV|8|14|meum est consilium et aequitas mea prudentia mea est fortitudo
PROV|8|15|per me reges regnant et legum conditores iusta decernunt
PROV|8|16|per me principes imperant et potentes decernunt iustitiam
PROV|8|17|ego diligentes me diligo et qui mane vigilant ad me invenient me
PROV|8|18|mecum sunt divitiae et gloria opes superbae et iustitia
PROV|8|19|melior est fructus meus auro et pretioso lapide et genimina mea argento electo
PROV|8|20|in viis iustitiae ambulo in medio semitarum iudicii
PROV|8|21|ut ditem diligentes me et thesauros eorum repleam
PROV|8|22|Dominus possedit me initium viarum suarum antequam quicquam faceret a principio
PROV|8|23|ab aeterno ordita sum et ex antiquis antequam terra fieret
PROV|8|24|necdum erant abyssi et ego iam concepta eram necdum fontes aquarum eruperant
PROV|8|25|necdum montes gravi mole constiterant ante colles ego parturiebar
PROV|8|26|adhuc terram non fecerat et flumina et cardines orbis terrae
PROV|8|27|quando praeparabat caelos aderam quando certa lege et gyro vallabat abyssos
PROV|8|28|quando aethera firmabat sursum et librabat fontes aquarum
PROV|8|29|quando circumdabat mari terminum suum et legem ponebat aquis ne transirent fines suos quando adpendebat fundamenta terrae
PROV|8|30|cum eo eram cuncta conponens et delectabar per singulos dies ludens coram eo omni tempore
PROV|8|31|ludens in orbe terrarum et deliciae meae esse cum filiis hominum
PROV|8|32|nunc ergo filii audite me beati qui custodiunt vias meas
PROV|8|33|audite disciplinam et estote sapientes et nolite abicere eam
PROV|8|34|beatus homo qui audit me qui vigilat ad fores meas cotidie et observat ad postes ostii mei
PROV|8|35|qui me invenerit inveniet vitam et hauriet salutem a Domino
PROV|8|36|qui autem in me peccaverit laedet animam suam omnes qui me oderunt diligunt mortem
PROV|9|1|sapientia aedificavit sibi domum excidit columnas septem
PROV|9|2|immolavit victimas suas miscuit vinum et proposuit mensam suam
PROV|9|3|misit ancillas suas ut vocarent ad arcem et ad moenia civitatis
PROV|9|4|si quis est parvulus veniat ad me et insipientibus locuta est
PROV|9|5|venite comedite panem meum et bibite vinum quod miscui vobis
PROV|9|6|relinquite infantiam et vivite et ambulate per vias prudentiae
PROV|9|7|qui erudit derisorem ipse sibi facit iniuriam et qui arguit impium generat maculam sibi
PROV|9|8|noli arguere derisorem ne oderit te argue sapientem et diliget te
PROV|9|9|da sapienti et addetur ei sapientia doce iustum et festinabit accipere
PROV|9|10|principium sapientiae timor Domini et scientia sanctorum prudentia
PROV|9|11|per me enim multiplicabuntur dies tui et addentur tibi anni vitae
PROV|9|12|si sapiens fueris tibimet ipsi eris si inlusor solus portabis malum
PROV|9|13|mulier stulta et clamosa plenaque inlecebris et nihil omnino sciens
PROV|9|14|sedit in foribus domus suae super sellam in excelso urbis loco
PROV|9|15|ut vocaret transeuntes viam et pergentes itinere suo
PROV|9|16|quis est parvulus declinet ad me et vecordi locuta est
PROV|9|17|aquae furtivae dulciores sunt et panis absconditus suavior
PROV|9|18|et ignoravit quod gigantes ibi sint et in profundis inferni convivae eius
PROV|10|1|parabolae Salomonis filius sapiens laetificat patrem filius vero stultus maestitia est matris suae
PROV|10|2|non proderunt thesauri impietatis iustitia vero liberabit a morte
PROV|10|3|non adfliget Dominus fame animam iusti et insidias impiorum subvertet
PROV|10|4|egestatem operata est manus remissa manus autem fortium divitias parat
PROV|10|5|qui congregat in messe filius sapiens est qui autem stertit aestate filius confusionis
PROV|10|6|benedictio super caput iusti os autem impiorum operit iniquitatem
PROV|10|7|memoria iusti cum laudibus et nomen impiorum putrescet
PROV|10|8|sapiens corde praecepta suscipiet stultus caeditur labiis
PROV|10|9|qui ambulat simpliciter ambulat confidenter qui autem depravat vias suas manifestus erit
PROV|10|10|qui annuit oculo dabit dolorem stultus labiis verberabitur
PROV|10|11|vena vitae os iusti et os impiorum operiet iniquitatem
PROV|10|12|odium suscitat rixas et universa delicta operit caritas
PROV|10|13|in labiis sapientis invenietur sapientia et virga in dorso eius qui indiget corde
PROV|10|14|sapientes abscondunt scientiam os autem stulti confusioni proximum est
PROV|10|15|substantia divitis urbs fortitudinis eius pavor pauperum egestas eorum
PROV|10|16|opus iusti ad vitam fructus impii ad peccatum
PROV|10|17|via vitae custodienti disciplinam qui autem increpationes relinquit errat
PROV|10|18|abscondunt odium labia mendacia qui profert contumeliam insipiens est
PROV|10|19|in multiloquio peccatum non deerit qui autem moderatur labia sua prudentissimus est
PROV|10|20|argentum electum lingua iusti cor impiorum pro nihilo
PROV|10|21|labia iusti erudiunt plurimos qui autem indocti sunt in cordis egestate morientur
PROV|10|22|benedictio Domini divites facit nec sociabitur ei adflictio
PROV|10|23|quasi per risum stultus operatur scelus sapientia autem est viro prudentia
PROV|10|24|quod timet impius veniet super eum desiderium suum iustis dabitur
PROV|10|25|quasi tempestas transiens non erit impius iustus autem quasi fundamentum sempiternum
PROV|10|26|sicut acetum dentibus et fumus oculis sic piger his qui miserunt eum
PROV|10|27|timor Domini adponet dies et anni impiorum breviabuntur
PROV|10|28|expectatio iustorum laetitia spes autem impiorum peribit
PROV|10|29|fortitudo simplicis via Domini et pavor his qui operantur malum
PROV|10|30|iustus in aeternum non commovebitur impii autem non habitabunt in terram
PROV|10|31|os iusti parturiet sapientiam lingua pravorum peribit
PROV|10|32|labia iusti considerant placita et os impiorum perversa
PROV|11|1|statera dolosa abominatio apud Dominum et pondus aequum voluntas eius
PROV|11|2|ubi fuerit superbia ibi erit et contumelia ubi autem humilitas ibi et sapientia
PROV|11|3|simplicitas iustorum diriget eos et subplantatio perversorum vastabit illos
PROV|11|4|non proderunt divitiae in die ultionis iustitia autem liberabit a morte
PROV|11|5|iustitia simplicis diriget viam eius et in impietate sua corruet impius
PROV|11|6|iustitia rectorum liberabit eos et in insidiis suis capientur iniqui
PROV|11|7|mortuo homine impio nulla erit ultra spes et expectatio sollicitorum peribit
PROV|11|8|iustus de angustia liberatus est et tradetur impius pro eo
PROV|11|9|simulator ore decipit amicum suum iusti autem liberabuntur scientia
PROV|11|10|in bonis iustorum exultabit civitas et in perditione impiorum erit laudatio
PROV|11|11|benedictione iustorum exaltabitur civitas et ore impiorum subvertetur
PROV|11|12|qui despicit amicum suum indigens corde est vir autem prudens tacebit
PROV|11|13|qui ambulat fraudulenter revelat arcana qui autem fidelis est animi celat commissum
PROV|11|14|ubi non est gubernator populus corruet salus autem ubi multa consilia
PROV|11|15|adfligetur malo qui fidem facit pro extraneo qui autem cavet laqueos securus erit
PROV|11|16|mulier gratiosa inveniet gloriam et robusti habebunt divitias
PROV|11|17|benefacit animae suae vir misericors qui autem crudelis est et propinquos abicit
PROV|11|18|impius facit opus instabile seminanti autem iustitiam merces fidelis
PROV|11|19|clementia praeparat vitam et sectatio malorum mortem
PROV|11|20|abominabile Domino pravum cor et voluntas eius in his qui simpliciter ambulant
PROV|11|21|manus in manu non erit innocens malus semen autem iustorum salvabitur
PROV|11|22|circulus aureus in naribus suis mulier pulchra et fatua
PROV|11|23|desiderium iustorum omne bonum est praestolatio impiorum furor
PROV|11|24|alii dividunt propria et ditiores fiunt alii rapiunt non sua et semper in egestate sunt
PROV|11|25|anima quae benedicit inpinguabitur et qui inebriat ipse quoque inebriabitur
PROV|11|26|qui abscondit frumenta maledicetur in populis benedictio autem super caput vendentium
PROV|11|27|bene consurgit diluculo qui quaerit bona qui autem investigator malorum est opprimetur ab eis
PROV|11|28|qui confidet in divitiis suis corruet iusti autem quasi virens folium germinabunt
PROV|11|29|qui conturbat domum suam possidebit ventos et qui stultus est serviet sapienti
PROV|11|30|fructus iusti lignum vitae et qui suscipit animas sapiens est
PROV|11|31|si iustus in terra recipit quanto magis impius et peccator
PROV|12|1|qui diligit disciplinam diligit scientiam qui autem odit increpationes insipiens est
PROV|12|2|qui bonus est hauriet a Domino gratiam qui autem confidit cogitationibus suis impie agit
PROV|12|3|non roborabitur homo ex impietate et radix iustorum non commovebitur
PROV|12|4|mulier diligens corona viro suo et putredo in ossibus eius quae confusione res dignas gerit
PROV|12|5|cogitationes iustorum iudicia et consilia impiorum fraudulentia
PROV|12|6|verba impiorum insidiantur sanguini os iustorum liberabit eos
PROV|12|7|verte impios et non erunt domus autem iustorum permanebit
PROV|12|8|doctrina sua noscetur vir qui autem vanus et excors est patebit contemptui
PROV|12|9|melior est pauper et sufficiens sibi quam gloriosus et indigens pane
PROV|12|10|novit iustus animas iumentorum suorum viscera autem impiorum crudelia
PROV|12|11|qui operatur terram suam saturabitur panibus qui autem sectatur otium stultissimus est
PROV|12|12|desiderium impii munimentum est pessimorum radix autem iustorum proficiet
PROV|12|13|propter peccata labiorum ruina proximat malo effugiet autem iustus de angustia
PROV|12|14|de fructu oris sui unusquisque replebitur bonis et iuxta opera manuum suarum retribuetur ei
PROV|12|15|via stulti recta in oculis eius qui autem sapiens est audit consilia
PROV|12|16|fatuus statim indicat iram suam qui autem dissimulat iniuriam callidus est
PROV|12|17|qui quod novit loquitur index iustitiae est qui autem mentitur testis est fraudulentus
PROV|12|18|est qui promittit et quasi gladio pungitur conscientiae lingua autem sapientium sanitas est
PROV|12|19|labium veritatis firmum erit in perpetuum qui autem testis est repentinus concinnat linguam mendacii
PROV|12|20|dolus in corde cogitantium mala qui autem ineunt pacis consilia sequitur eos gaudium
PROV|12|21|non contristabit iustum quicquid ei acciderit impii autem replebuntur malo
PROV|12|22|abominatio Domino labia mendacia qui autem fideliter agunt placent ei
PROV|12|23|homo versutus celat scientiam et cor insipientium provocabit stultitiam
PROV|12|24|manus fortium dominabitur quae autem remissa est tributis serviet
PROV|12|25|maeror in corde viri humiliabit illud et sermone bono laetificabitur
PROV|12|26|qui neglegit damnum propter amicum iustus est iter autem impiorum decipiet eos
PROV|12|27|non inveniet fraudulentus lucrum et substantia hominis erit auri pretium
PROV|12|28|in semita iustitiae vita iter autem devium ducit ad mortem
PROV|13|1|filius sapiens doctrina patris qui autem inlusor est non audit cum arguitur
PROV|13|2|de fructu oris homo saturabitur bonis anima autem praevaricatorum iniqua
PROV|13|3|qui custodit os suum custodit animam suam qui autem inconsideratus est ad loquendum sentiet mala
PROV|13|4|vult et non vult piger anima autem operantium inpinguabitur
PROV|13|5|verbum mendax iustus detestabitur impius confundit et confundetur
PROV|13|6|iustitia custodit innocentis viam impietas vero peccato subplantat
PROV|13|7|est quasi dives cum nihil habeat et est quasi pauper cum in multis divitiis sit
PROV|13|8|redemptio animae viri divitiae suae qui autem pauper est increpationem non sustinet
PROV|13|9|lux iustorum laetificat lucerna autem impiorum extinguetur
PROV|13|10|inter superbos semper iurgia sunt qui autem agunt cuncta consilio reguntur sapientia
PROV|13|11|substantia festinata minuetur quae autem paulatim colligitur manu multiplicabitur
PROV|13|12|spes quae differtur adfligit animam lignum vitae desiderium veniens
PROV|13|13|qui detrahit alicui rei ipse se in futurum obligat qui autem timet praeceptum in pace versabitur
PROV|13|14|lex sapientis fons vitae ut declinet a ruina mortis
PROV|13|15|doctrina bona dabit gratiam in itinere contemptorum vorago
PROV|13|16|astutus omnia agit cum consilio qui autem fatuus est aperit stultitiam
PROV|13|17|nuntius impii cadet in malum legatus fidelis sanitas
PROV|13|18|egestas et ignominia ei qui deserit disciplinam qui autem adquiescit arguenti glorificabitur
PROV|13|19|desiderium si conpleatur delectat animam detestantur stulti eos qui fugiunt mala
PROV|13|20|qui cum sapientibus graditur sapiens erit amicus stultorum efficietur similis
PROV|13|21|peccatores persequetur malum et iustis retribuentur bona
PROV|13|22|bonus relinquet heredes filios et nepotes et custoditur iusto substantia peccatoris
PROV|13|23|multi cibi in novalibus patrum et alii congregantur absque iudicio
PROV|13|24|qui parcit virgae suae odit filium suum qui autem diligit illum instanter erudit
PROV|13|25|iustus comedit et replet animam suam venter autem impiorum insaturabilis
PROV|14|1|sapiens mulier aedificavit domum suam insipiens instructam quoque destruet manibus
PROV|14|2|ambulans recto itinere et timens Deum despicitur ab eo qui infami graditur via
PROV|14|3|in ore stulti virga superbiae labia sapientium custodiunt eos
PROV|14|4|ubi non sunt boves praesepe vacuum est ubi autem plurimae segetes ibi manifesta fortitudo bovis
PROV|14|5|testis fidelis non mentietur profert mendacium testis dolosus
PROV|14|6|quaerit derisor sapientiam et non inveniet doctrina prudentium facilis
PROV|14|7|vade contra virum stultum et nescito labia prudentiae
PROV|14|8|sapientia callidi est intellegere viam suam et inprudentia stultorum errans
PROV|14|9|stultis inludet peccatum inter iustos morabitur gratia
PROV|14|10|cor quod novit amaritudinem animae suae in gaudio eius non miscebitur extraneus
PROV|14|11|domus impiorum delebitur tabernacula iustorum germinabunt
PROV|14|12|est via quae videtur homini iusta novissima autem eius deducunt ad mortem
PROV|14|13|risus dolore miscebitur et extrema gaudii luctus occupat
PROV|14|14|viis suis replebitur stultus et super eum erit vir bonus
PROV|14|15|innocens credit omni verbo astutus considerat gressus suos
PROV|14|16|sapiens timet et declinat malum stultus transilit et confidit
PROV|14|17|inpatiens operabitur stultitiam et vir versutus odiosus est
PROV|14|18|possidebunt parvuli stultitiam et astuti expectabunt scientiam
PROV|14|19|iacebunt mali ante bonos et impii ante portas iustorum
PROV|14|20|etiam proximo suo pauper odiosus erit amici vero divitum multi
PROV|14|21|qui despicit proximum suum peccat qui autem miseretur pauperi beatus erit
PROV|14|22|errant qui operantur malum misericordia et veritas praeparant bona
PROV|14|23|in omni opere erit abundantia ubi autem verba sunt plurima frequenter egestas
PROV|14|24|corona sapientium divitiae eorum fatuitas stultorum inprudentia
PROV|14|25|liberat animas testis fidelis et profert mendacia versipellis
PROV|14|26|in timore Domini fiducia fortitudinis et filiis eius erit spes
PROV|14|27|timor Domini fons vitae ut declinet a ruina mortis
PROV|14|28|in multitudine populi dignitas regis et in paucitate plebis ignominia principis
PROV|14|29|qui patiens est multa gubernatur prudentia qui autem inpatiens exaltat stultitiam suam
PROV|14|30|vita carnium sanitas cordis putredo ossuum invidia
PROV|14|31|qui calumniatur egentem exprobrat factori eius honorat autem eum qui miseretur pauperis
PROV|14|32|in malitia sua expelletur impius sperat autem iustus in morte sua
PROV|14|33|in corde prudentis requiescit sapientia et indoctos quoque erudiet
PROV|14|34|iustitia elevat gentem miseros facit populos peccatum
PROV|14|35|acceptus est regi minister intellegens iracundiam eius inutilis sustinebit
PROV|15|1|responsio mollis frangit iram sermo durus suscitat furorem
PROV|15|2|lingua sapientium ornat scientiam os fatuorum ebullit stultitiam
PROV|15|3|in omni loco oculi Domini contemplantur malos et bonos
PROV|15|4|lingua placabilis lignum vitae quae inmoderata est conteret spiritum
PROV|15|5|stultus inridet disciplinam patris sui qui autem custodit increpationes astutior fiet
PROV|15|6|domus iusti plurima fortitudo et in fructibus impii conturbatur
PROV|15|7|labia sapientium disseminabunt scientiam cor stultorum dissimile erit
PROV|15|8|victimae impiorum abominabiles Domino vota iustorum placabilia
PROV|15|9|abominatio est Domino via impii qui sequitur iustitiam diligetur ab eo
PROV|15|10|doctrina mala deserenti viam qui increpationes odit morietur
PROV|15|11|infernus et perditio coram Domino quanto magis corda filiorum hominum
PROV|15|12|non amat pestilens eum qui se corripit nec ad sapientes graditur
PROV|15|13|cor gaudens exhilarat faciem in maerore animi deicitur spiritus
PROV|15|14|cor sapientis quaerit doctrinam et os stultorum pascetur inperitia
PROV|15|15|omnes dies pauperis mali secura mens quasi iuge convivium
PROV|15|16|melius est parum cum timore Domini quam thesauri magni et insatiabiles
PROV|15|17|melius est vocare ad holera cum caritate quam ad vitulum saginatum cum odio
PROV|15|18|vir iracundus provocat rixas qui patiens est mitigat suscitatas
PROV|15|19|iter pigrorum quasi sepes spinarum via iustorum absque offendiculo
PROV|15|20|filius sapiens laetificat patrem et stultus homo despicit matrem suam
PROV|15|21|stultitia gaudium stulto et vir prudens dirigit gressus
PROV|15|22|dissipantur cogitationes ubi non est consilium ubi vero plures sunt consiliarii confirmantur
PROV|15|23|laetatur homo in sententia oris sui et sermo oportunus est optimus
PROV|15|24|semita vitae super eruditum ut declinet de inferno novissimo
PROV|15|25|domum superborum demolietur Dominus et firmos facit terminos viduae
PROV|15|26|abominatio Domini cogitationes malae et purus sermo pulcherrimus
PROV|15|27|conturbat domum suam qui sectatur avaritiam qui autem odit munera vivet
PROV|15|28|mens iusti meditatur oboedientiam os impiorum redundat malis
PROV|15|29|longe est Dominus ab impiis et orationes iustorum exaudiet
PROV|15|30|lux oculorum laetificat animam fama bona inpinguat ossa
PROV|15|31|auris quae audit increpationes vitae in medio sapientium commorabitur
PROV|15|32|qui abicit disciplinam despicit animam suam qui adquiescit increpationibus possessor est cordis
PROV|15|33|timor Domini disciplina sapientiae et gloriam praecedit humilitas
PROV|16|1|hominis est animum praeparare et Dei gubernare linguam
PROV|16|2|omnes viae hominum patent oculis eius spirituum ponderator est Dominus
PROV|16|3|revela Domino opera tua et dirigentur cogitationes tuae
PROV|16|4|universa propter semet ipsum operatus est Dominus impium quoque ad diem malum
PROV|16|5|abominatio Domini omnis arrogans etiam si manus ad manum fuerit non erit innocens
PROV|16|6|misericordia et veritate redimitur iniquitas et in timore Domini declinatur a malo
PROV|16|7|cum placuerint Domino viae hominis inimicos quoque eius convertet ad pacem
PROV|16|8|melius est parum cum iustitia quam multi fructus cum iniquitate
PROV|16|9|cor hominis disponet viam suam sed Domini est dirigere gressus eius
PROV|16|10|divinatio in labiis regis in iudicio non errabit os eius
PROV|16|11|pondus et statera iudicia Domini sunt et opera eius omnes lapides sacculi
PROV|16|12|abominabiles regi qui agunt impie quoniam iustitia firmatur solium
PROV|16|13|voluntas regum labia iusta qui recta loquitur diligetur
PROV|16|14|indignatio regis nuntii mortis et vir sapiens placabit eam
PROV|16|15|in hilaritate vultus regis vita et clementia eius quasi imber serotinus
PROV|16|16|posside sapientiam quia auro melior est et adquire prudentiam quia pretiosior est argento
PROV|16|17|semita iustorum declinat mala custos animae suae servat viam suam
PROV|16|18|contritionem praecedit superbia et ante ruinam exaltatur spiritus
PROV|16|19|melius est humiliari cum mitibus quam dividere spolia cum superbis
PROV|16|20|eruditus in verbo repperiet bona et qui in Domino sperat beatus est
PROV|16|21|qui sapiens corde est appellabitur prudens et qui dulcis eloquio maiora percipiet
PROV|16|22|fons vitae eruditio possidentis doctrina stultorum fatuitas
PROV|16|23|cor sapientis erudiet os eius et labiis illius addet gratiam
PROV|16|24|favus mellis verba conposita dulcedo animae et sanitas ossuum
PROV|16|25|est via quae videtur homini recta et novissimum eius ducit ad mortem
PROV|16|26|anima laborantis laborat sibi quia conpulit eum os suum
PROV|16|27|vir impius fodit malum et in labiis eius ignis ardescit
PROV|16|28|homo perversus suscitat lites et verbosus separat principes
PROV|16|29|vir iniquus lactat amicum suum et ducit eum per viam non bonam
PROV|16|30|qui adtonitis oculis cogitat prava mordens labia sua perficit malum
PROV|16|31|corona dignitatis senectus in viis iustitiae repperietur
PROV|16|32|melior est patiens viro forte et qui dominatur animo suo expugnatore urbium
PROV|16|33|sortes mittuntur in sinu sed a Domino temperantur
PROV|17|1|melior est buccella sicca cum gaudio quam domus plena victimis cum iurgio
PROV|17|2|servus sapiens dominabitur filiis stultis et inter fratres hereditatem dividet
PROV|17|3|sicut igne probatur argentum et aurum camino ita corda probat Dominus
PROV|17|4|malus oboedit linguae iniquae et fallax obtemperat labiis mendacibus
PROV|17|5|qui despicit pauperem exprobrat factori eius et qui in ruina laetatur alterius non erit inpunitus
PROV|17|6|corona senum filii filiorum et gloria filiorum patres sui
PROV|17|7|non decent stultum verba conposita nec principem labium mentiens
PROV|17|8|gemma gratissima expectatio praestolantis quocumque se verterit prudenter intellegit
PROV|17|9|qui celat delictum quaerit amicitias qui altero sermone repetit separat foederatos
PROV|17|10|plus proficit correptio apud prudentem quam centum plagae apud stultum
PROV|17|11|semper iurgia quaerit malus angelus autem crudelis mittetur contra eum
PROV|17|12|expedit magis ursae occurrere raptis fetibus quam fatuo confidenti sibi in stultitia sua
PROV|17|13|qui reddit mala pro bonis non recedet malum de domo eius
PROV|17|14|qui dimittit aquam caput est iurgiorum et antequam patiatur contumeliam iudicium deserit
PROV|17|15|et qui iustificat impium et qui condemnat iustum abominabilis est uterque apud Dominum
PROV|17|16|quid prodest habere divitias stultum cum sapientiam emere non possit
PROV|17|17|omni tempore diligit qui amicus est et frater in angustiis conprobatur
PROV|17|18|homo stultus plaudet manibus cum spoponderit pro amico suo
PROV|17|19|qui meditatur discordiam diligit rixas et qui exaltat ostium quaerit ruinam
PROV|17|20|qui perversi cordis est non inveniet bonum et qui vertit linguam incidet in malum
PROV|17|21|natus est stultus in ignominiam suam sed nec pater in fatuo laetabitur
PROV|17|22|animus gaudens aetatem floridam facit spiritus tristis exsiccat ossa
PROV|17|23|munera de sinu impius accipit ut pervertat semitas iudicii
PROV|17|24|in facie prudentis lucet sapientia oculi stultorum in finibus terrae
PROV|17|25|ira patris filius stultus et dolor matris quae genuit eum
PROV|17|26|non est bonum damnum inferre iusto nec percutere principem qui recta iudicat
PROV|17|27|qui moderatur sermones suos doctus et prudens est et pretiosi spiritus vir eruditus
PROV|17|28|stultus quoque si tacuerit sapiens putabitur et si conpresserit labia sua intellegens
PROV|18|1|occasiones quaerit qui vult recedere ab amico omni tempore erit exprobrabilis
PROV|18|2|non recipit stultus verba prudentiae nisi ea dixeris quae versantur in corde eius
PROV|18|3|impius cum in profundum venerit peccatorum contemnit sed sequitur eum ignominia et obprobrium
PROV|18|4|aqua profunda verba ex ore viri et torrens redundans fons sapientiae
PROV|18|5|accipere personam impii non est bonum ut declines a veritate iudicii
PROV|18|6|labia stulti inmiscunt se rixis et os eius iurgia provocat
PROV|18|7|os stulti contritio eius et labia illius ruina animae eius
PROV|18|8|verba bilinguis quasi simplicia et ipsa perveniunt usque ad interiora ventris
PROV|18|9|qui mollis et dissolutus est in opere suo frater est sua opera dissipantis
PROV|18|10|turris fortissima nomen Domini ad ipsum currit iustus et exaltabitur
PROV|18|11|substantia divitis urbs roboris eius et quasi murus validus circumdans eum
PROV|18|12|antequam conteratur exaltatur cor hominis et antequam glorificetur humiliatur
PROV|18|13|qui prius respondit quam audiat stultum se esse demonstrat et confusione dignum
PROV|18|14|spiritus viri sustentat inbecillitatem suam spiritum vero ad irascendum facilem quis poterit sustinere
PROV|18|15|cor prudens possidebit scientiam et auris sapientium quaerit doctrinam
PROV|18|16|donum hominis dilatat viam eius et ante principes spatium ei facit
PROV|18|17|iustus prior est accusator sui venit amicus eius et investigavit eum
PROV|18|18|contradictiones conprimit sors et inter potentes quoque diiudicat
PROV|18|19|frater qui adiuvatur a fratre quasi civitas firma et iudicia quasi vectes urbium
PROV|18|20|de fructu oris viri replebitur venter eius et genimina labiorum illius saturabunt eum
PROV|18|21|mors et vita in manu linguae qui diligunt eam comedent fructus eius
PROV|18|22|qui invenit mulierem invenit bonum et hauriet iucunditatem a Domino
PROV|18|23|cum obsecrationibus loquetur pauper et dives effabitur rigide
PROV|18|24|vir amicalis ad societatem magis amicus erit quam frater
PROV|19|1|melior est pauper qui ambulat in simplicitate sua quam torquens labia insipiens
PROV|19|2|ubi non est scientia animae non est bonum et qui festinus est pedibus offendit
PROV|19|3|stultitia hominis subplantat gressus eius et contra Deum fervet animo suo
PROV|19|4|divitiae addunt amicos plurimos a paupere autem et hii quos habuit separantur
PROV|19|5|testis falsus non erit inpunitus et qui mendacia loquitur non effugiet
PROV|19|6|multi colunt personam potentis et amici sunt dona tribuenti
PROV|19|7|fratres hominis pauperis oderunt eum insuper et amici procul recesserunt ab eo qui tantum verba sectatur nihil habebit
PROV|19|8|qui autem possessor est mentis diligit animam suam et custos prudentiae inveniet bona
PROV|19|9|testis falsus non erit inpunitus et qui loquitur mendacia peribit
PROV|19|10|non decent stultum deliciae nec servum dominari principibus
PROV|19|11|doctrina viri per patientiam noscitur et gloria eius est iniqua praetergredi
PROV|19|12|sicut fremitus leonis ita et regis ira et sicut ros super herbam ita hilaritas eius
PROV|19|13|dolor patris filius stultus et tecta iugiter perstillantia litigiosa mulier
PROV|19|14|domus et divitiae dantur a patribus a Domino autem proprie uxor prudens
PROV|19|15|pigredo inmittit soporem et anima dissoluta esuriet
PROV|19|16|qui custodit mandatum custodit animam suam qui autem neglegit vias suas mortificabitur
PROV|19|17|feneratur Domino qui miseretur pauperis et vicissitudinem suam reddet ei
PROV|19|18|erudi filium tuum ne desperes ad interfectionem autem eius ne ponas animam tuam
PROV|19|19|qui inpatiens est sustinebit damnum et cum rapuerit aliud adponet
PROV|19|20|audi consilium et suscipe disciplinam ut sis sapiens in novissimis tuis
PROV|19|21|multae cogitationes in corde viri voluntas autem Domini permanebit
PROV|19|22|homo indigens misericors est et melior pauper quam vir mendax
PROV|19|23|timor Domini ad vitam et in plenitudine commorabitur absque visitatione pessimi
PROV|19|24|abscondit piger manum suam sub ascella nec ad os suum adplicat eam
PROV|19|25|pestilente flagellato stultus sapientior erit sin autem corripueris sapientem intelleget disciplinam
PROV|19|26|qui adfligit patrem et fugat matrem ignominiosus est et infelix
PROV|19|27|non cesses fili audire doctrinam nec ignores sermones scientiae
PROV|19|28|testis iniquus deridet iudicium et os impiorum devorat iniquitatem
PROV|19|29|parata sunt derisoribus iudicia et mallei percutientes stultorum corporibus
PROV|20|1|luxuriosa res vinum et tumultuosa ebrietas quicumque his delectatur non erit sapiens
PROV|20|2|sicut rugitus leonis ita terror regis qui provocat eum peccat in animam suam
PROV|20|3|honor est homini qui separat se a contentionibus omnes autem stulti miscentur contumeliis
PROV|20|4|propter frigus piger arare noluit mendicabit ergo aestate et non dabitur ei
PROV|20|5|sicut aqua profunda sic consilium in corde viri sed homo sapiens exhauriet illud
PROV|20|6|multi homines misericordes vocantur virum autem fidelem quis inveniet
PROV|20|7|iustus qui ambulat in simplicitate sua beatos post se filios derelinquet
PROV|20|8|rex qui sedet in solio iudicii dissipat omne malum intuitu suo
PROV|20|9|quis potest dicere mundum est cor meum purus sum a peccato
PROV|20|10|pondus et pondus mensura et mensura utrumque abominabile est apud Deum
PROV|20|11|ex studiis suis intellegitur puer si munda et si recta sint opera eius
PROV|20|12|aurem audientem et oculum videntem Dominus fecit utrumque
PROV|20|13|noli diligere somnum ne te egestas opprimat aperi oculos tuos et saturare panibus
PROV|20|14|malum est malum est dicit omnis emptor et cum recesserit tunc gloriabitur
PROV|20|15|est aurum et multitudo gemmarum vas autem pretiosum labia scientiae
PROV|20|16|tolle vestimentum eius qui fideiussor extitit alieni et pro extraneis aufer pignus ab eo
PROV|20|17|suavis est homini panis mendacii et postea implebitur os eius calculo
PROV|20|18|cogitationes consiliis roborantur et gubernaculis tractanda sunt bella
PROV|20|19|ei qui revelat mysteria et ambulat fraudulenter et dilatat labia sua ne commiscearis
PROV|20|20|qui maledicit patri suo et matri extinguetur lucerna eius in mediis tenebris
PROV|20|21|hereditas ad quam festinatur in principio in novissimo benedictione carebit
PROV|20|22|ne dicas reddam malum expecta Dominum et liberabit te
PROV|20|23|abominatio est apud Deum pondus et pondus statera dolosa non est bona
PROV|20|24|a Domino diriguntur gressus viri quis autem hominum intellegere potest viam suam
PROV|20|25|ruina est hominis devorare sanctos et post vota tractare
PROV|20|26|dissipat impios rex sapiens et curvat super eos fornicem
PROV|20|27|lucerna Domini spiraculum hominis quae investigat omnia secreta ventris
PROV|20|28|misericordia et veritas custodiunt regem et roboratur clementia thronus eius
PROV|20|29|exultatio iuvenum fortitudo eorum et dignitas senum canities
PROV|20|30|livor vulneris absterget mala et plagae in secretioribus ventris
PROV|21|1|sicut divisiones aquarum ita cor regis in manu Domini quocumque voluerit inclinabit illud
PROV|21|2|omnis via viri recta sibi videtur adpendit autem corda Dominus
PROV|21|3|facere misericordiam et iudicium magis placent Domino quam victimae
PROV|21|4|exaltatio oculorum et dilatatio cordis lucerna impiorum peccatum
PROV|21|5|cogitationes robusti semper in abundantia omnis autem piger semper in egestate
PROV|21|6|qui congregat thesauros lingua mendacii vanus est et inpingetur ad laqueos mortis
PROV|21|7|rapinae impiorum detrahent eos quia noluerunt facere iudicium
PROV|21|8|perversa via viri aliena est qui autem mundus est rectum opus eius
PROV|21|9|melius est sedere in angulo domatis quam cum muliere litigiosa et in domo communi
PROV|21|10|anima impii desiderat malum non miserebitur proximo suo
PROV|21|11|multato pestilente sapientior erit parvulus et si sectetur sapientem sumet scientiam
PROV|21|12|excogitat iustus de domo impii ut detrahat impios in malum
PROV|21|13|qui obturat aurem suam ad clamorem pauperis et ipse clamabit et non exaudietur
PROV|21|14|munus absconditum extinguet iras et donum in sinu indignationem maximam
PROV|21|15|gaudium iusto est facere iudicium et pavor operantibus iniquitatem
PROV|21|16|vir qui erraverit a via doctrinae in coetu gigantum commorabitur
PROV|21|17|qui diligit epulas in egestate erit qui amat vinum et pinguia non ditabitur
PROV|21|18|pro iusto datur impius et pro rectis iniquus
PROV|21|19|melius est habitare in terra deserta quam cum muliere rixosa et iracunda
PROV|21|20|thesaurus desiderabilis et oleum in habitaculo iusti et inprudens homo dissipabit illud
PROV|21|21|qui sequitur iustitiam et misericordiam inveniet vitam et iustitiam et gloriam
PROV|21|22|civitatem fortium ascendit sapiens et destruxit robur fiduciae eius
PROV|21|23|qui custodit os suum et linguam suam custodit ab angustiis animam suam
PROV|21|24|superbus et arrogans vocatur indoctus qui in ira operatur superbiam
PROV|21|25|desideria occidunt pigrum noluerunt enim quicquam manus eius operari
PROV|21|26|tota die concupiscit et desiderat qui autem iustus est tribuet et non cessabit
PROV|21|27|hostiae impiorum abominabiles quia offeruntur ex scelere
PROV|21|28|testis mendax peribit vir oboediens loquitur victoriam
PROV|21|29|vir impius procaciter obfirmat vultum suum qui autem rectus est corrigit viam suam
PROV|21|30|non est sapientia non est prudentia non est consilium contra Dominum
PROV|21|31|equus paratur ad diem belli Dominus autem salutem tribuet
PROV|22|1|melius est nomen bonum quam divitiae multae super argentum et aurum gratia bona
PROV|22|2|dives et pauper obviaverunt sibi utriusque operator est Dominus
PROV|22|3|callidus vidit malum et abscondit se innocens pertransiit et adflictus est damno
PROV|22|4|finis modestiae timor Domini divitiae et gloria et vita
PROV|22|5|arma et gladii in via perversi custos animae suae longe recedit ab eis
PROV|22|6|proverbium est adulescens iuxta viam suam etiam cum senuerit non recedet ab ea
PROV|22|7|dives pauperibus imperat et qui accipit mutuum servus est fenerantis
PROV|22|8|qui seminat iniquitatem metet mala et virga irae suae consummabitur
PROV|22|9|qui pronus est ad misericordiam benedicetur de panibus enim suis dedit pauperi
PROV|22|10|eice derisorem et exibit cum eo iurgium cessabuntque causae et contumeliae
PROV|22|11|qui diligit cordis munditiam propter gratiam labiorum suorum habebit amicum regem
PROV|22|12|oculi Domini custodiunt scientiam et subplantantur verba iniqui
PROV|22|13|dicit piger leo foris in medio platearum occidendus sum
PROV|22|14|fovea profunda os alienae cui iratus est Dominus incidet in eam
PROV|22|15|stultitia conligata est in corde pueri et virga disciplinae fugabit eam
PROV|22|16|qui calumniatur pauperem ut augeat divitias suas dabit ipse ditiori et egebit
PROV|22|17|inclina aurem tuam et audi verba sapientium adpone autem cor ad doctrinam meam
PROV|22|18|quae pulchra erit tibi cum servaveris eam in ventre tuo et redundabit in labiis tuis
PROV|22|19|ut sit in Domino fiducia tua unde et ostendi eam tibi hodie
PROV|22|20|ecce descripsi eam tibi tripliciter in cogitationibus et scientia
PROV|22|21|ut ostenderem tibi firmitatem et eloquia veritatis respondere ex his illi qui misit te
PROV|22|22|non facias violentiam pauperi quia pauper est neque conteras egenum in porta
PROV|22|23|quia Dominus iudicabit causam eius et configet eos qui confixerint animam eius
PROV|22|24|noli esse amicus homini iracundo neque ambules cum viro furioso
PROV|22|25|ne forte discas semitas eius et sumas scandalum animae tuae
PROV|22|26|noli esse cum his qui defigunt manus suas et qui vades se offerunt pro debitis
PROV|22|27|si enim non habes unde restituas quid causae est ut tollat operimentum de cubili tuo
PROV|22|28|ne transgrediaris terminos antiquos quos posuerunt patres tui
PROV|22|29|vidisti virum velocem in opere suo coram regibus stabit nec erit ante ignobiles
PROV|23|1|quando sederis ut comedas cum principe diligenter adtende quae posita sunt ante faciem tuam
PROV|23|2|et statue cultrum in gutture tuo si tamen habes in potestate animam tuam
PROV|23|3|ne desideres de cibis eius in quo est panis mendacii
PROV|23|4|noli laborare ut diteris sed prudentiae tuae pone modum
PROV|23|5|ne erigas oculos tuos ad opes quas habere non potes quia facient sibi pinnas quasi aquilae et avolabunt in caelum
PROV|23|6|ne comedas cum homine invido et ne desideres cibos eius
PROV|23|7|quoniam in similitudinem arioli et coniectoris aestimat quod ignorat comede et bibe dicet tibi et mens eius non est tecum
PROV|23|8|cibos quos comederas evomes et perdes pulchros sermones tuos
PROV|23|9|in auribus insipientium ne loquaris quia despicient doctrinam eloquii tui
PROV|23|10|ne adtingas terminos parvulorum et agrum pupillorum ne introeas
PROV|23|11|propinquus enim eorum Fortis est et ipse iudicabit contra te causam illorum
PROV|23|12|ingrediatur ad doctrinam cor tuum et aures tuae ad verba scientiae
PROV|23|13|noli subtrahere a puero disciplinam si enim percusseris eum virga non morietur
PROV|23|14|tu virga percuties eum et animam eius de inferno liberabis
PROV|23|15|fili mi si sapiens fuerit animus tuus gaudebit tecum cor meum
PROV|23|16|et exultabunt renes mei cum locuta fuerint rectum labia tua
PROV|23|17|non aemuletur cor tuum peccatores sed in timore Domini esto tota die
PROV|23|18|quia habebis spem in novissimo et praestolatio tua non auferetur
PROV|23|19|audi fili mi et esto sapiens et dirige in via animum tuum
PROV|23|20|noli esse in conviviis potatorum nec in comesationibus eorum qui carnes ad vescendum conferunt
PROV|23|21|quia vacantes potibus et dantes symbola consumentur et vestietur pannis dormitatio
PROV|23|22|audi patrem tuum qui genuit te et ne contemnas cum senuerit mater tua
PROV|23|23|veritatem eme et noli vendere sapientiam et doctrinam et intellegentiam
PROV|23|24|exultat gaudio pater iusti qui sapientem genuit laetabitur in eo
PROV|23|25|gaudeat pater tuus et mater tua et exultet quae genuit te
PROV|23|26|praebe fili mi cor tuum mihi et oculi tui vias meas custodiant
PROV|23|27|fovea enim profunda est meretrix et puteus angustus aliena
PROV|23|28|insidiatur in via quasi latro et quos incautos viderit interficit
PROV|23|29|cui vae cuius patri vae cui rixae cui foveae cui sine causa vulnera cui suffusio oculorum
PROV|23|30|nonne his qui morantur in vino et student calicibus epotandis
PROV|23|31|ne intuearis vinum quando flavescit cum splenduerit in vitro color eius ingreditur blande
PROV|23|32|sed in novissimo mordebit ut coluber et sicut regulus venena diffundet
PROV|23|33|oculi tui videbunt extraneas et cor tuum loquetur perversa
PROV|23|34|et eris sicut dormiens in medio mari et quasi sopitus gubernator amisso clavo
PROV|23|35|et dices verberaverunt me sed non dolui traxerunt me et ego non sensi quando evigilabo et rursum vina repperiam
PROV|24|1|ne aemuleris viros malos nec desideres esse cum eis
PROV|24|2|quia rapinas meditatur mens eorum et fraudes labia eorum loquuntur
PROV|24|3|sapientia aedificabitur domus et prudentia roborabitur
PROV|24|4|in doctrina replebuntur cellaria universa substantia pretiosa et pulcherrima
PROV|24|5|vir sapiens et fortis est et vir doctus robustus et validus
PROV|24|6|quia cum dispositione initur bellum et erit salus ubi multa consilia sunt
PROV|24|7|excelsa stulto sapientia in porta non aperiet os suum
PROV|24|8|qui cogitat malefacere stultus vocabitur
PROV|24|9|cogitatio stulti peccatum est et abominatio hominum detractor
PROV|24|10|si desperaveris lassus in die angustiae inminuetur fortitudo tua
PROV|24|11|erue eos qui ducuntur ad mortem et qui trahuntur ad interitum liberare ne cesses
PROV|24|12|si dixeris vires non suppetunt qui inspector est cordis ipse intellegit et servatorem animae tuae nihil fallit reddetque homini iuxta opera sua
PROV|24|13|comede fili mi mel quia bonum est et favum dulcissimum gutturi tuo
PROV|24|14|sic et doctrina sapientiae animae tuae quam cum inveneris habebis in novissimis et spes tua non peribit
PROV|24|15|ne insidieris et quaeras impietatem in domo iusti neque vastes requiem eius
PROV|24|16|septies enim cadet iustus et resurget impii autem corruent in malum
PROV|24|17|cum ceciderit inimicus tuus ne gaudeas et in ruina eius ne exultet cor tuum
PROV|24|18|ne forte videat Dominus et displiceat ei et auferat ab eo iram suam
PROV|24|19|ne contendas cum pessimis nec aemuleris impios
PROV|24|20|quoniam non habent futurorum spem mali et lucerna impiorum extinguetur
PROV|24|21|time Dominum fili mi et regem et cum detractoribus non commiscearis
PROV|24|22|quoniam repente consurget perditio eorum et ruinam utriusque quis novit
PROV|24|23|haec quoque sapientibus cognoscere personam in iudicio non est bonum
PROV|24|24|qui dicit impio iustus es maledicent ei populi et detestabuntur eum tribus
PROV|24|25|qui arguunt laudabuntur et super ipsos veniet benedictio
PROV|24|26|labia deosculabitur qui recta verba respondet
PROV|24|27|praepara foris opus tuum et diligenter exerce agrum tuum ut postea aedifices domum tuam
PROV|24|28|ne sis testis frustra contra proximum tuum nec lactes quemquam labiis tuis
PROV|24|29|ne dicas quomodo fecit mihi sic faciam ei reddam unicuique secundum opus suum
PROV|24|30|per agrum hominis pigri transivi et per vineam viri stulti
PROV|24|31|et ecce totum repleverant urticae operuerant superficiem eius spinae et maceria lapidum destructa erat
PROV|24|32|quod cum vidissem posui in corde meo et exemplo didici disciplinam
PROV|24|33|parum inquam dormies modicum dormitabis pauxillum manus conseres ut quiescas
PROV|24|34|et veniet quasi cursor egestas tua et mendicitas quasi vir armatus
PROV|25|1|haec quoque parabolae Salomonis quas transtulerunt viri Ezechiae regis Iuda
PROV|25|2|gloria Dei celare verbum et gloria regum investigare sermonem
PROV|25|3|caelum sursum et terra deorsum et cor regum inscrutabile
PROV|25|4|aufer robiginem de argento et egredietur vas purissimum
PROV|25|5|aufer impietatem de vultu regis et firmabitur iustitia thronus eius
PROV|25|6|ne gloriosus appareas coram rege et in loco magnorum ne steteris
PROV|25|7|melius est enim ut dicatur tibi ascende huc quam ut humilieris coram principe
PROV|25|8|quae viderunt oculi tui ne proferas in iurgio cito ne postea emendare non possis cum dehonestaveris amicum tuum
PROV|25|9|causam tuam tracta cum amico tuo et secretum extraneo non reveles
PROV|25|10|ne forte insultet tibi cum audierit et exprobrare non cesset
PROV|25|11|mala aurea in lectis argenteis qui loquitur verbum in tempore suo
PROV|25|12|inauris aurea et margaritum fulgens qui arguit sapientem et aurem oboedientem
PROV|25|13|sicut frigus nivis in die messis ita legatus fidelis ei qui misit eum animam illius requiescere facit
PROV|25|14|nubes et ventus et pluviae non sequentes vir gloriosus et promissa non conplens
PROV|25|15|patientia lenietur princeps et lingua mollis confringet duritiam
PROV|25|16|mel invenisti comede quod sufficit tibi ne forte saturatus evomas illud
PROV|25|17|subtrahe pedem tuum de domo proximi tui nequando satiatus oderit te
PROV|25|18|iaculum et gladius et sagitta acuta homo qui loquitur contra proximum suum testimonium falsum
PROV|25|19|dens putridus et pes lapsus qui sperat super infideli in die angustiae
PROV|25|20|et amittit pallium in die frigoris acetum in nitro et qui cantat carmina cordi pessimo
PROV|25|21|si esurierit inimicus tuus ciba illum et si sitierit da ei aquam bibere
PROV|25|22|prunam enim congregabis super caput eius et Dominus reddet tibi
PROV|25|23|ventus aquilo dissipat pluvias et facies tristis linguam detrahentem
PROV|25|24|melius est sedere in angulo domatis quam cum muliere litigiosa et in domo communi
PROV|25|25|aqua frigida animae sitienti et nuntius bonus de terra longinqua
PROV|25|26|fons turbatus pede et vena corrupta iustus cadens coram impio
PROV|25|27|sicut qui mel multum comedit non est ei bonum sic qui scrutator est maiestatis opprimitur gloria
PROV|25|28|sicut urbs patens et absque murorum ambitu ita vir qui non potest in loquendo cohibere spiritum suum
PROV|26|1|quomodo nix aestate et pluvia in messe sic indecens est stulto gloria
PROV|26|2|sicut avis ad alia transvolans et passer quolibet vadens sic maledictum frustra prolatum in quempiam superveniet
PROV|26|3|flagellum equo et camus asino et virga dorso inprudentium
PROV|26|4|ne respondeas stulto iuxta stultitiam suam ne efficiaris ei similis
PROV|26|5|responde stulto iuxta stultitiam suam ne sibi sapiens esse videatur
PROV|26|6|claudus pedibus et iniquitatem bibens qui mittit verba per nuntium stultum
PROV|26|7|quomodo pulchras frustra habet claudus tibias sic indecens est in ore stultorum parabola
PROV|26|8|sicut qui mittit lapidem in acervum Mercurii ita qui tribuit insipienti honorem
PROV|26|9|quomodo si spina nascatur in manu temulenti sic parabola in ore stultorum
PROV|26|10|iudicium determinat causas et qui inponit stulto silentium iras mitigat
PROV|26|11|sicut canis qui revertitur ad vomitum suum sic inprudens qui iterat stultitiam suam
PROV|26|12|vidisti hominem sapientem sibi videri magis illo spem habebit stultus
PROV|26|13|dicit piger leaena in via leo in itineribus
PROV|26|14|sicut ostium vertitur in cardine suo ita piger in lectulo suo
PROV|26|15|abscondit piger manus sub ascellas suas et laborat si ad os suum eas converterit
PROV|26|16|sapientior sibi piger videtur septem viris loquentibus sententias
PROV|26|17|sicut qui adprehendit auribus canem sic qui transit et inpatiens commiscetur rixae alterius
PROV|26|18|sicut noxius est qui mittit lanceas et sagittas et mortem
PROV|26|19|sic vir qui fraudulenter nocet amico suo et cum fuerit deprehensus dicit ludens feci
PROV|26|20|cum defecerint ligna extinguetur ignis et susurrone subtracto iurgia conquiescunt
PROV|26|21|sicut carbones ad prunam et ligna ad ignem sic homo iracundus suscitat rixas
PROV|26|22|verba susurronis quasi simplicia et ipsa perveniunt ad intima ventris
PROV|26|23|quomodo si argento sordido ornare velis vas fictile sic labia tumentia cum pessimo corde sociata
PROV|26|24|labiis suis intellegitur inimicus cum in corde tractaverit dolos
PROV|26|25|quando submiserit vocem suam ne credideris ei quoniam septem nequitiae sunt in corde illius
PROV|26|26|qui operit odium fraudulenter revelabitur malitia eius in concilio
PROV|26|27|qui fodit foveam incidet in eam et qui volvit lapidem revertetur ad eum
PROV|26|28|lingua fallax non amat veritatem et os lubricum operatur ruinas
PROV|27|1|ne glorieris in crastinum ignorans quid superventura pariat dies
PROV|27|2|laudet te alienus et non os tuum extraneus et non labia tua
PROV|27|3|grave est saxum et onerosa harena sed ira stulti utroque gravior
PROV|27|4|ira non habet misericordiam nec erumpens furor et impetum concitati ferre quis poterit
PROV|27|5|melior est manifesta correptio quam amor absconditus
PROV|27|6|meliora sunt vulnera diligentis quam fraudulenta odientis oscula
PROV|27|7|anima saturata calcabit favum anima esuriens et amarum pro dulce sumet
PROV|27|8|sicut avis transmigrans de nido suo sic vir qui relinquit locum suum
PROV|27|9|unguento et variis odoribus delectatur cor et bonis amici consiliis anima dulcoratur
PROV|27|10|amicum tuum et amicum patris tui ne dimiseris et domum fratris tui ne ingrediaris in die adflictionis tuae melior est vicinus iuxta quam frater procul
PROV|27|11|stude sapientiae fili mi et laetifica cor meum ut possim exprobranti respondere sermonem
PROV|27|12|astutus videns malum absconditus est parvuli transeuntes sustinuere dispendia
PROV|27|13|tolle vestimentum eius qui spopondit pro extraneo et pro alienis auferto pignus
PROV|27|14|qui benedicit proximo suo voce grandi de nocte consurgens maledicenti similis erit
PROV|27|15|tecta perstillantia in die frigoris et litigiosa mulier conparantur
PROV|27|16|qui retinet eam quasi qui ventum teneat et oleum dexterae suae vocabit
PROV|27|17|ferrum ferro acuitur et homo exacuit faciem amici sui
PROV|27|18|qui servat ficum comedet fructus eius et qui custos est domini sui glorificabitur
PROV|27|19|quomodo in aquis resplendent vultus prospicientium sic corda hominum manifesta sunt prudentibus
PROV|27|20|infernus et perditio non replentur similiter et oculi hominum insatiabiles
PROV|27|21|quomodo probatur in conflatorio argentum et in fornace aurum sic probatur homo ore laudantis
PROV|27|22|si contuderis stultum in pila quasi tisanas feriente desuper pilo non auferetur ab eo stultitia eius
PROV|27|23|diligenter agnosce vultum pecoris tui tuosque greges considera
PROV|27|24|non enim habebis iugiter potestatem sed corona tribuetur in generatione generationum
PROV|27|25|aperta sunt prata et apparuerunt herbae virentes et collecta sunt faena de montibus
PROV|27|26|agni ad vestimentum tuum et hedi agri pretium
PROV|27|27|sufficiat tibi lac caprarum in cibos tuos in necessaria domus tuae et ad victum ancillis tuis
PROV|28|1|fugit impius nemine persequente iustus autem quasi leo confidens absque terrore erit
PROV|28|2|propter peccata terrae multi principes eius et propter hominis sapientiam et horum scientiam quae dicuntur vita ducis longior erit
PROV|28|3|vir pauper calumnians pauperes similis imbri vehementi in quo paratur fames
PROV|28|4|qui derelinquunt legem laudant impium qui custodiunt succenduntur contra eum
PROV|28|5|viri mali non cogitant iudicium qui autem requirunt Dominum animadvertunt omnia
PROV|28|6|melior est pauper ambulans in simplicitate sua quam dives pravis itineribus
PROV|28|7|qui custodit legem filius sapiens est qui pascit comesatores confundit patrem suum
PROV|28|8|qui coacervat divitias usuris et fenore liberali in pauperes congregat eas
PROV|28|9|qui declinat aurem suam ne audiat legem oratio eius erit execrabilis
PROV|28|10|qui decipit iustos in via mala in interitu suo corruet et simplices possidebunt bona
PROV|28|11|sapiens sibi videtur vir dives pauper autem prudens scrutabitur eum
PROV|28|12|in exultatione iustorum multa gloria regnantibus impiis ruinae hominum
PROV|28|13|qui abscondit scelera sua non dirigetur qui confessus fuerit et reliquerit ea misericordiam consequetur
PROV|28|14|beatus homo qui semper est pavidus qui vero mentis est durae corruet in malum
PROV|28|15|leo rugiens et ursus esuriens princeps impius super populum pauperem
PROV|28|16|dux indigens prudentia multos opprimet per calumniam qui autem odit avaritiam longi fient dies eius
PROV|28|17|hominem qui calumniatur animae sanguinem si usque ad lacum fugerit nemo sustentet
PROV|28|18|qui ambulat simpliciter salvus erit qui perversis ingreditur viis concidet semel
PROV|28|19|qui operatur terram suam saturabitur panibus qui sectatur otium replebitur egestate
PROV|28|20|vir fidelis multum laudabitur qui autem festinat ditari non erit innocens
PROV|28|21|qui cognoscit in iudicio faciem non facit bene iste et pro buccella panis deserit veritatem
PROV|28|22|vir qui festinat ditari et aliis invidet ignorat quod egestas superveniat ei
PROV|28|23|qui corripit hominem gratiam postea inveniet apud eum magis quam ille qui per linguae blandimenta decipit
PROV|28|24|qui subtrahit aliquid a patre suo et matre et dicit hoc non est peccatum particeps homicidae est
PROV|28|25|qui se iactat et dilatat iurgia concitat qui sperat in Domino saginabitur
PROV|28|26|qui confidit in corde suo stultus est qui autem graditur sapienter iste salvabitur
PROV|28|27|qui dat pauperi non indigebit qui despicit deprecantem sustinebit penuriam
PROV|28|28|cum surrexerint impii abscondentur homines cum illi perierint multiplicabuntur iusti
PROV|29|1|viro qui corripientem dura cervice contemnit repentinus superveniet interitus et eum sanitas non sequitur
PROV|29|2|in multiplicatione iustorum laetabitur vulgus cum impii sumpserint principatum gemet populus
PROV|29|3|vir qui amat sapientiam laetificat patrem suum qui autem nutrit scorta perdet substantiam
PROV|29|4|rex iustus erigit terram vir avarus destruet eam
PROV|29|5|homo qui blandis fictisque sermonibus loquitur amico suo rete expandit gressibus eius
PROV|29|6|peccantem virum iniquum involvet laqueus et iustus laudabit atque gaudebit
PROV|29|7|novit iustus causam pauperum impius ignorat scientiam
PROV|29|8|homines pestilentes dissipant civitatem sapientes avertunt furorem
PROV|29|9|vir sapiens si cum stulto contenderit sive irascatur sive rideat non inveniet requiem
PROV|29|10|viri sanguinum oderunt simplicem iusti quaerunt animam eius
PROV|29|11|totum spiritum suum profert stultus sapiens differt et reservat in posterum
PROV|29|12|princeps qui libenter audit verba mendacii omnes ministros habebit impios
PROV|29|13|pauper et creditor obviam fuerunt sibi utriusque inluminator est Dominus
PROV|29|14|rex qui iudicat in veritate pauperes thronus eius in aeternum firmabitur
PROV|29|15|virga atque correptio tribuet sapientiam puer autem qui dimittitur voluntati suae confundet matrem suam
PROV|29|16|in multiplicatione impiorum multiplicabuntur scelera et iusti ruinas eorum videbunt
PROV|29|17|erudi filium tuum et refrigerabit te et dabit delicias animae tuae
PROV|29|18|cum prophetia defecerit dissipabitur populus qui custodit legem beatus est
PROV|29|19|servus verbis non potest erudiri quia quod dicis intellegit et respondere contemnit
PROV|29|20|vidisti hominem velocem ad loquendum stulti magis speranda est quam illius correptio
PROV|29|21|qui delicate a pueritia nutrit servum suum postea illum sentiet contumacem
PROV|29|22|vir iracundus provocat rixas et qui ad indignandum facilis est erit ad peccata proclivior
PROV|29|23|superbum sequitur humilitas et humilem spiritu suscipiet gloria
PROV|29|24|qui cum fure partitur odit animam suam adiurantem audit et non indicat
PROV|29|25|qui timet hominem cito corruet qui sperat in Domino sublevabitur
PROV|29|26|multi requirunt faciem principis et a Domino iudicium egreditur singulorum
PROV|29|27|abominantur iusti virum impium et abominantur impii eos qui in recta sunt via
PROV|30|1|verba Congregantis filii Vomentis visio quam locutus est vir cum quo est Deus et qui Deo secum morante confortatus ait
PROV|30|2|stultissimus sum virorum et sapientia hominum non est mecum
PROV|30|3|non didici sapientiam et non novi sanctorum scientiam
PROV|30|4|quis ascendit in caelum atque descendit quis continuit spiritum manibus suis quis conligavit aquas quasi in vestimento quis suscitavit omnes terminos terrae quod nomen eius et quod nomen filii eius si nosti
PROV|30|5|omnis sermo Dei ignitus clypeus est sperantibus in se
PROV|30|6|ne addas quicquam verbis illius et arguaris inveniarisque mendax
PROV|30|7|duo rogavi te ne deneges mihi antequam moriar
PROV|30|8|vanitatem et verba mendacia longe fac a me mendicitatem et divitias ne dederis mihi tribue tantum victui meo necessaria
PROV|30|9|ne forte saturatus inliciar ad negandum et dicam quis est Dominus et egestate conpulsus furer et peierem nomen Dei mei
PROV|30|10|ne accuses servum ad dominum suum ne forte maledicat tibi et corruas
PROV|30|11|generatio quae patri suo maledicit et quae non benedicit matri suae
PROV|30|12|generatio quae sibi munda videtur et tamen non est lota a sordibus suis
PROV|30|13|generatio cuius excelsi sunt oculi et palpebrae eius in alta subrectae
PROV|30|14|generatio quae pro dentibus gladios habet et commandit molaribus suis ut comedat inopes de terra et pauperes ex hominibus
PROV|30|15|sanguisugae duae sunt filiae dicentes adfer adfer tria sunt insaturabilia et quartum quod numquam dicit sufficit
PROV|30|16|infernus et os vulvae et terra quae non satiatur aqua ignis vero numquam dicit sufficit
PROV|30|17|oculum qui subsannat patrem et qui despicit partum matris suae effodiant corvi de torrentibus et comedant illum filii aquilae
PROV|30|18|tria sunt difficilia mihi et quartum penitus ignoro
PROV|30|19|viam aquilae in caelo viam colubri super petram viam navis in medio mari et viam viri in adulescentula
PROV|30|20|talis est via mulieris adulterae quae comedit et tergens os suum dicit non sum operata malum
PROV|30|21|per tria movetur terra et quartum non potest sustinere
PROV|30|22|per servum cum regnaverit per stultum cum saturatus fuerit cibo
PROV|30|23|per odiosam mulierem cum in matrimonio fuerit adsumpta et per ancillam cum heres fuerit dominae suae
PROV|30|24|quattuor sunt minima terrae et ipsa sunt sapientiora sapientibus
PROV|30|25|formicae populus infirmus quae praeparant in messe cibum sibi
PROV|30|26|lepusculus plebs invalida quae conlocat in petra cubile suum
PROV|30|27|regem lucusta non habet et egreditur universa per turmas
PROV|30|28|stilio manibus nititur et moratur in aedibus regis
PROV|30|29|tria sunt quae bene gradiuntur et quartum quod incedit feliciter
PROV|30|30|leo fortissimus bestiarum ad nullius pavebit occursum
PROV|30|31|gallus succinctus lumbos et aries nec est rex qui resistat ei
PROV|30|32|et qui stultus apparuit postquam elatus est in sublime si enim intellexisset ori inposuisset manum
PROV|30|33|qui autem fortiter premit ubera ad eliciendum lac exprimit butyrum et qui vehementer emungitur elicit sanguinem et qui provocat iras producit discordias
PROV|31|1|verba Lamuhel regis visio qua erudivit eum mater sua
PROV|31|2|quid dilecte mi quid dilecte uteri mei quid dilecte votorum meorum
PROV|31|3|ne dederis mulieribus substantiam tuam et vias tuas ad delendos reges
PROV|31|4|noli regibus o Lamuhel noli regibus dare vinum quia nullum secretum est ubi regnat ebrietas
PROV|31|5|ne forte bibat et obliviscatur iudiciorum et mutet causam filiorum pauperis
PROV|31|6|date siceram maerentibus et vinum his qui amaro sunt animo
PROV|31|7|bibant ut obliviscantur egestatis suae et doloris non recordentur amplius
PROV|31|8|aperi os tuum muto et causis omnium filiorum qui pertranseunt
PROV|31|9|aperi os tuum decerne quod iustum est et iudica inopem et pauperem
PROV|31|10|aleph mulierem fortem quis inveniet procul et de ultimis finibus pretium eius
PROV|31|11|beth confidit in ea cor viri sui et spoliis non indigebit
PROV|31|12|gimel reddet ei bonum et non malum omnibus diebus vitae suae
PROV|31|13|deleth quaesivit lanam et linum et operata est consilio manuum suarum
PROV|31|14|he facta est quasi navis institoris de longe portat panem suum
PROV|31|15|vav et de nocte surrexit deditque praedam domesticis suis et cibaria ancillis suis
PROV|31|16|zai consideravit agrum et emit eum de fructu manuum suarum plantavit vineam
PROV|31|17|heth accinxit fortitudine lumbos suos et roboravit brachium suum
PROV|31|18|teth gustavit quia bona est negotiatio eius non extinguetur in nocte lucerna illius
PROV|31|19|ioth manum suam misit ad fortia et digiti eius adprehenderunt fusum
PROV|31|20|caph manum suam aperuit inopi et palmas suas extendit ad pauperem
PROV|31|21|lameth non timebit domui suae a frigoribus nivis omnes enim domestici eius vestiti duplicibus
PROV|31|22|mem stragulam vestem fecit sibi byssus et purpura indumentum eius
PROV|31|23|nun nobilis in portis vir eius quando sederit cum senatoribus terrae
PROV|31|24|samech sindonem fecit et vendidit et cingulum tradidit Chananeo
PROV|31|25|ain fortitudo et decor indumentum eius et ridebit in die novissimo
PROV|31|26|phe os suum aperuit sapientiae et lex clementiae in lingua eius
PROV|31|27|sade considerat semitas domus suae et panem otiosa non comedet
PROV|31|28|coph surrexerunt filii eius et beatissimam praedicaverunt vir eius et laudavit eam
PROV|31|29|res multae filiae congregaverunt divitias tu supergressa es universas
PROV|31|30|sin fallax gratia et vana est pulchritudo mulier timens Dominum ipsa laudabitur
PROV|31|31|thau date ei de fructu manuum suarum et laudent eam in portis opera eius
ECCL|1|1|verba Ecclesiastes filii David regis Hierusalem
ECCL|1|2|vanitas vanitatum dixit Ecclesiastes vanitas vanitatum omnia vanitas
ECCL|1|3|quid habet amplius homo de universo labore suo quod laborat sub sole
ECCL|1|4|generatio praeterit et generatio advenit terra vero in aeternum stat
ECCL|1|5|oritur sol et occidit et ad locum suum revertitur ibique renascens
ECCL|1|6|gyrat per meridiem et flectitur ad aquilonem lustrans universa circuitu pergit spiritus et in circulos suos regreditur
ECCL|1|7|omnia flumina intrant mare et mare non redundat ad locum unde exeunt flumina revertuntur ut iterum fluant
ECCL|1|8|cunctae res difficiles non potest eas homo explicare sermone non saturatur oculus visu nec auris impletur auditu
ECCL|1|9|quid est quod fuit ipsum quod futurum est quid est quod factum est ipsum quod fiendum est
ECCL|1|10|nihil sub sole novum nec valet quisquam dicere ecce hoc recens est iam enim praecessit in saeculis quae fuerunt ante nos
ECCL|1|11|non est priorum memoria sed nec eorum quidem quae postea futura sunt erit recordatio apud eos qui futuri sunt in novissimo
ECCL|1|12|ego Ecclesiastes fui rex Israhel in Hierusalem
ECCL|1|13|et proposui in animo meo quaerere et investigare sapienter de omnibus quae fiunt sub sole hanc occupationem pessimam dedit Deus filiis hominum ut occuparentur in ea
ECCL|1|14|vidi quae fiunt cuncta sub sole et ecce universa vanitas et adflictio spiritus
ECCL|1|15|perversi difficile corriguntur et stultorum infinitus est numerus
ECCL|1|16|locutus sum in corde meo dicens ecce magnus effectus sum et praecessi sapientia omnes qui fuerunt ante me in Hierusalem et mens mea contemplata est multa sapienter et didicit
ECCL|1|17|dedique cor meum ut scirem prudentiam atque doctrinam erroresque et stultitiam et agnovi quod in his quoque esset labor et adflictio spiritus
ECCL|1|18|eo quod in multa sapientia multa sit indignatio et qui addit scientiam addat et laborem
ECCL|2|1|dixi ego in corde meo vadam et affluam deliciis et fruar bonis et vidi quod hoc quoque esset vanitas
ECCL|2|2|risum reputavi errorem et gaudio dixi quid frustra deciperis
ECCL|2|3|cogitavi in corde meo abstrahere a vino carnem meam ut animum meum transferrem ad sapientiam devitaremque stultitiam donec viderem quid esset utile filiis hominum quod facto opus est sub sole numero dierum vitae suae
ECCL|2|4|magnificavi opera mea aedificavi mihi domos plantavi vineas
ECCL|2|5|feci hortos et pomeria et consevi ea cuncti generis arboribus
ECCL|2|6|extruxi mihi piscinas aquarum ut inrigarem silvam lignorum germinantium
ECCL|2|7|possedi servos et ancillas multamque familiam habui armenta quoque et magnos ovium greges ultra omnes qui fuerunt ante me in Hierusalem
ECCL|2|8|coacervavi mihi argentum et aurum et substantias regum ac provinciarum feci mihi cantores et cantrices et delicias filiorum hominum scyphos et urceos in ministerio ad vina fundenda
ECCL|2|9|et supergressus sum opibus omnes qui fuerunt ante me in Hierusalem sapientia quoque perseveravit mecum
ECCL|2|10|et omnia quae desideraverunt oculi mei non negavi eis nec prohibui cor quin omni voluptate frueretur et oblectaret se in his quae paraveram et hanc ratus sum partem meam si uterer labore meo
ECCL|2|11|cumque me convertissem ad universa opera quae fecerant manus meae et ad labores in quibus frustra sudaveram vidi in omnibus vanitatem et adflictionem animi et nihil permanere sub sole
ECCL|2|12|transivi ad contemplandam sapientiam erroresque et stultitiam quid est inquam homo ut sequi possit regem factorem suum
ECCL|2|13|et vidi quia tantum praecederet sapientia stultitiam quantum differt lux tenebris
ECCL|2|14|sapientis oculi in capite eius stultus in tenebris ambulat et didici quod unus utriusque esset interitus
ECCL|2|15|et dixi in corde meo si unus et stulti et meus occasus erit quid mihi prodest quod maiorem sapientiae dedi operam locutusque cum mente mea animadverti quod hoc quoque esset vanitas
ECCL|2|16|non enim erit memoria sapientis similiter ut stulti in perpetuum et futura tempora oblivione cuncta pariter obruent moritur doctus similiter et indoctus
ECCL|2|17|et idcirco taeduit me vitae meae videntem mala esse universa sub sole et cuncta vanitatem atque adflictionem spiritus
ECCL|2|18|rursum detestatus sum omnem industriam meam quae sub sole studiosissime laboravi habiturus heredem post me
ECCL|2|19|quem ignoro utrum sapiens an stultus futurus sit et dominabitur in laboribus meis quibus desudavi et sollicitus fui et est quicquam tam vanum
ECCL|2|20|unde cessavi renuntiavitque cor meum ultra laborare sub sole
ECCL|2|21|nam cum alius laboret in sapientia et doctrina et sollicitudine homini otioso quaesita dimittit et hoc ergo vanitas et magnum malum
ECCL|2|22|quid enim proderit homini de universo labore suo et adflictione spiritus qua sub sole cruciatus est
ECCL|2|23|cuncti dies eius doloribus et aerumnis pleni sunt nec per noctem mente requiescit et haec non vanitas est
ECCL|2|24|nonne melius est comedere et bibere et ostendere animae suae bona de laboribus suis et hoc de manu Dei est
ECCL|2|25|quis ita vorabit et deliciis affluet ut ego
ECCL|2|26|homini bono in conspectu suo dedit Deus sapientiam et scientiam et laetitiam peccatori autem dedit adflictionem et curam superfluam ut addat et congreget et tradat ei qui placuit Deo sed et hoc vanitas et cassa sollicitudo mentis
ECCL|3|1|omnia tempus habent et suis spatiis transeunt universa sub caelo
ECCL|3|2|tempus nascendi et tempus moriendi tempus plantandi et tempus evellendi quod plantatum est
ECCL|3|3|tempus occidendi et tempus sanandi tempus destruendi et tempus aedificandi
ECCL|3|4|tempus flendi et tempus ridendi tempus plangendi et tempus saltandi
ECCL|3|5|tempus spargendi lapides et tempus colligendi tempus amplexandi et tempus longe fieri a conplexibus
ECCL|3|6|tempus adquirendi et tempus perdendi tempus custodiendi et tempus abiciendi
ECCL|3|7|tempus scindendi et tempus consuendi tempus tacendi et tempus loquendi
ECCL|3|8|tempus dilectionis et tempus odii tempus belli et tempus pacis
ECCL|3|9|quid habet amplius homo de labore suo
ECCL|3|10|vidi adflictionem quam dedit Deus filiis hominum ut distendantur in ea
ECCL|3|11|cuncta fecit bona in tempore suo et mundum tradidit disputationi eorum ut non inveniat homo opus quod operatus est Deus ab initio usque ad finem
ECCL|3|12|et cognovi quod non esset melius nisi laetari et facere bene in vita sua
ECCL|3|13|omnis enim homo qui comedit et bibit et videt bonum de labore suo hoc donum Dei est
ECCL|3|14|didici quod omnia opera quae fecit Deus perseverent in perpetuum non possumus eis quicquam addere nec auferre quae fecit Deus ut timeatur
ECCL|3|15|quod factum est ipsum permanet quae futura sunt iam fuerunt et Deus instaurat quod abiit
ECCL|3|16|vidi sub sole in loco iudicii impietatem et in loco iustitiae iniquitatem
ECCL|3|17|et dixi in corde meo iustum et impium iudicabit Deus et tempus omni rei tunc erit
ECCL|3|18|dixi in corde meo de filiis hominum ut probaret eos Deus et ostenderet similes esse bestiis
ECCL|3|19|idcirco unus interitus est hominis et iumentorum et aequa utriusque condicio sicut moritur homo sic et illa moriuntur similiter spirant omnia et nihil habet homo iumento amplius cuncta subiacent vanitati
ECCL|3|20|et omnia pergunt ad unum locum de terra facta sunt et in terram pariter revertentur
ECCL|3|21|quis novit si spiritus filiorum Adam ascendat sursum et si spiritus iumentorum descendat deorsum
ECCL|3|22|et deprehendi nihil esse melius quam laetari hominem in opere suo et hanc esse partem illius quis enim eum adducet ut post se futura cognoscat
ECCL|4|1|verti me ad alia et vidi calumnias quae sub sole geruntur et lacrimas innocentum et consolatorem neminem nec posse resistere eorum violentiae cunctorum auxilio destitutos
ECCL|4|2|et laudavi magis mortuos quam viventes
ECCL|4|3|et feliciorem utroque iudicavi qui necdum natus est nec vidit mala quae sub sole fiunt
ECCL|4|4|rursum contemplatus omnes labores hominum et industrias animadverti patere invidiae proximi et in hoc ergo vanitas et cura superflua est
ECCL|4|5|stultus conplicat manus suas et comedit carnes suas dicens
ECCL|4|6|melior est pugillus cum requie quam plena utraque manus cum labore et adflictione animi
ECCL|4|7|considerans repperi et aliam vanitatem sub sole
ECCL|4|8|unus est et secundum non habet non filium non fratrem et tamen laborare non cessat nec satiantur oculi eius divitiis nec recogitat dicens cui laboro et fraudo animam meam bonis in hoc quoque vanitas est et adflictio pessima
ECCL|4|9|melius ergo est duos simul esse quam unum habent enim emolumentum societatis suae
ECCL|4|10|si unus ceciderit ab altero fulcietur vae soli quia cum ruerit non habet sublevantem
ECCL|4|11|et si dormierint duo fovebuntur mutuo unus quomodo calefiet
ECCL|4|12|et si quispiam praevaluerit contra unum duo resistent ei funiculus triplex difficile rumpitur
ECCL|4|13|melior est puer pauper et sapiens rege sene et stulto qui nescit providere in posterum
ECCL|4|14|quod et de carcere catenisque interdum quis egrediatur ad regnum et alius natus in regno inopia consumatur
ECCL|4|15|vidi cunctos viventes qui ambulant sub sole cum adulescente secundo qui consurgit pro eo
ECCL|4|16|infinitus numerus est populi omnium qui fuerunt ante eum et qui postea futuri sunt non laetabuntur in eo sed et hoc vanitas et adflictio spiritus
ECCL|4|17|custodi pedem tuum ingrediens domum Dei multo enim melior est oboedientia quam stultorum victimae qui nesciunt quid faciant mali
ECCL|5|1|ne temere quid loquaris neque cor tuum sit velox ad proferendum sermonem coram Deo Deus enim in caelo et tu super terram idcirco sint pauci sermones tui
ECCL|5|2|multas curas sequuntur somnia et in multis sermonibus invenitur stultitia
ECCL|5|3|si quid vovisti Deo ne moreris reddere displicet enim ei infidelis et stulta promissio sed quodcumque voveris redde
ECCL|5|4|multoque melius est non vovere quam post votum promissa non conplere
ECCL|5|5|ne dederis os tuum ut peccare faciat carnem tuam neque dicas coram angelo non est providentia ne forte iratus Deus super sermone tuo dissipet cuncta opera manuum tuarum
ECCL|5|6|ubi multa sunt somnia plurimae vanitates et sermones innumeri tu vero Deum time
ECCL|5|7|si videris calumnias egenorum et violenta iudicia et subverti iustitiam in provincia non mireris super hoc negotio quia excelso alius excelsior est et super hos quoque eminentiores sunt alii
ECCL|5|8|et insuper universae terrae rex imperat servienti
ECCL|5|9|avarus non implebitur pecunia et qui amat divitias fructus non capiet ex eis et hoc ergo vanitas
ECCL|5|10|ubi multae sunt opes multi et qui comedant eas et quid prodest possessori nisi quod cernit divitias oculis suis
ECCL|5|11|dulcis est somnus operanti sive parum sive multum comedat saturitas autem divitis non sinit dormire eum
ECCL|5|12|est et alia infirmitas pessima quam vidi sub sole divitiae conservatae in malum domini sui
ECCL|5|13|pereunt enim in adflictione pessima generavit filium qui in summa egestate erit
ECCL|5|14|sicut egressus est nudus de utero matris suae sic revertetur et nihil auferet secum de labore suo
ECCL|5|15|miserabilis prorsus infirmitas quomodo venit sic revertetur quid ergo prodest ei quod laboravit in ventum
ECCL|5|16|cunctis diebus vitae suae comedit in tenebris et in curis multis et in aerumna atque tristitia
ECCL|5|17|hoc itaque mihi visum est bonum ut comedat quis et bibat et fruatur laetitia ex labore suo quod laboravit ipse sub sole numerum dierum vitae suae quos dedit ei Deus et haec est pars illius
ECCL|5|18|et omni homini cui dedit Deus divitias atque substantiam potestatemque ei tribuit ut comedat ex eis et fruatur parte sua et laetetur de labore suo hoc est donum Dei
ECCL|5|19|non enim satis recordabitur dierum vitae suae eo quod Deus occupet deliciis cor eius
ECCL|6|1|est et aliud malum quod vidi sub sole et quidem frequens apud homines
ECCL|6|2|vir cui dedit Deus divitias et substantiam et honorem et nihil deest animae eius ex omnibus quae desiderat nec tribuit ei potestatem Deus ut comedat ex eo sed homo extraneus vorabit illud hoc vanitas et magna miseria est
ECCL|6|3|si genuerit quispiam centum et vixerit multos annos et plures dies aetatis habuerit et anima illius non utatur bonis substantiae suae sepulturaque careat de hoc ego pronuntio quod melior illo sit abortivus
ECCL|6|4|frustra enim venit et pergit ad tenebras et oblivione delebitur nomen eius
ECCL|6|5|non vidit solem neque cognovit distantiam boni et mali
ECCL|6|6|etiam si duobus milibus annis vixerit et non fuerit perfruitus bonis nonne ad unum locum properant omnia
ECCL|6|7|omnis labor hominis in ore eius sed anima illius non impletur
ECCL|6|8|quid habet amplius sapiens ab stulto et quid pauper nisi ut pergat illuc ubi est vita
ECCL|6|9|melius est videre quod cupias quam desiderare quod nescias sed et hoc vanitas est et praesumptio spiritus
ECCL|6|10|qui futurus est iam vocatum est nomen eius et scitur quod homo sit et non possit contra fortiorem se in iudicio contendere
ECCL|6|11|verba sunt plurima multa in disputando habentia vanitatem
ECCL|7|1|quid necesse est homini maiora se quaerere cum ignoret quid conducat sibi in vita sua numero dierum peregrinationis suae et tempore quo velut umbra praeterit aut quis ei poterit indicare quid post eum futurum sub sole sit
ECCL|7|2|melius est nomen bonum quam unguenta pretiosa et dies mortis die nativitatis
ECCL|7|3|melius est ire ad domum luctus quam ad domum convivii in illa enim finis cunctorum admonetur hominum et vivens cogitat quid futurum sit
ECCL|7|4|melior est ira risu quia per tristitiam vultus corrigitur animus delinquentis
ECCL|7|5|cor sapientium ubi tristitia est et cor stultorum ubi laetitia
ECCL|7|6|melius est a sapiente corripi quam stultorum adulatione decipi
ECCL|7|7|quia sicut sonitus spinarum ardentium sub olla sic risus stulti sed et hoc vanitas
ECCL|7|8|calumnia conturbat sapientem et perdet robur cordis illius
ECCL|7|9|melior est finis orationis quam principium melior est patiens arrogante
ECCL|7|10|ne velox sis ad irascendum quia ira in sinu stulti requiescit
ECCL|7|11|ne dicas quid putas causae est quod priora tempora meliora fuere quam nunc sunt stulta est enim huiuscemodi interrogatio
ECCL|7|12|utilior est sapientia cum divitiis et magis prodest videntibus solem
ECCL|7|13|sicut enim protegit sapientia sic protegit pecunia hoc autem plus habet eruditio et sapientia quod vitam tribuunt possessori suo
ECCL|7|14|considera opera Dei quod nemo possit corrigere quem ille despexerit
ECCL|7|15|in die bona fruere bonis et malam diem praecave sicut enim hanc sic et illam fecit Deus ut non inveniat homo contra eum iustas querimonias
ECCL|7|16|haec quoque vidi in diebus vanitatis meae iustus perit in iustitia sua et impius multo vivit tempore in malitia sua
ECCL|7|17|noli esse iustus multum neque plus sapias quam necesse est ne obstupescas
ECCL|7|18|ne impie agas multum et noli esse stultus ne moriaris in tempore non tuo
ECCL|7|19|bonum est te sustentare iustum sed et ab illo ne subtrahas manum tuam quia qui Deum timet nihil neglegit
ECCL|7|20|sapientia confortabit sapientem super decem principes civitatis
ECCL|7|21|non est enim homo iustus in terra qui faciat bonum et non peccet
ECCL|7|22|sed et cunctis sermonibus qui dicuntur ne accommodes cor tuum ne forte audias servum tuum maledicentem tibi
ECCL|7|23|scit enim tua conscientia quia et tu crebro maledixisti aliis
ECCL|7|24|cuncta temptavi in sapientia dixi sapiens efficiar et ipsa longius recessit a me
ECCL|7|25|multo magis quam erat et alta profunditas quis inveniet eam
ECCL|7|26|lustravi universa animo meo ut scirem et considerarem et quaererem sapientiam et rationem et ut cognoscerem impietatem stulti et errorem inprudentium
ECCL|7|27|et inveni amariorem morte mulierem quae laqueus venatorum est et sagena cor eius vincula sunt manus illius qui placet Deo effugiet eam qui autem peccator est capietur ab illa
ECCL|7|28|ecce hoc inveni dicit Ecclesiastes unum et alterum ut invenirem rationem
ECCL|7|29|quam adhuc quaerit anima mea et non inveni virum de mille unum repperi mulierem ex omnibus non inveni
ECCL|7|30|solummodo hoc inveni quod fecerit Deus hominem rectum et ipse se infinitis miscuerit quaestionibus quis talis ut sapiens est et quis cognovit solutionem verbi
ECCL|8|1|sapientia hominis lucet in vultu eius et potentissimus faciem illius commutavit
ECCL|8|2|ego os regis observo et praecepta iuramenti Dei
ECCL|8|3|ne festines recedere a facie eius neque permaneas in opere malo quia omne quod voluerit faciet
ECCL|8|4|et sermo illius potestate plenus est nec dicere ei quisquam potest quare ita facis
ECCL|8|5|qui custodit praeceptum non experietur quicquam mali tempus et responsionem cor sapientis intellegit
ECCL|8|6|omni negotio tempus est et oportunitas et multa hominis adflictio
ECCL|8|7|quia ignorat praeterita et ventura nullo scire potest nuntio
ECCL|8|8|non est in hominis dicione prohibere spiritum nec habet potestatem in die mortis nec sinitur quiescere ingruente bello neque salvabit impietas impium
ECCL|8|9|omnia haec consideravi et dedi cor meum in cunctis operibus quae fiunt sub sole interdum dominatur homo homini in malum suum
ECCL|8|10|vidi impios sepultos qui etiam cum adviverent in loco sancto erant et laudabantur in civitate quasi iustorum operum sed et hoc vanitas est
ECCL|8|11|etenim quia non profertur cito contra malos sententia absque ullo timore filii hominum perpetrant mala
ECCL|8|12|attamen ex eo quod peccator centies facit malum et per patientiam sustentatur ego cognovi quod erit bonum timentibus Deum qui verentur faciem eius
ECCL|8|13|non sit bonum impio nec prolongentur dies eius sed quasi umbra transeant qui non timent faciem Dei
ECCL|8|14|est et alia vanitas quae fit super terram sunt iusti quibus multa proveniunt quasi opera egerint impiorum et sunt impii qui ita securi sunt quasi iustorum facta habeant sed et hoc vanissimum iudico
ECCL|8|15|laudavi igitur laetitiam quod non esset homini bonum sub sole nisi quod comederet et biberet atque gauderet et hoc solum secum auferret de labore suo in diebus vitae quos dedit ei Deus sub sole
ECCL|8|16|et adposui cor meum ut scirem sapientiam et intellegerem distentionem quae versatur in terra est homo qui diebus ac noctibus somnum oculis non capit
ECCL|8|17|et intellexi quod omnium operum Dei nullam possit homo invenire rationem eorum quae fiunt sub sole et quanto plus laboraverit ad quaerendum tanto minus inveniat etiam si dixerit sapiens se nosse non poterit repperire
ECCL|9|1|omnia haec tractavi in corde meo ut curiose intellegerem sunt iusti atque sapientes et opera eorum in manu Dei et tamen nescit homo utrum amore an odio dignus sit
ECCL|9|2|sed omnia in futuro servantur incerta eo quod universa aeque eveniant iusto et impio bono et malo mundo et inmundo immolanti victimas et sacrificia contemnenti sicut bonus sic et peccator ut periurus ita et ille qui verum deierat
ECCL|9|3|hoc est pessimum inter omnia quae sub sole fiunt quia eadem cunctis eveniunt unde et corda filiorum hominum implentur malitia et contemptu in vita sua et post haec ad inferos deducentur
ECCL|9|4|nemo est qui semper vivat et qui huius rei habeat fiduciam melior est canis vivens leone mortuo
ECCL|9|5|viventes enim sciunt se esse morituros mortui vero nihil noverunt amplius nec habent ultra mercedem quia oblivioni tradita est memoria eorum
ECCL|9|6|amor quoque et odium et invidia simul perierunt nec habent partem in hoc saeculo et in opere quod sub sole geritur
ECCL|9|7|vade ergo et comede in laetitia panem tuum et bibe cum gaudio vinum tuum quia Deo placent opera tua
ECCL|9|8|omni tempore sint vestimenta tua candida et oleum de capite tuo non deficiat
ECCL|9|9|perfruere vita cum uxore quam diligis cunctis diebus vitae instabilitatis tuae qui dati sunt tibi sub sole omni tempore vanitatis tuae haec est enim pars in vita et in labore tuo quod laboras sub sole
ECCL|9|10|quodcumque potest manus tua facere instanter operare quia nec opus nec ratio nec scientia nec sapientia erunt apud inferos quo tu properas
ECCL|9|11|verti me alio vidique sub sole nec velocium esse cursum nec fortium bellum nec sapientium panem nec doctorum divitias nec artificum gratiam sed tempus casumque in omnibus
ECCL|9|12|nescit homo finem suum sed sicut pisces capiuntur hamo et sicut aves conprehenduntur laqueo sic capiuntur homines tempore malo cum eis extemplo supervenerit
ECCL|9|13|hanc quoque vidi sub sole sapientiam et probavi maximam
ECCL|9|14|civitas parva et pauci in ea viri venit contra eam rex magnus et vallavit eam extruxitque munitiones per gyrum et perfecta est obsidio
ECCL|9|15|inventusque in ea vir pauper et sapiens liberavit urbem per sapientiam suam et nullus deinceps recordatus est hominis illius pauperis
ECCL|9|16|et dicebam ego meliorem esse sapientiam fortitudine quomodo ergo sapientia pauperis contempta est et verba eius non sunt audita
ECCL|9|17|verba sapientium audiuntur in silentio plus quam clamor principis inter stultos
ECCL|9|18|melior est sapientia quam arma bellica et qui in uno peccaverit multa bona perdet
ECCL|10|1|muscae morientes perdunt suavitatem unguenti pretiosior est sapientia et gloria parva ad tempus stultitia
ECCL|10|2|cor sapientis in dextera eius et cor stulti in sinistra illius
ECCL|10|3|sed et in via stultus ambulans cum ipse insipiens sit omnes stultos aestimat
ECCL|10|4|si spiritus potestatem habentis ascenderit super te locum tuum ne dimiseris quia curatio cessare faciet peccata maxima
ECCL|10|5|est malum quod vidi sub sole quasi per errorem egrediens a facie principis
ECCL|10|6|positum stultum in dignitate sublimi et divites sedere deorsum
ECCL|10|7|vidi servos in equis et principes ambulantes quasi servos super terram
ECCL|10|8|qui fodit foveam incidet in eam et qui dissipat sepem mordebit eum coluber
ECCL|10|9|qui transfert lapides adfligetur in eis et qui scindit ligna vulnerabitur ab eis
ECCL|10|10|si retunsum fuerit ferrum et hoc non ut prius sed hebetatum erit multo labore exacuatur et post industriam sequitur sapientia
ECCL|10|11|si mordeat serpens in silentio nihil eo minus habet qui occulte detrahit
ECCL|10|12|verba oris sapientis gratia et labia insipientis praecipitabunt eum
ECCL|10|13|initium verborum eius stultitia et novissimum oris illius error pessimus
ECCL|10|14|stultus verba multiplicat ignorat homo quid ante se fuerit et quod post futurum est quis illi poterit indicare
ECCL|10|15|labor stultorum adfliget eos qui nesciunt in urbem pergere
ECCL|10|16|vae tibi terra cuius rex est puer et cuius principes mane comedunt
ECCL|10|17|beata terra cuius rex nobilis est et cuius principes vescuntur in tempore suo ad reficiendum et non ad luxuriam
ECCL|10|18|in pigritiis humiliabitur contignatio et in infirmitate manuum perstillabit domus
ECCL|10|19|in risu faciunt panem ac vinum ut epulentur viventes et pecuniae oboedient omnia
ECCL|10|20|in cogitatione tua regi ne detrahas et in secreto cubiculi tui ne maledixeris diviti quia avis caeli portabit vocem tuam et qui habet pinnas adnuntiabit sententiam
ECCL|11|1|mitte panem tuum super transeuntes aquas quia post multa tempora invenies illum
ECCL|11|2|da partem septem necnon et octo quia ignoras quid futurum sit mali super terram
ECCL|11|3|si repletae fuerint nubes imbrem super terram effundent si ceciderit lignum ad austrum aut ad aquilonem in quocumque loco ceciderit ibi erit
ECCL|11|4|qui observat ventum non seminat et qui considerat nubes numquam metet
ECCL|11|5|quomodo ignoras quae sit via spiritus et qua ratione conpingantur ossa in ventre praegnatis sic nescis opera Dei qui fabricator est omnium
ECCL|11|6|mane semina sementem tuam et vespere ne cesset manus tua quia nescis quid magis oriatur hoc an illud et si utrumque simul melius erit
ECCL|11|7|dulce lumen et delectabile est oculis videre solem
ECCL|11|8|si annis multis vixerit homo et in omnibus his laetatus fuerit meminisse debet tenebrosi temporis et dierum multorum qui cum venerint vanitatis arguentur praeterita
ECCL|11|9|laetare ergo iuvenis in adulescentia tua et in bono sit cor tuum in diebus iuventutis tuae et ambula in viis cordis tui et in intuitu oculorum tuorum et scito quod pro omnibus his adducet te Deus in iudicium
ECCL|11|10|aufer iram a corde tuo et amove malitiam a carne tua adulescentia enim et voluptas vana sunt
ECCL|12|1|memento creatoris tui in diebus iuventutis tuae antequam veniat tempus adflictionis et adpropinquent anni de quibus dicas non mihi placent
ECCL|12|2|antequam tenebrescat sol et lumen et luna et stellae et revertantur nubes post pluviam
ECCL|12|3|quando commovebuntur custodes domus et nutabuntur viri fortissimi et otiosae erunt molentes inminuto numero et tenebrescent videntes per foramina
ECCL|12|4|et claudent ostia in platea in humilitate vocis molentis et consurgent ad vocem volucris et obsurdescent omnes filiae carminis
ECCL|12|5|excelsa quoque timebunt et formidabunt in via florebit amigdalum inpinguabitur lucusta et dissipabitur capparis quoniam ibit homo in domum aeternitatis suae et circumibunt in platea plangentes
ECCL|12|6|antequam rumpatur funis argenteus et recurrat vitta aurea et conteratur hydria super fontem et confringatur rota super cisternam
ECCL|12|7|et revertatur pulvis in terram suam unde erat et spiritus redeat ad Deum qui dedit illum
ECCL|12|8|vanitas vanitatum dixit Ecclesiastes omnia vanitas
ECCL|12|9|cumque esset sapientissimus Ecclesiastes docuit populum et enarravit quae fecerit et investigans conposuit parabolas multas
ECCL|12|10|quaesivit verba utilia et conscripsit sermones rectissimos ac veritate plenos
ECCL|12|11|verba sapientium sicut stimuli et quasi clavi in altum defixi quae per magistrorum concilium data sunt a pastore uno
ECCL|12|12|his amplius fili mi ne requiras faciendi plures libros nullus est finis frequensque meditatio carnis adflictio est
ECCL|12|13|finem loquendi omnes pariter audiamus Deum time et mandata eius observa hoc est enim omnis homo
ECCL|12|14|et cuncta quae fiunt adducet Deus in iudicium pro omni errato sive bonum sive malum sit
SONG|1|1|osculetur me osculo oris sui quia meliora sunt ubera tua vino
SONG|1|2|fraglantia unguentis optimis oleum effusum nomen tuum ideo adulescentulae dilexerunt te
SONG|1|3|trahe me post te curremus introduxit me rex in cellaria sua exultabimus et laetabimur in te memores uberum tuorum super vinum recti diligunt te
SONG|1|4|nigra sum sed formonsa filiae Hierusalem sicut tabernacula Cedar sicut pelles Salomonis
SONG|1|5|nolite me considerare quod fusca sim quia decoloravit me sol filii matris meae pugnaverunt contra me posuerunt me custodem in vineis vineam meam non custodivi
SONG|1|6|indica mihi quem diligit anima mea ubi pascas ubi cubes in meridie ne vagari incipiam per greges sodalium tuorum
SONG|1|7|si ignoras te o pulchra inter mulieres egredere et abi post vestigia gregum et pasce hedos tuos iuxta tabernacula pastorum
SONG|1|8|equitatui meo in curribus Pharaonis adsimilavi te amica mea
SONG|1|9|pulchrae sunt genae tuae sicut turturis collum tuum sicut monilia
SONG|1|10|murenulas aureas faciemus tibi vermiculatas argento
SONG|1|11|dum esset rex in accubitu suo nardus mea dedit odorem suum
SONG|1|12|fasciculus murrae dilectus meus mihi inter ubera mea commorabitur
SONG|1|13|botrus cypri dilectus meus mihi in vineis Engaddi
SONG|1|14|ecce tu pulchra es amica mea ecce tu pulchra oculi tui columbarum
SONG|1|15|ecce tu pulcher es dilecte mi et decorus lectulus noster floridus
SONG|1|16|tigna domorum nostrarum cedrina laquearia nostra cypressina
SONG|2|1|ego flos campi et lilium convallium
SONG|2|2|sicut lilium inter spinas sic amica mea inter filias
SONG|2|3|sicut malum inter ligna silvarum sic dilectus meus inter filios sub umbra illius quam desideraveram sedi et fructus eius dulcis gutturi meo
SONG|2|4|introduxit me in cellam vinariam ordinavit in me caritatem
SONG|2|5|fulcite me floribus stipate me malis quia amore langueo
SONG|2|6|leva eius sub capite meo et dextera illius amplexabitur me
SONG|2|7|adiuro vos filiae Hierusalem per capreas cervosque camporum ne suscitetis neque evigilare faciatis dilectam quoadusque ipsa velit
SONG|2|8|vox dilecti mei ecce iste venit saliens in montibus transiliens colles
SONG|2|9|similis est dilectus meus capreae hinuloque cervorum en ipse stat post parietem nostrum despiciens per fenestras prospiciens per cancellos
SONG|2|10|et dilectus meus loquitur mihi surge propera amica mea formonsa mea et veni
SONG|2|11|iam enim hiemps transiit imber abiit et recessit
SONG|2|12|flores apparuerunt in terra tempus putationis advenit vox turturis audita est in terra nostra
SONG|2|13|ficus protulit grossos suos vineae florent dederunt odorem surge amica mea speciosa mea et veni
SONG|2|14|columba mea in foraminibus petrae in caverna maceriae ostende mihi faciem tuam sonet vox tua in auribus meis vox enim tua dulcis et facies tua decora
SONG|2|15|capite nobis vulpes vulpes parvulas quae demoliuntur vineas nam vinea nostra floruit
SONG|2|16|dilectus meus mihi et ego illi qui pascitur inter lilia
SONG|2|17|donec adspiret dies et inclinentur umbrae revertere similis esto dilecte mi capreae aut hinulo cervorum super montes Bether
SONG|3|1|in lectulo meo per noctes quaesivi quem diligit anima mea quaesivi illum et non inveni
SONG|3|2|surgam et circuibo civitatem per vicos et plateas quaeram quem diligit anima mea quaesivi illum et non inveni
SONG|3|3|invenerunt me vigiles qui custodiunt civitatem num quem dilexit anima mea vidistis
SONG|3|4|paululum cum pertransissem eos inveni quem diligit anima mea tenui eum nec dimittam donec introducam illum in domum matris meae et in cubiculum genetricis meae
SONG|3|5|adiuro vos filiae Hierusalem per capreas cervosque camporum ne suscitetis neque evigilare faciatis dilectam donec ipsa velit
SONG|3|6|quae est ista quae ascendit per desertum sicut virgula fumi ex aromatibus murrae et turis et universi pulveris pigmentarii
SONG|3|7|en lectulum Salomonis sexaginta fortes ambiunt ex fortissimis Israhel
SONG|3|8|omnes tenentes gladios et ad bella doctissimi uniuscuiusque ensis super femur suum propter timores nocturnos
SONG|3|9|ferculum fecit sibi rex Salomon de lignis Libani
SONG|3|10|columnas eius fecit argenteas reclinatorium aureum ascensum purpureum media caritate constravit propter filias Hierusalem
SONG|3|11|egredimini et videte filiae Sion regem Salomonem in diademate quo coronavit eum mater sua in die disponsionis illius et in die laetitiae cordis eius
SONG|4|1|quam pulchra es amica mea quam pulchra es oculi tui columbarum absque eo quod intrinsecus latet capilli tui sicut greges caprarum quae ascenderunt de monte Galaad
SONG|4|2|dentes tui sicut greges tonsarum quae ascenderunt de lavacro omnes gemellis fetibus et sterilis non est inter eas
SONG|4|3|sicut vitta coccinea labia tua et eloquium tuum dulce sicut fragmen mali punici ita genae tuae absque eo quod intrinsecus latet
SONG|4|4|sicut turris David collum tuum quae aedificata est cum propugnaculis mille clypei pendent ex ea omnis armatura fortium
SONG|4|5|duo ubera tua sicut duo hinuli capreae gemelli qui pascuntur in liliis
SONG|4|6|donec adspiret dies et inclinentur umbrae vadam ad montem murrae et ad collem turis
SONG|4|7|tota pulchra es amica mea et macula non est in te
SONG|4|8|veni de Libano sponsa veni de Libano veni coronaberis de capite Amana de vertice Sanir et Hermon de cubilibus leonum de montibus pardorum
SONG|4|9|vulnerasti cor meum soror mea sponsa vulnerasti cor meum in uno oculorum tuorum et in uno crine colli tui
SONG|4|10|quam pulchrae sunt mammae tuae soror mea sponsa pulchriora ubera tua vino et odor unguentorum tuorum super omnia aromata
SONG|4|11|favus distillans labia tua sponsa mel et lac sub lingua tua et odor vestimentorum tuorum sicut odor turis
SONG|4|12|hortus conclusus soror mea sponsa hortus conclusus fons signatus
SONG|4|13|emissiones tuae paradisus malorum punicorum cum pomorum fructibus cypri cum nardo
SONG|4|14|nardus et crocus fistula et cinnamomum cum universis lignis Libani murra et aloe cum omnibus primis unguentis
SONG|4|15|fons hortorum puteus aquarum viventium quae fluunt impetu de Libano
SONG|4|16|surge aquilo et veni auster perfla hortum meum et fluant aromata illius
SONG|5|1|veniat dilectus meus in hortum suum et comedat fructum pomorum suorum veni in hortum meum soror mea sponsa messui murram meam cum aromatibus meis comedi favum cum melle meo bibi vinum meum cum lacte meo comedite amici bibite et inebriamini carissimi
SONG|5|2|ego dormio et cor meum vigilat vox dilecti mei pulsantis aperi mihi soror mea amica mea columba mea inmaculata mea quia caput meum plenum est rore et cincinni mei guttis noctium
SONG|5|3|expoliavi me tunica mea quomodo induar illa lavi pedes meos quomodo inquinabo illos
SONG|5|4|dilectus meus misit manum suam per foramen et venter meus intremuit ad tactum eius
SONG|5|5|surrexi ut aperirem dilecto meo manus meae stillaverunt murra digiti mei pleni murra probatissima
SONG|5|6|pessulum ostii aperui dilecto meo at ille declinaverat atque transierat anima mea liquefacta est ut locutus est quaesivi et non inveni illum vocavi et non respondit mihi
SONG|5|7|invenerunt me custodes qui circumeunt civitatem percusserunt me vulneraverunt me tulerunt pallium meum mihi custodes murorum
SONG|5|8|adiuro vos filiae Hierusalem si inveneritis dilectum meum ut nuntietis ei quia amore langueo
SONG|5|9|qualis est dilectus tuus ex dilecto o pulcherrima mulierum qualis est dilectus tuus ex dilecto quia sic adiurasti nos
SONG|5|10|dilectus meus candidus et rubicundus electus ex milibus
SONG|5|11|caput eius aurum optimum comae eius sicut elatae palmarum nigrae quasi corvus
SONG|5|12|oculi eius sicut columbae super rivulos aquarum quae lacte sunt lotae et resident iuxta fluenta plenissima
SONG|5|13|genae illius sicut areolae aromatum consitae a pigmentariis labia eius lilia distillantia murram primam
SONG|5|14|manus illius tornatiles aureae plenae hyacinthis venter eius eburneus distinctus sapphyris
SONG|5|15|crura illius columnae marmoreae quae fundatae sunt super bases aureas species eius ut Libani electus ut cedri
SONG|5|16|guttur illius suavissimum et totus desiderabilis talis est dilectus meus et iste est amicus meus filiae Hierusalem
SONG|5|17|quo abiit dilectus tuus o pulcherrima mulierum quo declinavit dilectus tuus et quaeremus eum tecum
SONG|6|1|dilectus meus descendit in hortum suum ad areolam aromatis ut pascatur in hortis et lilia colligat
SONG|6|2|ego dilecto meo et dilectus meus mihi qui pascitur inter lilia
SONG|6|3|pulchra es amica mea suavis et decora sicut Hierusalem terribilis ut castrorum acies ordinata
SONG|6|4|averte oculos tuos a me quia ipsi me avolare fecerunt capilli tui sicut grex caprarum quae apparuerunt de Galaad
SONG|6|5|dentes tui sicut grex ovium quae ascenderunt de lavacro omnes gemellis fetibus et sterilis non est in eis
SONG|6|6|sicut cortex mali punici genae tuae absque occultis tuis
SONG|6|7|sexaginta sunt reginae et octoginta concubinae et adulescentularum non est numerus
SONG|6|8|una est columba mea perfecta mea una est matris suae electa genetrici suae viderunt illam filiae et beatissimam praedicaverunt reginae et concubinae et laudaverunt eam
SONG|6|9|quae est ista quae progreditur quasi aurora consurgens pulchra ut luna electa ut sol terribilis ut acies ordinata
SONG|6|10|descendi ad hortum nucum ut viderem poma convallis ut inspicerem si floruisset vinea et germinassent mala punica
SONG|6|11|nescivi anima mea conturbavit me propter quadrigas Aminadab
SONG|6|12|revertere revertere Sulamitis revertere revertere ut intueamur te
SONG|7|1|quid videbis in Sulamiten nisi choros castrorum quam pulchri sunt gressus tui in calciamentis filia principis iunctura feminum tuorum sicut monilia quae fabricata sunt manu artificis
SONG|7|2|umbilicus tuus crater tornatilis numquam indigens poculis venter tuus sicut acervus tritici vallatus liliis
SONG|7|3|duo ubera tua sicut duo hinuli gemelli capreae
SONG|7|4|collum tuum sicut turris eburnea oculi tui sicut piscinae in Esebon quae sunt in porta filiae multitudinis nasus tuus sicut turris Libani quae respicit contra Damascum
SONG|7|5|caput tuum ut Carmelus et comae capitis tui sicut purpura regis vincta canalibus
SONG|7|6|quam pulchra es et quam decora carissima in deliciis
SONG|7|7|statura tua adsimilata est palmae et ubera tua botris
SONG|7|8|dixi ascendam in palmam adprehendam fructus eius et erunt ubera tua sicut botri vineae et odor oris tui sicut malorum
SONG|7|9|guttur tuum sicut vinum optimum dignum dilecto meo ad potandum labiisque et dentibus illius ruminandum
SONG|7|10|ego dilecto meo et ad me conversio eius
SONG|7|11|veni dilecte mi egrediamur in agrum commoremur in villis
SONG|7|12|mane surgamus ad vineas videamus si floruit vinea si flores fructus parturiunt si floruerunt mala punica ibi dabo tibi ubera mea
SONG|7|13|mandragorae dederunt odorem in portis nostris omnia poma nova et vetera dilecte mi servavi tibi
SONG|8|1|quis mihi det te fratrem meum sugentem ubera matris meae ut inveniam te foris et deosculer et iam me nemo despiciat
SONG|8|2|adprehendam te et ducam in domum matris meae ibi me docebis et dabo tibi poculum ex vino condito et mustum malorum granatorum meorum
SONG|8|3|leva eius sub capite meo et dextera illius amplexabitur me
SONG|8|4|adiuro vos filiae Hierusalem ne suscitetis et evigilare faciatis dilectam donec ipsa velit
SONG|8|5|quae est ista quae ascendit de deserto deliciis affluens et nixa super dilectum suum sub arbore malo suscitavi te ibi corrupta est mater tua ibi violata est genetrix tua
SONG|8|6|pone me ut signaculum super cor tuum ut signaculum super brachium tuum quia fortis est ut mors dilectio dura sicut inferus aemulatio lampades eius lampades ignis atque flammarum
SONG|8|7|aquae multae non poterunt extinguere caritatem nec flumina obruent illam si dederit homo omnem substantiam domus suae pro dilectione quasi nihil despicient eum
SONG|8|8|soror nostra parva et ubera non habet quid faciemus sorori nostrae in die quando adloquenda est
SONG|8|9|si murus est aedificemus super eum propugnacula argentea si ostium est conpingamus illud tabulis cedrinis
SONG|8|10|ego murus et ubera mea sicut turris ex quo facta sum coram eo quasi pacem repperiens
SONG|8|11|vinea fuit Pacifico in ea quae habet populos tradidit eam custodibus vir adfert pro fructu eius mille argenteos
SONG|8|12|vinea mea coram me est mille tui Pacifice et ducenti his qui custodiunt fructus eius
SONG|8|13|quae habitas in hortis amici auscultant fac me audire vocem tuam
SONG|8|14|fuge dilecte mi et adsimilare capreae hinuloque cervorum super montes aromatum
ISA|1|1|visio Isaiae filii Amos quam vidit super Iudam et Hierusalem in diebus Oziae Ioatham Ahaz Ezechiae regum Iuda
ISA|1|2|audite caeli et auribus percipe terra quoniam Dominus locutus est filios enutrivi et exaltavi ipsi autem spreverunt me
ISA|1|3|cognovit bos possessorem suum et asinus praesepe domini sui Israhel non cognovit populus meus non intellexit
ISA|1|4|vae genti peccatrici populo gravi iniquitate semini nequam filiis sceleratis dereliquerunt Dominum blasphemaverunt Sanctum Israhel abalienati sunt retrorsum
ISA|1|5|super quo percutiam vos ultra addentes praevaricationem omne caput languidum et omne cor maerens
ISA|1|6|a planta pedis usque ad verticem non est in eo sanitas vulnus et livor et plaga tumens non est circumligata nec curata medicamine neque fota oleo
ISA|1|7|terra vestra deserta civitates vestrae succensae igni regionem vestram coram vobis alieni devorant et desolabitur sicut in vastitate hostili
ISA|1|8|et derelinquetur filia Sion ut umbraculum in vinea et sicut tugurium in cucumerario sicut civitas quae vastatur
ISA|1|9|nisi Dominus exercituum reliquisset nobis semen quasi Sodoma fuissemus et quasi Gomorra similes essemus
ISA|1|10|audite verbum Domini principes Sodomorum percipite auribus legem Dei nostri populus Gomorrae
ISA|1|11|quo mihi multitudinem victimarum vestrarum dicit Dominus plenus sum holocausta arietum et adipem pinguium et sanguinem vitulorum et agnorum et hircorum nolui
ISA|1|12|cum veneritis ante conspectum meum quis quaesivit haec de manibus vestris ut ambularetis in atriis meis
ISA|1|13|ne adferatis ultra sacrificium frustra incensum abominatio est mihi neomeniam et sabbatum et festivitates alias non feram iniqui sunt coetus vestri
ISA|1|14|kalendas vestras et sollemnitates vestras odivit anima mea facta sunt mihi molesta laboravi sustinens
ISA|1|15|et cum extenderitis manus vestras avertam oculos meos a vobis et cum multiplicaveritis orationem non audiam manus vestrae sanguine plenae sunt
ISA|1|16|lavamini mundi estote auferte malum cogitationum vestrarum ab oculis meis quiescite agere perverse
ISA|1|17|discite benefacere quaerite iudicium subvenite oppresso iudicate pupillo defendite viduam
ISA|1|18|et venite et arguite me dicit Dominus si fuerint peccata vestra ut coccinum quasi nix dealbabuntur et si fuerint rubra quasi vermiculus velut lana erunt
ISA|1|19|si volueritis et audieritis bona terrae comedetis
ISA|1|20|quod si nolueritis et me provocaveritis ad iracundiam gladius devorabit vos quia os Domini locutum est
ISA|1|21|quomodo facta est meretrix civitas fidelis plena iudicii iustitia habitavit in ea nunc autem homicidae
ISA|1|22|argentum tuum versum est in scoriam vinum tuum mixtum est aqua
ISA|1|23|principes tui infideles socii furum omnes diligunt munera sequuntur retributiones pupillo non iudicant et causa viduae non ingreditur ad eos
ISA|1|24|propter hoc ait Dominus exercituum Fortis Israhel heu consolabor super hostibus meis et vindicabor de inimicis meis
ISA|1|25|et convertam manum meam ad te et excoquam ad purum scoriam tuam et auferam omne stagnum tuum
ISA|1|26|et restituam iudices tuos ut fuerunt prius et consiliarios tuos sicut antiquitus post haec vocaberis civitas iusti urbs fidelis
ISA|1|27|Sion in iudicio redimetur et reducent eam in iustitia
ISA|1|28|et conteret scelestos et peccatores simul et qui dereliquerunt Dominum consumentur
ISA|1|29|confundentur enim ab idolis quibus sacrificaverunt et erubescetis super hortis quos elegeratis
ISA|1|30|cum fueritis velut quercus defluentibus foliis et velut hortus absque aqua
ISA|1|31|et erit fortitudo vestra ut favilla stuppae et opus vestrum quasi scintilla et succendetur utrumque simul et non erit qui extinguat
ISA|2|1|verbum quod vidit Isaias filius Amos super Iudam et Hierusalem
ISA|2|2|et erit in novissimis diebus praeparatus mons domus Domini in vertice montium et elevabitur super colles et fluent ad eum omnes gentes
ISA|2|3|et ibunt populi multi et dicent venite et ascendamus ad montem Domini et ad domum Dei Iacob et docebit nos vias suas et ambulabimus in semitis eius quia de Sion exibit lex et verbum Domini de Hierusalem
ISA|2|4|et iudicabit gentes et arguet populos multos et conflabunt gladios suos in vomeres et lanceas suas in falces non levabit gens contra gentem gladium nec exercebuntur ultra ad proelium
ISA|2|5|domus Iacob venite et ambulemus in lumine Domini
ISA|2|6|proiecisti enim populum tuum domum Iacob quia repleti sunt ut olim et augures habuerunt ut Philisthim et pueris alienis adheserunt
ISA|2|7|repleta est terra argento et auro et non est finis thesaurorum eius
ISA|2|8|et repleta est terra eius equis et innumerabiles quadrigae eius et repleta est terra eius idolis opus manuum suarum adoraverunt quod fecerunt digiti eorum
ISA|2|9|et incurvavit se homo et humiliatus est vir ne ergo dimittas eis
ISA|2|10|ingredere in petram abscondere fossa humo a facie timoris Domini et a gloria maiestatis eius
ISA|2|11|oculi sublimis hominis humiliati sunt et incurvabitur altitudo virorum exaltabitur autem Dominus solus in die illa
ISA|2|12|quia dies Domini exercituum super omnem superbum et excelsum et super omnem arrogantem et humiliabitur
ISA|2|13|et super omnes cedros Libani sublimes et erectas et super omnes quercus Basan
ISA|2|14|et super omnes montes excelsos et super omnes colles elevatos
ISA|2|15|et super omnem turrem excelsam et super omnem murum munitum
ISA|2|16|et super omnes naves Tharsis et super omne quod visu pulchrum est
ISA|2|17|et incurvabitur sublimitas hominum et humiliabitur altitudo virorum et elevabitur Dominus solus in die illa
ISA|2|18|et idola penitus conterentur
ISA|2|19|et introibunt in speluncas petrarum et in voragines terrae a facie formidinis Domini et a gloria maiestatis eius cum surrexerit percutere terram
ISA|2|20|in die illa proiciet homo idola argenti sui et simulacra auri sui quae fecerat sibi ut adoraret talpas et vespertiliones
ISA|2|21|et ingredietur fissuras petrarum et cavernas saxorum a facie formidinis Domini et a gloria maiestatis eius cum surrexerit percutere terram
ISA|2|22|quiescite ergo ab homine cuius spiritus in naribus eius quia excelsus reputatus est ipse
ISA|3|1|ecce enim Dominator Deus exercituum auferet ab Hierusalem et ab Iuda validum et fortem omne robur panis et omne robur aquae
ISA|3|2|fortem et virum bellatorem iudicem et prophetam et ariolum et senem
ISA|3|3|principem super quinquaginta et honorabilem vultu et consiliarium sapientem de architectis et prudentem eloquii mystici
ISA|3|4|et dabo pueros principes eorum et effeminati dominabuntur eis
ISA|3|5|et inruet populus vir ad virum unusquisque ad proximum suum tumultuabitur puer contra senem et ignobilis contra nobilem
ISA|3|6|adprehendet enim vir fratrem suum domesticum patris sui vestimentum tibi est princeps esto noster ruina autem haec sub manu tua
ISA|3|7|respondebit in die illa dicens non sum medicus et in domo mea non est panis neque vestimentum nolite constituere me principem populi
ISA|3|8|ruit enim Hierusalem et Iudas concidit quia lingua eorum et adinventiones eorum contra Dominum ut provocarent oculos maiestatis eius
ISA|3|9|agnitio vultus eorum respondit eis et peccatum suum quasi Sodomae praedicaverunt nec absconderunt vae animae eorum quoniam reddita sunt eis mala
ISA|3|10|dicite iusto quoniam bene quoniam fructum adinventionum suarum comedet
ISA|3|11|vae impio in malum retributio enim manuum eius fiet ei
ISA|3|12|populum meum exactores sui spoliaverunt et mulieres dominatae sunt eius popule meus qui beatum te dicunt ipsi te decipiunt et viam gressuum tuorum dissipant
ISA|3|13|stat ad iudicandum Dominus et stat ad iudicandos populos
ISA|3|14|Dominus ad iudicium veniet cum senibus populi sui et principibus eius vos enim depasti estis vineam meam et rapina pauperis in domo vestra
ISA|3|15|quare adteritis populum meum et facies pauperum commolitis dicit Dominus Deus exercituum
ISA|3|16|et dixit Dominus pro eo quod elevatae sunt filiae Sion et ambulaverunt extento collo et nutibus oculorum ibant et plaudebant ambulabant et in pedibus suis conposito gradu incedebant
ISA|3|17|decalvabit Dominus verticem filiarum Sion et Dominus crinem earum nudabit
ISA|3|18|in die illa auferet Dominus ornatum calciamentorum et lunulas
ISA|3|19|et torques et monilia et armillas et mitras
ISA|3|20|discriminalia et periscelidas et murenulas et olfactoriola et inaures
ISA|3|21|et anulos et gemmas in fronte pendentes
ISA|3|22|et mutatoria et pallia et linteamina et acus
ISA|3|23|et specula et sindones et vittas et theristra
ISA|3|24|et erit pro suavi odore fetor et pro zona funiculus et pro crispanti crine calvitium et pro fascia pectorali cilicium
ISA|3|25|pulcherrimi quoque viri tui gladio cadent et fortes tui in proelio
ISA|3|26|et maerebunt atque lugebunt portae eius et desolata in terra sedebit
ISA|4|1|et adprehendent septem mulieres virum unum in die illa dicentes panem nostrum comedemus et vestimentis nostris operiemur tantummodo vocetur nomen tuum super nos aufer obprobrium nostrum
ISA|4|2|in die illa erit germen Domini in magnificentia et in gloria et fructus terrae sublimis et exultatio his qui salvati fuerint de Israhel
ISA|4|3|et erit omnis qui relictus fuerit in Sion et residuus in Hierusalem sanctus vocabitur omnis qui scriptus est in vita in Hierusalem
ISA|4|4|si abluerit Dominus sordem filiarum Sion et sanguinem Hierusalem laverit de medio eius spiritu iudicii et spiritu ardoris
ISA|4|5|et creabit Dominus super omnem locum montis Sion et ubi invocatus est nubem per diem et fumum et splendorem ignis flammantis in nocte super omnem enim gloriam protectio
ISA|4|6|et tabernaculum erit in umbraculum diei ab aestu et in securitatem et absconsionem a turbine et a pluvia
ISA|5|1|cantabo dilecto meo canticum patruelis mei vineae suae vinea facta est dilecto meo in cornu filio olei
ISA|5|2|et sepivit eam et lapides elegit ex illa et plantavit eam electam et aedificavit turrem in medio eius et torcular extruxit in ea et expectavit ut faceret uvas et fecit labruscas
ISA|5|3|nunc ergo habitator Hierusalem et vir Iuda iudicate inter me et inter vineam meam
ISA|5|4|quid est quod debui ultra facere vineae meae et non feci ei an quod expectavi ut faceret uvas et fecit labruscas
ISA|5|5|et nunc ostendam vobis quid ego faciam vineae meae auferam sepem eius et erit in direptionem diruam maceriam eius et erit in conculcationem
ISA|5|6|et ponam eam desertam non putabitur et non fodietur et ascendent vepres et spinae et nubibus mandabo ne pluant super eam imbrem
ISA|5|7|vinea enim Domini exercituum domus Israhel et vir Iuda germen delectabile eius et expectavi ut faceret iudicium et ecce iniquitas et iustitiam et ecce clamor
ISA|5|8|vae qui coniungitis domum ad domum et agrum agro copulatis usque ad terminum loci numquid habitabitis soli vos in medio terrae
ISA|5|9|in auribus meis sunt haec Domini exercituum nisi domus multae desertae fuerint grandes et pulchrae absque habitatore
ISA|5|10|decem enim iuga vinearum facient lagunculam unam et triginta modii sementis facient modios tres
ISA|5|11|vae qui consurgitis mane ad ebrietatem sectandam et potandum usque ad vesperam ut vino aestuetis
ISA|5|12|cithara et lyra et tympanum et tibia et vinum in conviviis vestris et opus Domini non respicitis nec opera manuum eius consideratis
ISA|5|13|propterea captivus ductus est populus meus quia non habuit scientiam et nobiles eius interierunt fame et multitudo eius siti exaruit
ISA|5|14|propterea dilatavit infernus animam suam et aperuit os suum absque ullo termino et descendent fortes eius et populus eius et sublimes gloriosique eius ad eum
ISA|5|15|et incurvabitur homo et humiliabitur vir et oculi sublimium deprimentur
ISA|5|16|et exaltabitur Dominus exercituum in iudicio et Deus sanctus sanctificabitur in iustitia
ISA|5|17|et pascentur agni iuxta ordinem suum et deserta in ubertatem versa advenae comedent
ISA|5|18|vae qui trahitis iniquitatem in funiculis vanitatis et quasi vinculum plaustri peccatum
ISA|5|19|qui dicitis festinet et cito veniat opus eius ut videamus et adpropiet et veniat consilium Sancti Israhel et sciemus illud
ISA|5|20|vae qui dicitis malum bonum et bonum malum ponentes tenebras lucem et lucem tenebras ponentes amarum in dulce et dulce in amarum
ISA|5|21|vae qui sapientes estis in oculis vestris et coram vobismet ipsis prudentes
ISA|5|22|vae qui potentes estis ad bibendum vinum et viri fortes ad miscendam ebrietatem
ISA|5|23|qui iustificatis impium pro muneribus et iustitiam iusti aufertis ab eo
ISA|5|24|propter hoc sicut devorat stipulam lingua ignis et calor flammae exurit sic radix eorum quasi favilla erit et germen eorum ut pulvis ascendet abiecerunt enim legem Domini exercituum et eloquium Sancti Israhel blasphemaverunt
ISA|5|25|ideo iratus est furor Domini in populo suo et extendit manum suam super eum et percussit eum et conturbati sunt montes et facta sunt morticina eorum quasi stercus in medio platearum in omnibus his non est aversus furor eius sed adhuc manus eius extenta
ISA|5|26|et levabit signum nationibus procul et sibilabit ad eum de finibus terrae et ecce festinus velociter veniet
ISA|5|27|non est deficiens neque laborans in eo non dormitabit neque dormiet neque solvetur cingulum renum eius nec rumpetur corrigia calciamenti eius
ISA|5|28|sagittae eius acutae et omnes arcus eius extenti ungulae equorum eius ut silex et rotae eius quasi impetus tempestatis
ISA|5|29|rugitus eius ut leonis rugiet ut catuli leonum et frendet et tenebit praedam et amplexabitur et non erit qui eruat
ISA|5|30|et sonabit super eum in die illa sicut sonitus maris aspiciemus in terram et ecce tenebrae tribulationis et lux obtenebrata est in caligine eius
ISA|6|1|in anno quo mortuus est rex Ozias vidi Dominum sedentem super solium excelsum et elevatum et ea quae sub eo erant implebant templum
ISA|6|2|seraphin stabant super illud sex alae uni et sex alae alteri duabus velabant faciem eius et duabus velabant pedes eius et duabus volabant
ISA|6|3|et clamabant alter ad alterum et dicebant sanctus sanctus sanctus Dominus exercituum plena est omnis terra gloria eius
ISA|6|4|et commota sunt superliminaria cardinum a voce clamantis et domus impleta est fumo
ISA|6|5|et dixi vae mihi quia tacui quia vir pollutus labiis ego sum et in medio populi polluta labia habentis ego habito et Regem Dominum exercituum vidi oculis meis
ISA|6|6|et volavit ad me unus de seraphin et in manu eius calculus quem forcipe tulerat de altari
ISA|6|7|et tetigit os meum et dixit ecce tetigit hoc labia tua et auferetur iniquitas tua et peccatum tuum mundabitur
ISA|6|8|et audivi vocem Domini dicentis quem mittam et quis ibit nobis et dixi ecce ego sum mitte me
ISA|6|9|et dixit vade et dices populo huic audite audientes et nolite intellegere et videte visionem et nolite cognoscere
ISA|6|10|excaeca cor populi huius et aures eius adgrava et oculos eius claude ne forte videat oculis suis et auribus suis audiat et corde suo intellegat et convertatur et sanem eum
ISA|6|11|et dixi usquequo Domine et dixit donec desolentur civitates absque habitatore et domus sine homine et terra relinquetur deserta
ISA|6|12|et longe faciet Dominus homines et multiplicabitur quae derelicta fuerat in medio terrae
ISA|6|13|et adhuc in ea decimatio et convertetur et erit in ostensionem sicut terebinthus et sicuti quercus quae expandit ramos suos semen sanctum erit id quod steterit in ea
ISA|7|1|et factum est in diebus Ahaz filii Ioatham filii Oziae regis Iuda ascendit Rasin rex Syriae et Phacee filius Romeliae rex Israhel in Hierusalem ad proeliandum contra eam et non potuerunt debellare eam
ISA|7|2|et nuntiaverunt domui David dicentes requievit Syria super Ephraim et commotum est cor eius et cor populi eius sicut moventur ligna silvarum a facie venti
ISA|7|3|et dixit Dominus ad Isaiam egredere in occursum Ahaz tu et qui derelictus est Iasub filius tuus ad extremum aquaeductus piscinae superioris in via agri Fullonis
ISA|7|4|et dices ad eum vide ut sileas noli timere et cor tuum ne formidet a duobus caudis titionum fumigantium istorum in ira furoris Rasin et Syriae et filii Romeliae
ISA|7|5|eo quod consilium inierit contra te Syria malum Ephraim et filius Romeliae dicentes
ISA|7|6|ascendamus ad Iudam et suscitemus eum et avellamus eum ad nos et ponamus regem in medio eius filium Tabeel
ISA|7|7|haec dicit Dominus Deus non stabit et non erit istud
ISA|7|8|sed caput Syriae Damascus et caput Damasci Rasin et adhuc sexaginta et quinque anni et desinet Ephraim esse populus
ISA|7|9|et caput Ephraim Samaria et caput Samariae filius Romeliae si non credideritis non permanebitis
ISA|7|10|et adiecit Dominus loqui ad Ahaz dicens
ISA|7|11|pete tibi signum a Domino Deo tuo in profundum inferni sive in excelsum supra
ISA|7|12|et dixit Ahaz non petam et non temptabo Dominum
ISA|7|13|et dixit audite ergo domus David numquid parum vobis est molestos esse hominibus quia molesti estis et Deo meo
ISA|7|14|propter hoc dabit Dominus ipse vobis signum ecce virgo concipiet et pariet filium et vocabitis nomen eius Emmanuhel
ISA|7|15|butyrum et mel comedet ut sciat reprobare malum et eligere bonum
ISA|7|16|quia antequam sciat puer reprobare malum et eligere bonum derelinquetur terra quam tu detestaris a facie duum regum suorum
ISA|7|17|adducet Dominus super te et super populum tuum et super domum patris tui dies qui non venerunt a diebus separationis Ephraim a Iuda cum rege Assyriorum
ISA|7|18|et erit in die illa sibilabit Dominus muscae quae est in extremo fluminum Aegypti et api quae est in terra Assur
ISA|7|19|et venient et requiescent omnes in torrentibus vallium et cavernis petrarum et in omnibus frutectis et in universis foraminibus
ISA|7|20|in die illa radet Dominus in novacula conducta in his qui trans Flumen sunt in rege Assyriorum caput et pilos pedum et barbam universam
ISA|7|21|et erit in die illa nutriet homo vaccam boum et duas oves
ISA|7|22|et prae ubertate lactis comedet butyrum butyrum enim et mel manducabit omnis qui relictus fuerit in medio terrae
ISA|7|23|et erit in die illa omnis locus ubi fuerint mille vites mille argenteis et in spinas et in vepres erunt
ISA|7|24|cum sagittis et arcu ingredientur illuc vepres enim et spinae erunt in universa terra
ISA|7|25|et omnes montes qui in sarculo sarientur non veniet illuc terror spinarum et veprium et erit in pascua bovis et in conculcationem pecoris
ISA|8|1|et dixit Dominus ad me sume tibi librum grandem et scribe in eo stilo hominis Velociter spolia detrahe Cito praedare
ISA|8|2|et adhibui mihi testes fideles Uriam sacerdotem et Zacchariam filium Barachiae
ISA|8|3|et accessi ad prophetissam et concepit et peperit filium et dixit Dominus ad me voca nomen eius Adcelera spolia detrahere Festina praedari
ISA|8|4|quia antequam sciat puer vocare patrem suum et matrem suam auferetur fortitudo Damasci et spolia Samariae coram rege Assyriorum
ISA|8|5|et adiecit Dominus loqui ad me adhuc dicens
ISA|8|6|pro eo quod abiecit populus iste aquas Siloae quae vadunt cum silentio et adsumpsit magis Rasin et filium Romeliae
ISA|8|7|propter hoc ecce Dominus adducet super eos aquas Fluminis fortes et multas regem Assyriorum et omnem gloriam eius et ascendet super omnes rivos eius et fluet super universas ripas eius
ISA|8|8|et ibit per Iudam inundans et transiens usque ad collum veniet et erit extensio alarum eius implens latitudinem terrae tuae o Emmanuhel
ISA|8|9|congregamini populi et vincimini et audite universae procul terrae confortamini et vincimini accingite vos et vincimini
ISA|8|10|inite consilium et dissipabitur loquimini verbum et non fiet quia nobiscum Deus
ISA|8|11|haec enim ait Dominus ad me sicut in forti manu erudivit me ne irem in via populi huius dicens
ISA|8|12|non dicatis coniuratio omnia enim quae loquitur populus iste coniuratio est et timorem eius ne timeatis neque paveatis
ISA|8|13|Dominum exercituum ipsum sanctificate ipse pavor vester et ipse terror vester
ISA|8|14|et erit vobis in sanctificationem in lapidem autem offensionis et in petram scandali duabus domibus Israhel in laqueum et in ruinam habitantibus Hierusalem
ISA|8|15|et offendent ex eis plurimi et cadent et conterentur et inretientur et capientur
ISA|8|16|liga testimonium signa legem in discipulis meis
ISA|8|17|et expectabo Dominum qui abscondit faciem suam a domo Iacob et praestolabor eum
ISA|8|18|ecce ego et pueri quos mihi dedit Dominus in signum et in portentum Israhelis a Domino exercituum qui habitat in monte Sion
ISA|8|19|et cum dixerint ad vos quaerite a pythonibus et a divinis qui stridunt in incantationibus suis numquid non populus a Deo suo requirit pro vivis a mortuis
ISA|8|20|ad legem magis et ad testimonium quod si non dixerint iuxta verbum hoc non erit eis matutina lux
ISA|8|21|et transibit per eam corruet et esuriet et cum esurierit irascetur et maledicet regi suo et Deo suo et suspiciet sursum
ISA|8|22|et ad terram intuebitur et ecce tribulatio et tenebrae dissolutio angustia et caligo persequens et non poterit avolare de angustia sua
ISA|9|1|primo tempore adleviata est terra Zabulon et terra Nepthalim et novissimo adgravata est via maris trans Iordanem Galileae gentium
ISA|9|2|populus qui ambulabat in tenebris vidit lucem magnam habitantibus in regione umbrae mortis lux orta est eis
ISA|9|3|multiplicasti gentem non magnificasti laetitiam laetabuntur coram te sicut laetantur in messe sicut exultant quando dividunt spolia
ISA|9|4|iugum enim oneris eius et virgam umeri eius et sceptrum exactoris eius superasti sicut in die Madian
ISA|9|5|quia omnis violenta praedatio cum tumultu et vestimentum mixtum sanguine erit in conbustionem et cibus ignis
ISA|9|6|parvulus enim natus est nobis filius datus est nobis et factus est principatus super umerum eius et vocabitur nomen eius Admirabilis consiliarius Deus fortis Pater futuri saeculi Princeps pacis
ISA|9|7|multiplicabitur eius imperium et pacis non erit finis super solium David et super regnum eius ut confirmet illud et corroboret in iudicio et iustitia amodo et usque in sempiternum zelus Domini exercituum faciet hoc
ISA|9|8|verbum misit Dominus in Iacob et cecidit in Israhel
ISA|9|9|et sciet populus omnis Ephraim et habitantes Samariam in superbia et magnitudine cordis dicentes
ISA|9|10|lateres ceciderunt sed quadris lapidibus aedificabimus sycomoros succiderunt sed cedros inmutabimus
ISA|9|11|et elevabit Dominus hostes Rasin super eum et inimicos eius in tumultum vertet
ISA|9|12|Syriam ab oriente et Philisthim ab occidente et devorabunt Israhel toto ore in omnibus his non est aversus furor eius sed adhuc manus eius extenta
ISA|9|13|et populus non est reversus ad percutientem se et Dominum exercituum non inquisierunt
ISA|9|14|et disperdet Dominus ab Israhel caput et caudam incurvantem et refrenantem die una
ISA|9|15|longevus et honorabilis ipse est caput et propheta docens mendacium ipse cauda est
ISA|9|16|et erunt qui beatificant populum istum seducentes et qui beatificantur praecipitati
ISA|9|17|propter hoc super adulescentulis eius non laetabitur Dominus et pupillorum eius et viduarum non miserebitur quia omnis hypocrita est et nequam et universum os locutum est stultitiam in omnibus his non est aversus furor eius sed adhuc manus eius extenta
ISA|9|18|succensa est enim quasi ignis impietas veprem et spinam vorabit et succendetur in densitate saltus et convolvetur superbia fumi
ISA|9|19|in ira Domini exercituum conturbata est terra et erit populus quasi esca ignis vir fratri suo non parcet
ISA|9|20|et declinabit ad dexteram et esuriet et comedet ad sinistram et non saturabitur unusquisque carnem brachii sui vorabit Manasses Ephraim et Ephraim Manassen simul ipsi contra Iudam
ISA|9|21|in omnibus his non est aversus furor eius sed adhuc manus eius extenta
ISA|10|1|vae qui condunt leges iniquas et scribentes iniustitiam scripserunt
ISA|10|2|ut opprimerent in iudicio pauperes et vim facerent causae humilium populi mei ut essent viduae praeda eorum et pupillos diriperent
ISA|10|3|quid facietis in die visitationis et calamitatis de longe venientis ad cuius fugietis auxilium et ubi derelinquetis gloriam vestram
ISA|10|4|ne incurvemini sub vinculo et cum interfectis cadatis super omnibus his non est aversus furor eius sed adhuc manus eius extenta
ISA|10|5|vae Assur virga furoris mei et baculus ipse in manu eorum indignatio mea
ISA|10|6|ad gentem fallacem mittam eum et contra populum furoris mei mandabo illi ut auferat spolia et diripiat praedam et ponat illum in conculcationem quasi lutum platearum
ISA|10|7|ipse autem non sic arbitrabitur et cor eius non ita aestimabit sed ad conterendum erit cor eius et ad internicionem gentium non paucarum
ISA|10|8|dicet enim
ISA|10|9|numquid non principes mei simul reges sunt numquid non ut Charchamis sic Chalanno et ut Arfad sic Emath numquid non ut Damascus sic Samaria
ISA|10|10|quomodo invenit manus mea regna idoli sic et simulacra eorum de Hierusalem et de Samaria
ISA|10|11|numquid non sicut feci Samariae et idolis eius sic faciam Hierusalem et simulacris eius
ISA|10|12|et erit cum impleverit Dominus cuncta opera sua in monte Sion et in Hierusalem visitabo super fructum magnifici cordis regis Assur et super gloriam altitudinis oculorum eius
ISA|10|13|dixit enim in fortitudine manus meae feci et in sapientia mea intellexi et abstuli terminos populorum et principes eorum depraedatus sum et detraxi quasi potens in sublime residentes
ISA|10|14|et invenit quasi nidum manus mea fortitudinem populorum et sicut colliguntur ova quae derelicta sunt sic universam terram ego congregavi et non fuit qui moveret pinnam et aperiret os et ganniret
ISA|10|15|numquid gloriabitur securis contra eum qui secat in ea aut exaltabitur serra contra eum a quo trahitur quomodo si elevetur virga contra levantem se et exaltetur baculus qui utique lignum est
ISA|10|16|propter hoc mittet Dominator Deus exercituum in pinguibus eius tenuitatem et subtus gloriam eius succensa ardebit quasi conbustio ignis
ISA|10|17|et erit lumen Israhel in igne et Sanctus eius in flamma et succendetur et devorabitur spina eius et vepres in die una
ISA|10|18|et gloria saltus eius et Carmeli eius ab anima usque ad carnem consumetur et erit terrore profugus
ISA|10|19|et reliquiae ligni saltus eius pro paucitate numerabuntur et puer scribet eos
ISA|10|20|et erit in die illa non adiciet residuum Israhel et hii qui fugerint de domo Iacob inniti super eo qui percutit eos sed innitetur super Dominum Sanctum Israhel in veritate
ISA|10|21|reliquiae convertentur reliquiae inquam Iacob ad Deum fortem
ISA|10|22|si enim fuerit populus tuus Israhel quasi harena maris reliquiae convertentur ex eo consummatio adbreviata inundabit iustitiam
ISA|10|23|consummationem enim et adbreviationem Dominus Deus exercituum faciet in medio omnis terrae
ISA|10|24|propter hoc haec dicit Dominus Deus exercituum noli timere populus meus habitator Sion ab Assur in virga percutiet te et baculum suum levabit super te in via Aegypti
ISA|10|25|adhuc enim paululum modicumque et consummabitur indignatio et furor meus super scelus eorum
ISA|10|26|et suscitabit super eum Dominus exercituum flagellum iuxta plagam Madian in petra Oreb et virgam suam super mare et levabit eam in via Aegypti
ISA|10|27|et erit in die illa auferetur onus eius de umero tuo et iugum eius de collo tuo et conputrescet iugum a facie olei
ISA|10|28|veniet in Aiath transibit in Magron apud Machmas commendabit vasa sua
ISA|10|29|transierunt cursim Gabee sedes nostra obstipuit Rama Gabaath Saulis fugit
ISA|10|30|hinni voce tua filia Gallim adtende Laisa paupercula Anathoth
ISA|10|31|migravit Medemena habitatores Gebim confortamini
ISA|10|32|adhuc dies est ut in Nob stetur agitabit manum suam super montem filiae Sion collem Hierusalem
ISA|10|33|ecce Dominator Dominus exercituum confringet lagunculam in terrore et excelsi statura succidentur et sublimes humiliabuntur
ISA|10|34|et subvertentur condensa saltus ferro et Libanus cum excelsis cadet
ISA|11|1|et egredietur virga de radice Iesse et flos de radice eius ascendet
ISA|11|2|et requiescet super eum spiritus Domini spiritus sapientiae et intellectus spiritus consilii et fortitudinis spiritus scientiae et pietatis
ISA|11|3|et replebit eum spiritus timoris Domini non secundum visionem oculorum iudicabit neque secundum auditum aurium arguet
ISA|11|4|sed iudicabit in iustitia pauperes et arguet in aequitate pro mansuetis terrae et percutiet terram virga oris sui et spiritu labiorum suorum interficiet impium
ISA|11|5|et erit iustitia cingulum lumborum eius et fides cinctorium renis eius
ISA|11|6|habitabit lupus cum agno et pardus cum hedo accubabit vitulus et leo et ovis simul morabuntur et puer parvulus minabit eos
ISA|11|7|vitulus et ursus pascentur simul requiescent catuli eorum et leo quasi bos comedet paleas
ISA|11|8|et delectabitur infans ab ubere super foramine aspidis et in caverna reguli qui ablactatus fuerit manum suam mittet
ISA|11|9|non nocebunt et non occident in universo monte sancto meo quia repleta est terra scientia Domini sicut aquae maris operientes
ISA|11|10|in die illa radix Iesse qui stat in signum populorum ipsum gentes deprecabuntur et erit sepulchrum eius gloriosum
ISA|11|11|et erit in die illa adiciet Dominus secundo manum suam ad possidendum residuum populi sui quod relinquetur ab Assyriis et ab Aegypto et a Fetros et ab Aethiopia et ab Aelam et a Sennaar et ab Emath et ab insulis maris
ISA|11|12|et levabit signum in nationes et congregabit profugos Israhel et dispersos Iuda colliget a quattuor plagis terrae
ISA|11|13|et auferetur zelus Ephraim et hostes Iuda peribunt Ephraim non aemulabitur Iudam et Iudas non pugnabit contra Ephraim
ISA|11|14|et volabunt in umeros Philisthim per mare simul praedabuntur filios orientis Idumea et Moab praeceptum manus eorum et filii Ammon oboedientes erunt
ISA|11|15|et desolabit Dominus linguam maris Aegypti et levabit manum suam super Flumen in fortitudine spiritus sui et percutiet eum in septem rivis ita ut transeant per eum calciati
ISA|11|16|et erit via residuo populo meo qui relinquetur ab Assyriis sicut fuit Israhel in die qua ascendit de terra Aegypti
ISA|12|1|et dices in illa die confitebor tibi Domine quoniam iratus es mihi conversus est furor tuus et consolatus es me
ISA|12|2|ecce Deus salvator meus fiducialiter agam et non timebo quia fortitudo mea et laus mea Dominus Deus et factus est mihi in salutem
ISA|12|3|haurietis aquas in gaudio de fontibus salvatoris
ISA|12|4|et dicetis in illa die confitemini Domino et invocate nomen eius notas facite in populis adinventiones eius mementote quoniam excelsum est nomen eius
ISA|12|5|cantate Domino quoniam magnifice fecit adnuntiate hoc in universa terra
ISA|12|6|exulta et lauda habitatio Sion quia magnus in medio tui Sanctus Israhel
ISA|13|1|onus Babylonis quod vidit Isaias filius Amos
ISA|13|2|super montem caligosum levate signum exaltate vocem levate manum et ingrediantur portas duces
ISA|13|3|ego mandavi sanctificatis meis et vocavi fortes meos in ira mea exultantes in gloria mea
ISA|13|4|vox multitudinis in montibus quasi populorum frequentium vox sonitus regum gentium congregatarum Dominus exercituum praecepit militiae belli
ISA|13|5|venientibus de terra procul a summitate caeli Dominus et vasa furoris eius ut disperdat omnem terram
ISA|13|6|ululate quia prope est dies Domini quasi vastitas a Domino veniet
ISA|13|7|propter hoc omnes manus dissolventur et omne cor hominis tabescet
ISA|13|8|et conteretur tortiones et dolores tenebunt quasi parturiens dolebunt unusquisque ad proximum suum stupebit facies conbustae vultus eorum
ISA|13|9|ecce dies Domini venit crudelis et indignationis plenus et irae furorisque ad ponendam terram in solitudine et peccatores eius conterendos de ea
ISA|13|10|quoniam stellae caeli et splendor earum non expandent lumen suum obtenebratus est sol in ortu suo et luna non splendebit in lumine suo
ISA|13|11|et visitabo super orbis mala et contra impios iniquitatem eorum et quiescere faciam superbiam infidelium et arrogantiam fortium humiliabo
ISA|13|12|pretiosior erit vir auro et homo mundo obrizo
ISA|13|13|super hoc caelum turbabo et movebitur terra de loco suo propter indignationem Domini exercituum et propter diem irae furoris eius
ISA|13|14|et erit quasi dammula fugiens et quasi ovis et non erit qui congreget unusquisque ad populum suum convertetur et singuli ad terram suam fugient
ISA|13|15|omnis qui inventus fuerit occidetur et omnis qui supervenerit cadet in gladio
ISA|13|16|infantes eorum adlident in oculis eorum diripientur domus eorum et uxores eorum violabuntur
ISA|13|17|ecce ego suscitabo super eos Medos qui argentum non quaerant nec aurum velint
ISA|13|18|sed sagittis parvulos interficiant et lactantibus uteri non misereantur et super filios non parcat oculus eorum
ISA|13|19|et erit Babylon illa gloriosa in regnis inclita in superbia Chaldeorum sicut subvertit Deus Sodomam et Gomorram
ISA|13|20|non habitabitur usque in finem et non fundabitur usque ad generationem et generationem nec ponet ibi tentoria Arabs nec pastores requiescent ibi
ISA|13|21|sed requiescent ibi bestiae et replebuntur domus eorum draconibus et habitabunt ibi strutiones et pilosi saltabunt ibi
ISA|13|22|et respondebunt ibi ululae in aedibus eius et sirenae in delubris voluptatis
ISA|14|1|prope est ut veniat tempus eius et dies eius non elongabuntur miserebitur enim Dominus Iacob et eliget adhuc de Israhel et requiescere eos faciet super humum suam adiungetur advena ad eos et adherebit domui Iacob
ISA|14|2|et tenebunt eos populi et adducent eos in locum suum et possidebit eos domus Israhel super terram Domini in servos et ancillas et erunt capientes eos qui se ceperant et subicient exactores suos
ISA|14|3|et erit in die illa cum requiem dederit tibi Deus a labore tuo et a concussione tua et a servitute dura qua ante servisti
ISA|14|4|sumes parabolam istam contra regem Babylonis et dices quomodo cessavit exactor quievit tributum
ISA|14|5|contrivit Dominus baculum impiorum virgam dominantium
ISA|14|6|caedentem populos in indignatione plaga insanabili subicientem in furore gentes persequentem crudeliter
ISA|14|7|conquievit et siluit omnis terra gavisa est et exultavit
ISA|14|8|abietes quoque laetatae sunt super te et cedri Libani ex quo dormisti non ascendit qui succidat nos
ISA|14|9|infernus subter conturbatus est in occursum adventus tui suscitavit tibi gigantas omnes principes terrae surrexerunt de soliis suis omnes principes nationum
ISA|14|10|universi respondebunt et dicent tibi et tu vulneratus es sicut nos nostri similis effectus es
ISA|14|11|detracta est ad inferos superbia tua concidit cadaver tuum subter te sternetur tinea et operimentum tuum erunt vermes
ISA|14|12|quomodo cecidisti de caelo lucifer qui mane oriebaris corruisti in terram qui vulnerabas gentes
ISA|14|13|qui dicebas in corde tuo in caelum conscendam super astra Dei exaltabo solium meum sedebo in monte testamenti in lateribus aquilonis
ISA|14|14|ascendam super altitudinem nubium ero similis Altissimo
ISA|14|15|verumtamen ad infernum detraheris in profundum laci
ISA|14|16|qui te viderint ad te inclinabuntur teque prospicient numquid iste est vir qui conturbavit terram qui concussit regna
ISA|14|17|qui posuit orbem desertum et urbes eius destruxit vinctis eius non aperuit carcerem
ISA|14|18|omnes reges gentium universi dormierunt in gloria vir in domo sua
ISA|14|19|tu autem proiectus es de sepulchro tuo quasi stirps inutilis pollutus et obvolutus qui interfecti sunt gladio et descenderunt ad fundamenta laci quasi cadaver putridum
ISA|14|20|non habebis consortium neque cum eis in sepultura tu enim terram disperdisti tu populum occidisti non vocabitur in aeternum semen pessimorum
ISA|14|21|praeparate filios eius occisioni in iniquitate patrum eorum non consurgent nec hereditabunt terram neque implebunt faciem orbis civitatum
ISA|14|22|et consurgam super eos dicit Dominus exercituum et perdam Babylonis nomen et reliquias et germen et progeniem ait Dominus
ISA|14|23|et ponam eam in possessionem ericii et in paludes aquarum et scopabo eam in scopa terens dicit Dominus exercituum
ISA|14|24|iuravit Dominus exercituum dicens si non ut putavi ita erit et quomodo mente tractavi
ISA|14|25|sic eveniet ut conteram Assyrium in terra mea et in montibus meis conculcem eum et auferetur ab eis iugum eius et onus illius ab umero eorum tolletur
ISA|14|26|hoc consilium quod cogitavi super omnem terram et haec est manus extenta super universas gentes
ISA|14|27|Dominus enim exercituum decrevit et quis poterit infirmare et manus eius extenta et quis avertet eam
ISA|14|28|in anno quo mortuus est rex Ahaz factum est onus istud
ISA|14|29|ne laeteris Philisthea omnis tu quoniam comminuta est virga percussoris tui de radice enim colubri egredietur regulus et semen eius absorbens volucrem
ISA|14|30|et pascentur primogeniti pauperum et pauperes fiducialiter requiescent et interire faciam in fame radicem tuam et reliquias tuas interficiam
ISA|14|31|ulula porta clama civitas prostrata est Philisthea omnis ab aquilone enim fumus venit et non est qui effugiat agmen eius
ISA|14|32|et quid respondebitur nuntiis gentis quia Dominus fundavit Sion et in ipsa sperabunt pauperes populi eius
ISA|15|1|onus Moab quia nocte vastata est Ar Moab conticuit quia nocte vastatus est murus Moab conticuit
ISA|15|2|ascendit domus et Dibon ad excelsa in planctum super Nabo et super Medaba Moab ululabit in cunctis capitibus eius calvitium omnis barba radetur
ISA|15|3|in triviis eius accincti sunt sacco super tecta eius et in plateis eius omnis ululat descendit in fletum
ISA|15|4|clamavit Esebon et Eleale usque Iasa audita est vox eorum super hoc expediti Moab ululabunt anima eius ululabit sibi
ISA|15|5|cor meum ad Moab clamabit vectes eius usque ad Segor vitulam conternantem per ascensum enim Luith flens ascendet et in via Oronaim clamorem contritionis levabunt
ISA|15|6|aquae enim Nemrim desertae erunt quia aruit herba defecit germen viror omnis interiit
ISA|15|7|secundum magnitudinem operis et visitatio eorum ad torrentem salicum ducent eos
ISA|15|8|quoniam circumiit clamor terminum Moab usque ad Gallim ululatus eius et usque ad puteum Helim clamor eius
ISA|15|9|quia aquae Dibon repletae sunt sanguine ponam enim super Dibon additamenta his qui fugerint de Moab leonem et reliquiis terrae
ISA|16|1|emitte agnum dominatorem terrae de Petra deserti ad montem filiae Sion
ISA|16|2|et erit sicut avis fugiens et pulli de nido avolantes sic erunt filiae Moab in transcensu Arnon
ISA|16|3|ini consilium coge concilium pone quasi noctem umbram tuam in meridie absconde fugientes et vagos ne prodas
ISA|16|4|habitabunt apud te profugi mei Moab esto latibulum eorum a facie vastatoris finitus est enim pulvis consummatus est miser defecit qui conculcabat terram
ISA|16|5|et praeparabitur in misericordia solium et sedebit super eum in veritate in tabernaculo David iudicans et quaerens iudicium et velociter reddens quod iustum est
ISA|16|6|audivimus superbiam Moab superbus est valde superbia eius et arrogantia eius et indignatio eius plus quam fortitudo eius
ISA|16|7|idcirco ululabit Moab ad Moab universus ululabit his qui laetantur super muro cocti lateris loquimini plagas suas
ISA|16|8|quoniam suburbana Esebon deserta sunt et vinea Sabama domini gentium exciderunt flagella eius usque ad Iazer pervenerunt erraverunt in deserto propagines eius relictae sunt transierunt mare
ISA|16|9|super hoc plorabo in fletu Iazer vineam Sabama inebriabo te lacrima mea Esebon et Eleale quoniam super vindemiam tuam et super messem tuam vox calcantium inruit
ISA|16|10|et auferetur laetitia et exultatio de Carmelo et in vineis non exultabit neque iubilabit vinum in torculari non calcabit qui calcare consueverat vocem calcantium abstuli
ISA|16|11|super hoc venter meus ad Moab quasi cithara sonabit et viscera mea ad murum cocti lateris
ISA|16|12|et erit cum apparuerit quod laboravit Moab super excelsis suis ingredietur ad sancta sua ut obsecret et non valebit
ISA|16|13|hoc verbum quod locutus est Dominus ad Moab ex tunc
ISA|16|14|et nunc locutus est Dominus dicens in tribus annis quasi anni mercennarii auferetur gloria Moab super omni populo multo et relinquetur parvus et modicus nequaquam multus
ISA|17|1|onus Damasci ecce Damascus desinet esse civitas et erit sicut acervus lapidum in ruina
ISA|17|2|derelictae civitates Aroer gregibus erunt et requiescent ibi et non erit qui exterreat
ISA|17|3|et cessabit adiutorium ab Ephraim et regnum a Damasco et reliquiae Syriae sicut gloria filiorum Israhel erunt dicit Dominus exercituum
ISA|17|4|et erit in die illa adtenuabitur gloria Iacob et pingue carnis eius marcescet
ISA|17|5|et erit sicut congregans in messe quod restiterit et brachium eius spicas leget et erit sicut quaerens spicas in valle Rafaim
ISA|17|6|et relinquetur in eo sicut racemus et sicut excussio oleae duarum aut trium olivarum in summitate rami sive quattuor aut quinque in cacuminibus eius fructus eius dicit Dominus Deus Israhel
ISA|17|7|in die illa inclinabitur homo ad factorem suum et oculi eius ad Sanctum Israhel respicient
ISA|17|8|et non inclinabitur ad altaria quae fecerunt manus eius et quae operati sunt digiti eius non respiciet lucos et delubra
ISA|17|9|in die illa erunt civitates fortitudinis eius derelictae sicut aratra et segetes quae derelictae sunt a facie filiorum Israhel et erit deserta
ISA|17|10|quia oblita es Dei salvatoris tui et Fortis adiutoris tui non es recordata propterea plantabis plantationem fidelem et germen alienum seminabis
ISA|17|11|in die plantationis tuae labrusca et mane semen tuum florebit ablata est messis in die hereditatis et dolebit graviter
ISA|17|12|vae multitudo populorum multorum ut multitudo maris sonantis et tumultus turbarum sicut sonitus aquarum multarum
ISA|17|13|sonabunt populi sicut sonitus aquarum inundantium et increpabit eum et fugiet procul et rapietur sicut pulvis montium a facie venti et sicut turbo coram tempestate
ISA|17|14|in tempore vespere et ecce turbatio in matutino et non subsistet haec est pars eorum qui vastaverunt nos et sors diripientium nos
ISA|18|1|vae terrae cymbalo alarum quae est trans flumina Aethiopiae
ISA|18|2|qui mittit in mari legatos et in vasis papyri super aquas ite angeli veloces ad gentem convulsam et dilaceratam ad populum terribilem post quem non est alius gentem expectantem expectantem et conculcatam cuius diripuerunt flumina terram eius
ISA|18|3|omnes habitatores orbis qui moramini in terra cum elevatum fuerit signum in montibus videbitis et clangorem tubae audietis
ISA|18|4|quia haec dicit Dominus ad me quiescam et considerabo in loco meo sicut meridiana lux clara est et sicut nubes roris in die messis
ISA|18|5|ante messem enim totus effloruit et inmatura perfectio germinabit et praecidentur ramusculi eius falcibus et quae derelicta fuerint abscidentur excutientur
ISA|18|6|et relinquentur simul avibus montium et bestiis terrae et aestate perpetua erunt super eum volucres et omnes bestiae terrae super illum hiemabunt
ISA|18|7|in tempore illo deferetur munus Domino exercituum a populo divulso et dilacerato a populo terribili post quem non fuit alius a gente expectante expectante et conculcata cuius diripuerunt flumina terram eius ad locum nominis Domini exercituum montem Sion
ISA|19|1|onus Aegypti ecce Dominus ascendet super nubem levem et ingredietur Aegyptum et movebuntur simulacra Aegypti a facie eius et cor Aegypti tabescet in medio eius
ISA|19|2|et concurrere faciam Aegyptios adversum Aegyptios et pugnabit vir contra fratrem suum et vir contra amicum suum civitas adversus civitatem regnum adversus regnum
ISA|19|3|et disrumpetur spiritus Aegypti in visceribus eius et consilium eius praecipitabo et interrogabunt simulacra sua et divinos suos et pythones et ariolos
ISA|19|4|et tradam Aegyptum in manu dominorum crudelium et rex fortis dominabitur eorum ait Dominus Deus exercituum
ISA|19|5|et arescet aqua de mari et fluvius desolabitur atque siccabitur
ISA|19|6|et deficient flumina adtenuabuntur et siccabuntur rivi aggerum calamus et iuncus marcescet
ISA|19|7|nudabitur alveus rivi a fonte suo et omnis sementis inrigua siccabitur arescet et non erit
ISA|19|8|et maerebunt piscatores et lugebunt omnes mittentes in flumen hamum et expandentes rete super faciem aquae marcescent
ISA|19|9|confundentur qui operabantur linum pectentes et texentes subtilia
ISA|19|10|et erunt inrigua eius flaccentia omnes qui faciebant lacunas ad capiendos pisces
ISA|19|11|stulti principes Taneos sapientes consiliarii Pharao dederunt consilium insipiens quomodo dicetis Pharaoni filius sapientium ego filius regum antiquorum
ISA|19|12|ubi sunt nunc sapientes tui adnuntient tibi et indicent quid cogitaverit Dominus exercituum super Aegyptum
ISA|19|13|stulti facti sunt principes Taneos emarcuerunt principes Mempheos deceperunt Aegyptum angulum populorum eius
ISA|19|14|Dominus miscuit in medio eius spiritum vertiginis et errare fecerunt Aegyptum in omni opere suo sicut errat ebrius et vomens
ISA|19|15|et non erit Aegypto opus quod faciat caput et caudam incurvantem et refrenantem
ISA|19|16|in die illa erit Aegyptus quasi mulieres et stupebunt et timebunt a facie commotionis manus Domini exercituum quam ipse movebit super eam
ISA|19|17|et erit terra Iuda Aegypto in festivitatem omnis qui illius fuerit recordatus pavebit a facie consilii Domini exercituum quod ipse cogitavit super eam
ISA|19|18|in die illa erunt quinque civitates in terra Aegypti loquentes lingua Chanaan et iurantes per Dominum exercituum civitas Solis vocabitur una
ISA|19|19|in die illa erit altare Domini in medio terrae Aegypti et titulus iuxta terminum eius Domini
ISA|19|20|et erit in signum et in testimonium Domino exercituum in terra Aegypti clamabunt enim ad Dominum a facie tribulantis et mittet eis salvatorem et propugnatorem qui liberet eos
ISA|19|21|et cognoscetur Dominus ab Aegypto et cognoscent Aegyptii Dominum in die illa et colent eum in hostiis et muneribus et vota vovebunt Domino et solvent
ISA|19|22|et percutiet Dominus Aegyptum plaga et sanabit eam et revertentur ad Dominum et placabitur eis et sanabit eos
ISA|19|23|in die illa erit via de Aegypto in Assyrios et intrabit Assyrius Aegyptum et Aegyptius in Assyrios et servient Aegyptii Assur
ISA|19|24|in die illa erit Israhel tertius Aegyptio et Assyrio benedictio in medio terrae
ISA|19|25|cui benedixit Dominus exercituum dicens benedictus populus meus Aegypti et opus manuum mearum Assyrio hereditas autem mea Israhel
ISA|20|1|in anno quo ingressus est Tharthan in Azotum cum misisset eum Sargon rex Assyriorum et pugnasset contra Azotum et cepisset eam
ISA|20|2|in tempore illo locutus est Dominus in manu Isaiae filii Amos dicens vade et solve saccum de lumbis tuis et calciamenta tua tolle de pedibus tuis et fecit sic vadens nudus et disculciatus
ISA|20|3|et dixit Dominus sicut ambulavit servus meus Isaias nudus et disculciatus trium annorum signum et portentum erit super Aegyptum et super Aethiopiam
ISA|20|4|sic minabit rex Assyriorum captivitatem Aegypti et transmigrationem Aethiopiae iuvenum et senum nudam et disculciatam discopertis natibus ignominiam Aegypti
ISA|20|5|et timebunt et confundentur ab Aethiopia spe sua et ab Aegypto gloria sua
ISA|20|6|et dicet habitator insulae huius in die illa ecce haec erat spes nostra ad quos confugimus in auxilium ut liberaret nos a facie regis Assyriorum et quomodo effugere poterimus nos
ISA|21|1|onus deserti maris sicut turbines ab africo veniunt de deserto venit de terra horribili
ISA|21|2|visio dura nuntiata est mihi qui incredulus est infideliter agit et qui depopulator est vastat ascende Aelam obside Mede omnem gemitum eius cessare feci
ISA|21|3|propterea repleti sunt lumbi mei dolore angustia possedit me sicut angustia parientis corrui cum audirem conturbatus sum cum viderem
ISA|21|4|emarcuit cor meum tenebrae stupefecerunt me Babylon dilecta mea posita est mihi in miraculum
ISA|21|5|pone mensam contemplare in specula comedentes bibentes surgite principes arripite clypeum
ISA|21|6|haec enim dixit mihi Dominus vade et pone speculatorem et quodcumque viderit adnuntiet
ISA|21|7|et vidit currum duorum equitum ascensorem asini et ascensorem cameli et contemplatus est diligenter multo intuitu
ISA|21|8|et clamavit leo super specula Domini ego sum stans iugiter per diem et super custodiam meam ego sum stans totis noctibus
ISA|21|9|ecce iste venit ascensor vir bigae equitum et respondit et dixit cecidit cecidit Babylon et omnia sculptilia deorum eius contrita sunt in terram
ISA|21|10|tritura mea et fili areae meae quae audivi a Domino exercituum Deo Israhel adnuntiavi vobis
ISA|21|11|onus Duma ad me clamat ex Seir custos quid de nocte custos quid de nocte
ISA|21|12|dixit custos venit mane et nox si quaeritis quaerite convertimini venite
ISA|21|13|onus in Arabia in saltu ad vesperam dormietis in semitis Dodanim
ISA|21|14|occurrentes sitienti ferte aquam qui habitatis terram austri cum panibus occurrite fugienti
ISA|21|15|a facie enim gladiorum fugerunt a facie gladii inminentis a facie arcus extenti a facie gravis proelii
ISA|21|16|quoniam haec dicit Dominus ad me adhuc in uno anno quasi in anno mercennarii et auferetur omnis gloria Cedar
ISA|21|17|et reliquiae numeri sagittariorum fortium de filiis Cedar inminuentur Dominus enim Deus Israhel locutus est
ISA|22|1|onus vallis Visionis quidnam tibi quoque est quia ascendisti et tu omnis in tecta
ISA|22|2|clamoris plena urbs frequens civitas exultans interfecti tui non interfecti gladio nec mortui in bello
ISA|22|3|cuncti principes tui fugerunt simul dureque ligati sunt omnes qui inventi sunt vincti sunt pariter procul fugerunt
ISA|22|4|propterea dixi recedite a me amare flebo nolite incumbere ut consolemini me super vastitate filiae populi mei
ISA|22|5|dies enim interfectionis et conculcationis et fletuum Domino Deo exercituum in valle Visionis scrutans murum et magnificus super montem
ISA|22|6|et Aelam sumpsit faretram currum hominis equitis et parietem nudavit clypeus
ISA|22|7|et erunt electae valles tuae plenae quadrigarum et equites ponent sedes suas in porta
ISA|22|8|et revelabitur operimentum Iudae et videbis in die illa armamentarium domus saltus
ISA|22|9|et scissuras civitatis David videbitis quia multiplicatae sunt et congregastis aquas piscinae inferioris
ISA|22|10|et domos Hierusalem numerastis et destruxistis domos ad muniendum murum
ISA|22|11|et lacum fecistis inter duos muros et aquam piscinae veteris et non suspexistis ad eum qui fecerat eam et operatorem eius de longe non vidistis
ISA|22|12|et vocavit Dominus Deus exercituum in die illa ad fletum et ad planctum ad calvitium et ad cingulum sacci
ISA|22|13|et ecce gaudium et laetitia occidere vitulos et iugulare arietes comedere carnes et bibere vinum comedamus et bibamus cras enim moriemur
ISA|22|14|et revelata est in auribus meis Domini exercituum si dimittetur iniquitas haec vobis donec moriamini dicit Dominus Deus exercituum
ISA|22|15|haec dicit Dominus Deus exercituum vade ingredere ad eum qui habitat in tabernaculo ad Sobnam praepositum templi
ISA|22|16|quid tu hic aut quasi quis hic quia excidisti tibi hic sepulchrum excidisti in excelso memoriam diligenter in petra tabernaculum tibi
ISA|22|17|ecce Dominus asportari te faciet sicut asportatur gallus gallinacius et quasi amictum sic sublevabit te
ISA|22|18|coronans coronabit te tribulatione quasi pilam mittet te in terram latam et spatiosam ibi morieris et ibi erit currus gloriae tuae ignominia domus Domini tui
ISA|22|19|et expellam te de statione tua et de ministerio tuo deponam te
ISA|22|20|et erit in die illa vocabo servum meum Eliachim filium Helciae
ISA|22|21|et induam illum tunicam tuam et cingulo tuo confortabo eum et potestatem tuam dabo in manu eius et erit quasi pater habitantibus Hierusalem et domui Iuda
ISA|22|22|et dabo clavem domus David super umerum eius et aperiet et non erit qui claudat et claudet et non erit qui aperiat
ISA|22|23|et figam illum paxillum in loco fideli et erit in solium gloriae domui patris sui
ISA|22|24|et suspendent super eum omnem gloriam domus patris eius vasorum diversa genera omne vas parvulum a vasis craterarum usque ad omne vas musicorum
ISA|22|25|in die illo dicit Dominus exercituum auferetur paxillus qui fixus fuerat in loco fideli et frangetur et cadet et peribit quod pependerat in eo quia Dominus locutus est
ISA|23|1|onus Tyri ululate naves maris quia vastata est domus unde venire consueverant de terra Cetthim revelatum est eis
ISA|23|2|tacete qui habitatis in insula negotiatio Sidonis transfretantes mare repleverunt te
ISA|23|3|in aquis multis semen Nili messis fluminis fruges eius et facta est negotiatio gentium
ISA|23|4|erubesce Sidon ait enim mare fortitudo maris dicens non parturivi et non peperi et non enutrivi iuvenes nec ad incrementum perduxi virgines
ISA|23|5|cum auditum fuerit in Aegypto dolebunt cum audierint de Tyro
ISA|23|6|transite maria ululate qui habitatis in insula
ISA|23|7|numquid non haec vestra est quae gloriabatur a diebus pristinis in antiquitate sua ducent eam pedes sui longe ad peregrinandum
ISA|23|8|quis cogitavit hoc super Tyrum quondam coronatam cuius negotiatores principes institores eius incliti terrae
ISA|23|9|Dominus exercituum cogitavit hoc ut detraheret superbiam omnis gloriae et ad ignominiam deduceret universos inclitos terrae
ISA|23|10|transi terram tuam quasi flumen filia maris non est cingulum ultra tibi
ISA|23|11|manum suam extendit super mare conturbavit regna Dominus mandavit adversum Chanaan ut contereret fortes eius
ISA|23|12|et dixit non adicies ultra ut glorieris calumniam sustinens virgo filia Sidonis in Cetthim consurgens transfreta ibi quoque non erit requies tibi
ISA|23|13|ecce terra Chaldeorum talis populus non fuit Assur fundavit eam in captivitatem transduxerunt robustos eius suffoderunt domos eius posuerunt eam in ruinam
ISA|23|14|ululate naves maris quia devastata est fortitudo vestra
ISA|23|15|et erit in die illa in oblivione eris o Tyre septuaginta annis sicut dies regis unius post septuaginta autem annos erit Tyro quasi canticum meretricis
ISA|23|16|sume citharam circui civitatem meretrix oblivioni tradita bene cane frequenta canticum ut memoria tui sit
ISA|23|17|et erit post septuaginta annos visitabit Dominus Tyrum et reducet eam ad mercedes suas et rursum fornicabitur cum universis regnis terrae super faciem terrae
ISA|23|18|et erunt negotiatio eius et mercedes eius sanctificatae Domino non condentur neque reponentur quia his qui habitaverint coram Domino erit negotiatio eius ut manducent in saturitatem et vestiantur usque ad vetustatem
ISA|24|1|ecce Dominus dissipabit terram et nudabit eam et adfliget faciem eius et disperget habitatores eius
ISA|24|2|et erit sicut populus sic sacerdos et sicut servus sic dominus eius sicut ancilla sic domina eius sicut emens sic ille qui vendit sicut fenerator sic is qui mutuum accipit sicut qui repetit sic qui debet
ISA|24|3|dissipatione dissipabitur terra et direptione praedabitur Dominus enim locutus est verbum hoc
ISA|24|4|luxit et defluxit terra et infirmata est defluxit orbis infirmata est altitudo populi terrae
ISA|24|5|et terra interfecta est ab habitatoribus suis quia transgressi sunt leges mutaverunt ius dissipaverunt foedus sempiternum
ISA|24|6|propter hoc maledictio vorabit terram et peccabunt habitatores eius ideoque insanient cultores eius et relinquentur homines pauci
ISA|24|7|luxit vindemia infirmata est vitis ingemuerunt omnes qui laetabantur corde
ISA|24|8|cessavit gaudium tympanorum quievit sonitus laetantium conticuit dulcedo citharae
ISA|24|9|cum cantico non bibent vinum amara erit potio bibentibus illam
ISA|24|10|adtrita est civitas vanitatis clausa est omnis domus nullo introeunte
ISA|24|11|clamor erit super vino in plateis deserta est omnis laetitia translatum est gaudium terrae
ISA|24|12|relicta est in urbe solitudo et calamitas opprimet portas
ISA|24|13|quia haec erunt in medio terrae in medio populorum quomodo si paucae olivae quae remanserunt excutiantur ex olea et racemi cum fuerit finita vindemia
ISA|24|14|hii levabunt vocem suam atque laudabunt cum glorificatus fuerit Dominus hinnient de mari
ISA|24|15|propter hoc in doctrinis glorificate Dominum in insulis maris nomen Domini Dei Israhel
ISA|24|16|a finibus terrae laudes audivimus gloriam iusti et dixi secretum meum mihi secretum meum mihi vae mihi praevaricantes praevaricati sunt et praevaricatione transgressorum praevaricati sunt
ISA|24|17|formido et fovea et laqueus super te qui habitator es terrae
ISA|24|18|et erit qui fugerit a voce formidinis cadet in foveam et qui se explicuerit de fovea tenebitur laqueo quia cataractae de excelsis apertae sunt et concutientur fundamenta terrae
ISA|24|19|confractione confringetur terra contritione conteretur terra commotione commovebitur terra
ISA|24|20|agitatione agitabitur terra sicut ebrius et auferetur quasi tabernaculum unius noctis et gravabit eam iniquitas sua et corruet et non adiciet ut resurgat
ISA|24|21|et erit in die illa visitabit Dominus super militiam caeli in excelso et super reges terrae qui sunt super terram
ISA|24|22|et congregabuntur in congregationem unius fascis in lacum et cludentur ibi in carcerem et post multos dies visitabuntur
ISA|24|23|et erubescet luna et confundetur sol cum regnaverit Dominus exercituum in monte Sion et in Hierusalem et in conspectu senum suorum fuerit glorificatus
ISA|25|1|Domine Deus meus es tu exaltabo te confitebor nomini tuo quoniam fecisti mirabilia cogitationes antiquas fideles amen
ISA|25|2|quia posuisti civitatem in tumulum urbem fortem in ruinam domum alienorum ut non sit civitas et in sempiternum non aedificetur
ISA|25|3|super hoc laudabit te populus fortis civitas gentium robustarum timebit te
ISA|25|4|quia factus es fortitudo pauperi fortitudo egeno in tribulatione sua spes a turbine umbraculum ab aestu spiritus enim robustorum quasi turbo inpellens parietem
ISA|25|5|sicut aestum in siti tumultum alienorum humiliabis et quasi calore sub nube torrente propaginem fortium marcescere facies
ISA|25|6|et faciet Dominus exercituum omnibus populis in monte hoc convivium pinguium convivium vindemiae pinguium medullatorum vindemiae defecatae
ISA|25|7|et praecipitabit in monte isto faciem vinculi conligati super omnes populos et telam quam orditus est super universas nationes
ISA|25|8|praecipitabit mortem in sempiternum et auferet Dominus Deus lacrimam ab omni facie et obprobrium populi sui auferet de universa terra quia Dominus locutus est
ISA|25|9|et dicet in die illa ecce Deus noster iste expectavimus eum et salvabit nos iste Dominus sustinuimus eum exultabimus et laetabimur in salutari eius
ISA|25|10|quia requiescet manus Domini in monte isto et triturabitur Moab sub eo sicuti teruntur paleae in plaustro
ISA|25|11|et extendet manus suas sub eo sicut extendit natans ad natandum et humiliabit gloriam eius cum adlisione manuum eius
ISA|25|12|et munimenta sublimium murorum tuorum concident et humiliabuntur et detrahentur in terram usque ad pulverem
ISA|26|1|in die illa cantabitur canticum istud in terra Iuda urbs fortitudinis nostrae salvator ponetur in ea murus et antemurale
ISA|26|2|aperite portas et ingrediatur gens iusta custodiens veritatem
ISA|26|3|vetus error abiit servabis pacem pacem quia in te speravimus
ISA|26|4|sperastis in Domino in saeculis aeternis in Domino Deo forti in perpetuum
ISA|26|5|quia incurvabit habitantes in excelso civitatem sublimem humiliabit humiliabit eam usque ad terram detrahet eam usque ad pulverem
ISA|26|6|conculcabit eam pes pedes pauperis gressus egenorum
ISA|26|7|semita iusti recta est rectus callis iusti ad ambulandum
ISA|26|8|et in semita iudiciorum tuorum Domine sustinuimus te nomen tuum et memoriale tuum in desiderio animae
ISA|26|9|anima mea desideravit te in nocte sed et spiritu meo in praecordiis meis de mane vigilabo ad te cum feceris iudicia tua in terra iustitiam discent habitatores orbis
ISA|26|10|misereamur impio et non discet iustitiam in terra sanctorum inique gessit et non videbit gloriam Domini
ISA|26|11|Domine exaltetur manus tua et non videant videant et confundantur zelantes populi et ignis hostes tuos devoret
ISA|26|12|Domine dabis pacem nobis omnia enim opera nostra operatus es nobis
ISA|26|13|Domine Deus noster possederunt nos domini absque te tantum in te recordemur nominis tui
ISA|26|14|morientes non vivant gigantes non resurgant propterea visitasti et contrivisti eos et perdidisti omnem memoriam eorum
ISA|26|15|indulsisti genti Domine indulsisti genti numquid glorificatus es elongasti omnes terminos terrae
ISA|26|16|Domine in angustia requisierunt te in tribulatione murmuris doctrina tua eis
ISA|26|17|sicut quae concipit cum adpropinquaverit ad partum dolens clamat in doloribus suis sic facti sumus a facie tua Domine
ISA|26|18|concepimus et quasi parturivimus et peperimus spiritum salutes non fecimus in terra ideo non ceciderunt habitatores terrae
ISA|26|19|vivent mortui tui interfecti mei resurgent expergiscimini et laudate qui habitatis in pulvere quia ros lucis ros tuus et terram gigantum detrahes in ruinam
ISA|26|20|vade populus meus intra in cubicula tua claude ostia tua super te abscondere modicum ad momentum donec pertranseat indignatio
ISA|26|21|ecce enim Dominus egreditur de loco suo ut visitet iniquitatem habitatoris terrae contra eum et revelabit terra sanguinem suum et non operiet ultra interfectos suos
ISA|27|1|in die illo visitabit Dominus in gladio suo duro et grandi et forti super Leviathan serpentem vectem et super Leviathan serpentem tortuosum et occidet cetum qui in mari est
ISA|27|2|in die illa vinea meri cantabit ei
ISA|27|3|ego Dominus qui servo eam repente propinabo ei ne forte visitetur contra eam nocte et die servo eam
ISA|27|4|indignatio non est mihi quis dabit me spinam et veprem in proelio gradiar super eam succendam eam pariter
ISA|27|5|an potius tenebit fortitudinem meam faciet pacem mihi pacem faciet mihi
ISA|27|6|qui egrediuntur impetu ad Iacob florebit et germinabit Israhel et implebunt faciem orbis semine
ISA|27|7|numquid iuxta plagam percutientis se percussit eum aut sicut occidit interfectos eius sic occisus est
ISA|27|8|in mensura contra mensuram cum abiecta fuerit iudicabis eam meditata est in spiritu suo duro per diem aestus
ISA|27|9|idcirco super hoc dimittetur iniquitas domui Iacob et iste omnis fructus ut auferatur peccatum eius cum posuerit omnes lapides altaris sicut lapides cineris adlisos non stabunt luci et delubra
ISA|27|10|civitas enim munita desolata erit speciosa relinquetur et dimittetur quasi desertum ibi pascetur vitulus et ibi accubabit et consumet summitates eius
ISA|27|11|in siccitate messis illius conterentur mulieres venientes et docentes eam non est enim populus sapiens propterea non miserebitur eius qui fecit eum et qui formavit eum non parcet ei
ISA|27|12|et erit in die illa percutiet Dominus ab alveo Fluminis usque ad torrentem Aegypti et vos congregabimini unus et unus filii Israhel
ISA|27|13|et erit in die illa clangetur in tuba magna et venient qui perditi fuerant de terra Assyriorum et qui eiecti erant in terra Aegypti et adorabunt Dominum in monte sancto in Hierusalem
ISA|28|1|vae coronae superbiae ebriis Ephraim et flori decidenti gloriae exultationis eius qui erant in vertice vallis pinguissimae errantes a vino
ISA|28|2|ecce validus et fortis Domini sicut impetus grandinis turbo confringens sicut impetus aquarum multarum inundantium et emissarum super terram spatiosam
ISA|28|3|pedibus conculcabitur corona superbiae ebriorum Ephraim
ISA|28|4|et erit flos decidens gloriae exultationis eius qui est super verticem vallis pinguium quasi temporaneum ante maturitatem autumni quod cum aspexerit videns statim ut manu tenuerit devorabit illud
ISA|28|5|in die illa erit Dominus exercituum corona gloriae et sertum exultationis residuo populi sui
ISA|28|6|et spiritus iudicii sedenti super iudicium et fortitudo revertentibus de bello ad portam
ISA|28|7|verum hii quoque prae vino nescierunt et prae ebrietate erraverunt sacerdos et propheta nescierunt prae ebrietate absorti sunt a vino erraverunt in ebrietate nescierunt videntem ignoraverunt iudicium
ISA|28|8|omnes enim mensae repletae sunt vomitu sordiumque ita ut non esset ultra locus
ISA|28|9|quem docebit scientiam et quem intellegere faciet auditum ablactatos a lacte apulsos ab uberibus
ISA|28|10|quia manda remanda manda remanda expecta reexpecta expecta reexpecta modicum ibi modicum ibi
ISA|28|11|in loquella enim labii et lingua altera loquetur ad populum istum
ISA|28|12|cui dixit haec requies reficite lassum et hoc est meum refrigerium et noluerunt audire
ISA|28|13|et erit eis verbum Domini manda remanda manda remanda expecta reexpecta expecta reexpecta modicum ibi modicum ibi ut vadant et cadant retrorsum et conterantur et inlaqueentur et capiantur
ISA|28|14|propter hoc audite verbum Domini viri inlusores qui dominamini super populum meum qui est in Hierusalem
ISA|28|15|dixistis enim percussimus foedus cum morte et cum inferno fecimus pactum flagellum inundans cum transierit non veniet super nos quia posuimus mendacium spem nostram et mendacio protecti sumus
ISA|28|16|idcirco haec dicit Dominus Deus ecce ego mittam in fundamentis Sion lapidem lapidem probatum angularem pretiosum in fundamento fundatum qui crediderit non festinet
ISA|28|17|et ponam iudicium in pondere et iustitiam in mensura et subvertet grando spem mendacii et protectionem aquae inundabunt
ISA|28|18|et delebitur foedus vestrum cum morte et pactum vestrum cum inferno non stabit flagellum inundans cum transierit eritis ei in conculcationem
ISA|28|19|quandocumque pertransierit tollet vos quoniam mane diluculo pertransibit in die et in nocte et tantummodo sola vexatio intellectum dabit auditui
ISA|28|20|coangustatum est enim stratum ita ut alter decidat et pallium breve utrumque operire non potest
ISA|28|21|sicut enim in monte Divisionum stabit Dominus sicut in valle quae est in Gabao irascetur ut faciat opus suum alienum opus eius ut operetur opus suum peregrinum est opus ab eo
ISA|28|22|et nunc nolite inludere ne forte constringantur vincula vestra consummationem enim et adbreviationem audivi a Domino Deo exercituum super universam terram
ISA|28|23|auribus percipite et audite vocem meam adtendite et audite eloquium meum
ISA|28|24|numquid tota die arabit arans ut serat proscindet et sariet humum suam
ISA|28|25|nonne cum adaequaverit faciem eius seret gith et cyminum sparget et ponet triticum per ordinem et hordeum et milium et viciam in finibus suis
ISA|28|26|et erudiet eum illud in iudicio Deus suus docebit eum illud
ISA|28|27|non enim in serris triturabitur gith nec rota plaustri super cyminum circumiet sed in virga excutietur gith et cyminum in baculo
ISA|28|28|panis autem comminuetur verum non in perpetuum triturans triturabit illum neque vexabit eum rota plaustri nec in ungulis suis comminuet eum
ISA|28|29|et hoc a Domino Deo exercituum exivit ut mirabile faceret consilium et magnificaret iustitiam
ISA|29|1|vae Arihel Arihel civitas quam circumdedit David additus est annus ad annum sollemnitates evolutae sunt
ISA|29|2|et circumvallabo Arihel et erit tristis et maerens et erit mihi quasi Arihel
ISA|29|3|et circumdabo quasi spheram in circuitu tuo et iaciam contra te aggerem et munimenta ponam in obsidionem tuam
ISA|29|4|humiliaberis de terra loqueris et de humo audietur eloquium tuum et erit quasi pythonis de terra vox tua et de humo eloquium tuum mussitabit
ISA|29|5|et erit sicut pulvis tenuis multitudo ventilantium te et sicut favilla pertransiens multitudo eorum qui contra te praevaluerunt
ISA|29|6|eritque repente confestim a Domino exercituum visitabitur in tonitru et commotione terrae et voce magna turbinis et tempestatis et flammae ignis devorantis
ISA|29|7|et erit sicut somnium visionis nocturnae multitudo omnium gentium quae dimicaverunt contra Arihel et omnes qui militaverunt et obsederunt et praevaluerunt adversus eam
ISA|29|8|et sicuti somniat esuriens et comedit cum autem fuerit expertus vacua est anima eius et sicut somniat sitiens et bibit et postquam fuerit expergefactus lassus adhuc sitit et anima eius vacua est sic erit multitudo omnium gentium quae dimicaverunt contra montem Sion
ISA|29|9|obstupescite et admiramini fluctuate et vacillate inebriamini et non a vino movemini et non ebrietate
ISA|29|10|quoniam miscuit vobis Dominus spiritum soporis claudet oculos vestros prophetas et principes vestros qui vident visiones operiet
ISA|29|11|et erit vobis visio omnium sicut verba libri signati quem cum dederint scienti litteras dicent lege istum et respondebit non possum signatus est enim
ISA|29|12|et dabitur liber nescienti litteras diceturque ei lege et respondebit nescio litteras
ISA|29|13|et dixit Dominus eo quod adpropinquat populus iste ore suo et labiis suis glorificat me cor autem eius longe est a me et timuerunt me mandato hominum et doctrinis
ISA|29|14|ideo ecce ego addam ut admirationem faciam populo huic miraculo grandi et stupendo peribit enim sapientia a sapientibus eius et intellectus prudentium eius abscondetur
ISA|29|15|vae qui profundi estis corde ut a Domino abscondatis consilium quorum sunt in tenebris opera et dicunt quis videt nos et quis novit nos
ISA|29|16|perversa est haec vestra cogitatio quasi lutum contra figulum cogitet et dicat opus factori suo non fecisti me et figmentum dicat fictori suo non intellegis
ISA|29|17|nonne adhuc in modico et in brevi convertetur Libanus in Chermel et Chermel in saltum reputabitur
ISA|29|18|et audient in die illa surdi verba libri et de tenebris et caligine oculi caecorum videbunt
ISA|29|19|et addent mites in Domino laetitiam et pauperes homines in Sancto Israhel exultabunt
ISA|29|20|quoniam defecit qui praevalebat consummatus est inlusor et succisi sunt omnes qui vigilabant super iniquitatem
ISA|29|21|qui peccare faciebant homines in verbo et arguentem in porta subplantabant et declinaverunt frustra a iusto
ISA|29|22|propter hoc haec dicit Dominus ad domum Iacob qui redemit Abraham non modo confundetur Iacob nec modo vultus eius erubescet
ISA|29|23|sed cum viderit filios suos opera manuum mearum in medio sui sanctificantes nomen meum et sanctificabunt Sanctum Iacob et Deum Israhel praedicabunt
ISA|29|24|et scient errantes spiritu intellectum et mussitatores discent legem
ISA|30|1|vae filii desertores dicit Dominus ut faceretis consilium et non ex me et ordiremini telam et non per spiritum meum ut adderetur peccatum super peccatum
ISA|30|2|qui ambulatis ut descendatis in Aegyptum et os meum non interrogastis sperantes auxilium in fortitudine Pharao et habentes fiduciam in umbra Aegypti
ISA|30|3|et erit vobis fortitudo Pharaonis in confusionem et fiducia umbrae Aegypti in ignominiam
ISA|30|4|erant enim in Tanis principes tui et nuntii tui usque ad Anes pervenerunt
ISA|30|5|omnes confusi sunt super populo qui eis prodesse non potuit non fuerunt in auxilium et in aliquam utilitatem sed in confusionem et obprobrium
ISA|30|6|onus iumentorum austri in terra tribulationis et angustiae leaena et leo ex eis vipera et regulus volans portantes super umeros iumentorum divitias suas et super gibbum camelorum thesauros suos ad populum qui eis prodesse non poterit
ISA|30|7|Aegyptus enim frustra et vane auxiliabitur ideo clamavi super hoc superbia tantum est quiesce
ISA|30|8|nunc ingressus scribe eis super buxum et in libro diligenter exara illud et erit in die novissimo in testimonium usque ad aeternum
ISA|30|9|populus enim ad iracundiam provocans est et filii mendaces filii nolentes audire legem Domini
ISA|30|10|qui dicunt videntibus nolite videre et aspicientibus nolite aspicere nobis ea quae recta sunt loquimini nobis placentia videte nobis errores
ISA|30|11|auferte a me viam declinate a me semitam cesset a facie nostra Sanctus Israhel
ISA|30|12|propterea haec dicit Sanctus Israhel pro eo quod reprobastis verbum hoc et sperastis in calumniam et tumultum et innixi estis super eo
ISA|30|13|propterea erit vobis iniquitas haec sicut interruptio cadens et requisita in muro excelso quoniam subito dum non speratur veniet contritio eius
ISA|30|14|et comminuetur sicut conteritur lagoena figuli contritione pervalida et non invenietur de fragmentis eius testa in qua portetur igniculus de incendio aut hauriatur parum aquae de fovea
ISA|30|15|quia haec dicit Dominus Deus Sanctus Israhel si revertamini et quiescatis salvi eritis in silentio et in spe erit fortitudo vestra et noluistis
ISA|30|16|et dixistis nequaquam sed ad equos fugiemus ideo fugietis et super veloces ascendemus ideo veloces erunt qui persequentur vos
ISA|30|17|mille homines a facie terroris unius et a facie terroris quinque fugietis donec relinquamini quasi malus navis in vertice montis et quasi signum super collem
ISA|30|18|propterea expectat Dominus ut misereatur vestri et ideo exaltabitur parcens vobis quia Deus iudicii Dominus beati omnes qui expectant eum
ISA|30|19|populus enim Sion habitabit in Hierusalem plorans nequaquam plorabis miserans miserebitur tui ad vocem clamoris tui statim ut audierit respondebit tibi
ISA|30|20|et dabit vobis Dominus panem artum et aquam brevem et non faciet avolare a te ultra doctorem tuum et erunt oculi tui videntes praeceptorem tuum
ISA|30|21|et aures tuae audient verbum post tergum monentis haec via ambulate in ea neque ad dexteram neque ad sinistram
ISA|30|22|et contaminabis lamminas sculptilium argenti tui et vestimentum conflatilis auri tui et disperges ea sicut inmunditiam menstruatae egredere dices ei
ISA|30|23|et dabitur pluvia semini tuo ubicumque seminaveris in terra et panis frugum terrae erit uberrimus et pinguis pascetur in possessione tua in die illo agnus spatiose
ISA|30|24|et tauri tui et pulli asinorum qui operantur terram commixtum migma comedent sic in area ut ventilatum est
ISA|30|25|et erunt super omnem montem excelsum et super omnem collem elevatum rivi currentium aquarum in die interfectionis multorum cum ceciderint turres
ISA|30|26|et erit lux lunae sicut lux solis et lux solis erit septempliciter sicut lux septem dierum in die qua alligaverit Dominus vulnus populi sui et percussuram plagae eius sanaverit
ISA|30|27|ecce nomen Domini venit de longinquo ardens furor eius et gravis ad portandum labia eius repleta sunt indignatione et lingua eius quasi ignis devorans
ISA|30|28|spiritus eius velut torrens inundans usque ad medium colli ad perdendas gentes in nihilum et frenum erroris quod erat in maxillis populorum
ISA|30|29|canticum erit vobis sicut nox sanctificatae sollemnitatis et laetitia cordis sicut qui pergit cum tibia ut intret in montem Domini ad Fortem Israhel
ISA|30|30|et auditam faciet Dominus gloriam vocis suae et terrorem brachii sui ostendet in comminatione furoris et flamma ignis devorantis adlidet in turbine et in lapide grandinis
ISA|30|31|a voce enim Domini pavebit Assur virga percussus
ISA|30|32|et erit transitus virgae fundatus quam requiescere faciet Dominus super eum in tympanis et in citharis et in bellis praecipuis expugnabit eos
ISA|30|33|praeparata est enim ab heri Thofeth a rege praeparata profunda et dilatata nutrimenta eius ignis et ligna multa flatus Domini sicut torrens sulphuris succendens eam
ISA|31|1|vae qui descendunt in Aegyptum ad auxilium in equis sperantes et habentes fiduciam super quadrigis quia multae sunt et super equitibus quia praevalidi nimis et non sunt confisi super Sanctum Israhel et Dominum non requisierunt
ISA|31|2|ipse autem sapiens adduxit malum et verba sua non abstulit et consurget contra domum pessimorum et contra auxilium operantium iniquitatem
ISA|31|3|Aegyptus homo et non deus et equi eorum caro et non spiritus et Dominus inclinabit manum suam et corruet auxiliator et cadet cui praestatur auxilium simulque omnes consumentur
ISA|31|4|quia haec dicit Dominus ad me quomodo si rugiat leo et catulus leonis super praedam suam cum occurrerit ei multitudo pastorum a voce eorum non formidabit et a multitudine eorum non pavebit sic descendet Dominus exercituum ut proelietur super montem Sion et super collem eius
ISA|31|5|sicut aves volantes sic proteget Dominus exercituum Hierusalem protegens et liberans transiens et salvans
ISA|31|6|convertimini sicut in profundum recesseratis filii Israhel
ISA|31|7|in die enim illa abiciet vir idola argenti sui et idola auri sui quae fecerunt vobis manus vestrae in peccatum
ISA|31|8|et cadet Assur in gladio non viri et gladius non hominis vorabit eum et fugiet non a facie gladii et iuvenes eius vectigales erunt
ISA|31|9|et fortitudo eius a terrore transibit et pavebunt fugientes principes eius dixit Dominus cuius ignis est in Sion et caminus eius in Hierusalem
ISA|32|1|ecce in iustitia regnabit rex et principes in iudicio praeerunt
ISA|32|2|et erit vir sicut qui absconditur a vento et celat se a tempestate sicut rivi aquarum in siti et umbra petrae prominentis in terra deserta
ISA|32|3|non caligabunt oculi videntium et aures audientium diligenter auscultabunt
ISA|32|4|et cor stultorum intelleget scientiam et lingua balborum velociter loquetur et plane
ISA|32|5|non vocabitur ultra is qui insipiens est princeps neque fraudulentus appellabitur maior
ISA|32|6|stultus enim fatua loquetur et cor eius faciet iniquitatem ut perficiat simulationem et loquatur ad Dominum fraudulenter et vacuefaciat animam esurientis et potum sitienti auferat
ISA|32|7|fraudulenti vasa pessima sunt ipse enim cogitationes concinnavit ad perdendos mites in sermone mendacii cum loqueretur pauper iudicium
ISA|32|8|princeps vero ea quae digna sunt principe cogitavit et ipse super duces stabit
ISA|32|9|mulieres opulentae surgite et audite vocem meam filiae confidentes percipite auribus eloquium meum
ISA|32|10|post dies et annum et vos conturbabimini confidentes consummata est enim vindemia collectio ultra non veniet
ISA|32|11|obstupescite opulentae conturbamini confidentes exuite vos et confundimini accingite lumbos vestros
ISA|32|12|super ubera plangite super regione desiderabili super vinea fertili
ISA|32|13|super humum populi mei spina et vepres ascendent quanto magis super omnes domos gaudii civitatis exultantis
ISA|32|14|domus enim dimissa est multitudo urbis relicta est tenebrae et palpatio factae sunt super speluncas usque in aeternum gaudium onagrorum pascua gregum
ISA|32|15|donec effundatur super nos spiritus de excelso et erit desertum in Chermel et Chermel in saltum reputabitur
ISA|32|16|et habitabit in solitudine iudicium et iustitia in Chermel sedebit
ISA|32|17|et erit opus iustitiae pax et cultus iustitiae silentium et securitas usque in sempiternum
ISA|32|18|et sedebit populus meus in pulchritudine pacis et in tabernaculis fiduciae et in requie opulenta
ISA|32|19|grando autem in descensione saltus et humilitate humiliabitur civitas
ISA|32|20|beati qui seminatis super omnes aquas inmittentes pedem bovis et asini
ISA|33|1|vae qui praedaris nonne et ipse praedaberis et qui spernis nonne et ipse sperneris cum consummaveris depraedationem depraedaberis cum fatigatus desiveris contemnere contemneris
ISA|33|2|Domine miserere nostri te expectavimus esto brachium eorum in mane et salus nostra in tempore tribulationis
ISA|33|3|a voce angeli fugerunt populi ab exaltatione tua dispersae sunt gentes
ISA|33|4|et congregabuntur spolia vestra sicut colligitur brucus velut cum fossae plenae fuerint de eo
ISA|33|5|magnificatus est Dominus quoniam habitavit in excelso implevit Sion iudicio et iustitia
ISA|33|6|et erit fides in temporibus tuis divitiae salutis sapientia et scientia timor Domini ipse thesaurus eius
ISA|33|7|ecce videntes clamabunt foris angeli pacis amare flebunt
ISA|33|8|dissipatae sunt viae cessavit transiens per semitam irritum factum est pactum proiecit civitates non reputavit homines
ISA|33|9|luxit et elanguit terra confusus est Libanus et obsorduit et factus est Saron sicut desertum et concussa est Basan et Carmelus
ISA|33|10|nunc consurgam dicit Dominus nunc exaltabor nunc sublevabor
ISA|33|11|concipietis ardorem parietis stipulam spiritus vester ut ignis vorabit vos
ISA|33|12|et erunt populi quasi de incendio cinis spinae congregatae igni conburentur
ISA|33|13|audite qui longe estis quae fecerim et cognoscite vicini fortitudinem meam
ISA|33|14|conterriti sunt in Sion peccatores possedit tremor hypocritas quis poterit habitare de vobis cum igne devorante quis habitabit ex vobis cum ardoribus sempiternis
ISA|33|15|qui ambulat in iustitiis et loquitur veritates qui proicit avaritiam ex calumnia et excutit manus suas ab omni munere qui obturat aures suas ne audiat sanguinem et claudit oculos suos ne videat malum
ISA|33|16|iste in excelsis habitabit munimenta saxorum sublimitas eius panis ei datus est aquae eius fideles sunt
ISA|33|17|regem in decore suo videbunt oculi eius cernent terram de longe
ISA|33|18|cor tuum meditabitur timorem ubi est litteratus ubi legis verba ponderans ubi doctor parvulorum
ISA|33|19|populum inpudentem non videbis populum alti sermonis ita ut non possis intellegere disertitudinem linguae eius in quo nulla est sapientia
ISA|33|20|respice Sion civitatem sollemnitatis nostrae oculi tui videbunt Hierusalem habitationem opulentam tabernaculum quod nequaquam transferri poterit nec auferentur clavi eius in sempiternum et omnes funiculi eius non rumpentur
ISA|33|21|quia solummodo ibi magnificus Dominus noster locus fluviorum rivi latissimi et patentes non transibit per eum navis remigum neque trieris magna transgredietur eum
ISA|33|22|Dominus enim iudex noster Dominus legifer noster Dominus rex noster ipse salvabit nos
ISA|33|23|laxati sunt funiculi tui sed non praevalebunt sic erit malus tuus ut dilatare signum non queas tunc dividentur spolia praedarum multarum claudi diripient rapinam
ISA|33|24|nec dicet vicinus elangui populus qui habitat in ea auferetur ab eo iniquitas
ISA|34|1|accedite gentes et audite et populi adtendite audiat terra et plenitudo eius orbis et omne germen eius
ISA|34|2|quia indignatio Domini super omnes gentes et furor super universam militiam eorum interfecit eos et dedit eos in occisionem
ISA|34|3|interfecti eorum proicientur et de cadaveribus eorum ascendet fetor tabescent montes sanguine eorum
ISA|34|4|et tabescet omnis militia caelorum et conplicabuntur sicut liber caeli et omnis militia eorum defluet sicut defluit folium de vinea et de ficu
ISA|34|5|quoniam inebriatus est in caelo gladius meus ecce super Idumeam descendet et super populum interfectionis meae ad iudicium
ISA|34|6|gladius Domini repletus est sanguine incrassatus est adipe de sanguine agnorum et hircorum de sanguine medullatorum arietum victima enim Domini in Bosra et interfectio magna in terra Edom
ISA|34|7|et descendent unicornes cum eis et tauri cum potentibus inebriabitur terra eorum sanguine et humus eorum adipe pinguium
ISA|34|8|quia dies ultionis Domini annus retributionum iudicii Sion
ISA|34|9|et convertentur torrentes eius in picem et humus eius in sulphur et erit terra eius in picem ardentem
ISA|34|10|nocte et die non extinguetur in sempiternum ascendet fumus eius a generatione in generationem desolabitur in saeculum saeculorum non erit transiens per eam
ISA|34|11|et possidebunt illam onocrotalus et ericius et ibis et corvus habitabunt in ea et extendetur super eam mensura ut redigatur ad nihilum et perpendiculum in desolationem
ISA|34|12|nobiles eius non erunt ibi regem potius invocabunt et omnes principes eius erunt in nihilum
ISA|34|13|et orientur in domibus eius spinae et urticae et paliurus in munitionibus eius et erit cubile draconum et pascua strutionum
ISA|34|14|et occurrent daemonia onocentauris et pilosus clamabit alter ad alterum ibi cubavit lamia et invenit sibi requiem
ISA|34|15|ibi habuit foveam ericius et enutrivit catulos et circumfodit et fovit in umbra eius illuc congregati sunt milvi alter ad alterum
ISA|34|16|requirite diligenter in libro Domini et legite unum ex eis non defuit alter ad alterum non quaesivit quia quod ex ore meo procedit ille mandavit et spiritus eius ipse congregavit ea
ISA|34|17|et ipse misit eis sortem et manus eius divisit eam illis in mensuram usque in aeternum possidebunt eam in generatione et generatione habitabunt in ea
ISA|35|1|laetabitur deserta et invia et exultabit solitudo et florebit quasi lilium
ISA|35|2|germinans germinabit et exultabit laetabunda et laudans gloria Libani data est ei decor Carmeli et Saron ipsi videbunt gloriam Domini et decorem Dei nostri
ISA|35|3|confortate manus dissolutas et genua debilia roborate
ISA|35|4|dicite pusillanimis confortamini nolite timere ecce Deus vester ultionem adducet retributionis Deus ipse veniet et salvabit vos
ISA|35|5|tunc aperientur oculi caecorum et aures surdorum patebunt
ISA|35|6|tunc saliet sicut cervus claudus et aperta erit lingua mutorum quia scissae sunt in deserto aquae et torrentes in solitudine
ISA|35|7|et quae erat arida in stagnum et sitiens in fontes aquarum in cubilibus in quibus prius dracones habitabant orietur viror calami et iunci
ISA|35|8|et erit ibi semita et via et via sancta vocabitur non transibit per eam pollutus et haec erit nobis directa via ita ut stulti non errent per eam
ISA|35|9|non erit ibi leo et mala bestia non ascendet per eam nec invenietur ibi et ambulabunt qui liberati fuerint
ISA|35|10|et redempti a Domino convertentur et venient in Sion cum laude et laetitia sempiterna super caput eorum gaudium et laetitiam obtinebunt et fugiet dolor et gemitus
ISA|36|1|et factum est in quartodecimo anno regis Ezechiae ascendit Sennacherib rex Assyriorum super omnes civitates Iuda munitas et cepit eas
ISA|36|2|et misit rex Assyriorum Rabsacen de Lachis in Hierusalem ad regem Ezechiam in manu gravi et stetit in aquaeductu piscinae superioris in via agri Fullonis
ISA|36|3|et egressus est ad eum Eliachim filius Helciae qui erat super domum et Sobna scriba et Ioae filius Asaph a commentariis
ISA|36|4|et dixit ad eos Rabsaces dicite Ezechiae haec dicit rex magnus rex Assyriorum quae est ista fiducia qua confidis
ISA|36|5|aut quo consilio vel fortitudine rebellare disponis super quem habes fiduciam quia recessisti a me
ISA|36|6|ecce confidis super baculum harundineum confractum istum super Aegyptum cui si innisus fuerit homo intrabit in manu eius et perforabit eam sic Pharao rex Aegypti omnibus qui confidunt in eo
ISA|36|7|quod si responderis mihi in Domino Deo nostro confidimus nonne ipse est cuius abstulit Ezechias excelsa et altaria et dixit Iudae et Hierusalem coram altari isto adorabitis
ISA|36|8|et nunc trade te domino meo regi Assyriorum et dabo tibi duo milia equorum nec poteris ex te praebere ascensores eorum
ISA|36|9|et quomodo sustinebis faciem iudicis unius loci ex servis domini mei minoribus quod si confidis in Aegypto in quadriga et in equitibus
ISA|36|10|et nunc numquid sine Domino ascendi ad terram istam ut disperderem eam Dominus dixit ad me ascende super terram istam et disperde eam
ISA|36|11|et dixit Eliachim et Sobna et Ioae ad Rabsacen loquere ad servos tuos syra lingua intellegimus enim ne loquaris ad nos iudaice in auribus populi qui est super murum
ISA|36|12|et dixit ad eos Rabsaces numquid ad dominum tuum et ad te misit me dominus meus ut loquerer omnia verba ista et non potius ad viros qui sedent in muro ut comedant stercora sua et bibant urinam pedum suorum vobiscum
ISA|36|13|et stetit Rabsaces et clamavit voce magna iudaice et dixit audite verba regis magni regis Assyriorum
ISA|36|14|haec dicit rex non seducat vos Ezechias quia non poterit eruere vos
ISA|36|15|et non vobis tribuat fiduciam Ezechias super Domino dicens eruens liberabit nos Dominus non dabitur civitas ista in manu regis Assyriorum
ISA|36|16|nolite audire Ezechiam haec enim dicit rex Assyriorum facite mecum benedictionem et egredimini ad me et comedite unusquisque vineam suam et unusquisque ficum suam et bibite unusquisque aquam cisternae suae
ISA|36|17|donec veniam et tollam vos ad terram quae est ut terra vestra terram frumenti et vini terram panum et vinearum
ISA|36|18|ne conturbet vos Ezechias dicens Dominus liberabit nos numquid liberaverunt dii gentium unusquisque terram suam de manu regis Assyriorum
ISA|36|19|ubi est deus Emath et Arfad ubi est deus Seffarvaim numquid liberaverunt Samariam de manu mea
ISA|36|20|quis est ex omnibus diis terrarum istarum qui eruerit terram suam de manu mea ut eruat Dominus Hierusalem de manu mea
ISA|36|21|et siluerunt et non responderunt ei verbum mandaverat enim rex dicens ne respondeatis ei
ISA|36|22|et ingressus est Eliachim filius Helciae qui erat super domum et Sobna scriba et Ioae filius Asaph a commentariis ad Ezechiam scissis vestibus et nuntiaverunt ei verba Rabsacis
ISA|37|1|et factum est cum audisset rex Ezechias scidit vestimenta sua et obvolutus est sacco et intravit in domum Domini
ISA|37|2|et misit Eliachim qui erat super domum et Sobnam scribam et seniores de sacerdotibus opertos saccis ad Isaiam filium Amos prophetam
ISA|37|3|et dixerunt ad eum haec dicit Ezechias dies tribulationis et correptionis et blasphemiae dies haec quia venerunt filii usque ad partum et virtus non est parienti
ISA|37|4|si quo modo audiat Dominus Deus tuus verba Rabsaces quem misit rex Assyriorum dominus suus ad blasphemandum Deum viventem et obprobrandum sermonibus quos audivit Dominus Deus tuus leva ergo orationem pro reliquiis quae reppertae sunt
ISA|37|5|et venerunt servi regis Ezechiae ad Isaiam
ISA|37|6|et dixit ad eos Isaias haec dicetis domino vestro haec dicit Dominus ne timeas a facie verborum quae audisti quibus blasphemaverunt pueri regis Assyriorum me
ISA|37|7|ecce ego dabo ei spiritum et audiet nuntium et revertetur ad terram suam et corruere eum faciam gladio in terra sua
ISA|37|8|reversus est autem Rabsaces et invenit regem Assyriorum proeliantem adversus Lobna audierat enim quia profectus esset de Lachis
ISA|37|9|et audivit de Tharaca rege Aethiopiae dicentes egressus est ut pugnet contra te quod cum audisset misit nuntios ad Ezechiam dicens
ISA|37|10|haec dicetis Ezechiae regi Iudae loquentes non te decipiat Deus tuus in quo tu confidis dicens non dabitur Hierusalem in manu regis Assyriorum
ISA|37|11|ecce tu audisti omnia quae fecerunt reges Assyriorum omnibus terris quas subverterunt et tu poteris liberari
ISA|37|12|numquid eruerunt eos dii gentium quos subverterunt patres mei Gozan et Aran et Reseph et filios Eden qui erant in Thalassar
ISA|37|13|ubi est rex Emath et rex Arfad et rex urbis Seffarvaim Anahe et Ava
ISA|37|14|et tulit Ezechias libros de manu nuntiorum et legit eos et ascendit in domum Domini et expandit eos Ezechias coram Domino
ISA|37|15|et oravit Ezechias ad Dominum dicens
ISA|37|16|Domine exercituum Deus Israhel qui sedes super cherubin tu es Deus solus omnium regnorum terrae tu fecisti caelum et terram
ISA|37|17|inclina Domine aurem tuam et audi aperi Domine oculos tuos et vide et audi omnia verba Sennacherib quae misit ad blasphemandum Deum viventem
ISA|37|18|vere enim Domine desertas fecerunt reges Assyriorum terras et regiones earum
ISA|37|19|et dederunt deos earum igni non enim erant dii sed opera manuum hominum lignum et lapis et comminuerunt eos
ISA|37|20|et nunc Domine Deus noster salva nos de manu eius et cognoscant omnia regna terrae quia tu es Dominus solus
ISA|37|21|et misit Isaias filius Amos ad Ezechiam dicens haec dicit Dominus Deus Israhel pro quibus rogasti me de Sennacherib rege Assyriorum
ISA|37|22|hoc est verbum quod locutus est Dominus super eum despexit te subsannavit te virgo filia Sion post te caput movit filia Hierusalem
ISA|37|23|cui exprobrasti et quem blasphemasti et super quem exaltasti vocem et levasti altitudinem oculorum tuorum ad Sanctum Israhel
ISA|37|24|in manu servorum tuorum exprobrasti Domino et dixisti in multitudine quadrigarum mearum ego ascendi altitudinem montium iuga Libani et succidam excelsa cedrorum eius electas abietes illius et introibo altitudinem summitatis eius saltum Carmeli eius
ISA|37|25|ego fodi et bibi aquam et exsiccavi vestigio pedis mei omnes rivos aggerum
ISA|37|26|numquid non audisti quae olim fecerim ei ex diebus antiquis ego plasmavi illud et nunc adduxi et factum est in eradicationem collium conpugnantium et civitatum munitarum
ISA|37|27|habitatores earum breviata manu contremuerunt et confusi sunt facti sunt sicut faenum agri et gramen pascuae et herba tectorum quae exaruit antequam maturesceret
ISA|37|28|habitationem tuam et egressum tuum et introitum tuum cognovi et insaniam tuam contra me
ISA|37|29|cum fureres adversum me superbia tua ascendit in aures meas ponam ergo circulum in naribus tuis et frenum in labiis tuis et reducam te in viam per quam venisti
ISA|37|30|tibi autem hoc erit signum comede hoc anno quae sponte nascuntur et in anno secundo pomis vescere in anno autem tertio seminate et metite et plantate vineas et comedite fructum earum
ISA|37|31|et mittet id quod salvatum fuerit de domo Iuda et quod reliquum est radicem deorsum et faciet fructum sursum
ISA|37|32|quia de Hierusalem exibunt reliquiae et salvatio de monte Sion zelus Domini exercituum faciet istud
ISA|37|33|propterea haec dicit Dominus de rege Assyriorum non introibit civitatem hanc et non iaciet ibi sagittam et non occupabit eam clypeus et non mittet in circuitu eius aggerem
ISA|37|34|in via qua venit per eam revertetur et civitatem hanc non ingredietur dicit Dominus
ISA|37|35|et protegam civitatem istam ut salvem eam propter me et propter David servum meum
ISA|37|36|egressus est autem angelus Domini et percussit in castris Assyriorum centum octoginta quinque milia et surrexerunt mane et ecce omnes cadavera mortuorum
ISA|37|37|et egressus est et abiit et reversus est Sennacherib rex Assyriorum et habitavit in Nineve
ISA|37|38|et factum est cum adoraret in templo Nesrach deum suum Adramelech et Sarasar filii eius percusserunt eum gladio fugeruntque in terram Ararat et regnavit Asoraddon filius eius pro eo
ISA|38|1|in diebus illis aegrotavit Ezechias usque ad mortem et introivit ad eum Isaias filius Amos propheta et dixit ei haec dicit Dominus dispone domui tuae quia morieris tu et non vives
ISA|38|2|et convertit Ezechias faciem suam ad parietem et oravit ad Dominum
ISA|38|3|et dixit obsecro Domine memento quaeso quomodo ambulaverim coram te in veritate et in corde perfecto et quod bonum est in oculis tuis fecerim et flevit Ezechias fletu magno
ISA|38|4|et factum est verbum Domini ad Isaiam dicens
ISA|38|5|vade et dic Ezechiae haec dicit Dominus Deus David patris tui audivi orationem tuam vidi lacrimam tuam ecce ego adiciam super dies tuos quindecim annos
ISA|38|6|et de manu regis Assyriorum eruam te et civitatem istam et protegam eam
ISA|38|7|hoc autem tibi erit signum a Domino quia faciet Dominus verbum hoc quod locutus est
ISA|38|8|ecce ego reverti faciam umbram linearum per quas descenderat in horologio Ahaz in sole retrorsum decem lineis et reversus est sol decem lineis per gradus quos descenderat
ISA|38|9|scriptura Ezechiae regis Iuda cum aegrotasset et convaluisset de infirmitate sua
ISA|38|10|ego dixi in dimidio dierum meorum vadam ad portas inferi quaesivi residuum annorum meorum
ISA|38|11|dixi non videbo Dominum Dominum in terra viventium non aspiciam hominem ultra et habitatorem quievit
ISA|38|12|generatio mea ablata est et convoluta est a me quasi tabernaculum pastorum praecisa est velut a texente vita mea dum adhuc ordirer succidit me de mane usque ad vesperam finies me
ISA|38|13|sperabam usque ad mane quasi leo sic contrivit omnia ossa mea de mane usque ad vesperam finies me
ISA|38|14|sicut pullus hirundinis sic clamabo meditabor ut columba adtenuati sunt oculi mei suspicientes in excelsum Domine vim patior sponde pro me
ISA|38|15|quid dicam aut quid respondebit mihi cum ipse fecerit recogitabo omnes annos meos in amaritudine animae meae
ISA|38|16|Domine sic vivitur et in talibus vita spiritus mei corripies me et vivificabis me
ISA|38|17|ecce in pace amaritudo mea amarissima tu autem eruisti animam meam ut non periret proiecisti post tergum tuum omnia peccata mea
ISA|38|18|quia non infernus confitebitur tibi neque mors laudabit te non expectabunt qui descendunt in lacum veritatem tuam
ISA|38|19|vivens vivens ipse confitebitur tibi sicut et ego hodie pater filiis notam faciet veritatem tuam
ISA|38|20|Domine salvum me fac et psalmos nostros cantabimus cunctis diebus vitae nostrae in domo Domini
ISA|38|21|et iussit Isaias ut tollerent massam de ficis et cataplasmarent super vulnus et sanaretur
ISA|38|22|et dixit Ezechias quod erit signum quia ascendam in domo Domini
ISA|39|1|in tempore illo misit Marodach Baladan filius Baladan rex Babylonis libros et munera ad Ezechiam audierat enim quod aegrotasset et convaluisset
ISA|39|2|laetatus est autem super eis Ezechias et ostendit eis cellam aromatum et argenti et auri et odoramentorum et unguenti optimi et omnes apothecas supellectilis suae et universa quae inventa sunt in thesauris eius non fuit verbum quod non ostenderet eis Ezechias in domo sua et in omni potestate sua
ISA|39|3|introiit autem Isaias propheta ad regem Ezechiam et dixit ei quid dixerunt viri isti et unde venerunt ad te et dixit Ezechias de terra longinqua venerunt ad me de Babylone
ISA|39|4|et dixit quid viderunt in domo tua et dixit Ezechias omnia quae in domo mea sunt viderunt non fuit res quam non ostenderim eis in thesauris meis
ISA|39|5|et dixit Isaias ad Ezechiam audi verbum Domini exercituum
ISA|39|6|ecce dies venient et auferentur omnia quae in domo tua sunt et quae thesaurizaverunt patres tui usque ad diem hanc in Babylonem non relinquetur quicquam dicit Dominus
ISA|39|7|et de filiis tuis qui exibunt de te quos genueris tollent et erunt eunuchi in palatio regis Babylonis
ISA|39|8|et dixit Ezechias ad Isaiam bonum verbum Domini quod locutus est et dixit fiat tantum pax et veritas in diebus meis
ISA|40|1|consolamini consolamini populus meus dicit Deus vester
ISA|40|2|loquimini ad cor Hierusalem et avocate eam quoniam conpleta est malitia eius dimissa est iniquitas illius suscepit de manu Domini duplicia pro omnibus peccatis suis
ISA|40|3|vox clamantis in deserto parate viam Domini rectas facite in solitudine semitas Dei nostri
ISA|40|4|omnis vallis exaltabitur et omnis mons et collis humiliabitur et erunt prava in directa et aspera in vias planas
ISA|40|5|et revelabitur gloria Domini et videbit omnis caro pariter quod os Domini locutum est
ISA|40|6|vox dicentis clama et dixi quid clamabo omnis caro faenum et omnis gloria eius quasi flos agri
ISA|40|7|exsiccatum est faenum et cecidit flos quia spiritus Domini sufflavit in eo vere faenum est populus
ISA|40|8|exsiccatum est faenum cecidit flos verbum autem Dei nostri stabit in aeternum
ISA|40|9|super montem excelsum ascende tu quae evangelizas Sion exalta in fortitudine vocem tuam quae evangelizas Hierusalem exalta noli timere dic civitatibus Iudae ecce Deus vester
ISA|40|10|ecce Dominus Deus in fortitudine veniet et brachium eius dominabitur ecce merces eius cum eo et opus illius coram eo
ISA|40|11|sicut pastor gregem suum pascet in brachio suo congregabit agnos et in sinu suo levabit fetas ipse portabit
ISA|40|12|quis mensus est pugillo aquas et caelos palmo ponderavit quis adpendit tribus digitis molem terrae et libravit in pondere montes et colles in statera
ISA|40|13|quis adiuvit spiritum Domini aut quis consiliarius eius fuit et ostendit illi
ISA|40|14|cum quo iniit consilium et instruxit eum et docuit eum semitam iustitiae et erudivit eum scientiam et viam prudentiae ostendit illi
ISA|40|15|ecce gentes quasi stilla situlae et quasi momentum staterae reputatae sunt ecce insulae quasi pulvis exiguus
ISA|40|16|et Libanus non sufficiet ad succendendum et animalia eius non sufficient ad holocaustum
ISA|40|17|omnes gentes quasi non sint sic sunt coram eo et quasi nihilum et inane reputatae sunt ei
ISA|40|18|cui ergo similem fecistis Deum aut quam imaginem ponetis ei
ISA|40|19|numquid sculptile conflavit faber aut aurifex auro figuravit illud et lamminis argenteis argentarius
ISA|40|20|forte lignum et inputribile elegit artifex sapiens quaerit quomodo statuat simulacrum quod non moveatur
ISA|40|21|numquid non scietis numquid non audietis numquid non adnuntiatum est ab initio vobis numquid non intellexistis fundamenta terrae
ISA|40|22|qui sedet super gyrum terrae et habitatores eius sunt quasi lucustae qui extendit velut nihilum caelos et expandit eos sicut tabernaculum ad inhabitandum
ISA|40|23|qui dat secretorum scrutatores quasi non sint iudices terrae velut inane fecit
ISA|40|24|et quidem neque plantatos neque satos neque radicato in terra trunco eorum repente flavit in eos et aruerunt et turbo quasi stipulam auferet eos
ISA|40|25|et cui adsimilastis me et adaequastis dicit Sanctus
ISA|40|26|levate in excelsum oculos vestros et videte quis creavit haec qui educit in numero militiam eorum et omnes ex nomine vocat prae multitudine fortitudinis et roboris virtutisque eius neque unum reliquum fuit
ISA|40|27|quare dicis Iacob et loqueris Israhel abscondita est via mea a Domino et a Deo meo iudicium meum transibit
ISA|40|28|numquid nescis aut non audisti Deus sempiternus Dominus qui creavit terminos terrae non deficiet neque laborabit nec est investigatio sapientiae eius
ISA|40|29|qui dat lasso virtutem et his qui non sunt fortitudinem et robur multiplicat
ISA|40|30|deficient pueri et laborabunt et iuvenes in infirmitate cadent
ISA|40|31|qui autem sperant in Domino mutabunt fortitudinem adsument pinnas sicut aquilae current et non laborabunt ambulabunt et non deficient
ISA|41|1|taceant ad me insulae et gentes mutent fortitudinem accedant et tunc loquantur simul ad iudicium propinquemus
ISA|41|2|quis suscitavit ab oriente iustum vocavit eum ut sequeretur se dabit in conspectu eius gentes et reges obtinebit dabit quasi pulverem gladio eius sicut stipulam vento raptam arcui eius
ISA|41|3|persequetur eos transibit in pace semita in pedibus eius non apparebit
ISA|41|4|quis haec operatus est et fecit vocans generationes ab exordio ego Dominus primus et novissimus ego sum
ISA|41|5|viderunt insulae et timuerunt extrema terrae obstipuerunt adpropinquaverunt et accesserunt
ISA|41|6|unusquisque proximo suo auxiliatur et fratri suo dicit confortare
ISA|41|7|confortabit faber aerarius percutiens malleo eum qui cudebat tunc temporis dicens glutino bonum est et confortavit eum in clavis ut non moveatur
ISA|41|8|et tu Israhel serve meus Iacob quem elegi semen Abraham amici mei
ISA|41|9|in quo adprehendi te ab extremis terrae et a longinquis eius vocavi te et dixi tibi servus meus es tu elegi te et non abieci te
ISA|41|10|ne timeas quia tecum sum ego ne declines quia ego Deus tuus confortavi te et auxiliatus sum tui et suscepi te dextera iusti mei
ISA|41|11|ecce confundentur et erubescent omnes qui pugnant adversum te erunt quasi non sint et peribunt viri qui contradicunt tibi
ISA|41|12|quaeres eos et non invenies viros rebelles tuos erunt quasi non sint et veluti consumptio homines bellantes adversum te
ISA|41|13|quia ego Dominus Deus tuus adprehendens manum tuam dicensque tibi ne timeas ego adiuvi te
ISA|41|14|noli timere vermis Iacob qui mortui estis ex Israhel ego auxiliatus sum tui dicit Dominus et redemptor tuus Sanctus Israhel
ISA|41|15|ego posui te quasi plaustrum triturans novum habens rostra serrantia triturabis montes et comminues et colles quasi pulverem pones
ISA|41|16|ventilabis eos et ventus tollet et turbo disperget eos et tu exultabis in Domino in Sancto Israhel laetaberis
ISA|41|17|egeni et pauperes quaerunt aquas et non sunt lingua eorum siti aruit ego Dominus exaudiam eos Deus Israhel non derelinquam eos
ISA|41|18|aperiam in supinis collibus flumina et in medio camporum fontes ponam desertum in stagna aquarum et terram inviam in rivos aquarum
ISA|41|19|dabo in solitudine cedrum et spinam et myrtum et lignum olivae ponam in deserto abietem ulmum et buxum simul
ISA|41|20|ut videant et sciant et recogitent et intellegant pariter quia manus Domini fecit hoc et Sanctus Israhel creavit illud
ISA|41|21|prope facite iudicium vestrum dicit Dominus adferte si quid forte habetis dixit Rex Iacob
ISA|41|22|accedant et nuntient nobis quaecumque ventura sunt priora quae fuerint nuntiate et ponemus cor nostrum et sciemus novissima eorum et quae ventura sunt indicate nobis
ISA|41|23|adnuntiate quae ventura sunt in futurum et sciemus quia dii estis vos bene quoque aut male si potestis facite et loquamur et videamus simul
ISA|41|24|ecce vos estis ex nihilo et opus vestrum ex eo quod non est abominatio est qui elegit vos
ISA|41|25|suscitavi ab aquilone et venit ab ortu solis vocabit nomen meum et adducet magistratus quasi lutum et velut plastes conculcans humum
ISA|41|26|quis adnuntiavit ab exordio ut sciamus et a principio ut dicamus iustus es non est neque adnuntians neque praedicens neque audiens sermones vestros
ISA|41|27|primus ad Sion dicet ecce adsunt et Hierusalem evangelistam dabo
ISA|41|28|et vidi et non erat neque ex istis quisquam qui iniret consilium et interrogatus responderet verbum
ISA|41|29|ecce omnes iniusti et vana opera eorum ventus et inane simulacra eorum
ISA|42|1|ecce servus meus suscipiam eum electus meus conplacuit sibi in illo anima mea dedi spiritum meum super eum iudicium gentibus proferet
ISA|42|2|non clamabit neque accipiet personam nec audietur foris vox eius
ISA|42|3|calamum quassatum non conteret et linum fumigans non extinguet in veritate educet iudicium
ISA|42|4|non erit tristis neque turbulentus donec ponat in terra iudicium et legem eius insulae expectabunt
ISA|42|5|haec dicit Dominus Deus creans caelos et extendens eos firmans terram et quae germinant ex ea dans flatum populo qui est super eam et spiritum calcantibus eam
ISA|42|6|ego Dominus vocavi te in iustitia et adprehendi manum tuam et servavi et dedi te in foedus populi in lucem gentium
ISA|42|7|ut aperires oculos caecorum et educeres de conclusione vinctum de domo carceris sedentes in tenebris
ISA|42|8|ego Dominus hoc est nomen meum gloriam meam alteri non dabo et laudem meam sculptilibus
ISA|42|9|quae prima fuerant ecce venerunt nova quoque ego adnuntio antequam oriantur audita vobis faciam
ISA|42|10|cantate Domino canticum novum laus eius ab extremis terrae qui descenditis in mare et plenitudo eius insulae et habitatores earum
ISA|42|11|sublevetur desertum et civitates eius in domibus habitabit Cedar laudate habitatores Petrae de vertice montium clamabunt
ISA|42|12|ponent Domino gloriam et laudem eius in insulis nuntiabunt
ISA|42|13|Dominus sicut fortis egredietur sicut vir proeliator suscitabit zelum vociferabitur et clamabit super inimicos suos confortabitur
ISA|42|14|tacui semper silui patiens fui sicut pariens loquar dissipabo et absorbebo simul
ISA|42|15|desertos faciam montes et colles et omne gramen eorum exsiccabo et ponam flumina in insulas et stagna arefaciam
ISA|42|16|et ducam caecos in via quam nesciunt in semitis quas ignoraverunt ambulare eos faciam ponam tenebras coram eis in lucem et prava in recta haec verba feci eis et non dereliqui eos
ISA|42|17|conversi sunt retrorsum confundantur confusione qui confidunt in sculptili qui dicunt conflatili vos dii nostri
ISA|42|18|surdi audite et caeci intuemini ad videndum
ISA|42|19|quis caecus nisi servus meus et surdus nisi ad quem nuntios meos misi quis caecus nisi qui venundatus est quis caecus nisi servus Domini
ISA|42|20|qui vides multa nonne custodies qui apertas habes aures nonne audies
ISA|42|21|et Dominus voluit ut sanctificaret eum et magnificaret legem et extolleret
ISA|42|22|ipse autem populus direptus et vastatus laqueus iuvenum omnes et in domibus carcerum absconditi sunt facti sunt in rapinam nec est qui eruat in direptionem et non est qui dicat redde
ISA|42|23|quis est in vobis qui audiat hoc adtendat et auscultet futura
ISA|42|24|quis dedit in direptionem Iacob et Israhel vastantibus nonne Dominus ipse cui peccavimus et noluerunt in viis eius ambulare et non audierunt legem eius
ISA|42|25|et effudit super eum indignationem furoris sui et forte bellum et conbusit eum in circuitu et non cognovit et succendit eum et non intellexit
ISA|43|1|et nunc haec dicit Dominus creans te Iacob et formans te Israhel noli timere quia redemi te et vocavi nomine tuo meus es tu
ISA|43|2|cum transieris per aquas tecum ero et flumina non operient te cum ambulaveris in igne non conbureris et flamma non ardebit in te
ISA|43|3|quia ego Dominus Deus tuus Sanctus Israhel salvator tuus dedi propitiationem tuam Aegyptum Aethiopiam et Saba pro te
ISA|43|4|ex quo honorabilis factus es in oculis meis et gloriosus ego dilexi te et dabo homines pro te et populos pro anima tua
ISA|43|5|noli timere quoniam tecum ego sum ab oriente adducam semen tuum et ab occidente congregabo te
ISA|43|6|dicam aquiloni da et austro noli prohibere adfer filios meos de longinquo et filias meas ab extremis terrae
ISA|43|7|et omnem qui invocat nomen meum in gloriam meam creavi eum et formavi eum et feci eum
ISA|43|8|educ foras populum caecum et oculos habentem surdum et aures ei sunt
ISA|43|9|omnes gentes congregatae sunt simul et collectae sunt tribus quis in vobis adnuntiet istud et quae prima sunt audire nos faciat dent testes eorum et iustificentur et audiant et dicant vere
ISA|43|10|vos testes mei dicit Dominus et servus meus quem elegi ut sciatis et credatis mihi et intellegatis quia ego ipse sum ante me non est formatus deus et post me non erit
ISA|43|11|ego sum ego sum Dominus et non est absque me salvator
ISA|43|12|ego adnuntiavi et salvavi auditum feci et non fuit in vobis alienus vos testes mei dicit Dominus et ego Deus
ISA|43|13|et ab initio ego ipse et non est qui de manu mea eruat operabor et quis avertet illud
ISA|43|14|haec dicit Dominus redemptor vester Sanctus Israhel propter vos emisi Babylonem et detraxi vectes universos et Chaldeos in navibus suis gloriantes
ISA|43|15|ego Dominus Sanctus vester creans Israhel Rex vester
ISA|43|16|haec dicit Dominus qui dedit in mari viam et in aquis torrentibus semitam
ISA|43|17|qui eduxit quadrigam et equum agmen et robustum simul obdormierunt nec resurgent contriti sunt quasi linum et extincti sunt
ISA|43|18|ne memineritis priorum et antiqua ne intueamini
ISA|43|19|ecce ego facio nova et nunc orientur utique cognoscetis ea ponam in deserto viam et in invio flumina
ISA|43|20|glorificabit me bestia agri dracones et strutiones quia dedi in deserto aquas flumina in invio ut darem potum populo meo electo meo
ISA|43|21|populum istum formavi mihi laudem meam narrabit
ISA|43|22|non me invocasti Iacob nec laborasti in me Israhel
ISA|43|23|non obtulisti mihi arietem holocausti tui et victimis tuis non glorificasti me non te servire feci in oblatione nec laborem tibi praebui in ture
ISA|43|24|non emisti mihi argento calamum et adipe victimarum tuarum non inebriasti me verumtamen servire me fecisti in peccatis tuis praebuisti mihi laborem in iniquitatibus tuis
ISA|43|25|ego sum ego sum ipse qui deleo iniquitates tuas propter me et peccatorum tuorum non recordabor
ISA|43|26|reduc me in memoriam et iudicemur simul narra si quid habes ut iustificeris
ISA|43|27|pater tuus primus peccavit et interpretes tui praevaricati sunt in me
ISA|43|28|et contaminavi principes sanctos dedi ad internicionem Iacob et Israhel in blasphemiam
ISA|44|1|et nunc audi Iacob serve meus et Israhel quem elegi
ISA|44|2|haec dicit Dominus faciens et formans te ab utero auxiliator tuus noli timere serve meus Iacob et Rectissime quem elegi
ISA|44|3|effundam enim aquas super sitientem et fluenta super aridam effundam spiritum meum super semen tuum et benedictionem meam super stirpem tuam
ISA|44|4|et germinabunt inter herbas quasi salices iuxta praeterfluentes aquas
ISA|44|5|iste dicet Domini ego sum et ille vocabit in nomine Iacob et hic scribet manu sua Domino et in nomine Israhel adsimilabitur
ISA|44|6|haec dicit Dominus rex Israhel et redemptor eius Dominus exercituum ego primus et ego novissimus et absque me non est deus
ISA|44|7|quis similis mei vocet et adnuntiet et ordinem exponat mihi ex quo constitui populum antiquum ventura et quae futura sunt adnuntient eis
ISA|44|8|nolite timere neque conturbemini ex tunc audire te feci et adnuntiavi vos estis testes mei numquid est deus absque me et formator quem ego non noverim
ISA|44|9|plastae idoli omnes nihil sunt et amantissima eorum non proderunt eis ipsi sunt testes eorum quia non vident neque intellegunt ut confundantur
ISA|44|10|quis formavit deum et sculptile conflavit ad nihil utile
ISA|44|11|ecce omnes participes eius confundentur fabri enim sunt ex hominibus convenient omnes stabunt et pavebunt et confundentur simul
ISA|44|12|faber ferrarius lima operatus est in prunis et in malleis formavit illud et operatus est in brachio fortitudinis suae esuriet et deficiet non bibet aquam et lassescet
ISA|44|13|artifex lignarius extendit normam formavit illud in runcina fecit illud in angularibus et in circino tornavit illud et fecit imaginem viri quasi speciosum hominem habitantem in domo
ISA|44|14|succidit cedros tulit ilicem et quercum quae steterat inter ligna saltus plantavit pinum quam pluvia nutrivit
ISA|44|15|et facta est hominibus in focum sumpsit ex eis et calefactus est et succendit et coxit panes de reliquo autem operatus est deum et adoravit fecit sculptile et curvatus est ante illud
ISA|44|16|medium eius conbusit igni et de medio eius carnes comedit coxit pulmentum et saturatus est et calefactus est et dixit va calefactus sum vidi focum
ISA|44|17|reliquum autem eius deum fecit sculptile sibi curvatur ante illud et adorat illud et obsecrat dicens libera me quia deus meus es tu
ISA|44|18|nescierunt neque intellexerunt lutati enim sunt ne videant oculi eorum et ne intellegant corde suo
ISA|44|19|non recogitant in mente sua neque cognoscunt neque sentiunt ut dicant medietatem eius conbusi igne et coxi super carbones eius panes coxi carnes et comedi et de reliquo eius idolum faciam ante truncum ligni procidam
ISA|44|20|pars eius cinis est cor insipiens adoravit illud et non liberabit animam suam neque dicet forte mendacium est in dextera mea
ISA|44|21|memento horum Iacob et Israhel quoniam servus meus es tu formavi te servus meus es tu Israhel non oblivisceris mei
ISA|44|22|delevi ut nubem iniquitates tuas et quasi nebulam peccata tua revertere ad me quoniam redemi te
ISA|44|23|laudate caeli quoniam fecit Dominus iubilate extrema terrae resonate montes laudationem saltus et omne lignum eius quoniam redemit Dominus Iacob et Israhel gloriabitur
ISA|44|24|haec dicit Dominus redemptor tuus et formator tuus ex utero ego sum Dominus faciens omnia extendens caelos solus stabiliens terram et nullus mecum
ISA|44|25|irrita faciens signa divinorum et ariolos in furorem vertens convertens sapientes retrorsum et scientiam eorum stultam faciens
ISA|44|26|suscitans verbum servi sui et consilium nuntiorum suorum conplens qui dico Hierusalem habitaberis et civitatibus Iuda aedificabimini et deserta eius suscitabo
ISA|44|27|qui dico profundo desolare et flumina tua arefaciam
ISA|44|28|qui dico Cyro pastor meus es et omnem voluntatem meam conplebis qui dico Hierusalem aedificaberis et templo fundaberis
ISA|45|1|haec dicit Dominus christo meo Cyro cuius adprehendi dexteram ut subiciam ante faciem eius gentes et dorsa regum vertam et aperiam coram eo ianuas et portae non cludentur
ISA|45|2|ego ante te ibo et gloriosos terrae humiliabo portas aereas conteram et vectes ferreos confringam
ISA|45|3|et dabo tibi thesauros absconditos et arcana secretorum ut scias quia ego Dominus qui voco nomen tuum Deus Israhel
ISA|45|4|propter servum meum Iacob et Israhel electum meum et vocavi te in nomine tuo adsimilavi te et non cognovisti me
ISA|45|5|ego Dominus et non est amplius extra me non est deus accinxi te et non cognovisti me
ISA|45|6|ut sciant hii qui ab ortu solis et qui ab occidente quoniam absque me non est ego Dominus et non est alter
ISA|45|7|formans lucem et creans tenebras faciens pacem et creans malum ego Dominus faciens omnia haec
ISA|45|8|rorate caeli desuper et nubes pluant iustum aperiatur terra et germinet salvatorem et iustitia oriatur simul ego Dominus creavi eum
ISA|45|9|vae qui contradicit fictori suo testa de samiis terrae numquid dicet lutum figulo suo quid facis et opus tuum absque manibus est
ISA|45|10|vae qui dicit patri quid generas et mulieri quid parturis
ISA|45|11|haec dicit Dominus Sanctus Israhel plastes eius ventura interrogate me super filios meos et super opus manuum mearum mandastis mihi
ISA|45|12|ego feci terram et hominem super eam creavi ego manus meae tetenderunt caelos et omni militiae eorum mandavi
ISA|45|13|ego suscitavi eum ad iustitiam et omnes vias eius dirigam ipse aedificabit civitatem meam et captivitatem meam dimittet non in pretio neque in muneribus dicit Dominus Deus exercituum
ISA|45|14|haec dicit Dominus labor Aegypti et negotiatio Aethiopiae et Sabaim viri sublimes ad te transibunt et tui erunt post te ambulabunt vincti manicis pergent et te adorabunt teque deprecabuntur tantum in te est Deus et non est absque te deus
ISA|45|15|vere tu es Deus absconditus Deus Israhel salvator
ISA|45|16|confusi sunt et erubuerunt omnes simul abierunt in confusione fabricatores errorum
ISA|45|17|Israhel salvatus est in Domino salute aeterna non confundemini et non erubescetis usque in saeculum saeculi
ISA|45|18|quia haec dicit Dominus creans caelos ipse Deus formans terram et faciens eam ipse plastes eius non in vanum creavit eam ut habitetur formavit eam ego Dominus et non est alius
ISA|45|19|non in abscondito locutus sum in loco terrae tenebroso non dixi semini Iacob frustra quaerite me ego Dominus loquens iustitiam adnuntians recta
ISA|45|20|congregamini et venite et accedite simul qui salvati estis ex gentibus nescierunt qui levant lignum sculpturae suae et rogant deum non salvantem
ISA|45|21|adnuntiate et venite et consiliamini simul quis auditum fecit hoc ab initio ex tunc praedixit illud numquid non ego Dominus et non est ultra Deus absque me Deus iustus et salvans non est praeter me
ISA|45|22|convertimini ad me et salvi eritis omnes fines terrae quia ego Deus et non est alius
ISA|45|23|in memet ipso iuravi egredietur de ore meo iustitiae verbum et non revertetur quia mihi curvabunt omnia genu et iurabit omnis lingua
ISA|45|24|ergo in Domino dicet meae sunt iustitiae et imperium ad eum venient et confundentur omnes qui repugnant ei
ISA|45|25|in Domino iustificabitur et laudabitur omne semen Israhel
ISA|46|1|conflatus est Bel contritus est Nabo facta sunt simulacra eorum bestiis et iumentis onera vestra gravi pondere usque ad lassitudinem
ISA|46|2|contabuerunt et contrita sunt simul non potuerunt salvare portantem et anima eorum in captivitatem ibit
ISA|46|3|audite me domus Iacob et omne residuum domus Israhel qui portamini a meo utero qui gestamini a mea vulva
ISA|46|4|usque ad senectam ego ipse et usque ad canos ego portabo ego feci et ego feram et ego portabo et salvabo
ISA|46|5|cui adsimilastis me et adaequastis et conparastis me et fecistis similem
ISA|46|6|qui confertis aurum de sacculo et argentum statera ponderatis conducentes aurificem ut faciat deum et procidunt et adorant
ISA|46|7|portant illud in umeris gestantes et ponentes in loco suo et stabit ac de loco suo non movebitur sed et cum clamaverint ad eum non audiet de tribulatione non salvabit eos
ISA|46|8|mementote istud et fundamini redite praevaricatores ad cor
ISA|46|9|recordamini prioris saeculi quoniam ego sum Deus et non est ultra Deus nec est similis mei
ISA|46|10|adnuntians ab exordio novissimum et ab initio quae necdum facta sunt dicens consilium meum stabit et omnis voluntas mea fiet
ISA|46|11|vocans ab oriente avem et de terra longinqua virum voluntatis meae et locutus sum et adducam illud creavi et faciam illud
ISA|46|12|audite me duro corde qui longe estis a iustitia
ISA|46|13|prope feci iustitiam meam non elongabitur et salus mea non morabitur dabo in Sion salutem et Israheli gloriam meam
ISA|47|1|descende sede in pulverem virgo filia Babylon sede in terra non est solium filiae Chaldeorum quia ultra non vocaberis mollis et tenera
ISA|47|2|tolle molam et mole farinam denuda turpitudinem tuam discoperi umerum revela crus transi flumina
ISA|47|3|revelabitur ignominia tua et videbitur obprobrium tuum ultionem capiam et non resistet mihi homo
ISA|47|4|redemptor noster Dominus exercituum nomen illius Sanctus Israhel
ISA|47|5|sede tace et intra in tenebras filia Chaldeorum quia non vocaberis ultra domina regnorum
ISA|47|6|iratus sum super populum meum contaminavi hereditatem meam et dedi eos in manu tua non posuisti eis misericordias super senem adgravasti iugum tuum valde
ISA|47|7|et dixisti in sempiternum ero domina non posuisti haec super cor tuum neque recordata es novissimi tui
ISA|47|8|et nunc audi haec delicata et habitans confidenter quae dicis in corde tuo ego sum et non est praeter me amplius non sedebo vidua et ignorabo sterilitatem
ISA|47|9|venient tibi duo haec subito in die una sterilitas et viduitas universa venerunt super te propter multitudinem maleficiorum tuorum et propter duritiam incantatorum tuorum vehementem
ISA|47|10|et fiduciam habuisti in malitia tua et dixisti non est qui videat me sapientia tua et scientia tua haec decepit te et dixisti in corde tuo ego sum et praeter me non est altera
ISA|47|11|veniet super te malum et nescies ortum eius et inruet super te calamitas quam non poteris expiare veniet super te repente miseria quam nescies
ISA|47|12|sta cum incantatoribus tuis et cum multitudine maleficiorum tuorum in quibus laborasti ab adulescentia tua si forte quid prosit tibi aut si possis fieri fortior
ISA|47|13|defecisti in multitudine consiliorum tuorum stent et salvent te augures caeli qui contemplabantur sidera et supputabant menses ut ex eis adnuntiarent ventura tibi
ISA|47|14|ecce facti sunt quasi stipula ignis conbusit eos non liberabunt animam suam de manu flammae non sunt prunae quibus calefiant nec focus ut sedeant ad eum
ISA|47|15|sic facta sunt tibi in quibuscumque laboraveras negotiatores tui ab adulescentia tua unusquisque in via sua erraverunt non est qui salvet te
ISA|48|1|audite hoc domus Iacob qui vocamini nomine Israhel et de aquis Iuda existis qui iuratis in nomine Domini et Dei Israhel recordamini non in veritate neque in iustitia
ISA|48|2|de civitate enim sancta vocati sunt et super Deum Israhel constabiliti sunt Dominus exercituum nomen eius
ISA|48|3|priora ex tunc adnuntiavi et ex ore meo exierunt et audita feci ea repente operatus sum et venerunt
ISA|48|4|scivi enim quia durus es tu et nervus ferreus cervix tua et frons tua aerea
ISA|48|5|praedixi tibi ex tunc antequam venirent indicavi tibi ne forte diceres idola mea fecerunt haec et sculptilia mea et conflatilia mandaverunt ista
ISA|48|6|quae audisti vide omnia vos autem non adnuntiastis audita feci tibi nova ex nunc et conservata quae nescis
ISA|48|7|nunc creata sunt et non ex tunc et ante diem et non audisti ea ne forte dicas ecce cognovi ea
ISA|48|8|neque audisti neque cognovisti neque ex tunc aperta est auris tua scio enim quia praevaricans praevaricabis et transgressorem ex ventre vocavi te
ISA|48|9|propter nomen meum longe faciam furorem meum et laude mea infrenabo te ne intereas
ISA|48|10|ecce excoxi te sed non quasi argentum elegi te in camino paupertatis
ISA|48|11|propter me propter me faciam ut non blasphemer et gloriam meam alteri non dabo
ISA|48|12|audi me Iacob et Israhel quem ego voco ego ipse ego primus et ego novissimus
ISA|48|13|manus quoque mea fundavit terram et dextera mea mensa est caelos ego vocabo eos et stabunt simul
ISA|48|14|congregamini omnes vos et audite quis de eis adnuntiavit haec Dominus dilexit eum faciet voluntatem suam in Babylone et brachium suum in Chaldeis
ISA|48|15|ego ego locutus sum et vocavi eum adduxi eum et directa est via eius
ISA|48|16|accedite ad me et audite hoc non a principio in abscondito locutus sum ex tempore antequam fieret ibi eram et nunc Dominus Deus misit me et spiritus eius
ISA|48|17|haec dicit Dominus redemptor tuus Sanctus Israhel ego Dominus Deus tuus docens te utilia gubernans te in via qua ambulas
ISA|48|18|utinam adtendisses mandata mea facta fuisset sicut flumen pax tua et iustitia tua sicut gurgites maris
ISA|48|19|et fuisset quasi harena semen tuum et stirps uteri tui ut lapilli eius non interisset et non fuisset adtritum nomen eius a facie mea
ISA|48|20|egredimini de Babylone fugite a Chaldeis in voce exultationis adnuntiate auditum facite hoc efferte illud usque ad extrema terrae dicite redemit Dominus servum suum Iacob
ISA|48|21|non sitierunt in deserto cum educeret eos aquam de petra produxit eis et scidit petram et fluxerunt aquae
ISA|48|22|non est pax dicit Dominus impiis
ISA|49|1|audite insulae et adtendite populi de longe Dominus ab utero vocavit me de ventre matris meae recordatus est nominis mei
ISA|49|2|et posuit os meum quasi gladium acutum in umbra manus suae protexit me et posuit me sicut sagittam electam in faretra sua abscondit me
ISA|49|3|et dixit mihi servus meus es tu Israhel quia in te gloriabor
ISA|49|4|et ego dixi in vacuum laboravi sine causa et vane fortitudinem meam consumpsi ergo iudicium meum cum Domino et opus meum cum Deo meo
ISA|49|5|et nunc dicit Dominus formans me ex utero servum sibi ut reducam Iacob ad eum et Israhel non congregabitur et glorificatus sum in oculis Domini et Deus meus factus est fortitudo mea
ISA|49|6|et dixit parum est ut sis mihi servus ad suscitandas tribus Iacob et feces Israhel convertendas dedi te in lucem gentium ut sis salus mea usque ad extremum terrae
ISA|49|7|haec dicit Dominus redemptor Israhel Sanctus eius ad contemptibilem animam ad abominatam gentem ad servum dominorum reges videbunt et consurgent principes et adorabunt propter Dominum quia fidelis est et Sanctum Israhel qui elegit te
ISA|49|8|haec dicit Dominus in tempore placito exaudivi te et in die salutis auxiliatus sum tui et servavi te et dedi te in foedus populi ut suscitares terram et possideres hereditates dissipatas
ISA|49|9|ut diceres his qui vincti sunt exite et his qui in tenebris revelamini super vias pascentur et in omnibus planis pascua eorum
ISA|49|10|non esurient neque sitient et non percutiet eos aestus et sol quia miserator eorum reget eos et ad fontes aquarum portabit eos
ISA|49|11|et ponam omnes montes meos in viam et semitae meae exaltabuntur
ISA|49|12|ecce isti de longe venient et ecce illi ab aquilone et mari et isti de terra australi
ISA|49|13|laudate caeli et exulta terra iubilate montes laudem quia consolatus est Dominus populum suum et pauperum suorum miserebitur
ISA|49|14|et dixit Sion dereliquit me Dominus et Dominus oblitus est mei
ISA|49|15|numquid oblivisci potest mulier infantem suum ut non misereatur filio uteri sui et si illa oblita fuerit ego tamen non obliviscar tui
ISA|49|16|ecce in manibus meis descripsi te muri tui coram oculis meis semper
ISA|49|17|venerunt structores tui destruentes te et dissipantes a te exibunt
ISA|49|18|leva in circuitu oculos tuos et vide omnes isti congregati sunt venerunt tibi vivo ego dicit Dominus quia omnibus his velut ornamento vestieris et circumdabis tibi eos quasi sponsa
ISA|49|19|quia deserta tua et solitudines tuae et terra ruinae tuae nunc angusta erunt prae habitatoribus et longe fugabuntur qui absorbebant te
ISA|49|20|adhuc dicent in auribus tuis filii sterilitatis tuae angustus mihi est locus fac spatium mihi ut habitem
ISA|49|21|et dices in corde tuo quis genuit mihi istos ego sterilis et non pariens transmigrata et captiva et istos quis enutrivit ego destituta et sola et isti ubi hic erant
ISA|49|22|haec dicit Dominus Deus ecce levo ad gentes manum meam et ad populos exaltabo signum meum et adferent filios tuos in ulnis et filias tuas super umeros portabunt
ISA|49|23|et erunt reges nutricii tui et reginae nutrices tuae vultu in terra dimisso adorabunt te et pulverem pedum tuorum lingent et scies quia ego Dominus super quo non confundentur qui expectant eum
ISA|49|24|numquid tolletur a forte praeda aut quod captum fuerit a robusto salvum esse poterit
ISA|49|25|quia haec dicit Dominus equidem et captivitas a forte tolletur et quod ablatum fuerit a robusto salvabitur eos vero qui iudicaverunt te ego iudicabo et filios tuos ego salvabo
ISA|49|26|et cibabo hostes tuos carnibus suis et quasi musto sanguine suo inebriabuntur et sciet omnis caro quia ego Dominus salvans te et redemptor tuus Fortis Iacob
ISA|50|1|haec dicit Dominus quis est hic liber repudii matris vestrae quo dimisi eam aut quis est creditor meus cui vendidi vos ecce in iniquitatibus vestris venditi estis et in sceleribus vestris dimisi matrem vestram
ISA|50|2|quia veni et non erat vir vocavi et non erat qui audiret numquid adbreviata et parvula facta est manus mea ut non possim redimere aut non est in me virtus ad liberandum ecce in increpatione mea desertum faciam mare ponam flumina in siccum conputrescent pisces sine aqua et morientur in siti
ISA|50|3|induam caelos tenebris et saccum ponam operimentum eorum
ISA|50|4|Dominus dedit mihi linguam eruditam ut sciam sustentare eum qui lassus est verbo erigit mane mane erigit mihi aurem ut audiam quasi magistrum
ISA|50|5|Dominus Deus aperuit mihi aurem ego autem non contradico retrorsum non abii
ISA|50|6|corpus meum dedi percutientibus et genas meas vellentibus faciem meam non averti ab increpantibus et conspuentibus
ISA|50|7|Dominus Deus auxiliator meus ideo non sum confusus ideo posui faciem meam ut petram durissimam et scio quoniam non confundar
ISA|50|8|iuxta est qui iustificat me quis contradicet mihi stemus simul quis est adversarius meus accedat ad me
ISA|50|9|ecce Dominus Deus auxiliator meus quis est qui condemnet me ecce omnes quasi vestimentum conterentur tinea comedet eos
ISA|50|10|quis ex vobis timens Dominum audiens vocem servi sui qui ambulavit in tenebris et non est lumen ei speret in nomine Domini et innitatur super Deum suum
ISA|50|11|ecce omnes vos accendentes ignem accincti flammis ambulate in lumine ignis vestri et in flammis quas succendistis de manu mea factum est hoc vobis in doloribus dormietis
ISA|51|1|audite me qui sequimini quod iustum est et quaeritis Dominum adtendite ad petram unde excisi estis et ad cavernam laci de qua praecisi estis
ISA|51|2|adtendite ad Abraham patrem vestrum et ad Sarram quae peperit vos quia unum vocavi eum et benedixi ei et multiplicavi eum
ISA|51|3|consolabitur ergo Dominus et Sion consolabitur omnes ruinas eius et ponet desertum eius quasi delicias et solitudinem eius quasi hortum Domini gaudium et laetitia invenietur in ea gratiarum actio et vox laudis
ISA|51|4|adtendite ad me populus meus et tribus mea me audite quia lex a me exiet et iudicium meum in lucem populorum requiescet
ISA|51|5|prope est iustus meus egressus est salvator meus et brachia mea populos iudicabunt me insulae expectabunt et brachium meum sustinebunt
ISA|51|6|levate in caelum oculos vestros et videte sub terra deorsum quia caeli sicut fumus liquescent et terra sicut vestimentum adteretur et habitatores eius sicut haec interibunt salus autem mea in sempiternum erit et iustitia mea non deficiet
ISA|51|7|audite me qui scitis iustum populus lex mea in corde eorum nolite timere obprobrium hominum et blasphemias eorum ne metuatis
ISA|51|8|sicut enim vestimentum sic comedet eos vermis et sicut lanam sic devorabit eos tinea salus autem mea in sempiternum erit et iustitia mea in generationes generationum
ISA|51|9|consurge consurge induere fortitudinem brachium Domini consurge sicut in diebus antiquis in generationibus saeculorum numquid non tu percussisti superbum vulnerasti draconem
ISA|51|10|numquid non tu siccasti mare aquam abyssi vehementis qui posuisti profundum maris viam ut transirent liberati
ISA|51|11|et nunc qui redempti sunt a Domino revertentur et venient in Sion laudantes et laetitia sempiterna super capita eorum gaudium et laetitiam tenebunt fugiet dolor et gemitus
ISA|51|12|ego ego ipse consolabor vos quis tu ut timeres ab homine mortali et a filio hominis qui quasi faenum ita arescet
ISA|51|13|et oblitus es Domini factoris tui qui tetendit caelos et fundavit terram et formidasti iugiter tota die a facie furoris eius qui te tribulabat et paraverat ad perdendum ubi nunc est furor tribulantis
ISA|51|14|cito veniet gradiens ad aperiendum et non interficiet usque ad internicionem nec deficiet panis eius
ISA|51|15|ego autem sum Dominus Deus tuus qui conturbo mare et intumescunt fluctus eius Dominus exercituum nomen meum
ISA|51|16|posui verba mea in ore tuo et in umbra manus meae protexi te ut plantes caelos et fundes terram et dicas ad Sion populus meus es tu
ISA|51|17|elevare elevare consurge Hierusalem quae bibisti de manu Domini calicem irae eius usque ad fundum calicis soporis bibisti et epotasti usque ad feces
ISA|51|18|non est qui sustentet eam ex omnibus filiis quos genuit et non est qui adprehendat manum eius ex omnibus filiis quos enutrivit
ISA|51|19|duo sunt quae occurrerunt tibi quis contristabitur super te vastitas et contritio et fames et gladius quis consolabitur te
ISA|51|20|filii tui proiecti sunt dormierunt in capite omnium viarum sicut bestia inlaqueata pleni indignatione Domini increpatione Dei tui
ISA|51|21|idcirco audi hoc paupercula et ebria non a vino
ISA|51|22|haec dicit Dominator tuus Dominus et Deus tuus qui pugnavit pro populo suo ecce tuli de manu tua calicem soporis fundum calicis indignationis meae non adicies ut bibas illud ultra
ISA|51|23|et ponam illud in manu eorum qui te humiliaverunt et dixerunt animae tuae incurvare ut transeamus et posuisti ut terram corpus tuum et quasi viam transeuntibus
ISA|52|1|consurge consurge induere fortitudine tua Sion induere vestimentis gloriae tuae Hierusalem civitas sancti quia non adiciet ultra ut pertranseat per te incircumcisus et inmundus
ISA|52|2|excutere de pulvere consurge sede Hierusalem solve vincula colli tui captiva filia Sion
ISA|52|3|quia haec dicit Dominus gratis venundati estis et sine argento redimemini
ISA|52|4|quia haec dicit Dominus Deus in Aegyptum descendit populus meus in principio ut colonus esset ibi et Assur absque ulla causa calumniatus est eum
ISA|52|5|et nunc quid mihi est hic dicit Dominus quoniam ablatus est populus meus gratis dominatores eius inique agunt dicit Dominus et iugiter tota die nomen meum blasphematur
ISA|52|6|propter hoc sciet populus meus nomen meum in die illa quia ego ipse qui loquebar ecce adsum
ISA|52|7|quam pulchri super montes pedes adnuntiantis et praedicantis pacem adnuntiantis bonum praedicantis salutem dicentis Sion regnavit Deus tuus
ISA|52|8|vox speculatorum tuorum levaverunt vocem simul laudabunt quia oculum ad oculum videbunt cum converterit Dominus Sion
ISA|52|9|gaudete et laudate simul deserta Hierusalem quia consolatus est Dominus populum suum redemit Hierusalem
ISA|52|10|paravit Dominus brachium sanctum suum in oculis omnium gentium et videbunt omnes fines terrae salutare Dei nostri
ISA|52|11|recedite recedite exite inde pollutum nolite tangere exite de medio eius mundamini qui fertis vasa Domini
ISA|52|12|quoniam non in tumultu exibitis nec in fuga properabitis praecedet enim vos Dominus et congregabit vos Deus Israhel
ISA|52|13|ecce intelleget servus meus exaltabitur et elevabitur et sublimis erit valde
ISA|52|14|sicut obstipuerunt super te multi sic inglorius erit inter viros aspectus eius et forma eius inter filios hominum
ISA|52|15|iste asperget gentes multas super ipsum continebunt reges os suum quia quibus non est narratum de eo viderunt et qui non audierunt contemplati sunt
ISA|53|1|quis credidit auditui nostro et brachium Domini cui revelatum est
ISA|53|2|et ascendet sicut virgultum coram eo et sicut radix de terra sitienti non est species ei neque decor et vidimus eum et non erat aspectus et desideravimus eum
ISA|53|3|despectum et novissimum virorum virum dolorum et scientem infirmitatem et quasi absconditus vultus eius et despectus unde nec reputavimus eum
ISA|53|4|vere languores nostros ipse tulit et dolores nostros ipse portavit et nos putavimus eum quasi leprosum et percussum a Deo et humiliatum
ISA|53|5|ipse autem vulneratus est propter iniquitates nostras adtritus est propter scelera nostra disciplina pacis nostrae super eum et livore eius sanati sumus
ISA|53|6|omnes nos quasi oves erravimus unusquisque in viam suam declinavit et Dominus posuit in eo iniquitatem omnium nostrum
ISA|53|7|oblatus est quia ipse voluit et non aperuit os suum sicut ovis ad occisionem ducetur et quasi agnus coram tondente obmutescet et non aperiet os suum
ISA|53|8|de angustia et de iudicio sublatus est generationem eius quis enarrabit quia abscisus est de terra viventium propter scelus populi mei percussit eum
ISA|53|9|et dabit impios pro sepultura et divitem pro morte sua eo quod iniquitatem non fecerit neque dolus fuerit in ore eius
ISA|53|10|et Dominus voluit conterere eum in infirmitate si posuerit pro peccato animam suam videbit semen longevum et voluntas Domini in manu eius dirigetur
ISA|53|11|pro eo quod laboravit anima eius videbit et saturabitur in scientia sua iustificabit ipse iustus servus meus multos et iniquitates eorum ipse portabit
ISA|53|12|ideo dispertiam ei plurimos et fortium dividet spolia pro eo quod tradidit in morte animam suam et cum sceleratis reputatus est et ipse peccatum multorum tulit et pro transgressoribus rogavit
ISA|54|1|lauda sterilis quae non paris decanta laudem et hinni quae non pariebas quoniam multi filii desertae magis quam eius quae habebat virum dicit Dominus
ISA|54|2|dilata locum tentorii tui et pelles tabernaculorum tuorum extende ne parcas longos fac funiculos tuos et clavos tuos consolida
ISA|54|3|ad dexteram enim et ad levam penetrabis et semen tuum gentes hereditabit et civitates desertas inhabitabit
ISA|54|4|noli timere quia non confunderis neque erubescas non enim te pudebit quia confusionis adulescentiae tuae oblivisceris et obprobrii viduitatis tuae non recordaberis amplius
ISA|54|5|quia dominabitur tui qui fecit te Dominus exercituum nomen eius et redemptor tuus Sanctus Israhel Deus omnis terrae vocabitur
ISA|54|6|quia ut mulierem derelictam et maerentem spiritu vocavit te Dominus et uxorem ab adulescentia abiectam dixit Deus tuus
ISA|54|7|ad punctum in modico dereliqui te et in miserationibus magnis congregabo te
ISA|54|8|in momento indignationis abscondi faciem meam parumper a te et in misericordia sempiterna misertus sum tui dixit redemptor tuus Dominus
ISA|54|9|sicut in diebus Noe istud mihi est cui iuravi ne inducerem aquas Noe ultra super terram sic iuravi ut non irascar tibi et non increpem te
ISA|54|10|montes enim commovebuntur et colles contremescent misericordia autem mea non recedet et foedus pacis meae non movebitur dixit miserator tuus Dominus
ISA|54|11|paupercula tempestate convulsa absque ulla consolatione ecce ego sternam per ordinem lapides tuos et fundabo te in sapphyris
ISA|54|12|et ponam iaspidem propugnacula tua et portas tuas in lapides sculptos et omnes terminos tuos in lapides desiderabiles
ISA|54|13|universos filios tuos doctos a Domino et multitudinem pacis filiis tuis
ISA|54|14|et in iustitia fundaberis recede procul a calumnia quia non timebis et a pavore quia non adpropinquabit tibi
ISA|54|15|ecce accola veniet qui non erat mecum advena quondam tuus adiungetur tibi
ISA|54|16|ecce ego creavi fabrum sufflantem in igne prunas et proferentem vas in opus suum et ego creavi interfectorem ad disperdendum
ISA|54|17|omne vas quod fictum est contra te non dirigetur et omnem linguam resistentem tibi in iudicio iudicabis haec hereditas servorum Domini et iustitia eorum apud me dicit Dominus
ISA|55|1|o omnes sitientes venite ad aquas et qui non habetis argentum properate emite et comedite venite emite absque argento et absque ulla commutatione vinum et lac
ISA|55|2|quare adpenditis argentum non in panibus et laborem vestrum non in saturitate audite audientes me et comedite bonum et delectabitur in crassitudine anima vestra
ISA|55|3|inclinate aurem vestram et venite ad me audite et vivet anima vestra et feriam vobis pactum sempiternum misericordias David fideles
ISA|55|4|ecce testem populis dedi eum ducem ac praeceptorem gentibus
ISA|55|5|ecce gentem quam nesciebas vocabis et gentes quae non cognoverunt te ad te current propter Dominum Deum tuum et Sanctum Israhel quia glorificavit te
ISA|55|6|quaerite Dominum dum inveniri potest invocate eum dum prope est
ISA|55|7|derelinquat impius viam suam et vir iniquus cogitationes suas et revertatur ad Dominum et miserebitur eius et ad Deum nostrum quoniam multus est ad ignoscendum
ISA|55|8|non enim cogitationes meae cogitationes vestrae neque viae vestrae viae meae dicit Dominus
ISA|55|9|quia sicut exaltantur caeli a terra sic exaltatae sunt viae meae a viis vestris et cogitationes meae a cogitationibus vestris
ISA|55|10|et quomodo descendit imber et nix de caelo et illuc ultra non revertitur sed inebriat terram et infundit eam et germinare eam facit et dat semen serenti et panem comedenti
ISA|55|11|sic erit verbum meum quod egredietur de ore meo non revertetur ad me vacuum sed faciet quaecumque volui et prosperabitur in his ad quae misi illud
ISA|55|12|quia in laetitia egrediemini et in pace deducemini montes et colles cantabunt coram vobis laudem et omnia ligna regionis plaudent manu
ISA|55|13|pro saliunca ascendet abies et pro urtica crescet myrtus et erit Dominus nominatus in signum aeternum quod non auferetur
ISA|56|1|haec dicit Dominus custodite iudicium et facite iustitiam quia iuxta est salus mea ut veniat et iustitia mea ut reveletur
ISA|56|2|beatus vir qui facit hoc et filius hominis qui adprehendit istud custodiens sabbatum ne polluat illud custodiens manus suas ne faciat omne malum
ISA|56|3|et non dicat filius advenae qui adheret Domino dicens separatione dividet me Dominus a populo suo et non dicat eunuchus ecce ego lignum aridum
ISA|56|4|quia haec dicit Dominus eunuchis qui custodierint sabbata mea et elegerint quae volui et tenuerint foedus meum
ISA|56|5|dabo eis in domo mea et in muris meis locum et nomen melius a filiis et filiabus nomen sempiternum dabo eis quod non peribit
ISA|56|6|et filios advenae qui adherent Domino ut colant eum et diligant nomen eius ut sint ei in servos omnem custodientem sabbatum ne polluat illud et tenentem foedus meum
ISA|56|7|adducam eos in montem sanctum meum et laetificabo eos in domo orationis meae holocausta eorum et victimae eorum placebunt mihi super altari meo quia domus mea domus orationis vocabitur cunctis populis
ISA|56|8|ait Dominus Deus qui congregat dispersos Israhel adhuc congregabo ad eum congregatos eius
ISA|56|9|omnes bestiae agri venite ad devorandum universae bestiae saltus
ISA|56|10|speculatores eius caeci omnes nescierunt universi canes muti non valentes latrare videntes vana dormientes et amantes somnia
ISA|56|11|et canes inpudentissimi nescierunt saturitatem ipsi pastores ignoraverunt intellegentiam omnes in viam suam declinaverunt unusquisque ad avaritiam suam a summo usque ad novissimum
ISA|56|12|venite sumamus vinum et impleamur ebrietate et erit sicut hodie sic et cras et multo amplius
ISA|57|1|iustus perit et nemo est qui recogitet in corde suo et viri misericordiae colliguntur quia non est qui intellegat a facie enim malitiae collectus est iustus
ISA|57|2|veniat pax requiescat in cubili suo qui ambulavit in directione sua
ISA|57|3|vos autem accedite huc filii auguratricis semen adulteri et fornicariae
ISA|57|4|super quem lusistis super quem dilatastis os et eiecistis linguam numquid non vos filii scelesti semen mendax
ISA|57|5|qui consolamini in diis subter omne lignum frondosum immolantes parvulos in torrentibus subter inminentes petras
ISA|57|6|in partibus torrentis pars tua haec est sors tua et ipsis effudisti libamen obtulisti sacrificium numquid super his non indignabor
ISA|57|7|super montem excelsum et sublimem posuisti cubile tuum et illuc ascendisti ut immolares hostias
ISA|57|8|et post ostium et retro postem posuisti memoriale tuum quia iuxta me discoperuisti et suscepisti adulterum dilatasti cubile tuum et pepigisti cum eis dilexisti stratum eorum manu aperta
ISA|57|9|et ornasti te regi unguento et multiplicasti pigmenta tua misisti legatos tuos procul et humiliata es usque ad inferos
ISA|57|10|in multitudine viae tuae laborasti non dixisti quiescam vitam manus tuae invenisti propterea non rogasti
ISA|57|11|pro quo sollicita timuisti quia mentita es et mei non es recordata neque cogitasti in corde tuo quia ego tacens et quasi non videns et mei oblita es
ISA|57|12|ego adnuntiabo iustitiam tuam et opera tua non proderunt tibi
ISA|57|13|cum clamaveris liberent te congregati tui et omnes eos auferet ventus tollet aura qui autem fiduciam habet mei hereditabit terram et possidebit montem sanctum meum
ISA|57|14|et dicam viam facite praebete iter declinate de semita auferte offendicula de via populi mei
ISA|57|15|quia haec dicit Excelsus et Sublimis habitans aeternitatem et sanctum nomen eius in excelso et in sancto habitans et cum contrito et humili spiritu ut vivificet spiritum humilium et vivificet cor contritorum
ISA|57|16|non enim in sempiternum litigabo neque usque ad finem irascar quia spiritus a facie mea egredietur et flatus ego faciam
ISA|57|17|propter iniquitatem avaritiae eius iratus sum et percussi eum abscondi et indignatus sum et abiit vagus in via cordis sui
ISA|57|18|vias eius vidi et dimisi eum et reduxi eum et reddidi consolationes ipsi et lugentibus eius
ISA|57|19|creavi fructum labiorum pacem pacem ei qui longe est et qui prope dixit Dominus et sanavi eum
ISA|57|20|impii autem quasi mare fervens quod quiescere non potest et redundant fluctus eius in conculcationem et lutum
ISA|57|21|non est pax dixit Deus meus impiis
ISA|58|1|clama ne cesses quasi tuba exalta vocem tuam et adnuntia populo meo scelera eorum et domui Iacob peccata eorum
ISA|58|2|me etenim de die in diem quaerunt et scire vias meas volunt quasi gens quae iustitiam fecerit et quae iudicium Dei sui non reliquerit rogant me iudicia iustitiae adpropinquare Deo volunt
ISA|58|3|quare ieiunavimus et non aspexisti humiliavimus animam nostram et nescisti ecce in die ieiunii vestri invenitur voluntas et omnes debitores vestros repetitis
ISA|58|4|ecce ad lites et contentiones ieiunatis et percutitis pugno impie nolite ieiunare sicut usque ad hanc diem ut audiatur in excelso clamor vester
ISA|58|5|numquid tale est ieiunium quod elegi per diem adfligere hominem animam suam numquid contorquere quasi circulum caput suum et saccum et cinerem sternere numquid istud vocabis ieiunium et diem acceptabilem Domino
ISA|58|6|nonne hoc est magis ieiunium quod elegi dissolve conligationes impietatis solve fasciculos deprimentes dimitte eos qui confracti sunt liberos et omne onus disrumpe
ISA|58|7|frange esurienti panem tuum et egenos vagosque induc in domum tuam cum videris nudum operi eum et carnem tuam ne despexeris
ISA|58|8|tunc erumpet quasi mane lumen tuum et sanitas tua citius orietur et anteibit faciem tuam iustitia tua et gloria Domini colliget te
ISA|58|9|tunc invocabis et Dominus exaudiet clamabis et dicet ecce adsum si abstuleris de medio tui catenam et desieris digitum extendere et loqui quod non prodest
ISA|58|10|cum effuderis esurienti animam tuam et animam adflictam repleveris orietur in tenebris lux tua et tenebrae tuae erunt sicut meridies
ISA|58|11|et requiem tibi dabit Dominus semper et implebit splendoribus animam tuam et ossa tua liberabit et eris quasi hortus inriguus et sicut fons aquarum cuius non deficient aquae
ISA|58|12|et aedificabuntur in te deserta saeculorum fundamenta generationis et generationis suscitabis et vocaberis aedificator sepium avertens semitas in quietem
ISA|58|13|si averteris a sabbato pedem tuum facere voluntatem tuam in die sancto meo et vocaveris sabbatum delicatum et sanctum Domini gloriosum et glorificaveris eum dum non facis vias tuas et non invenitur voluntas tua ut loquaris sermonem
ISA|58|14|tunc delectaberis super Domino et sustollam te super altitudines terrae et cibabo te hereditate Iacob patris tui os enim Domini locutum est
ISA|59|1|ecce non est adbreviata manus Domini ut salvare nequeat neque adgravata est auris eius ut non exaudiat
ISA|59|2|sed iniquitates vestrae diviserunt inter vos et Deum vestrum et peccata vestra absconderunt faciem eius a vobis ne exaudiret
ISA|59|3|manus enim vestrae pollutae sunt sanguine et digiti vestri iniquitate labia vestra locuta sunt mendacium et lingua vestra iniquitatem fatur
ISA|59|4|non est qui invocet iustitiam neque est qui iudicet vere sed confidunt in nihili et loquuntur vanitates conceperunt laborem et pepererunt iniquitatem
ISA|59|5|ova aspidum ruperunt et telas araneae texuerunt qui comederit de ovis eorum morietur et quod confotum est erumpet in regulum
ISA|59|6|telae eorum non erunt in vestimentum neque operientur operibus suis opera eorum opera inutilia et opus iniquitatis in manibus eorum
ISA|59|7|pedes eorum ad malum currunt et festinant ut effundant sanguinem innocentem cogitationes eorum cogitationes inutiles vastitas et contritio in viis eorum
ISA|59|8|viam pacis nescierunt et non est iudicium in gressibus eorum semitae eorum incurvatae sunt eis omnis qui calcat in ea ignorat pacem
ISA|59|9|propter hoc elongatum est iudicium a nobis et non adprehendet nos iustitia expectavimus lucem et ecce tenebrae splendorem et in tenebris ambulavimus
ISA|59|10|palpavimus sicut caeci parietem et quasi absque oculis adtrectavimus inpegimus meridie quasi in tenebris in caligosis quasi mortui
ISA|59|11|rugiemus quasi ursi omnes et quasi columbae meditantes gememus expectavimus iudicium et non est salutem et elongata est a nobis
ISA|59|12|multiplicatae sunt enim iniquitates nostrae coram te et peccata nostra responderunt nobis quia scelera nostra nobiscum et iniquitates nostras cognovimus
ISA|59|13|peccare et mentiri contra Dominum et aversi sumus ne iremus post tergum Dei nostri ut loqueremur calumniam et transgressionem concepimus et locuti sumus de corde verba mendacii
ISA|59|14|et conversum est retrorsum iudicium et iustitia longe stetit quia corruit in platea veritas et aequitas non potuit ingredi
ISA|59|15|et facta est veritas in oblivione et qui recessit a malo praedae patuit et vidit Dominus et malum apparuit in oculis eius quia non est iudicium
ISA|59|16|et vidit quia non est vir et aporiatus est quia non est qui occurrat et salvavit sibi brachium suum et iustitia eius ipsa confirmavit eum
ISA|59|17|indutus est iustitia ut lorica et galea salutis in capite eius indutus est vestimentis ultionis et opertus est quasi pallio zeli
ISA|59|18|sicut ad vindictam quasi ad retributionem indignationis hostibus suis et vicissitudinem inimicis suis insulis vicem reddet
ISA|59|19|et timebunt qui ab occidente nomen Domini et qui ab ortu solis gloriam eius cum venerit quasi fluvius violentus quem spiritus Domini cogit
ISA|59|20|et venerit Sion redemptor et eis qui redeunt ab iniquitate in Iacob dicit Dominus
ISA|59|21|hoc foedus meum cum eis dicit Dominus spiritus meus qui est in te et verba mea quae posui in ore tuo non recedent de ore tuo et de ore seminis tui et de ore seminis seminis tui dixit Dominus amodo et usque in sempiternum
ISA|60|1|surge inluminare quia venit lumen tuum et gloria Domini super te orta est
ISA|60|2|quia ecce tenebrae operient terram et caligo populos super te autem orietur Dominus et gloria eius in te videbitur
ISA|60|3|et ambulabunt gentes in lumine tuo et reges in splendore ortus tui
ISA|60|4|leva in circuitu oculos tuos et vide omnes isti congregati sunt venerunt tibi filii tui de longe venient et filiae tuae in latere sugent
ISA|60|5|tunc videbis et afflues et mirabitur et dilatabitur cor tuum quando conversa fuerit ad te multitudo maris fortitudo gentium venerit tibi
ISA|60|6|inundatio camelorum operiet te dromedariae Madian et Efa omnes de Saba venient aurum et tus deferentes et laudem Domino adnuntiantes
ISA|60|7|omne pecus Cedar congregabitur tibi arietes Nabaioth ministrabunt tibi offerentur super placabili altari meo et domum maiestatis meae glorificabo
ISA|60|8|qui sunt isti qui ut nubes volant et quasi columbae ad fenestras suas
ISA|60|9|me enim insulae expectant et naves maris in principio ut adducam filios tuos de longe argentum eorum et aurum eorum cum eis nomini Domini Dei tui et Sancto Israhel quia glorificavit te
ISA|60|10|et aedificabunt filii peregrinorum muros tuos et reges eorum ministrabunt tibi in indignatione enim mea percussi te et in reconciliatione mea misertus sum tui
ISA|60|11|et aperientur portae tuae iugiter die et nocte non claudentur ut adferatur ad te fortitudo gentium et reges earum adducantur
ISA|60|12|gens enim et regnum quod non servierit tibi peribit et gentes solitudine vastabuntur
ISA|60|13|gloria Libani ad te veniet abies et buxus et pinus simul ad ornandum locum sanctificationis meae et locum pedum meorum glorificabo
ISA|60|14|et venient ad te curvi filii eorum qui humiliaverunt te et adorabunt vestigia pedum tuorum omnes qui detrahebant tibi et vocabunt te civitatem Domini Sion Sancti Israhel
ISA|60|15|pro eo quod fuisti derelicta et odio habita et non erat qui per te transiret ponam te in superbiam saeculorum gaudium in generationem et generationem
ISA|60|16|et suges lac gentium et mamilla regum lactaberis et scies quia ego Dominus salvans te et redemptor tuus Fortis Iacob
ISA|60|17|pro aere adferam aurum et pro ferro adferam argentum et pro lignis aes et pro lapidibus ferrum et ponam visitationem tuam pacem et praepositos tuos iustitiam
ISA|60|18|non audietur ultra iniquitas in terra tua vastitas et contritio in terminis tuis et occupabit salus muros tuos et portas tuas laudatio
ISA|60|19|non erit tibi amplius sol ad lucendum per diem nec splendor lunae inluminabit te sed erit tibi Dominus in lucem sempiternam et Deus tuus in gloriam tuam
ISA|60|20|non occidet ultra sol tuus et luna tua non minuetur quia Dominus erit in lucem sempiternam et conplebuntur dies luctus tui
ISA|60|21|populus autem tuus omnes iusti in perpetuum hereditabunt terram germen plantationis meae opus manus meae ad glorificandum
ISA|60|22|minimus erit in mille et parvulus in gentem fortissimam ego Dominus in tempore eius subito faciam istud
ISA|61|1|spiritus Domini super me eo quod unxerit Dominus me ad adnuntiandum mansuetis misit me ut mederer contritis corde et praedicarem captivis indulgentiam et clausis apertionem
ISA|61|2|ut praedicarem annum placabilem Domini et diem ultionis Deo nostro ut consolarer omnes lugentes
ISA|61|3|ut ponerem lugentibus Sion et darem eis coronam pro cinere oleum gaudii pro luctu pallium laudis pro spiritu maeroris et vocabuntur in ea fortes iustitiae plantatio Domini ad glorificandum
ISA|61|4|et aedificabunt deserta a saeculo et ruinas antiquas erigent et instaurabunt civitates desertas dissipatas in generationem et generationem
ISA|61|5|et stabunt alieni et pascent pecora vestra et filii peregrinorum agricolae et vinitores vestri erunt
ISA|61|6|vos autem sacerdotes Domini vocabimini ministri Dei nostri dicetur vobis fortitudinem gentium comedetis et in gloria earum superbietis
ISA|61|7|pro confusione vestra duplici et rubore laudabunt partem eorum propter hoc in terra sua duplicia possidebunt laetitia sempiterna erit eis
ISA|61|8|quia ego Dominus diligens iudicium odio habens rapinam in holocausto et dabo opus eorum in veritate et foedus perpetuum feriam eis
ISA|61|9|et scietur in gentibus semen eorum et germen eorum in medio populorum omnes qui viderint eos cognoscent eos quia isti sunt semen cui benedixit Dominus
ISA|61|10|gaudens gaudebo in Domino et exultabit anima mea in Deo meo quia induit me vestimentis salutis et indumento iustitiae circumdedit me quasi sponsum decoratum corona et quasi sponsam ornatam monilibus suis
ISA|61|11|sicut enim terra profert germen suum et sicut hortus semen suum germinat sic Dominus Deus germinabit iustitiam et laudem coram universis gentibus
ISA|62|1|propter Sion non tacebo et propter Hierusalem non quiescam donec egrediatur ut splendor iustus eius et salvator eius ut lampas accendatur
ISA|62|2|et videbunt gentes iustum tuum et cuncti reges inclitum tuum et vocabitur tibi nomen novum quod os Domini nominabit
ISA|62|3|et eris corona gloriae in manu Domini et diadema regni in manu Dei tui
ISA|62|4|non vocaberis ultra Derelicta et terra tua non vocabitur amplius Desolata sed vocaberis Voluntas mea in ea et terra tua Inhabitata quia conplacuit Domino in te et terra tua inhabitabitur
ISA|62|5|habitabit enim iuvenis cum virgine et habitabunt in te filii tui et gaudebit sponsus super sponsam gaudebit super te Deus tuus
ISA|62|6|super muros tuos Hierusalem constitui custodes tota die et tota nocte perpetuo non tacebunt qui reminiscimini Domini ne taceatis
ISA|62|7|et ne detis silentium ei donec stabiliat et donec ponat Hierusalem laudem in terra
ISA|62|8|iuravit Dominus in dextera sua et in brachio fortitudinis suae si dedero triticum tuum ultra cibum inimicis tuis et si biberint filii alieni vinum tuum in quo laborasti
ISA|62|9|quia qui congregabunt illud comedent et laudabunt Dominum et qui conportant illud bibent in atriis sanctis meis
ISA|62|10|transite transite per portas praeparate viam populo planum facite iter et eligite lapides elevate signum ad populos
ISA|62|11|ecce Dominus auditum fecit in extremis terrae dicite filiae Sion ecce salvator tuus venit ecce merces eius cum eo et opus eius coram illo
ISA|62|12|et vocabunt eos Populus sanctus Redempti a Domino tu autem vocaberis Quaesita civitas et non Derelicta
ISA|63|1|quis est iste qui venit de Edom tinctis vestibus de Bosra iste formonsus in stola sua gradiens in multitudine fortitudinis suae ego qui loquor iustitiam et propugnator sum ad salvandum
ISA|63|2|quare ergo rubrum est indumentum tuum et vestimenta tua sicut calcantium in torculari
ISA|63|3|torcular calcavi solus et de gentibus non est vir mecum calcavi eos in furore meo et conculcavi eos in ira mea et aspersus est sanguis eorum super vestimenta mea et omnia indumenta mea inquinavi
ISA|63|4|dies enim ultionis in corde meo annus redemptionis meae venit
ISA|63|5|circumspexi et non erat auxiliator quaesivi et non fuit qui adiuvaret et salvavit mihi brachium meum et indignatio mea ipsa auxiliata est mihi
ISA|63|6|et conculcavi populos in furore meo et inebriavi eos in indignatione mea et detraxi in terra virtutem eorum
ISA|63|7|miserationum Domini recordabor laudem Domini super omnibus quae reddidit nobis Dominus et super multitudinem bonorum domui Israhel quae largitus est eis secundum indulgentiam suam et secundum multitudinem misericordiarum suarum
ISA|63|8|et dixit verumtamen populus meus est filii non negantes et factus est eis salvator
ISA|63|9|in omni tribulatione eorum non est tribulatus et angelus faciei eius salvavit eos in dilectione sua et in indulgentia sua ipse redemit eos et portavit eos et levavit eos cunctis diebus saeculi
ISA|63|10|ipsi autem ad iracundiam provocaverunt et adflixerunt spiritum Sancti eius et conversus est eis in inimicum et ipse debellavit eos
ISA|63|11|et recordatus est dierum saeculi Mosi populi sui ubi est qui eduxit eos de mari cum pastoribus gregis sui ubi est qui posuit in medio eius spiritum Sancti sui
ISA|63|12|qui eduxit ad dexteram Mosen brachio maiestatis suae qui scidit aquas ante eos ut faceret sibi nomen sempiternum
ISA|63|13|qui duxit eos per abyssos quasi equum in deserto non inpingentem
ISA|63|14|quasi animal in campo descendens spiritus Domini ductor eius fuit sic adduxisti populum tuum ut faceres tibi nomen gloriae
ISA|63|15|adtende de caelo et vide de habitaculo sancto tuo et gloriae tuae ubi est zelus tuus et fortitudo tua multitudo viscerum tuorum et miserationum tuarum super me continuerunt se
ISA|63|16|tu enim pater noster et Abraham nescivit nos et Israhel ignoravit nos tu Domine pater noster redemptor noster a saeculo nomen tuum
ISA|63|17|quare errare nos fecisti Domine de viis tuis indurasti cor nostrum ne timeremus te convertere propter servos tuos tribus hereditatis tuae
ISA|63|18|quasi nihilum possederunt populum sanctum tuum hostes nostri conculcaverunt sanctificationem tuam
ISA|63|19|facti sumus quasi in principio cum non dominareris nostri neque invocaretur nomen tuum super nos
ISA|64|1|utinam disrumperes caelos et descenderes a facie tua montes defluerent
ISA|64|2|sicut exustio ignis tabescerent aquae arderent igni ut notum fieret nomen tuum inimicis tuis a facie tua gentes turbarentur
ISA|64|3|cum feceris mirabilia non sustinebimus descendisti et a facie tua montes defluxerunt
ISA|64|4|a saeculo non audierunt neque auribus perceperunt oculus non vidit Deus absque te quae praeparasti expectantibus te
ISA|64|5|occurristi laetanti et facienti iustitiam in viis tuis recordabuntur tui ecce tu iratus es et peccavimus in ipsis fuimus semper et salvabimur
ISA|64|6|et facti sumus ut inmundus omnes nos quasi pannus menstruatae universae iustitiae nostrae et cecidimus quasi folium universi et iniquitates nostrae quasi ventus abstulerunt nos
ISA|64|7|non est qui invocet nomen tuum qui consurgat et teneat te abscondisti faciem tuam a nobis et adlisisti nos in manu iniquitatis nostrae
ISA|64|8|et nunc Domine pater noster es tu nos vero lutum et fictor noster et opera manuum tuarum omnes nos
ISA|64|9|ne irascaris Domine satis et ne ultra memineris iniquitatis ecce respice populus tuus omnes nos
ISA|64|10|civitas sancti tui facta est deserta Sion deserta facta est Hierusalem desolata
ISA|64|11|domus sanctificationis nostrae et gloriae nostrae ubi laudaverunt te patres nostri facta est in exustionem ignis et omnia desiderabilia nostra versa sunt in ruinas
ISA|64|12|numquid super his continebis te Domine tacebis et adfliges nos vehementer
ISA|65|1|quaesierunt me qui ante non interrogabant invenerunt qui non quaesierunt me dixi ecce ego ecce ego ad gentem quae non vocabat nomen meum
ISA|65|2|expandi manus meas tota die ad populum incredulum qui graditur in via non bona post cogitationes suas
ISA|65|3|populus qui ad iracundiam provocat me ante faciem meam semper qui immolant in hortis et sacrificant super lateres
ISA|65|4|qui habitant in sepulchris et in delubris idolorum dormiunt qui comedunt carnem suillam et ius profanum in vasis eorum
ISA|65|5|qui dicunt recede a me non adpropinques mihi quia inmundus es isti fumus erunt in furore meo ignis ardens tota die
ISA|65|6|ecce scriptum est coram me non tacebo sed reddam et retribuam in sinu eorum
ISA|65|7|iniquitates vestras et iniquitates patrum vestrorum simul dicit Dominus qui sacrificaverunt super montes et super colles exprobraverunt mihi et remetiar opus eorum primum in sinu eorum
ISA|65|8|haec dicit Dominus quomodo si inveniatur granum in botro et dicatur ne dissipes illud quoniam benedictio est sic faciam propter servos meos ut non disperdam totum
ISA|65|9|et educam de Iacob semen et de Iuda possidentem montes meos et hereditabunt eam electi mei et servi mei habitabunt ibi
ISA|65|10|et erunt campestria in caulas gregum et vallis Achor in cubile armentorum populo meo qui requisierunt me
ISA|65|11|et vos qui dereliquistis Dominum qui obliti estis montem sanctum meum qui ponitis Fortunae mensam et libatis super eam
ISA|65|12|numerabo vos in gladio et omnes in caede corruetis pro eo quod vocavi et non respondistis locutus sum et non audistis et faciebatis malum in oculis meis et quae nolui elegistis
ISA|65|13|propter hoc haec dicit Dominus Deus ecce servi mei comedent et vos esurietis ecce servi mei bibent et vos sitietis
ISA|65|14|ecce servi mei laetabuntur et vos confundemini ecce servi mei laudabunt prae exultatione cordis et vos clamabitis prae dolore cordis et prae contritione spiritus ululabitis
ISA|65|15|et dimittetis nomen vestrum in iuramentum electis meis et interficiet te Dominus Deus et servos suos vocabit nomine alio
ISA|65|16|in quo qui benedictus est super terram benedicetur in Deo amen et qui iurat in terra iurabit in Deo amen quia oblivioni traditae sunt angustiae priores et quia absconditae sunt ab oculis nostris
ISA|65|17|ecce enim ego creo caelos novos et terram novam et non erunt in memoria priora et non ascendent super cor
ISA|65|18|sed gaudebitis et exultabitis usque in sempiternum in his quae ego creo quia ecce ego creo Hierusalem exultationem et populum eius gaudium
ISA|65|19|et exultabo in Hierusalem et gaudebo in populo meo et non audietur in eo ultra vox fletus et vox clamoris
ISA|65|20|non erit ibi amplius infans dierum et senex qui non impleat dies suos quoniam puer centum annorum morietur et peccator centum annorum maledictus erit
ISA|65|21|et aedificabunt domos et habitabunt et plantabunt vineas et comedent fructum earum
ISA|65|22|non aedificabunt et alius habitabit non plantabunt et alius comedet secundum dies enim ligni erunt dies populi mei et opera manuum eorum inveterabunt
ISA|65|23|electis meis non laborabunt frustra neque generabunt in conturbatione quia semen benedictorum Domini est et nepotes eorum cum eis
ISA|65|24|eritque antequam clament ego exaudiam adhuc illis loquentibus ego audiam
ISA|65|25|lupus et agnus pascentur simul et leo et bos comedent paleas et serpenti pulvis panis eius non nocebunt neque occident in omni monte sancto meo dicit Dominus
ISA|66|1|haec dicit Dominus caelum sedis mea et terra scabillum pedum meorum quae ista domus quam aedificabitis mihi et quis iste locus quietis meae
ISA|66|2|omnia haec manus mea fecit et facta sunt universa ista dicit Dominus ad quem autem respiciam nisi ad pauperculum et contritum spiritu et trementem sermones meos
ISA|66|3|qui immolat bovem quasi qui interficiat virum qui mactat pecus quasi qui excerebret canem qui offert oblationem quasi qui sanguinem suillum offerat qui recordatur turis quasi qui benedicat idolo haec omnia elegerunt in viis suis et in abominationibus suis anima eorum delectata est
ISA|66|4|unde et ego eligam inlusiones eorum et quae timebant adducam eis quia vocavi et non erat qui responderet locutus sum et non audierunt feceruntque malum in oculis meis et quae nolui elegerunt
ISA|66|5|audite verbum Domini qui tremetis ad verbum eius dixerunt fratres vestri odientes vos et abicientes propter nomen meum glorificetur Dominus et videbimus in laetitia vestra ipsi autem confundentur
ISA|66|6|vox populi de civitate vox de templo vox Domini reddentis retributionem inimicis suis
ISA|66|7|antequam parturiret peperit antequam veniret partus eius peperit masculum
ISA|66|8|quis audivit umquam tale et quis vidit huic simile numquid parturiet terra in die una aut parietur gens simul quia parturivit et peperit Sion filios suos
ISA|66|9|numquid ego qui alios parere facio ipse non pariam dicit Dominus si ego qui generationem ceteris tribuo sterilis ero ait Dominus Deus tuus
ISA|66|10|laetamini cum Hierusalem et exultate in ea omnes qui diligitis eam gaudete cum ea gaudio universi qui lugetis super eam
ISA|66|11|ut sugatis et repleamini ab ubere consolationis eius ut mulgeatis et deliciis affluatis ab omnimoda gloria eius
ISA|66|12|quia haec dicit Dominus ecce ego declinabo super eam quasi fluvium pacis et quasi torrentem inundantem gloriam gentium quam sugetis ad ubera portabimini et super genua blandientur vobis
ISA|66|13|quomodo si cui mater blandiatur ita ego consolabor vos et in Hierusalem consolabimini
ISA|66|14|videbitis et gaudebit cor vestrum et ossa vestra quasi herba germinabunt et cognoscetur manus Domini servis eius et indignabitur inimicis suis
ISA|66|15|quia ecce Dominus in igne veniet et quasi turbo quadrigae eius reddere in indignatione furorem suum et increpationem suam in flamma ignis
ISA|66|16|quia in igne Dominus diiudicatur et in gladio suo ad omnem carnem et multiplicabuntur interfecti a Domino
ISA|66|17|qui sanctificabantur et mundos se putabant in hortis post unam intrinsecus qui comedebant carnem suillam et abominationem et murem simul consumentur dicit Dominus
ISA|66|18|ego autem opera eorum et cogitationes eorum venio ut congregem cum omnibus gentibus et linguis et venient et videbunt gloriam meam
ISA|66|19|et ponam in eis signum et mittam ex eis qui salvati fuerint ad gentes in mari in Africa in Lydia tenentes sagittam in Italiam et Graeciam ad insulas longe ad eos qui non audierunt de me et non viderunt gloriam meam et adnuntiabunt gloriam meam gentibus
ISA|66|20|et adducent omnes fratres vestros de cunctis gentibus donum Domino in equis et in quadrigis et in lecticis et in mulis et in carrucis ad montem sanctum meum Hierusalem dicit Dominus quomodo si inferant filii Israhel munus in vase mundo in domum Domini
ISA|66|21|et adsumam ex eis in sacerdotes et in Levitas dicit Dominus
ISA|66|22|quia sicut caeli novi et terra nova quae ego facio stare coram me dicit Dominus sic stabit semen vestrum et nomen vestrum
ISA|66|23|et erit mensis ex mense et sabbatum ex sabbato veniet omnis caro ut adoret coram facie mea dicit Dominus
ISA|66|24|et egredientur et videbunt cadavera virorum qui praevaricati sunt in me vermis eorum non morietur et ignis eorum non extinguetur et erunt usque ad satietatem visionis omni carni
JER|1|1|verba Hieremiae filii Helciae de sacerdotibus qui fuerunt in Anathoth in terra Beniamin
JER|1|2|quod factum est verbum Domini ad eum in diebus Iosiae filii Amon regis Iuda in tertiodecimo anno regni eius
JER|1|3|et factum est in diebus Ioachim filii Iosiae regis Iuda usque ad consummationem undecimi anni Sedeciae filii Iosiae regis Iuda usque ad transmigrationem Hierusalem in mense quinto
JER|1|4|et factum est verbum Domini ad me dicens
JER|1|5|priusquam te formarem in utero novi te et antequam exires de vulva sanctificavi te prophetam gentibus dedi te
JER|1|6|et dixi a a a Domine Deus ecce nescio loqui quia puer ego sum
JER|1|7|et dixit Dominus ad me noli dicere puer sum quoniam ad omnia quae mittam te ibis et universa quaecumque mandavero tibi loqueris
JER|1|8|ne timeas a facie eorum quia tecum ego sum ut eruam te dicit Dominus
JER|1|9|et misit Dominus manum suam et tetigit os meum et dixit Dominus ad me ecce dedi verba mea in ore tuo
JER|1|10|ecce constitui te hodie super gentes et super regna ut evellas et destruas et disperdas et dissipes et aedifices et plantes
JER|1|11|et factum est verbum Domini ad me dicens quid tu vides Hieremia et dixi virgam vigilantem ego video
JER|1|12|et dixit Dominus ad me bene vidisti quia vigilabo ego super verbo meo ut faciam illud
JER|1|13|et factum est verbum Domini secundo ad me dicens quid tu vides et dixi ollam succensam ego video et faciem eius a facie aquilonis
JER|1|14|et dixit Dominus ad me ab aquilone pandetur malum super omnes habitatores terrae
JER|1|15|quia ecce ego convocabo omnes cognationes regnorum aquilonis ait Dominus et venient et ponent unusquisque solium suum in introitu portarum Hierusalem et super omnes muros eius in circuitu et super universas urbes Iuda
JER|1|16|et loquar iudicia mea cum eis super omni malitia eorum qui dereliquerunt me et libaverunt diis alienis et adoraverunt opus manuum suarum
JER|1|17|tu ergo accinge lumbos tuos et surge et loquere ad eos omnia quae ego praecipio tibi ne formides a facie eorum nec enim timere te faciam vultum eorum
JER|1|18|ego quippe dedi te hodie in civitatem munitam et in columnam ferream et in murum aereum super omnem terram regibus Iuda principibus eius et sacerdotibus et populo terrae
JER|1|19|et bellabunt adversum te et non praevalebunt quia tecum ego sum ait Dominus ut liberem te
JER|2|1|et factum est verbum Domini ad me dicens
JER|2|2|vade et clama in auribus Hierusalem dicens haec dicit Dominus recordatus sum tui miserans adulescentiam tuam et caritatem disponsationis tuae quando secuta me es in deserto in terra quae non seminatur
JER|2|3|sanctus Israhel Domino primitiae frugum eius omnes qui devorant eum delinquunt mala venient super eos dicit Dominus
JER|2|4|audite verbum Domini domus Iacob et omnes cognationes domus Israhel
JER|2|5|haec dicit Dominus quid invenerunt patres vestri in me iniquitatis quia elongaverunt a me et ambulaverunt post vanitatem et vani facti sunt
JER|2|6|et non dixerunt ubi est Dominus qui ascendere nos fecit de terra Aegypti qui transduxit nos per desertum per terram inhabitabilem et inviam per terram sitis et imaginem mortis per terram in qua non ambulavit vir neque habitavit homo
JER|2|7|et induxi vos in terram Carmeli ut comederetis fructum eius et optima illius et ingressi contaminastis terram meam et hereditatem meam posuistis in abominationem
JER|2|8|sacerdotes non dixerunt ubi est Dominus et tenentes legem nescierunt me et pastores praevaricati sunt in me et prophetae prophetaverunt in Baal et idola secuti sunt
JER|2|9|propterea adhuc iudicio contendam vobiscum ait Dominus et cum filiis vestris disceptabo
JER|2|10|transite ad insulas Cetthim et videte et in Cedar mittite et considerate vehementer et videte si factum est huiuscemodi
JER|2|11|si mutavit gens deos et certe ipsi non sunt dii populus vero meus mutavit Gloriam suam in idolum
JER|2|12|obstupescite caeli super hoc et portae eius desolamini vehementer dicit Dominus
JER|2|13|duo enim mala fecit populus meus me dereliquerunt fontem aquae vivae ut foderent sibi cisternas cisternas dissipatas quae continere non valent aquas
JER|2|14|numquid servus est Israhel aut vernaculus quare ergo est factus in praedam
JER|2|15|super eum rugierunt leones et dederunt vocem suam posuerunt terram eius in solitudinem civitates eius exustae sunt et non est qui habitet in eis
JER|2|16|filii quoque Memfeos et Tafnes constupraverunt te usque ad verticem
JER|2|17|numquid non istud factum est tibi quia dereliquisti Dominum Deum tuum eo tempore quo ducebat te per viam
JER|2|18|et nunc quid tibi vis in via Aegypti ut bibas aquam turbidam et quid tibi cum via Assyriorum ut bibas aquam Fluminis
JER|2|19|arguet te malitia tua et aversio tua increpabit te scito et vide quia malum et amarum est reliquisse te Dominum Deum tuum et non esse timorem mei apud te dicit Dominus Deus exercituum
JER|2|20|a saeculo confregisti iugum meum rupisti vincula mea et dixisti non serviam in omni enim colle sublimi et sub omni ligno frondoso tu prosternebaris meretrix
JER|2|21|ego autem plantavi te vineam electam omne semen verum quomodo ergo conversa es in pravum vinea aliena
JER|2|22|si laveris te nitro et multiplicaveris tibi herbam borith maculata es in iniquitate tua coram me dicit Dominus Deus
JER|2|23|quomodo dicis non sum polluta post Baalim non ambulavi vide vias tuas in convalle scito quid feceris cursor levis explicans vias tuas
JER|2|24|onager adsuetus in solitudine in desiderio animae suae adtraxit ventum amoris sui nullus avertet eam omnes qui quaerunt eam non deficient in menstruis eius invenient eam
JER|2|25|prohibe pedem tuum a nuditate et guttur tuum a siti et dixisti desperavi nequaquam faciam adamavi quippe alienos et post eos ambulabo
JER|2|26|quomodo confunditur fur quando deprehenditur sic confusi sunt domus Israhel ipsi et reges eorum principes et sacerdotes et prophetae eorum
JER|2|27|dicentes ligno pater meus es tu et lapidi tu me genuisti verterunt ad me tergum et non faciem et in tempore adflictionis suae dicent surge et libera nos
JER|2|28|ubi sunt dii tui quos fecisti tibi surgant et liberent te in tempore adflictionis tuae secundum numerum quippe civitatum tuarum erant dii tui Iuda
JER|2|29|quid vultis mecum iudicio contendere omnes dereliquistis me dicit Dominus
JER|2|30|frustra percussi filios vestros disciplinam non receperunt devoravit gladius vester prophetas vestros quasi leo vastator
JER|2|31|generatio vestra videte verbum Domini numquid solitudo factus sum Israheli aut terra serotina quare ergo dixit populus meus recessimus non veniemus ultra ad te
JER|2|32|numquid obliviscitur virgo ornamenti sui sponsa fasciae pectoralis suae populus vero meus oblitus est mei diebus innumeris
JER|2|33|quid niteris bonam ostendere viam tuam ad quaerendam dilectionem quae insuper et malitias tuas docuisti vias tuas
JER|2|34|et in alis tuis inventus est sanguis animarum pauperum et innocentium non in fossis inveni eos sed in omnibus quae supra memoravi
JER|2|35|et dixisti absque peccato et innocens ego sum et propterea avertatur furor tuus a me ecce ego iudicio contendam tecum eo quod dixeris non peccavi
JER|2|36|quam vilis es facta nimis iterans vias tuas et ab Aegypto confunderis sicut confusa es ab Assur
JER|2|37|nam et ab ista egredieris et manus tuae erunt super caput tuum quoniam obtrivit Dominus confidentiam tuam et nihil habebis prosperum
JER|3|1|vulgo dicitur si dimiserit vir uxorem suam et recedens ab eo duxerit virum alterum numquid revertetur ad eam ultra numquid non polluta et contaminata erit mulier illa tu autem fornicata es cum amatoribus multis tamen revertere ad me dicit Dominus
JER|3|2|leva oculos tuos in directum et vide ubi non prostrata sis in viis sedebas expectans eos quasi latro in solitudine et polluisti terram in fornicationibus tuis et in malitiis tuis
JER|3|3|quam ob rem prohibitae sunt stillae pluviarum et serotinus imber non fuit frons mulieris meretricis facta est tibi noluisti erubescere
JER|3|4|ergo saltim amodo voca me pater meus dux virginitatis meae tu es
JER|3|5|numquid irasceris in perpetuum aut perseverabis in finem ecce locuta es et fecisti mala et potuisti
JER|3|6|et dixit Dominus ad me in diebus Iosiae regis numquid vidisti quae fecerit aversatrix Israhel abiit sibimet super omnem montem excelsum et sub omne lignum frondosum et fornicata est ibi
JER|3|7|et dixi cum fecisset haec omnia ad me convertere et non est reversa et vidit praevaricatrix soror eius Iuda
JER|3|8|quia pro eo quod moechata esset aversatrix Israhel dimisissem eam et dedissem ei libellum repudii et non timuit praevaricatrix Iuda soror eius sed abiit et fornicata est etiam ipsa
JER|3|9|et facilitate fornicationis suae contaminavit terram et moechata est cum lapide et cum ligno
JER|3|10|et in omnibus his non est reversa ad me praevaricatrix soror eius Iuda in toto corde suo sed in mendacio ait Dominus
JER|3|11|et dixit Dominus ad me iustificavit animam suam aversatrix Israhel conparatione praevaricatricis Iuda
JER|3|12|vade et clama sermones istos contra aquilonem et dices revertere aversatrix Israhel ait Dominus et non avertam faciem meam a vobis quia sanctus ego sum dicit Dominus et non irascar in perpetuum
JER|3|13|tamen scito iniquitatem tuam quia in Dominum Deum tuum praevaricata es et dispersisti vias tuas alienis sub omni ligno frondoso et vocem meam non audisti ait Dominus
JER|3|14|convertimini filii revertentes dicit Dominus quia ego vir vester et adsumam vos unum de civitate et duos de cognatione et introducam vos in Sion
JER|3|15|et dabo vobis pastores iuxta cor meum et pascent vos scientia et doctrina
JER|3|16|cumque multiplicati fueritis et creveritis in terra in diebus illis ait Dominus non dicent ultra arca testamenti Domini neque ascendet super cor neque recordabuntur illius nec visitabitur nec fiet ultra
JER|3|17|in tempore illo vocabunt Hierusalem solium Domini et congregabuntur ad eam omnes gentes in nomine Domini in Hierusalem et non ambulabunt post pravitatem cordis sui pessimi
JER|3|18|in diebus illis ibit domus Iuda ad domum Israhel et venient simul de terra aquilonis ad terram quam dedi patribus vestris
JER|3|19|ego autem dixi quomodo ponam te in filiis et tribuam tibi terram desiderabilem hereditatem praeclaram exercituum gentium et dixi patrem vocabis me et post me ingredi non cessabis
JER|3|20|sed quomodo si contemnat mulier amatorem suum sic contempsit me domus Israhel dicit Dominus
JER|3|21|vox in viis audita est ploratus et ululatus filiorum Israhel quoniam iniquam fecerunt viam suam obliti sunt Domini Dei sui
JER|3|22|convertimini filii revertentes et sanabo aversiones vestras ecce nos venimus ad te tu enim es Dominus Deus noster
JER|3|23|vere mendaces erant colles multitudo montium vere in Domino Deo nostro salus Israhel
JER|3|24|confusio comedit laborem patrum nostrorum ab adulescentia nostra greges eorum et armenta eorum filios eorum et filias eorum
JER|3|25|dormiemus in confusione nostra et operiet nos ignominia nostra quoniam Domino Deo nostro peccavimus nos et patres nostri ab adulescentia nostra usque ad hanc diem et non audivimus vocem Domini Dei nostri
JER|4|1|si converteris Israhel ait Dominus ad me convertere si abstuleris offendicula tua a facie mea non commoveberis
JER|4|2|et iurabis vivit Dominus in veritate et in iudicio et in iustitia et benedicent eum gentes ipsumque laudabunt
JER|4|3|haec enim dicit Dominus viro Iuda et Hierusalem novate vobis novale et nolite serere super spinas
JER|4|4|circumcidimini Domino et auferte praeputia cordium vestrorum vir Iuda et habitatores Hierusalem ne forte egrediatur ut ignis indignatio mea et succendatur et non sit qui extinguat propter malitiam cogitationum vestrarum
JER|4|5|adnuntiate in Iuda et in Hierusalem auditum facite loquimini et canite tuba in terra clamate fortiter dicite congregamini et ingrediamur civitates munitas
JER|4|6|levate signum in Sion confortamini nolite stare quia malum ego adduco ab aquilone et contritionem magnam
JER|4|7|ascendit leo de cubili suo et praedo gentium se levavit egressus est de loco suo ut ponat terram tuam in desolationem civitates tuae vastabuntur remanentes absque habitatore
JER|4|8|super hoc accingite vos ciliciis plangite et ululate quia non est aversa ira furoris Domini a nobis
JER|4|9|et erit in die illa dicit Dominus peribit cor regis et cor principum et obstupescent sacerdotes et prophetae consternabuntur
JER|4|10|et dixi heu heu heu Domine Deus ergone decepisti populum istum et Hierusalem dicens pax erit vobis et ecce pervenit gladius usque ad animam
JER|4|11|in tempore illo dicetur populo huic et Hierusalem ventus urens in viis quae sunt in deserto viae filiae populi mei non ad ventilandum et ad purgandum
JER|4|12|spiritus plenus ex his veniet mihi et nunc ego sed loquar iudicia mea cum eis
JER|4|13|ecce quasi nubes ascendet et quasi tempestas currus eius velociores aquilis equi illius vae nobis quoniam vastati sumus
JER|4|14|lava a malitia cor tuum Hierusalem ut salva fias usquequo morabuntur in te cogitationes noxiae
JER|4|15|vox enim adnuntiantis a Dan et notum facientis idolum de monte Ephraim
JER|4|16|concitate gentes ecce auditum est in Hierusalem custodes venire de terra longinqua et dare super civitates Iuda vocem suam
JER|4|17|quasi custodes agrorum facti sunt super eam in gyro quia me ad iracundiam provocavit ait Dominus
JER|4|18|viae tuae et cogitationes tuae fecerunt haec tibi ista malitia tua quia amara quia tetigit cor tuum
JER|4|19|ventrem meum ventrem meum doleo sensus cordis mei turbati sunt in me non tacebo quoniam vocem bucinae audivit anima mea clamorem proelii
JER|4|20|contritio super contritionem vocata est et vastata est omnis terra repente vastata sunt tabernacula mea subito pelles meae
JER|4|21|usquequo videbo fugientem audiam vocem bucinae
JER|4|22|quia stultus populus meus me non cognovit filii insipientes sunt et vecordes sapientes sunt ut faciant mala bene autem facere nescierunt
JER|4|23|aspexi terram et ecce vacua erat et nihili et caelos et non erat lux in eis
JER|4|24|vidi montes et ecce movebantur et omnes colles conturbati sunt
JER|4|25|intuitus sum et non erat homo et omne volatile caeli recessit
JER|4|26|aspexi et ecce Carmelus desertus et omnes urbes eius destructae sunt a facie Domini et a facie irae furoris eius
JER|4|27|haec enim dicit Dominus deserta erit omnis terra sed tamen consummationem non faciam
JER|4|28|lugebit terra et maerebunt caeli desuper eo quod locutus sum cogitavi et non paenituit me nec aversus sum ab eo
JER|4|29|a voce equitis et mittentis sagittam fugit omnis civitas ingressi sunt ardua et ascenderunt rupes universae urbes derelictae sunt et non habitat in eis homo
JER|4|30|tu autem vastata quid facies cum vestieris te coccino cum ornata fueris monili aureo et pinxeris stibio oculos tuos frustra conponeris contempserunt te amatores tui animam tuam quaerent
JER|4|31|vocem enim quasi parturientis audivi angustias ut puerperae vox filiae Sion intermorientis expandentisque manus suas vae mihi quia defecit anima mea propter interfectos
JER|5|1|circuite vias Hierusalem et aspicite et considerate et quaerite in plateis eius an inveniatis virum facientem iudicium et quaerentem fidem et propitius ero eius
JER|5|2|quod si etiam vivit Dominus dixerint et hoc falso iurabunt
JER|5|3|Domine oculi tui respiciunt fidem percussisti eos et non doluerunt adtrivisti eos et rennuerunt accipere disciplinam induraverunt facies suas super petram noluerunt reverti
JER|5|4|ego autem dixi forsitan pauperes sunt et stulti ignorantes viam Domini iudicium Dei sui
JER|5|5|ibo igitur ad optimates et loquar eis ipsi enim cognoverunt viam Domini iudicium Dei sui et ecce magis hii simul confregerunt iugum ruperunt vincula
JER|5|6|idcirco percussit eos leo de silva lupus ad vesperam vastavit eos pardus vigilans super civitates eorum omnis qui egressus fuerit ex eis capietur quia multiplicatae sunt praevaricationes eorum confortatae sunt aversiones eorum
JER|5|7|super quo propitius tibi esse potero filii tui dereliquerunt me et iurant in his qui non sunt dii saturavi eos et moechati sunt et in domo meretricis luxuriabantur
JER|5|8|equi amatores et admissarii facti sunt unusquisque ad uxorem proximi sui hinniebat
JER|5|9|numquid super his non visitabo dicit Dominus et in gente tali non ulciscetur anima mea
JER|5|10|ascendite muros eius et dissipate consummationem autem nolite facere auferte propagines eius quia non sunt Domini
JER|5|11|praevaricatione enim praevaricata est in me domus Israhel et domus Iuda ait Dominus
JER|5|12|negaverunt Dominum et dixerunt non est ipse neque veniet super nos malum gladium et famem non videbimus
JER|5|13|prophetae fuerunt in ventum et responsum non fuit in eis haec ergo evenient illis
JER|5|14|haec dicit Dominus Deus exercituum quia locuti estis verbum istud ecce ego do verba mea in ore tuo in ignem et populum istum ligna et vorabit eos
JER|5|15|ecce ego adducam super vos gentem de longinquo domus Israhel ait Dominus gentem robustam gentem antiquam gentem cuius ignorabis linguam nec intelleges quid loquatur
JER|5|16|faretra eius quasi sepulchrum patens universi fortes
JER|5|17|et comedet segetes tuas et panem tuum devorabit filios tuos et filias tuas comedet gregem tuum et armenta tua comedet vineam tuam et ficum tuam et conteret urbes munitas tuas in quibus tu habes fiduciam gladio
JER|5|18|verumtamen et diebus illis ait Dominus non faciam vos in consummationem
JER|5|19|quod si dixeritis quare fecit Dominus Deus noster nobis haec omnia dices ad eos sicut dereliquistis me et servistis deo alieno in terra vestra sic servietis alienis in terra non vestra
JER|5|20|adnuntiate hoc domui Iacob et auditum facite in Iuda dicentes
JER|5|21|audi populus stulte qui non habes cor qui habentes oculos non videtis et aures et non auditis
JER|5|22|me ergo non timebitis ait Dominus et a facie mea non dolebitis qui posui harenam terminum mari praeceptum sempiternum quod non praeteribit et commovebuntur et non poterunt et intumescent fluctus eius et non transibunt illud
JER|5|23|populo autem huic factum est cor incredulum et exasperans recesserunt et abierunt
JER|5|24|et non dixerunt in corde suo metuamus Dominum Deum nostrum qui dat nobis pluviam temporaneam et serotinam in tempore suo plenitudinem annuae messis custodientem nobis
JER|5|25|iniquitates nostrae declinaverunt haec et peccata nostra prohibuerunt bonum a nobis
JER|5|26|quia inventi sunt in populo meo impii insidiantes quasi aucupes laqueos ponentes et pedicas ad capiendos viros
JER|5|27|sicut decipula plena avibus sic domus eorum plenae dolo ideo magnificati sunt et ditati
JER|5|28|incrassati sunt et inpinguati et praeterierunt sermones meos pessime causam non iudicaverunt causam pupilli non direxerunt et iudicium pauperum non iudicaverunt
JER|5|29|numquid super his non visitabo dicit Dominus aut super gentem huiuscemodi non ulciscetur anima mea
JER|5|30|stupor et mirabilia facta sunt in terra
JER|5|31|prophetae prophetabant mendacium et sacerdotes adplaudebant manibus suis et populus meus dilexit talia quid igitur fiet in novissimo eius
JER|6|1|confortamini filii Beniamin in medio Hierusalem et in Thecua clangite bucina et super Bethaccharem levate vexillum quia malum visum est ab aquilone et contritio magna
JER|6|2|speciosae et delicatae adsimilavi filiam Sion
JER|6|3|ad eam venient pastores et greges eorum fixerunt in ea tentoria in circuitu pascet unusquisque eos qui sub manu sua sunt
JER|6|4|sanctificate super eam bellum consurgite et ascendamus in meridie vae nobis quia declinavit dies quia longiores factae sunt umbrae vesperi
JER|6|5|surgite et ascendamus in nocte et dissipemus domos eius
JER|6|6|quia haec dicit Dominus exercituum caedite lignum eius et fundite circa Hierusalem aggerem haec est civitas visitationis omnis calumnia in medio eius
JER|6|7|sicut frigidam facit cisterna aquam suam sic frigidam fecit malitiam suam iniquitas et vastitas audietur in ea coram me semper infirmitas et plaga
JER|6|8|erudire Hierusalem ne forte recedat anima mea a te ne forte ponam te desertam terram inhabitabilem
JER|6|9|haec dicit Dominus exercituum usque ad racemum colligent quasi in vinea reliquias Israhel converte manum tuam quasi vindemiator ad cartallum
JER|6|10|cui loquar et quem contestabor ut audiant ecce incircumcisae aures eorum et audire non possunt ecce verbum Domini factum est eis in obprobrium et non suscipient illud
JER|6|11|idcirco furore Domini plenus sum laboravi sustinens effunde super parvulum foris et super concilium iuvenum simul vir enim cum muliere capietur senex cum pleno dierum
JER|6|12|et transibunt domus eorum ad alteros agri et uxores pariter quia extendam manum meam super habitantes terram dicit Dominus
JER|6|13|a minore quippe usque ad maiorem omnes avaritiae student et a propheta usque ad sacerdotem cuncti faciunt dolum
JER|6|14|et curabant contritionem filiae populi mei cum ignominia dicentes pax pax et non erat pax
JER|6|15|confusi sunt quia abominationem fecerunt quin potius confusione non sunt confusi et erubescere nescierunt quam ob rem cadent inter ruentes in tempore visitationis suae corruent dicit Dominus
JER|6|16|haec dicit Dominus state super vias et videte et interrogate de semitis antiquis quae sit via bona et ambulate in ea et invenietis refrigerium animabus vestris et dixerunt non ambulabimus
JER|6|17|et constitui super vos speculatores audite vocem tubae et dixerunt non audiemus
JER|6|18|ideo audite gentes et cognosce congregatio quanta ego faciam eis
JER|6|19|audi terra ecce ego adducam mala super populum istum fructum cogitationum eius quia verba mea non audierunt et legem meam proiecerunt
JER|6|20|ut quid mihi tus de Saba adfertis et calamum suave olentem de terra longinqua holocaustomata vestra non sunt accepta et victimae vestrae non placuerunt mihi
JER|6|21|propterea haec dicit Dominus ecce ego dabo in populum istum ruinas et ruent in eis patres et filii simul vicinus et proximus et peribunt
JER|6|22|haec dicit Dominus ecce populus venit de terra aquilonis et gens magna consurget a finibus terrae
JER|6|23|sagittam et scutum arripiet crudelis est et non miserebitur vox eius quasi mare sonabit et super equos ascendent praeparati quasi vir ad proelium adversum te filia Sion
JER|6|24|audivimus famam eius dissolutae sunt manus nostrae tribulatio adprehendit nos dolores ut parturientem
JER|6|25|nolite exire ad agros et in via ne ambuletis quoniam gladius inimici pavor in circuitu
JER|6|26|filia populi mei accingere cilicio et conspergere cinere luctum unigeniti fac tibi planctum amarum quia repente veniet vastator super nos
JER|6|27|probatorem dedi te in populo meo robustum et scies et probabis viam eorum
JER|6|28|omnes isti principes declinantum ambulantes fraudulenter aes et ferrum universi corrupti sunt
JER|6|29|defecit sufflatorium in igne consumptum est plumbum frustra conflavit conflator malitiae enim eorum non sunt consumptae
JER|6|30|argentum reprobum vocate eos quia Dominus proiecit illos
JER|7|1|verbum quod factum est ad Hieremiam a Domino dicens
JER|7|2|sta in porta domus Domini et praedica ibi verbum istud et dic audite verbum Domini omnis Iuda qui ingredimini per portas has ut adoretis Dominum
JER|7|3|haec dicit Dominus exercituum Deus Israhel bonas facite vias vestras et studia vestra et habitabo vobiscum in loco isto
JER|7|4|nolite confidere in verbis mendacii dicentes templum Domini templum Domini templum Domini est
JER|7|5|quoniam si bene direxeritis vias vestras et studia vestra si feceritis iudicium inter virum et proximum eius
JER|7|6|advenae et pupillo et viduae non feceritis calumniam nec sanguinem innocentem effuderitis in loco hoc et post deos alienos non ambulaveritis in malum vobismet ipsis
JER|7|7|habitabo vobiscum in loco isto in terra quam dedi patribus vestris a saeculo usque in saeculum
JER|7|8|ecce vos confiditis vobis in sermonibus mendacii qui non proderunt vobis
JER|7|9|furari occidere adulterare iurare mendaciter libare Baali et ire post deos alienos quos ignoratis
JER|7|10|et venistis et stetistis coram me in domo hac in qua invocatum est nomen meum et dixistis liberati sumus eo quod fecerimus omnes abominationes istas
JER|7|11|ergo spelunca latronum facta est domus ista in qua invocatum est nomen meum in oculis vestris ego ego sum ego vidi dicit Dominus
JER|7|12|ite ad locum meum in Silo ubi habitavit nomen meum a principio et videte quae fecerim ei propter malitiam populi mei Israhel
JER|7|13|et nunc quia fecistis omnia opera haec dicit Dominus et locutus sum ad vos mane consurgens et loquens et non audistis et vocavi vos et non respondistis
JER|7|14|faciam domui huic in qua invocatum est nomen meum et in qua vos habetis fiduciam et loco quem dedi vobis et patribus vestris sicut feci Silo
JER|7|15|et proiciam vos a facie mea sicut proieci omnes fratres vestros universum semen Ephraim
JER|7|16|tu ergo noli orare pro populo hoc nec adsumas pro eis laudem et orationem et non obsistas mihi quia non exaudiam te
JER|7|17|nonne vides quid isti faciant in civitatibus Iuda et in plateis Hierusalem
JER|7|18|filii colligunt ligna et patres succendunt ignem et mulieres conspergunt adipem ut faciant placentas Reginae caeli et libent diis alienis et me ad iracundiam provocent
JER|7|19|numquid me ad iracundiam provocant dicit Dominus nonne semet ipsos in confusionem vultus sui
JER|7|20|ideo haec dicit Dominus Deus ecce furor meus et indignatio mea conflatur super locum istum super viros et super iumenta et super lignum regionis et super fruges terrae et succendetur et non extinguetur
JER|7|21|haec dicit Dominus exercituum Deus Israhel holocaustomata vestra addite victimis vestris et comedite carnes
JER|7|22|quia non sum locutus cum patribus vestris et non praecepi eis in die qua eduxi eos de terra Aegypti de verbo holocaustomatum et victimarum
JER|7|23|sed hoc verbum praecepi eis dicens audite vocem meam et ero vobis Deus et vos eritis mihi populus et ambulate in omni via quam mandavi vobis ut bene sit vobis
JER|7|24|et non audierunt nec inclinaverunt aurem suam sed abierunt in voluntatibus et pravitate cordis sui mali factique sunt retrorsum et non in ante
JER|7|25|a die qua egressi sunt patres eorum de terra Aegypti usque ad diem hanc et misi ad vos omnes servos meos prophetas per diem consurgens diluculo et mittens
JER|7|26|et non audierunt me nec inclinaverunt aurem suam sed induraverunt cervicem et peius operati sunt quam patres eorum
JER|7|27|et loqueris ad eos omnia verba haec et non audient te et vocabis eos et non respondebunt tibi
JER|7|28|et dices ad eos haec est gens quae non audivit vocem Domini Dei sui nec recepit disciplinam periit fides et ablata est de ore eorum
JER|7|29|tonde capillum tuum et proice et sume in directum planctum quia proiecit Dominus et reliquit generationem furoris sui
JER|7|30|quia fecerunt filii Iuda malum in oculis meis dicit Dominus posuerunt offendicula sua in domo in qua invocatum est nomen meum ut polluerent eam
JER|7|31|et aedificaverunt excelsa Thofeth qui est in valle filii Ennom ut incenderent filios suos et filias suas igni quae non praecepi nec cogitavi in corde meo
JER|7|32|ideo ecce dies venient dicit Dominus et non dicetur amplius Thofeth et vallis filii Ennom sed vallis Interfectionis et sepelient in Thofeth eo quod non sit locus
JER|7|33|et erit morticinum populi huius in cibum volucribus caeli et bestiis terrae et non erit qui abigat
JER|7|34|et quiescere faciam de urbibus Iuda et de plateis Hierusalem vocem gaudii et vocem laetitiae vocem sponsi et vocem sponsae in desolatione enim erit terra
JER|8|1|in tempore illo ait Dominus eicient ossa regis Iuda et ossa principum eius et ossa sacerdotum et ossa prophetarum et ossa eorum qui habitaverunt Hierusalem de sepulchris suis
JER|8|2|et pandent ea ad solem et lunam et omnem militiam caeli quae dilexerunt et quibus servierunt et post quae ambulaverunt et quae quaesierunt et adoraverunt non colligentur et non sepelientur in sterquilinium super faciem terrae erunt
JER|8|3|et eligent magis mortem quam vitam omnes qui residui fuerint de cognatione hac pessima in universis locis quae derelicta sunt ad quae eieci eos dicit Dominus exercituum
JER|8|4|et dices ad eos haec dicit Dominus numquid qui cadet non resurget et qui aversus est non revertetur
JER|8|5|quare ergo aversus est populus iste in Hierusalem aversione contentiosa adprehenderunt mendacium et noluerunt reverti
JER|8|6|adtendi et auscultavi nemo quod bonum est loquitur nullus est qui agat paenitentiam super peccato suo dicens quid feci omnes conversi sunt ad cursum suum quasi equus impetu vadens in proelio
JER|8|7|milvus in caelo cognovit tempus suum turtur et hirundo et ciconia custodierunt tempus adventus sui populus autem meus non cognovit iudicium Domini
JER|8|8|quomodo dicitis sapientes nos sumus et lex Domini nobiscum est vere mendacium operatus est stilus mendax scribarum
JER|8|9|confusi sunt sapientes perterriti et capti sunt verbum enim Domini proiecerunt et sapientia nulla est in eis
JER|8|10|propterea dabo mulieres eorum exteris agros eorum heredibus quia a minimo usque ad maximum omnes avaritiam sequuntur a propheta usque ad sacerdotem cuncti faciunt mendacium
JER|8|11|et sanabant contritionem filiae populi mei ad ignominiam dicentes pax pax cum non esset pax
JER|8|12|confusi sunt quia abominationem fecerunt quinimmo confusione non sunt confusi et erubescere nescierunt idcirco cadent inter corruentes in tempore visitationis suae corruent dicit Dominus
JER|8|13|congregans congregabo eos ait Dominus non est uva in vitibus et non sunt ficus in ficulnea folium defluxit et dedi eis quae praetergressa sunt
JER|8|14|quare sedemus convenite et ingrediamur civitatem munitam et sileamus ibi quia Dominus noster silere nos fecit et potum dedit nobis aquam fellis peccavimus enim Domino
JER|8|15|expectavimus pacem et non erat bonum tempus medellae et ecce formido
JER|8|16|a Dan auditus est fremitus equorum eius a voce hinnituum pugnatorum eius commota est omnis terra et venerunt et devoraverunt terram et plenitudinem eius urbem et habitatores eius
JER|8|17|quia ecce ego mittam vobis serpentes regulos quibus non est incantatio et mordebunt vos ait Dominus
JER|8|18|dolor meus super dolorem in me cor meum maerens
JER|8|19|ecce vox clamoris filiae populi mei de terra longinqua numquid Dominus non est in Sion aut rex eius non est in ea quare ergo me ad iracundiam concitaverunt in sculptilibus suis et in vanitatibus alienis
JER|8|20|transiit messis finita est aestas et nos salvati non sumus
JER|8|21|super contritionem filiae populi mei contritus sum et contristatus stupor obtinuit me
JER|8|22|numquid resina non est in Galaad aut medicus non est ibi quare igitur non est obducta cicatrix filiae populi mei
JER|9|1|quis dabit capiti meo aquam et oculis meis fontem lacrimarum et plorabo die et nocte interfectos filiae populi mei
JER|9|2|quis dabit me in solitudine diversorium viatorum et derelinquam populum meum et recedam ab eis quia omnes adulteri sunt coetus praevaricatorum
JER|9|3|et extenderunt linguam suam quasi arcum mendacii et non veritatis confortati sunt in terra quia de malo ad malum egressi sunt et me non cognoverunt dicit Dominus
JER|9|4|unusquisque se a proximo suo custodiat et in omni fratre suo non habeat fiduciam quia omnis frater subplantans subplantabit et omnis amicus fraudulenter incedet
JER|9|5|et vir fratrem suum deridebit et veritatem non loquentur docuerunt enim linguam suam loqui mendacium ut inique agerent laboraverunt
JER|9|6|habitatio tua in medio doli in dolo rennuerunt scire me dicit Dominus
JER|9|7|propterea haec dicit Dominus exercituum ecce ego conflabo et probabo eos quid enim aliud faciam a facie filiae populi mei
JER|9|8|sagitta vulnerans lingua eorum dolum locuta est in ore suo pacem cum amico suo loquitur et occulte ponit ei insidias
JER|9|9|numquid super his non visitabo dicit Dominus aut in gentem huiuscemodi non ulciscetur anima mea
JER|9|10|super montes adsumam fletum ac lamentum et super speciosa deserti planctum quoniam incensa sunt eo quod non sit vir pertransiens et non audierunt vocem possidentis a volucre caeli usque ad pecora transmigraverunt et recesserunt
JER|9|11|et dabo Hierusalem in acervos harenae et cubilia draconum et civitates Iuda dabo in desolationem eo quod non sit habitator
JER|9|12|quis est vir sapiens qui intellegat hoc et ad quem verbum oris Domini fiat ut adnuntiet istud quare perierit terra exusta sit quasi desertum eo quod non sit qui pertranseat
JER|9|13|et dixit Dominus quia dereliquerunt legem meam quam dedi eis et non audierunt vocem meam et non ambulaverunt in ea
JER|9|14|et abierunt post pravitatem cordis sui et post Baalim quos didicerunt a patribus suis
JER|9|15|idcirco haec dicit Dominus exercituum Deus Israhel ecce ego cibabo eos populum istum absinthio et potum dabo eis aquam fellis
JER|9|16|et dispergam eos in gentibus quas non noverunt ipsi et patres eorum et mittam post eos gladium donec consumantur
JER|9|17|haec dicit Dominus exercituum contemplamini et vocate lamentatrices et veniant et ad eas quae sapientes sunt mittite et properent
JER|9|18|festinent et adsumant super nos lamentum deducant oculi nostri lacrimas et palpebrae nostrae defluant aquis
JER|9|19|quia vox lamentationis audita est de Sion quomodo vastati sumus et confusi vehementer quia dereliquimus terram quoniam deiecta sunt tabernacula nostra
JER|9|20|audite ergo mulieres verbum Domini et adsumat auris vestra sermonem oris eius et docete filias vestras lamentum et unaquaeque proximam suam planctum
JER|9|21|quia ascendit mors per fenestras nostras ingressa est domos nostras disperdere parvulos de foris iuvenes de plateis
JER|9|22|loquere haec dicit Dominus et cadet morticinum hominis quasi stercus super faciem regionis et quasi faenum post tergum metentis et non est qui colligat
JER|9|23|haec dicit Dominus non glorietur sapiens in sapientia sua et non glorietur fortis in fortitudine sua et non glorietur dives in divitiis suis
JER|9|24|sed in hoc glorietur qui gloriatur scire et nosse me quia ego sum Dominus qui facio misericordiam et iudicium et iustitiam in terra haec enim placent mihi ait Dominus
JER|9|25|ecce dies veniunt dicit Dominus et visitabo super omnem qui circumcisum habet praeputium
JER|9|26|super Aegyptum et super Iudam et super Edom et super filios Ammon et super Moab et super omnes qui adtonsi sunt in comam habitantes in deserto quia omnes gentes habent praeputium omnis autem domus Israhel incircumcisi sunt corde
JER|10|1|audite verbum quod locutus est Dominus super vos domus Israhel
JER|10|2|haec dicit Dominus iuxta vias gentium nolite discere et a signis caeli nolite metuere quae timent gentes
JER|10|3|quia leges populorum vanae sunt quia lignum de saltu praecidit opus manuum artificis in ascia
JER|10|4|argento et auro decoravit illud clavis et malleis conpegit ut non dissolvatur
JER|10|5|in similitudinem palmae fabricata sunt et non loquentur portata tollentur quia incedere non valent nolite ergo timere ea quia nec male possunt facere nec bene
JER|10|6|non est similis tui Domine magnus tu et magnum nomen tuum in fortitudine
JER|10|7|quis non timebit te o rex gentium tuum est enim decus inter cunctos sapientes gentium et in universis regnis eorum nullus est similis tui
JER|10|8|pariter insipientes et fatui probabuntur doctrina vanitatis eorum lignum est
JER|10|9|argentum involutum de Tharsis adfertur et aurum de Ofaz opus artificis et manus aerarii hyacinthus et purpura indumentum eorum opus artificum universa haec
JER|10|10|Dominus autem Deus verus est ipse Deus vivens et rex sempiternus ab indignatione eius commovebitur terra et non sustinebunt gentes comminationem eius
JER|10|11|sic ergo dicetis eis dii qui caelos et terram non fecerunt pereant de terra et de his quae sub caelis sunt
JER|10|12|qui facit terram in fortitudine sua praeparat orbem in sapientia sua et prudentia sua extendit caelos
JER|10|13|ad vocem suam dat multitudinem aquarum in caelo et elevat nebulas ab extremitatibus terrae fulgura in pluviam facit et educit ventum de thesauris suis
JER|10|14|stultus factus est omnis homo ab scientia confusus est omnis artifex in sculptili quoniam falsum est quod conflavit et non est spiritus in eis
JER|10|15|vana sunt et opus risu dignum in tempore visitationis suae peribunt
JER|10|16|non est his similis pars Iacob qui enim formavit omnia ipse est et Israhel virga hereditatis eius Dominus exercituum nomen illi
JER|10|17|congrega de terra confusionem tuam quae habitas in obsidione
JER|10|18|quia haec dicit Dominus ecce ego longe proiciam habitatores terrae in hac vice et tribulabo eos ita ut inveniantur
JER|10|19|vae mihi super contritione mea pessima plaga mea ego autem dixi plane haec infirmitas mea est et portabo illam
JER|10|20|tabernaculum meum vastatum est omnes funiculi mei disrupti sunt filii mei exierunt a me et non subsistunt non est qui extendat ultra tentorium meum et erigat pelles meas
JER|10|21|quia stulte egerunt pastores et Dominum non quaesierunt propterea non intellexerunt et omnis grex eorum dispersus est
JER|10|22|vox auditionis ecce venit et commotio magna de terra aquilonis ut ponat civitates Iuda solitudinem et habitaculum draconum
JER|10|23|scio Domine quia non est hominis via eius nec viri est ut ambulet et dirigat gressus suos
JER|10|24|corripe me Domine verumtamen in iudicio et non in furore tuo ne forte ad nihilum redigas me
JER|10|25|effunde indignationem tuam super gentes quae non cognoverunt te et super provincias quae nomen tuum non invocaverunt quia comederunt Iacob et devoraverunt eum et consumpserunt illum et decus eius dissipaverunt
JER|11|1|verbum quod factum est ad Hieremiam a Domino dicens
JER|11|2|audite verba pacti huius et loquimini ad viros Iuda et habitatores Hierusalem
JER|11|3|et dices ad eos haec dicit Dominus Deus Israhel maledictus vir qui non audierit verba pacti huius
JER|11|4|quod praecepi patribus vestris in die qua eduxi eos de terra Aegypti de fornace ferrea dicens audite vocem meam et facite omnia quae praecipio vobis et eritis mihi in populum et ego ero vobis in Deum
JER|11|5|ut suscitem iuramentum quod iuravi patribus vestris daturum me eis terram fluentem lacte et melle sicut est dies haec et respondi et dixi amen Domine
JER|11|6|et dixit Dominus ad me vociferare omnia verba haec in civitatibus Iuda et foris Hierusalem dicens audite verba pacti huius et facite illa
JER|11|7|quia contestans contestatus sum patres vestros in die qua eduxi eos de terra Aegypti usque ad diem hanc mane surgens contestatus sum et dixi audite vocem meam
JER|11|8|et non audierunt nec inclinaverunt aurem suam sed abierunt unusquisque in pravitate cordis sui mali et induxi super eos omnia verba pacti huius quod praecepi ut facerent et non fecerunt
JER|11|9|et dixit Dominus ad me inventa est coniuratio in viris Iuda et in habitatoribus Hierusalem
JER|11|10|reversi sunt ad iniquitates patrum suorum priores qui noluerunt audire verba mea et hii ergo abierunt post deos alienos ut servirent eis irritum fecerunt domus Israhel et domus Iuda pactum meum quod pepigi cum patribus eorum
JER|11|11|quam ob rem haec dicit Dominus ecce ego inducam super eos mala de quibus exire non poterunt et clamabunt ad me et non exaudiam eos
JER|11|12|et ibunt civitates Iuda et habitatores Hierusalem et clamabunt ad deos quibus libant et non salvabunt eos in tempore adflictionis eorum
JER|11|13|secundum numerum enim civitatum tuarum erant dii tui Iuda et secundum numerum viarum Hierusalem posuistis aras confusionis aras ad libandum Baali
JER|11|14|tu ergo noli orare pro populo hoc et ne adsumas pro eis laudem et orationem quia non exaudiam in tempore clamoris eorum ad me in tempore adflictionis eorum
JER|11|15|quid est quod dilectus meus in domo mea fecit scelera multa numquid carnes sanctae auferent a te malitias tuas in quibus gloriata es
JER|11|16|olivam uberem pulchram fructiferam speciosam vocavit Dominus nomen tuum ad vocem loquellae grandis exarsit ignis in ea et conbusta sunt frutecta eius
JER|11|17|et Dominus exercituum qui plantavit te locutus est super te malum pro malis domus Israhel et domus Iuda quae fecerunt sibi ad inritandum me libantes Baali
JER|11|18|tu autem Domine demonstrasti mihi et cognovi tunc ostendisti mihi studia eorum
JER|11|19|et ego quasi agnus mansuetus qui portatur ad victimam et non cognovi quia super me cogitaverunt consilia mittamus lignum in panem eius et eradamus eum de terra viventium et nomen eius non memoretur amplius
JER|11|20|tu autem Domine Sabaoth qui iudicas iuste et probas renes et cor videam ultionem tuam ex eis tibi enim revelavi causam meam
JER|11|21|propterea haec dicit Dominus ad viros Anathoth qui quaerunt animam tuam et dicunt non prophetabis in nomine Domini et non morieris in manibus nostris
JER|11|22|propterea haec dicit Dominus exercituum ecce ego visitabo super eos iuvenes morientur in gladio filii eorum et filiae eorum morientur in fame
JER|11|23|et reliquiae non erunt ex eis inducam enim malum super viros Anathoth annum visitationis eorum
JER|12|1|iustus quidem tu es Domine si disputem tecum verumtamen iusta loquar ad te quare via impiorum prosperatur bene est omnibus qui praevaricantur et inique agunt
JER|12|2|plantasti eos et radicem miserunt proficiunt et faciunt fructum prope es tu ori eorum et longe a renibus eorum
JER|12|3|et tu Domine nosti me vidisti me et probasti cor meum tecum congrega eos quasi gregem ad victimam et sanctifica eos in die occisionis
JER|12|4|usquequo lugebit terra et herba omnis regionis siccabitur propter malitiam habitantium in ea consumptum est animal et volucre quoniam dixerunt non videbit novissima nostra
JER|12|5|si cum peditibus currens laborasti quomodo contendere poteris cum equis cum autem in terra pacis secura fueris quid facies in superbia Iordanis
JER|12|6|nam et fratres tui et domus patris tui etiam ipsi pugnaverunt adversum te et clamaverunt post te plena voce ne credas eis cum locuti fuerint tibi bona
JER|12|7|reliqui domum meam dimisi hereditatem meam dedi dilectam animam meam in manu inimicorum eius
JER|12|8|facta est mihi hereditas mea quasi leo in silva dedit contra me vocem ideo odivi eam
JER|12|9|numquid avis discolor hereditas mea mihi numquid avis tincta per totum venite congregamini omnes bestiae terrae properate ad devorandum
JER|12|10|pastores multi demoliti sunt vineam meam conculcaverunt partem meam dederunt portionem meam desiderabilem in desertum solitudinis
JER|12|11|posuerunt eam in dissipationem luxitque super me desolatione desolata est omnis terra quia nullus est qui recogitet corde
JER|12|12|super omnes vias deserti venerunt vastatores quia gladius Domini devoravit ab extremo terrae usque ad extremum eius non est pax universae carni
JER|12|13|seminaverunt triticum et spinas messuerunt hereditatem acceperunt et non eis proderit confundemini a fructibus vestris propter iram furoris Domini
JER|12|14|haec dicit Dominus adversum omnes vicinos meos pessimos qui tangunt hereditatem quam distribui populo meo Israhel ecce ego evellam eos de terra eorum et domum Iuda evellam de medio eorum
JER|12|15|et cum evellero eos convertar et miserebor eorum et reducam eos virum ad hereditatem suam et virum in terram suam
JER|12|16|et erit si eruditi didicerint vias populi mei ut iurent in nomine meo vivit Dominus sicut docuerunt populum meum iurare in Baal aedificabuntur in medio populi mei
JER|12|17|quod si non audierint evellam gentem illam evulsione et perditione ait Dominus
JER|13|1|haec dicit Dominus ad me vade et posside tibi lumbare lineum et pones illud super lumbos tuos et in aquam non inferes illud
JER|13|2|et possedi lumbare iuxta verbum Domini et posui circa lumbos meos
JER|13|3|et factus est sermo Domini ad me secundo dicens
JER|13|4|tolle lumbare quod possedisti quod est circa lumbos tuos et surgens vade ad Eufraten et absconde illud ibi in foramine petrae
JER|13|5|et abii et abscondi illud in Eufraten sicut praeceperat mihi Dominus
JER|13|6|et factum est post dies plurimos dixit Dominus ad me surge vade ad Eufraten et tolle inde lumbare quod praecepi tibi ut absconderes illud ibi
JER|13|7|et abii ad Eufraten et fodi et tuli lumbare de loco ubi absconderam illud et ecce conputruerat lumbare ita ut nullo usui aptum esset
JER|13|8|et factum est verbum Domini ad me dicens
JER|13|9|haec dicit Dominus sic putrescere faciam superbiam Iuda et superbiam Hierusalem multam
JER|13|10|populum istum pessimum qui nolunt audire verba mea et ambulant in pravitate cordis sui abieruntque post deos alienos ut servirent eis et adorarent eos et erunt sicut lumbare istud quod nullo usui aptum est
JER|13|11|sicut enim adheret lumbare ad lumbos viri sic adglutinavi mihi omnem domum Israhel et omnem domum Iuda dicit Dominus ut esset mihi in populum et in nomen et in laudem et in gloriam et non audierunt
JER|13|12|dices ergo ad eos sermonem istum haec dicit Dominus Deus Israhel omnis laguncula implebitur vino et dicent ad te numquid ignoramus quia omnis laguncula implebitur vino
JER|13|13|et dices ad eos haec dicit Dominus ecce ego implebo omnes habitatores terrae huius et reges qui sedent de stirpe David super thronum eius et sacerdotes et prophetas et omnes habitatores Hierusalem ebrietate
JER|13|14|et dispergam eos virum a fratre suo et patres et filios pariter ait Dominus non parcam et non concedam neque miserebor ut non disperdam eos
JER|13|15|audite et auribus percipite nolite elevari quia Dominus locutus est
JER|13|16|date Domino Deo vestro gloriam antequam contenebrescat et antequam offendant pedes vestri ad montes caligosos expectabitis lucem et ponet eam in umbram mortis et in caliginem
JER|13|17|quod si hoc non audieritis in abscondito plorabit anima mea a facie superbiae plorans plorabit et deducet oculus meus lacrimam quia captus est grex Domini
JER|13|18|dic regi et dominatrici humiliamini sedete quoniam descendit de capite vestro corona gloriae vestrae
JER|13|19|civitates austri clausae sunt et non est qui aperiat translata est omnis Iudaea transmigratione perfecta
JER|13|20|levate oculos vestros et videte qui venitis ab aquilone ubi est grex qui datus est tibi pecus inclitum tuum
JER|13|21|quid dices cum visitaverit te tu enim docuisti eos adversum te et erudisti in caput tuum numquid non dolores adprehendent te quasi mulierem parturientem
JER|13|22|quod si dixeris in corde tuo quare venerunt mihi haec propter multitudinem iniquitatis tuae revelata sunt verecundiora tua pollutae sunt plantae tuae
JER|13|23|si mutare potest Aethiops pellem suam aut pardus varietates suas et vos poteritis bene facere cum didiceritis malum
JER|13|24|et disseminabo eos quasi stipulam quae vento raptatur in deserto
JER|13|25|haec sors tua parsque mensurae tuae a me dicit Dominus quia oblita es mei et confisa es in mendacio
JER|13|26|unde et ego nudavi femora tua contra faciem tuam et apparuit ignominia tua
JER|13|27|adulteria tua et hinnitus tuus scelus fornicationis tuae super colles in agro vidi abominationes tuas vae tibi Hierusalem non mundaberis post me usquequo adhuc
JER|14|1|quod factum est verbum Domini ad Hieremiam de sermonibus siccitatis
JER|14|2|luxit Iudaea et portae eius corruerunt et obscuratae sunt in terra et clamor Hierusalem ascendit
JER|14|3|maiores miserunt minores suos ad aquam venerunt ad hauriendum non invenerunt aquam reportaverunt vasa sua vacua confusi sunt et adflicti et operuerunt capita sua
JER|14|4|propter terrae vastitatem quia non venit pluvia in terra confusi sunt agricolae operuerunt capita sua
JER|14|5|nam et cerva in agro peperit et reliquit quia non erat herba
JER|14|6|et onagri steterunt in rupibus traxerunt ventum quasi dracones defecerunt oculi eorum quia non erat herba
JER|14|7|si iniquitates nostrae responderunt nobis Domine fac propter nomen tuum quoniam multae sunt aversiones nostrae tibi peccavimus
JER|14|8|expectatio Israhel salvator eius in tempore tribulationis quare quasi colonus futurus es in terra et quasi viator declinans ad manendum
JER|14|9|quare futurus es velut vir vagus ut fortis qui non potest salvare tu autem in nobis es Domine et nomen tuum super nos invocatum est ne derelinquas nos
JER|14|10|haec dicit Dominus populo huic qui dilexit movere pedes suos et non quievit et Domino non placuit nunc recordabitur iniquitatum eorum et visitabit peccata eorum
JER|14|11|et dixit Dominus ad me noli orare pro populo isto in bonum
JER|14|12|cum ieiunaverint non exaudiam preces eorum et si obtulerint holocaustomata et victimas non suscipiam ea quoniam gladio et fame et peste ego consumam eos
JER|14|13|et dixi a a a Domine Deus prophetae dicunt eis non videbitis gladium et famis non erit in vobis sed pacem veram dabit vobis in loco isto
JER|14|14|et dixit Dominus ad me falso prophetae vaticinantur in nomine meo non misi eos et non praecepi eis neque locutus sum ad eos visionem mendacem et divinationem et fraudulentiam et seductionem cordis sui prophetant vobis
JER|14|15|ideo haec dicit Dominus de prophetis qui prophetant in nomine meo quos ego non misi dicentes gladius et famis non erit in terra hac in gladio et fame consumentur prophetae illi
JER|14|16|et populi quibus prophetant erunt proiecti in viis Hierusalem prae fame et gladio et non erit qui sepeliat eos ipsi et uxores eorum filii et filiae eorum et effundam super eos malum suum
JER|14|17|et dices ad eos verbum istud deducant oculi mei lacrimam per noctem et diem et non taceant quoniam contritione magna contrita est virgo filia populi mei plaga pessima vehementer
JER|14|18|si egressus fuero ad agros ecce occisi gladio et si introiero in civitatem ecce adtenuati fame propheta quoque et sacerdos abierunt in terram quam ignorabant
JER|14|19|numquid proiciens abiecisti Iudam aut Sion abominata est anima tua quare ergo percussisti nos ita ut nulla sit sanitas expectavimus pacem et non est bonum et tempus curationis et ecce turbatio
JER|14|20|cognovimus Domine impietates nostras iniquitatem patrum nostrorum quia peccavimus tibi
JER|14|21|ne nos des in obprobrium propter nomen tuum neque facias nobis contumeliam solii gloriae tuae recordare ne irritum facias foedus tuum nobiscum
JER|14|22|numquid sunt in sculptilibus gentium qui pluant aut caeli possunt dare imbres nonne tu es Domine Deus noster quem expectavimus tu enim fecisti omnia haec
JER|15|1|et dixit Dominus ad me si steterit Moses et Samuhel coram me non est anima mea ad populum istum eice illos a facie mea et egrediantur
JER|15|2|quod si dixerint ad te quo egrediemur dices ad eos haec dicit Dominus qui ad mortem ad mortem et qui ad gladium ad gladium et qui ad famem ad famem et qui ad captivitatem ad captivitatem
JER|15|3|et visitabo super eos quattuor species dicit Dominus gladium ad occisionem et canes ad lacerandum et volatilia caeli et bestias terrae ad devorandum et dissipandum
JER|15|4|et dabo eos in fervorem universis regnis terrae propter Manassem filium Ezechiae regis Iuda super omnibus quae fecit in Hierusalem
JER|15|5|quis enim miserebitur tui Hierusalem aut quis contristabitur pro te aut quis ibit ad rogandum pro pace tua
JER|15|6|tu reliquisti me dicit Dominus retrorsum abisti et extendam manum meam super te et interficiam te laboravi rogans
JER|15|7|et dispergam eos ventilabro in portis terrae interfeci et perdidi populum meum et tamen a viis suis non sunt reversi
JER|15|8|multiplicatae sunt mihi viduae eius super harenam maris induxi eis super matrem adulescentis vastatorem meridie misi super civitates repente terrorem
JER|15|9|infirmata est quae peperit septem defecit anima eius occidit ei sol cum adhuc esset dies confusa est et erubuit et residuos eius in gladium dabo in conspectu inimicorum eorum ait Dominus
JER|15|10|vae mihi mater mea quare genuisti me virum rixae virum discordiae in universa terra non feneravi nec feneravit mihi quisquam omnes maledicunt mihi
JER|15|11|dicit Dominus si non reliquiae tuae in bonum si non occurri tibi in tempore adflictionis et in tempore tribulationis adversum inimicum
JER|15|12|numquid foederabitur ferrum ferro ab aquilone et aes
JER|15|13|divitias tuas et thesauros tuos in direptionem dabo gratis in omnibus peccatis tuis et in omnibus terminis tuis
JER|15|14|et adducam inimicos tuos de terra qua nescis quia ignis succensus est in furore meo super vos ardebit
JER|15|15|tu scis Domine recordare mei et visita me et tuere me ab his qui persequuntur me noli in patientia tua suscipere me scito quoniam sustinui pro te obprobrium
JER|15|16|inventi sunt sermones tui et comedi eos et factum est mihi verbum tuum in gaudium et in laetitiam cordis mei quoniam invocatum est nomen tuum super me Domine Deus exercituum
JER|15|17|non sedi in concilio ludentium et gloriatus sum a facie manus tuae solus sedebam quoniam comminatione replesti me
JER|15|18|quare factus est dolor meus perpetuus et plaga mea desperabilis rennuit curari facta est mihi quasi mendacium aquarum infidelium
JER|15|19|propter hoc haec dicit Dominus si converteris convertam te et ante faciem meam stabis et si separaveris pretiosum a vili quasi os meum eris convertentur ipsi ad te et tu non converteris ad eos
JER|15|20|et dabo te populo huic in murum aereum fortem et bellabunt adversum te et non praevalebunt quia ego tecum sum ut salvem te et eruam dicit Dominus
JER|15|21|et liberabo te de manu pessimorum et redimam te de manu fortium
JER|16|1|et factum est verbum Domini ad me dicens
JER|16|2|non accipies uxorem et non erunt tibi filii et filiae in loco isto
JER|16|3|quia haec dicit Dominus super filios et filias qui generantur in loco isto et super matres eorum quae genuerunt eos et super patres eorum de quorum stirpe sunt nati in terra hac
JER|16|4|mortibus aegrotationum morientur non plangentur et non sepelientur in sterquilinium super faciem terrae erunt et gladio et fame consumentur et erit cadaver eorum in escam volatilibus caeli et bestiis terrae
JER|16|5|haec enim dicit Dominus ne ingrediaris domum convivii neque vadas ad plangendum neque consoleris eos quia abstuli pacem meam a populo isto dicit Dominus misericordiam et miserationes
JER|16|6|et morientur grandes et parvi in terra ista non sepelientur neque plangentur et non se incident neque calvitium fiet pro eis
JER|16|7|et non frangent inter eos lugenti panem ad consolandum super mortuo et non dabunt eis potum calicis ad consolandum super patre suo et matre
JER|16|8|et domum convivii non ingredieris ut sedeas cum eis et comedas et bibas
JER|16|9|quia haec dicit Dominus exercituum Deus Israhel ecce ego auferam de loco isto in oculis vestris et in diebus vestris vocem gaudii et vocem laetitiae vocem sponsi et vocem sponsae
JER|16|10|et cum adnuntiaveris populo huic omnia verba haec et dixerint tibi quare locutus est Dominus super nos omne malum grande istud quae iniquitas nostra et quod peccatum nostrum quod peccavimus Domino Deo nostro
JER|16|11|dices ad eos quia dereliquerunt patres vestri me ait Dominus et abierunt post deos alienos et servierunt eis et adoraverunt eos et me dereliquerunt et legem meam non custodierunt
JER|16|12|sed et vos peius operati estis quam patres vestri ecce enim ambulat unusquisque post pravitatem cordis sui mali ut me non audiat
JER|16|13|et eiciam vos de terra hac in terram quam ignoratis vos et patres vestri et servietis ibi diis alienis die ac nocte qui non dabunt vobis requiem
JER|16|14|propterea ecce dies veniunt dicit Dominus et non dicetur ultra vivit Dominus qui eduxit filios Israhel de terra Aegypti
JER|16|15|sed vivit Dominus qui eduxit filios Israhel de terra aquilonis et de universis terris ad quas eieci eos et reducam eos in terram suam quam dedi patribus eorum
JER|16|16|ecce ego mittam piscatores multos dicit Dominus et piscabuntur eos et post haec mittam eis multos venatores et venabuntur eos de omni monte et de omni colle et de cavernis petrarum
JER|16|17|quia oculi mei super omnes vias eorum non sunt absconditae a facie mea et non fuit occulta iniquitas eorum ab oculis meis
JER|16|18|et reddam primum duplices iniquitates et peccata eorum quia contaminaverunt terram meam in morticinis idolorum suorum et abominationibus suis impleverunt hereditatem meam
JER|16|19|Domine fortitudo mea et robur meum et refugium meum in die tribulationis ad te gentes venient ab extremis terrae et dicent vere mendacium possederunt patres nostri vanitatem quae eis non profuit
JER|16|20|numquid faciet sibi homo deos et ipsi non sunt dii
JER|16|21|idcirco ecce ego ostendam eis per vicem hanc ostendam eis manum meam et virtutem meam et scient quia nomen mihi Dominus
JER|17|1|peccatum Iuda scriptum est stilo ferreo in ungue adamantino exaratum super latitudinem cordis eorum et in cornibus ararum eorum
JER|17|2|cum recordati fuerint filii eorum ararum suarum et lucorum lignorumque frondentium in montibus excelsis
JER|17|3|sacrificantes in agro fortitudinem tuam et omnes thesauros tuos in direptionem dabo excelsa tua propter peccata in universis finibus tuis
JER|17|4|et relinqueris sola ab hereditate tua quam dedi tibi et servire te faciam inimicis tuis in terra quam ignoras quoniam ignem succendisti in furore meo usque in aeternum ardebit
JER|17|5|haec dicit Dominus maledictus homo qui confidit in homine et ponit carnem brachium suum et a Domino recedit cor eius
JER|17|6|erit enim quasi myrice in deserto et non videbit cum venerit bonum sed habitabit in siccitate in deserto in terra salsuginis et inhabitabili
JER|17|7|benedictus vir qui confidit in Domino et erit Dominus fiducia eius
JER|17|8|et erit quasi lignum quod transplantatur super aquas quod ad humorem mittit radices suas et non timebit cum venerit aestus et erit folium eius viride et in tempore siccitatis non erit sollicitum nec aliquando desinet facere fructum
JER|17|9|pravum est cor omnium et inscrutabile quis cognoscet illud
JER|17|10|ego Dominus scrutans cor et probans renes qui do unicuique iuxta viam et iuxta fructum adinventionum suarum
JER|17|11|perdix fovit quae non peperit fecit divitias et non in iudicio in dimidio dierum suorum derelinquet eas et in novissimo suo erit insipiens
JER|17|12|solium gloriae altitudinis a principio locus sanctificationis nostrae
JER|17|13|expectatio Israhel Domine omnes qui te derelinquunt confundentur recedentes in terra scribentur quoniam dereliquerunt venam aquarum viventium Dominum
JER|17|14|sana me Domine et sanabor salvum me fac et salvus ero quoniam laus mea tu es
JER|17|15|ecce ipsi dicunt ad me ubi est verbum Domini veniat
JER|17|16|et ego non sum turbatus te pastorem sequens et diem hominis non desideravi tu scis quod egressum est de labiis meis rectum in conspectu tuo fuit
JER|17|17|non sis mihi tu formidini spes mea tu in die adflictionis
JER|17|18|confundantur qui persequuntur me et non confundar ego paveant illi et non paveam ego induc super eos diem adflictionis et duplici contritione contere eos
JER|17|19|haec dicit Dominus ad me vade et sta in porta filiorum populi per quam ingrediuntur reges Iuda et egrediuntur et in cunctis portis Hierusalem
JER|17|20|et dices ad eos audite verbum Domini reges Iuda et omnis Iudaea cunctique habitatores Hierusalem qui ingredimini per portas istas
JER|17|21|haec dicit Dominus custodite animas vestras et nolite portare pondera in die sabbati nec inferatis per portas Hierusalem
JER|17|22|et nolite eicere onera de domibus vestris in die sabbati et omne opus non facietis sanctificate diem sabbati sicut praecepi patribus vestris
JER|17|23|et non audierunt nec inclinaverunt aurem suam sed induraverunt cervicem suam ne audirent me et ne acciperent disciplinam
JER|17|24|et erit si audieritis me dicit Dominus ut non inferatis onera per portas civitatis huius in die sabbati et si sanctificaveritis diem sabbati ne faciatis in ea omne opus
JER|17|25|ingredientur per portas civitatis huius reges et principes sedentes super solium David et ascendentes in curribus et equis ipsi et principes eorum vir Iuda et habitatores Hierusalem et habitabitur civitas haec in sempiternum
JER|17|26|et venient de civitate Iuda et de circuitu Hierusalem et de terra Beniamin et de campestribus et de montuosis et ab austro portantes holocaustum et victimam et sacrificium et tus et inferent oblationem in domum Domini
JER|17|27|si autem non audieritis me ut sanctificetis diem sabbati et ne portetis onus et ne inferatis per portas Hierusalem in die sabbati succendam ignem in portis eius et devorabit domos Hierusalem et non extinguetur
JER|18|1|verbum quod factum est ad Hieremiam a Domino dicens
JER|18|2|surge et descende in domum figuli et ibi audies verba mea
JER|18|3|et descendi in domum figuli et ecce ipse faciebat opus super rotam
JER|18|4|et dissipatum est vas quod ipse faciebat e luto manibus suis conversusque fecit illud vas alterum sicut placuerat in oculis eius ut faceret
JER|18|5|et factum est verbum Domini ad me dicens
JER|18|6|numquid sicut figulus iste non potero facere vobis domus Israhel ait Dominus ecce sicut lutum in manu figuli sic vos in manu mea domus Israhel
JER|18|7|repente loquar adversum gentem et adversum regnum ut eradicem et destruam et disperdam illud
JER|18|8|si paenitentiam egerit gens illa a malo suo quod locutus sum adversum eam agam et ego paenitentiam super malo quod cogitavi ut facerem ei
JER|18|9|et subito loquar de gente et regno ut aedificem et ut plantem illud
JER|18|10|si fecerit malum in oculis meis ut non audiat vocem meam paenitentiam agam super bono quod locutus sum ut facerem ei
JER|18|11|nunc ergo dic viro Iudae et habitatoribus Hierusalem dicens haec dicit Dominus ecce ego fingo contra vos malum et cogito contra vos cogitationem revertatur unusquisque a via sua mala et dirigite vias vestras et studia vestra
JER|18|12|qui dixerunt desperavimus post cogitationes enim nostras ibimus et unusquisque pravitatem cordis sui mali faciemus
JER|18|13|ideo haec dicit Dominus interrogate gentes quis audivit talia horribilia quae fecit nimis virgo Israhel
JER|18|14|numquid deficiet de petra agri nix Libani aut evelli possunt aquae erumpentes frigidae et defluentes
JER|18|15|quia oblitus est mei populus meus frustra libantes et inpingentes in viis suis in semitis saeculi ut ambularent per eas in itinere non trito
JER|18|16|ut fieret terra eorum in desolationem et in sibilum sempiternum omnis qui praeterit per eam obstupescet et movebit caput suum
JER|18|17|sicut ventus urens dispergam eos coram inimico dorsum et non faciem ostendam eis in die perditionis eorum
JER|18|18|et dixerunt venite et cogitemus contra Hieremiam cogitationes non enim peribit lex a sacerdote neque consilium a sapiente nec sermo a propheta venite et percutiamus eum lingua et non adtendamus ad universos sermones eius
JER|18|19|adtende Domine ad me et audi vocem adversariorum meorum
JER|18|20|numquid redditur pro bono malum quia foderunt foveam animae meae recordare quod steterim in conspectu tuo ut loquerer pro eis bonum et averterem indignationem tuam ab eis
JER|18|21|propterea da filios eorum in famem et deduc eos in manus gladii fiant uxores eorum absque liberis et viduae et viri earum interficiantur morte iuvenes eorum confodiantur gladio in proelio
JER|18|22|audiatur clamor de domibus eorum adduces enim super eos latronem repente quia foderunt foveam ut caperent me et laqueos absconderunt pedibus meis
JER|18|23|tu autem Domine scis omne consilium eorum adversum me in mortem ne propitieris iniquitati eorum et peccatum eorum a facie tua non deleatur fiant corruentes in conspectu tuo in tempore furoris tui abutere eis
JER|19|1|haec dicit Dominus vade et accipe lagunculam figuli testeam a senioribus populi et a senioribus sacerdotum
JER|19|2|et egredere ad vallem filii Ennom quae est iuxta introitum portae Fictilis et praedicabis ibi verba quae ego loquar ad te
JER|19|3|et dices audite verbum Domini reges Iuda et habitatores Hierusalem haec dicit Dominus exercituum Deus Israhel ecce ego inducam adflictionem super locum istum ita ut omnis qui audierit illam tinniant aures eius
JER|19|4|eo quod dereliquerint me et alienum fecerint locum istum et libaverint in eo diis alienis quos nescierunt ipsi et patres eorum et reges Iuda et repleverunt locum istum sanguine innocentium
JER|19|5|et aedificaverunt excelsa Baali ad conburendos filios suos igni in holocaustum Baali quae non praecepi nec locutus sum nec ascenderunt in cor meum
JER|19|6|propterea ecce dies veniunt dicit Dominus et non vocabitur locus iste amplius Thofeth et vallis filii Ennom sed vallis Occisionis
JER|19|7|et dissipabo consilium Iudae et Hierusalem in loco isto et subvertam eos gladio in conspectu inimicorum suorum et in manu quaerentium animas eorum et dabo cadavera eorum escam volatilibus caeli et bestiis terrae
JER|19|8|et ponam civitatem hanc in stuporem et in sibilum omnis qui praeterierit per eam obstupescet et sibilabit super universa plaga eius
JER|19|9|et cibabo eos carnibus filiorum suorum et carnibus filiarum suarum et unusquisque carnes amici sui comedet in obsidione et in angustia in qua concludent eos inimici eorum et qui quaerunt animas eorum
JER|19|10|et conteres lagunculam in oculis virorum qui ibunt tecum
JER|19|11|et dices ad eos haec dicit Dominus exercituum sic conteram populum istum et civitatem istam sicut conteritur vas figuli quod non potest ultra instaurari et in Thofeth sepelientur eo quod non sit alius locus ad sepeliendum
JER|19|12|sic faciam loco huic ait Dominus et habitatoribus eius ut ponam civitatem istam sicut Thofeth
JER|19|13|et erunt domus Hierusalem et domus regum Iuda sicut locus Thofeth inmundae omnes domus in quarum domatibus sacrificaverunt omni militiae caeli et libaverunt libamina diis alienis
JER|19|14|venit autem Hieremias de Thofeth quo miserat eum Dominus ad prophetandum et stetit in atrio domus Domini et dixit ad omnem populum
JER|19|15|haec dicit Dominus exercituum Deus Israhel ecce ego inducam super civitatem hanc et super omnes urbes eius universa mala quae locutus sum adversum eam quoniam induraverunt cervicem suam ut non audirent sermones meos
JER|20|1|et audivit Phassur filius Emmer sacerdos qui constitutus erat princeps in domo Domini Hieremiam prophetantem sermones istos
JER|20|2|et percussit Phassur Hieremiam prophetam et misit eum in nervum quod erat in porta Beniamin superiori in domo Domini
JER|20|3|cumque inluxisset in crastinum eduxit Phassur Hieremiam de nervo et dixit ad eum Hieremias non Phassur vocavit Dominus nomen tuum sed Pavorem undique
JER|20|4|quia haec dicit Dominus ecce ego dabo te in pavorem te et omnes amicos tuos et corruent gladio inimicorum suorum et oculi tui videbunt et omnem Iudam dabo in manu regis Babylonis et traducet eos in Babylonem et percutiet eos gladio
JER|20|5|et dabo universam substantiam civitatis huius et omnem laborem eius omneque pretium et cunctos thesauros regum Iuda dabo in manu inimicorum eorum et diripient eos et tollent et ducent in Babylonem
JER|20|6|tu autem Phassur et omnes habitatores domus tuae ibitis in captivitatem et in Babylonem venies et ibi morieris ibique sepelieris tu et omnes amici tui quibus prophetasti mendacium
JER|20|7|seduxisti me Domine et seductus sum fortior me fuisti et invaluisti factus sum in derisum tota die omnes subsannant me
JER|20|8|quia iam olim loquor vociferans iniquitatem et vastitatem clamito et factus est mihi sermo Domini in obprobrium et in derisum tota die
JER|20|9|et dixi non recordabor eius neque loquar ultra in nomine illius et factus est in corde meo quasi ignis exaestuans claususque in ossibus meis et defeci ferre non sustinens
JER|20|10|audivi enim contumelias multorum et terrorem in circuitu persequimini et persequamur eum ab omnibus viris qui erant pacifici mei et custodientes latus meum si quo modo decipiatur et praevaleamus adversus eum et consequamur ultionem ex eo
JER|20|11|Dominus autem mecum est quasi bellator fortis idcirco qui persequuntur me cadent et infirmi erunt confundentur vehementer quia non intellexerunt obprobrium sempiternum quod numquam delebitur
JER|20|12|et tu Domine exercituum probator iusti qui vides renes et cor videam quaeso ultionem tuam ex eis tibi enim revelavi causam meam
JER|20|13|cantate Domino laudate Dominum quia liberavit animam pauperis de manu malorum
JER|20|14|maledicta dies in qua natus sum dies in qua peperit me mater mea non sit benedicta
JER|20|15|maledictus vir qui adnuntiavit patri meo dicens natus est tibi puer masculus et quasi gaudio laetificavit eum
JER|20|16|sit homo ille ut sunt civitates quas subvertit Dominus et non paenituit eum audiat clamorem mane et ululatum in tempore meridiano
JER|20|17|qui non me interfecit a vulva ut fieret mihi mater mea sepulchrum et vulva eius conceptus aeternus
JER|20|18|quare de vulva egressus sum ut viderem laborem et dolorem et consumerentur in confusione dies mei
JER|21|1|verbum quod factum est ad Hieremiam a Domino quando misit ad eum rex Sedecias Phassur filium Melchiae et Sophoniam filium Maasiae sacerdotem dicens
JER|21|2|interroga pro nobis Dominum quia Nabuchodonosor rex Babylonis proeliatur adversum nos si forte faciat Dominus nobiscum secundum omnia mirabilia sua et recedat a nobis
JER|21|3|et dixit Hieremias ad eos sic dicetis Sedeciae
JER|21|4|haec dicit Dominus Deus Israhel ecce ego convertam vasa belli quae in manibus vestris sunt et quibus vos pugnatis adversum regem Babylonis et Chaldeos qui obsident vos in circuitu murorum et congregabo ea in medio civitatis huius
JER|21|5|et debellabo ego vos in manu extenta et brachio forti et in furore et in indignatione et in ira grandi
JER|21|6|et percutiam habitatores civitatis huius homines et bestiae pestilentia magna morientur
JER|21|7|et post haec ait Dominus dabo Sedeciam regem Iuda et servos eius et populum eius et qui derelicti sunt in civitate hac a peste et gladio et fame in manu Nabuchodonosor regis Babylonis et in manu inimicorum eorum et in manu quaerentium animam eorum et percutiet eos in ore gladii et non movebitur neque parcet nec miserebitur
JER|21|8|et ad populum hunc dices haec dicit Dominus ecce ego do coram vobis viam vitae et viam mortis
JER|21|9|qui habitaverit in urbe hac morietur gladio et fame et peste qui autem egressus fuerit et transfugerit ad Chaldeos qui obsident vos vivet et erit ei anima sua quasi spolium
JER|21|10|posui enim faciem meam super civitatem hanc in malum et non in bonum ait Dominus in manu regis Babylonis dabitur et exuret eam igni
JER|21|11|et domui regis Iuda audite verbum Domini
JER|21|12|domus David haec dicit Dominus iudicate mane iudicium et eruite vi oppressum de manu calumniantis ne forte egrediatur ut ignis indignatio mea et succendatur et non sit qui extinguat propter malitiam studiorum vestrorum
JER|21|13|ecce ego ad te habitatricem vallis solidae atque campestris ait Dominus qui dicitis quis percutiet nos et quis ingredietur domos nostras
JER|21|14|et visitabo super vos iuxta fructum studiorum vestrorum dicit Dominus et succendam ignem in saltu eius et devorabit omnia in circuitu eius
JER|22|1|haec dicit Dominus descende in domum regis Iuda et loqueris ibi verbum hoc
JER|22|2|et dices audi verbum Domini rex Iuda qui sedes super solium David tu et servi tui et populus tuus qui ingredimini per portas istas
JER|22|3|haec dicit Dominus facite iudicium et iustitiam et liberate vi oppressum de manu calumniatoris et advenam et pupillum et viduam nolite contristare neque opprimatis inique et sanguinem innocentem ne effundatis in loco isto
JER|22|4|si enim facientes feceritis verbum istud ingredientur per portas domus huius reges sedentes de genere David super thronum eius et ascendentes currus et equos ipsi et servi et populus eorum
JER|22|5|quod si non audieritis verba haec in memet ipso iuravi dicit Dominus quia in solitudinem erit domus haec
JER|22|6|quia haec dicit Dominus super domum regis Iuda Galaad tu mihi caput Libani si non posuero te solitudinem urbes inhabitabiles
JER|22|7|et sanctificabo super te interficientem virum et arma eius et succident electam cedrum tuam et praecipitabunt in ignem
JER|22|8|et pertransibunt gentes multae per civitatem hanc et dicet unusquisque proximo suo quare fecit Dominus sic civitati huic grandi
JER|22|9|et respondebunt eo quod dereliquerint pactum Domini Dei sui et adoraverint deos alienos et servierint eis
JER|22|10|nolite flere mortuum neque lugeatis super eum fletu plangite eum qui egreditur quia non revertetur ultra nec videbit terram nativitatis suae
JER|22|11|quia haec dicit Dominus ad Sellum filium Iosiae regem Iuda qui regnavit pro Iosia patre suo qui egressus est de loco isto non revertetur huc amplius
JER|22|12|sed in loco ad quem transtuli eum ibi morietur et terram istam non videbit amplius
JER|22|13|vae qui aedificat domum suam in iniustitia et cenacula sua non in iudicio amicum suum opprimet frustra et mercedem eius non reddet ei
JER|22|14|qui dicit aedificabo mihi domum latam et cenacula spatiosa qui aperit sibi fenestras et facit laquearia cedrina pingitque sinopide
JER|22|15|numquid regnabis quoniam confers te cedro pater tuus numquid non comedit et bibit et fecit iudicium et iustitiam tunc cum bene erat ei
JER|22|16|iudicavit causam pauperis et egeni in bonum suum numquid non ideo quia cognovit me dicit Dominus
JER|22|17|tui vero oculi et cor ad avaritiam et ad sanguinem innocentem fundendum et ad calumniam et ad cursum mali operis
JER|22|18|propterea haec dicit Dominus ad Ioachim filium Iosiae regem Iuda non plangent eum vae frater et vae fratres non concrepabunt ei vae domine et vae inclite
JER|22|19|sepultura asini sepelietur putrefactus et proiectus extra portas Hierusalem
JER|22|20|ascende Libanum et clama et in Basan da vocem tuam et clama ad transeuntes quia contriti sunt omnes amatores tui
JER|22|21|locutus sum ad te in abundantia tua dixisti non audiam haec est via tua ab adulescentia tua quia non audisti vocem meam
JER|22|22|omnes pastores tuos pascet ventus et amatores tui in captivitatem ibunt et tunc confunderis et erubesces ab omni malitia tua
JER|22|23|quae sedes in Libano et nidificas in cedris quomodo congemuisti cum venissent tibi dolores quasi dolores parturientis
JER|22|24|vivo ego dicit Dominus quia si fuerit Iechonias filius Ioachim regis Iuda anulus in manu dextera mea inde avellam eum
JER|22|25|et dabo te in manu quaerentium animam tuam et in manu quorum tu formidas faciem et in manu Nabuchodonosor regis Babylonis et in manu Chaldeorum
JER|22|26|et mittam te et matrem tuam quae genuit te in terram alienam in qua nati non estis ibique moriemini
JER|22|27|et in terram ad quam ipsi levant animam suam ut revertantur illuc non revertentur
JER|22|28|numquid vas fictile atque contritum vir iste Iechonias numquid vas absque omni voluptate quare abiecti sunt ipse et semen eius et proiecti in terram quam ignoraverunt
JER|22|29|terra terra terra audi sermonem Domini
JER|22|30|haec dicit Dominus scribe virum istum sterilem virum qui in diebus suis non prosperabitur nec enim erit de semine eius vir qui sedeat super solium David et potestatem habeat ultra in Iuda
JER|23|1|vae pastoribus qui disperdunt et dilacerant gregem pascuae meae dicit Dominus
JER|23|2|ideo haec dicit Dominus Deus Israhel ad pastores qui pascunt populum meum vos dispersistis gregem meum eiecistis eos et non visitastis eos ecce ego visitabo super vos malitiam studiorum vestrorum ait Dominus
JER|23|3|et ego congregabo reliquias gregis mei de omnibus terris ad quas eiecero eos illuc et convertam eos ad rura sua et crescent et multiplicabuntur
JER|23|4|et suscitabo super eos pastores et pascent eos non formidabunt ultra et non pavebunt et nullus quaeretur ex numero dicit Dominus
JER|23|5|ecce dies veniunt ait Dominus et suscitabo David germen iustum et regnabit rex et sapiens erit et faciet iudicium et iustitiam in terra
JER|23|6|in diebus illius salvabitur Iuda et Israhel habitabit confidenter et hoc est nomen quod vocabunt eum Dominus iustus noster
JER|23|7|propter hoc ecce dies veniunt dicit Dominus et non dicent ultra vivit Dominus qui eduxit filios Israhel de terra Aegypti
JER|23|8|sed vivit Dominus qui eduxit et adduxit semen domus Israhel de terra aquilonis et de cunctis terris ad quas eieceram eos illuc et habitabunt in terra sua
JER|23|9|ad prophetas contritum est cor meum in medio mei contremuerunt omnia ossa mea factus sum quasi vir ebrius et quasi homo madidus a vino a facie Domini et a facie verborum sanctorum eius
JER|23|10|quia adulteris repleta est terra quia a facie maledictionis luxit terra arefacta sunt arva deserti factus est cursus eorum malus et fortitudo eorum dissimilis
JER|23|11|propheta namque et sacerdos polluti sunt et in domo mea inveni malum eorum ait Dominus
JER|23|12|idcirco via eorum erit quasi lubricum in tenebris inpellentur enim et corruent in ea adferam enim super eos mala annum visitationis eorum ait Dominus
JER|23|13|et in prophetis Samariae vidi fatuitatem prophetabant in Baal et decipiebant populum meum Israhel
JER|23|14|et in prophetis Hierusalem vidi similitudinem adulterium et iter mendacii et confortaverunt manus pessimorum ut non converteretur unusquisque a malitia sua facti sunt mihi omnes Sodoma et habitatores eius quasi Gomorra
JER|23|15|propterea haec dicit Dominus exercituum ad prophetas ecce ego cibabo eos absinthio et potabo eos felle a prophetis enim Hierusalem est egressa pollutio super omnem terram
JER|23|16|haec dicit Dominus exercituum nolite audire verba prophetarum qui prophetant vobis et decipiunt vos visionem cordis sui loquuntur non de ore Domini
JER|23|17|dicunt his qui blasphemant me locutus est Dominus pax erit vobis et omni qui ambulat in pravitate cordis sui dixerunt non veniet super vos malum
JER|23|18|quis enim adfuit in consilio Domini et vidit et audivit sermonem eius quis consideravit verbum illius et audivit
JER|23|19|ecce turbo dominicae indignationis egredietur et tempestas erumpens super caput impiorum veniet
JER|23|20|non revertetur furor Domini usque dum faciat et usque dum conpleat cogitationem cordis sui in novissimis diebus intellegetis consilium eius
JER|23|21|non mittebam prophetas et ipsi currebant non loquebar ad eos et ipsi prophetabant
JER|23|22|si stetissent in consilio meo et nota fecissent verba mea populo meo avertissem utique eos a via sua mala et a pessimis cogitationibus suis
JER|23|23|putasne Deus e vicino ego sum dicit Dominus et non Deus de longe
JER|23|24|si occultabitur vir in absconditis et ego non videbo eum dicit Dominus numquid non caelum et terram ego impleo ait Dominus
JER|23|25|audivi quae dixerunt prophetae prophetantes in nomine meo mendacium atque dicentes somniavi somniavi
JER|23|26|usquequo istud in corde est prophetarum vaticinantium mendacium et prophetantium seductiones cordis sui
JER|23|27|qui volunt facere ut obliviscatur populus meus nominis mei propter somnia eorum quae narrant unusquisque ad proximum suum sicut obliti sunt patres eorum nominis mei propter Baal
JER|23|28|propheta qui habet somnium narret somnium et qui habet sermonem meum loquatur sermonem meum vere quid paleis ad triticum dicit Dominus
JER|23|29|numquid non verba mea sunt quasi ignis ait Dominus et quasi malleus conterens petram
JER|23|30|propterea ecce ego ad prophetas ait Dominus qui furantur verba mea unusquisque a proximo suo
JER|23|31|ecce ego ad prophetas ait Dominus qui adsumunt linguas suas et aiunt dicit Dominus
JER|23|32|ecce ego ad prophetas somniantes mendacium ait Dominus qui narraverunt ea et seduxerunt populum meum in mendacio suo et in miraculis suis cum ego non misissem eos nec mandassem eis qui nihil profuerunt populo huic dicit Dominus
JER|23|33|si igitur interrogaverit te populus iste vel propheta aut sacerdos dicens quod est onus Domini dices ad eos ut quid vobis onus proiciam quippe vos dicit Dominus
JER|23|34|et prophetes et sacerdos et populus qui dicit onus Domini visitabo super virum illum et super domum eius
JER|23|35|haec dicetis unusquisque ad proximum et ad fratrem suum quid respondit Dominus et quid locutus est Dominus
JER|23|36|et onus Domini ultra non memorabitur quia onus erit unicuique sermo suus et pervertitis verba Dei viventis Domini exercituum Dei nostri
JER|23|37|haec dices ad prophetam quid respondit tibi Dominus et quid locutus est Dominus
JER|23|38|si autem onus Domini dixeritis propter hoc haec dicit Dominus quia dixistis sermonem istum onus Domini et misi ad vos dicens nolite dicere onus Domini
JER|23|39|propterea ecce ego tollam vos portans et derelinquam vos et civitatem quam dedi vobis et patribus vestris a facie mea
JER|23|40|et dabo vos in obprobrium sempiternum et in ignominiam aeternam quae numquam oblivione delebitur
JER|24|1|ostendit mihi Dominus et ecce duo calathi pleni ficis positi ante templum Domini postquam transtulit Nabuchodonosor rex Babylonis Iechoniam filium Ioachim regem Iuda et principes eius et fabrum et inclusorem de Hierusalem et adduxit eos in Babylonem
JER|24|2|calathus unus ficus bonas habebat nimis ut solent ficus esse primi temporis et calathus unus ficus habebat malas nimis quae comedi non poterant eo quod essent malae
JER|24|3|et dixit Dominus ad me quid tu vides Hieremia et dixi ficus ficus bonas bonas valde et malas malas valde quae comedi non possunt eo quod sint malae
JER|24|4|et factum est verbum Domini ad me dicens
JER|24|5|haec dicit Dominus Deus Israhel sicut ficus hae bonae sic cognoscam transmigrationem Iuda quam emisi de loco isto in terram Chaldeorum in bonum
JER|24|6|et ponam oculos meos super eos ad placandum et reducam eos in terram hanc et aedificabo eos et non destruam et plantabo eos et non evellam
JER|24|7|et dabo eis cor ut sciant me quia ego sum Dominus et erunt mihi in populum et ego ero eis in Deum quia revertentur ad me in toto corde suo
JER|24|8|et sicut ficus pessimae quae comedi non possunt eo quod sint malae haec dicit Dominus sic dabo Sedeciam regem Iuda et principes eius et reliquos de Hierusalem qui remanserunt in urbe hac et qui habitant in terra Aegypti
JER|24|9|et dabo eos in vexationem adflictionemque omnibus regnis terrae in obprobrium et in parabolam et in proverbium et in maledictionem in universis locis ad quos eieci eos
JER|24|10|et mittam in eis gladium et famem et pestem donec consumantur de terra quam dedi eis et patribus eorum
JER|25|1|verbum quod factum est ad Hieremiam de omni populo Iudae in anno quarto Ioachim filii Iosiae regis Iuda ipse est annus primus Nabuchodonosor regis Babylonis
JER|25|2|quae locutus est Hieremias propheta ad omnem populum Iuda et ad universos habitatores Hierusalem dicens
JER|25|3|a tertiodecimo anno Iosiae filii Amon regis Iuda usque ad diem hanc iste est tertius et vicesimus annus factum est verbum Domini ad me et locutus sum ad vos de nocte consurgens et loquens et non audistis
JER|25|4|et misit Dominus ad vos omnes servos suos prophetas consurgens diluculo mittensque et non audistis neque inclinastis aures vestras ut audiretis
JER|25|5|cum diceret revertimini unusquisque a via sua mala et a pessimis cogitationibus vestris et habitabitis in terram quam dedit Dominus vobis et patribus vestris a saeculo et usque in saeculum
JER|25|6|et nolite ire post deos alienos ut serviatis eis adoretisque eos neque me ad iracundiam provocetis in operibus manuum vestrarum et non adfligam vos
JER|25|7|et non audistis me dicit Dominus ut me ad iracundiam provocaretis in operibus manuum vestrarum in malum vestrum
JER|25|8|propterea haec dicit Dominus exercituum pro eo quod non audistis verba mea
JER|25|9|ecce ego mittam et adsumam universas cognationes aquilonis ait Dominus et ad Nabuchodonosor regem Babylonis servum meum et adducam eos super terram istam et super habitatores eius et super omnes nationes quae in circuitu illius sunt et interficiam eos et ponam eos in stuporem et in sibilum et in solitudines sempiternas
JER|25|10|perdamque ex eis vocem gaudii et vocem laetitiae vocem sponsae et vocem sponsi vocem molae et lumen lucernae
JER|25|11|et erit universa terra eius in solitudinem et in stuporem et servient omnes gentes istae regi Babylonis septuaginta annis
JER|25|12|cumque impleti fuerint anni septuaginta visitabo super regem Babylonis et super gentem illam dicit Dominus iniquitatem eorum et super terram Chaldeorum et ponam illam in solitudines sempiternas
JER|25|13|et adducam super terram illam omnia verba mea quae locutus sum contra eam omne quod scriptum est in libro isto quaecumque prophetavit Hieremias adversum omnes gentes
JER|25|14|quia servierunt eis cum essent gentes multae et reges magni et reddam eis secundum opera eorum et secundum facta manuum suarum
JER|25|15|quia sic dicit Dominus exercituum Deus Israhel sume calicem vini furoris huius de manu mea et propinabis de illo cunctis gentibus ad quas ego mittam te
JER|25|16|et bibent et turbabuntur et insanient a facie gladii quem ego mittam inter eos
JER|25|17|et accepi calicem de manu Domini et propinavi cunctis gentibus ad quas misit me Dominus
JER|25|18|Hierusalem et civitatibus Iudae et regibus eius et principibus eius ut darem eos in solitudinem et in stuporem in sibilum et in maledictionem sicut est dies ista
JER|25|19|Pharaoni regi Aegypti et servis eius et principibus eius et omni populo eius
JER|25|20|et universis generaliter cunctis regibus terrae Ausitidis et cunctis regibus terrae Philisthim et Ascaloni et Gazae et Accaroni et reliquiis Azoti
JER|25|21|Idumeae et Moab et filiis Ammon
JER|25|22|et cunctis regibus Tyri et cunctis regibus Sidonis et regibus terrae insularum qui sunt trans mare
JER|25|23|et Dedan et Theman et Buz et universis qui adtonsi sunt in comam
JER|25|24|et cunctis regibus Arabiae et cunctis regibus occidentis qui habitant in deserto
JER|25|25|et cunctis regibus Zambri et cunctis regibus Aelam et cunctis regibus Medorum
JER|25|26|et cunctis regibus aquilonis de prope et de longe unicuique contra fratrem suum et omnibus regnis terrae quae super faciem eius sunt et rex Sesach bibet post eos
JER|25|27|et dices ad eos haec dicit Dominus exercituum Deus Israhel bibite et inebriamini et vomite et cadite neque surgatis a facie gladii quem ego mittam inter vos
JER|25|28|cumque noluerint accipere calicem de manu ut bibant dices ad eos haec dicit Dominus exercituum bibentes bibetis
JER|25|29|quia ecce in civitate in qua invocatum est nomen meum ego incipio adfligere et vos quasi innocentes inmunes eritis non eritis inmunes gladium enim ego voco super omnes habitatores terrae dicit Dominus exercituum
JER|25|30|et tu prophetabis ad eos omnia verba haec et dices ad illos Dominus de excelso rugiet et de habitaculo sancto suo dabit vocem suam rugiens rugiet super decorem suum celeuma quasi calcantium concinetur adversus omnes habitatores terrae
JER|25|31|pervenit sonitus usque ad extrema terrae quia iudicium Domino cum gentibus iudicatur ipse cum omni carne impios tradidit gladio dicit Dominus
JER|25|32|haec dicit Dominus exercituum ecce adflictio egredietur de gente in gentem et turbo magnus egredietur a summitatibus terrae
JER|25|33|et erunt interfecti Domini in die illa a summo terrae usque ad summum eius non plangentur et non colligentur neque sepelientur in sterquilinium super faciem terrae iacebunt
JER|25|34|ululate pastores et clamate et aspergite vos cinere optimates gregis quia conpleti sunt dies vestri ut interficiamini et dissipationes vestrae et cadetis quasi vasa pretiosa
JER|25|35|et peribit fuga a pastoribus et salvatio ab optimatibus gregis
JER|25|36|vox clamoris pastorum et ululatus optimatium gregis quia vastavit Dominus pascuam eorum
JER|25|37|et conticuerunt arva pacis a facie irae furoris Domini
JER|25|38|dereliquit quasi leo umbraculum suum facta est terra eorum in desolationem a facie irae columbae et a facie irae furoris Domini
JER|26|1|in principio regis Ioachim filii Iosiae regis Iuda factum est verbum istud a Domino dicens
JER|26|2|haec dicit Dominus sta in atrio domus Domini et loqueris ad omnes civitates Iuda de quibus veniunt ut adorent in domo Domini universos sermones quos ego mandavi tibi ut loquaris ad eos noli subtrahere verbum
JER|26|3|si forte audiant et convertantur unusquisque a via sua mala et paeniteat me mali quod cogito facere eis propter malitias studiorum eorum
JER|26|4|et dices ad eos haec dicit Dominus si non audieritis me ut ambuletis in lege mea quam dedi vobis
JER|26|5|ut audiatis sermones servorum meorum prophetarum quos ego misi ad vos de nocte consurgens et dirigens et non audistis
JER|26|6|dabo domum istam sicut Silo et urbem hanc dabo in maledictionem cunctis gentibus terrae
JER|26|7|et audierunt sacerdotes et prophetae et omnis populus Hieremiam loquentem verba haec in domo Domini
JER|26|8|cumque conplesset Hieremias loquens omnia quae praeceperat ei Dominus ut loqueretur ad universum populum adprehenderunt eum sacerdotes et prophetae et omnis populus dicens morte morietur
JER|26|9|quare prophetavit in nomine Domini dicens sicut Silo erit domus haec et urbs ista desolabitur eo quod non sit habitator et congregatus est omnis populus adversum Hieremiam in domum Domini
JER|26|10|et audierunt principes Iuda verba haec et ascenderunt de domo regis in domum Domini et sederunt in introitu portae Domini novae
JER|26|11|et locuti sunt sacerdotes et prophetae ad principes et ad omnem populum dicentes iudicium mortis est viro huic quia prophetavit adversum civitatem istam sicut audistis auribus vestris
JER|26|12|et ait Hieremias ad omnes principes et ad universum populum dicens Dominus misit me ut prophetarem ad domum istam et ad civitatem hanc omnia verba quae audistis
JER|26|13|nunc ergo bonas facite vias vestras et studia vestra et audite vocem Domini Dei vestri et paenitebit Dominum mali quod locutus est adversum vos
JER|26|14|ego autem ecce in manibus vestris sum facite mihi ut bonum et rectum est in oculis vestris
JER|26|15|verumtamen scitote et cognoscite quod si occideritis me sanguinem innocentem traditis contra vosmet ipsos et contra civitatem istam et habitatores eius in veritate enim misit me Dominus ad vos ut loquerer in auribus vestris omnia verba haec
JER|26|16|et dixerunt principes et omnis populus ad sacerdotes et prophetas non est viro huic iudicium mortis quia in nomine Domini Dei nostri locutus est ad nos
JER|26|17|surrexerunt ergo viri de senioribus terrae et dixerunt ad omnem coetum populi loquentes
JER|26|18|Michas de Morasthim fuit propheta in diebus Ezechiae regis Iudae et ait ad omnem populum Iudae dicens haec dicit Dominus exercituum Sion quasi ager arabitur et Hierusalem in acervum lapidum erit et mons domus in excelsa silvarum
JER|26|19|numquid morte condemnavit eum Ezechias rex Iuda et omnis Iuda numquid non timuerunt Dominum et deprecati sunt faciem Domini et paenituit Dominum mali quod locutus erat adversum eos itaque nos facimus malum grande contra animas nostras
JER|26|20|fuit quoque vir prophetans in nomine Domini Urias filius Semei de Cariathiarim et prophetavit adversum civitatem istam et adversum terram hanc iuxta universa verba Hieremiae
JER|26|21|et audivit rex Ioachim et omnes potentes et principes eius verba haec et quaesivit rex interficere eum et audivit Urias et timuit fugitque et ingressus est Aegyptum
JER|26|22|et misit rex Ioachim viros in Aegyptum Elnathan filium Achobor et viros cum eo in Aegyptum
JER|26|23|et eduxerunt Uriam de Aegypto et adduxerunt eum ad regem Ioachim et percussit eum gladio et proiecit cadaver eius in sepulchris vulgi ignobilis
JER|26|24|igitur manus Ahicam filii Saphan fuit cum Hieremia ut non traderetur in manu populi et interficerent eum
JER|27|1|in principio regni Ioachim filii Iosiae regis Iuda factum est verbum istud ad Hieremiam a Domino dicens
JER|27|2|haec dicit Dominus ad me fac tibi vincula et catenas et pones eas in collo tuo
JER|27|3|et mittes eas ad regem Edom et ad regem Moab et ad regem filiorum Ammon et ad regem Tyri et ad regem Sidonis in manu nuntiorum qui venerunt Hierusalem ad Sedeciam regem Iuda
JER|27|4|et praecipies eis ut ad dominos suos loquantur haec dicit Dominus exercituum Deus Israhel haec dicetis ad dominos vestros
JER|27|5|ego feci terram et hominem et iumenta quae sunt super faciem terrae in fortitudine mea magna et in brachio meo extento et dedi eam ei qui placuit in oculis meis
JER|27|6|et nunc itaque ego dedi omnes terras istas in manu Nabuchodonosor regis Babylonis servi mei insuper et bestias agri dedi ei ut serviant illi
JER|27|7|et servient ei omnes gentes et filio eius et filio filii eius donec veniat tempus terrae eius et ipsius et servient ei gentes multae et reges magni
JER|27|8|gens autem et regnum quod non servierit Nabuchodonosor regi Babylonis et quicumque non curvaverit collum suum sub iugo regis Babylonis in gladio et in fame et in peste visitabo super gentem illam ait Dominus donec consumam eos in manu eius
JER|27|9|vos ergo nolite audire prophetas vestros et divinos et somniatores et augures et maleficos qui dicunt vobis non servietis regi Babylonis
JER|27|10|quia mendacium prophetant vobis ut longe faciant vos de terra vestra et eiciant vos et pereatis
JER|27|11|porro gens quae subiecerit cervicem suam sub iugo regis Babylonis et servierit ei dimittam eam in terra sua dicit Dominus et colet eam et habitabit in ea
JER|27|12|et ad Sedeciam regem Iuda locutus sum secundum omnia verba haec dicens subicite colla vestra sub iugo regis Babylonis et servite ei et populo eius et vivetis
JER|27|13|quare moriemini tu et populus tuus gladio fame et peste sicut locutus est Dominus ad gentem quae servire noluerit regi Babylonis
JER|27|14|nolite audire verba prophetarum dicentium vobis non servietis regi Babylonis quia mendacium ipsi loquuntur vobis
JER|27|15|quia non misi eos ait Dominus et ipsi prophetant in nomine meo mendaciter ut eiciant vos et pereatis tam vos quam prophetae qui vaticinantur vobis
JER|27|16|et ad sacerdotes et ad populum istum locutus sum dicens haec dicit Dominus nolite audire verba prophetarum vestrorum qui prophetant vobis dicentes ecce vasa Domini revertentur de Babylone nunc cito mendacium enim prophetant vobis
JER|27|17|nolite ergo audire eos sed servite regi Babylonis ut vivatis quare datur haec civitas in solitudinem
JER|27|18|et si prophetae sunt et est verbum Domini in eis occurrant Domino exercituum ut non veniant vasa quae derelicta fuerant in domum Domini et in domum regis Iuda et in Hierusalem in Babylonem
JER|27|19|quia haec dicit Dominus exercituum ad columnas et ad mare et ad bases et ad reliqua vasorum quae remanserunt in civitate hac
JER|27|20|quae non tulit Nabuchodonosor rex Babylonis cum transferret Iechoniam filium Ioachim regem Iuda de Hierusalem in Babylonem et omnes optimates Iuda et Hierusalem
JER|27|21|quia haec dicit Dominus exercituum Deus Israhel ad vasa quae derelicta sunt in domum Domini et in domum regis Iuda et Hierusalem
JER|27|22|in Babylonem transferentur et ibi erunt usque ad diem visitationis suae dicit Dominus et adferri faciam ea et restitui in loco isto
JER|28|1|et factum est in anno illo in principio regni Sedeciae regis Iuda in anno quarto in mense quinto dixit ad me Ananias filius Azur propheta de Gabaon in domo Domini coram sacerdotibus et omni populo dicens
JER|28|2|haec dicit Dominus exercituum Deus Israhel contrivi iugum regis Babylonis
JER|28|3|adhuc duo anni dierum et ego referri faciam ad locum istum omnia vasa Domini quae tulit Nabuchodonosor rex Babylonis de loco isto et transtulit ea in Babylonem
JER|28|4|et Iechoniam filium Ioachim regem Iuda et omnem transmigrationem Iudae qui ingressi sunt in Babylonem ego convertam ad locum istum ait Dominus conteram enim iugum regis Babylonis
JER|28|5|et dixit Hieremias propheta ad Ananiam prophetam in oculis sacerdotum et in oculis omnis populi qui stabant in domo Domini
JER|28|6|et ait Hieremias propheta amen sic faciat Dominus suscitet Dominus verba tua quae prophetasti ut referantur vasa in domum Domini et omnis transmigratio de Babylone ad locum istum
JER|28|7|verumtamen audi verbum hoc quod ego loquor in auribus tuis et in auribus universi populi
JER|28|8|prophetae qui fuerunt ante me et te ab initio et prophetaverunt super terras multas et super regna magna de proelio et de adflictione et de fame
JER|28|9|propheta qui vaticinatus est pacem cum venerit verbum eius scietur propheta quem misit Dominus in veritate
JER|28|10|et tulit Ananias propheta catenam de collo Hieremiae prophetae et confregit eam
JER|28|11|et ait Ananias in conspectu omnis populi dicens haec dicit Dominus sic confringam iugum Nabuchodonosor regis Babylonis post duos annos dierum de collo omnium gentium
JER|28|12|et abiit Hieremias prophetes in viam suam et factum est verbum Domini ad Hieremiam postquam confregit Ananias propheta catenam de collo Hieremiae prophetae dicens
JER|28|13|vade et dices Ananiae haec dicit Dominus catenas ligneas contrivisti et facies pro eis catenas ferreas
JER|28|14|quia haec dicit Dominus exercituum Deus Israhel iugum ferreum posui super collum cunctarum gentium istarum ut serviant Nabuchodonosor regi Babylonis et servient ei insuper et bestias terrae dedi ei
JER|28|15|et dixit Hieremias propheta ad Ananiam prophetam audi Anania non misit te Dominus et tu confidere fecisti populum istum in mendacio
JER|28|16|idcirco haec dicit Dominus ecce emittam te a facie terrae hoc anno morieris adversum Dominum enim locutus es
JER|28|17|et mortuus est Ananias propheta in anno illo mense septimo
JER|29|1|et haec sunt verba libri quae misit Hieremias propheta de Hierusalem ad reliquias seniorum transmigrationis et ad sacerdotes et ad prophetas et ad omnem populum quem transduxerat Nabuchodonosor de Hierusalem in Babylonem
JER|29|2|postquam egressus est Iechonias rex et domina et eunuchi et principes Iuda et Hierusalem et faber et inclusor de Hierusalem
JER|29|3|in manu Ellasa filii Saphan et Gamaliae filii Helciae quos misit Sedecias rex Iuda ad Nabuchodonosor regem Babylonis in Babylonem dicens
JER|29|4|haec dicit Dominus exercituum Deus Israhel omni transmigrationi quam transtuli de Hierusalem in Babylonem
JER|29|5|aedificate domos et habitate et plantate hortos et comedite fructum eorum
JER|29|6|accipite uxores et generate filios et filias date filiis vestris uxores et filias vestras date viris et pariant filios et filias et multiplicamini ibi et nolite esse pauci numero
JER|29|7|et quaerite pacem civitatis ad quam transmigrare vos feci et orate pro ea ad Dominum quia in pace illius erit pax vobis
JER|29|8|haec enim dicit Dominus exercituum Deus Israhel non vos inducant prophetae vestri qui sunt in medio vestrum et divini vestri et ne adtendatis ad somnia vestra quae vos somniatis
JER|29|9|quia falso ipsi prophetant vobis in nomine meo et non misi eos dicit Dominus
JER|29|10|quia haec dicit Dominus cum coeperint impleri in Babylone septuaginta anni visitabo vos et suscitabo super vos verbum meum bonum ut reducam vos ad locum istum
JER|29|11|ego enim scio cogitationes quas cogito super vos ait Dominus cogitationes pacis et non adflictionis ut dem vobis finem et patientiam
JER|29|12|et invocabitis me et ibitis et orabitis me et exaudiam vos
JER|29|13|quaeretis me et invenietis cum quaesieritis me in toto corde vestro
JER|29|14|et inveniar a vobis ait Dominus et reducam captivitatem vestram et congregabo vos de universis gentibus et de cunctis locis ad quae expuli vos dicit Dominus et reverti vos faciam de loco ad quem transmigrare vos feci
JER|29|15|quia dixistis suscitavit nobis Dominus prophetas in Babylone
JER|29|16|quia haec dicit Dominus ad regem qui sedet super solium David et ad omnem populum habitatorem urbis huius ad fratres vestros qui non sunt egressi vobiscum in transmigrationem
JER|29|17|haec dicit Dominus exercituum ecce mittam in eis gladium et famem et pestem et ponam eos quasi ficus malas quae comedi non possunt eo quod pessimae sint
JER|29|18|et persequar eos in gladio in fame et in pestilentia et dabo eos in vexationem universis regnis terrae in maledictionem et in stuporem et in sibilum et in obprobrium cunctis gentibus ad quas ego eieci eos
JER|29|19|eo quod non audierint verba mea dicit Dominus quae misi ad eos per servos meos prophetas de nocte consurgens et mittens et non audistis dicit Dominus
JER|29|20|vos ergo audite verbum Domini omnis transmigratio quam emisi de Hierusalem in Babylonem
JER|29|21|haec dicit Dominus exercituum Deus Israhel ad Ahab filium Culia et ad Sedeciam filium Maasiae qui prophetant vobis in nomine meo mendaciter ecce ego tradam eos in manu Nabuchodonosor regis Babylonis et percutiet eos in oculis vestris
JER|29|22|et adsumetur ex eis maledictio omni transmigrationi Iuda quae est in Babylone dicentium ponat te Dominus sicut Sedeciam et sicut Ahab quos frixit rex Babylonis in igne
JER|29|23|pro eo quod fecerint stultitiam in Israhel et moechati sunt in uxores amicorum suorum et locuti sunt verbum in nomine meo mendaciter quod non mandavi eis ego sum iudex et testis dicit Dominus
JER|29|24|et ad Semeiam Neelamiten dices
JER|29|25|haec dicit Dominus exercituum Deus Israhel pro eo quod misisti in nomine tuo libros ad omnem populum qui est in Hierusalem et ad Sophoniam filium Maasiae sacerdotem et ad universos sacerdotes dicens
JER|29|26|Dominus dedit te sacerdotem pro Ioiadae sacerdote ut sis dux in domo Domini super omnem virum arrepticium et prophetantem ut mittas eum in nervum et in carcerem
JER|29|27|et nunc quare non increpasti Hieremiam Anathothiten qui prophetat vobis
JER|29|28|quia super hoc misit ad nos in Babylonem dicens longum est aedificate domos et habitate et plantate hortos et comedite fructum eorum
JER|29|29|legit ergo Sophonias sacerdos librum istum in auribus Hieremiae prophetae
JER|29|30|et factum est verbum Domini ad Hieremiam dicens
JER|29|31|mitte ad omnem transmigrationem dicens haec dicit Dominus ad Semeiam Neelamiten pro eo quod prophetavit vobis Semeias et ego non misi eum et fecit vos confidere in mendacio
JER|29|32|idcirco haec dicit Dominus ecce ego visitabo super Semeiam Neelamiten et super semen eius non erit ei vir sedens in medio populi huius et non videbit bonum quod ego faciam populo meo ait Dominus quia praevaricationem locutus est adversum Dominum
JER|30|1|hoc verbum quod factum est ad Hieremiam a Domino dicens
JER|30|2|haec dicit Dominus Deus Israhel dicens scribe tibi omnia verba quae locutus sum ad te in libro
JER|30|3|ecce enim dies veniunt dicit Dominus et convertam conversionem populi mei Israhel et Iuda ait Dominus et convertam eos ad terram quam dedi patribus eorum et possidebunt eam
JER|30|4|et haec verba quae locutus est Dominus ad Israhel et ad Iudam
JER|30|5|quoniam haec dicit Dominus vocem terroris audivimus formido et non est pax
JER|30|6|interrogate et videte si generat masculus quare ergo vidi omnis viri manum super lumbum suum quasi parientis et conversae sunt universae facies in auruginem
JER|30|7|vae quia magna dies illa nec est similis eius tempusque tribulationis est Iacob et ex ipso salvabitur
JER|30|8|et erit in die illa ait Dominus exercituum conteram iugum eius de collo tuo et vincula illius disrumpam et non dominabuntur ei amplius alieni
JER|30|9|sed servient Domino Deo suo et David regi suo quem suscitabo eis
JER|30|10|tu ergo ne timeas serve meus Iacob ait Dominus neque paveas Israhel quia ecce ego salvo te de terra longinqua et semen tuum de terra captivitatis eorum et revertetur Iacob et quiescet et cunctis affluet et non erit quem formidet
JER|30|11|quoniam tecum ego sum ait Dominus ut salvem te faciam enim consummationem in cunctis gentibus in quibus dispersi te te autem non faciam in consummationem sed castigabo te in iudicio ut non tibi videaris innoxius
JER|30|12|quia haec dicit Dominus insanabilis fractura tua pessima plaga tua
JER|30|13|non est qui iudicet iudicium tuum ad alligandum curationum utilitas non est tibi
JER|30|14|omnes amatores tui obliti sunt tui te non quaerent plaga enim inimici percussi te castigatione crudeli propter multitudinem iniquitatis tuae dura facta sunt peccata tua
JER|30|15|quid clamas super contritione tua insanabilis est dolor tuus propter multitudinem iniquitatis tuae et dura peccata tua feci haec tibi
JER|30|16|propterea omnes qui comedunt te devorabuntur et universi hostes tui in captivitatem ducentur et qui te vastant vastabuntur cunctosque praedatores tuos dabo in praedam
JER|30|17|obducam enim cicatricem tibi et a vulneribus tuis sanabo te dicit Dominus quia Eiectam vocaverunt te Sion haec est quae non habebat requirentem
JER|30|18|haec dicit Dominus ecce ego convertam conversionem tabernaculorum Iacob et tectis eius miserebor et aedificabitur civitas in excelso suo et templum iuxta ordinem suum fundabitur
JER|30|19|et egredietur de eis laus voxque ludentium et multiplicabo eos et non inminuentur et glorificabo eos et non adtenuabuntur
JER|30|20|et erunt filii eius sicut a principio et coetus eius coram me permanebit et visitabo adversum omnes qui tribulant eum
JER|30|21|et erit dux eius ex eo et princeps de medio eius producetur et adplicabo eum et accedet ad me quis enim iste est qui adplicet cor suum ut adpropinquet mihi ait Dominus
JER|30|22|et eritis mihi in populum et ego ero vobis in Deum
JER|30|23|ecce turbo Domini furor egrediens procella ruens in capite impiorum conquiescet
JER|30|24|non avertet iram indignationis Dominus donec faciat et conpleat cogitationem cordis sui in novissimo dierum intellegetis ea
JER|31|1|in tempore illo dicit Dominus ero Deus universis cognationibus Israhel et ipsi erunt mihi in populum
JER|31|2|haec dicit Dominus invenit gratiam in deserto populus qui remanserat gladio vadet ad requiem suam Israhel
JER|31|3|longe Dominus apparuit mihi et in caritate perpetua dilexi te ideo adtraxi te miserans
JER|31|4|rursumque aedificabo te et aedificaberis virgo Israhel adhuc ornaberis tympanis tuis et egredieris in choro ludentium
JER|31|5|adhuc plantabis vineas in montibus Samariae plantabunt plantantes et donec tempus veniat non vindemiabunt
JER|31|6|quia erit dies in qua clamabunt custodes in monte Ephraim surgite et ascendamus in Sion ad Dominum Deum nostrum
JER|31|7|quia haec dicit Dominus exultate in laetitia Iacob et hinnite contra caput gentium personate canite et dicite salva Domine populum tuum reliquias Israhel
JER|31|8|ecce ego adducam eos de terra aquilonis et congregabo eos ab extremis terrae inter quos erunt caecus et claudus et praegnans et pariens simul coetus magnus revertentium huc
JER|31|9|in fletu venient et in precibus deducam eos et adducam eos per torrentes aquarum in via recta et non inpingent in ea quia factus sum Israheli pater et Ephraim primogenitus meus est
JER|31|10|audite verbum Domini gentes et adnuntiate insulis quae procul sunt et dicite qui dispersit Israhel congregabit eum et custodiet eum sicut pastor gregem suum
JER|31|11|redemit enim Dominus Iacob et liberavit eum de manu potentioris
JER|31|12|et venient et laudabunt in monte Sion et confluent ad bona Domini super frumento et vino et oleo et fetu pecorum et armentorum eritque anima eorum quasi hortus inriguus et ultra non esurient
JER|31|13|tunc laetabitur virgo in choro iuvenes et senes simul et convertam luctum eorum in gaudium et consolabor eos et laetificabo a dolore suo
JER|31|14|et inebriabo animam sacerdotum pinguedine et populus meus bonis meis adimplebitur ait Dominus
JER|31|15|haec dicit Dominus vox in excelso audita est lamentationis fletus et luctus Rachel plorantis filios suos et nolentis consolari super eis quia non sunt
JER|31|16|haec dicit Dominus quiescat vox tua a ploratu et oculi tui a lacrimis quia est merces operi tuo ait Dominus et revertentur de terra inimici
JER|31|17|et est spes novissimis tuis ait Dominus et revertentur filii ad terminos suos
JER|31|18|audiens audivi Ephraim transmigrantem castigasti me et eruditus sum quasi iuvenculus indomitus converte me et revertar quia tu Dominus Deus meus
JER|31|19|postquam enim convertisti me egi paenitentiam et postquam ostendisti mihi percussi femur meum confusus sum et erubui quoniam sustinui obprobrium adulescentiae meae
JER|31|20|si filius honorabilis mihi Ephraim si puer delicatus quia ex quo locutus sum de eo adhuc recordabor eius idcirco conturbata sunt viscera mea super eum miserans miserebor eius ait Dominus
JER|31|21|statue tibi speculam pone tibi amaritudines dirige cor tuum in viam directam in qua ambulasti revertere virgo Israhel revertere ad civitates tuas istas
JER|31|22|usquequo deliciis dissolveris filia vaga quia creavit Dominus novum super terram femina circumdabit virum
JER|31|23|haec dicit Dominus exercituum Deus Israhel adhuc dicent verbum istud in terra Iuda et in urbibus eius cum convertero captivitatem eorum benedicat tibi Dominus pulchritudo iustitiae mons sanctus
JER|31|24|et habitabunt in eo Iudas et omnes civitates eius simul agricolae et minantes greges
JER|31|25|quia inebriavi animam lassam et omnem animam esurientem saturavi
JER|31|26|ideo quasi de somno suscitatus sum et vidi et somnus meus dulcis mihi
JER|31|27|ecce dies veniunt dicit Dominus et seminabo domum Israhel et domum Iuda semine hominis et semine iumentorum
JER|31|28|et sicut vigilavi super eos ut evellerem et demolirer et dissiparem et disperderem et adfligerem sic vigilabo super eos ut aedificem et plantem ait Dominus
JER|31|29|in diebus illis non dicent ultra patres comederunt uvam acerbam et dentes filiorum obstipuerunt
JER|31|30|sed unusquisque in iniquitate sua morietur omnis homo qui comederit uvam acerbam obstupescent dentes eius
JER|31|31|ecce dies veniunt dicit Dominus et feriam domui Israhel et domui Iuda foedus novum
JER|31|32|non secundum pactum quod pepigi cum patribus vestris in die qua adprehendi manum eorum ut educerem eos de terra Aegypti pactum quod irritum fecerunt et ego dominatus sum eorum dicit Dominus
JER|31|33|sed hoc erit pactum quod feriam cum domo Israhel post dies illos dicit Dominus dabo legem meam in visceribus eorum et in corde eorum scribam eam et ero eis in Deum et ipsi erunt mihi in populum
JER|31|34|et non docebunt ultra vir proximum suum et vir fratrem suum dicens cognoscite Dominum omnes enim cognoscent me a minimo eorum usque ad maximum ait Dominus quia propitiabor iniquitati eorum et peccati eorum non ero memor amplius
JER|31|35|haec dicit Dominus qui dat solem in lumine diei ordinem lunae et stellarum in lumine noctis qui turbat mare et sonant fluctus eius Dominus exercituum nomen illi
JER|31|36|si defecerint leges istae coram me dicit Dominus tunc et semen Israhel deficiet ut non sit gens coram me cunctis diebus
JER|31|37|haec dicit Dominus si mensurari potuerint caeli sursum et investigari fundamenta terrae deorsum et ego abiciam universum semen Israhel propter omnia quae fecerunt dicit Dominus
JER|31|38|ecce dies veniunt dicit Dominus et aedificabitur civitas Domino a turre Ananehel usque ad portam Anguli
JER|31|39|et exibit ultra norma mensurae in conspectu eius super collem Gareb et circuibit Goatha
JER|31|40|et omnem vallem cadaverum et cineris et universam regionem mortis usque ad torrentem Cedron et usque ad angulum portae Equorum orientalis sanctum Domini non evelletur et non destruetur ultra in perpetuum
JER|32|1|verbum quod factum est ad Hieremiam a Domino in anno decimo Sedeciae regis Iuda ipse est annus octavusdecimus Nabuchodonosor
JER|32|2|tunc exercitus regis Babylonis obsidebat Hierusalem et Hieremias propheta erat clausus in atrio carceris qui erat in domo regis Iuda
JER|32|3|clauserat enim eum Sedecias rex Iuda dicens quare vaticinaris dicens haec dicit Dominus ecce ego dabo civitatem istam in manu regis Babylonis et capiet eam
JER|32|4|et Sedecias rex Iuda non effugiet de manu Chaldeorum sed tradetur in manu regis Babylonis et loquetur os eius cum ore illius et oculi eius oculos illius videbunt
JER|32|5|et in Babylonem ducet Sedeciam et ibi erit donec visitem eum ait Dominus si autem dimicaveritis adversum Chaldeos nihil prosperum habebitis
JER|32|6|et dixit Hieremias factum est verbum Domini ad me dicens
JER|32|7|ecce Anamehel filius Sellum patruelis tuus veniet ad te dicens eme tibi agrum meum qui est in Anathoth tibi enim conpetit ex propinquitate ut emas
JER|32|8|et venit ad me Anamehel filius patrui mei secundum verbum Domini ad vestibulum carceris et ait ad me posside agrum meum qui est in Anathoth in terra Beniamin quia tibi conpetit hereditas et tu propinquus ut possideas intellexi autem quod verbum Domini esset
JER|32|9|et emi agrum ab Anamehel filio patrui mei qui est in Anathoth et adpendi ei argentum septem stateres et decem argenteos
JER|32|10|et scripsi in libro et signavi et adhibui testes et adpendi argentum in statera
JER|32|11|et accepi librum possessionis signatum stipulationes et rata et signa forinsecus
JER|32|12|et dedi librum possessionis Baruch filio Neri filii Maasiae in oculis Anamehel patruelis mei et in oculis testium qui scripti erant in libro emptionis in oculis omnium Iudaeorum qui sedebant in atrio carceris
JER|32|13|et praecepi Baruch coram eis dicens
JER|32|14|haec dicit Dominus exercituum Deus Israhel sume libros istos librum emptionis hunc signatum et librum hunc qui apertus est et pones illos in vase fictili ut permanere possint diebus multis
JER|32|15|haec enim dicit Dominus exercituum Deus Israhel adhuc possidebuntur domus et agri et vineae in terra ista
JER|32|16|et oravi ad Dominum postquam tradidi librum possessionis Baruch filio Neri dicens
JER|32|17|heu heu heu Domine Deus ecce tu fecisti caelum et terram in fortitudine tua magna et in brachio tuo extento non erit tibi difficile omne verbum
JER|32|18|qui facis misericordiam in milibus et reddes iniquitatem patrum in sinu filiorum eorum post eos fortissime magne potens Dominus exercituum nomen tibi
JER|32|19|magnus consilio et inconprehensibilis cogitatu cuius oculi aperti sunt super omnes vias filiorum Adam ut reddas unicuique secundum vias suas et secundum fructum adinventionum eius
JER|32|20|qui posuisti signa et portenta in terra Aegypti usque ad diem hanc et in Israhel et in hominibus et fecisti tibi nomen sicut est dies haec
JER|32|21|et eduxisti populum tuum Israhel de terra Aegypti in signis et in portentis et in manu robusta et in brachio extento et in terrore magno
JER|32|22|et dedisti eis terram hanc quam iurasti patribus eorum ut dares eis terram fluentem lacte et melle
JER|32|23|et ingressi sunt et possederunt eam et non oboedierunt voci tuae et in lege tua non ambulaverunt omnia quae mandasti eis ut facerent non fecerunt et evenerunt eis omnia mala haec
JER|32|24|ecce munitiones extructae sunt adversum civitatem ut capiatur et urbs data est in manu Chaldeorum qui proeliantur adversum eam a facie gladii et famis et pestilentiae et quaecumque locutus es acciderunt ut ipse tu cernis
JER|32|25|et tu dicis mihi Domine Deus eme agrum argento et adhibe testes cum urbs data sit in manu Chaldeorum
JER|32|26|et factum est verbum Domini ad Hieremiam dicens
JER|32|27|ecce ego Dominus Deus universae carnis numquid mihi difficile erit omne verbum
JER|32|28|propterea haec dicit Dominus ecce ego tradam civitatem istam in manu Chaldeorum et in manu regis Babylonis et capiet eam
JER|32|29|et venient Chaldei proeliantes adversum urbem hanc et succendent eam igni et conburent eam et domos in quarum domatibus sacrificabant Baal et libabant diis alienis libamina ad inritandum me
JER|32|30|erant enim filii Israhel et filii Iuda iugiter facientes malum in oculis meis ab adulescentia sua filii Israhel qui usque nunc exacerbant me in opere manuum suarum dicit Dominus
JER|32|31|quia in furore et in indignatione mea facta est mihi civitas haec a die qua aedificaverunt eam usque ad diem istam qua aufertur de conspectu meo
JER|32|32|propter malitiam filiorum Israhel et filiorum Iuda quam fecerunt ad iracundiam me provocantes ipsi et reges eorum principes eorum et sacerdotes et prophetae eorum vir Iuda et habitatores Hierusalem
JER|32|33|et verterunt ad me terga et non facies cum docerem eos diluculo et erudirem et nollent audire ut acciperent disciplinam
JER|32|34|et posuerunt idola sua in domo in qua invocatum est nomen meum ut polluerent eam
JER|32|35|et aedificaverunt excelsa Baal quae sunt in valle filii Ennom ut initiarent filios suos et filias suas Moloch quod non mandavi eis nec ascendit in cor meum ut facerent abominationem hanc et in peccatum deducerent Iudam
JER|32|36|et nunc propter ista haec dicit Dominus Deus Israhel ad civitatem hanc de qua vos dicitis quod tradatur in manu regis Babylonis in gladio et in fame et in peste
JER|32|37|ecce ego congregabo eos de universis terris ad quas eieci eos in furore meo et in ira mea et in indignatione grandi et reducam eos ad locum istum et habitare eos faciam confidenter
JER|32|38|et erunt mihi in populum et ego ero eis in Deum
JER|32|39|et dabo eis cor unum et viam unam ut timeant me universis diebus et bene sit eis et filiis eorum post eos
JER|32|40|et feriam eis pactum sempiternum et non desinam eis benefacere et timorem meum dabo in corde eorum ut non recedant a me
JER|32|41|et laetabor super eis cum bene eis fecero et plantabo eos in terra ista in veritate in toto corde meo et in tota anima mea
JER|32|42|quia haec dicit Dominus sicut adduxi super populum istum omne malum hoc grande sic adducam super eos omne bonum quod ego loquor ad eos
JER|32|43|et possidebuntur agri in terra ista de qua vos dicitis quod deserta sit eo quod non remanserit homo et iumentum et data sit in manu Chaldeorum
JER|32|44|agri pecunia ementur et scribentur in libro et inprimetur signum et testis adhibebitur in terra Beniamin et in circuitu Hierusalem in civitatibus Iuda et in civitatibus montanis et in civitatibus campestribus et in civitatibus quae ad austrum sunt quia convertam captivitatem eorum ait Dominus
JER|33|1|et factum est verbum Domini ad Hieremiam secundo cum adhuc clausus esset in atrio carceris dicens
JER|33|2|haec dicit Dominus qui facturus est Dominus et formaturus illud et paraturus Dominus nomen eius
JER|33|3|clama ad me et exaudiam te et adnuntiabo tibi grandia et firma quae nescis
JER|33|4|quia haec dicit Dominus Deus Israhel ad domos urbis huius et ad domos regis Iuda quae destructae sunt et ad munitiones et gladium
JER|33|5|venientium ut dimicent cum Chaldeis et impleant eas cadaveribus hominum quas percussi in furore meo et in indignatione mea abscondens faciem meam a civitate hac propter omnem malitiam eorum
JER|33|6|ecce ego obducam ei cicatricem et sanitatem et curabo eos et revelabo illis deprecationem pacis et veritatis
JER|33|7|et convertam conversionem Iuda et conversionem Hierusalem et aedificabo eos sicut a principio
JER|33|8|et emundabo illos ab omni iniquitate sua in qua peccaverunt mihi et propitius ero cunctis iniquitatibus eorum in quibus deliquerunt mihi et spreverunt me
JER|33|9|et erit mihi in nomen et in gaudium et in laudem et in exultationem cunctis gentibus terrae quae audierint omnia bona quae ego facturus sum eis et pavebunt et turbabuntur in universis bonis et in omni pace quam ego faciam ei
JER|33|10|haec dicit Dominus adhuc audietur in loco isto quem vos dicitis esse desertum eo quod non sit homo et iumentum in civitatibus Iuda et foris Hierusalem quae desolatae sunt absque homine et absque habitatore et absque pecore
JER|33|11|vox gaudii et vox laetitiae vox sponsi et vox sponsae vox dicentium confitemini Domino exercituum quoniam bonus Dominus quoniam in aeternum misericordia eius et portantium vota in domum Domini reducam enim conversionem terrae sicut a principio dicit Dominus
JER|33|12|haec dicit Dominus exercituum adhuc erit in loco isto deserto absque homine et absque iumento et in cunctis civitatibus eius habitaculum pastorum accubantium gregum
JER|33|13|in civitatibus montuosis et in civitatibus campestribus et in civitatibus quae ad austrum sunt et in terra Beniamin et in circuitu Hierusalem et in civitatibus Iuda adhuc transibunt greges ad manum numerantis ait Dominus
JER|33|14|ecce dies veniunt dicit Dominus et suscitabo verbum bonum quod locutus sum ad domum Israhel et ad domum Iuda
JER|33|15|in diebus illis et in tempore illo germinare faciam David germen iustitiae et faciet iudicium et iustitiam in terra
JER|33|16|in diebus illis salvabitur Iuda et Hierusalem habitabit confidenter et hoc est quod vocabit eam Dominus iustus noster
JER|33|17|quia haec dicit Dominus non interibit de David vir qui sedeat super thronum domus Israhel
JER|33|18|et de sacerdotibus et Levitis non interibit vir a facie mea qui offerat holocaustomata et incendat sacrificium et caedat victimas cunctis diebus
JER|33|19|et factum est verbum Domini ad Hieremiam dicens
JER|33|20|haec dicit Dominus si irritum fieri potest pactum meum cum die et pactum meum cum nocte ut non sit dies et nox in tempore suo
JER|33|21|et pactum meum irritum esse poterit cum David servo meo ut non sit ex eo filius qui regnet in throno eius et Levitae et sacerdotes ministri mei
JER|33|22|sicuti numerari non possunt stellae caeli et metiri harena maris sic multiplicabo semen David servi mei et Levitas ministros meos
JER|33|23|et factum est verbum Domini ad Hieremiam dicens
JER|33|24|numquid non vidisti quid populus hic locutus sit dicens duae cognationes quas elegerat Dominus abiectae sunt et populum meum despexerunt eo quod non sit ultra gens coram eis
JER|33|25|haec dicit Dominus si pactum meum inter diem et noctem et leges caelo et terrae non posui
JER|33|26|equidem et semen Iacob et David servi mei proiciam ut non adsumam de semine eius principes seminis Abraham et Isaac et Iacob reducam enim conversionem eorum et miserebor eis
JER|34|1|verbum quod factum est ad Hieremiam a Domino quando Nabuchodonosor rex Babylonis et omnis exercitus eius universaque regna terrae quae erant sub potestate manus eius et omnes populi bellabant contra Hierusalem et contra omnes urbes eius dicens
JER|34|2|haec dicit Dominus Deus Israhel vade et loquere ad Sedeciam regem Iuda et dices ad eum haec dicit Dominus ecce ego tradam civitatem hanc in manu regis Babylonis et succendet eam igni
JER|34|3|et tu non effugies de manu eius sed conprehensione capieris et in manu eius traderis et oculi tui oculos regis Babylonis videbunt et os eius cum ore tuo loquetur et Babylonem introibis
JER|34|4|attamen audi verbum Domini Sedecia rex Iuda haec dicit Dominus ad te non morieris in gladio
JER|34|5|sed in pace morieris et secundum conbustiones patrum tuorum regum priorum qui fuerunt ante te sic conburent te et vae domine plangent te quia verbum ego locutus sum dicit Dominus
JER|34|6|et locutus est Hieremias propheta ad Sedeciam regem Iuda universa verba haec in Hierusalem
JER|34|7|et exercitus regis Babylonis pugnabat contra Hierusalem et contra omnes civitates Iuda quae reliquae erant contra Lachis et contra Azeca haec enim supererant de civitatibus Iuda urbes munitae
JER|34|8|verbum quod factum est ad Hieremiam a Domino postquam percussit rex Sedecias foedus cum omni populo in Hierusalem praedicans
JER|34|9|ut dimitteret unusquisque servum suum et unusquisque ancillam suam hebraeum et hebraeam liberos et nequaquam dominarentur eis id est in Iudaeo et fratre suo
JER|34|10|audierunt ergo omnes principes et universus populus qui inierant pactum ut dimitteret unusquisque servum suum et unusquisque ancillam suam liberos et ultra non dominarentur in eis audierunt igitur et dimiserunt
JER|34|11|et conversi sunt deinceps et retraxerunt servos et ancillas suas quos dimiserant liberos et subiugaverunt in famulos et in famulas
JER|34|12|et factum est verbum Domini ad Hieremiam a Domino dicens
JER|34|13|haec dicit Dominus Deus Israhel ego percussi foedus cum patribus vestris in die qua eduxi eos de terra Aegypti de domo servitutis dicens
JER|34|14|cum conpleti fuerint septem anni dimittat unusquisque fratrem suum hebraeum qui venditus est ei et serviet tibi sex annis et dimittes eum a te liberum et non audierunt patres vestri me nec inclinaverunt aurem suam
JER|34|15|et conversi estis vos hodie et fecistis quod rectum est in oculis meis ut praedicaretis libertatem unusquisque ad amicum suum et inistis pactum in conspectu meo in domo in qua invocatum est nomen meum super eam
JER|34|16|et reversi estis et commaculastis nomen meum et reduxistis unusquisque servum suum et unusquisque ancillam suam quos dimiseratis ut essent liberi et suae potestatis et subiugastis eos ut sint vobis servi et ancillae
JER|34|17|propterea haec dicit Dominus vos non audistis me ut praedicaretis libertatem unusquisque fratri suo et unusquisque amico suo ecce ego praedico libertatem ait Dominus ad gladium et pestem et famem et dabo vos in commotionem cunctis regnis terrae
JER|34|18|et dabo viros qui praevaricantur foedus meum et non observaverunt verba foederis quibus adsensi sunt in conspectu meo vitulum quem ceciderunt in duas partes et transierunt inter divisiones eius
JER|34|19|principes Iuda et principes Hierusalem eunuchi et sacerdotes et omnis populus terrae qui transierunt inter divisiones vituli
JER|34|20|et dabo eos in manu inimicorum suorum et in manu quaerentium animam eorum et erit morticinum eorum in escam volucribus caeli et bestiis terrae
JER|34|21|et Sedeciam regem Iuda et principes eius dabo in manu inimicorum suorum et in manu quaerentium animam eorum et in manu exercituum regis Babylonis qui recesserunt a vobis
JER|34|22|ecce ego praecipio dicit Dominus et reducam eos in civitatem hanc et proeliabuntur adversum eam et capient eam et incendent igni et civitates Iuda dabo in solitudinem eo quod non sit habitator
JER|35|1|verbum quod factum est ad Hieremiam a Domino in diebus Ioachim filii Iosiae regis Iuda dicens
JER|35|2|vade ad domum Rechabitarum et loquere eis et introduces eos in domum Domini in unam exedram thesaurorum et dabis eis bibere vinum
JER|35|3|et adsumpsi Iezoniam filium Hieremiae filii Absaniae et fratres eius et omnes filios eius et universam domum Rechabitarum
JER|35|4|et introduxi eos in domum Domini ad gazofilacium filiorum Anan filii Hiegedeliae hominis Dei quod erat iuxta gazofilacium principum super thesaurum Maasiae filii Sellum qui erat custos vestibuli
JER|35|5|et posui coram filiis domus Rechabitarum scyphos plenos vino et calices et dixi ad eos bibite vinum
JER|35|6|qui responderunt non bibemus vinum quia Ionadab filius Rechab pater noster praecepit nobis dicens non bibetis vinum vos et filii vestri usque in sempiternum
JER|35|7|et domum non aedificabitis et sementem non seretis et vineas non plantabitis nec habebitis sed in tabernaculis habitabitis cunctis diebus vestris ut vivatis diebus multis super faciem terrae in qua vos peregrinamini
JER|35|8|oboedivimus ergo voci Ionadab filii Rechab patris nostri in omnibus quae praecepit nobis ita ut non biberemus vinum cunctis diebus nostris nos et mulieres nostrae filii et filiae nostrae
JER|35|9|et non aedificaremus domos ad habitandum et vineam et agrum et sementem non habuimus
JER|35|10|sed habitavimus in tabernaculis et oboedientes fecimus iuxta omnia quae praecepit nobis Ionadab pater noster
JER|35|11|cum autem ascendisset Nabuchodonosor rex Babylonis ad terram nostram diximus venite et ingrediamur Hierusalem a facie exercitus Chaldeorum et a facie exercitus Syriae et mansimus in Hierusalem
JER|35|12|et factum est verbum Domini ad Hieremiam dicens
JER|35|13|haec dicit Dominus exercituum Deus Israhel vade et dic viris Iuda et habitatoribus Hierusalem numquid non recipietis disciplinam ut oboediatis verbis meis dicit Dominus
JER|35|14|praevaluerunt sermones Ionadab filii Rechab quos praecepit filiis suis ut non biberent vinum et non biberunt usque ad diem hanc quia oboedierunt praecepto patris sui ego autem locutus sum ad vos de mane consurgens et loquens et non oboedistis mihi
JER|35|15|misique ad vos omnes servos meos prophetas consurgens diluculo mittensque et dicens convertimini unusquisque a via sua pessima et bona facite studia vestra et nolite sequi deos alienos neque colatis eos et habitabitis in terra quam dedi vobis et patribus vestris et non inclinastis aurem vestram neque audistis me
JER|35|16|firmaverunt igitur filii Ionadab filii Rechab praeceptum patris sui quod praeceperat eis populus autem iste non oboedivit mihi
JER|35|17|idcirco haec dicit Dominus exercituum Deus Israhel ecce ego adduco super Iudam et super omnes habitatores Hierusalem universam adflictionem quam locutus sum adversum eos eo quod locutus sum ad illos et non audierunt vocavi illos et non responderunt mihi
JER|35|18|domui autem Rechabitarum dixit Hieremias haec dicit Dominus exercituum Deus Israhel pro eo quod oboedistis praecepto Ionadab patris vestri et custodistis omnia mandata eius et fecistis universa quae praecepit vobis
JER|35|19|propterea haec dicit Dominus exercituum Deus Israhel non deficiet vir de stirpe Ionadab filii Rechab stans in conspectu meo cunctis diebus
JER|36|1|et factum est in anno quarto Ioachim filii Iosiae regis Iuda factum est verbum hoc ad Hieremiam a Domino dicens
JER|36|2|tolle volumen libri et scribes in eo omnia verba quae locutus sum tibi adversum Israhel et Iudam et adversum omnes gentes a die qua locutus sum ad te ex diebus Iosiae usque ad diem hanc
JER|36|3|si forte audiente domo Iuda universa mala quae ego cogito facere eis revertatur unusquisque a via sua pessima et propitius ero iniquitati et peccato eorum
JER|36|4|vocavit ergo Hieremias Baruch filium Neriae et scripsit Baruch ex ore Hieremiae omnes sermones Domini quos locutus est ad eum in volumine libri
JER|36|5|et praecepit Hieremias Baruch dicens ego clausus sum nec valeo ingredi domum Domini
JER|36|6|ingredere ergo tu et lege de volumine in quo scripsisti ex ore meo verba Domini audiente populo in domo Domini in die ieiunii insuper et audiente universo Iuda qui veniunt de civitatibus suis leges eis
JER|36|7|si forte cadat oratio eorum in conspectu Domini et revertatur unusquisque a via sua pessima quoniam magnus furor et indignatio quam locutus est Dominus adversum populum hunc
JER|36|8|et fecit Baruch filius Neriae iuxta omnia quae praeceperat ei Hieremias propheta legens ex volumine sermones Domini in domo Domini
JER|36|9|factum est autem in anno quinto Ioachim filii Iosiae regis Iuda in mense nono praedicaverunt ieiunium in conspectu Domini omni populo in Hierusalem et universae multitudini quae confluxerat de civitatibus Iuda in Hierusalem
JER|36|10|legitque Baruch ex volumine sermones Hieremiae in domo Domini in gazofilacio Gamariae filii Saphan scribae in vestibulo superiori in introitu portae novae domus Domini audiente omni populo
JER|36|11|cumque audisset Micheas filius Gamariae filii Saphan omnes sermones Domini ex libro
JER|36|12|descendit in domum regis ad gazofilacium scribae et ecce ibi omnes principes sedebant Elisama scriba et Dalaias filius Semeiae et Elnathan filius Achobor et Gamarias filius Saphan et Sedecias filius Ananiae et universi principes
JER|36|13|et nuntiavit eis Micheas omnia verba quae audivit legente Baruch ex volumine in auribus populi
JER|36|14|miserunt itaque omnes principes ad Baruch Iudi filium Nathaniae filii Selemiae filii Chusi dicentes volumen ex quo legisti audiente populo sume in manu tua et veni tulit ergo Baruch filius Neriae volumen in manu sua et venit ad eos
JER|36|15|et dixerunt ad eum sede et lege haec in auribus nostris et legit Baruch in auribus eorum
JER|36|16|igitur cum audissent omnia verba obstipuerunt unusquisque ad proximum suum et dixerunt ad Baruch nuntiare debemus regi omnes sermones istos
JER|36|17|et interrogaverunt eum dicentes indica nobis quomodo scripsisti omnes sermones istos ex ore eius
JER|36|18|dixit autem eis Baruch ex ore suo loquebatur quasi legens ad me omnes sermones istos et ego scribebam in volumine atramento
JER|36|19|et dixerunt principes ad Baruch vade et abscondere tu et Hieremias et nemo sciat ubi sitis
JER|36|20|et ingressi sunt ad regem in atrium porro volumen commendaverunt in gazofilacio Elisamae scribae et nuntiaverunt audiente rege omnes sermones
JER|36|21|misitque rex Iudi ut sumeret volumen qui tollens illud de gazofilacio Elisamae scribae legit audiente rege et universis principibus qui stabant circa regem
JER|36|22|rex autem sedebat in domo hiemali in mense nono et posita erat arula coram eo plena prunis
JER|36|23|cumque legisset Iudi tres pagellas vel quattuor scidit illud scalpello scribae et proiecit in igne qui erat super arulam donec consumeretur omne volumen igni qui erat in arula
JER|36|24|et non timuerunt neque sciderunt vestimenta sua rex et omnes servi eius qui audierunt universos sermones istos
JER|36|25|verumtamen Elnathan et Dalaias et Gamarias contradixerunt regi ne conbureret librum et non audivit eos
JER|36|26|et praecepit rex Hieremahel filio Ammelech et Saraiae filio Ezrihel et Selemiae filio Abdehel ut conprehenderent Baruch scribam et Hieremiam prophetam abscondit autem eos Dominus
JER|36|27|et factum est verbum Domini ad Hieremiam postquam conbuserat rex volumen et sermones quos scripserat Baruch ex ore Hieremiae dicens
JER|36|28|rursum tolle volumen aliud et scribe in eo omnes sermones priores qui erant in volumine primo quod conbusit Ioachim rex Iuda
JER|36|29|et ad Ioachim regem Iuda dices haec dicit Dominus tu conbusisti volumen illud dicens quare scripsisti in eo adnuntians festinus veniet rex Babylonis et vastabit terram hanc et cessare faciet ex illa hominem et iumentum
JER|36|30|propterea haec dicit Dominus contra Ioachim regem Iuda non erit ex eo qui sedeat super solium David et cadaver eius proicietur ad aestum per diem et ad gelu per noctem
JER|36|31|et visitabo contra eum et contra semen eius et contra servos eius iniquitates suas et adducam super eos et super habitatores Hierusalem et super viros Iuda omne malum quod locutus sum ad eos et non audierunt
JER|36|32|Hieremias autem tulit volumen aliud et dedit illud Baruch filio Neriae scribae qui scripsit in eo ex ore Hieremiae omnes sermones libri quem conbuserat Ioachim rex Iuda igni et insuper additi sunt sermones multo plures quam ante fuerant
JER|37|1|et regnavit rex Sedecias filius Iosiae pro Iechonia filio Ioachim quem constituit regem Nabuchodonosor rex Babylonis in terra Iuda
JER|37|2|et non oboedivit ipse et servi eius et populus terrae verbis Domini quae locutus est in manu Hieremiae prophetae
JER|37|3|et misit rex Sedecias Iuchal filium Selemiae et Sophoniam filium Maasiae sacerdotem ad Hieremiam prophetam dicens ora pro nobis Dominum Deum nostrum
JER|37|4|Hieremias autem libere ambulabat in medio populi non enim miserant eum in custodiam carceris igitur exercitus Pharao egressus est Aegyptum et audientes Chaldei qui obsidebant Hierusalem huiuscemodi nuntium recesserunt ab Hierusalem
JER|37|5|et factum est verbum Domini ad Hieremiam prophetam dicens
JER|37|6|haec dicit Dominus Deus Israhel sic dicetis regi Iuda qui misit vos ad me ad interrogandum ecce exercitus Pharaonis qui egressus est vobis in auxilium revertetur in terram suam in Aegyptum
JER|37|7|et redient Chaldei et bellabunt contra civitatem hanc et capient eam et incendent igni
JER|37|8|haec dicit Dominus nolite decipere animas vestras dicentes euntes abibunt et recedent a nobis Chaldei quia non abibunt
JER|37|9|sed et si percusseritis omnem exercitum Chaldeorum qui proeliantur adversum vos et derelicti fuerint ex eis aliqui vulnerati singuli de tentorio suo consurgent et incendent civitatem hanc igni
JER|37|10|ergo cum recessisset exercitus Chaldeorum ab Hierusalem propter exercitum Pharaonis
JER|37|11|egressus est Hieremias de Hierusalem ut iret in terram Beniamin et divideret ibi possessionem in conspectu civium
JER|37|12|cumque pervenisset ad portam Beniamin erat ibi custos portae per vices nomine Hierias filius Selemiae filii Ananiae et adprehendit Hieremiam prophetam dicens ad Chaldeos profugis
JER|37|13|et respondit Hieremias falsum est non fugio ad Chaldeos et non audivit eum sed conprehendit Hierias Hieremiam et adduxit eum ad principes
JER|37|14|quam ob rem irati principes contra Hieremiam caesum eum miserunt in carcerem qui erat in domo Ionathan scribae ipse enim praepositus erat super carcerem
JER|37|15|itaque ingressus est Hieremias in domum laci et in ergastula et sedit ibi Hieremias diebus multis
JER|37|16|mittens autem rex Sedecias tulit eum et interrogavit in domo sua abscondite et dixit putasne est sermo a Domino et dixit Hieremias est et ait in manu regis Babylonis traderis
JER|37|17|et dixit Hieremias ad regem Sedeciam quid peccavi tibi et servis tuis et populo tuo quia misisti me in domum carceris
JER|37|18|ubi sunt prophetae vestri qui prophetabant vobis et dicebant non veniet rex Babylonis super vos et super terram hanc
JER|37|19|nunc ergo audi obsecro domine mi rex valeat deprecatio mea in conspectu tuo et ne me remittas in domum Ionathan scribae ne moriar ibi
JER|37|20|praecepit ergo rex Sedecias ut traderetur Hieremias in vestibulo carceris et daretur ei torta panis cotidie excepto pulmento donec consumerentur omnes panes de civitate et mansit Hieremias in vestibulo carceris
JER|38|1|audivit autem Saphatias filius Matthan et Gedelias filius Phassur et Iuchal filius Selemiae et Phassur filius Melchiae sermones quos Hieremias loquebatur ad omnem populum dicens
JER|38|2|haec dicit Dominus quicumque manserit in civitate hac morietur gladio et fame et peste qui autem profugerit ad Chaldeos vivet et erit anima eius sospes et vivens
JER|38|3|haec dicit Dominus tradenda tradetur civitas haec in manu exercitus regis Babylonis et capiet eam
JER|38|4|et dixerunt principes regi rogamus ut occidatur homo iste de industria enim dissolvit manus virorum bellantium qui remanserunt in civitate hac et manus universi populi loquens ad eos iuxta verba haec siquidem homo hic non quaerit pacem populi huius sed malum
JER|38|5|et dixit rex Sedecias ecce ipse in manibus vestris est nec enim fas est regem vobis quicquam negare
JER|38|6|tulerunt ergo Hieremiam et proiecerunt eum in lacu Melchiae filii Ammelech qui erat in vestibulo carceris et submiserunt Hieremiam in funibus et in lacum non erat aqua sed lutum descendit itaque Hieremias in caenum
JER|38|7|audivit autem Abdemelech Aethiops vir eunuchus qui erat in domo regis quod misissent Hieremiam in lacum porro rex sedebat in porta Beniamin
JER|38|8|et egressus est Abdemelech de domo regis et locutus est ad regem dicens
JER|38|9|domine mi rex malefecerunt viri isti omnia quaecumque perpetrarunt contra Hieremiam prophetam mittentes eum in lacum ut moriatur ibi fame non sunt enim panes ultra in civitate
JER|38|10|praecepit itaque rex Abdemelech Aethiopi dicens tolle tecum hinc triginta viros et leva Hieremiam prophetam de lacu antequam moriatur
JER|38|11|adsumptis ergo Abdemelech secum viris ingressus est domum regis quae erat sub cellario et tulit inde veteres pannos et antiqua quae conputruerant et submisit ea ad Hieremiam in lacum per funiculos
JER|38|12|dixitque Abdemelech Aethiops ad Hieremiam pone veteres pannos et haec scissa et putrida sub cubitu manuum tuarum et subter funes fecit ergo Hieremias sic
JER|38|13|et extraxerunt Hieremiam funibus et eduxerunt eum de lacu mansit autem Hieremias in vestibulo carceris
JER|38|14|et misit rex Sedecias et tulit ad se Hieremiam prophetam ad ostium tertium quod erat in domo Domini et dixit rex ad Hieremiam interrogo ego te sermonem ne abscondas a me aliquid
JER|38|15|dixit autem Hieremias ad Sedeciam si adnuntiavero tibi numquid non interficies me et si consilium tibi dedero non me audies
JER|38|16|iuravit ergo rex Sedecias Hieremiae clam dicens vivit Dominus qui fecit nobis animam hanc si occidero te et si tradidero te in manu virorum istorum qui quaerunt animam tuam
JER|38|17|et dixit Hieremias ad Sedeciam haec dicit Dominus exercituum Deus Israhel si profectus exieris ad principes regis Babylonis vivet anima tua et civitas haec non succendetur igni et salvus eris tu et domus tua
JER|38|18|si autem non exieris ad principes regis Babylonis tradetur civitas haec in manu Chaldeorum et succendent eam igni et tu non effugies de manu eorum
JER|38|19|et dixit rex Sedecias ad Hieremiam sollicitus sum propter Iudaeos qui transfugerunt ad Chaldeos ne forte tradar in manus eorum et inludant mihi
JER|38|20|respondit autem Hieremias non te tradent audi quaeso vocem Domini quam ego loquor ad te et bene tibi erit et vivet anima tua
JER|38|21|quod si nolueris egredi iste est sermo quem ostendit mihi Dominus
JER|38|22|ecce omnes mulieres quae remanserunt in domo regis Iuda educentur ad principes regis Babylonis et ipsae dicent seduxerunt te et praevaluerunt adversum te viri pacifici tui demerserunt in caeno et lubrico pedes tuos et recesserunt a te
JER|38|23|et omnes uxores tuae et filii tui educentur ad Chaldeos et non effugies manus eorum sed in manu regis Babylonis capieris et civitatem hanc conburet igni
JER|38|24|dixit ergo Sedecias ad Hieremiam nullus sciat verba haec et non morieris
JER|38|25|si autem audierint principes quia locutus sum tecum et venerint ad te et dixerint tibi indica nobis quid locutus sis cum rege ne celes nos et non te interficiemus et quid locutus est tecum rex
JER|38|26|dices ad eos prostravi ego preces meas coram rege ne me reduci iuberet in domum Ionathan et ibi morerer
JER|38|27|venerunt ergo omnes principes ad Hieremiam et interrogaverunt eum et locutus est eis iuxta omnia verba quae praeceperat ei rex et cessaverunt ab eo nihil enim fuerat auditum
JER|38|28|mansit vero Hieremias in vestibulo carceris usque ad diem quo capta est Hierusalem et factum est ut caperetur Hierusalem
JER|39|1|anno nono Sedeciae regis Iuda mense decimo venit Nabuchodonosor rex Babylonis et omnis exercitus eius ad Hierusalem et obsidebant eam
JER|39|2|undecimo autem anno Sedeciae mense quarto quinta mensis aperta est civitas
JER|39|3|et ingressi sunt omnes principes regis Babylonis et sederunt in porta media Neregel Sereser Semegar Nabu Sarsachim Rabsares Neregel Sereser Rebmag et omnes reliqui principes regis Babylonis
JER|39|4|cumque vidisset eos Sedecias rex Iuda et omnes viri bellatores fugerunt et egressi sunt nocte de civitate per viam horti regis et per portam quae erat inter duos muros et egressi sunt ad viam deserti
JER|39|5|persecutus est autem eos exercitus Chaldeorum et conprehenderunt Sedeciam in campo solitudinis hiericuntinae et captum adduxerunt ad Nabuchodonosor regem Babylonis in Reblatha quae est in terra Emath et locutus est ad eum iudicia
JER|39|6|et occidit rex Babylonis filios Sedeciae in Reblatha in oculis eius et omnes nobiles Iuda occidit rex Babylonis
JER|39|7|oculos quoque Sedeciae eruit et vinxit eum conpedibus ut duceretur in Babylonem
JER|39|8|domum quoque regis et domum vulgi succenderunt Chaldei igni et murum Hierusalem subverterunt
JER|39|9|et reliquias populi quae remanserunt in civitate et perfugas qui transfugerant ad eum et superfluos vulgi qui remanserant transtulit Nabuzardan magister militum in Babylonem
JER|39|10|et de plebe pauperum qui nihil penitus habebant dimisit Nabuzardan magister militum in terra Iuda et dedit eis vineas et cisternas in die illa
JER|39|11|praeceperat autem Nabuchodonosor rex Babylonis de Hieremia Nabuzardan magistro militiae dicens
JER|39|12|tolle illum et pone super eum oculos tuos nihilque ei mali facias sed ut voluerit sic facies ei
JER|39|13|misit ergo Nabuzardan princeps militiae et Nabu et Sesban et Rabsares et Neregel et Sereser et Rebmag et omnes optimates regis Babylonis
JER|39|14|miserunt et tulerunt Hieremiam de vestibulo carceris et tradiderunt eum Godoliae filio Ahicam filii Saphan ut intraret domum et habitaret in populo
JER|39|15|ad Hieremiam autem factus fuerat sermo Domini cum clausus esset in vestibulo carceris dicens
JER|39|16|vade et dic Abdemelech Aethiopi dicens haec dicit Dominus exercituum Deus Israhel ecce ego inducam sermones meos super civitatem hanc in malum et non in bonum et erunt in conspectu tuo in die illa
JER|39|17|et liberabo te in die illa ait Dominus et non traderis in manus virorum quos tu formidas
JER|39|18|sed eruens liberabo te et gladio non cades sed erit tibi anima tua in salutem quia in me habuisti fiduciam ait Dominus
JER|40|1|sermo qui factus est ad Hieremiam a Domino postquam dimissus est a Nabuzardan magistro militiae de Rama quando tulit eum vinctum catenis in medio omnium qui migrabant de Hierusalem et Iuda et ducebantur in Babylonem
JER|40|2|tollens ergo princeps militiae Hieremiam dixit ad eum Dominus Deus tuus locutus est malum hoc super locum istum
JER|40|3|et adduxit et fecit Dominus sicut locutus est quia peccastis Domino et non audistis vocem eius et factus est vobis sermo hic
JER|40|4|nunc ergo ecce solvi te hodie de catenis quae sunt in manibus tuis si placet tibi ut venias mecum in Babylonem veni et ponam oculos meos super te si autem displicet tibi venire mecum in Babylonem reside ecce omnis terra in conspectu tuo quod elegeris et quo placuerit tibi ut vadas illuc perge
JER|40|5|et mecum noli venire sed habita apud Godoliam filium Ahicam filii Saphan quem praeposuit rex Babylonis civitatibus Iudaeae habita ergo cum eo in medio populi vel quocumque placuerit tibi ut vadas vade dedit quoque ei magister militiae cibaria et munuscula et dimisit eum
JER|40|6|venit autem Hieremias ad Godoliam filium Ahicam in Masphat et habitavit cum eo in medio populi qui relictus fuerat in terra
JER|40|7|cum ergo audissent omnes principes exercitus qui dispersi fuerant per regiones ipsi et socii eorum quod praefecisset rex Babylonis Godoliam filium Ahicam terrae et quod commendasset ei viros et mulieres et parvulos et de pauperibus terrae qui non fuerant translati in Babylonem
JER|40|8|venerunt ad Godoliam in Masphat et Ismahel filius Nathaniae et Iohanan et Ionathan filii Caree et Sareas filius Thenoemeth et filii Offi qui erat de Nethophathi et Iezonias filius Maachathi ipsi et viri eorum
JER|40|9|et iuravit eis Godolias filius Ahicam filii Saphan et comitibus eorum dicens nolite timere servire Chaldeis habitate in terra et servite regi Babylonis et bene erit vobis
JER|40|10|ecce ego habito in Masphat ut respondeam praecepto Chaldeorum qui mittuntur ad nos vos autem colligite vindemiam et messem et oleum et condite in vasis vestris et manete in urbibus vestris quas tenetis
JER|40|11|sed et omnes Iudaei qui erant in Moab et in filiis Ammon et in Idumea et in universis regionibus audito quod dedisset rex Babylonis reliquias in Iudaeam et quod praeposuisset super eos Godoliam filium Ahicam filii Saphan
JER|40|12|reversi sunt inquam omnes Iudaei de universis locis ad quae profugerant et venerunt in terram Iuda ad Godoliam in Masphat et collegerunt vinum et messem multam nimis
JER|40|13|Iohanan autem filius Caree et omnes principes exercitus qui dispersi erant in regionibus venerunt ad Godoliam in Masphat
JER|40|14|et dixerunt ei scito quia Baalis rex filiorum Ammon misit Ismahel filium Nathaniae percutere animam tuam et non credidit eis Godolias filius Ahicam
JER|40|15|Iohanan vero filius Caree dixit ad Godoliam seorsum in Masphat loquens ibo et percutiam Ismahel filium Nathaniae nullo sciente ne interficiat animam tuam et dissipentur omnes Iudaei qui congregati sunt ad te et peribunt reliquiae Iuda
JER|40|16|et ait Godolias filius Ahicam ad Iohanan filium Caree noli facere verbum hoc falsum enim tu loqueris de Ismahel
JER|41|1|et factum est in mense septimo venit Ismahel filius Nathaniae filii Elisama de semine regali et optimates regis et decem viri cum eo ad Godoliam filium Ahicam in Masphat et comederunt ibi panes simul in Masphat
JER|41|2|surrexit autem Ismahel filius Nathaniae et decem viri qui erant cum eo et percusserunt Godoliam filium Ahicam filii Saphan gladio et interfecerunt eum quem praefecerat rex Babylonis terrae
JER|41|3|omnes quoque Iudaeos qui erant cum Godolia in Masphat et Chaldeos qui repperti sunt ibi et viros bellatores percussit Ismahel
JER|41|4|secundo autem die postquam occiderat Godoliam nullo adhuc sciente
JER|41|5|venerunt viri de Sychem et de Silo et de Samaria octoginta viri rasi barbam et scissis vestibus et squalentes munera et tus habebant in manu ut offerrent in domo Domini
JER|41|6|egressus ergo Ismahel filius Nathaniae in occursum eorum de Masphat incedens et plorans ibat cum autem occurrisset eis dixit ad eos venite ad Godoliam filium Ahicam
JER|41|7|qui cum venissent ad medium civitatis interfecit eos Ismahel filius Nathaniae circa medium laci ipse et viri qui erant cum eo
JER|41|8|decem autem viri repperti sunt inter eos qui dixerunt ad Ismahel noli occidere nos quia habemus thesauros in agro frumenti et hordei et olei et mellis et cessavit et non interfecit eos cum fratribus suis
JER|41|9|lacus autem in quem proiecerat Ismahel omnia cadavera virorum quos percussit propter Godoliam ipse est quem fecit rex Asa propter Baasa regem Israhel ipsum replevit Ismahel filius Nathaniae occisis
JER|41|10|et captivas duxit Ismahel omnes reliquias populi qui erant in Masphat filias regis et universum populum qui remanserat in Masphat quos commendarat Nabuzardan princeps militiae Godoliae filio Ahicam et cepit eos Ismahel filius Nathaniae et abiit ut transiret ad filios Ammon
JER|41|11|audivit autem Iohanan filius Caree et omnes principes bellatorum qui erant cum eo omne malum quod fecerat Ismahel filius Nathaniae
JER|41|12|et adsumptis universis viris profecti sunt ut bellarent adversum Ismahel filium Nathaniae et invenerunt eum ad aquas Multas quae sunt in Gabaon
JER|41|13|cumque vidisset omnis populus qui erat cum Ismahel Iohanan filium Caree et universos principes bellatorum qui erant cum eo laetati sunt
JER|41|14|et reversus est omnis populus quem ceperat Ismahel in Masphat reversusque abiit ad Iohanan filium Caree
JER|41|15|Ismahel autem filius Nathaniae fugit cum octo viris a facie Iohanan et abiit ad filios Ammon
JER|41|16|tulit ergo Iohanan filius Caree et omnes principes bellatorum qui erant cum eo universas reliquias vulgi quas reduxerat ab Ismahel filio Nathaniae de Masphat postquam percussit Godoliam filium Ahicam fortes viros ad proelium et mulieres et pueros et eunuchos quos reduxerat de Gabaon
JER|41|17|et abierunt et sederunt peregrinantes in Chamaam quae est iuxta Bethleem ut pergerent et introirent Aegyptum
JER|41|18|a facie Chaldeorum timebant enim eos quia percusserat Ismahel filius Nathaniae Godoliam filium Ahicam quem praeposuerat rex Babylonis in terra Iuda
JER|42|1|et accesserunt omnes principes bellatorum et Iohanan filius Caree et Iezonias filius Osaiae et reliquum vulgus a parvo usque ad magnum
JER|42|2|dixeruntque ad Hieremiam prophetam cadat oratio nostra in conspectu tuo et ora pro nobis ad Dominum Deum tuum pro universis reliquiis istis quia derelicti sumus pauci de pluribus sicut oculi tui nos intuentur
JER|42|3|et adnuntiet nobis Dominus Deus tuus viam per quam pergamus et verbum quod faciamus
JER|42|4|dixit autem ad eos Hieremias propheta audivi ecce ego oro ad Dominum Deum vestrum secundum verba vestra omne verbum quodcumque responderit mihi indicabo vobis nec celabo vos quicquam
JER|42|5|et illi dixerunt ad Hieremiam sit Dominus inter nos testis veritatis et fidei si non iuxta omne verbum in quo miserit te Dominus Deus tuus ad nos sic faciemus
JER|42|6|sive bonum est sive malum voci Domini Dei nostri ad quem mittimus te oboediemus ut bene sit nobis cum audierimus vocem Domini Dei nostri
JER|42|7|cum autem conpleti essent decem dies factum est verbum Domini ad Hieremiam
JER|42|8|vocavitque Iohanan filium Caree et omnes principes bellatorum qui erant cum eo et universum populum a minimo usque ad magnum
JER|42|9|et dixit ad eos haec dicit Dominus Deus Israhel ad quem misistis me ut prosternerem preces vestras in conspectu eius
JER|42|10|si quiescentes manseritis in terra hac aedificabo vos et non destruam plantabo et non evellam iam enim placatus sum super malo quod feci vobis
JER|42|11|nolite timere a facie regis Babylonis quem vos pavidi formidatis nolite eum metuere dicit Dominus quia vobiscum sum ego ut salvos faciam vos et eruam de manu eius
JER|42|12|et dabo vobis misericordiam et miserebor vestri et habitare vos faciam in terra vestra
JER|42|13|si autem dixeritis vos non habitabimus in terra ista nec audiemus vocem Domini Dei nostri
JER|42|14|dicentes nequaquam sed ad terram Aegypti pergemus ubi non videbimus bellum et clangorem tubae non audiemus et famem non sustinebimus et ibi habitabimus
JER|42|15|propter hoc nunc audite verbum Domini reliquiae Iuda haec dicit Dominus exercituum Deus Israhel si posueritis faciem vestram ut ingrediamini Aegyptum et intraveritis ut ibi habitetis
JER|42|16|gladium quem vos formidatis ibi conprehendet vos in terra Aegypti et fames pro qua estis solliciti adherebit vobis in Aegypto et ibi moriemini
JER|42|17|omnesque viri qui posuerint faciem suam ut ingrediantur Aegyptum et habitent ibi morientur gladio et fame et peste nullus de eis remanebit nec effugient a facie mali quod ego adferam super eos
JER|42|18|quia haec dicit Dominus exercituum Deus Israhel sicut conflatus est furor meus et indignatio mea super habitatores Hierusalem sic conflabitur indignatio mea super vos cum ingressi fueritis Aegyptum et eritis in iusiurandum et in stuporem et in maledictum et in obprobrium et nequaquam ultra videbitis locum istum
JER|42|19|verbum Domini super vos reliquiae Iuda nolite intrare Aegyptum scientes scietis quia obtestatus sum vobis hodie
JER|42|20|quia decepistis animas vestras vos enim misistis me ad Dominum Deum nostrum dicentes ora pro nobis ad Dominum Deum nostrum et iuxta omnia quaecumque dixerit tibi Dominus Deus noster sic adnuntia nobis et faciemus
JER|42|21|et adnuntiavi vobis hodie et non audistis vocem Domini Dei vestri super universis pro quibus misit me ad vos
JER|42|22|nunc ergo scientes scietis quia gladio et fame et peste moriemini in loco ad quem voluistis intrare ut habitaretis ibi
JER|43|1|factum est autem cum conplesset Hieremias loquens ad populum universos sermones Domini Dei eorum pro quibus miserat eum Dominus Deus eorum ad illos omnia verba haec
JER|43|2|dixit Azarias filius Osaiae et Iohanan filius Caree et omnes viri superbi dicentes ad Hieremiam mendacium tu loqueris non misit te Dominus Deus noster dicens ne ingrediamini Aegyptum ut habitetis illuc
JER|43|3|sed Baruch filius Neriae incitat te adversum nos ut tradat nos in manibus Chaldeorum ut interficiat nos et transduci faciat in Babylonem
JER|43|4|et non audivit Iohanan filius Caree et omnes principes bellatorum et universus populus vocem Domini ut maneret in terra Iuda
JER|43|5|sed tollens Iohanan filius Caree et universi principes bellatorum universos reliquiarum Iuda qui reversi fuerant de cunctis gentibus ad quas fuerant ante dispersi ut habitarent in terra Iuda
JER|43|6|viros et mulieres et parvulos et filias regis et omnem animam quam reliquerat Nabuzardan princeps militiae cum Godolia filio Ahicam filii Saphan et Hieremiam prophetam et Baruch filium Neriae
JER|43|7|et ingressi sunt terram Aegypti quia non oboedierunt voci Domini et venerunt usque ad Tafnas
JER|43|8|et factus est sermo Domini ad Hieremiam in Tafnis dicens
JER|43|9|sume in manu tua lapides grandes et absconde eos in crypta quae est sub muro latericio in porta domus Pharaonis in Tafnis cernentibus viris iudaeis
JER|43|10|et dices ad eos haec dicit Dominus exercituum Deus Israhel ecce ego mittam et adsumam Nabuchodonosor regem Babylonis servum meum et ponam thronum eius super lapides istos quos abscondi et statuet solium suum super eos
JER|43|11|veniensque percutiet terram Aegypti quos in morte in morte et quos in captivitate in captivitate et quos in gladio in gladio
JER|43|12|et succendet ignem in delubris deorum Aegypti et conburet ea et captivos ducet illos et amicietur terra Aegypti sicut amicitur pastor pallio suo et egredietur inde in pace
JER|43|13|et conteret statuas domus Solis quae sunt in terra Aegypti et delubra deorum Aegypti conburet igni
JER|44|1|verbum quod factum est ad Hieremiam ad omnes Iudaeos qui habitant in terra Aegypti habitantes in Magdolo et in Tafnis et in Memphis et in terra Fatures dicens
JER|44|2|haec dicit Dominus exercituum Deus Israhel vos vidistis omne malum istud quod adduxi super Hierusalem et super omnes urbes Iuda et ecce sunt desertae hodie et non est in eis habitator
JER|44|3|propter malitiam quam fecerunt ut me ad iracundiam provocarent et irent et sacrificarent et colerent deos alienos quos nesciebant et illi et vos et patres vestri
JER|44|4|et misi ad vos omnes servos meos prophetas de nocte consurgens mittensque et dicens nolite facere verbum abominationis huius quam odi
JER|44|5|et non audierunt nec inclinaverunt aurem suam ut converterentur a malis suis et non sacrificarent diis alienis
JER|44|6|et conflata est indignatio mea et furor meus et succensa est in civitatibus Iuda et in plateis Hierusalem et versae sunt in solitudinem et vastitatem secundum diem hanc
JER|44|7|et nunc haec dicit Dominus exercituum Deus Israhel quare vos facitis malum grande contra animas vestras ut intereat ex vobis vir et mulier parvulus et lactans de medio Iudae nec relinquatur vobis quicquam residuum
JER|44|8|provocantes me in operibus manuum vestrarum sacrificando diis alienis in terra Aegypti in quam ingressi estis ut habitetis ibi et dispereatis et sitis in maledictionem et in obprobrium cunctis gentibus terrae
JER|44|9|numquid obliti estis mala patrum vestrorum et mala regum Iuda et mala uxorum eius et mala vestra et mala uxorum vestrarum quae fecerunt in terra Iuda et in regionibus Hierusalem
JER|44|10|non sunt mundati usque ad diem hanc et non timuerunt et non ambulaverunt in lege et in praeceptis meis quae dedi coram vobis et coram patribus vestris
JER|44|11|ideo haec dicit Dominus exercituum Deus Israhel ecce ego pono faciem meam in vobis in malum et disperdam omnem Iudam
JER|44|12|et adsumam reliquias Iudae qui posuerunt facies suas ut ingrederentur terram Aegypti et habitarent ibi et consumentur omnes in terra Aegypti cadent in gladio et in fame consumentur a minimo usque ad maximum in gladio et in fame morientur et erunt in iusiurandum et in miraculum et in maledictionem et in obprobrium
JER|44|13|et visitabo habitatores terrae Aegypti sicut visitavi super Hierusalem in gladio et in fame et in peste
JER|44|14|et non erit qui effugiat et sit residuus de reliquiis Iudaeorum qui vadunt ut peregrinentur in terra Aegypti et revertantur in terram Iuda ad quam ipsi elevant animas suas ut revertantur et habitent ibi non revertentur nisi qui fugerint
JER|44|15|responderunt autem Hieremiae omnes viri scientes quod sacrificarent uxores eorum diis alienis et universae mulieres quarum stabat multitudo grandis et omnis populus habitantium in terra Aegypti in Fatures dicens
JER|44|16|sermonem quem locutus es ad nos in nomine Domini non audiemus ex te
JER|44|17|sed facientes faciemus omne verbum quod egreditur de ore nostro ut sacrificemus Reginae caeli et libemus ei libamina sicut fecimus nos et patres nostri reges nostri et principes nostri in urbibus Iuda et in plateis Hierusalem et saturati sumus panibus et bene nobis erat malumque non vidimus
JER|44|18|ex eo autem quo cessavimus sacrificare Reginae caeli et libare ei libamina indigemus omnibus et gladio et fame consumpti sumus
JER|44|19|quod si nos sacrificamus Reginae caeli et libamus ei libamina numquid sine viris nostris fecimus ei placentas ad colendum eam et liba libandi
JER|44|20|et dixit Hieremias ad omnem populum adversum viros et adversum mulieres et adversum universam plebem qui responderant ei verbum dicens
JER|44|21|numquid non sacrificium quod sacrificastis in civitatibus Iuda et in plateis Hierusalem vos et patres vestri reges vestri et principes vestri et populus terrae horum recordatus est Dominus et ascendit super cor eius
JER|44|22|et non poterat Dominus ultra portare propter malitiam studiorum vestrorum et propter abominationes quas fecistis et facta est terra vestra in desolationem et in stuporem et in maledictum eo quod non sit habitator sicut est dies haec
JER|44|23|propterea quod sacrificaveritis idolis et peccaveritis Domino et non audieritis vocem Domini et in lege et in praeceptis et in testimoniis eius non ambulaveritis idcirco evenerunt vobis mala haec sicut est dies haec
JER|44|24|dixit autem Hieremias ad omnem populum et ad universas mulieres audite verbum Domini omnis Iuda qui estis in terra Aegypti
JER|44|25|haec inquit Dominus exercituum Deus Israhel dicens vos et uxores vestrae locuti estis ore vestro et manibus vestris implestis dicentes faciamus vota nostra quae vovimus ut sacrificemus Reginae caeli et libemus ei libamina implestis vota vestra et opere perpetrastis ea
JER|44|26|ideo audite verbum Domini omnis Iuda qui habitatis in terra Aegypti ecce ego iuravi in nomine meo magno ait Dominus quia nequaquam ultra nomen meum vocabitur ex ore omnis viri iudaei dicentis vivit Dominus Deus in omni terra Aegypti
JER|44|27|ecce ego vigilabo super eos in malum et non in bonum et consumentur omnes viri Iuda qui sunt in terra Aegypti gladio et fame donec penitus consumantur
JER|44|28|et qui fugerint gladium revertentur de terra Aegypti in terram Iuda viri pauci et scient omnes reliquiae Iuda ingredientium terram Aegypti ut habitent ibi cuius sermo conpleatur meus an illorum
JER|44|29|et hoc vobis signum ait Dominus quod visitem ego super vos in loco isto ut sciatis quia vere conplebuntur sermones mei contra vos in malum
JER|44|30|haec dicit Dominus ecce ego tradam Pharaonem Efree regem Aegypti in manu inimicorum eius et in manu quaerentium animam illius sicut tradidi Sedeciam regem Iuda in manu Nabuchodonosor regis Babylonis inimici sui et quaerentis animam eius
JER|45|1|verbum quod locutus est Hieremias propheta ad Baruch filium Neri cum scripsisset verba haec in libro de ore Hieremiae anno quarto Ioachim filii Iosiae regis Iuda dicens
JER|45|2|haec dicit Dominus Deus Israhel ad te Baruch
JER|45|3|dixisti vae misero mihi quoniam addidit Dominus dolorem dolori meo laboravi in gemitu meo et requiem non inveni
JER|45|4|haec dices ad eum sic dicit Dominus ecce quos aedificavi ego destruo et quos plantavi ego evello et universam terram hanc
JER|45|5|et tu quaeris tibi grandia noli quaerere quia ecce ego adducam malum super omnem carnem ait Dominus et dabo tibi animam tuam in salutem in omnibus locis ad quaecumque perrexeris
JER|46|1|quod factum est verbum Domini ad Hieremiam prophetam contra gentes
JER|46|2|ad Aegyptum adversum exercitum Pharaonis Nechao regis Aegypti qui erat iuxta flumen Eufraten in Charchamis quem percussit Nabuchodonosor rex Babylonis in quarto anno Ioachim filii Iosiae regis Iuda
JER|46|3|praeparate scutum et clypeum et procedite ad bellum
JER|46|4|iungite equos et ascendite equites state in galeis polite lanceas induite vos loricis
JER|46|5|quid igitur vidi ipsos pavidos et terga vertentes fortes eorum caesos fugerunt conciti nec respexerunt terror undique ait Dominus
JER|46|6|non fugiat velox nec salvari se putet fortis ad aquilonem iuxta flumen Eufraten victi sunt et ruerunt
JER|46|7|quis est iste qui quasi flumen ascendit et veluti fluviorum intumescunt gurgites eius
JER|46|8|Aegyptus fluminis instar ascendet et velut flumina movebuntur fluctus eius et dicet ascendens operiam terram perdam civitatem et habitatores eius
JER|46|9|ascendite equos et exultate in curribus et procedant fortes Aethiopia et Lybies tenentes scutum et Lydii arripientes et iacientes sagittas
JER|46|10|dies autem ille Domini Dei exercituum dies ultionis ut sumat vindictam de inimicis suis devorabit gladius et saturabitur et inebriabitur sanguine eorum victima enim Domini exercituum in terra aquilonis iuxta flumen Eufraten
JER|46|11|ascende in Galaad et tolle resinam virgo filia Aegypti frustra multiplicas medicamina sanitas non erit tibi
JER|46|12|audierunt gentes ignominiam tuam et ululatus tuus replevit terram quia fortis inpegit in fortem ambo pariter conciderunt
JER|46|13|verbum quod locutus est Dominus ad Hieremiam prophetam super eo quod venturus esset Nabuchodonosor rex Babylonis et percussurus terram Aegypti
JER|46|14|adnuntiate Aegypto et auditum facite Magdolo et resonet in Memphis et in Tafnis dicite sta et praepara te quia devoravit gladius ea quae per circuitum tuum sunt
JER|46|15|quare conputruit fortis tuus non stetit quoniam Dominus subvertit eum
JER|46|16|multiplicavit ruentes ceciditque vir ad proximum suum et dicent surge et revertamur ad populum nostrum et ad terram nativitatis nostrae a facie gladii columbae
JER|46|17|vocate nomen Pharao regis Aegypti Tumultum adduxit tempus
JER|46|18|vivo ego inquit Rex Dominus exercituum nomen eius quoniam sicut Thabor in montibus et sicut Carmelus in mari veniet
JER|46|19|vasa transmigrationis fac tibi habitatrix filia Aegypti quia Memphis in solitudinem erit et deseretur inhabitabilis
JER|46|20|vitula eligans atque formonsa Aegyptus stimulator ab aquilone veniet ei
JER|46|21|mercennarii quoque eius qui versabantur in medio eius quasi vituli saginati versi sunt et fugerunt simul nec stare potuerunt quia dies interfectionis eorum venit super eos tempus visitationis eorum
JER|46|22|vox eius quasi aeris sonabit quoniam cum exercitu properabunt et cum securibus venient ei quasi ligna caedentes
JER|46|23|succiderunt saltum eius ait Dominus qui supputari non potest multiplicati sunt super lucustas et non est eis numerus
JER|46|24|confusa est filia Aegypti et tradita in manu populi aquilonis
JER|46|25|dixit Dominus exercituum Deus Israhel ecce ego visitabo super tumultum Alexandriae et super Pharao et super Aegyptum et super deos eius et super reges eius et super Pharao et super eos qui confidunt in eo
JER|46|26|et dabo eos in manu quaerentium animam eorum et in manu Nabuchodonosor regis Babylonis et in manu servorum eius et post haec habitabitur sicut diebus pristinis ait Dominus
JER|46|27|et tu ne timeas serve meus Iacob et ne paveas Israhel quia ecce ego salvum te faciam de longinquo et semen tuum de terra captivitatis suae et revertetur Iacob et quiescet et prosperabitur et non erit qui exterreat eum
JER|46|28|et tu noli timere serve meus Iacob ait Dominus quia tecum ego sum quia consumam ego cunctas gentes ad quas eieci te te vero non consumam sed castigabo te in iudicio nec quasi innocenti parcam tibi
JER|47|1|quod factum est verbum Domini ad Hieremiam prophetam contra Palestinos antequam percuteret Pharao Gazam
JER|47|2|haec dicit Dominus ecce aquae ascendunt ab aquilone et erunt quasi torrens inundans et operient terram et plenitudinem eius urbem et habitatores eius clamabunt homines et ululabit omnis habitator terrae
JER|47|3|ab strepitu pompae armorum et bellatorum eius a commotione quadrigarum eius et multitudine rotarum illius non respexerunt patres filios manibus dissolutis
JER|47|4|pro adventu diei in quo vastabuntur omnes Philisthim et dissipabitur Tyrus et Sidon cum omnibus reliquis auxiliis suis depopulatus est enim Dominus Palestinos reliquias insulae Cappadociae
JER|47|5|venit calvitium super Gazam conticuit Ascalon et reliquiae vallis earum usquequo concideris
JER|47|6|o mucro Domini usquequo non quiescis ingredere in vaginam tuam refrigerare et sile
JER|47|7|quomodo quiescet cum Dominus praeceperit ei adversus Ascalonem et adversus maritimas eius regiones ibique condixerit illi
JER|48|1|ad Moab haec dicit Dominus exercituum Deus Israhel vae super Nabo quoniam vastata est et confusa capta est Cariathaim confusa est fortis et tremuit
JER|48|2|non est ultra exultatio in Moab contra Esebon cogitaverunt malum venite et disperdamus eam de gente ergo silens conticesces sequeturque te gladius
JER|48|3|vox clamoris de Oronaim vastitas et contritio magna
JER|48|4|contrita est Moab adnuntiate clamorem parvulis eius
JER|48|5|per ascensum enim Luaith plorans ascendet in fletu quoniam in descensu Oronaim hostes ululatum contritionis audierunt
JER|48|6|fugite salvate animas vestras et eritis quasi myrice in deserto
JER|48|7|pro eo enim quod habuisti fiduciam in munitionibus tuis et in thesauris tuis tu quoque capieris et ibit Chamos in transmigrationem sacerdotes eius et principes eius simul
JER|48|8|et veniet praedo ad omnem urbem et urbs nulla salvabitur et peribit vallis et dissipabuntur campestria quoniam dixit Dominus
JER|48|9|date florem Moab quia floriens egredietur et civitates eius desertae erunt et inhabitabiles
JER|48|10|maledictus qui facit opus Domini fraudulenter et maledictus qui prohibet gladium suum a sanguine
JER|48|11|fertilis fuit Moab ab adulescentia sua et requievit in fecibus suis nec transfusus est de vase in vas et in transmigrationem non abiit idcirco permansit gustus eius in eo et odor eius non est inmutatus
JER|48|12|propterea ecce dies veniunt dicit Dominus et mittam ei ordinatores et stratores laguncularum et sternent eum et vasa eius exhaurient et lagoenas eorum conlident
JER|48|13|et confundetur Moab a Chamos sicut confusa est domus Israhel a Bethel in qua habebat fiduciam
JER|48|14|quomodo dicitis fortes sumus et viri robusti ad proeliandum
JER|48|15|vastata est Moab et civitates illius ascenderunt et electi iuvenes eius descenderunt in occisionem ait Rex Dominus exercituum nomen ei
JER|48|16|prope est interitus Moab ut veniat et malum eius velociter adcurret nimis
JER|48|17|consolamini eum omnes qui estis in circuitu eius et universi qui scitis nomen eius dicite quomodo confracta est virga fortis baculus gloriosus
JER|48|18|descende de gloria et sede in siti habitatio filiae Dibon quoniam vastator Moab ascendet ad te dissipabit munitiones tuas
JER|48|19|in via sta et prospice habitatio Aroer interroga fugientem et eum qui evasit dic quid accidit
JER|48|20|confusus est Moab quoniam victus est ululate et clamate adnuntiate in Arnon quoniam vastata est Moab
JER|48|21|et iudicium venit ad terram campestrem super Helon et super Iaesa et super Mefath
JER|48|22|et super Dibon et super Nabo et super domum Deblathaim
JER|48|23|et super Cariathaim et super Bethgamul et super Bethmaon
JER|48|24|et super Carioth et super Bosra et super omnes civitates terrae Moab quae longe et quae prope sunt
JER|48|25|abscisum est cornu Moab et brachium eius contritum est ait Dominus
JER|48|26|inebriate eum quoniam contra Dominum erectus est et adlidet manum Moab in vomitu suo et erit in derisum etiam ipse
JER|48|27|fuit enim in derisum tibi Israhel quasi inter fures repperisses eum propter verba ergo tua quae adversum illum locutus es captivus duceris
JER|48|28|relinquite civitates et habitate in petra habitatores Moab et estote quasi columba nidificans in summo ore foraminis
JER|48|29|audivimus superbiam Moab superbus est valde sublimitatem eius et arrogantiam et superbiam et altitudinem cordis illius
JER|48|30|ego scio ait Dominus iactantiam eius et quod non sit iuxta eam virtus eius nec iuxta quod poterat conata sit facere
JER|48|31|ideo super Moab heiulabo et ad Moab universam clamabo ad viros muri fictilis lamentantes
JER|48|32|de planctu Iazer plorabo tibi vinea Sobema propagines tuae transierunt mare usque ad mare Iazer pervenerunt super messem tuam et vindemiam tuam praedo inruit
JER|48|33|ablata est laetitia et exultatio de Carmelo et de terra Moab et vinum de torcularibus sustuli nequaquam calcator uvae solitum celeuma cantabit
JER|48|34|de clamore Esebon usque Eleale et Iaesa dederunt vocem suam a Segor usque ad Oronaim vitula conternante aquae quoque Namrim pessimae erunt
JER|48|35|et auferam de Moab ait Dominus offerentem in excelsis et sacrificantem diis eius
JER|48|36|propterea cor meum ad Moab quasi tibiae resonabit et cor meum ad viros muri fictilis dabit sonitum tibiarum quia plus fecit quam potuit idcirco perierunt
JER|48|37|omne enim caput calvitium et omnis barba rasa erit in cunctis manibus conligatio et super omne dorsum cilicium
JER|48|38|super omnia tecta Moab et in plateis eius omnis planctus quia contrivi Moab sicut vas inutile ait Dominus
JER|48|39|quomodo victa est et ululaverunt quomodo deiecit cervicem Moab et confusus est eritque Moab in derisum et in exemplum omnibus in circuitu suo
JER|48|40|haec dicit Dominus ecce quasi aquila evolabit et extendet alas suas ad Moab
JER|48|41|capta est Carioth et munitiones conprehensae sunt et erit cor fortium Moab in die illa sicut cor mulieris parturientis
JER|48|42|et cessabit Moab esse populus quoniam contra Dominum gloriatus est
JER|48|43|pavor et fovea et laqueus super te o habitator Moab ait Dominus
JER|48|44|qui fugit a facie pavoris cadet in foveam et qui conscenderit de fovea capietur laqueo adducam enim super Moab annum visitationis eorum dicit Dominus
JER|48|45|in umbra Esebon steterunt de laqueo fugientes quia ignis egressus est de Esebon et flamma de medio Seon et devorabit partem Moab et verticem filiorum tumultus
JER|48|46|vae tibi Moab peristi popule Chamos quia conprehensi sunt filii tui et filiae tuae in captivitatem
JER|48|47|et convertam captivitatem Moab in novissimis diebus ait Dominus hucusque iudicia Moab
JER|49|1|ad filios Ammon haec dicit Dominus numquid filii non sunt Israhel aut heres non est ei cur igitur hereditate possedit Melchom Gad et populus eius in urbibus eius habitavit
JER|49|2|ideo ecce dies veniunt dicit Dominus et auditum faciam super Rabbath filiorum Ammon fremitum proelii et erit in tumulum dissipata filiaeque eius igni succendentur et possidebit Israhel possessores suos dicit Dominus
JER|49|3|ulula Esebon quoniam vastata est Ahi clamate filiae Rabbath accingite vos ciliciis plangite et circuite per sepes quia Melchom in transmigratione ducetur sacerdotes eius et principes eius simul
JER|49|4|quid gloriaris in vallibus defluxit vallis tua filia delicata quae confidebas in thesauris tuis et dicebas quis veniet ad me
JER|49|5|ecce ego inducam super te terrorem ait Dominus Deus exercituum ab omnibus qui sunt in circuitu tuo et dispergemini singuli a conspectu vestro nec erit qui congreget fugientem
JER|49|6|et post haec reverti faciam captivos filiorum Ammon ait Dominus
JER|49|7|ad Idumeam haec dicit Dominus exercituum numquid non est ultra sapientia in Theman periit consilium a filiis inutilis facta est sapientia eorum
JER|49|8|fugite terga vertite descendite in voragine habitatores Dedan quoniam perditionem Esau adduxi super eum tempus visitationis eius
JER|49|9|si vindemiatores venissent super te non reliquissent racemum si fures in nocte rapuissent quod sufficeret sibi
JER|49|10|ego vero discoperui Esau revelavi abscondita eius et celari non poterit vastatum est semen eius et fratres eius et vicini eius et non erit
JER|49|11|relinque pupillos tuos ego eos faciam vivere et viduae tuae in me sperabunt
JER|49|12|quia haec dicit Dominus ecce quibus non erat iudicium ut biberent calicem bibentes bibent et tu quasi innocens relinqueris non eris innocens sed bibens bibes
JER|49|13|quia per memet ipsum iuravi dicit Dominus quod in solitudinem et in obprobrium et in desertum et in maledictionem erit Bosra et omnes civitates eius erunt in solitudines sempiternas
JER|49|14|auditum audivi a Domino et legatus ad gentes missus est congregamini et venite contra eam et consurgamus in proelium
JER|49|15|ecce enim parvulum dedi te in gentibus contemptibilem inter homines
JER|49|16|arrogantia tua decepit te et superbia cordis tui qui habitas in cavernis petrae et adprehendere niteris altitudinem collis cum exaltaveris quasi aquila nidum tuum inde detraham te dicit Dominus
JER|49|17|et erit Idumea deserta omnis qui transibit per eam stupebit et sibilabit super omnes plagas eius
JER|49|18|sicuti subversa est Sodoma et Gomorra et vicinae eius ait Dominus non habitabit ibi vir et non incolet eam filius hominis
JER|49|19|ecce quasi leo ascendet de superbia Iordanis ad pulchritudinem robustam quia subito currere eum faciam ad illam et quis erit electus quem praeponam ei quis enim similis mei et quis sustinebit me et quis est iste pastor qui resistat vultui meo
JER|49|20|propterea audite consilium Domini quod iniit de Edom et cogitationes eius quas cogitavit de habitatoribus Theman si non deiecerint eos parvuli gregis nisi dissipaverint cum eis habitaculum eorum
JER|49|21|a voce ruinae eorum commota est terra clamor in mari Rubro auditus est vocis eius
JER|49|22|ecce quasi aquila ascendet et evolabit et expandet alas suas super Bosram et erit cor fortium Idumeae in die illa quasi cor mulieris parturientis
JER|49|23|ad Damascum confusa est Emath et Arfad quia auditum pessimum audierunt turbati sunt in mari sollicitudine quiescere non potuit
JER|49|24|dissoluta est Damascus versa in fugam tremor adprehendit eam angustia et dolores tenuerunt eam quasi parturientem
JER|49|25|quomodo dereliquerunt civitatem laudabilem urbem laetitiae
JER|49|26|ideo cadent iuvenes eius in plateis eius et omnes viri proelii conticescent in die illa ait Dominus exercituum
JER|49|27|et succendam ignem in muro Damasci et devorabit moenia Benadad
JER|49|28|ad Cedar et ad regna Asor quae percussit Nabuchodonosor rex Babylonis haec dicit Dominus surgite ascendite ad Cedar et vastate filios orientis
JER|49|29|tabernacula eorum et greges eorum capient pelles eorum et omnia vasa eorum et camelos eorum tollent sibi et vocabunt super eos formidinem in circuitu
JER|49|30|fugite abite vehementer in voraginibus sedete qui habitatis Asor ait Dominus iniit enim contra vos Nabuchodonosor rex Babylonis consilium et cogitavit adversum vos cogitationes
JER|49|31|consurgite et ascendite ad gentem quietam et habitantem confidenter ait Dominus non ostia non vectes ei soli habitant
JER|49|32|et erunt cameli eorum in direptionem et multitudo iumentorum in praedam et dispergam eos in omnem ventum qui sunt adtonsi in comam et ex omni confinio eorum adducam interitum super eos ait Dominus
JER|49|33|et erit Asor in habitaculum draconum deserta usque in aeternum non manebit ibi vir nec incolet eam filius hominis
JER|49|34|quod factum est verbum Domini ad Hieremiam prophetam adversus Aelam in principio regni Sedeciae regis Iuda dicens
JER|49|35|haec dicit Dominus exercituum ecce ego confringam arcum Aelam summam fortitudinem eorum
JER|49|36|et inducam super Aelam quattuor ventos a quattuor plagis caeli et ventilabo eos in omnes ventos istos et non erit gens ad quam non perveniant profugi Aelam
JER|49|37|et pavere faciam Aelam coram inimicis suis et in conspectu quaerentium animam eorum et adducam super eos malum iram furoris mei dicit Dominus et emittam post eos gladium donec consumam eos
JER|49|38|et ponam solium meum in Aelam et perdam inde reges et principes ait Dominus
JER|49|39|in novissimis autem diebus reverti faciam captivos Aelam dicit Dominus
JER|50|1|verbum quod locutus est Dominus de Babylone et de terra Chaldeorum in manu Hieremiae prophetae
JER|50|2|adnuntiate in gentibus et auditum facite levate signum praedicate et nolite celare dicite capta est Babylon confusus est Bel victus est Marodach confusa sunt sculptilia eius superata sunt idola eorum
JER|50|3|quoniam ascendit contra eam gens ab aquilone quae ponet terram eius in solitudinem et non erit qui habitet in ea ab homine usque ad pecus et moti sunt et abierunt
JER|50|4|in diebus illis et in tempore illo ait Dominus venient filii Israhel ipsi et filii Iuda simul ambulantes et flentes properabunt et Dominum Deum suum quaerent
JER|50|5|in Sion interrogabunt viam huc facies eorum venient et adponentur ad Dominum foedere sempiterno quod nulla oblivione delebitur
JER|50|6|grex perditus factus est populus meus pastores eorum seduxerunt eos feceruntque vagari in montibus de monte in collem transierunt obliti sunt cubilis sui
JER|50|7|omnes qui invenerunt comederunt eos et hostes eorum dixerunt non peccavimus pro eo quod peccaverunt Domino decori iustitiae et expectationi patrum eorum Domino
JER|50|8|recedite de medio Babylonis et de terra Chaldeorum egredimini et estote quasi hedi ante greges
JER|50|9|quoniam ecce ego suscito et adducam in Babylonem congregationem gentium magnarum de terra aquilonis et praeparabuntur adversum eam et inde capietur sagitta eius quasi viri fortis interfectoris non revertetur vacua
JER|50|10|et erit Chaldea in praedam omnes vastantes eam replebuntur ait Dominus
JER|50|11|quoniam exultatis et magna loquimini diripientes hereditatem meam quoniam effusi estis sicut vitulus super herbam et mugistis ut tauri
JER|50|12|confusa est mater vestra nimis et adaequata pulveri quae genuit vos ecce novissima erit in gentibus deserta invia et arens
JER|50|13|ab ira Domini non habitabitur sed redigetur tota in solitudinem omnis qui transit per Babylonem stupebit et sibilabit super universis plagis eius
JER|50|14|praeparamini contra Babylonem per circuitum omnes qui intenditis arcum debellate eam non parcatis iaculis quia Domino peccavit
JER|50|15|clamate adversus eam ubique dedit manum ceciderunt fundamenta eius destructi sunt muri eius quoniam ultio Domini est ultionem accipite de ea sicut fecit facite ei
JER|50|16|disperdite satorem de Babylone et tenentem falcem in tempore messis a facie gladii columbae unusquisque ad populum suum convertetur et singuli ad terram suam fugient
JER|50|17|grex dispersus Israhel leones eiecerunt eum primus comedit eum rex Assur iste novissimus exossavit eum Nabuchodonosor rex Babylonis
JER|50|18|propterea haec dicit Dominus exercituum Deus Israhel ecce ego visitabo regem Babylonis et terram eius sicut visitavi regem Assur
JER|50|19|et reducam Israhel ad habitaculum suum et pascetur Carmelum et Basan et in monte Ephraim et Galaad saturabitur anima eius
JER|50|20|in diebus illis et in tempore illo ait Dominus quaeretur iniquitas Israhel et non erit et peccatum Iuda et non invenietur quoniam propitius ero eis quos reliquero
JER|50|21|super terram dominantium ascende et super habitatores eius visita dissipa et interfice quae post eos sunt ait Dominus et fac iuxta omnia quae praecepi tibi
JER|50|22|vox belli in terra et contritio magna
JER|50|23|quomodo confractus est et contritus est malleus universae terrae quomodo versa est in desertum Babylon in gentibus
JER|50|24|inlaqueavi te et capta es Babylon et nesciebas inventa es et adprehensa quoniam Dominum provocasti
JER|50|25|aperuit Dominus thesaurum suum et protulit vasa irae suae quoniam opus est Domino Deo exercituum in terra Chaldeorum
JER|50|26|venite ad eam ab extremis finibus aperite ut exeant qui conculcent eam tollite de via lapides et redigite in acervos et interficite eam nec sit quicquam reliquum
JER|50|27|dissipate universos fortes eius descendant in occisionem vae eis quia venit dies eorum tempus visitationis eorum
JER|50|28|vox fugientium et eorum qui evaserunt de terra Babylonis ut adnuntient in Sion ultionem Domini Dei nostri ultionem templi eius
JER|50|29|adnuntiate in Babylonem plurimis omnibus qui tendunt arcum consistite adversum eam per gyrum et nullus evadat reddite ei secundum opus suum iuxta omnia quae fecit facite illi quia contra Dominum erecta est adversum Sanctum Israhel
JER|50|30|idcirco cadent iuvenes eius in plateis eius et omnes viri bellatores eius conticescent in die illa ait Dominus
JER|50|31|ecce ego ad te superbe dicit Dominus Deus exercituum quia venit dies tuus tempus visitationis tuae
JER|50|32|et cadet superbus et corruet et non erit qui suscitet eum et succendam ignem in urbibus eius et devorabit omnia in circuitu eius
JER|50|33|haec dicit Dominus exercituum calumniam sustinent filii Israhel et filii Iuda simul omnes qui ceperunt eos tenent nolunt dimittere eos
JER|50|34|redemptor eorum Fortis Dominus exercituum nomen eius iudicio defendet causam eorum ut exterreat terram et commoveat habitatores Babylonis
JER|50|35|gladius ad Chaldeos ait Dominus et ad habitatores Babylonis et ad principes et ad sapientes eius
JER|50|36|gladius ad divinos eius qui stulti erunt gladius ad fortes illius qui timebunt
JER|50|37|gladius ad equos eius et ad currus eius et ad omne vulgus quod est in medio eius et erunt quasi mulieres gladius ad thesauros eius qui diripientur
JER|50|38|siccitas super aquas eius erit et arescent quia terra sculptilium est et in portentis gloriantur
JER|50|39|propterea habitabunt dracones cum fatuis ficariis et habitabunt in ea strutiones et non habitabitur ultra usque ad sempiternum nec extruetur usque ad generationem et generationem
JER|50|40|sicut subvertit Deus Sodomam et Gomorram et vicinas eius ait Dominus non habitabit ibi vir nec incolet eam filius hominis
JER|50|41|ecce populus venit ab aquilone et gens magna et reges multi consurgent a finibus terrae
JER|50|42|arcum et scutum adprehendent crudeles sunt et inmisericordes vox eorum quasi mare sonabit et super equos ascendent sicut vir paratus ad proelium contra te filia Babylon
JER|50|43|audivit rex Babylonis famam eorum et dissolutae sunt manus eius angustia adprehendit eum dolor quasi parturientem
JER|50|44|ecce quasi leo ascendet de superbia Iordanis ad pulchritudinem robustam quia subito currere eum faciam ad illam et quis erit electus quem praeponam ei quis enim similis mei et quis sustinebit me et quis est iste pastor qui resistat vultui meo
JER|50|45|propterea audite consilium Domini quod mente concepit adversum Babylonem et cogitationes eius quas cogitavit super terram Chaldeorum nisi detraxerint eos parvuli gregum nisi dissipatum fuerit cum ipsis habitaculum eorum
JER|50|46|a voce captivitatis Babylonis commota est terra et clamor inter gentes auditus est
JER|51|1|haec dicit Dominus ecce ego suscitabo super Babylonem et super habitatores eius qui cor suum levaverunt contra me quasi ventum pestilentem
JER|51|2|et mittam in Babylonem ventilatores et ventilabunt eam et demolientur terram eius quoniam venerunt super eam undique in die adflictionis eius
JER|51|3|non tendat qui tendit arcum suum et non ascendat loricatus nolite parcere iuvenibus eius interficite omnem militiam eius
JER|51|4|et cadent interfecti in terra Chaldeorum et vulnerati in regionibus eius
JER|51|5|quoniam non fuit viduatus Israhel et Iuda a Deo suo Domino exercituum terra autem eorum repleta est delicto a Sancto Israhel
JER|51|6|fugite de medio Babylonis et salvet unusquisque animam suam nolite tacere super iniquitatem eius quoniam tempus ultionis est Domino vicissitudinem ipse retribuet ei
JER|51|7|calix aureus Babylon in manu Domini inebrians omnem terram de vino eius biberunt gentes et ideo commotae sunt
JER|51|8|subito cecidit Babylon et contrita est ululate super eam tollite resinam ad dolorem eius si forte sanetur
JER|51|9|curavimus Babylonem et non est sanata derelinquamus eam et eamus unusquisque in terram suam quoniam pervenit usque ad caelos iudicium eius et elevatum est usque ad nubes
JER|51|10|protulit Dominus iustitias nostras venite et narremus in Sion opus Domini Dei nostri
JER|51|11|acuite sagittas implete faretras suscitavit Dominus spiritum regum Medorum et contra Babylonem mens eius ut perdat eam quoniam ultio Domini est ultio templi sui
JER|51|12|super muros Babylonis levate signum augete custodiam levate custodes praeparate insidias quia cogitavit Dominus et fecit quaecumque locutus est contra habitatores Babylonis
JER|51|13|quae habitas super aquas multas locuples in thesauris venit finis tuus pedalis praecisionis tuae
JER|51|14|iuravit Dominus exercituum per animam suam quoniam replebo te hominibus quasi brucho et super te celeuma cantabitur
JER|51|15|qui fecit terram in fortitudine sua praeparavit orbem in sapientia sua et prudentia sua extendit caelos
JER|51|16|dante eo vocem multiplicantur aquae in caelo qui levat nubes ab extremo terrae fulgura in pluviam fecit et produxit ventum de thesauris suis
JER|51|17|stultus factus est omnis homo ab scientia confusus est omnis conflator in sculptili quia mendax conflatio eius nec est spiritus in eis
JER|51|18|vana sunt opera et risu digna in tempore visitationis suae peribunt
JER|51|19|non sicut haec pars Iacob quia qui fecit omnia ipse est et Israhel sceptrum hereditatis eius Dominus exercituum nomen eius
JER|51|20|conlidis tu mihi vasa belli et ego conlidam in te gentes et disperdam in te regna
JER|51|21|et conlidam in te equum et equitem eius et conlidam in te currum et ascensorem eius
JER|51|22|et conlidam in te virum et mulierem et conlidam in te senem et puerum et conlidam in te iuvenem et virginem
JER|51|23|et conlidam in te pastorem et gregem eius et conlidam in te agricolam et iugales eius et conlidam in te duces et magistratus
JER|51|24|et reddam Babyloni et cunctis habitatoribus Chaldeae omne malum suum quod fecerunt in Sion in oculis vestris ait Dominus
JER|51|25|ecce ego ad te mons pestifer ait Dominus qui corrumpis universam terram et extendam manum meam super te et evolvam te de petris et dabo te in montem conbustionis
JER|51|26|et non tollent de te lapidem in angulum et lapidem in fundamenta sed perditus in aeternum eris ait Dominus
JER|51|27|levate signum in terra clangite bucina in gentibus sanctificate super eam gentes adnuntiate contra illam regibus Ararat Menni et Aschenez numerate contra eam Thapsar adducite equum quasi bruchum aculeatum
JER|51|28|sanctificate contra eam gentes reges Mediae duces eius et universos magistratus eius cunctamque terram potestatis eius
JER|51|29|et commovebitur terra et turbabitur quia evigilavit contra Babylonem cogitatio Domini ut ponat terram Babylonis desertam et inhabitabilem
JER|51|30|cessaverunt fortes Babylonis a proelio habitaverunt in praesidiis devoratum est robur eorum et facti sunt quasi mulieres incensa sunt tabernacula eius contriti sunt vectes eius
JER|51|31|currens obviam currenti veniet et nuntius obvius nuntianti ut adnuntiet regi Babylonis quia capta est civitas eius a summo usque ad summum
JER|51|32|et vada praeoccupata sunt et paludes incensae sunt igni et viri bellatores conturbati sunt
JER|51|33|quia haec dicit Dominus exercituum Deus Israhel filia Babylon quasi area tempus triturae eius adhuc modicum et veniet tempus messionis eius
JER|51|34|comedit me devoravit me Nabuchodonosor rex Babylonis reddidit me quasi vas inane absorbuit me sicut draco replevit ventrem suum teneritudine mea et eiecit me
JER|51|35|iniquitas adversum me et caro mea super Babylonem dicit habitatio Sion et sanguis meus super habitatores Chaldeae dicit Hierusalem
JER|51|36|propterea haec dicit Dominus ecce ego iudicabo causam tuam et ulciscar ultionem tuam et desertum faciam mare eius et siccabo venam eius
JER|51|37|et erit Babylon in tumulos habitatio draconum stupor et sibilus eo quod non sit habitator
JER|51|38|simul ut leones rugient excutient comas velut catuli leonum
JER|51|39|in calore eorum ponam potus eorum et inebriabo eos ut sopiantur et dormiant somnum sempiternum et non consurgant dicit Dominus
JER|51|40|deducam eos quasi agnos ad victimam quasi arietes cum hedis
JER|51|41|quomodo capta est Sesach et conprehensa est inclita universae terrae quomodo facta est in stuporem Babylon inter gentes
JER|51|42|ascendit super Babylonem mare multitudine fluctuum eius operta est
JER|51|43|factae sunt civitates eius in stuporem terra inhabitabilis et deserta terra in qua nullus habitet nec transeat per eam filius hominis
JER|51|44|et visitabo super Bel in Babylone et eiciam quod absorbuerat de ore eius et non confluent ad eum ultra gentes siquidem et murus Babylonis corruit
JER|51|45|egredimini de medio eius populus meus ut salvet unusquisque animam suam ab ira furoris Domini
JER|51|46|et ne forte mollescat cor vestrum et timeatis auditum qui audietur in terra et veniet in anno auditio et post hunc annum auditio et iniquitas in terra et dominator super dominatorem
JER|51|47|propterea ecce dies veniunt et visitabo super sculptilia Babylonis et omnis terra eius confundetur et universi interfecti eius cadent in medio eius
JER|51|48|et laudabunt super Babylonem caeli et terra et omnia quae in eis sunt quia ab aquilone venient ei praedones ait Dominus
JER|51|49|et quomodo fecit Babylon ut caderent occisi in Israhel sic de Babylone cadent occisi in universa terra
JER|51|50|qui fugistis gladium venite nolite stare recordamini procul Domini et Hierusalem ascendat super cor vestrum
JER|51|51|confusi sumus quoniam audivimus obprobrium operuit ignominia facies nostras quia venerunt alieni super sanctificationem domus Domini
JER|51|52|propterea ecce dies veniunt ait Dominus et visitabo super sculptilia eius et in omni terra eius mugiet vulneratus
JER|51|53|si ascenderit Babylon in caelum et firmaverit in excelso robur suum a me venient vastatores eius ait Dominus
JER|51|54|vox clamoris de Babylone et contritio magna de terra Chaldeorum
JER|51|55|quoniam vastavit Dominus Babylonem et perdidit ex ea vocem magnam et sonabunt fluctus eorum quasi aquae multae dedit sonitum vox eorum
JER|51|56|quia venit super eam id est super Babylonem praedo et adprehensi sunt fortes eius et emarcuit arcus eorum quia fortis ultor Dominus reddens retribuet
JER|51|57|et inebriabo principes eius et sapientes eius duces eius et magistratus eius et fortes eius et dormient somnum sempiternum et non expergiscentur ait Rex Dominus exercituum nomen eius
JER|51|58|haec dicit Dominus exercituum murus Babylonis ille latissimus suffossione suffodietur et portae eius excelsae igni conburentur et labores populorum ad nihilum et gentium in igne erunt et disperibunt
JER|51|59|verbum quod praecepit Hieremias prophetes Saraiae filio Neriae filii Maasiae cum pergeret cum Sedecia rege in Babylonem in anno quarto regni eius Saraias autem erat princeps prophetiae
JER|51|60|et scripsit Hieremias omne malum quod venturum erat super Babylonem in libro uno omnia verba haec quae scripta sunt contra Babylonem
JER|51|61|et dixit Hieremias ad Saraiam cum veneris Babylonem et videris et legeris omnia verba haec
JER|51|62|dices Domine tu locutus es contra locum istum ut disperderes eum ne sit qui in eo habitet ab homine usque ad pecus et ut sit perpetua solitudo
JER|51|63|cumque conpleveris legere librum istum ligabis ad eum lapidem et proicies illum in medio Eufraten
JER|51|64|et dices sic submergetur Babylon et non consurget a facie adflictionis quam ego adduco super eam et dissolventur hucusque verba Hieremiae
JER|52|1|filius viginti et unius anni Sedecias cum regnare coepisset et undecim annis regnavit in Hierusalem et nomen matris eius Amithal filia Hieremiae de Lobna
JER|52|2|et fecit malum in oculis Domini iuxta omnia quae fecerat Ioachim
JER|52|3|quoniam furor Domini erat in Hierusalem et in Iuda usquequo proiceret eos a facie sua et recessit Sedecias a rege Babylonis
JER|52|4|factum est autem in anno nono regni eius in mense decimo decima mensis venit Nabuchodonosor rex Babylonis ipse et omnis exercitus eius adversum Hierusalem et obsederunt eam et aedificaverunt contra eam munitiones in circuitu
JER|52|5|et fuit civitas obsessa usque ad undecimum annum regis Sedeciae
JER|52|6|mense autem quarto nona mensis obtinuit fames in civitate et non erant alimenta populo terrae
JER|52|7|et disrupta est civitas et omnes viri bellatores fugerunt et exierunt de civitate nocte per viam portae quae est inter duos muros et ducit ad hortum regis Chaldeis obsidentibus urbem in gyro et abierunt per viam quae ducit in heremum
JER|52|8|persecutus est autem exercitus Chaldeorum regem et adprehenderunt Sedeciam in deserto quod est iuxta Hiericho et omnis comitatus eius diffugit ab eo
JER|52|9|cumque conprehendissent regem adduxerunt eum ad regem Babylonis in Reblatha quae est in terra Emath et locutus est ad eum iudicia
JER|52|10|et iugulavit rex Babylonis filios Sedeciae in oculis eius sed et omnes principes Iudae occidit in Reblatha
JER|52|11|et oculos Sedeciae eruit et vinxit eum conpedibus et adduxit eum rex Babylonis in Babylonem et posuit eum in domo carceris usque ad diem mortis eius
JER|52|12|in mense autem quinto decima mensis ipse est annus nonusdecimus Nabuchodonosor regis Babylonis venit Nabuzardan princeps militiae qui stabat coram rege Babylonis in Hierusalem
JER|52|13|et incendit domum Domini et domum regis et omnes domos Hierusalem et omnem domum magnam igne conbusit
JER|52|14|et totum murum Hierusalem per circuitum destruxit cunctus exercitus Chaldeorum qui erat cum magistro militiae
JER|52|15|de pauperibus autem populi et de reliquo vulgo quod remanserat in civitate et de perfugis qui transfugerant ad regem Babylonis et ceteros de multitudine transtulit Nabuzardan princeps militiae
JER|52|16|de pauperibus vero terrae reliquit Nabuzardan princeps militiae in vinitores et in agricolas
JER|52|17|columnas quoque aereas quae erant in domo Domini et bases et mare aereum quod erat in domo Domini confregerunt Chaldei et tulerunt omne aes eorum in Babylonem
JER|52|18|et lebetas et creagras et psalteria et fialas et mortariola et omnia vasa aerea quae in ministerio fuerant tulerunt
JER|52|19|et hydrias et thymiamateria et urceos et pelves et candelabra et mortaria et cyatos quotquot aurea aurea et quotquot argentea argentea tulit magister militiae
JER|52|20|columnas duas et mare unum vitulos duodecim aereos qui erant sub basibus quas fecerat rex Salomon in domo Domini non erat pondus aeris omnium vasorum horum
JER|52|21|de columnis autem decem et octo cubiti altitudinis erant in columna una et funiculus duodecim cubitorum circuibat eam porro grossitudo eius quattuor digitorum et intrinsecus cava erat
JER|52|22|et capitella super utramque aerea altitudo capitelli unius quinque cubitorum et retiacula et mala granata
JER|52|23|nonaginta sex dependentia omnia mala granata centum retiaculis circumdabantur
JER|52|24|et tulit magister militiae Saraiam sacerdotem primum et Sophoniam sacerdotem secundum et tres custodes vestibuli
JER|52|25|et de civitate tulit eunuchum unum qui erat praepositus super viros bellatores et septem viros de his qui videbant faciem regis qui inventi sunt in civitate et scribam principem militum qui probabat tirones et sexaginta viros de populo terrae qui inventi sunt in medio civitatis
JER|52|26|tulit autem eos Nabuzardan magister militiae et duxit eos ad regem Babylonis in Reblatha
JER|52|27|et percussit eos rex Babylonis et interfecit eos in Reblatha in terra Emath et translatus est Iuda de terra sua
JER|52|28|iste est populus quem transtulit Nabuchodonosor in anno septimo Iudaeos tria milia et viginti tres
JER|52|29|in anno octavodecimo Nabuchodonosor de Hierusalem animas octingentas triginta duas
JER|52|30|in anno vicesimo tertio Nabuchodonosor transtulit Nabuzardan magister militiae Iudaeorum animas septingentas quadraginta quinque omnes ergo animae quattuor milia sescentae
JER|52|31|et factum est in tricesimo septimo anno transmigrationis Ioachim regis Iudae duodecimo mense vicesima quinta mensis elevavit Evilmerodach rex Babylonis ipso anno regni sui caput Ioachim regis Iudae et eduxit eum de domo carceris
JER|52|32|et locutus est cum eo bona et posuit thronum eius super thronos regum qui erant post se in Babylone
JER|52|33|et mutavit vestimenta carceris eius et comedebat panem coram eo semper cunctis diebus vitae suae
JER|52|34|et cibaria eius cibaria perpetua dabantur ei a rege Babylonis statuta per singulos dies usque ad diem mortis suae cunctis diebus vitae eius
LAM|1|1|ALEPH quomodo sedit sola civitas plena populo facta est quasi vidua domina gentium princeps provinciarum facta est sub tributo
LAM|1|2|BETH plorans ploravit in nocte et lacrimae eius in maxillis eius non est qui consoletur eam ex omnibus caris eius omnes amici eius spreverunt eam et facti sunt ei inimici
LAM|1|3|GIMEL migravit Iuda propter adflictionem et multitudinem servitutis habitavit inter gentes nec invenit requiem omnes persecutores eius adprehenderunt eam inter angustias
LAM|1|4|DELETH viae Sion lugent eo quod non sint qui veniant ad sollemnitatem omnes portae eius destructae sacerdotes eius gementes virgines eius squalidae et ipsa oppressa amaritudine
LAM|1|5|HE facti sunt hostes eius in capite inimici illius locupletati sunt quia Dominus locutus est super eam propter multitudinem iniquitatum eius parvuli eius ducti sunt captivi ante faciem tribulantis
LAM|1|6|VAV et egressus est a filia Sion omnis decor eius facti sunt principes eius velut arietes non invenientes pascuam et abierunt absque fortitudine ante faciem subsequentis
LAM|1|7|ZAI recordata est Hierusalem dierum adflictionis suae et praevaricationis omnium desiderabilium suorum quae habuerat a diebus antiquis cum caderet populus eius in manu hostili et non esset auxiliator viderunt eam hostes et deriserunt sabbata eius
LAM|1|8|HETH peccatum peccavit Hierusalem propterea instabilis facta est omnes qui glorificabant eam spreverunt illam quia viderunt ignominiam eius ipsa autem gemens et conversa retrorsum
LAM|1|9|TETH sordes eius in pedibus eius nec recordata est finis sui deposita est vehementer non habens consolatorem vide Domine adflictionem meam quoniam erectus est inimicus
LAM|1|10|IOTH manum suam misit hostis ad omnia desiderabilia eius quia vidit gentes ingressas sanctuarium suum de quibus praeceperas ne intrarent in ecclesiam tuam
LAM|1|11|CAPH omnis populus eius gemens et quaerens panem dederunt pretiosa quaeque pro cibo ad refocilandam animam vide Domine considera quoniam facta sum vilis
LAM|1|12|LAMED o vos omnes qui transitis per viam adtendite et videte si est dolor sicut dolor meus quoniam vindemiavit me ut locutus est Dominus in die irae furoris sui
LAM|1|13|MEM de excelso misit ignem in ossibus meis et erudivit me expandit rete pedibus meis convertit me retrorsum posuit me desolatam tota die maerore confectam
LAM|1|14|NUN vigilavit iugum iniquitatum mearum in manu eius convolutae sunt et inpositae collo meo infirmata est virtus mea dedit me Dominus in manu de qua non potero surgere
LAM|1|15|SAMECH abstulit omnes magnificos meos Dominus de medio mei vocavit adversum me tempus ut contereret electos meos torcular calcavit Dominus virgini filiae Iuda
LAM|1|16|AIN idcirco ego plorans et oculus meus deducens aquam quia longe factus est a me consolator convertens animam meam facti sunt filii mei perditi quoniam invaluit inimicus
LAM|1|17|FE expandit Sion manus suas non est qui consoletur eam mandavit Dominus adversum Iacob in circuitu eius hostes eius facta est Hierusalem quasi polluta menstruis inter eos
LAM|1|18|SADE iustus est Dominus quia os eius ad iracundiam provocavi audite obsecro universi populi et videte dolorem meum virgines meae et iuvenes mei abierunt in captivitatem
LAM|1|19|COPH vocavi amicos meos et ipsi deceperunt me sacerdotes mei et senes mei in urbe consumpti sunt quia quaesierunt cibum sibi ut refocilarent animam suam
LAM|1|20|RES vide Domine quoniam tribulor venter meus conturbatus est subversum est cor meum in memet ipsa quoniam amaritudine plena sum foris interfecit gladius et domi mors similis est
LAM|1|21|SEN audierunt quia ingemesco ego et non est qui consoletur me omnes inimici mei audierunt malum meum laetati sunt quoniam tu fecisti adduxisti diem consolationis et fient similes mei
LAM|1|22|THAU ingrediatur omne malum eorum coram te et devindemia eos sicut vindemiasti me propter omnes iniquitates meas multi enim gemitus mei et cor meum maerens
LAM|2|1|ALEPH quomodo obtexit caligine in furore suo Dominus filiam Sion proiecit de caelo terram inclitam Israhel et non recordatus est scabilli pedum suorum in die furoris sui
LAM|2|2|BETH praecipitavit Dominus nec pepercit omnia speciosa Iacob destruxit in furore suo munitiones virginis Iuda deiecit in terram polluit regnum et principes eius
LAM|2|3|GIMEL confregit in ira furoris omne cornu Israhel avertit retrorsum dexteram suam a facie inimici et succendit in Iacob quasi ignem flammae devorantis in gyro
LAM|2|4|DELETH tetendit arcum suum quasi inimicus firmavit dexteram suam quasi hostis et occidit omne quod pulchrum erat visu in tabernaculo filiae Sion effudit quasi ignem indignationem suam
LAM|2|5|HE factus est Dominus velut inimicus praecipitavit Israhel praecipitavit omnia moenia eius dissipavit munitiones eius et replevit in filia Iuda humiliatum et humiliatam
LAM|2|6|VAV et dissipavit quasi hortum tentorium suum demolitus est tabernaculum suum oblivioni tradidit Dominus in Sion festivitatem et sabbatum et obprobrio in indignatione furoris sui regem et sacerdotem
LAM|2|7|ZAI reppulit Dominus altare suum maledixit sanctificationi suae tradidit in manu inimici muros turrium eius vocem dederunt in domo Domini sicut in die sollemni
LAM|2|8|HETH cogitavit Dominus dissipare murum filiae Sion tetendit funiculum suum et non avertit manum suam a perditione luxitque antemurale et murus pariter dissipatus est
LAM|2|9|TETH defixae sunt in terra portae eius perdidit et contrivit vectes eius regem eius et principes eius in gentibus non est lex et prophetae eius non invenerunt visionem a Domino
LAM|2|10|IOTH sederunt in terra conticuerunt senes filiae Sion consperserunt cinere capita sua accincti sunt ciliciis abiecerunt in terra capita sua virgines Hierusalem
LAM|2|11|CAPH defecerunt prae lacrimis oculi mei conturbata sunt viscera mea effusum est in terra iecur meum super contritione filiae populi mei cum deficeret parvulus et lactans in plateis oppidi
LAM|2|12|LAMED matribus suis dixerunt ubi est triticum et vinum cum deficerent quasi vulnerati in plateis civitatis cum exhalarent animas suas in sinu matrum suarum
LAM|2|13|MEM cui conparabo te vel cui adsimilabo te filia Hierusalem cui exaequabo te et consolabor te virgo filia Sion magna enim velut mare contritio tua quis medebitur tui
LAM|2|14|NUN prophetae tui viderunt tibi falsa et stulta nec aperiebant iniquitatem tuam ut te ad paenitentiam provocarent viderunt autem tibi adsumptiones falsas et eiectiones
LAM|2|15|SAMECH plauserunt super te manibus omnes transeuntes per viam sibilaverunt et moverunt caput suum super filiam Hierusalem haecine est urbs dicentes perfecti decoris gaudium universae terrae
LAM|2|16|FE aperuerunt super te os suum omnes inimici tui sibilaverunt et fremuerunt dentibus dixerunt devoravimus en ista est dies quam expectabamus invenimus vidimus
LAM|2|17|AIN fecit Dominus quae cogitavit conplevit sermonem suum quem praeceperat a diebus antiquis destruxit et non pepercit et laetificavit super te inimicum et exaltavit cornu hostium tuorum
LAM|2|18|SADE clamavit cor eorum ad Dominum super muros filiae Sion deduc quasi torrentem lacrimas per diem et per noctem non des requiem tibi neque taceat pupilla oculi tui
LAM|2|19|COPH consurge lauda in nocte in principio vigiliarum effunde sicut aqua cor tuum ante conspectum Domini leva ad eum manus tuas pro anima parvulorum tuorum qui defecerunt in fame in capite omnium conpetorum
LAM|2|20|RES vide Domine et considera quem vindemiaveris ita ergone comedent mulieres fructum suum parvulos ad mensuram palmae si occidetur in sanctuario Domini sacerdos et propheta
LAM|2|21|SEN iacuerunt in terra foris puer et senex virgines meae et iuvenes mei ceciderunt in gladio interfecisti in die furoris tui percussisti nec misertus es
LAM|2|22|THAU vocasti quasi ad diem sollemnem qui terrerent me de circuitu et non fuit in die furoris Domini qui effugeret et relinqueretur quos educavi et enutrivi inimicus meus consumpsit eos
LAM|3|1|ALEPH ego vir videns paupertatem meam in virga indignationis eius
LAM|3|2|ALEPH me minavit et adduxit in tenebris et non in lucem
LAM|3|3|ALEPH tantum in me vertit et convertit manum suam tota die
LAM|3|4|BETH vetustam fecit pellem meam et carnem meam contrivit ossa mea
LAM|3|5|BETH aedificavit in gyro meo et circumdedit me felle et labore
LAM|3|6|BETH in tenebrosis conlocavit me quasi mortuos sempiternos
LAM|3|7|GIMEL circumaedificavit adversum me ut non egrediar adgravavit conpedem meam
LAM|3|8|GIMEL sed et cum clamavero et rogavero exclusit orationem meam
LAM|3|9|GIMEL conclusit vias meas lapidibus quadris semitas meas subvertit
LAM|3|10|DELETH ursus insidians factus est mihi leo in absconditis
LAM|3|11|DELETH semitas meas subvertit et confregit me posuit me desolatam
LAM|3|12|DELETH tetendit arcum suum et posuit me quasi signum ad sagittam
LAM|3|13|HE misit in renibus meis filias faretrae suae
LAM|3|14|HE factus sum in derisu omni populo meo canticum eorum tota die
LAM|3|15|HE replevit me amaritudinibus inebriavit me absinthio
LAM|3|16|VAV et fregit ad numerum dentes meos cibavit me cinere
LAM|3|17|VAV et repulsa est anima mea oblitus sum bonorum
LAM|3|18|VAV et dixi periit finis meus et spes mea a Domino
LAM|3|19|ZAI recordare paupertatis et transgressionis meae absinthii et fellis
LAM|3|20|ZAI memoria memor ero et tabescet in me anima mea
LAM|3|21|ZAI hoc recolens in corde meo ideo sperabo
LAM|3|22|HETH misericordiae Domini quia non sumus consumpti quia non defecerunt miserationes eius
LAM|3|23|HETH novae diluculo multa est fides tua
LAM|3|24|HETH pars mea Dominus dixit anima mea propterea expectabo eum
LAM|3|25|TETH bonus est Dominus sperantibus in eum animae quaerenti illum
LAM|3|26|TETH bonum est praestolari cum silentio salutare Domini
LAM|3|27|TETH bonum est viro cum portaverit iugum ab adulescentia sua
LAM|3|28|IOTH sedebit solitarius et tacebit quia levavit super se
LAM|3|29|IOTH ponet in pulvere os suum si forte sit spes
LAM|3|30|IOTH dabit percutienti se maxillam saturabitur obprobriis
LAM|3|31|CAPH quia non repellet in sempiternum Dominus
LAM|3|32|CAPH quia si abiecit et miserebitur secundum multitudinem misericordiarum suarum
LAM|3|33|CAPH non enim humiliavit ex corde suo et abiecit filios hominis
LAM|3|34|LAMED ut contereret sub pedibus suis omnes vinctos terrae
LAM|3|35|LAMED ut declinaret iudicium viri in conspectu vultus Altissimi
LAM|3|36|LAMED ut perverteret hominem in iudicio suo Dominus ignoravit
LAM|3|37|MEM quis est iste qui dixit ut fieret Domino non iubente
LAM|3|38|MEM ex ore Altissimi non egredientur nec mala nec bona
LAM|3|39|MEM quid murmuravit homo vivens vir pro peccatis suis
LAM|3|40|NUN scrutemur vias nostras et quaeramus et revertamur ad Dominum
LAM|3|41|NUN levemus corda nostra cum manibus ad Dominum in caelos
LAM|3|42|NUN nos inique egimus et ad iracundiam provocavimus idcirco tu inexorabilis es
LAM|3|43|SAMECH operuisti in furore et percussisti nos occidisti nec pepercisti
LAM|3|44|SAMECH opposuisti nubem tibi ne transeat oratio
LAM|3|45|SAMECH eradicationem et abiectionem posuisti me in medio populorum
LAM|3|46|FE aperuerunt super nos os suum omnes inimici
LAM|3|47|FE formido et laqueus facta est nobis vaticinatio et contritio
LAM|3|48|FE divisiones aquarum deduxit oculus meus in contritione filiae populi mei
LAM|3|49|AIN oculus meus adflictus est nec tacuit eo quod non esset requies
LAM|3|50|AIN donec respiceret et videret Dominus de caelis
LAM|3|51|AIN oculus meus depraedatus est animam meam in cunctis filiabus urbis meae
LAM|3|52|SADE venatione ceperunt me quasi avem inimici mei gratis
LAM|3|53|SADE lapsa est in lacu vita mea et posuerunt lapidem super me
LAM|3|54|SADE inundaverunt aquae super caput meum dixi perii
LAM|3|55|COPH invocavi nomen tuum Domine de lacis novissimis
LAM|3|56|COPH vocem meam audisti ne avertas aurem tuam a singultu meo et clamoribus
LAM|3|57|COPH adpropinquasti in die quando invocavi te dixisti ne timeas
LAM|3|58|RES iudicasti Domine causam animae meae redemptor vitae meae
LAM|3|59|RES vidisti Domine iniquitatem adversum me iudica iudicium meum
LAM|3|60|RES vidisti omnem furorem universas cogitationes eorum adversum me
LAM|3|61|SEN audisti obprobria eorum Domine omnes cogitationes eorum adversum me
LAM|3|62|SEN labia insurgentium mihi et meditationes eorum adversum me tota die
LAM|3|63|SEN sessionem eorum et resurrectionem eorum vide ego sum psalmus eorum
LAM|3|64|THAU reddes eis vicem Domine iuxta opera manuum suarum
LAM|3|65|THAU dabis eis scutum cordis laborem tuum
LAM|3|66|THAU persequeris in furore et conteres eos sub caelis Domine
LAM|4|1|ALEPH quomodo obscuratum est aurum mutatus est color optimus dispersi sunt lapides sanctuarii in capite omnium platearum
LAM|4|2|BETH filii Sion incliti et amicti auro primo quomodo reputati sunt in vasa testea opus manuum figuli
LAM|4|3|GIMEL sed et lamiae nudaverunt mammam lactaverunt catulos suos filia populi mei crudelis quasi strutio in deserto
LAM|4|4|DELETH adhesit lingua lactantis ad palatum eius in siti parvuli petierunt panem et non erat qui frangeret eis
LAM|4|5|HE qui vescebantur voluptuose interierunt in viis qui nutriebantur in croceis amplexati sunt stercora
LAM|4|6|VAV et maior effecta est iniquitas filiae populi mei peccato Sodomorum quae subversa est in momento et non ceperunt in ea manus
LAM|4|7|ZAI candidiores nazarei eius nive nitidiores lacte rubicundiores ebore antiquo sapphyro pulchriores
LAM|4|8|HETH denigrata est super carbones facies eorum et non sunt cogniti in plateis adhesit cutis eorum ossibus aruit et facta est quasi lignum
LAM|4|9|TETH melius fuit occisis gladio quam interfectis fame quoniam isti extabuerunt consumpti ab sterilitate terrae
LAM|4|10|IOTH manus mulierum misericordium coxerunt filios suos facti sunt cibus earum in contritione filiae populi mei
LAM|4|11|CAPH conplevit Dominus furorem suum effudit iram indignationis suae et succendit ignem in Sion et devoravit fundamenta eius
LAM|4|12|LAMED non crediderunt reges terrae et universi habitatores orbis quoniam ingrederetur hostis et inimicus per portas Hierusalem
LAM|4|13|MEM propter peccata prophetarum eius iniquitates sacerdotum eius qui effuderunt in medio eius sanguinem iustorum
LAM|4|14|NUN erraverunt caeci in plateis polluti sunt sanguine cumque non possent tenuerunt lacinias suas
LAM|4|15|SAMECH recedite polluti clamaverunt eis recedite abite nolite tangere iurgati quippe sunt et commoti dixerunt inter gentes non addet ultra ut habitet in eis
LAM|4|16|FE facies Domini divisit eos non addet ut respiciat eos facies sacerdotum non erubuerunt neque senum miserti sunt
LAM|4|17|AIN cum adhuc subsisteremus defecerunt oculi nostri ad auxilium nostrum vanum cum respiceremus adtenti ad gentem quae salvare non poterat
LAM|4|18|SADE lubricaverunt vestigia nostra in itinere platearum nostrarum adpropinquavit finis noster conpleti sunt dies nostri quia venit finis noster
LAM|4|19|COPH velociores fuerunt persecutores nostri aquilis caeli super montes persecuti sunt nos in deserto insidiati sunt nobis
LAM|4|20|RES spiritus oris nostri christus dominus captus est in peccatis nostris cui diximus in umbra tua vivemus in gentibus
LAM|4|21|SEN gaude et laetare filia Edom quae habitas in terra Hus ad te quoque perveniet calix inebriaberis atque nudaberis
LAM|4|22|THAU conpleta est iniquitas tua filia Sion non addet ultra ut transmigret te visitavit iniquitatem tuam filia Edom discoperuit peccata tua
LAM|5|1|recordare Domine quid acciderit nobis intuere et respice obprobrium nostrum
LAM|5|2|hereditas nostra versa est ad alienos domus nostrae ad extraneos
LAM|5|3|pupilli facti sumus absque patre matres nostrae quasi viduae
LAM|5|4|aquam nostram pecunia bibimus ligna nostra pretio conparavimus
LAM|5|5|cervicibus minabamur lassis non dabatur requies
LAM|5|6|Aegypto dedimus manum et Assyriis ut saturaremur pane
LAM|5|7|patres nostri peccaverunt et non sunt et nos iniquitates eorum portavimus
LAM|5|8|servi dominati sunt nostri non fuit qui redimeret de manu eorum
LAM|5|9|in animabus nostris adferebamus panem nobis a facie gladii in deserto
LAM|5|10|pellis nostra quasi clibanus exusta est a facie tempestatum famis
LAM|5|11|mulieres in Sion humiliaverunt virgines in civitatibus Iuda
LAM|5|12|principes manu suspensi sunt facies senum non erubuerunt
LAM|5|13|adulescentibus inpudice abusi sunt et pueri in ligno corruerunt
LAM|5|14|senes de portis defecerunt iuvenes de choro psallentium
LAM|5|15|defecit gaudium cordis nostri versus est in luctu chorus noster
LAM|5|16|cecidit corona capitis nostri vae nobis quia peccavimus
LAM|5|17|propterea maestum factum est cor nostrum ideo contenebrati sunt oculi nostri
LAM|5|18|propter montem Sion quia disperiit vulpes ambulaverunt in eo
LAM|5|19|tu autem Domine in aeternum permanebis solium tuum in generatione et generatione
LAM|5|20|quare in perpetuum oblivisceris nostri derelinques nos in longitudinem dierum
LAM|5|21|converte nos Domine ad te et convertemur innova dies nostros sicut a principio
LAM|5|22|sed proiciens reppulisti nos iratus es contra nos vehementer
EZEK|1|1|et factum est in tricesimo anno in quarto mense in quinta mensis cum essem in medio captivorum iuxta fluvium Chobar aperti sunt caeli et vidi visiones Dei
EZEK|1|2|in quinta mensis ipse est annus quintus transmigrationis regis Ioachin
EZEK|1|3|factum est verbum Domini ad Hiezecihel filium Buzi sacerdotem in terra Chaldeorum secus flumen Chobar et facta est super eum ibi manus Domini
EZEK|1|4|et vidi et ecce ventus turbinis veniebat ab aquilone et nubes magna et ignis involvens et splendor in circuitu eius et de medio eius quasi species electri id est de medio ignis
EZEK|1|5|et ex medio eorum similitudo quattuor animalium et hic aspectus eorum similitudo hominis in eis
EZEK|1|6|et quattuor facies uni et quattuor pinnae uni
EZEK|1|7|et pedes eorum pedes recti et planta pedis eorum quasi planta pedis vituli et scintillae quasi aspectus aeris candentis
EZEK|1|8|et manus hominis sub pinnis eorum in quattuor partibus et facies et pinnas per quattuor partes habebant
EZEK|1|9|iunctaeque erant pinnae eorum alterius ad alterum non revertebantur cum incederent sed unumquodque ante faciem suam gradiebatur
EZEK|1|10|similitudo autem vultus eorum facies hominis et facies leonis a dextris ipsorum quattuor facies autem bovis a sinistris ipsorum quattuor et facies aquilae ipsorum quattuor
EZEK|1|11|et facies eorum et pinnae eorum extentae desuper duae pinnae singulorum iungebantur et duae tegebant corpora eorum
EZEK|1|12|et unumquodque coram facie sua ambulabat ubi erat impetus spiritus illuc gradiebantur nec revertebantur cum ambularent
EZEK|1|13|et similitudo animalium aspectus eorum quasi carbonum ignis ardentium et quasi aspectus lampadarum haec erat visio discurrens in medio animalium splendor ignis et de igne fulgor egrediens
EZEK|1|14|et animalia ibant et revertebantur in similitudinem fulguris coruscantis
EZEK|1|15|cumque aspicerem animalia apparuit rota una super terram iuxta animalia habens quattuor facies
EZEK|1|16|et aspectus rotarum et opus earum quasi visio maris et una similitudo ipsarum quattuor et aspectus earum et opera quasi sit rota in medio rotae
EZEK|1|17|per quattuor partes earum euntes ibant et non revertebantur cum ambularent
EZEK|1|18|statura quoque erat rotis et altitudo et horribilis aspectus et totum corpus plenum oculis in circuitu ipsarum quattuor
EZEK|1|19|cumque ambularent animalia ambulabant pariter et rotae iuxta ea et cum elevarentur animalia de terra elevabantur simul et rotae
EZEK|1|20|quocumque ibat spiritus illuc eunte spiritu et rotae pariter levabantur sequentes eum spiritus enim vitae erat in rotis
EZEK|1|21|cum euntibus ibant et cum stantibus stabant et cum elevatis a terra pariter elevabantur et rotae sequentes ea quia spiritus vitae erat in rotis
EZEK|1|22|et similitudo super caput animalium firmamenti quasi aspectus cristalli horribilis et extenti super capita eorum desuper
EZEK|1|23|sub firmamento autem pinnae eorum rectae alterius ad alterum unumquodque duabus alis velabat corpus suum et alterum similiter velabatur
EZEK|1|24|et audiebam sonum alarum quasi sonum aquarum multarum quasi sonum sublimis Dei cum ambularent quasi sonus erat multitudinis ut sonus castrorum cumque starent dimittebantur pinnae eorum
EZEK|1|25|nam cum fieret vox supra firmamentum quod erat super caput eorum stabant et submittebant alas suas
EZEK|1|26|et super firmamentum quod erat inminens capiti eorum quasi aspectus lapidis sapphyri similitudo throni et super similitudinem throni similitudo quasi aspectus hominis desuper
EZEK|1|27|et vidi quasi speciem electri velut aspectum ignis intrinsecus eius per circuitum a lumbis eius et desuper et a lumbis eius usque deorsum vidi quasi speciem ignis splendentis in circuitu
EZEK|1|28|velut aspectum arcus cum fuerit in nube in die pluviae hic erat aspectus splendoris per gyrum
EZEK|2|1|haec visio similitudinis gloriae Domini et vidi et cecidi in faciem meam et audivi vocem loquentis et dixit ad me fili hominis sta supra pedes tuos et loquar tecum
EZEK|2|2|et ingressus est in me spiritus postquam locutus est mihi et statuit me supra pedes meos et audivi loquentem ad me
EZEK|2|3|et dicentem fili hominis mitto ego te ad filios Israhel ad gentes apostatrices quae recesserunt a me patres eorum praevaricati sunt pactum meum usque ad diem hanc
EZEK|2|4|et filii dura facie et indomabili corde sunt ad quos ego mitto te et dices ad eos haec dicit Dominus Deus
EZEK|2|5|si forte vel ipsi audiant et si forte quiescant quoniam domus exasperans est et scient quia propheta fuerit in medio eorum
EZEK|2|6|tu ergo fili hominis ne timeas eos neque sermones eorum metuas quoniam increduli et subversores sunt tecum et cum scorpionibus habitas verba eorum ne timeas et vultus eorum ne formides quia domus exasperans est
EZEK|2|7|loqueris ergo verba mea ad eos si forte audiant et quiescant quoniam inritatores sunt
EZEK|2|8|tu autem fili hominis audi quaecumque loquor ad te et noli esse exasperans sicut domus exasperatrix est aperi os tuum et comede quaecumque ego do tibi
EZEK|2|9|et vidi et ecce manus missa ad me in qua erat involutus liber et expandit illum coram me qui erat scriptus intus et foris et scriptae erant in eo lamentationes et carmen et vae
EZEK|3|1|et dixit ad me fili hominis quodcumque inveneris comede comede volumen istud et vadens loquere ad filios Israhel
EZEK|3|2|et aperui os meum et cibavit me volumine illo
EZEK|3|3|et dixit ad me fili hominis venter tuus comedet et viscera tua conplebuntur volumine isto quod ego do tibi et comedi illud et factum est in ore meo sicut mel dulce
EZEK|3|4|et dixit ad me fili hominis vade ad domum Israhel et loqueris verba mea ad eos
EZEK|3|5|non enim ad populum profundi sermonis et ignotae linguae tu mitteris ad domum Israhel
EZEK|3|6|neque ad populos multos profundi sermonis et ignotae linguae quorum non possis audire sermones et si ad illos mittereris ipsi audirent te
EZEK|3|7|domus autem Israhel nolent audire te quia nolunt audire me omnis quippe domus Israhel adtrita fronte est et duro corde
EZEK|3|8|ecce dedi faciem tuam valentiorem faciebus eorum et frontem tuam duriorem frontibus eorum
EZEK|3|9|ut adamantem et ut silicem dedi faciem tuam ne timeas eos neque metuas a facie eorum quia domus exasperans est
EZEK|3|10|et dixit ad me fili hominis omnes sermones meos quos loquor ad te adsume in corde tuo et auribus tuis audi
EZEK|3|11|et vade ingredere ad transmigrationem ad filios populi tui et loqueris ad eos et dices eis haec dicit Dominus Deus si forte audiant et quiescant
EZEK|3|12|et adsumpsit me spiritus et audivi post me vocem commotionis magnae benedicta gloria Domini de loco suo
EZEK|3|13|et vocem alarum animalium percutientium alteram ad alteram et vocem rotarum sequentium animalia et vocem commotionis magnae
EZEK|3|14|spiritus quoque levavit me et adsumpsit me et abii amarus in indignatione spiritus mei manus enim Domini erat mecum confortans me
EZEK|3|15|et veni ad transmigrationem acervum novarum frugum ad eos qui habitabant iuxta flumen Chobar et sedi ubi illi sedebant et mansi ibi septem diebus maerens in medio eorum
EZEK|3|16|cum autem pertransissent septem dies factum est verbum Domini ad me dicens
EZEK|3|17|fili hominis speculatorem dedi te domui Israhel et audies de ore meo verbum et adnuntiabis eis ex me
EZEK|3|18|si dicente me ad impium morte morieris non adnuntiaveris ei neque locutus fueris ut avertatur a via sua impia et vivat ipse impius in iniquitate sua morietur sanguinem autem eius de manu tua requiram
EZEK|3|19|si autem tu adnuntiaveris impio et ille non fuerit conversus ab impietate sua et via sua impia ipse quidem in iniquitate sua morietur tu autem animam tuam liberasti
EZEK|3|20|sed et si conversus iustus a iustitia sua fecerit iniquitatem ponam offendiculum coram eo ipse morietur quia non adnuntiasti ei in peccato suo morietur et non erunt in memoria iustitiae eius quas fecit sanguinem vero eius de manu tua requiram
EZEK|3|21|si autem tu adnuntiaveris iusto ut non peccet iustus et ille non peccaverit vivens vivet quia adnuntiasti ei et tu animam tuam liberasti
EZEK|3|22|et facta est super me manus Domini et dixit ad me surgens egredere in campum et ibi loquar tecum
EZEK|3|23|et surgens egressus sum in campum et ecce ibi gloria Domini stabat quasi gloria quam vidi iuxta fluvium Chobar et cecidi in faciem meam
EZEK|3|24|et ingressus est in me spiritus et statuit me super pedes meos et locutus est mihi et dixit ad me ingredere et includere in medio domus tuae
EZEK|3|25|et tu fili hominis ecce data sunt super te vincula et ligabunt te in eis et non egredieris in medio eorum
EZEK|3|26|et linguam tuam adherescere faciam palato tuo et eris mutus nec quasi vir obiurgans quia domus exasperans est
EZEK|3|27|cum autem locutus fuero tibi aperiam os tuum et dices ad eos haec dicit Dominus Deus qui audit audiat et qui quiescit quiescat quia domus exasperans est
EZEK|4|1|et tu fili hominis sume tibi laterem et pones eum coram te et describes in eo civitatem Hierusalem
EZEK|4|2|et ordinabis adversus eam obsidionem et aedificabis munitiones et conportabis aggerem et dabis contra eam castra et pones arietes in gyro
EZEK|4|3|et tu sume tibi sartaginem ferream et pones eam murum ferreum inter te et inter civitatem et obfirmabis faciem tuam ad eam et erit in obsidionem et circumdabis eam signum est domui Israhel
EZEK|4|4|et tu dormies super latus tuum sinistrum et pones iniquitates domus Israhel super eo numero dierum quibus dormies super illud et adsumes iniquitatem eorum
EZEK|4|5|ego autem dedi tibi annos iniquitatis eorum numero dierum trecentos et nonaginta dies et portabis iniquitatem domus Israhel
EZEK|4|6|et cum conpleveris haec dormies super latus tuum dextrum secundo et adsumes iniquitatem domus Iuda quadraginta diebus diem pro anno diem inquam pro anno dedi tibi
EZEK|4|7|et ad obsidionem Hierusalem convertes faciem tuam et brachium tuum erit exertum et prophetabis adversus eam
EZEK|4|8|ecce circumdedi te vinculis et non te convertes a latere tuo in latus aliud donec conpleas dies obsidionis tuae
EZEK|4|9|et tu sume tibi frumentum et hordeum et fabam et lentem et milium et viciam et mittes ea in vas unum et facies tibi panes numero dierum quibus dormies super latus tuum trecentis et nonaginta diebus comedes illud
EZEK|4|10|cibus autem tuus quo vesceris erit in pondere viginti stateres in die a tempore usque ad tempus comedes illud
EZEK|4|11|et aquam in mensura bibes sextam partem hin a tempore usque ad tempus bibes illud
EZEK|4|12|et quasi subcinericium hordiacium comedes illud et stercore quod egredietur de homine operies illud in oculis eorum
EZEK|4|13|et dixit Dominus sic comedent filii Israhel panem suum pollutum inter gentes ad quas eiciam eos
EZEK|4|14|et dixi ha ha ha Domine Deus ecce anima mea non est polluta et morticinum et laceratum a bestiis non comedi ab infantia mea usque nunc et non est ingressa os meum omnis caro inmunda
EZEK|4|15|et dixit ad me ecce dedi tibi fimum boum pro stercoribus humanis et facies panem tuum in eo
EZEK|4|16|et dixit ad me fili hominis ecce ego conteram baculum panis in Hierusalem et comedent panem in pondere et in sollicitudine et aquam in mensura et in angustia bibent
EZEK|4|17|ut deficientibus pane et aqua corruat unusquisque ad fratrem suum et contabescant in iniquitatibus suis
EZEK|5|1|et tu fili hominis sume tibi gladium acutum radentem pilos adsumes eum et duces per caput tuum et per barbam tuam et adsumes tibi stateram ponderis et divides eos
EZEK|5|2|tertiam partem igni conbures in medio civitatis iuxta conpletionem dierum obsidionis et adsumens tertiam partem concides gladio in circuitu eius tertiam vero aliam disperges in ventum et gladium nudabo post eos
EZEK|5|3|et sumes inde parvum numerum et ligabis eos in summitate pallii tui
EZEK|5|4|et ex eis rursum tolles et proicies in medio ignis et conbures eos igni ex eo egredietur ignis in omnem domum Israhel
EZEK|5|5|haec dicit Dominus Deus ista est Hierusalem in medio gentium posui eam et in circuitu eius terras
EZEK|5|6|et contempsit iudicia mea ut plus esset impia quam gentes et praecepta mea ultra quam terrae quae in circuitu eius sunt iudicia enim mea proiecerunt et in praeceptis meis non ambulaverunt
EZEK|5|7|idcirco haec dicit Dominus Deus quia superastis gentes quae in circuitu vestro sunt in praeceptis meis non ambulastis et iudicia mea non fecistis et iuxta iudicia gentium quae in circuitu vestro sunt non estis operati
EZEK|5|8|ideo haec dicit Dominus Deus ecce ego ad te et ipse ego faciam in medio tui iudicia in oculis gentium
EZEK|5|9|et faciam in te quae non feci et quibus similia ultra non faciam propter omnes abominationes tuas
EZEK|5|10|ideo patres comedent filios in medio tui et filii comedent patres suos et faciam in te iudicia et ventilabo universas reliquias tuas in omnem ventum
EZEK|5|11|idcirco vivo ego dicit Dominus Deus nisi pro eo quod sanctum meum violasti in omnibus offensionibus tuis et in omnibus abominationibus tuis ego quoque confringam et non parcet oculus meus et non miserebor
EZEK|5|12|tertia tui pars peste morietur et fame consumetur in medio tui et tertia tui pars gladio cadet in circuitu tuo tertiam vero partem tuam in omnem ventum dispergam et gladium evaginabo post eos
EZEK|5|13|et conpleam furorem meum et requiescere faciam indignationem meam in eis et consolabor et scient quia ego Dominus locutus sum in zelo meo cum implevero indignationem meam in eis
EZEK|5|14|et dabo te in desertum et in obprobrium in gentibus quae in circuitu tuo sunt in conspectu omnis praetereuntis
EZEK|5|15|et eris obprobrium et blasphemia exemplum et stupor in gentibus quae in circuitu tuo sunt cum fecero in te iudicia in furore et in indignatione et in increpationibus irae
EZEK|5|16|ego Dominus locutus sum quando misero sagittas famis pessimas in eos quae erunt mortiferae et quas mittam ut disperdam vos et famem congregabo super vos et conteram vobis baculum panis
EZEK|5|17|et inmittam in vos famem et bestias pessimas usque ad internicionem et pestilentia et sanguis transibunt per te et gladium inducam super te ego Dominus locutus sum
EZEK|6|1|et factus est sermo Domini ad me dicens
EZEK|6|2|fili hominis pone faciem tuam ad montes Israhel et prophetabis ad eos
EZEK|6|3|et dices montes Israhel audite verbum Domini Dei haec dicit Dominus Deus montibus et collibus rupibus et vallibus ecce ego inducam super vos gladium et disperdam excelsa vestra
EZEK|6|4|et demoliar aras vestras et confringentur simulacra vestra et deiciam interfectos vestros ante idola vestra
EZEK|6|5|et dabo cadavera filiorum Israhel ante faciem simulacrorum vestrorum et dispergam ossa vestra circum aras vestras
EZEK|6|6|in omnibus habitationibus vestris urbes desertae erunt et excelsa demolientur et dissipabuntur et interibunt arae vestrae et confringentur et cessabunt idola vestra et conterentur delubra vestra et delebuntur opera vestra
EZEK|6|7|et cadet interfectus in medio vestri et scietis quoniam ego Dominus
EZEK|6|8|et relinquam in vobis eos qui fugerint gladium in gentibus cum dispersero vos in terris
EZEK|6|9|et recordabuntur mei liberati vestri in gentibus ad quas captivi ducti sunt quia contrivi cor eorum fornicans et recedens a me et oculos eorum fornicantes post idola sua et displicebunt sibimet super malis quae fecerunt in universis abominationibus suis
EZEK|6|10|et scient quia ego Dominus non frustra locutus sum ut facerem eis malum hoc
EZEK|6|11|haec dicit Dominus Deus percute manu tua et adlide pedem tuum et dic eheu ad omnes abominationes malorum domus Israhel qui gladio fame peste ruituri sunt
EZEK|6|12|qui longe est peste morietur qui autem prope gladio corruet et qui relictus fuerit et obsessus fame morietur et conpleam indignationem meam in eis
EZEK|6|13|et scietis quia ego Dominus cum fuerint interfecti vestri in medio idolorum vestrorum in circuitu ararum vestrarum in omni colle excelso in cunctis summitatibus montium et subtus omne lignum nemorosum et subtus universam quercum frondosam locum ubi accenderunt tura redolentia universis idolis suis
EZEK|6|14|et extendam manum meam super eos et faciam terram desolatam et destitutam a deserto Deblatha in omnibus habitationibus eorum et scient quia ego Dominus
EZEK|7|1|et factus est sermo Domini ad me dicens
EZEK|7|2|et tu fili hominis haec dicit Dominus Deus terrae Israhel finis venit finis super quattuor plagas terrae
EZEK|7|3|nunc finis super te et emittam furorem meum in te et iudicabo te iuxta vias tuas et ponam contra te omnes abominationes tuas
EZEK|7|4|et non parcet oculus meus super te et non miserebor sed vias tuas ponam super te et abominationes tuae in medio tui erunt et scietis quia ego Dominus
EZEK|7|5|haec dicit Dominus Deus adflictio una adflictio ecce venit
EZEK|7|6|finis venit venit finis evigilavit adversum te ecce venit
EZEK|7|7|venit contractio super te qui habitas in terra venit tempus prope est dies occisionis et non gloriae montium
EZEK|7|8|nunc de propinquo effundam iram meam super te et conpleam furorem meum in te et iudicabo te iuxta vias tuas et inponam tibi omnia scelera tua
EZEK|7|9|et non parcet oculus meus neque miserebor sed vias tuas inponam tibi et abominationes tuae in medio tui erunt et scietis quia ego sum Dominus percutiens
EZEK|7|10|ecce dies ecce venit egressa est contractio floruit virga germinavit superbia
EZEK|7|11|iniquitas surrexit in virga impietatis non ex eis et non ex populo neque ex sonitu eorum et non erit requies in eis
EZEK|7|12|venit tempus adpropinquavit dies qui emit non laetetur et qui vendit non lugeat quia ira super omnem populum eius
EZEK|7|13|quia qui vendit ad id quod vendidit non revertetur et adhuc in viventibus vita eorum visio enim ad omnem multitudinem eius non regredietur et vir in iniquitate vitae suae non confortabitur
EZEK|7|14|canite tuba praeparentur omnes et non est qui vadat ad proelium ira enim mea super universum populum eius
EZEK|7|15|gladius foris pestis et fames intrinsecus qui in agro est gladio morietur et qui in civitate pestilentia et fame devorabuntur
EZEK|7|16|et salvabuntur qui fugerint ex eis et erunt in montibus quasi columbae convallium omnes trepidi unusquisque in iniquitate sua
EZEK|7|17|omnes manus dissolventur et omnia genua fluent aquis
EZEK|7|18|et accingent se ciliciis et operiet eos formido et in omni facie confusio et in universis capitibus eorum calvitium
EZEK|7|19|argentum eorum foris proicietur et aurum eorum in sterquilinium erit argentum eorum et aurum eorum non valebit liberare eos in die furoris Domini animam suam non saturabunt et ventres eorum non implebuntur quia scandalum iniquitatis eorum factum est
EZEK|7|20|et ornamentum monilium suorum in superbiam posuerunt et imagines abominationum suarum et simulacrorum fecerunt ex eo propter hoc dedi eis illud in inmunditiam
EZEK|7|21|et dabo illud in manus alienorum ad diripiendum et impiis terrae in praedam et contaminabunt illud
EZEK|7|22|et avertam faciem meam ab eis et violabunt arcanum meum et introibunt in illud emissarii et contaminabunt illud
EZEK|7|23|fac conclusionem quoniam terra plena est iudicio sanguinum et civitas plena iniquitate
EZEK|7|24|et adducam pessimos de gentibus et possidebunt domos eorum et quiescere faciam superbiam potentium et possidebunt sanctuaria eorum
EZEK|7|25|angustia superveniente requirent pacem et non erit
EZEK|7|26|conturbatio super conturbationem veniet et auditus super auditum et quaerent visionem de propheta et lex peribit a sacerdote et consilium a senioribus
EZEK|7|27|rex lugebit et princeps induetur maerore et manus populi terrae conturbabuntur secundum viam eorum faciam eis et secundum iudicia eorum iudicabo eos et scient quia ego Dominus
EZEK|8|1|et factum est in anno sexto in sexto mense in quinta mensis ego sedebam in domo mea et senes Iuda sedebant coram me et cecidit super me ibi manus Domini Dei
EZEK|8|2|et vidi et ecce similitudo quasi aspectus ignis ab aspectu lumborum eius et deorsum ignis et a lumbis eius et sursum quasi aspectus splendoris ut visio electri
EZEK|8|3|et emissa similitudo manus adprehendit me in cincinno capitis mei et elevavit me spiritus inter terram et caelum et adduxit in Hierusalem in visione Dei iuxta ostium interius quod respiciebat aquilonem ubi erat statutum idolum zeli ad provocandam aemulationem
EZEK|8|4|et ecce ibi gloria Dei Israhel secundum visionem quam videram in campo
EZEK|8|5|et dixit ad me fili hominis leva oculos tuos ad viam aquilonis et levavi oculos meos ad viam aquilonis et ecce ab aquilone portae altaris idolum zeli in ipso introitu
EZEK|8|6|et dixit ad me fili hominis putasne vides tu quid isti faciant abominationes magnas quas domus Israhel facit hic ut procul recedam a sanctuario meo et adhuc conversus videbis abominationes maiores
EZEK|8|7|et introduxit me ad ostium atrii et vidi et ecce foramen unum in pariete
EZEK|8|8|et dixit ad me fili hominis fode parietem et cum perfodissem parietem apparuit ostium unum
EZEK|8|9|et dixit ad me ingredere et vide abominationes pessimas quas isti faciunt hic
EZEK|8|10|et ingressus vidi et ecce omnis similitudo reptilium et animalium abominatio et universa idola domus Israhel depicta erant in pariete in circuitu per totum
EZEK|8|11|et septuaginta viri de senioribus domus Israhel et Hiezonias filius Saphan stabat in medio eorum stantium ante picturas et unusquisque habebat turibulum in manu sua et vapor nebulae de ture consurgebat
EZEK|8|12|et dixit ad me certe vides fili hominis quae seniores domus Israhel faciunt in tenebris unusquisque in abscondito cubiculi sui dicunt enim non videt Dominus nos dereliquit Dominus terram
EZEK|8|13|et dixit ad me adhuc conversus videbis abominationes maiores quas isti faciunt
EZEK|8|14|et introduxit me per ostium portae domus Domini quod respiciebat ad aquilonem et ecce ibi mulieres sedebant plangentes Adonidem
EZEK|8|15|et dixit ad me certe vidisti fili hominis adhuc conversus videbis abominationes maiores his
EZEK|8|16|et introduxit me in atrium domus Domini interius et ecce in ostio templi Domini inter vestibulum et altare quasi viginti quinque viri dorsa habentes contra templum Domini et facies ad orientem et adorabant ad ortum solis
EZEK|8|17|et dixit ad me certe vidisti fili hominis numquid leve est hoc domui Iuda ut facerent abominationes istas quas fecerunt hic quia replentes terram iniquitate conversi sunt ad inritandum me et ecce adplicant ramum ad nares suas
EZEK|8|18|ergo et ego faciam in furore non parcet oculus meus nec miserebor et cum clamaverint ad aures meas voce magna non exaudiam eos
EZEK|9|1|et clamavit in auribus meis voce magna dicens adpropinquaverunt visitationes urbis et unusquisque vas interfectionis habet in manu sua
EZEK|9|2|et ecce sex viri veniebant de via portae superioris quae respicit ad aquilonem et uniuscuiusque vas interitus in manu eius vir quoque unus in medio eorum vestitus lineis et atramentarium scriptoris ad renes eius et ingressi sunt et steterunt iuxta altare aereum
EZEK|9|3|et gloria Domini Israhel adsumpta est de cherub quae erat super eum ad limen domus et vocavit virum qui indutus erat lineis et atramentarium scriptoris habebat in lumbis suis
EZEK|9|4|et dixit Dominus ad eum transi per mediam civitatem in medio Hierusalem et signa thau super frontes virorum gementium et dolentium super cunctis abominationibus quae fiunt in medio eius
EZEK|9|5|et illis dixit audiente me transite per civitatem sequentes eum et percutite non parcat oculus vester neque misereamini
EZEK|9|6|senem adulescentulum et virginem parvulum et mulieres interficite usque ad internicionem omnem autem super quem videritis thau ne occidatis et a sanctuario meo incipite coeperunt ergo a viris senioribus qui erant ante faciem domus
EZEK|9|7|et dixit ad eos contaminate domum et implete atria interfectis egredimini et egressi sunt et percutiebant eos qui erant in civitate
EZEK|9|8|et caede conpleta remansi ego ruique super faciem meam et clamans aio heu heu heu Domine Deus ergone disperdes omnes reliquias Israhel effundens furorem tuum super Hierusalem
EZEK|9|9|et dixit ad me iniquitas domus Israhel et Iuda magna est nimis valde et repleta est terra sanguinibus et civitas repleta est aversione dixerunt enim dereliquit Dominus terram et Dominus non videt
EZEK|9|10|igitur et meus non parcet oculus neque miserebor viam eorum super caput eorum reddam
EZEK|9|11|et ecce vir qui indutus erat lineis qui habebat atramentarium in dorso suo respondit verbum dicens feci sicut praecepisti mihi
EZEK|10|1|et vidi et ecce in firmamento quod erat super caput cherubin quasi lapis sapphyrus quasi species similitudinis solii apparuit super ea
EZEK|10|2|et dixit ad virum qui indutus erat lineis et ait ingredere in medio rotarum quae sunt subtus cherub et imple manum tuam prunis ignis quae sunt inter cherubin et effunde super civitatem ingressusque est in conspectu meo
EZEK|10|3|cherubin autem stabant a dextris domus cum ingrederetur vir et nubes implevit atrium interius
EZEK|10|4|et elevata est gloria Domini desuper cherub ad limen domus et repleta est domus nube et atrium repletum est splendore gloriae Domini
EZEK|10|5|et sonitus alarum cherubin audiebatur usque ad atrium exterius quasi vox Dei omnipotentis loquentis
EZEK|10|6|cumque praecepisset viro qui indutus erat lineis dicens sume ignem de medio rotarum quae sunt inter cherubin ingressus ille stetit iuxta rotam
EZEK|10|7|et extendit cherub manum de medio cherubin ad ignem qui erat inter cherubin et sumpsit et dedit in manus eius qui indutus erat lineis qui accipiens egressus est
EZEK|10|8|et apparuit in cherubin similitudo manus hominis subtus pinnas eorum
EZEK|10|9|et vidi et ecce quattuor rotae iuxta cherubin rota una iuxta cherub unum et rota alia iuxta cherub unum species autem erat rotarum quasi visio lapidis chrysoliti
EZEK|10|10|et aspectus earum similitudo una quattuor quasi sit rota in medio rotae
EZEK|10|11|cumque ambularent in quattuor partes gradiebantur non revertebantur ambulantes sed ad locum ad quem ire declinabat quae prima erat sequebantur et ceterae nec convertebantur
EZEK|10|12|et omne corpus earum et colla et manus et pinnae et circuli plena erant oculis in circuitu quattuor rotarum
EZEK|10|13|et rotas istas vocavit volubiles audiente me
EZEK|10|14|quattuor autem facies habebat unum facies una facies cherub et facies secunda facies hominis et in tertio facies leonis et in quarto facies aquilae
EZEK|10|15|et elevata sunt cherubin ipsum est animal quod videram iuxta flumen Chobar
EZEK|10|16|cumque ambularent cherubin ibant pariter et rotae iuxta ea et cum levarent cherubin alas suas ut exaltarentur de terra non residebant rotae sed et ipsae iuxta erant
EZEK|10|17|stantibus illis stabant et cum elevatis elevabantur spiritus enim vitae erat in eis
EZEK|10|18|et egressa est gloria Domini a limine templi et stetit super cherubin
EZEK|10|19|et elevantia cherubin alas suas exaltata sunt a terra coram me et illis egredientibus rotae quoque subsecutae sunt et stetit in introitu portae domus Domini orientalis et gloria Dei Israhel erat super ea
EZEK|10|20|ipsum est animal quod vidi subter Deum Israhel iuxta fluvium Chobar et intellexi quia cherubin essent
EZEK|10|21|quattuor per quattuor vultus uni et quattuor alae uni et similitudo manus hominis sub alis eorum
EZEK|10|22|et similitudo vultuum eorum ipsi vultus quos videram iuxta fluvium Chobar et intuitus eorum et impetus singulorum ante faciem suam ingredi
EZEK|11|1|et elevavit me spiritus et introduxit me ad portam domus Domini orientalem quae respicit solis ortum et ecce in introitu portae viginti quinque viri et vidi in medio eorum Hiezoniam filium Azur et Pheltiam filium Banaiae principes populi
EZEK|11|2|dixitque ad me fili hominis hii viri qui cogitant iniquitatem et tractant consilium pessimum in urbe ista
EZEK|11|3|dicentes nonne dudum aedificatae sunt domus haec est lebes nos autem carnes
EZEK|11|4|idcirco vaticinare de eis vaticinare fili hominis
EZEK|11|5|et inruit in me spiritus Domini et dixit ad me loquere haec dicit Dominus sic locuti estis domus Israhel et cogitationes cordis vestri ego novi
EZEK|11|6|plurimos occidistis in urbe hac et implestis vias eius interfectis
EZEK|11|7|propterea haec dicit Dominus Deus interfecti vestri quos posuistis in medio eius hii sunt carnes et haec est lebes et educam vos de medio eius
EZEK|11|8|gladium metuistis et gladium inducam super vos ait Dominus Deus
EZEK|11|9|et eiciam vos de medio eius daboque vos in manu hostium et faciam in vobis iudicia
EZEK|11|10|gladio cadetis in finibus Israhel iudicabo vos et scietis quia ego Dominus
EZEK|11|11|haec non erit vobis in lebetem et vos non eritis in medio eius in carnes in finibus Israhel iudicabo vos
EZEK|11|12|et scietis quia ego Dominus qui in praeceptis meis non ambulastis et iudicia mea non fecistis sed iuxta iudicia gentium quae in circuitu vestro sunt estis operati
EZEK|11|13|et factum est cum prophetarem Pheltias filius Banaiae mortuus est et cecidi in faciem meam clamans voce magna et dixi heu heu heu Domine Deus consummationem tu facis reliquiarum Israhel
EZEK|11|14|et factum est verbum Domini ad me dicens
EZEK|11|15|fili hominis fratres tui fratres tui viri propinqui tui et omnis domus Israhel universi quibus dixerunt habitatores Hierusalem longe recedite a Domino nobis data est terra in possessionem
EZEK|11|16|propterea haec dicit Dominus Deus quia longe feci eos in gentibus et quia dispersi eos in terris ero eis in sanctificationem modicam in terris ad quas venerunt
EZEK|11|17|propterea loquere haec dicit Dominus Deus congregabo vos de populis et adunabo de terris in quibus dispersi estis daboque vobis humum Israhel
EZEK|11|18|et ingredientur illuc et auferent omnes offensiones cunctasque abominationes eius de illa
EZEK|11|19|et dabo eis cor unum et spiritum novum tribuam in visceribus eorum et auferam cor lapideum de carne eorum et dabo eis cor carneum
EZEK|11|20|ut in praeceptis meis ambulent et iudicia mea custodiant faciantque ea et sint mihi in populum et ego sim eis in Deum
EZEK|11|21|quorum cor post offendicula et abominationes suas ambulat horum viam in capite suo ponam dicit Dominus Deus
EZEK|11|22|et elevaverunt cherubin alas suas et rotae cum eis et gloria Dei Israhel erat super ea
EZEK|11|23|et ascendit gloria Domini de medio civitatis stetitque super montem qui est ad orientem urbis
EZEK|11|24|et spiritus levavit me adduxitque in Chaldeam ad transmigrationem in visione in spiritu Dei et sublata est a me visio quam videram
EZEK|11|25|et locutus sum ad transmigrationem omnia verba Domini quae ostenderat mihi
EZEK|12|1|et factus est sermo Domini ad me dicens
EZEK|12|2|fili hominis in medio domus exasperantis tu habitas qui oculos habent ad videndum et non vident et aures ad audiendum et non audiunt quia domus exasperans est
EZEK|12|3|tu ergo fili hominis fac tibi vasa transmigrationis et transmigrabis per diem coram eis transmigrabis autem de loco tuo ad locum alterum in conspectu eorum si forte aspiciant quia domus exasperans est
EZEK|12|4|et efferes foras vasa tua quasi vasa transmigrantis per diem in conspectu eorum tu autem egredieris vespere coram eis sicut egreditur migrans
EZEK|12|5|ante oculos eorum perfodi tibi parietem et egredieris per eum
EZEK|12|6|in conspectu eorum in umeris portaberis in caligine effereris faciem tuam velabis et non videbis terram quia portentum dedi te domui Israhel
EZEK|12|7|feci ergo sicut praeceperat mihi vasa mea protuli quasi vasa transmigrantis per diem et vespere perfodi mihi parietem manu in caligine egressus sum et in umeris portatus in conspectu eorum
EZEK|12|8|et factus est sermo Domini ad me mane dicens
EZEK|12|9|fili hominis numquid non dixerunt ad te domus Israhel domus exasperans quid tu facis
EZEK|12|10|dic ad eos haec dicit Dominus Deus super ducem onus istud qui est in Hierusalem et super omnem domum Israhel quae est in medio eorum
EZEK|12|11|dic ego portentum vestrum quomodo feci sic fiet illis in transmigrationem et captivitatem ibunt
EZEK|12|12|et dux qui est in medio eorum in umeris portabitur in caligine egredietur parietem perfodient ut educant eum facies eius operietur ut non videat oculo terram
EZEK|12|13|et extendam rete meum super illum et capietur in sagena mea et adducam eum in Babylonem in terram Chaldeorum et ipsam non videbit ibique morietur
EZEK|12|14|et omnes qui circa eum sunt praesidium eius et agmina eius dispergam in omnem ventum et gladium evaginabo post eos
EZEK|12|15|et scient quia ego Dominus quando dispersero illos in gentibus et disseminavero eos in terris
EZEK|12|16|et relinquam ex eis viros paucos a gladio et fame et pestilentia ut narrent omnia scelera eorum in gentibus ad quas ingredientur et scient quia ego Dominus
EZEK|12|17|et factus est sermo Domini ad me dicens
EZEK|12|18|fili hominis panem tuum in conturbatione comede sed et aquam tuam in festinatione et maerore bibe
EZEK|12|19|et dices ad populum terrae haec dicit Dominus Deus ad eos qui habitant in Hierusalem in terra Israhel panem suum in sollicitudine comedent et aquam suam in desolatione bibent ut desoletur terra a multitudine sua propter iniquitatem omnium qui habitant in ea
EZEK|12|20|et civitates quae nunc habitantur desolatae erunt terraque deserta et scietis quia ego Dominus
EZEK|12|21|et factus est sermo Domini ad me dicens
EZEK|12|22|fili hominis quod est proverbium istud vobis in terra Israhel dicentium in longum differentur dies et peribit omnis visio
EZEK|12|23|ideo dic ad eos haec dicit Dominus Deus quiescere faciam proverbium istud neque vulgo dicetur ultra in Israhel et loquere ad eos quod adpropinquaverint dies et sermo omnis visionis
EZEK|12|24|non enim erit ultra omnis visio cassa neque divinatio ambigua in medio filiorum Israhel
EZEK|12|25|quia ego Dominus loquar quodcumque locutus fuero verbum et fiet non prolongabitur amplius sed in diebus vestris domus exasperans loquar verbum et faciam illud dicit Dominus Deus
EZEK|12|26|et factus est sermo Domini ad me dicens
EZEK|12|27|fili hominis ecce domus Israhel dicentium visio quam hic videt in dies multos et in tempora longa iste prophetat
EZEK|12|28|propterea dic ad eos haec dicit Dominus Deus non prolongabitur ultra omnis sermo meus verbum quod locutus fuero conplebitur dicit Dominus Deus
EZEK|13|1|et factus est sermo Domini ad me dicens
EZEK|13|2|fili hominis vaticinare ad prophetas Israhel qui prophetant et dices prophetantibus de corde suo audite verbum Domini
EZEK|13|3|haec dicit Dominus Deus vae prophetis insipientibus qui sequuntur spiritum suum et nihil vident
EZEK|13|4|quasi vulpes in desertis prophetae tui Israhel erant
EZEK|13|5|non ascendistis ex adverso neque opposuistis murum pro domo Israhel ut staretis in proelio in die Domini
EZEK|13|6|vident vana et divinant mendacium dicentes ait Dominus cum Dominus non miserit eos et perseveraverunt confirmare sermonem
EZEK|13|7|numquid non visionem cassam vidistis et divinationem mendacem locuti estis et dicitis ait Dominus cum ego non sim locutus
EZEK|13|8|propterea haec dicit Dominus Deus quia locuti estis vana et vidistis mendacium ideo ecce ego ad vos ait Dominus Deus
EZEK|13|9|et erit manus mea super prophetas qui vident vana et divinant mendacium in concilio populi mei non erunt et in scriptura domus Israhel non scribentur nec in terra Israhel ingredientur et scietis quia ego Dominus Deus
EZEK|13|10|eo quod deceperint populum meum dicentes pax et non est pax et ipse aedificabat parietem illi autem liniebant eum luto absque paleis
EZEK|13|11|dic ad eos qui liniunt absque temperatura quod casurus sit erit enim imber inundans et dabo lapides praegrandes desuper inruentes et ventum procellae dissipantem
EZEK|13|12|siquidem ecce cecidit paries numquid non dicetur vobis ubi est litura quam levistis
EZEK|13|13|propterea haec dicit Dominus Deus et erumpere faciam spiritum tempestatum in indignatione mea et imber inundans in furore meo erit et lapides grandes in ira in consummationem
EZEK|13|14|et destruam parietem quem levistis absque temperamento et adaequabo eum terrae et revelabitur fundamentum eius et cadet et consumetur in medio eius et scietis quia ego sum Dominus
EZEK|13|15|et conplebo indignationem meam in parietem et in his qui linunt eum absque temperamento dicamque vobis non est paries et non sunt qui linunt eum
EZEK|13|16|prophetae Israhel qui prophetant ad Hierusalem et vident ei visionem pacis et non est pax ait Dominus Deus
EZEK|13|17|et tu fili hominis pone faciem tuam contra filias populi tui quae prophetant de corde suo et vaticinare super eas
EZEK|13|18|et dic haec ait Dominus Deus vae quae consuunt pulvillos sub omni cubito manus et faciunt cervicalia sub capite universae aetatis ad capiendas animas cum caperent animas populi mei vivificabant animas eorum
EZEK|13|19|et violabant me ad populum meum propter pugillum hordei et fragmen panis ut interficerent animas quae non moriuntur et vivificarent animas quae non vivunt mentientes populo meo credenti mendaciis
EZEK|13|20|propter hoc haec dicit Dominus Deus ecce ego ad pulvillos vestros quibus vos capitis animas volantes et disrumpam eos de brachiis vestris et dimittam animas quas vos capitis animas ad volandum
EZEK|13|21|et disrumpam cervicalia vestra et liberabo populum meum de manu vestra neque erunt ultra in manibus vestris ad praedandum et scietis quia ego Dominus
EZEK|13|22|pro eo quod maerere fecistis cor iusti mendaciter quem ego non contristavi et confortastis manus impii ut non reverteretur a via sua mala et viveret
EZEK|13|23|propterea vana non videbitis et divinationes non divinabitis amplius et eruam populum meum de manu vestra et scietis quoniam ego Dominus
EZEK|14|1|et venerunt ad me viri seniorum Israhel et sederunt coram me
EZEK|14|2|et factus est sermo Domini ad me dicens
EZEK|14|3|fili hominis viri isti posuerunt inmunditias suas in cordibus suis et scandalum iniquitatis suae statuerunt contra faciem suam numquid interrogatus respondebo eis
EZEK|14|4|propter hoc loquere eis et dices ad eos haec dicit Dominus Deus homo homo de domo Israhel qui posuerit inmunditias suas in corde suo et scandalum iniquitatis suae statuerit contra faciem suam et venerit ad prophetam interrogans per eum me ego Dominus respondebo ei in multitudine inmunditiarum suarum
EZEK|14|5|ut capiatur domus Israhel in corde suo quo recesserunt a me in cunctis idolis suis
EZEK|14|6|propterea dic ad domum Israhel haec dicit Dominus Deus convertimini et recedite ab idolis vestris et ab universis contaminationibus vestris avertite facies vestras
EZEK|14|7|quia homo homo de domo Israhel et de proselytis quicumque advena fuerit in Israhel si alienatus fuerit a me et posuerit idola sua in corde suo et scandalum iniquitatis suae statuerit contra faciem suam et venerit ad prophetam ut interroget per eum me ego Dominus respondebo ei per me
EZEK|14|8|et ponam faciem meam super hominem illum et faciam eum in exemplum et in proverbium et disperdam eum de medio populi mei et scietis quia ego Dominus
EZEK|14|9|et propheta cum erraverit et locutus fuerit verbum ego Dominus decepi prophetam illum et extendam manum meam super eum et delebo eum de medio populi mei Israhel
EZEK|14|10|et portabunt iniquitatem suam iuxta iniquitatem interrogantis sic iniquitas prophetae erit
EZEK|14|11|ut non erret ultra domus Israhel a me neque polluatur in universis praevaricationibus suis sed sit mihi in populum et ego sim eis in Deum ait Dominus exercituum
EZEK|14|12|et factus est sermo Domini ad me dicens
EZEK|14|13|fili hominis terra cum peccaverit mihi ut praevaricetur praevaricans extendam manum meam super eam et conteram virgam panis eius et inmittam in eam famem et interficiam de ea hominem et iumentum
EZEK|14|14|et si fuerint tres viri isti in medio eius Noe Danihel et Iob ipsi iustitia sua liberabunt animas suas ait Dominus exercituum
EZEK|14|15|quod si et bestias pessimas induxero super terram ut vastem eam et fuerit invia eo quod non sit pertransiens propter bestias
EZEK|14|16|tres viri isti qui fuerint in ea vivo ego dicit Dominus Deus quia nec filios nec filias liberabunt sed ipsi soli liberabuntur terra autem desolabitur
EZEK|14|17|vel si gladium induxero super terram illam et dixero gladio transi per terram et interfecero de ea hominem et iumentum
EZEK|14|18|et tres viri isti fuerint in medio eius vivo ego dicit Dominus Deus non liberabunt filios neque filias sed ipsi soli liberabuntur
EZEK|14|19|si autem et pestilentiam inmisero super terram illam et effudero indignationem meam super eam in sanguine ut auferam ex ea hominem et iumentum
EZEK|14|20|et Noe et Danihel et Iob fuerint in medio eius vivo ego dicit Dominus Deus quia filium et filiam non liberabunt sed ipsi iustitia sua liberabunt animas suas
EZEK|14|21|quoniam haec dicit Dominus Deus quod si et quattuor iudicia mea pessima gladium et famem et bestias malas et pestilentiam misero in Hierusalem ut interficiam de ea hominem et pecus
EZEK|14|22|tamen relinquetur in ea salvatio educentium filios et filias ecce ipsi egredientur ad vos et videbitis viam eorum et adinventiones eorum et consolabimini super malo quod induxi in Hierusalem in omnibus quae inportavi super eam
EZEK|14|23|et consolabuntur vos cum videritis viam eorum et adinventiones eorum et cognoscetis quod non frustra fecerim omnia quae feci in ea ait Dominus Deus
EZEK|15|1|et factus est sermo Domini ad me dicens
EZEK|15|2|fili hominis quid fiet ligno vitis ex omnibus lignis nemorum quae sunt inter ligna silvarum
EZEK|15|3|numquid tolletur de ea lignum ut fiat opus aut fabricabitur de ea paxillus ut dependeat in eo quodcumque vas
EZEK|15|4|ecce igni datum est in escam utramque partem eius consumpsit ignis et medietas eius redacta est in favillam numquid utile erit ad opus
EZEK|15|5|etiam cum esset integrum non erat aptum ad opus quanto magis cum ignis illud devoraverit et conbuserit nihil ex eo fiet operis
EZEK|15|6|propterea haec dicit Dominus Deus quomodo lignum vitis inter ligna silvarum quod dedi igni ad devorandum sic tradidi habitatores Hierusalem
EZEK|15|7|et ponam faciem meam in eos de igne egredientur et ignis consumet eos et scietis quia ego Dominus cum posuero faciem meam in eos
EZEK|15|8|et dedero terram inviam et desolatam eo quod praevaricatores extiterint dicit Dominus Deus
EZEK|16|1|et factus est sermo Domini ad me dicens
EZEK|16|2|fili hominis notas fac Hierusalem abominationes suas
EZEK|16|3|et dices haec dicit Dominus Deus Hierusalem radix tua et generatio tua de terra chananea pater tuus Amorreus et mater tua Cetthea
EZEK|16|4|et quando nata es in die ortus tui non est praecisus umbilicus tuus et in aqua non es lota in salutem nec sale salita nec involuta pannis
EZEK|16|5|non pepercit super te oculus ut facerem tibi unum de his miseratus tui sed proiecta es super faciem terrae in abiectione animae tuae in die qua nata es
EZEK|16|6|transiens autem per te vidi te conculcari in sanguine tuo et dixi tibi cum esses in sanguine tuo vive dixi inquam tibi in sanguine tuo vive
EZEK|16|7|multiplicatam quasi germen agri dedi te et multiplicata es et grandis effecta et ingressa es et pervenisti ad mundum muliebrem ubera tua intumuerunt et pilus tuus germinavit et eras nuda et confusionis plena
EZEK|16|8|et transivi per te et vidi te et ecce tempus tuum tempus amantium et expandi amictum meum super te et operui ignominiam tuam et iuravi tibi et ingressus sum pactum tecum ait Dominus Deus et facta es mihi
EZEK|16|9|et lavi te aqua et emundavi sanguinem tuum ex te et unxi te oleo
EZEK|16|10|et vestivi te discoloribus et calciavi te ianthino et cinxi te bysso et indui te subtilibus
EZEK|16|11|et ornavi te ornamento et dedi armillas in manibus tuis et torquem circa collum tuum
EZEK|16|12|et dedi inaurem super os tuum et circulos auribus tuis et coronam decoris in capite tuo
EZEK|16|13|et ornata es auro et argento et vestita es bysso et polymito et multicoloribus similam et mel et oleum comedisti et decora facta es vehementer nimis et profecisti in regnum
EZEK|16|14|et egressum est nomen tuum in gentes propter speciem tuam quia perfecta eras in decore meo quem posueram super te dicit Dominus Deus
EZEK|16|15|et habens fiduciam in pulchritudine tua fornicata es in nomine tuo et exposuisti fornicationem tuam omni transeunti ut eius fieres
EZEK|16|16|et sumens de vestimentis meis fecisti tibi excelsa hinc inde consuta et fornicata es super eis sicut non est factum neque futurum est
EZEK|16|17|et tulisti vasa decoris tui de auro meo et argento meo quae dedi tibi et fecisti tibi imagines masculinas et fornicata es in eis
EZEK|16|18|et sumpsisti vestimenta tua multicoloria et vestita es eis et oleum meum et thymiama meum posuisti coram eis
EZEK|16|19|et panem meum quem dedi tibi similam et oleum et mel quibus enutrivi te posuisti in conspectu eorum in odorem suavitatis et factum est ait Dominus Deus
EZEK|16|20|et tulisti filios tuos et filias tuas quas generasti mihi et immolasti eis ad devorandum numquid parva est fornicatio tua
EZEK|16|21|immolantis filios meos et dedisti illos consecrans eis
EZEK|16|22|et post omnes abominationes tuas et fornicationes non es recordata dierum adulescentiae tuae quando eras nuda et confusione plena conculcata in sanguine tuo
EZEK|16|23|et accidit post omnem malitiam tuam vae vae tibi ait Dominus Deus
EZEK|16|24|et aedificasti tibi lupanar et fecisti tibi prostibulum in cunctis plateis
EZEK|16|25|ad omne caput viae aedificasti signum prostitutionis tuae et abominabilem fecisti decorem tuum et divisisti pedes tuos omni transeunti et multiplicasti fornicationes tuas
EZEK|16|26|et fornicata es cum filiis Aegypti vicinis tuis magnarum carnium et multiplicasti fornicationem tuam ad inritandum me
EZEK|16|27|ecce ego extendi manum meam super te et auferam ius tuum et dabo te in animam odientium te filiarum Palestinarum quae erubescunt in via tua scelerata
EZEK|16|28|et fornicata es in filiis Assyriorum eo quod necdum fueris expleta et postquam fornicata es nec sic es satiata
EZEK|16|29|et multiplicasti fornicationem tuam in terra Chanaan cum Chaldeis et nec sic satiata es
EZEK|16|30|in quo mundabo cor tuum ait Dominus Deus cum facias omnia haec opera mulieris meretricis et procacis
EZEK|16|31|quia fabricasti lupanar tuum in capite omnis viae et excelsum tuum fecisti in omni platea nec facta es quasi meretrix fastidio augens pretium
EZEK|16|32|sed quasi mulier adultera quae super virum suum inducit alienos
EZEK|16|33|omnibus meretricibus dantur mercedes tu autem dedisti mercedes cunctis amatoribus tuis et donabas eis ut intrarent ad te undique ad fornicandum tecum
EZEK|16|34|factumque in te est contra consuetudinem mulierum in fornicationibus tuis et post te non erit fornicatio in eo enim quod dedisti mercedes et mercedes non accepisti factum est in te contrarium
EZEK|16|35|propterea meretrix audi verbum Domini
EZEK|16|36|haec dicit Dominus Deus quia effusum est aes tuum et revelata est ignominia tua in fornicationibus tuis super amatores tuos et super idola abominationum tuarum in sanguine filiorum tuorum quos dedisti eis
EZEK|16|37|ecce ego congregabo omnes amatores tuos quibus commixta es et omnes quos dilexisti cum universis quos oderas et congregabo eos super te undique et nudabo ignominiam tuam coram eis et videbunt omnem turpitudinem tuam
EZEK|16|38|et iudicabo te iudiciis adulterarum et effundentium sanguinem et dabo te in sanguinem furoris et zeli
EZEK|16|39|et dabo te in manus eorum et destruent lupanar tuum et demolientur prostibulum tuum et denudabunt te vestimentis tuis et auferent vasa decoris tui et derelinquent te nudam plenamque ignominia
EZEK|16|40|et adducent super te multitudinem et lapidabunt te lapidibus et trucidabunt te gladiis suis
EZEK|16|41|et conburent domos tuas igni et facient in te iudicia in oculis mulierum plurimarum et desines fornicari et mercedes ultra non dabis
EZEK|16|42|et requiescet indignatio mea in te et auferetur zelus meus a te et quiescam nec irascar amplius
EZEK|16|43|eo quod non fueris recordata dierum adulescentiae tuae et provocasti me in omnibus his quapropter et ego vias tuas in capite tuo dedi ait Dominus Deus et non feci iuxta scelera tua in omnibus abominationibus tuis
EZEK|16|44|ecce omnis qui dicit vulgo proverbium in te adsumet illud dicens sicut mater ita et filia eius
EZEK|16|45|filia matris tuae es tu quae proiecit virum suum et filios suos et soror sororum tuarum tu quae proiecerunt viros suos et filios suos mater vestra Cetthea et pater vester Amorreus
EZEK|16|46|et soror tua maior Samaria ipsa et filiae eius quae habitat ad sinistram tuam soror autem tua minor te quae habitat a dextris tuis Sodoma et filiae eius
EZEK|16|47|sed nec in viis earum ambulasti neque secundum scelera earum fecisti pauxillum minus paene sceleratiora fecisti illis in omnibus viis tuis
EZEK|16|48|vivo ego dicit Dominus Deus quia non fecit Sodoma soror tua ipsa et filiae eius sicut fecisti tu et filiae tuae
EZEK|16|49|ecce haec fuit iniquitas Sodomae sororis tuae superbia saturitas panis et abundantia et otium ipsius et filiarum eius et manum egeno et pauperi non porrigebant
EZEK|16|50|et elevatae sunt et fecerunt abominationes coram me et abstuli eas sicut vidisti
EZEK|16|51|et Samaria dimidium peccatorum tuorum non peccavit sed vicisti eas sceleribus tuis et iustificasti sorores tuas in omnibus abominationibus tuis quas operata es
EZEK|16|52|ergo et tu porta confusionem tuam quae vicisti sorores tuas peccatis tuis sceleratius agens ab eis iustificatae sunt enim a te ergo et tu confundere et porta ignominiam tuam quae iustificasti sorores tuas
EZEK|16|53|et convertam restituens eas conversione Sodomorum cum filiabus suis et conversione Samariae et filiarum eius et convertam reversionem tuam in medio earum
EZEK|16|54|ut portes ignominiam tuam et confundaris in omnibus quae fecisti consolans eas
EZEK|16|55|et soror tua Sodoma et filiae eius revertentur ad antiquitatem suam et Samaria et filiae eius revertentur ad antiquitatem suam et tu et filiae tuae revertimini ad antiquitatem vestram
EZEK|16|56|non fuit autem Sodoma soror tua audita in ore tuo in die superbiae tuae
EZEK|16|57|antequam revelaretur malitia tua sicut hoc tempore in obprobrium filiarum Syriae et cunctarum in circuitu tuo filiarum Palestinarum quae ambiunt te per gyrum
EZEK|16|58|scelus tuum et ignominiam tuam tu portasti ait Dominus Deus
EZEK|16|59|quia haec dicit Dominus Deus et faciam tibi sicut dispexisti iuramentum ut irritum faceres pactum
EZEK|16|60|et recordabor ego pacti mei tecum in diebus adulescentiae tuae et suscitabo tibi pactum sempiternum
EZEK|16|61|et recordaberis viarum tuarum et confunderis cum receperis sorores tuas te maiores cum minoribus tuis et dabo eas tibi in filias sed non ex pacto tuo
EZEK|16|62|et suscitabo ego pactum meum tecum et scies quia ego Dominus
EZEK|16|63|ut recorderis et confundaris et non sit tibi ultra aperire os prae confusione tua cum placatus fuero tibi in omnibus quae fecisti ait Dominus Deus
EZEK|17|1|et factum est verbum Domini ad me dicens
EZEK|17|2|fili hominis propone enigma et narra parabolam ad domum Israhel
EZEK|17|3|et dices haec dicit Dominus Deus aquila grandis magnarum alarum longo membrorum ductu plena plumis et varietate venit ad Libanum et tulit medullam cedri
EZEK|17|4|summitatem frondium eius avellit et transportavit eam in terram Chanaan in urbem negotiatorum posuit illam
EZEK|17|5|et tulit de semente terrae et posuit illud in terra pro semine ut firmaret radicem super aquas multas in superficie posuit illud
EZEK|17|6|cumque germinasset crevit in vineam latiorem humili statura respicientibus ramis eius ad eam et radices eius sub illa erunt facta est ergo vinea et fructificavit in palmites et emisit propagines
EZEK|17|7|et facta est aquila altera grandis magnis alis multisque plumis et ecce vinea ista quasi mittens radices suas ad eam palmites suos extendit ad illam ut inrigaret eam de areolis germinis sui
EZEK|17|8|in terra bona super aquas multas plantata est ut faciat frondes et portet fructum et sit in vineam grandem
EZEK|17|9|dic haec dicit Dominus Deus ergone prosperabitur nonne radices eius evellet et fructum eius distringet et siccabit omnes palmites germinis eius et arescet et non in brachio grandi neque in populo multo ut evelleret eam radicitus
EZEK|17|10|ecce plantata est ergone prosperabitur nonne cum tetigerit eam ventus urens siccabitur et in areis germinis sui arescet
EZEK|17|11|et factum est verbum Domini ad me dicens
EZEK|17|12|dic ad domum exasperantem nescitis quid ista significent dic ecce venit rex Babylonis Hierusalem et adsumet regem et principes eius et adducet eos ad semet ipsum in Babylonem
EZEK|17|13|et tollet de semine regni ferietque cum eo foedus et accipiet ab eo iusiurandum sed et fortes terrae tollet
EZEK|17|14|ut sit regnum humile et non elevetur sed custodiat pactum eius et servet illud
EZEK|17|15|qui recedens ab eo misit nuntios ad Aegyptum ut daret sibi equos et populum multum numquid prosperabitur vel consequetur salutem qui fecit haec et qui dissolvit pactum numquid effugiet
EZEK|17|16|vivo ego dicit Dominus Deus quoniam in loco regis qui constituit eum regem cuius fecit irritum iuramentum et solvit pactum quod habebat cum eo in medio Babylonis morietur
EZEK|17|17|et non in exercitu grandi neque in populo multo faciet contra eum Pharao proelium in iactu aggeris et in extructione vallorum ut interficiat animas multas
EZEK|17|18|spreverat enim iuramentum ut solveret foedus et ecce dedit manum suam et cum omnia haec fecerit non effugiet
EZEK|17|19|propterea haec dicit Dominus Deus vivo ego quoniam iuramentum quod sprevit et foedus quod praevaricatus est ponam in caput eius
EZEK|17|20|et expandam super eum rete meum et conprehendetur sagena mea et adducam eum in Babylonem et iudicabo illum ibi in praevaricatione qua despexit me
EZEK|17|21|et omnes profugi eius cum universo agmine gladio cadent residui autem in omnem ventum dispergentur et scietis quia ego Dominus locutus sum
EZEK|17|22|haec dicit Dominus Deus et sumam ego de medulla cedri sublimis et ponam de vertice ramorum eius tenerum distringam et plantabo super montem excelsum et eminentem
EZEK|17|23|in monte sublimi Israhel plantabo illud et erumpet in germen et faciet fructum et erit in cedrum magnam et habitabunt sub eo omnes volucres universum volatile sub umbra frondium eius nidificabit
EZEK|17|24|et scient omnia ligna regionis quia ego Dominus humiliavi lignum sublime et exaltavi lignum humile et siccavi lignum viride et frondere feci lignum aridum ego Dominus locutus sum et feci
EZEK|18|1|et factus est sermo Domini ad me dicens
EZEK|18|2|quid est quod inter vos parabolam vertitis in proverbium istud in terra Israhel dicentes patres comederunt uvam acerbam et dentes filiorum obstupescunt
EZEK|18|3|vivo ego dicit Dominus Deus si erit vobis ultra parabola haec in proverbium in Israhel
EZEK|18|4|ecce omnes animae meae sunt ut anima patris ita et anima filii mea est anima quae peccaverit ipsa morietur
EZEK|18|5|et vir si fuerit iustus et fecerit iudicium et iustitiam
EZEK|18|6|in montibus non comederit et oculos suos non levaverit ad idola domus Israhel et uxorem proximi sui non violaverit et ad mulierem menstruatam non accesserit
EZEK|18|7|et hominem non contristaverit pignus debitori reddiderit per vim nihil rapuerit panem suum esurienti dederit et nudum operuerit vestimento
EZEK|18|8|ad usuram non commodaverit et amplius non acceperit ab iniquitate averterit manum suam iudicium verum fecerit inter virum et virum
EZEK|18|9|in praeceptis meis ambulaverit et iudicia mea custodierit ut faciat veritatem hic iustus est vita vivet ait Dominus Deus
EZEK|18|10|quod si genuerit filium latronem effundentem sanguinem et fecerit unum de istis
EZEK|18|11|et haec quidem omnia non facientem sed in montibus comedentem et uxorem proximi sui polluentem
EZEK|18|12|egenum et pauperem contristantem rapientem rapinas pignus non reddentem et ad idola levantem oculos suos abominationem facientem
EZEK|18|13|ad usuram dantem et amplius accipientem numquid vivet non vivet cum universa detestanda haec fecerit morte morietur sanguis eius in ipso erit
EZEK|18|14|quod si genuerit filium qui videns omnia peccata patris sui quae fecit timuerit et non fecerit simile eis
EZEK|18|15|super montes non comederit et oculos suos non levaverit ad idola domus Israhel et uxorem proximi sui non violaverit
EZEK|18|16|et virum non contristaverit pignus non retinuerit et rapinam non rapuerit panem suum esurienti dederit et nudum operuerit vestimento
EZEK|18|17|a pauperis iniuria averterit manum suam usuram et superabundantiam non acceperit iudicia mea fecerit in praeceptis meis ambulaverit hic non morietur in iniquitate patris sui sed vita vivet
EZEK|18|18|pater eius quia calumniatus est et vim fecit fratri et malum operatus est in medio populi sui ecce mortuus est in iniquitate sua
EZEK|18|19|et dicitis quare non portavit filius iniquitatem patris videlicet quia filius iudicium et iustitiam operatus est omnia praecepta mea custodivit et fecit illa vita vivet
EZEK|18|20|anima quae peccaverit ipsa morietur filius non portabit iniquitatem patris et pater non portabit iniquitatem filii iustitia iusti super eum erit et impietas impii erit super eum
EZEK|18|21|si autem impius egerit paenitentiam ab omnibus peccatis suis quae operatus est et custodierit universa praecepta mea et fecerit iudicium et iustitiam vita vivet non morietur
EZEK|18|22|omnium iniquitatum eius quas operatus est non recordabor in iustitia sua quam operatus est vivet
EZEK|18|23|numquid voluntatis meae est mors impii dicit Dominus Deus et non ut convertatur a viis suis et vivat
EZEK|18|24|si autem averterit se iustus a iustitia sua et fecerit iniquitatem secundum omnes abominationes quas operari solet impius numquid vivet omnes iustitiae eius quas fecerat non recordabuntur in praevaricatione qua praevaricatus est et in peccato suo quod peccavit in ipsis morietur
EZEK|18|25|et dixistis non est aequa via Domini audite domus Israhel numquid via mea non est aequa et non magis viae vestrae pravae sunt
EZEK|18|26|cum enim averterit se iustus a iustitia sua et fecerit iniquitatem morietur in eis in iniustitia quam operatus est morietur
EZEK|18|27|et cum averterit se impius ab impietate sua quam operatus est et fecerit iudicium et iustitiam ipse animam suam vivificabit
EZEK|18|28|considerans enim et avertens se ab omnibus iniquitatibus suis quas operatus est vita vivet et non morietur
EZEK|18|29|et dicunt filii Israhel non est aequa via Domini numquid viae meae non sunt aequae domus Israhel et non magis viae vestrae pravae
EZEK|18|30|idcirco unumquemque iuxta vias suas iudicabo domus Israhel ait Dominus Deus convertimini et agite paenitentiam ab omnibus iniquitatibus vestris et non erit vobis in ruinam iniquitas
EZEK|18|31|proicite a vobis omnes praevaricationes vestras in quibus praevaricati estis et facite vobis cor novum et spiritum novum et quare moriemini domus Israhel
EZEK|18|32|quia nolo mortem morientis dicit Dominus Deus revertimini et vivite
EZEK|19|1|et tu adsume planctum super principes Israhel
EZEK|19|2|et dices quare mater tua leaena inter leones cubavit in medio leunculorum enutrivit catulos suos
EZEK|19|3|et eduxit unum de leunculis suis leo factus est et didicit capere praedam hominemque comedere
EZEK|19|4|et audierunt de eo gentes et non absque vulneribus suis ceperunt eum et adduxerunt eum in catenis in terram Aegypti
EZEK|19|5|quae cum vidisset quoniam infirmata est et periit expectatio eius tulit unum de leunculis suis leonem constituit eum
EZEK|19|6|qui incedebat inter leones et factus est leo didicit praedam capere et homines devorare
EZEK|19|7|didicit viduas facere et civitates eorum in desertum adducere et desolata est terra et plenitudo eius a voce rugitus illius
EZEK|19|8|et convenerunt adversum eum gentes undique de provinciis et expanderunt super eum rete suum in vulneribus earum captus est
EZEK|19|9|et miserunt eum in caveam in catenis adduxerunt eum ad regem Babylonis miseruntque eum in carcerem ne audiretur vox eius ultra super montes Israhel
EZEK|19|10|mater tua quasi vinea in sanguine tuo super aquam plantata fructus eius et frondes eius creverunt ex aquis multis
EZEK|19|11|et factae sunt ei virgae solidae in sceptra dominantium et exaltata est statura eius inter frondes et vidit altitudinem suam in multitudine palmitum suorum
EZEK|19|12|et evulsa est in ira in terramque proiecta et ventus urens siccavit fructum eius marcuerunt et arefactae sunt virgae roboris eius ignis comedit eam
EZEK|19|13|et nunc transplantata est in desertum in terra invia et sitienti
EZEK|19|14|et egressus est ignis de virga ramorum eius qui fructum eius comedit et non fuit in ea virga fortis sceptrum dominantium planctus est et erit in planctum
EZEK|20|1|et factum est in anno septimo in quinto mense in decima mensis venerunt viri de senioribus Israhel ut interrogarent Dominum et sederunt coram me
EZEK|20|2|et factus est sermo Domini ad me dicens
EZEK|20|3|fili hominis loquere senioribus Israhel et dices ad eos haec dicit Dominus Deus num ad interrogandum me vos venistis vivo ego quia non respondebo vobis ait Dominus Deus
EZEK|20|4|si iudicas eos si iudicas fili hominis abominationes patrum eorum ostende eis
EZEK|20|5|et dices ad eos haec dicit Dominus Deus in die qua elegi Israhel et levavi manum meam pro stirpe domus Iacob et apparui eis in terra Aegypti et levavi manum meam pro eis dicens ego Dominus Deus vester
EZEK|20|6|in die illa levavi manum meam pro eis ut educerem eos de terra Aegypti in terram quam provideram eis fluentem lacte et melle quae est egregia inter omnes terras
EZEK|20|7|et dixi ad eos unusquisque offensiones oculorum suorum abiciat et in idolis Aegypti nolite pollui ego Dominus Deus vester
EZEK|20|8|et inritaverunt me nolueruntque audire unusquisque abominationes oculorum suorum non proiecit nec idola Aegypti reliquerunt et dixi ut effunderem indignationem meam super eos et implerem iram meam in eis in medio terrae Aegypti
EZEK|20|9|et feci propter nomen meum ut non violaretur coram gentibus in quarum medio erant et inter quas apparui eis ut educerem eos de terra Aegypti
EZEK|20|10|eieci ergo eos de terra Aegypti et eduxi in desertum
EZEK|20|11|et dedi eis praecepta mea et iudicia mea ostendi eis quae faciat homo et vivat in eis
EZEK|20|12|insuper et sabbata mea dedi eis ut esset signum inter me et eos et scirent quia ego Dominus sanctificans eos
EZEK|20|13|et inritaverunt me domus Israhel in deserto in praeceptis meis non ambulaverunt et iudicia mea proiecerunt quae faciens homo vivet in eis et sabbata mea violaverunt vehementer dixi ergo ut effunderem furorem meum super eos in deserto et consumerem eos
EZEK|20|14|et feci propter nomen meum ne violaretur coram gentibus de quibus eieci eos in conspectu earum
EZEK|20|15|ego igitur levavi manum meam super eos in deserto ne inducerem eos in terram quam dedi eis fluentem lacte et melle praecipuam terrarum omnium
EZEK|20|16|quia iudicia mea proiecerunt et in praeceptis meis non ambulaverunt et sabbata mea violaverunt post idola enim cor eorum gradiebatur
EZEK|20|17|et pepercit oculus meus super eos ut non interficerem eos nec consumpsi eos in deserto
EZEK|20|18|dixi autem ad filios eorum in solitudine in praeceptis patrum vestrorum nolite incedere nec iudicia eorum custodiatis nec in idolis eorum polluamini
EZEK|20|19|ego Dominus Deus vester in praeceptis meis ambulate et iudicia mea custodite et facite ea
EZEK|20|20|et sabbata mea sanctificate ut sit signum inter me et vos et sciatur quia ego Dominus Deus vester
EZEK|20|21|et exacerbaverunt me filii in praeceptis meis non ambulaverunt et iudicia mea non custodierunt ut facerent ea quae cum fecerit homo vivet in eis et sabbata mea violaverunt et comminatus sum ut effunderem furorem meum super eos et implerem iram meam in eis in deserto
EZEK|20|22|averti autem manum meam et feci propter nomen meum ut non violaretur coram gentibus de quibus eieci eos in oculis earum
EZEK|20|23|iterum levavi manum meam in eos in solitudine ut dispergerem illos in nationes et ventilarem in terras
EZEK|20|24|eo quod iudicia mea non fecissent et praecepta mea reprobassent et sabbata mea violassent et post idola patrum suorum fuissent oculi eorum
EZEK|20|25|ergo et ego dedi eis praecepta non bona et iudicia in quibus non vivent
EZEK|20|26|et pollui eos in muneribus suis cum offerrent omne quod aperit vulvam propter delicta sua et scient quia ego Dominus
EZEK|20|27|quam ob rem loquere ad domum Israhel fili hominis et dices ad eos haec dicit Dominus Deus adhuc et in hoc blasphemaverunt me patres vestri cum sprevissent me contemnentes
EZEK|20|28|et induxissem eos in terram super quam levavi manum meam ut darem eis viderunt omnem collem excelsum et omne lignum nemorosum et immolaverunt ibi victimas suas et dederunt ibi inritationem oblationis suae et posuerunt ibi odorem suavitatis suae et libaverunt libationes suas
EZEK|20|29|et dixi ad eos quid est excelsum ad quod vos ingredimini et vocatum est nomen eius Excelsum usque ad hanc diem
EZEK|20|30|propterea dic ad domum Israhel haec dicit Dominus Deus certe in via patrum vestrorum vos polluimini et post offendicula eorum vos fornicamini
EZEK|20|31|et in oblatione donorum vestrorum cum transducitis filios vestros per ignem vos polluimini in omnibus idolis vestris usque hodie et ego respondebo vobis domus Israhel vivo ego dicit Dominus Deus quia non respondebo vobis
EZEK|20|32|neque cogitatio mentis vestrae fiet dicentium erimus sicut gentes et sicut cognationes terrae ut colamus ligna et lapides
EZEK|20|33|vivo ego dicit Dominus Deus quoniam in manu forti et brachio extento et in furore effuso regnabo super vos
EZEK|20|34|et educam vos de populis et congregabo vos de terris in quibus dispersi estis in manu valida et brachio extento et in furore effuso regnabo super vos
EZEK|20|35|et adducam vos in desertum populorum et iudicabor vobiscum ibi facie ad faciem
EZEK|20|36|sicut iudicio contendi adversum patres vestros in deserto terrae Aegypti sic iudicabo vos dicit Dominus Deus
EZEK|20|37|et subiciam vos sceptro meo et inducam vos in vinculis foederis
EZEK|20|38|et eligam de vobis transgressores et impios et de terra incolatus eorum educam eos et terram Israhel non ingredientur et scietis quia ego Dominus
EZEK|20|39|et vos domus Israhel haec dicit Dominus Deus singuli post idola vestra ambulate et servite eis quod si et in hoc non audieritis me et nomen meum sanctum pollueritis ultra in muneribus vestris et in idolis vestris
EZEK|20|40|in monte sancto meo in monte excelso Israhel ait Dominus Deus ibi serviet mihi omnis domus Israhel omnes inquam in terra in qua placebunt mihi et ibi quaeram primitias vestras et initium decimarum vestrarum in omnibus sanctificationibus vestris
EZEK|20|41|in odorem suavitatis suscipiam vos cum eduxero vos de populis et congregavero vos de terris in quas dispersi estis et sanctificabor in vobis in oculis nationum
EZEK|20|42|et scietis quia ego Dominus cum induxero vos ad terram Israhel in terram pro qua levavi manum meam ut darem eam patribus vestris
EZEK|20|43|et recordabimini ibi viarum vestrarum et omnium scelerum vestrorum quibus polluti estis in eis et displicebitis vobis in conspectu vestro in omnibus malitiis vestris quas fecistis
EZEK|20|44|et scietis quia ego Dominus cum benefecero vobis propter nomen meum non secundum vias vestras malas neque secundum scelera vestra pessima domus Israhel ait Dominus Deus
EZEK|20|45|et factus est sermo Domini ad me dicens
EZEK|20|46|fili hominis pone faciem tuam contra viam austri et stilla ad africum et propheta ad saltum agri meridiani
EZEK|20|47|et dices saltui meridiano audi verbum Domini haec dicit Dominus Deus ecce ego succendam in te ignem et conburam in te omne lignum viride et omne lignum aridum non extinguetur flamma succensionis et conburetur in ea omnis facies ab austro usque ad aquilonem
EZEK|20|48|et videbit universa caro quia ego Dominus succendi eam nec extinguetur
EZEK|20|49|et dixi ha ha ha Domine Deus ipsi dicunt de me numquid non per parabolas loquitur iste
EZEK|21|1|et factus est sermo Domini ad me dicens
EZEK|21|2|fili hominis pone faciem tuam ad Hierusalem et stilla ad sanctuaria et propheta contra humum Israhel
EZEK|21|3|et dices terrae Israhel haec dicit Dominus Deus ecce ego ad te et eiciam gladium meum de vagina sua et occidam in te iustum et impium
EZEK|21|4|pro eo autem quod occidi in te iustum et impium idcirco egredietur gladius meus de vagina sua ad omnem carnem ab austro ad aquilonem
EZEK|21|5|ut sciat omnis caro quia ego Dominus eduxi gladium meum de vagina sua inrevocabilem
EZEK|21|6|et tu fili hominis ingemesce in contritione lumborum et in amaritudinibus ingemesce coram eis
EZEK|21|7|cumque dixerint ad te quare tu gemis dices pro auditu quia venit et tabescet omne cor et dissolventur universae manus et infirmabitur omnis spiritus et per cuncta genua fluent aquae ecce venit et fiet ait Dominus Deus
EZEK|21|8|et factus est sermo Domini ad me dicens
EZEK|21|9|fili hominis propheta et dices haec dicit Dominus Deus loquere gladius gladius exacutus est et limatus
EZEK|21|10|ut caedat victimas exacutus est ut splendeat limatus est qui moves sceptrum filii mei succidisti omne lignum
EZEK|21|11|et dedi eum ad levigandum ut teneatur manu iste exacutus est gladius et iste limatus ut sit in manu interficientis
EZEK|21|12|clama et ulula fili hominis quia hic factus est in populo meo hic in cunctis ducibus Israhel qui fugerant gladio traditi sunt cum populo meo idcirco plaude super femur
EZEK|21|13|quia probatus est et hoc cum sceptrum subverterit et non erit dicit Dominus Deus
EZEK|21|14|tu ergo fili hominis propheta et percute manu ad manum et duplicetur gladius ac triplicetur gladius interfectorum hic est gladius occisionis magnae qui obstupescere eos facit
EZEK|21|15|et corde tabescere et multiplicat ruinas in omnibus portis eorum dedi conturbationem gladii acuti et limati ad fulgendum amicti ad caedem
EZEK|21|16|exacuere vade ad dextram sive ad sinistram quocumque faciei tuae est appetitus
EZEK|21|17|quin et ego plaudam manu ad manum et implebo indignationem meam ego Dominus locutus sum
EZEK|21|18|et factus est sermo Domini ad me dicens
EZEK|21|19|et tu fili hominis pone tibi duas vias ut veniat gladius regis Babylonis de terra una egredientur ambo et manu capiet coniecturam in capite viae civitatis coniciet
EZEK|21|20|viam pones ut veniat gladius ad Rabbath filiorum Ammon et ad Iudam in Hierusalem munitissimam
EZEK|21|21|stetit enim rex Babylonis in bivio in capite duarum viarum divinationem quaerens commiscens sagittas interrogavit idola exta consuluit
EZEK|21|22|ad dextram eius facta est divinatio super Hierusalem ut ponat arietes ut aperiat os in caede ut elevet vocem in ululatu ut ponat arietes contra portas ut conportet aggerem ut aedificet munitiones
EZEK|21|23|eritque quasi consulens frustra oraculum in oculis eorum et sabbatorum otium imitans ipse autem recordabitur iniquitatis ad capiendum
EZEK|21|24|idcirco haec dicit Dominus Deus pro eo quod recordati estis iniquitatis vestrae et revelastis praevaricationes vestras et apparuerunt peccata vestra in omnibus cogitationibus vestris pro eo inquam quod recordati estis manu capiemini
EZEK|21|25|tu autem profane impie dux Israhel cuius venit dies in tempore iniquitatis praefinita
EZEK|21|26|haec dicit Dominus Deus aufer cidarim tolle coronam nonne haec est quae humilem sublevavit et sublimem humiliavit
EZEK|21|27|iniquitatem iniquitatem iniquitatem ponam eam et hoc nunc factum est donec veniret cuius est iudicium et tradam ei
EZEK|21|28|et tu fili hominis propheta et dic haec dicit Dominus Deus ad filios Ammon et ad obprobrium eorum et dices mucro mucro evaginate ad occidendum limate ut interficias et fulgeas
EZEK|21|29|cum tibi viderentur vana et divinarentur mendacia ut dareris super colla vulneratorum impiorum quorum venit dies in tempore iniquitatis praefinita
EZEK|21|30|revertere ad vaginam tuam in loco in quo creatus es in terra nativitatis tuae iudicabo te
EZEK|21|31|et effundam super te indignationem meam in igne furoris mei sufflabo in te daboque te in manus hominum insipientium et fabricantium interitum
EZEK|21|32|igni eris cibus sanguis tuus erit in medio terrae oblivioni traderis quia ego Dominus locutus sum
EZEK|22|1|et factum est verbum Domini ad me dicens
EZEK|22|2|et tu fili hominis num iudicas num iudicas civitatem sanguinum
EZEK|22|3|et ostendes ei omnes abominationes suas et dices haec dicit Dominus Deus civitas effundens sanguinem in medio sui ut veniat tempus eius et quae fecit idola contra semet ipsam ut pollueretur
EZEK|22|4|in sanguine tuo qui a te effusus est deliquisti et in idolis tuis quae fecisti polluta es et adpropinquare fecisti dies tuos et adduxisti tempus annorum tuorum propterea dedi te obprobrium gentibus et inrisionem universis terris
EZEK|22|5|quae iuxta sunt et quae procul a te triumphabunt de te sordida nobilis grandis interitu
EZEK|22|6|ecce principes Israhel singuli in brachio suo fuerunt in te ad effundendum sanguinem
EZEK|22|7|patrem et matrem contumeliis adfecerunt in te advenam calumniati sunt in medio tui pupillum et viduam contristaverunt apud te
EZEK|22|8|sanctuaria mea sprevistis et sabbata mea polluistis
EZEK|22|9|viri detractores fuerunt in te ad effundendum sanguinem et super montes comederunt in te scelus operati sunt in medio tui
EZEK|22|10|verecundiora patris discoperuerunt in te inmunditiam menstruatae humiliaverunt in te
EZEK|22|11|et unusquisque in uxorem proximi sui operatus est abominationem et socer nurum suam polluit nefarie frater sororem suam filiam patris sui oppressit in te
EZEK|22|12|munera acceperunt apud te ad effundendum sanguinem usuram et superabundantiam accepisti et avare proximos tuos calumniabaris meique oblita es ait Dominus Deus
EZEK|22|13|ecce conplosi manus meas super avaritiam tuam quam fecisti et super sanguinem qui effusus est in medio tui
EZEK|22|14|numquid sustinebit cor tuum aut praevalebunt manus tuae in diebus quos ego faciam tibi ego Dominus locutus sum et faciam
EZEK|22|15|et dispergam te in nationes et ventilabo te in terras et deficere faciam inmunditiam tuam a te
EZEK|22|16|et possidebo te in conspectu gentium et scies quia ego Dominus
EZEK|22|17|et factum est verbum Domini ad me dicens
EZEK|22|18|fili hominis versa est mihi domus Israhel in scoriam omnes isti aes et stagnum et ferrum et plumbum in medio fornacis scoria argenti facti sunt
EZEK|22|19|propterea haec dicit Dominus Deus eo quod versi estis omnes in scoriam propterea ecce ego congregabo vos in medium Hierusalem
EZEK|22|20|congregatione argenti et aeris et ferri et stagni et plumbi in medium fornacis ut succendam in eam ignem ad conflandum sic congregabo in furore meo et in ira mea et requiescam et conflabo vos
EZEK|22|21|et congregabo vos et succendam vos in igne furoris mei et conflabimini in medio eius
EZEK|22|22|ut conflatur argentum in medio fornacis sic eritis in medio eius et scietis quia ego Dominus effuderim indignationem meam super vos
EZEK|22|23|et factum est verbum Domini ad me dicens
EZEK|22|24|fili hominis dic ei tu es terra inmunda et non conpluta in die furoris
EZEK|22|25|coniuratio prophetarum in medio eius sicut leo rugiens capiensque praedam animam devoraverunt opes et pretium acceperunt viduas eius multiplicaverunt in medio illius
EZEK|22|26|sacerdotes eius contempserunt legem meam et polluerunt sanctuaria mea inter sanctum et profanum non habuere distantiam et inter pollutum et mundum non intellexerunt et a sabbatis meis averterunt oculos suos et coinquinabar in medio eorum
EZEK|22|27|principes eius in medio illius quasi lupi rapientes praedam ad effundendum sanguinem et perdendas animas et avare sectanda lucra
EZEK|22|28|prophetae autem eius liniebant eos absque temperamento videntes vana et divinantes eis mendacium dicentes haec dicit Dominus Deus cum Dominus non sit locutus
EZEK|22|29|populi terrae calumniabantur calumniam et rapiebant violenter egenum et pauperem adfligebant et advenam opprimebant calumnia absque iudicio
EZEK|22|30|et quaesivi de eis virum qui interponeret sepem et staret oppositus contra me pro terra ne dissiparem eam et non inveni
EZEK|22|31|et effudi super eos indignationem meam in igne irae meae consumpsi eos viam eorum in caput eorum reddidi ait Dominus Deus
EZEK|23|1|et factus est sermo Domini ad me dicens
EZEK|23|2|fili hominis duae mulieres filiae matris unius fuerunt
EZEK|23|3|et fornicatae sunt in Aegypto in adulescentia sua fornicatae sunt ibi subacta sunt ubera earum et fractae sunt mammae pubertatis earum
EZEK|23|4|nomina autem earum Oolla maior et Ooliba soror eius et habui eas et pepererunt filios et filias porro earum nomina Samaria Oolla et Hierusalem Ooliba
EZEK|23|5|fornicata est igitur Oolla super me et insanivit in amatores suos in Assyrios propinquantes
EZEK|23|6|vestitos hyacintho principes et magistratus iuvenes cupidinis universos equites ascensores equorum
EZEK|23|7|et dedit fornicationes suas super eos electos filios Assyriorum universos et in omnibus in quos insanivit in inmunditiis eorum polluta est
EZEK|23|8|insuper et fornicationes suas quas habuerat in Aegypto non reliquit nam et illi dormierant cum ea in adulescentia eius et illi confregerant ubera pubertatis eius et effuderant fornicationem suam super eam
EZEK|23|9|propterea tradidi eam in manu amatorum suorum in manus filiorum Assur super quorum insanivit libidinem
EZEK|23|10|ipsi discoperuerunt ignominiam eius filios et filias illius tulerunt et ipsam occiderunt gladio et factae sunt famosae mulieres et iudicia perpetrarunt in ea
EZEK|23|11|quod cum vidisset soror eius Ooliba plus quam illa insanivit libidine et fornicationem suam super fornicationem sororis suae
EZEK|23|12|ad filios Assyriorum praebuit inpudenter ducibus et magistratibus ad se venientibus indutis veste varia equitibus qui vectabantur equis et adulescentibus forma cunctis egregia
EZEK|23|13|et vidi quod polluta esset via una ambarum
EZEK|23|14|et auxit fornicationes suas cumque vidisset viros depictos in pariete imagines Chaldeorum expressas coloribus
EZEK|23|15|et accinctos balteis renes et tiaras tinctas in capitibus eorum formam ducum omnium similitudinem filiorum Babylonis terraeque Chaldeorum in qua orti sunt
EZEK|23|16|et insanivit super eos concupiscentia oculorum suorum et misit nuntios ad eos in Chaldeam
EZEK|23|17|cumque venissent ad eam filii Babylonis ad cubile mammarum polluerunt eam stupris suis et polluta est ab eis et saturata est anima eius ab illis
EZEK|23|18|denudavit quoque fornicationes suas et discoperuit ignominiam suam et recessit anima mea ab ea sicut recesserat anima mea a sorore eius
EZEK|23|19|multiplicavit enim fornicationes suas recordans dies adulescentiae suae quibus fornicata est in terra Aegypti
EZEK|23|20|et insanivit libidine super concubitu eorum quorum carnes sunt ut carnes asinorum et sicut fluxus equorum fluxus eorum
EZEK|23|21|et visitasti scelus adulescentiae tuae quando subacta sunt in Aegypto ubera tua et confractae mammae pubertatis tuae
EZEK|23|22|propterea Ooliba haec dicit Dominus Deus ecce ego suscitabo omnes amatores tuos contra te de quibus satiata est anima tua et congregabo eos adversum te in circuitu
EZEK|23|23|filios Babylonis et universos Chaldeos nobiles tyrannosque et principes omnes filios Assyriorum iuvenes forma egregia duces et magistratus universos principes principum et nominatos ascensores equorum
EZEK|23|24|et venient super te instructi curru et rota multitudo populorum lorica et clypeo et galea armabuntur contra te undique et dabo coram eis iudicium et iudicabunt te iudiciis suis
EZEK|23|25|et ponam zelum meum in te quem exercent tecum in furore nasum tuum et aures tuas praecident et quae remanserint gladio concident ipsi filios tuos et filias tuas capient et novissimum tuum devorabitur igni
EZEK|23|26|et denudabunt te vestimentis tuis et tollent vasa gloriae tuae
EZEK|23|27|et requiescere faciam scelus tuum de te et fornicationem tuam de terra Aegypti nec levabis oculos tuos ad eos et Aegypti non recordaberis amplius
EZEK|23|28|quia haec dicit Dominus Deus ecce ego tradam te in manu eorum quos odisti in manu de quibus satiata est anima tua
EZEK|23|29|et agent tecum in odio et tollent omnes labores tuos et dimittent te nudam et ignominia plenam revelabitur ignominia fornicationum tuarum scelus tuum et fornicationes tuae
EZEK|23|30|fecerunt haec tibi quia fornicata es post gentes inter quas polluta es in idolis eorum
EZEK|23|31|in via sororis tuae ambulasti et dabo calicem eius in manu tua
EZEK|23|32|haec dicit Dominus Deus calicem sororis tuae bibes profundum et latum eris in derisum et in subsannationem quae es capacissima
EZEK|23|33|ebrietate et dolore repleberis calice maeroris et tristitiae calice sororis tuae Samariae
EZEK|23|34|et bibes illum et epotabis usque ad feces et fragmenta eius devorabis et ubera tua lacerabis quia ego locutus sum ait Dominus Deus
EZEK|23|35|propterea haec dicit Dominus Deus quia oblita es mei et proiecisti me post corpus tuum tu quoque porta scelus tuum et fornicationes tuas
EZEK|23|36|et ait Dominus ad me dicens fili hominis numquid iudicas Oollam et Oolibam et adnuntias eis scelera earum
EZEK|23|37|quia adulterae sunt et sanguis in manibus earum et cum idolis suis fornicatae sunt insuper et filios suos quos genuerunt mihi obtulerunt eis ad devorandum
EZEK|23|38|sed et hoc fecerunt mihi polluerunt sanctuarium meum in die illa et sabbata mea profanaverunt
EZEK|23|39|cumque immolarent filios suos idolis suis et ingrederentur sanctuarium meum in die illa ut polluerent illud etiam haec fecerunt in medio domus meae
EZEK|23|40|miserunt ad viros venientes de longe ad quos nuntium miserant itaque ecce venerunt quibus te lavisti et circumlevisti stibio oculos tuos et ornata es mundo muliebri
EZEK|23|41|sedisti in lecto pulcherrimo et mensa ordinata est ante te thymiama meum et unguentum meum posuisti super eam
EZEK|23|42|et vox multitudinis exultantis erat in ea et in viris qui de multitudine hominum adducebantur et veniebant de deserto posuerunt armillas in manibus eorum et coronas speciosas in capitibus eorum
EZEK|23|43|et dixi ei quae adtrita est in adulteriis nunc fornicabitur in fornicatione sua etiam haec
EZEK|23|44|et ingressi sunt ad eam quasi ad mulierem meretricem sic ingrediebantur ad Oollam et ad Oolibam mulieres nefarias
EZEK|23|45|viri ergo iusti sunt hii iudicabunt eas iudicio adulterarum et iudicio effundentium sanguinem quia adulterae sunt et sanguis in manibus earum
EZEK|23|46|haec enim dicit Dominus Deus adduc ad eas multitudinem et trade eas in tumultum et in rapinam
EZEK|23|47|et lapidentur lapidibus populorum et confodiantur gladiis eorum filios et filias earum interficient et domos earum igne succendent
EZEK|23|48|et auferam scelus de terra et discent omnes mulieres ne faciant secundum scelus earum
EZEK|23|49|et dabunt scelus vestrum super vos et peccata idolorum vestrorum portabitis et scietis quia ego Dominus Deus
EZEK|24|1|et factum est verbum Domini ad me in anno nono in mense decimo decima mensis dicens
EZEK|24|2|fili hominis scribe tibi nomen diei huius in qua confirmatus est rex Babylonis adversum Hierusalem hodie
EZEK|24|3|et dices per proverbium ad domum inritatricem parabolam et loqueris ad eos haec dicit Dominus Deus pone ollam pone inquam et mitte in ea aquam
EZEK|24|4|congere frusta eius in ea omnem partem bonam femur et armum electa et ossibus plena
EZEK|24|5|pinguissimum pecus adsume conpone quoque struices ossuum sub ea efferbuit coctio eius et discocta sunt ossa illius in medio eius
EZEK|24|6|propterea haec dicit Dominus Deus vae civitati sanguinum ollae cuius rubigo in ea est et rubigo eius non exivit de ea per partes et per partes suas eice eam non cecidit super eam sors
EZEK|24|7|sanguis enim eius in medio eius est super limpidissimam petram effudit illum non effudit illum super terram ut possit operiri pulvere
EZEK|24|8|ut superducerem indignationem meam et vindicta ulciscerer dedi sanguinem eius super petram limpidissimam ne operiretur
EZEK|24|9|propterea haec dicit Dominus Deus vae civitati sanguinum cuius ego grandem faciam pyram
EZEK|24|10|congere ossa quae igne succendam consumentur carnes et concoquetur universa conpositio et ossa tabescent
EZEK|24|11|pone quoque eam super prunas vacuam ut incalescat et liquefiat aes eius et confletur in medio eius inquinamentum eius et consumatur rubigo eius
EZEK|24|12|multo labore sudatum est et non exibit de ea nimia rubigo eius neque per ignem
EZEK|24|13|inmunditia tua execrabilis quia mundare te volui et non es mundata a sordibus tuis sed nec mundaberis prius donec quiescere faciam indignationem meam in te
EZEK|24|14|ego Dominus locutus sum venit et faciam non transeam nec parcam nec placabor iuxta vias tuas et iuxta adinventiones tuas iudicavi te dicit Dominus
EZEK|24|15|et factum est verbum Domini ad me dicens
EZEK|24|16|fili hominis ecce ego tollo a te desiderabile oculorum tuorum in plaga et non planges neque plorabis neque fluent lacrimae tuae
EZEK|24|17|ingemesce tacens mortuorum luctum non facies corona tua circumligata sit tibi et calciamenta tua erunt in pedibus tuis nec amictu ora velabis nec cibos lugentium comedes
EZEK|24|18|locutus sum ergo ad populum mane et mortua est uxor mea vesperi fecique mane sicut praeceperat mihi
EZEK|24|19|et dixit ad me populus quare non indicas nobis quid ista significent quae tu facis
EZEK|24|20|et dixi ad eos sermo Domini factus est ad me dicens
EZEK|24|21|loquere domui Israhel haec dicit Dominus Deus ecce ego polluam sanctuarium meum superbiam imperii vestri et desiderabile oculorum vestrorum et super quo pavet anima vestra et filii vestri et filiae quas reliquistis gladio cadent
EZEK|24|22|et facietis sicut feci ora amictu non velabitis et cibos lugentium non comedetis
EZEK|24|23|coronas habebitis in capitibus vestris et calciamenta in pedibus non plangetis neque flebitis sed tabescetis in iniquitatibus vestris et unusquisque gemet ad fratrem suum
EZEK|24|24|eritque Hiezecihel vobis in portentum iuxta omnia quae fecit facietis cum venerit istud et scietis quia ego Dominus Deus
EZEK|24|25|et tu fili hominis ecce in die quo tollam ab eis fortitudinem eorum et gaudium dignitatis et desiderium oculorum eorum super quo requiescunt animae eorum filios et filias eorum
EZEK|24|26|in die illa cum venerit fugiens ad te ut adnuntiet tibi
EZEK|24|27|in die inquam illa aperietur os tuum cum eo qui fugit et loqueris et non silebis ultra erisque eis in portentum et scietis quia ego Dominus
EZEK|25|1|et factus est sermo Domini ad me dicens
EZEK|25|2|fili hominis pone faciem tuam contra filios Ammon et prophetabis de eis
EZEK|25|3|et dices filiis Ammon audite verbum Domini Dei haec dicit Dominus Deus pro eo quod dixisti euge euge super sanctuarium meum quia pollutum est et super terram Israhel quoniam desolata est et super domum Iuda quoniam ducti sunt in captivitatem
EZEK|25|4|idcirco ego tradam te filiis orientalibus in hereditatem et conlocabunt caulas suas in te et ponent in te tentoria sua ipsi comedent fruges tuas et ipsi bibent lac tuum
EZEK|25|5|daboque Rabbath in habitaculum camelorum et filios Ammon in cubile pecorum et scietis quia ego Dominus
EZEK|25|6|quia haec dicit Dominus Deus pro eo quod plausisti manu et percussisti pede et gavisa es ex toto affectu super terram Israhel
EZEK|25|7|idcirco ecce ego extendam manum meam super te et tradam te in direptionem gentium et interficiam te de populis et perdam de terris et conteram et scies quia ego Dominus
EZEK|25|8|haec dicit Dominus Deus pro eo quod dixerunt Moab et Seir ecce sicut omnes gentes domus Iuda
EZEK|25|9|idcirco ecce ego aperiam umerum Moab de civitatibus de civitatibus inquam eius et de finibus eius inclitas terrae Bethiesimoth et Beelmeon et Cariathaim
EZEK|25|10|filiis orientis cum filiis Ammon et dabo eam in hereditatem ut non sit memoria ultra filiorum Ammon in gentibus
EZEK|25|11|et in Moab faciam iudicia et scient quia ego Dominus
EZEK|25|12|haec dicit Dominus Deus pro eo quod fecit Idumea ultionem ut se vindicaret de filiis Iuda peccavitque delinquens et vindictam expetivit de eis
EZEK|25|13|idcirco haec dicit Dominus Deus extendam manum meam super Idumeam et auferam de ea hominem et iumentum et faciam eam desertum ab austro et qui sunt in Daedan gladio cadent
EZEK|25|14|et dabo ultionem meam super Idumeam per manum populi mei Israhel et facient in Edom iuxta iram meam et furorem meum et scient vindictam meam dicit Dominus Deus
EZEK|25|15|haec dicit Dominus Deus pro eo quod fecerunt Palestini in vindictam et ulti se sunt toto animo interficientes et implentes inimicitias veteres
EZEK|25|16|propterea haec dicit Dominus Deus ecce ego extendam manum meam super Palestinos et interficiam interfectores et perdam reliquias maritimae regionis
EZEK|25|17|faciamque in eis ultiones magnas arguens in furore et scient quia ego Dominus cum dedero vindictam meam super eos
EZEK|26|1|et factum est in undecimo anno prima mensis factus est sermo Domini ad me dicens
EZEK|26|2|fili hominis pro eo quod dixit Tyrus de Hierusalem euge confractae sunt portae populorum conversa est ad me implebor deserta est
EZEK|26|3|propterea haec dicit Dominus Deus ecce ego super te Tyre et ascendere faciam ad te gentes multas sicut ascendit mare fluctuans
EZEK|26|4|et dissipabunt muros Tyri et destruent turres eius et radam pulverem eius de ea et dabo eam in limpidissimam petram
EZEK|26|5|siccatio sagenarum erit in medio maris quia ego locutus sum ait Dominus Deus et erit in direptionem gentibus
EZEK|26|6|filiae quoque eius quae sunt in agro gladio interficientur et scient quia ego Dominus
EZEK|26|7|quia haec dicit Dominus Deus ecce ego adducam ad Tyrum Nabuchodonosor regem Babylonis ab aquilone regem regum cum equis et curribus et equitibus et coetu populoque magno
EZEK|26|8|filias tuas quae sunt in agro gladio interficiet et circumdabit te munitionibus et conportabit aggerem in gyro et levabit contra te clypeum
EZEK|26|9|et vineas et arietes temperabit in muros tuos et turres tuas destruet in armatura sua
EZEK|26|10|inundatione equorum eius operiet te pulvis eorum a sonitu equitum et rotarum et curruum movebuntur muri tui dum ingressus fuerit portas tuas quasi per introitus urbis dissipatae
EZEK|26|11|ungulis equorum suorum conculcabit omnes plateas tuas populum tuum gladio caedet et statuae tuae nobiles in terram corruent
EZEK|26|12|vastabunt opes tuas diripient negotiationes tuas et destruent muros tuos et domos tuas praeclaras subvertent et lapides tuos et ligna tua et pulverem tuum in medio aquarum ponent
EZEK|26|13|et quiescere faciam multitudinem canticorum tuorum et sonitus cithararum tuarum non audietur amplius
EZEK|26|14|et dabo te in limpidissimam petram siccatio sagenarum eris nec aedificaberis ultra quia ego locutus sum dicit Dominus Deus
EZEK|26|15|haec dicit Dominus Deus Tyro numquid non a sonitu ruinae tuae et gemitu interfectorum tuorum cum occisi fuerint in medio tui commovebuntur insulae
EZEK|26|16|et descendent de sedibus suis omnes principes maris et auferent exuvias suas et vestimenta sua varia abicient et induentur stupore in terra sedebunt et adtoniti super repentino casu tuo admirabuntur
EZEK|26|17|et adsumentes super te lamentum dicent tibi quomodo peristi quae habitas in mari urbs inclita quae fuisti fortis in mari cum habitatoribus tuis quos formidabant universi
EZEK|26|18|nunc stupebunt naves in die pavoris tui et turbabuntur insulae in mari eo quod nullus egrediatur ex te
EZEK|26|19|quia haec dicit Dominus Deus cum dedero te urbem desolatam sicut civitates quae non habitantur et adduxero super te abyssum et operuerint te aquae multae
EZEK|26|20|et detraxero te cum his qui descendunt in lacum ad populum sempiternum et conlocavero te in terra novissima sicut solitudines veteres cum his qui deducuntur in lacum ut non habiteris porro dedero gloriam in terra viventium
EZEK|26|21|in nihilum redigam te et non eris et requisita non invenieris ultra in sempiternum dicit Dominus Deus
EZEK|27|1|et factum est verbum Domini ad me dicens
EZEK|27|2|tu ergo fili hominis adsume super Tyrum lamentum
EZEK|27|3|et dices Tyro quae habitat in introitu maris negotiationi populorum ad insulas multas haec dicit Dominus Deus o Tyre tu dixisti perfecti decoris ego sum
EZEK|27|4|et in corde maris sita finitimi tui qui te aedificaverunt impleverunt decorem tuum
EZEK|27|5|abietibus de Sanir extruxerunt te cum omnibus tabulatis maris cedrum de Libano tulerunt ut facerent tibi malum
EZEK|27|6|quercus de Basan dolaverunt in remos tuos transtra tua fecerunt tibi ex ebore indico et praetoriola de insulis Italiae
EZEK|27|7|byssus varia de Aegypto texta est tibi in velum ut poneretur in malo hyacinthus et purpura de insulis Elisa facta sunt operimentum tuum
EZEK|27|8|habitatores Sidonis et Aradii fuerunt remiges tui sapientes tui Tyre facti sunt gubernatores tui
EZEK|27|9|senes Bibli et prudentes eius habuerunt nautas ad ministerium variae supellectilis tuae omnes naves maris et nautae earum fuerunt in populo negotiationis tuae
EZEK|27|10|Persae et Lydi et Lybies erant in exercitu tuo viri bellatores tui clypeum et galeam suspenderunt in te pro ornatu tuo
EZEK|27|11|filii Aradii cum exercitu tuo erant super muros tuos in circuitu sed et Pigmei qui erant in turribus tuis faretras suas suspenderunt in muris tuis per gyrum ipsi conpleverunt pulchritudinem tuam
EZEK|27|12|Carthaginienses negotiatores tui a multitudine cunctarum divitiarum argento ferro stagno plumboque repleverunt nundinas tuas
EZEK|27|13|Graecia Thubal et Mosoch ipsi institores tui mancipia et vasa aerea adduxerunt populo tuo
EZEK|27|14|de domo Thogorma equos et equites et mulos adduxerunt ad forum tuum
EZEK|27|15|filii Dadan negotiatores tui insulae multae negotiatio manus tuae dentes eburneos et hebeninos commutaverunt in pretio tuo
EZEK|27|16|Syrus negotiator tuus propter multitudinem operum tuorum gemmam purpuram et scutulata et byssum et sericum et chodchod proposuerunt in mercatu tuo
EZEK|27|17|Iuda et terra Israhel ipsi institores tui in frumento primo balsamum et mel et oleum et resinam proposuerunt in nundinis tuis
EZEK|27|18|Damascenus negotiator tuus in multitudine operum tuorum in multitudine diversarum opum in vino pingui in lanis coloris optimi
EZEK|27|19|Dan et Graecia et Mozel in nundinis tuis proposuerunt ferrum fabrefactum stacte et calamus in negotiatione tua
EZEK|27|20|Dadan institores tui in tapetibus ad sedendum
EZEK|27|21|Arabia et universi principes Cedar ipsi negotiatores manus tuae cum agnis et arietibus et hedis venerunt ad te negotiatores tui
EZEK|27|22|venditores Saba et Reema ipsi negotiatores tui cum universis primis aromatibus et lapide pretioso et auro quod proposuerunt in mercatu tuo
EZEK|27|23|Aran et Chenne et Eden negotiatores Saba Assur Chelmad venditores tui
EZEK|27|24|ipsi negotiatores tui multifariam involucris hyacinthi et polymitorum gazarumque pretiosarum quae obvolutae et adstrictae erant funibus cedros quoque habebant in negotiationibus tuis
EZEK|27|25|naves maris principes tuae in negotiatione tua et repleta es et glorificata nimis in corde maris
EZEK|27|26|in aquis multis adduxerunt te remiges tui ventus auster contrivit te in corde maris
EZEK|27|27|divitiae tuae et thesauri tui et multiplex instrumentum tuum nautae tui et gubernatores tui qui tenebant supellectilem tuam et populo tuo praeerant viri quoque bellatores tui qui erant in te cum universa multitudine tua quae est in medio tui cadent in corde maris in die ruinae tuae
EZEK|27|28|a sonitu clamoris gubernatorum tuorum conturbabuntur classes
EZEK|27|29|et descendent de navibus suis omnes qui tenebant remum nautae et universi gubernatores maris in terra stabunt
EZEK|27|30|et heiulabunt super te voce magna et clamabunt amare et superiacient pulverem capitibus suis et cinere conspergentur
EZEK|27|31|et radent super te calvitium et accingentur ciliciis et plorabunt te in amaritudine animae ploratu amarissimo
EZEK|27|32|et adsument super te carmen lugubre et plangent te quae est ut Tyrus quae obmutuit in medio maris
EZEK|27|33|quae in exitu negotiationum tuarum de mari implesti populos multos in multitudine divitiarum tuarum et populorum tuorum ditasti reges terrae
EZEK|27|34|nunc contrita es a mari in profundis aquarum opes tuae et omnis multitudo tua quae erat in medio tui ceciderunt
EZEK|27|35|universi habitatores insularum obstipuerunt super te et reges earum omnes tempestate perculsi mutaverunt vultus
EZEK|27|36|negotiatores populorum sibilaverunt super te ad nihilum deducta es et non eris usque in perpetuum
EZEK|28|1|et factus est sermo Domini ad me dicens
EZEK|28|2|fili hominis dic principi Tyri haec dicit Dominus Deus eo quod elevatum est cor tuum et dixisti Deus ego sum et in cathedra Dei sedi in corde maris cum sis homo et non Deus et dedisti cor tuum quasi cor Dei
EZEK|28|3|ecce sapientior es tu Danihele omne secretum non est absconditum a te
EZEK|28|4|in sapientia et prudentia tua fecisti tibi fortitudinem et adquisisti aurum et argentum in thesauris tuis
EZEK|28|5|in multitudine sapientiae tuae et in negotiatione tua multiplicasti tibi fortitudinem et elevatum est cor tuum in robore tuo
EZEK|28|6|propterea haec dicit Dominus Deus eo quod elevatum est cor tuum quasi cor Dei
EZEK|28|7|idcirco ecce ego adducam super te alienos robustissimos gentium et nudabunt gladios suos super pulchritudinem sapientiae tuae et polluent decorem tuum
EZEK|28|8|interficient et detrahent te et morieris interitu occisorum in corde maris
EZEK|28|9|numquid dicens loqueris Deus ego sum coram interficientibus te cum sis homo et non Deus in manu occidentium te
EZEK|28|10|morte incircumcisorum morieris in manu alienorum quia ego locutus sum ait Dominus Deus
EZEK|28|11|et factus est sermo Domini ad me dicens fili hominis leva planctum super regem Tyri
EZEK|28|12|et dices ei haec dicit Dominus Deus tu signaculum similitudinis plenus sapientia et perfectus decore
EZEK|28|13|in deliciis paradisi Dei fuisti omnis lapis pretiosus operimentum tuum sardius topazius et iaspis chrysolitus et onyx et berillus sapphyrus et carbunculus et zmaragdus aurum opus decoris tui et foramina tua in die qua conditus es praeparata sunt
EZEK|28|14|tu cherub extentus et protegens et posui te in monte sancto Dei in medio lapidum ignitorum ambulasti
EZEK|28|15|perfectus in viis tuis a die conditionis tuae donec inventa est iniquitas in te
EZEK|28|16|in multitudine negotiationis tuae repleta sunt interiora tua iniquitate et peccasti et eieci te de monte Dei et perdidi te o cherub protegens de medio lapidum ignitorum
EZEK|28|17|elevatum est cor tuum in decore tuo perdidisti sapientiam tuam in decore tuo in terram proieci te ante faciem regum dedi te ut cernerent te
EZEK|28|18|in multitudine iniquitatum tuarum et iniquitate negotiationis tuae polluisti sanctificationem tuam producam ergo ignem de medio tui qui comedat te et dabo te in cinerem super terram in conspectu omnium videntium te
EZEK|28|19|omnes qui viderint te in gentibus obstupescent super te nihili factus es et non eris in perpetuum
EZEK|28|20|et factus est sermo Domini ad me dicens
EZEK|28|21|fili hominis pone faciem tuam contra Sidonem et prophetabis de ea
EZEK|28|22|et dices haec dicit Dominus Deus ecce ego ad te Sidon et glorificabor in medio tui et scient quia ego Dominus cum fecero in ea iudicia et sanctificatus fuero in ea
EZEK|28|23|et inmittam ei pestilentiam et sanguinem in plateis eius et corruent interfecti in medio eius gladio per circuitum et scient quia ego Dominus
EZEK|28|24|et non erit ultra domui Israhel offendiculum amaritudinis et spina dolorem inferens undique per circuitum eorum qui adversantur eis et scient quia ego Dominus Deus
EZEK|28|25|haec dicit Dominus Deus quando congregavero domum Israhel de populis in quibus dispersi sunt sanctificabor in eis coram gentibus et habitabunt in terra sua quam dedi servo meo Iacob
EZEK|28|26|et habitabunt in ea securi et aedificabunt domos plantabuntque vineas et habitabunt confidenter cum fecero iudicia in omnibus qui adversantur eis per circuitum et scient quia ego Dominus Deus eorum
EZEK|29|1|in anno decimo in decimo mense undecima mensis factum est verbum Domini ad me dicens
EZEK|29|2|fili hominis pone faciem tuam contra Pharaonem regem Aegypti et prophetabis de eo et de Aegypto universa
EZEK|29|3|loquere et dices haec dicit Dominus Deus ecce ego ad te Pharao rex Aegypti draco magne qui cubas in medio fluminum tuorum et dicis meus est fluvius et ego feci memet ipsum
EZEK|29|4|et ponam frenum in maxillis tuis et adglutinabo pisces fluminum tuorum squamis tuis et extraham te de medio fluminum tuorum et universi pisces tui squamis tuis adherebunt
EZEK|29|5|et proiciam te in desertum et omnes pisces fluminis tui super faciem terrae cades non colligeris neque congregaberis bestiis terrae et volatilibus caeli dedi te ad devorandum
EZEK|29|6|et scient omnes habitatores Aegypti quia ego Dominus pro eo quod fuisti baculus harundineus domui Israhel
EZEK|29|7|quando adprehenderunt te manu et confractus es et lacerasti omnem umerum eorum et innitentibus eis super te comminutus es et dissolvisti omnes renes eorum
EZEK|29|8|propterea haec dicit Dominus Deus ecce ego adducam super te gladium et interficiam de te hominem et iumentum
EZEK|29|9|et erit terra Aegypti in desertum et solitudinem et scient quia ego Dominus eo quod dixerit fluvius meus est et ego feci
EZEK|29|10|idcirco ecce ego ad te et ad flumina tua daboque terram Aegypti in solitudines gladio dissipatam a turre Syenes usque ad terminos Aethiopiae
EZEK|29|11|non pertransibit eam pes hominis neque pes iumenti gradietur in ea et non habitabitur quadraginta annis
EZEK|29|12|daboque terram Aegypti desertam in medio terrarum desertarum et civitates eius in medio urbium subversarum erunt desolatae quadraginta annis et dispergam Aegyptios in nationes et ventilabo eos in terras
EZEK|29|13|quia haec dicit Dominus Deus post finem quadraginta annorum congregabo Aegyptum de populis in quibus dispersi fuerunt
EZEK|29|14|et reducam captivitatem Aegypti et conlocabo eos in terra Fatures in terra nativitatis suae et erunt ibi in regnum humile
EZEK|29|15|inter regna cetera erit humillima et non elevabitur ultra super nationes et inminuam eos ne imperent gentibus
EZEK|29|16|neque erunt ultra domui Israhel in confidentia docentes iniquitatem ut fugiant et sequantur eos et scient quia ego Dominus Deus
EZEK|29|17|et factum est in vicesimo et septimo anno in primo in una mensis factum est verbum Domini ad me dicens
EZEK|29|18|fili hominis Nabuchodonosor rex Babylonis servire fecit exercitum suum servitute magna adversum Tyrum omne caput decalvatum et omnis umerus depilatus est et merces non est reddita ei neque exercitui eius de Tyro pro servitute qua servivit mihi adversum eam
EZEK|29|19|propterea haec dicit Dominus Deus ecce ego dabo Nabuchodonosor regem Babylonis in terra Aegypti et accipiet multitudinem eius et depraedabitur manubias eius et diripiet spolia eius et erit merces exercitui illius
EZEK|29|20|et operi pro quo servivit adversum eam dedi ei terram Aegypti pro eo quod laboraverunt mihi ait Dominus Deus
EZEK|29|21|in die illo pullulabit cornu domui Israhel et tibi dabo apertum os in medio eorum et scient quoniam ego Dominus
EZEK|30|1|et factum est verbum Domini ad me dicens
EZEK|30|2|fili hominis propheta et dic haec dicit Dominus Deus ululate vae vae diei
EZEK|30|3|quia iuxta est dies et adpropinquavit dies Domini dies nubis tempus gentium erit
EZEK|30|4|et veniet gladius in Aegyptum et erit pavor in Aethiopia cum ceciderint vulnerati in Aegypto et ablata fuerit multitudo illius et destructa fundamenta eius
EZEK|30|5|Aethiopia et Lybia et Lydii et omne reliquum vulgus et Chub et filii terrae foederis cum eis gladio cadent
EZEK|30|6|haec dicit Dominus Deus et corruent fulcientes Aegyptum et destruetur superbia imperii eius a turre Syenes gladio cadent in ea ait Dominus exercituum
EZEK|30|7|et dissipabuntur in medio terrarum desolatarum et urbes eius in medio civitatum desertarum erunt
EZEK|30|8|et scient quoniam ego Dominus cum dedero ignem in Aegyptum et adtriti fuerint omnes auxiliatores eius
EZEK|30|9|in die illa egredientur nuntii a facie mea in trieribus ad conterendam Aethiopiae confidentiam et erit pavor in eis in die Aegypti quia absque dubio veniet
EZEK|30|10|haec dicit Dominus Deus et cessare faciam multitudinem Aegypti in manu Nabuchodonosor regis Babylonis
EZEK|30|11|ipse et populus eius cum eo fortissimi gentium adducentur ad disperdendam terram et evaginabunt gladios suos super Aegyptum et implebunt terram interfectis
EZEK|30|12|et faciam alveos fluminum aridos et tradam terram in manu pessimorum et dissipabo terram et plenitudinem eius in manu alienorum ego Dominus locutus sum
EZEK|30|13|haec dicit Dominus Deus et disperdam simulacra et cessare faciam idola de Memphis et dux de terra Aegypti non erit amplius et dabo terrorem in terra Aegypti
EZEK|30|14|et disperdam terram Fatures et dabo ignem in Tafnis et faciam iudicia in Alexandriam
EZEK|30|15|et effundam indignationem meam super Pelusium robur Aegypti et interficiam multitudinem Alexandriae
EZEK|30|16|et dabo ignem in Aegypto quasi parturiens dolebit Pelusium et Alexandria erit dissipata et in Memphis angustiae cotidianae
EZEK|30|17|iuvenes Eliupoleos et Bubasti gladio cadent et ipsae captivae ducentur
EZEK|30|18|et in Tafnis nigrescet dies cum contrivero ibi sceptra Aegypti et defecerit in ea superbia potentiae eius ipsam nubes operiet filiae autem eius in captivitatem ducentur
EZEK|30|19|et faciam iudicia in Aegypto et scient quia ego Dominus
EZEK|30|20|et factum est in undecimo anno in primo in septima mensis factum est verbum Domini ad me dicens
EZEK|30|21|fili hominis brachium Pharao regis Aegypti confregi et ecce non est obvolutum ut restitueretur ei sanitas ut ligaretur pannis et farciretur linteolis et recepto robore posset tenere gladium
EZEK|30|22|propterea haec dicit Dominus Deus ecce ego ad Pharao regem Aegypti et comminuam brachium eius forte sed confractum et deiciam gladium de manu eius
EZEK|30|23|et dispergam Aegyptum in gentibus et ventilabo eos in terris
EZEK|30|24|et confortabo brachia regis Babylonis daboque gladium meum in manu eius et confringam brachia Pharaonis et gement gemitibus interfecti coram facie eius
EZEK|30|25|et confortabo brachia regis Babylonis et brachia Pharaonis concident et scient quia ego Dominus cum dedero gladium meum in manu regis Babylonis et extenderit eum super terram Aegypti
EZEK|30|26|et dispergam Aegyptum in nationes et ventilabo eos in terris et scient quia ego Dominus
EZEK|31|1|et factum est in undecimo anno tertio una mensis factum est verbum Domini ad me dicens
EZEK|31|2|fili hominis dic Pharaoni regi Aegypti et populo eius cui similis factus es in magnitudine tua
EZEK|31|3|ecce Assur quasi cedrus in Libano pulcher ramis et frondibus nemorosus excelsusque altitudine et inter condensas frondes elevatum est cacumen eius
EZEK|31|4|aquae nutrierunt illum abyssus exaltavit eum flumina eius manabant in circuitu radicum eius et rivos suos emisit ad universa ligna regionis
EZEK|31|5|propterea elevata est altitudo eius super omnia ligna regionis et multiplicata sunt arbusta eius et elevati sunt rami eius prae aquis multis
EZEK|31|6|cumque extendisset umbram suam in ramis eius fecerunt nidos omnia volatilia caeli et sub frondibus eius genuerunt omnes bestiae saltuum et sub umbraculo illius habitabat coetus gentium plurimarum
EZEK|31|7|eratque pulcherrimus in magnitudine sua et in dilatatione arbustorum suorum erat enim radix illius iuxta aquas multas
EZEK|31|8|cedri non fuerunt altiores illo in paradiso Dei abietes non adaequaverunt summitatem eius et platani non fuerunt aequae frondibus illius omne lignum paradisi Dei non est adsimilatum illi et pulchritudini eius
EZEK|31|9|quoniam speciosum feci eum et multis condensisque frondibus et aemulata sunt eum omnia ligna voluptatis quae erant in paradiso Dei
EZEK|31|10|propterea haec dicit Dominus Deus pro eo quod sublimatus est in altitudine et dedit summitatem suam virentem atque condensam et elevatum est cor eius in altitudine sua
EZEK|31|11|tradidi eum in manu fortissimi gentium faciens faciet ei iuxta impietatem eius eieci eum
EZEK|31|12|et succident illum alieni et crudelissimi nationum et proicient eum super montes et in cunctis convallibus corruent rami eius et confringentur arbusta eius in universis rupibus terrae et recedent de umbraculo eius omnes populi terrae et relinquent eum
EZEK|31|13|in ruina eius habitaverunt omnia volatilia caeli et in ramis eius fuerunt universae bestiae regionis
EZEK|31|14|quam ob rem non elevabuntur in altitudine sua omnia ligna aquarum neque ponent sublimitatem suam inter nemorosa atque frondosa nec stabunt in sublimitate eorum omnia quae inrigantur aquis quia omnes traditi sunt in mortem ad terram ultimam in medio filiorum hominum ad eos qui descendunt in lacum
EZEK|31|15|haec dicit Dominus Deus in die quando descendit ad inferos indixi luctum operui eum abysso et prohibui flumina eius et coercui aquas multas contristatus est super eum Libanus et omnia ligna agri concussa sunt
EZEK|31|16|a sonitu ruinae eius commovi gentes cum deducerem eum ad infernum cum his qui descendebant in lacum et consolata sunt in terra infima omnia ligna voluptatis egregia atque praeclara in Libano universa quae inrigabantur aquis
EZEK|31|17|nam et ipsi cum ea descendent ad infernum ad interfectos gladio et brachium uniuscuiusque sedebit sub umbraculo eius in medio nationum
EZEK|31|18|cui adsimilatus es o inclite atque sublimis inter ligna voluptatis ecce deductus es cum lignis voluptatis ad terram ultimam in medio incircumcisorum dormies cum his qui interfecti sunt gladio ipse est Pharao et omnis multitudo eius dicit Dominus Deus
EZEK|32|1|et factum est duodecimo anno in mense duodecimo in una mensis factum est verbum Domini ad me dicens
EZEK|32|2|fili hominis adsume lamentum super Pharao regem Aegypti et dices ad eum leoni gentium adsimilatus es et draconi qui est in mari et ventilabas cornu in fluminibus tuis et conturbabas aquas pedibus tuis et conculcabas flumina eorum
EZEK|32|3|propterea haec dicit Dominus Deus expandam super te rete meum in multitudine populorum multorum et extrahent te in sagena mea
EZEK|32|4|et proiciam te in terram super faciem agri abiciam te et habitare faciam super te omnia volatilia caeli et saturabo de te bestias universae terrae
EZEK|32|5|et dabo carnes tuas super montes et implebo colles tuos sanie tua
EZEK|32|6|et inrigabo terram pedore sanguinis tui super montes et valles implebuntur ex te
EZEK|32|7|et operiam cum extinctus fueris caelos et nigrescere faciam stellas eius solem nube tegam et luna non dabit lumen suum
EZEK|32|8|omnia luminaria caeli maerere faciam super te et dabo tenebras super terram tuam dicit Dominus Deus
EZEK|32|9|et inritabo cor populorum multorum cum induxero contritionem tuam in gentibus super terras quas nescis
EZEK|32|10|et stupescere faciam super te populos multos et reges eorum horrore nimio formidabunt super te cum volare coeperit gladius meus super facies eorum et obstupescent repente singuli pro anima sua in die ruinae suae
EZEK|32|11|quia haec dicit Dominus Deus gladius regis Babylonis veniet tibi
EZEK|32|12|in gladiis fortium deiciam multitudinem tuam inexpugnabiles gentes omnes heae et vastabunt superbiam Aegypti et dissipabitur multitudo eius
EZEK|32|13|et perdam omnia iumenta eius quae erant super aquas plurimas et non conturbabit eas pes hominis ultra neque ungula iumentorum turbabit eas
EZEK|32|14|tunc purissimas reddam aquas eorum et flumina eorum quasi oleum adducam ait Dominus Deus
EZEK|32|15|cum dedero terram Aegypti desolatam deseretur autem terra a plenitudine sua quando percussero omnes habitatores eius et scient quia ego Dominus
EZEK|32|16|planctus est et plangent eum filiae gentium plangent eum super Aegypto et super multitudine eius plangent eum ait Dominus Deus
EZEK|32|17|et factum est in duodecimo anno in quintadecima mensis factum est verbum Domini ad me dicens
EZEK|32|18|fili hominis cane lugubre super multitudine Aegypti et detrahe eam ipsam et filias gentium robustarum ad terram ultimam cum his qui descendunt in lacum
EZEK|32|19|quo pulchrior es descende et dormi cum incircumcisis
EZEK|32|20|in medio interfectorum gladio cadent gladius datus est adtraxerunt eam et omnes populos eius
EZEK|32|21|loquentur ei potentissimi robustorum de medio inferni qui cum auxiliatoribus eius descenderunt et dormierunt incircumcisi interfecti gladio
EZEK|32|22|ibi Assur et omnis multitudo eius in circuitu illius sepulchra eius omnes interfecti et qui ceciderunt gladio
EZEK|32|23|quorum data sunt sepulchra in novissimis laci et facta est multitudo eius per gyrum sepulchri eius universi interfecti cadentesque gladio qui dederant quondam formidinem in terra viventium
EZEK|32|24|ibi Aelam et omnis multitudo eius per gyrum sepulchri sui omnes hii interfecti ruentesque gladio qui descenderunt incircumcisi ad terram ultimam qui posuerunt terrorem suum in terra viventium et portaverunt ignominiam suam cum his qui descendunt in lacum
EZEK|32|25|in medio interfectorum posuerunt cubile eius in universis populis eius in circuitu eius sepulchrum illius omnes hii incircumcisi interfectique gladio dederant enim terrorem in terra viventium et portaverunt ignominiam suam cum his qui descendunt in lacum in medio interfectorum positi sunt
EZEK|32|26|ibi Mosoch et Thubal et omnis multitudo eius in circuitu illius sepulchra eius omnes hii incircumcisi interfectique et cadentes gladio quia dederunt formidinem suam in terra viventium
EZEK|32|27|et non dormient cum fortibus cadentibusque et incircumcisis qui descenderunt ad infernum cum armis suis et posuerunt gladios suos sub capitibus suis et fuerunt iniquitates eorum in ossibus eorum quia terror fortium facti sunt in terra viventium
EZEK|32|28|et tu ergo in medio incircumcisorum contereris et dormies cum interfectis gladio
EZEK|32|29|ibi Idumea et reges eius omnes duces eius qui dati sunt cum exercitu suo cum interfectis gladio et qui cum incircumcisis dormierunt et cum his qui descenderunt in lacum
EZEK|32|30|ibi principes aquilonis omnes et universi venatores qui deducti sunt cum interfectis paventes et in sua fortitudine confusi qui dormierunt incircumcisi cum interfectis gladio et portaverunt confusionem suam cum his qui descendunt in lacum
EZEK|32|31|vidit eos Pharao et consolatus est super universa multitudine sua quae interfecta est gladio Pharao et omnis exercitus eius ait Dominus Deus
EZEK|32|32|quia dedi terrorem meum in terra viventium et dormivit in medio incircumcisorum cum interfectis gladio Pharao et omnis multitudo eius ait Dominus Deus
EZEK|33|1|et factum est verbum Domini ad me dicens
EZEK|33|2|fili hominis loquere ad filios populi tui et dices ad eos terra cum induxero super eam gladium et tulerit populus terrae virum unum de novissimis suis et constituerit eum super se speculatorem
EZEK|33|3|et ille viderit gladium venientem super terram et cecinerit bucina et adnuntiaverit populo
EZEK|33|4|audiens autem quisquis ille est sonum bucinae non se observaverit veneritque gladius et tulerit eum sanguis ipsius super caput eius erit
EZEK|33|5|sonum bucinae audivit et non se observavit sanguis eius in ipso erit si autem custodierit animam suam salvavit
EZEK|33|6|quod si speculator viderit gladium venientem et non insonuerit bucina et populus non se custodierit veneritque gladius et tulerit de eis animam ille quidem in iniquitate sua captus est sanguinem autem eius de manu speculatoris requiram
EZEK|33|7|et tu fili hominis speculatorem dedi te domui Israhel audiens ergo ex ore meo sermonem adnuntiabis eis ex me
EZEK|33|8|si me dicente ad impium impie morte morieris non fueris locutus ut se custodiat impius a via sua ipse impius in iniquitate sua morietur sanguinem autem eius de manu tua requiram
EZEK|33|9|si autem adnuntiante te ad impium ut a viis suis convertatur non fuerit conversus a via sua ipse in iniquitate sua morietur porro tu animam tuam liberasti
EZEK|33|10|tu ergo fili hominis dic ad domum Israhel sic locuti estis dicentes iniquitates nostrae et peccata nostra super nos sunt et in ipsis nos tabescimus quomodo ergo vivere poterimus
EZEK|33|11|dic ad eos vivo ego dicit Dominus Deus nolo mortem impii sed ut revertatur impius a via sua et vivat convertimini a viis vestris pessimis et quare moriemini domus Israhel
EZEK|33|12|tu itaque fili hominis dic ad filios populi tui iustitia iusti non liberabit eum in quacumque die peccaverit et impietas impii non nocebit ei in quacumque die conversus fuerit ab impietate sua et iustus non poterit vivere in iustitia sua in quacumque die peccaverit
EZEK|33|13|etiam si dixero iusto quod vita vivat et confisus in iustitia sua fecerit iniquitatem omnes iustitiae eius oblivioni tradentur et in iniquitate sua quam operatus est in ipsa morietur
EZEK|33|14|sin autem dixero impio morte morieris et egerit paenitentiam a peccato suo feceritque iudicium et iustitiam
EZEK|33|15|pignus restituerit ille impius rapinamque reddiderit in mandatis vitae ambulaverit nec fecerit quicquam iniustum vita vivet et non morietur
EZEK|33|16|omnia peccata eius quae peccavit non inputabuntur ei iudicium et iustitiam fecit vita vivet
EZEK|33|17|et dixerunt filii populi tui non est aequi ponderis via Domini et ipsorum via iniusta est
EZEK|33|18|cum enim recesserit iustus a iustitia sua feceritque iniquitatem morietur in eis
EZEK|33|19|et cum recesserit impius ab impietate sua feceritque iudicium et iustitiam vivet in eis
EZEK|33|20|et dicitis non est recta via Domini unumquemque iuxta vias suas iudicabo de vobis domus Israhel
EZEK|33|21|et factum est in duodecimo anno in duodecimo mense in quinta mensis transmigrationis nostrae venit ad me qui fugerat de Hierusalem dicens vastata est civitas
EZEK|33|22|manus autem Domini facta fuerat ad me vespere antequam veniret qui fugerat aperuitque os meum donec veniret ad me mane et aperto ore meo non silui amplius
EZEK|33|23|et factum est verbum Domini ad me dicens
EZEK|33|24|fili hominis qui habitant in ruinosis his super humum Israhel loquentes aiunt unus erat Abraham et hereditate possedit terram nos autem multi nobis data est terra in possessionem
EZEK|33|25|idcirco dices ad eos haec dicit Dominus Deus qui in sanguine comeditis et oculos vestros levatis ad inmunditias vestras et sanguinem funditis numquid terram hereditate possidebitis
EZEK|33|26|stetistis in gladiis vestris fecistis abominationes et unusquisque uxorem proximi sui polluit et terram hereditate possidebitis
EZEK|33|27|haec dices ad eos sic dicit Dominus Deus vivo ego quia qui in ruinosis habitant gladio cadent et qui in agro est bestiis tradetur ad devorandum qui autem in praesidiis et in speluncis sunt peste morientur
EZEK|33|28|et dabo terram in solitudinem et desertum et deficiet superba fortitudo eius et desolabuntur montes Israhel eo quod nullus sit qui per eos transeat
EZEK|33|29|et scient quia ego Dominus cum dedero terram desolatam et desertam propter universas abominationes suas quas operati sunt
EZEK|33|30|et tu fili hominis filii populi tui qui loquuntur de te iuxta muros et in ostiis domorum et dicunt unus ad alterum vir ad proximum suum loquentes venite et audiamus qui sit sermo egrediens a Domino
EZEK|33|31|et veniunt ad te quasi si ingrediatur populus et sedent coram te populus meus et audiunt sermones tuos et non faciunt eos quia in canticum oris sui vertunt illos et avaritiam suam sequitur cor eorum
EZEK|33|32|et es eis quasi carmen musicum quod suavi dulcique sono canitur et audient verba tua et non facient ea
EZEK|33|33|et cum venerit quod praedictum est ecce enim venit tunc scient quod prophetes fuerit inter eos
EZEK|34|1|et factum est verbum Domini ad me dicens
EZEK|34|2|fili hominis propheta de pastoribus Israhel propheta et dices pastoribus haec dicit Dominus Deus vae pastoribus Israhel qui pascebant semet ipsos nonne greges pascuntur a pastoribus
EZEK|34|3|lac comedebatis et lanis operiebamini et quod crassum erat occidebatis gregem autem meum non pascebatis
EZEK|34|4|quod infirmum fuit non consolidastis et quod aegrotum non sanastis quod fractum est non alligastis et quod abiectum est non reduxistis quod perierat non quaesistis sed cum austeritate imperabatis eis et cum potentia
EZEK|34|5|et dispersae sunt oves meae eo quod non esset pastor et factae sunt in devorationem omnium bestiarum agri et dispersae sunt
EZEK|34|6|erraverunt greges mei in cunctis montibus et in universo colle excelso et super omnem faciem terrae dispersi sunt greges mei et non erat qui requireret non erat inquam qui requireret
EZEK|34|7|propterea pastores audite verbum Domini
EZEK|34|8|vivo ego dicit Dominus Deus quia pro eo quod facti sunt greges mei in rapinam et oves meae in devorationem omnium bestiarum agri eo quod non esset pastor neque enim quaesierunt pastores gregem meum sed pascebant pastores semet ipsos et greges meos non pascebant
EZEK|34|9|propterea pastores audite verbum Domini
EZEK|34|10|haec dicit Dominus Deus ecce ego ipse super pastores requiram gregem meum de manu eorum et cessare eos faciam ut ultra non pascant gregem nec pascant amplius pastores semet ipsos et liberabo gregem meum de ore eorum et non erunt ultra eis in escam
EZEK|34|11|quia haec dicit Dominus Deus ecce ego ipse requiram oves meas et visitabo eas
EZEK|34|12|sicut visitat pastor gregem suum in die quando fuerit in medio ovium suarum dissipatarum sic visitabo oves meas et liberabo eas de omnibus locis quo dispersae fuerant in die nubis et caliginis
EZEK|34|13|et educam eas de populis et congregabo eas de terris et inducam eas in terram suam et pascam eas in montibus Israhel in rivis et in cunctis sedibus terrae
EZEK|34|14|in pascuis uberrimis pascam eas et in montibus excelsis Israhel erunt pascuae eorum ibi requiescent in herbis virentibus et in pascuis pinguibus pascentur super montes Israhel
EZEK|34|15|ego pascam oves meas et ego eas accubare faciam dicit Dominus Deus
EZEK|34|16|quod perierat requiram et quod abiectum erat reducam et quod confractum fuerat alligabo et quod infirmum erat consolidabo et quod pingue et forte custodiam et pascam illas in iudicio
EZEK|34|17|vos autem greges mei haec dicit Dominus Deus ecce ego iudico inter pecus et pecus arietum et hircorum
EZEK|34|18|nonne satis vobis erat pascuam bonam depasci insuper et reliquias pascuarum vestrarum conculcastis pedibus vestris et cum purissimam aquam biberetis reliquam pedibus vestris turbabatis
EZEK|34|19|et oves meae his quae conculcata pedibus vestris fuerant pascebantur et quae pedes vestri turbaverant haec bibebant
EZEK|34|20|propterea haec dicit Dominus Deus ad eos ecce ego ipse iudico inter pecus pingue et macilentum
EZEK|34|21|pro eo quod lateribus et umeris inpingebatis et cornibus vestris ventilabatis omnia infirma pecora donec dispergerentur foras
EZEK|34|22|salvabo gregem meum et non erit ultra in rapinam et iudicabo inter pecus et pecus
EZEK|34|23|et suscitabo super ea pastorem unum qui pascat ea servum meum David ipse pascet ea et ipse erit eis in pastorem
EZEK|34|24|ego autem Dominus ero eis in Deum et servus meus David princeps in medio eorum ego Dominus locutus sum
EZEK|34|25|et faciam cum eis pactum pacis et cessare faciam bestias pessimas de terra et qui habitant in deserto securi dormient in saltibus
EZEK|34|26|et ponam eos in circuitu collis mei benedictionem et deducam imbrem in tempore suo pluviae benedictionis erunt
EZEK|34|27|et dabit lignum agri fructum suum et terra dabit germen suum et erunt in terra sua absque timore et scient quia ego Dominus cum contrivero catenas iugi eorum et eruero eos de manu imperantium sibi
EZEK|34|28|et non erunt ultra in rapinam gentibus neque bestiae terrae devorabunt eos sed habitabunt confidenter absque ullo terrore
EZEK|34|29|et suscitabo eis germen nominatum et non erunt ultra inminuti fame in terra neque portabunt amplius obprobria gentium
EZEK|34|30|et scient quia ego Dominus Deus eorum cum eis et ipsi populus meus domus Israhel ait Dominus Deus
EZEK|34|31|vos autem greges mei greges pascuae meae homines estis et ego Dominus Deus vester dicit Dominus Deus
EZEK|35|1|et factus est sermo Domini ad me dicens
EZEK|35|2|fili hominis pone faciem tuam adversum montem Seir et prophetabis de eo et dices illi
EZEK|35|3|haec dicit Dominus Deus ecce ego ad te mons Seir et extendam manum meam super te et dabo te desolatum atque desertum
EZEK|35|4|urbes tuas demoliar et tu desertus eris et scies quia ego Dominus
EZEK|35|5|eo quod fueris inimicus sempiternus et concluseris filios Israhel in manus gladii in tempore adflictionis eorum in tempore iniquitatis extremae
EZEK|35|6|propterea vivo ego dicit Dominus Deus quoniam sanguini tradam te et sanguis te persequetur et cum sanguinem oderis sanguis persequetur te
EZEK|35|7|et dabo montem Seir desolatum et desertum et auferam de eo euntem et redeuntem
EZEK|35|8|et implebo montes eius occisorum suorum in collibus tuis et in vallibus tuis atque in torrentibus interfecti gladio cadent
EZEK|35|9|in solitudines sempiternas tradam te et civitates tuae non habitabuntur et scietis quoniam ego Dominus
EZEK|35|10|eo quod dixeris duae gentes et duae terrae meae erunt et hereditate possidebo eas cum Dominus esset ibi
EZEK|35|11|propterea vivo ego dicit Dominus Deus quia faciam iuxta iram tuam et secundum zelum tuum quem fecisti odio habens eos et notus efficiar per eos cum te iudicavero
EZEK|35|12|et scies quia ego Dominus audivi universa obprobria tua quae locutus es de montibus Israhel dicens deserti nobis dati sunt ad devorandum
EZEK|35|13|et insurrexistis super me ore vestro et rogastis adversum me verba vestra ego audivi
EZEK|35|14|haec dicit Dominus Deus laetante universa terra in solitudinem te redigam
EZEK|35|15|sicuti gavisus es super hereditatem domus Israhel eo quod fuerit dissipata sic faciam tibi dissipatus eris mons Seir et Idumea omnis et scient quia ego Dominus
EZEK|36|1|tu autem fili hominis propheta super montes Israhel et dices montes Israhel audite verbum Domini
EZEK|36|2|haec dicit Dominus Deus eo quod dixerit inimicus de vobis euge altitudines sempiternae in hereditatem datae sunt nobis
EZEK|36|3|propterea vaticinare et dic haec dicit Dominus Deus pro eo quod desolati estis et conculcati per circuitum et facti in hereditatem reliquis gentibus et ascendistis super labium linguae et obprobrium populi
EZEK|36|4|propterea montes Israhel audite verbum Domini Dei haec dicit Dominus Deus montibus et collibus torrentibus vallibusque et desertis parietinis et urbibus derelictis quae depopulatae sunt et subsannatae a reliquis gentibus per circuitum
EZEK|36|5|propterea haec dicit Dominus Deus quoniam in igne zeli mei locutus sum de reliquis gentibus et de Idumea universa qui dederunt terram meam sibi in hereditatem cum gaudio et toto corde ex animo et eiecerunt eam ut vastarent
EZEK|36|6|idcirco vaticinare super humum Israhel et dices montibus et collibus iugis et vallibus haec dicit Dominus Deus ecce ego in zelo meo et in furore meo locutus sum eo quod confusionem gentium sustinueritis
EZEK|36|7|idcirco haec dicit Dominus Deus ego levavi manum meam ut gentes quae in circuitu vestro sunt ipsae confusionem suam portent
EZEK|36|8|vos autem montes Israhel ramos vestros germinetis et fructum vestrum adferatis populo meo Israhel prope est enim ut veniat
EZEK|36|9|quia ecce ego ad vos et convertar ad vos et arabimini et accipietis sementem
EZEK|36|10|et multiplicabo in vobis homines omnemque domum Israhel et habitabuntur civitates et ruinosa instaurabuntur
EZEK|36|11|et replebo vos hominibus et iumentis et multiplicabuntur et crescent et habitari vos faciam sicut a principio bonisque donabo maioribus quam habuistis ab initio et scietis quia ego Dominus
EZEK|36|12|et adducam super vos homines populum meum Israhel et hereditate possidebunt te et eris eis in hereditatem et non addes ultra ut absque eis sis
EZEK|36|13|haec dicit Dominus Deus pro eo quod dicunt de vobis devoratrix hominum es et suffocans gentem tuam
EZEK|36|14|propterea homines non comedes amplius et gentem tuam non necabis ultra ait Dominus Deus
EZEK|36|15|nec auditam faciam in te amplius confusionem gentium et obprobrium populorum nequaquam portabis et gentem tuam non amittes amplius ait Dominus Deus
EZEK|36|16|et factum est verbum Domini ad me dicens
EZEK|36|17|fili hominis domus Israhel habitaverunt in humo sua et polluerunt eam in viis suis et in studiis suis iuxta inmunditiam menstruatae facta est via eorum coram me
EZEK|36|18|et effudi indignationem meam super eos pro sanguine quem fuderunt super terram et in idolis suis polluerunt eam
EZEK|36|19|et dispersi eos in gentes et ventilati sunt in terris iuxta vias eorum et adinventiones iudicavi eos
EZEK|36|20|et ingressi sunt ad gentes ad quas introierunt et polluerunt nomen sanctum meum cum diceretur de eis populus Domini iste est et de terra eius egressi sunt
EZEK|36|21|et peperci nomini meo sancto quod polluerat domus Israhel in gentibus ad quas ingressi sunt
EZEK|36|22|idcirco dices domui Israhel haec dicit Dominus Deus non propter vos ego faciam domus Israhel sed propter nomen sanctum meum quod polluistis in gentibus ad quas intrastis
EZEK|36|23|et sanctificabo nomen meum magnum quod pollutum est inter gentes quod polluistis in medio earum ut sciant gentes quia ego Dominus ait Dominus exercituum cum sanctificatus fuero in vobis coram eis
EZEK|36|24|tollam quippe vos de gentibus et congregabo de universis terris et adducam vos in terram vestram
EZEK|36|25|et effundam super vos aquam mundam et mundabimini ab omnibus inquinamentis vestris et ab universis idolis vestris mundabo vos
EZEK|36|26|et dabo vobis cor novum et spiritum novum ponam in medio vestri et auferam cor lapideum de carne vestra et dabo vobis cor carneum
EZEK|36|27|et spiritum meum ponam in medio vestri et faciam ut in praeceptis meis ambuletis et iudicia mea custodiatis et operemini
EZEK|36|28|et habitabitis in terra quam dedi patribus vestris et eritis mihi in populum et ego ero vobis in Deum
EZEK|36|29|et salvabo vos ex universis inquinamentis vestris et vocabo frumentum et multiplicabo illud et non inponam in vobis famem
EZEK|36|30|et multiplicabo fructum ligni et genimina agri ut non portetis ultra obprobrium famis in gentibus
EZEK|36|31|et recordabimini viarum vestrarum pessimarum studiorumque non bonorum et displicebunt vobis iniquitates vestrae et scelera vestra
EZEK|36|32|non propter vos ego faciam ait Dominus Deus notum sit vobis confundimini et erubescite super viis vestris domus Israhel
EZEK|36|33|haec dicit Dominus Deus in die qua mundavero vos ex omnibus iniquitatibus vestris et habitari fecero urbes et instauravero ruinosa
EZEK|36|34|et terra deserta fuerit exculta quae quondam erat desolata in oculis omnis viatoris
EZEK|36|35|dicent terra illa inculta facta est ut hortus voluptatis et civitates desertae et destitutae atque suffossae munitae sederunt
EZEK|36|36|et scient gentes quaecumque derelictae fuerint in circuitu vestro quia ego Dominus aedificavi dissipata plantavique inculta ego Dominus locutus sum et fecerim
EZEK|36|37|haec dicit Dominus Deus adhuc in hoc invenient me domus Israhel ut faciam eis multiplicabo eos sicut gregem hominum
EZEK|36|38|ut gregem sanctum ut gregem Hierusalem in sollemnitatibus eius sic erunt civitates desertae plenaeque gregibus hominum et scient quia ego Dominus
EZEK|37|1|facta est super me manus Domini et eduxit me in spiritu Domini et dimisit me in medio campi qui erat plenus ossibus
EZEK|37|2|et circumduxit me per ea in gyro erant autem multa valde super faciem campi siccaque vehementer
EZEK|37|3|et dixit ad me fili hominis putasne vivent ossa ista et dixi Domine Deus tu nosti
EZEK|37|4|et dixit ad me vaticinare de ossibus istis et dices eis ossa arida audite verbum Domini
EZEK|37|5|haec dicit Dominus Deus ossibus his ecce ego intromittam in vos spiritum et vivetis
EZEK|37|6|et dabo super vos nervos et succrescere faciam super vos carnes et superextendam in vobis cutem et dabo vobis spiritum et vivetis et scietis quia ego Dominus
EZEK|37|7|et prophetavi sicut praeceperat mihi factus est autem sonitus prophetante me et ecce commotio et accesserunt ossa ad ossa unumquodque ad iuncturam suam
EZEK|37|8|et vidi et ecce super ea nervi et carnes ascenderunt et extenta est in eis cutis desuper et spiritum non habebant
EZEK|37|9|et dixit ad me vaticinare ad spiritum vaticinare fili hominis et dices ad spiritum haec dicit Dominus Deus a quattuor ventis veni spiritus et insufla super interfectos istos et revivescant
EZEK|37|10|et prophetavi sicut praeceperat mihi et ingressus est in ea spiritus et vixerunt steteruntque super pedes suos exercitus grandis nimis valde
EZEK|37|11|et dixit ad me fili hominis ossa haec universa domus Israhel est ipsi dicunt aruerunt ossa nostra et periit spes nostra et abscisi sumus
EZEK|37|12|propterea vaticinare et dices ad eos haec dicit Dominus Deus ecce ego aperiam tumulos vestros et educam vos de sepulchris vestris populus meus et inducam vos in terram Israhel
EZEK|37|13|et scietis quia ego Dominus cum aperuero sepulchra vestra et eduxero vos de tumulis vestris populus meus
EZEK|37|14|et dedero spiritum meum in vobis et vixeritis et requiescere vos faciam super humum vestram et scietis quia ego Dominus locutus sum et feci ait Dominus Deus
EZEK|37|15|et factus est sermo Domini ad me dicens
EZEK|37|16|et tu fili hominis sume tibi lignum unum et scribe super illud Iudae et filiorum Israhel sociis eius et tolle lignum alterum et scribe super eum Ioseph lignum Ephraim et cunctae domui Israhel sociorumque eius
EZEK|37|17|et adiunge illa unum ad alterum tibi in lignum unum et erunt in unionem in manu tua
EZEK|37|18|cum autem dixerint ad te filii populi tui loquentes nonne indicas nobis quid in his tibi velis
EZEK|37|19|loqueris ad eos haec dicit Dominus Deus ecce ego adsumam lignum Ioseph quod est in manu Ephraim et tribus Israhel quae iunctae sunt ei et dabo eas pariter cum ligno Iuda et faciam eas in lignum unum et erunt unum in manu eius
EZEK|37|20|erunt autem ligna super quae scripseris in manu tua in oculis eorum
EZEK|37|21|et dices ad eos haec dicit Dominus Deus ecce ego adsumam filios Israhel de medio nationum ad quas abierunt et congregabo eos undique et adducam eos ad humum suam
EZEK|37|22|et faciam eos gentem unam in terra in montibus Israhel et rex unus erit omnibus imperans et non erunt ultra duae gentes nec dividentur amplius in duo regna
EZEK|37|23|neque polluentur ultra in idolis suis et abominationibus suis et in cunctis iniquitatibus suis et salvos eos faciam de universis sedibus suis in quibus peccaverunt et mundabo eos et erunt mihi populus et ego ero eis Deus
EZEK|37|24|et servus meus David rex super eos et pastor unus erit omnium eorum in iudiciis meis ambulabunt et mandata mea custodient et facient ea
EZEK|37|25|et habitabunt super terram quam dedi servo meo Iacob in qua habitaverunt patres vestri et habitabunt super eam ipsi et filii eorum et filii filiorum eorum usque in sempiternum et David servus meus princeps eorum in perpetuum
EZEK|37|26|et percutiam illis foedus pacis pactum sempiternum erit eis et fundabo eos et multiplicabo et dabo sanctificationem meam in medio eorum in perpetuum
EZEK|37|27|et erit tabernaculum meum in eis et ero eis Deus et ipsi erunt mihi populus
EZEK|37|28|et scient gentes quia ego Dominus sanctificator Israhel cum fuerit sanctificatio mea in medio eorum in perpetuum
EZEK|38|1|et factus est sermo Domini ad me dicens
EZEK|38|2|fili hominis pone faciem tuam contra Gog terram Magog principem capitis Mosoch et Thubal et vaticinare de eo
EZEK|38|3|et dices ad eum haec dicit Dominus Deus ecce ego ad te Gog principem capitis Mosoch et Thubal
EZEK|38|4|et circumagam te et ponam frenum in maxillis tuis et educam te et omnem exercitum tuum equos et equites vestitos loricis universos multitudinem magnam hastam et clypeum arripientium et gladium
EZEK|38|5|Persae Aethiopes et Lybies cum eis omnes scutati et galeati
EZEK|38|6|Gomer et universa agmina eius domus Thogorma latera aquilonis et totum robur eius populique multi tecum
EZEK|38|7|praepara et instrue te et omnem multitudinem tuam quae coacervata est ad te et esto eis in praeceptum
EZEK|38|8|post dies multos visitaberis in novissimo annorum venies ad terram quae reversa est a gladio congregata est de populis multis ad montes Israhel qui fuerunt deserti iugiter haec de populis educta est et habitaverunt in ea confidenter universi
EZEK|38|9|ascendens autem quasi tempestas venies et quasi nubes ut operias terram tu et omnia agmina tua et populi multi tecum
EZEK|38|10|haec dicit Dominus Deus in die illa ascendent sermones super cor tuum et cogitabis cogitationem pessimam
EZEK|38|11|et dices ascendam ad terram absque muro veniam ad quiescentes habitantesque secure omnes habitant sine muro vectes et portae non sunt eis
EZEK|38|12|ut diripias spolia et invadas praedam ut inferas manum tuam super eos qui deserti fuerant et postea restituti et super populum qui est congregatus ex gentibus qui possidere coepit et esse habitator umbilici terrae
EZEK|38|13|Seba et Dedan et negotiatores Tharsis et omnes leones eius dicent tibi numquid ad sumenda spolia tu venis ecce ad diripiendam praedam congregasti multitudinem tuam ut tollas argentum et aurum auferas supellectilem atque substantiam et diripias manubias infinitas
EZEK|38|14|propterea vaticinare fili hominis et dices ad Gog haec dicit Dominus Deus numquid non in die illo cum habitaverit populus meus Israhel confidenter scies
EZEK|38|15|et venies de loco tuo a lateribus aquilonis tu et populi multi tecum ascensores equorum universi coetus magnus et exercitus vehemens
EZEK|38|16|et ascendes super populum meum Israhel quasi nubes ut operias terram in novissimis diebus eris et adducam te super terram meam ut sciant gentes me cum sanctificatus fuero in te in oculis eorum o Gog
EZEK|38|17|haec dicit Dominus Deus tu ergo ille es de quo locutus sum in diebus antiquis in manu servorum meorum prophetarum Israhel qui prophetaverunt in diebus illorum temporum ut adducerem te super eos
EZEK|38|18|et erit in die illa in die adventus Gog super terram Israhel ait Dominus Deus ascendet indignatio mea in furore meo
EZEK|38|19|et in zelo meo in igne irae meae locutus sum quia in die illa erit commotio magna super terram Israhel
EZEK|38|20|et commovebuntur a facie mea pisces maris et volucres caeli et bestiae agri et omne reptile quod movetur super humum cunctique homines qui sunt super faciem terrae et subvertentur montes et cadent sepes et omnis murus in terra corruet
EZEK|38|21|et convocabo adversum eum in cunctis montibus meis gladium ait Dominus Deus gladius uniuscuiusque in fratrem suum dirigetur
EZEK|38|22|et iudicabo eum peste et sanguine et imbre vehementi et lapidibus inmensis ignem et sulphur pluam super eum et super exercitum eius et super populos multos qui sunt cum eo
EZEK|38|23|et magnificabor et sanctificabor et notus ero in oculis gentium multarum et scient quia ego Dominus
EZEK|39|1|tu autem fili hominis vaticinare adversum Gog et dices haec dicit Dominus Deus ecce ego super te Gog principem capitis Mosoch et Thubal
EZEK|39|2|et circumagam te et seducam te et ascendere faciam de lateribus aquilonis et adducam te super montes Israhel
EZEK|39|3|et percutiam arcum tuum in manu sinistra tua et sagittas tuas de manu dextera tua deiciam
EZEK|39|4|super montes Israhel cades tu et omnia agmina tua et populi qui sunt tecum feris avibus omnique volatili et bestiis terrae dedi te devorandum
EZEK|39|5|super faciem agri cades quia ego locutus sum ait Dominus Deus
EZEK|39|6|et emittam ignem in Magog et in his qui habitant in insulis confidenter et scient quia ego Dominus
EZEK|39|7|et nomen sanctum meum notum faciam in medio populi mei Israhel et non polluam nomen sanctum meum amplius et scient gentes quia ego Dominus Sanctus Israhel
EZEK|39|8|ecce venit et factum est ait Dominus Deus haec est dies de qua locutus sum
EZEK|39|9|et egredientur habitatores de civitatibus Israhel et succendent et conburent arma clypeum et hastas arcum et sagittas et baculos manus et contos et succendent ea igne septem annis
EZEK|39|10|et non portabunt ligna de regionibus neque succident de saltibus quoniam arma succendent igne et depraedabuntur eos quibus praedae fuerant et diripient vastatores suos ait Dominus Deus
EZEK|39|11|et erit in die illa dabo Gog locum nominatum sepulchrum in Israhel vallem Viatorum ad orientem maris quae obstupescere facit praetereuntes et sepelient ibi Gog et omnem multitudinem eius et vocabitur vallis Multitudinis Gog
EZEK|39|12|et sepelient eos domus Israhel ut mundent terram septem mensibus
EZEK|39|13|sepeliet autem omnis populus terrae et erit eis nominata dies in qua glorificatus sum ait Dominus Deus
EZEK|39|14|et viros iugiter constituent lustrantes terram qui sepeliant et requirant eos qui remanserant super faciem terrae ut emundent eam post menses autem septem quaerere incipient
EZEK|39|15|et circumibunt peragrantes terram cumque viderint os hominis statuent iuxta illud titulum donec sepeliant illud pollinctores in valle Multitudinis Gog
EZEK|39|16|nomen autem civitatis Amona et mundabunt terram
EZEK|39|17|tu ergo fili hominis haec dicit Dominus Deus dic omni volucri et universis avibus cunctisque bestiis agri convenite properate concurrite undique ad victimam meam quam ego immolo vobis victimam grandem super montes Israhel ut comedatis carnes et bibatis sanguinem
EZEK|39|18|carnes fortium comedetis et sanguinem principum terrae bibetis arietum agnorum et hircorum taurorumque altilium et pinguium omnium
EZEK|39|19|et comedetis adipem in saturitate et bibetis sanguinem in ebrietate de victima quam ego immolabo vobis
EZEK|39|20|et saturabimini super mensam meam de equo et de equite forti et de universis viris bellatoribus ait Dominus Deus
EZEK|39|21|et ponam gloriam meam in gentibus et videbunt omnes gentes iudicium meum quod fecerim et manum meam quam posuerim super eos
EZEK|39|22|et scient domus Israhel quia ego Dominus Deus eorum a die illa et deinceps
EZEK|39|23|et scient gentes quoniam in iniquitate sua capta sit domus Israhel eo quod reliquerint me et absconderim faciem meam ab eis et tradiderim eos in manu hostium et ceciderint in gladio universi
EZEK|39|24|iuxta inmunditiam eorum et scelus feci eis et abscondi faciem meam ab illis
EZEK|39|25|propterea haec dicit Dominus Deus nunc reducam captivitatem Iacob et miserebor omnis domus Israhel et adsumam zelum pro nomine sancto meo
EZEK|39|26|et portabunt confusionem suam et omnem praevaricationem quam praevaricati sunt in me cum habitaverint in terra sua confidenter neminem formidantes
EZEK|39|27|et reduxero eos de populis et congregavero de terris inimicorum suorum et sanctificatus fuero in eis in oculis gentium plurimarum
EZEK|39|28|et scient quia ego Dominus Deus eorum eo quod transtulerim eos in nationes et congregavero eos super terram suam et non dereliquerim quemquam ex eis ibi
EZEK|39|29|et non abscondam ultra faciem meam ab eis eo quod effuderim spiritum meum super omnem domum Israhel ait Dominus Deus
EZEK|40|1|in vicesimo et quinto anno transmigrationis nostrae in exordio anni decima mensis quartodecimo anno postquam percussa est civitas in ipsa hac die facta est super me manus Domini et adduxit me illuc
EZEK|40|2|in visionibus Dei adduxit me in terram Israhel et dimisit me super montem excelsum nimis super quem erat quasi aedificium civitatis vergentis ad austrum
EZEK|40|3|et introduxit me illuc et ecce vir cuius erat species quasi species aeris et funiculus lineus in manu eius et calamus mensurae in manu eius stabat autem in porta
EZEK|40|4|et locutus est ad me idem vir fili hominis vide oculis tuis et auribus tuis audi et pone cor tuum in omnia quae ego ostendam tibi quia ut ostendantur tibi adductus es huc adnuntia omnia quae tu vides domui Israhel
EZEK|40|5|et ecce murus forinsecus in circuitu domus undique et in manu viri calamus mensurae sex cubitorum et palmo et mensus est latitudinem aedificii calamo uno altitudinem quoque calamo uno
EZEK|40|6|et venit ad portam quae respiciebat viam orientalem et ascendit per gradus eius et mensus est limen portae calamo uno latitudinem id est limen unum calamo uno in latitudine
EZEK|40|7|et thalamum uno calamo in longum et uno calamo in latum et inter thalamos quinque cubitos
EZEK|40|8|et limen portae iuxta vestibulum portae intrinsecus calamo uno
EZEK|40|9|et mensus est vestibulum portae octo cubitorum et frontem eius duobus cubitis vestibulum autem portae erat intrinsecus
EZEK|40|10|porro thalami portae ad viam orientalem tres hinc et tres inde mensura una trium et mensura una frontium ex utraque parte
EZEK|40|11|et mensus est latitudinem liminis portae decem cubitorum et longitudinem portae tredecim cubitorum
EZEK|40|12|et marginem ante thalamos cubiti unius et cubitus unus finis utrimque thalami autem sex cubitorum erant hinc et inde
EZEK|40|13|et mensus est portam a tecto thalami usque ad tectum eius latitudinem viginti et quinque cubitorum ostium contra ostium
EZEK|40|14|et fecit frontes per sexaginta cubitos et ad frontem atrium portae undique per circuitum
EZEK|40|15|et ante faciem portae quae pertingebat usque ad faciem vestibuli portae interioris quinquaginta cubitos
EZEK|40|16|et fenestras obliquas in thalamis et in frontibus eorum quae erant intra portam undique per circuitum similiter autem erant et in vestibulis fenestrae per gyrum intrinsecus et ante frontes pictura palmarum
EZEK|40|17|et eduxit me ad atrium exterius et ecce gazofilacia et pavimentum stratum lapide in atrio per circuitum triginta gazofilacia in circuitu pavimenti
EZEK|40|18|et pavimentum in fronte portarum secundum longitudinem portarum erat inferius
EZEK|40|19|et mensus est latitudinem a facie portae inferioris usque ad frontem atrii interioris extrinsecus centum cubitos ad orientem et ad aquilonem
EZEK|40|20|portam quoque quae respiciebat viam aquilonis atrii exterioris mensus est tam in longitudine quam in latitudine
EZEK|40|21|et thalamos eius tres hinc et tres inde et frontem eius et vestibulum eius secundum mensuram portae prioris quinquaginta cubitorum longitudinem eius et latitudinem viginti quinque cubitorum
EZEK|40|22|fenestrae autem eius et vestibulum et scalpturae secundum mensuram portae quae respiciebat ad orientem et septem graduum erat ascensus eius et vestibulum ante eam
EZEK|40|23|et porta atrii interioris contra portam aquilonis et orientalem et mensus est a porta usque ad portam centum cubitos
EZEK|40|24|et duxit me ad viam australem et ecce porta quae respiciebat ad austrum et mensus est frontem eius et vestibulum eius iuxta mensuras superiores
EZEK|40|25|et fenestras eius et vestibula in circuitu sicut fenestras ceteras quinquaginta cubitorum longitudine et latitudine viginti quinque cubitorum
EZEK|40|26|et in gradibus septem ascendebatur ad eam et vestibulum ante fores eius et celatae palmae erant una hinc et altera inde in fronte eius
EZEK|40|27|et porta atrii interioris in via australi et mensus est a porta usque ad portam in via australi centum cubitos
EZEK|40|28|et introduxit me in atrium interius ad portam australem et mensus est portam iuxta mensuras superiores
EZEK|40|29|thalamum eius et frontem eius et vestibulum eius hisdem mensuris et fenestras eius et vestibulorum eius in circuitu quinquaginta cubitos longitudinis et latitudinis viginti quinque cubitos
EZEK|40|30|et vestibulum per gyrum longitudine viginti quinque cubitorum et latitudine quinque cubitorum
EZEK|40|31|et vestibulum eius ad atrium exterius et palmas eius in fronte et octo gradus erant quibus ascendebatur per eam
EZEK|40|32|et introduxit me in atrium interius per viam orientalem et mensus est portam secundum mensuras superiores
EZEK|40|33|thalamum eius et frontem eius et vestibula eius sicut supra et fenestras eius et vestibuli eius in circuitu longitudine quinquaginta cubitorum et latitudine viginti quinque cubitorum
EZEK|40|34|et vestibulum eius id est atrii exterioris et palmae celatae in fronte eius hinc et inde et in octo gradibus ascensus eius
EZEK|40|35|et introduxit me ad portam quae respiciebat ad aquilonem et mensus est secundum mensuras superiores
EZEK|40|36|thalamum eius frontem eius vestibulum eius et fenestras eius per circuitum longitudine quinquaginta cubitorum et latitudine viginti quinque cubitorum
EZEK|40|37|vestibulum eius in atrium exterius et celatura palmarum in fronte illius hinc et inde et in octo gradibus ascensus eius
EZEK|40|38|et per singula gazofilacia ostium in frontibus portarum ibi lavabunt holocaustum
EZEK|40|39|et in vestibulo portae duae mensae hinc et duae mensae inde ut immoletur super eas holocaustum et pro peccato et pro delicto
EZEK|40|40|et ad latus exterius quod ascendit ad ostium portae quae pergit ad aquilonem duae mensae et ad latus alterum ante vestibulum portae duae mensae
EZEK|40|41|quattuor mensae hinc et quattuor mensae inde per latera portae octo mensae erunt super quas immolabunt
EZEK|40|42|quattuor autem mensae ad holocaustum de lapidibus quadris extructae longitudine cubiti unius et dimidii et latitudine cubiti unius et dimidii et altitudine cubiti unius super quas ponant vasa in quibus immolatur holocaustum et victima
EZEK|40|43|et labia earum palmi unius reflexa intrinsecus per circuitum super mensas autem carnes oblationis
EZEK|40|44|et extra portam interiorem gazofilacia cantorum in atrio interiori quod erat in latere portae respicientis ad aquilonem et facies eorum contra viam australem una ex latere portae orientalis quae respiciebat ad viam aquilonis
EZEK|40|45|et dixit ad me hoc est gazofilacium quod respicit viam meridianam sacerdotum qui excubant in custodiis templi
EZEK|40|46|porro gazofilacium quod respicit ad viam aquilonis sacerdotum erit qui excubant ad ministerium altaris isti sunt filii Sadoc qui accedunt de filiis Levi ad Dominum ut ministrent ei
EZEK|40|47|et mensus est atrium longitudine centum cubitorum et latitudine centum cubitorum per quadrum et altare ante faciem templi
EZEK|40|48|et introduxit me in vestibulum templi et mensus est vestibulum quinque cubitis hinc et quinque cubitis inde et latitudinem portae trium cubitorum hinc et trium cubitorum inde
EZEK|40|49|longitudinem autem vestibuli viginti cubitorum et latitudinem undecim cubitorum et octo gradibus ascendebatur ad eam et columnae erant in frontibus una hinc et altera inde
EZEK|41|1|et introduxit me in templum et mensus est frontes sex cubitos latitudinis hinc et sex cubitos latitudinis inde latitudinem tabernaculi
EZEK|41|2|et latitudo portae decem cubitorum erat et latera portae quinque cubitis hinc et quinque cubitis inde et mensus est longitudinem eius quadraginta cubitorum et latitudinem viginti cubitorum
EZEK|41|3|et introgressus intrinsecus mensus est in fronte portae duos cubitos et portam sex cubitorum et latitudinem portae septem cubitorum
EZEK|41|4|et mensus est longitudinem eius viginti cubitorum et latitudinem viginti cubitorum ante faciem templi et dixit ad me hoc est sanctum sanctorum
EZEK|41|5|et mensus est parietem domus sex cubitorum et latitudinem lateris quattuor cubitorum undique per circuitum domus
EZEK|41|6|latera autem latus ad latus bis triginta tria et erant eminentia quae ingrederentur per parietem domus in lateribus per circuitum ut continerent et non adtingerent parietem templi
EZEK|41|7|et platea erat in rotundum ascendens sursum per cocleam et in cenaculum templi deferebat per gyrum idcirco latius erat templum in superioribus et sic de inferioribus ascendebatur ad superiora in medium
EZEK|41|8|et vidi in domo altitudinem per circuitum fundata latera ad mensuram calami sex cubitorum spatio
EZEK|41|9|et latitudinem per parietem lateris forinsecus quinque cubitorum et interior domus in lateribus domus
EZEK|41|10|et inter gazofilacia latitudinem viginti cubitorum in circuitu domus undique
EZEK|41|11|et ostium lateris ad orationem ostium unum ad viam aquilonis et ostium unum ad viam australem et latitudinem loci ad orationem quinque cubitorum in circuitu
EZEK|41|12|et aedificium quod erat separatum versumque ad viam respicientem ad mare latitudinis septuaginta cubitorum paries autem aedificii quinque cubitorum latitudinis per circuitum et longitudo eius nonaginta cubitorum
EZEK|41|13|et mensus est domus longitudinem centum cubitorum et quod separatum erat aedificium et parietes eius longitudinis centum cubitorum
EZEK|41|14|latitudo autem ante faciem domus et eius quod erat separatum contra orientem centum cubitorum
EZEK|41|15|et mensus est longitudinem aedificii contra faciem eius quod erat separatum ad dorsum ekthetas ex utraque parte centum cubitorum et templum interius et vestibula atrii
EZEK|41|16|limina et fenestras obliquas et ekthetas in circuitu per tres partes contra uniuscuiusque limen stratumque ligno per gyrum in circuitu terra autem usque ad fenestras et fenestrae clausae super ostia
EZEK|41|17|et usque ad domum interiorem et forinsecus per omnem parietem in circuitu intrinsecus et forinsecus ad mensuram
EZEK|41|18|et fabrefacta cherubin et palmae et palma inter cherub et cherub duasque facies habebat cherub
EZEK|41|19|faciem hominis iuxta palmam ex hac parte et faciem leonis iuxta palmam ex alia parte expressam per omnem domum in circuitu
EZEK|41|20|de terra usque ad superiora portae cherubin et palmae celatae erant in pariete templi
EZEK|41|21|limen quadrangulum et facies sanctuarii aspectus contra aspectum
EZEK|41|22|altaris lignei trium cubitorum altitudo et longitudo eius duo cubitorum et anguli eius et longitudo eius et parietes eius lignei et locutus est ad me haec est mensa coram Domino
EZEK|41|23|et duo ostia erant in templo et in sanctuario
EZEK|41|24|et in duobus ostiis ex utraque parte bina erant ostiola quae in se invicem plicabantur bina enim ostia erant ex utraque parte ostiorum
EZEK|41|25|et celata erant in ipsis ostiis templi cherubin et scalptura palmarum sicut in parietibus quoque expressa erat quam ob rem erant et grossiora ligna in vestibuli fronte forinsecus
EZEK|41|26|super quae fenestrae obliquae et similitudo palmarum hinc atque inde in umerulis vestibuli secundum latera domus latitudinemque parietum
EZEK|42|1|et eduxit me in atrium exterius per viam ducentem ad aquilonem et eduxit me in gazofilacium quod erat contra separatum aedificium et contra aedem vergentem ad aquilonem
EZEK|42|2|in facie longitudinis centum cubitos ostii aquilonis et latitudinis quinquaginta cubitos
EZEK|42|3|contra viginti cubitos atrii interioris et contra pavimentum stratum lapide atrii exterioris ubi erat porticus iuncta porticui triplici
EZEK|42|4|et ante gazofilacia deambulatio decem cubitorum latitudinis ad interiora respiciens viae cubiti unius et ostia earum ad aquilonem
EZEK|42|5|ubi erant gazofilacia in superioribus humiliora quia subportabant porticus quae ex illis eminebant de inferioribus et de mediis aedificii
EZEK|42|6|tristega enim erant et non habebant columnas sicut erant columnae atriorum propterea eminebant de inferioribus et de mediis a terra
EZEK|42|7|et peribolus exterior secundum gazofilacia quae erant in via atrii exterioris ante gazofilacia longitudo eius quinquaginta cubitorum
EZEK|42|8|quia longitudo erat gazofilaciorum atrii exterioris quinquaginta cubitorum et longitudo ante faciem templi centum cubitorum
EZEK|42|9|et erat subter gazofilacia haec introitus ab oriente ingredientium in ea de atrio exteriori
EZEK|42|10|in latitudine periboli atrii quod erat contra viam orientalem in facie aedificii separati et erant ante aedificium gazofilacia
EZEK|42|11|et via ante faciem eorum iuxta similitudinem gazofilaciorum quae erant in via aquilonis secundum longitudinem eorum sic et latitudo eorum et omnis introitus eorum et similitudines et ostia eorum
EZEK|42|12|secundum ostia gazofilaciorum quae erant in via respiciente ad notum ostium in capite viae quae via erat ante vestibulum separatum per viam orientalem ingredientibus
EZEK|42|13|et dixit ad me gazofilacia aquilonis et gazofilacia austri quae sunt ante aedificium separatum haec sunt gazofilacia sancta in quibus vescuntur sacerdotes qui adpropinquant ad Dominum in sancta sanctorum ibi ponent sancta sanctorum et oblationem pro peccato et pro delicto locus enim sanctus est
EZEK|42|14|cum autem ingressi fuerint sacerdotes non egredientur de sanctis in atrium exterius et ibi reponent vestimenta sua in quibus ministrant quia sancta sunt vestienturque vestimentis aliis et sic procedent ad populum
EZEK|42|15|cumque conplesset mensuras domus interioris eduxit me per viam portae quae respiciebat ad viam orientalem et mensus est eam undique per circuitum
EZEK|42|16|mensus autem est contra ventum orientalem calamo mensurae quingentos calamos in calamo mensurae per circuitum
EZEK|42|17|et mensus est contra ventum aquilonem quingentos calamos in calamo mensurae per gyrum
EZEK|42|18|et ad ventum australem mensus est quingentos calamos in calamo mensurae per circuitum
EZEK|42|19|et ad ventum occidentalem mensus est quingentos calamos in calamo mensurae
EZEK|42|20|per quattuor ventos mensus est illud murum eius undique per circuitum longitudine quingentorum cubitorum et latitudine quingentorum cubitorum dividentem inter sanctuarium et vulgi locum
EZEK|43|1|et duxit me ad portam quae respiciebat ad viam orientalem
EZEK|43|2|et ecce gloria Dei Israhel ingrediebatur per viam orientalem et vox erat ei quasi vox aquarum multarum et terra splendebat a maiestate eius
EZEK|43|3|et vidi visionem secundum speciem quam videram quando venit ut disperderet civitatem et species secundum aspectum quem videram iuxta fluvium Chobar et cecidi super faciem meam
EZEK|43|4|et maiestas Domini ingressa est templum per viam portae quae respiciebat ad orientem
EZEK|43|5|et levavit me spiritus et introduxit me in atrium interius et ecce repleta erat gloria Domini domus
EZEK|43|6|et audivi loquentem ad me de domo et vir qui stabat iuxta me
EZEK|43|7|dixit ad me fili hominis locus solii mei et locus vestigiorum pedum meorum ubi habito in medio filiorum Israhel in aeternum et non polluent ultra domus Israhel nomen sanctum meum ipsi et reges eorum in fornicationibus suis et in ruinis regum suorum et in excelsis
EZEK|43|8|qui fabricati sunt limen suum iuxta limen meum et postes suos iuxta postes meos et murus erat inter me et eos et polluerunt nomen sanctum meum in abominationibus quas fecerunt propter quod consumpsi eos in ira mea
EZEK|43|9|nunc ergo repellant procul fornicationem suam et ruinas regum suorum a me et habitabo in medio eorum semper
EZEK|43|10|tu autem fili hominis ostende domui Israhel templum et confundantur ab iniquitatibus suis et metiantur fabricam
EZEK|43|11|et erubescant ex omnibus quae fecerunt figuram domus et fabricae eius exitus et introitus et omnem descriptionem eius et universa praecepta eius cunctumque ordinem eius et omnes leges eius ostende eis et scribes in oculis eorum et custodiant omnes descriptiones eius et praecepta illius et faciant ea
EZEK|43|12|ista est lex domus in summitate montis omnes fines eius in circuitu sanctum sanctorum est haec ergo est lex domus
EZEK|43|13|istae autem mensurae altaris in cubito verissimo qui habebat cubitum et palmum in sinu eius erat cubitus et cubitus in latitudine et definitio usque ad labium eius in circuitu palmus unus haec quoque erat fossa altaris
EZEK|43|14|et de sinu terrae usque ad crepidinem novissimam duo cubiti et latitudo cubiti unius et a crepidine maiori usque ad crepidinem minorem quattuor cubiti et latitudo unius cubiti
EZEK|43|15|ipse autem arihel quattuor cubitorum et ab arihel usque sursum cornua quattuor
EZEK|43|16|et arihel duodecim cubitorum in longitudine per duodecim cubitos latitudinis quadrangulatum aequis lateribus
EZEK|43|17|et crepido quattuordecim cubitorum longitudinis per quattuordecim latitudinis in quattuor angulis eius et corona in circuitu eius dimidii cubitus et sinus eius unius cubiti per circuitum gradus autem eius versi ad orientem
EZEK|43|18|et dixit ad me fili hominis haec dicit Dominus Deus hii sunt ritus altaris in quacumque die fuerit fabricatum ut offeratur super illud holocaustum et effundatur sanguis
EZEK|43|19|et dabis sacerdotibus Levitis qui sunt de semine Sadoc qui accedunt ad me ait Dominus Deus ut offerant mihi vitulum de armento pro peccato
EZEK|43|20|et adsumens de sanguine eius pones super quattuor cornua eius et super quattuor angulos crepidinis et super coronam in circuitu et mundabis illud et expiabis
EZEK|43|21|et tolles vitulum qui oblatus fuerit pro peccato et conbures illum in separato loco domus extra sanctuarium
EZEK|43|22|et in die secunda offeres hircum caprarum inmaculatum pro peccato et expiabunt altare sicut expiaverunt in vitulo
EZEK|43|23|cumque conpleveris expians illud offeres vitulum de armento inmaculatum et arietem de grege inmaculatum
EZEK|43|24|et offeres eos in conspectu Domini et mittent sacerdotes super eos sal et offerent eos holocaustum Domino
EZEK|43|25|septem diebus facies hircum pro peccato cotidie et vitulum de armento et arietem de pecoribus inmaculatos offerent
EZEK|43|26|septem diebus expiabunt altare et mundabunt illud et implebunt manum eius
EZEK|43|27|expletis autem diebus in die octava et ultra facient sacerdotes super altare holocausta vestra et quae pro pace offerunt et placatus ero vobis ait Dominus Deus
EZEK|44|1|et convertit me ad viam portae sanctuarii exterioris quae respiciebat ad orientem et erat clausa
EZEK|44|2|et dixit Dominus ad me porta haec clausa erit non aperietur et vir non transiet per eam quoniam Dominus Deus Israhel ingressus est per eam eritque clausa
EZEK|44|3|principi princeps ipse sedebit in ea ut comedat panem coram Domino per viam vestibuli portae ingredietur et per viam eius egredietur
EZEK|44|4|et adduxit me per viam portae aquilonis in conspectu domus et vidi et ecce implevit gloria Domini domum Domini et cecidi in faciem meam
EZEK|44|5|et dixit ad me Dominus fili hominis pone cor tuum et vide oculis tuis et auribus tuis audi omnia quae ego loquor ad te de universis caerimoniis domus Domini et de cunctis legibus eius et pones cor tuum in viis templi per omnes exitus sanctuarii
EZEK|44|6|et dices ad exasperantem me domum Israhel haec dicit Dominus Deus sufficiant vobis omnia scelera vestra domus Israhel
EZEK|44|7|eo quod inducitis filios alienos incircumcisos corde et incircumcisos carne ut sint in sanctuario meo et polluant domum meam et offertis panes meos adipem et sanguinem et dissolvitis pactum meum in omnibus sceleribus vestris
EZEK|44|8|et non servastis praecepta sanctuarii mei et posuistis custodes observationum mearum in sanctuario meo vobismet ipsis
EZEK|44|9|haec dicit Dominus Deus omnis alienigena incircumcisus corde et incircumcisus carne non ingredietur sanctuarium meum omnis filius alienus qui est in medio filiorum Israhel
EZEK|44|10|sed et Levitae qui longe recesserunt a me in errore filiorum Israhel et erraverunt a me post idola sua et portaverunt iniquitatem suam
EZEK|44|11|erunt in sanctuario meo aeditui et ianitores portarum domus et ministri domus ipsi mactabunt holocaustosin et victimas populi et ipsi stabunt in conspectu eorum ut ministrent eis
EZEK|44|12|pro eo quod ministraverunt illis in conspectu idolorum suorum et facti sunt domui Israhel in offendiculum iniquitatis idcirco levavi manum meam super eos dicit Dominus Deus et portaverunt iniquitatem suam
EZEK|44|13|et non adpropinquabunt ad me ut sacerdotio fungantur mihi neque accedent ad omne sanctuarium meum iuxta sancta sanctorum sed portabunt confusionem suam et scelera sua quae fecerunt
EZEK|44|14|et dabo eos ianitores domus in omni ministerio eius et universis quae fiunt in ea
EZEK|44|15|sacerdotes autem Levitae filii Sadoc qui custodierunt caerimonias sanctuarii mei cum errarent filii Israhel a me ipsi accedent ad me ut ministrent mihi et stabunt in conspectu meo ut offerant mihi adipem et sanguinem ait Dominus Deus
EZEK|44|16|ipsi ingredientur sanctuarium meum et ipsi accedent ad mensam meam ut ministrent mihi et custodiant caerimonias meas
EZEK|44|17|cumque ingredientur portas atrii interioris vestibus lineis induentur nec ascendet super eos quicquam laneum quando ministrant in portis atrii interioris et intrinsecus
EZEK|44|18|vittae lineae erunt in capitibus eorum et feminalia linea erunt in lumbis eorum et non accingentur in sudore
EZEK|44|19|cumque egredientur atrium exterius ad populum exuent se vestimenta sua in quibus ministraverunt et reponent ea in gazofilacio sanctuarii et vestient se vestimentis aliis et non sanctificabunt populum in vestibus suis
EZEK|44|20|caput autem suum non radent neque comam nutrient sed tondentes adtondent capita sua
EZEK|44|21|et vinum non bibet omnis sacerdos quando ingressurus est atrium interius
EZEK|44|22|et viduam et repudiatam non accipient uxores sed virgines de semine domus Israhel sed et viduam quae fuerit vidua a sacerdote accipient
EZEK|44|23|et populum meum docebunt quid sit inter sanctum et pollutum et inter mundum et inmundum ostendent eis
EZEK|44|24|et cum fuerit controversia stabunt in iudiciis meis et iudicabunt leges meas et praecepta mea in omnibus sollemnitatibus meis custodient et sabbata mea sanctificabunt
EZEK|44|25|et ad mortuum hominem non ingredientur ne polluantur nisi ad patrem et matrem et filium et filiam et fratrem et sororem quae alterum virum non habuit in quibus contaminabuntur
EZEK|44|26|et postquam fuerit emundatus septem dies numerabuntur ei
EZEK|44|27|et in die introitus sui in sanctuarium ad atrium interius ut ministret mihi in sanctuario offeret pro peccato suo ait Dominus Deus
EZEK|44|28|erit autem eis hereditas ego hereditas eorum et possessionem non dabitis eis in Israhel ego enim possessio eorum
EZEK|44|29|victimam et pro peccato et pro delicto ipsi comedent et omne votum in Israhel ipsorum erit
EZEK|44|30|et primitiva omnium primogenitorum et omnia libamenta ex omnibus quae offeruntur sacerdotum erunt et primitiva ciborum vestrorum dabitis sacerdoti ut reponat benedictionem domui suae
EZEK|44|31|omne morticinum et captum a bestia de avibus et de pecoribus non comedent sacerdotes
EZEK|45|1|cumque coeperitis terram dividere sortito separate primitias Domino sanctificatum de terra longitudine viginti quinque milia et latitudine decem milia sanctificatum erit in omni termino eius per circuitum
EZEK|45|2|et erit ex omni parte sanctificatum quingentos per quingentos quadrifariam per circuitum et quinquaginta cubitis in suburbana eius per gyrum
EZEK|45|3|et a mensura ista mensurabis longitudinem viginti quinque milium et latitudinem decem milium et in ipso erit templum sanctumque sanctorum
EZEK|45|4|sanctificatum de terra erit sacerdotibus ministris sanctuarii qui accedunt ad ministerium Domini et erit eis locus in domos et in sanctuarium sanctitatis
EZEK|45|5|viginti quinque autem milia longitudinis et decem milia latitudinis erunt Levitis qui ministrant domui ipsi possidebunt viginti gazofilacia
EZEK|45|6|et possessionem civitatis dabitis quinque milia latitudinis et longitudinis viginti quinque milia secundum separationem sanctuarii omni domui Israhel
EZEK|45|7|principi quoque hinc et inde in separationem sanctuarii et in possessionem civitatis contra faciem separationis sanctuarii et contra faciem possessionis urbis a latere maris usque ad mare et a latere orientis usque ad orientem longitudinem autem iuxta unamquamque partium a termino occidentali usque ad terminum orientalem
EZEK|45|8|de terra erit ei possessio in Israhel et non depopulabuntur ultra principes populum meum sed terram dabunt domui Israhel secundum tribus eorum
EZEK|45|9|haec dicit Dominus Deus sufficiat vobis principes Israhel iniquitatem et rapinas intermittite et iudicium et iustitiam facite separate confinia vestra a populo meo ait Dominus Deus
EZEK|45|10|statera iusta et oephi iustum et batus iustus erit vobis
EZEK|45|11|oephi et batus aequalia et unius mensurae erunt ut capiat decimam partem chori batus et decimam partem chori oephi iuxta mensuram chori erit aequa libratio eorum
EZEK|45|12|siclus autem viginti obolos habeat porro viginti sicli et viginti quinque sicli et quindecim sicli minam facient
EZEK|45|13|et haec sunt primitiae quas tolletis sextam partem oephi de choro frumenti et sextam partem oephi de choro hordei
EZEK|45|14|mensura quoque olei batus olei decima pars chori est et decem bati chorum faciunt quia decem bati implent chorum
EZEK|45|15|et arietem unum de grege ducentorum de his quae nutriunt Israhel in sacrificium et in holocaustum et in pacifica ad expiandum pro eis ait Dominus Deus
EZEK|45|16|omnis populus terrae tenebitur primitiis his principi in Israhel
EZEK|45|17|et super principem erunt holocausta et sacrificium et libamina in sollemnitatibus et in kalendis et in sabbatis in universis sollemnitatibus domus Israhel ipse faciat pro peccato sacrificium et holocaustum et pacifica ad expiandum pro domo Israhel
EZEK|45|18|haec dicit Dominus Deus in primo mense una mensis sumes vitulum de armento inmaculatum et expiabis sanctuarium
EZEK|45|19|et tollet sacerdos de sanguine quod erit pro peccato et ponet in postibus domus et in quattuor angulis crepidinis altaris et in postibus portae atrii interioris
EZEK|45|20|et sic facies in septima mensis pro unoquoque qui ignoravit et errore deceptus est et expiabitis pro domo
EZEK|45|21|in primo mense quartadecima die mensis erit vobis paschae sollemnitas septem diebus azyma comedentur
EZEK|45|22|et faciet princeps in die illa pro se et pro universo populo terrae vitulum pro peccato
EZEK|45|23|et in septem dierum sollemnitate faciet holocaustum Domino septem vitulos et septem arietes inmaculatos cotidie septem diebus et pro peccato hircum caprarum cotidie
EZEK|45|24|et sacrificium oephi per vitulum et oephi per arietem faciet et olei hin per singula oephi
EZEK|45|25|septimo mense quintadecima die mensis in sollemnitate faciet sicut supra dicta sunt per septem dies tam pro peccato quam pro holocausto et in sacrificio et in oleo
EZEK|46|1|haec dicit Dominus Deus porta atrii interioris quae respicit ad orientem erit clausa sex diebus in quibus opus fit die autem sabbati aperietur sed et in die kalendarum aperietur
EZEK|46|2|et intrabit princeps per viam vestibuli portae de foris et stabit in limine portae et facient sacerdotes holocaustum eius et pacifica eius et adorabit super limen portae et egredietur porta autem non claudetur usque ad vesperam
EZEK|46|3|et adorabit populus terrae ad ostium portae illius in sabbatis et in kalendis coram Domino
EZEK|46|4|holocaustum autem hoc offeret princeps Domino in die sabbati sex agnos inmaculatos et arietem inmaculatum
EZEK|46|5|et sacrificium oephi per arietem agnis autem sacrificium quod dederit manus eius et olei hin per singula oephi
EZEK|46|6|in die autem kalendarum vitulum de armento inmaculatum et sex agni et arietes inmaculati erunt
EZEK|46|7|et oephi per vitulum oephi quoque per arietem faciet sacrificium agnis autem sicut invenerit manus eius et olei hin per singula oephi
EZEK|46|8|cumque ingressurus est princeps per viam vestibuli portae ingrediatur et per eandem viam exeat
EZEK|46|9|et cum intrabit populus terrae in conspectu Domini in sollemnitatibus qui ingreditur per portam aquilonis ut adoret egrediatur per viam portae meridianae porro qui ingreditur per viam portae meridianae egrediatur per viam portae aquilonis non revertetur per viam portae per quam ingressus est sed e regione illius egredietur
EZEK|46|10|princeps autem in medio eorum cum ingredientibus ingredietur et cum egredientibus egredietur
EZEK|46|11|et in nundinis et in sollemnitatibus erit sacrificium oephi per vitulum et oephi per arietem agnis autem erit sacrificium sicut invenerit manus eius et olei hin per singula oephi
EZEK|46|12|cum autem fecerit princeps spontaneum holocaustum aut pacifica voluntaria Domino aperietur ei porta quae respicit ad orientem et faciet holocaustum suum et pacifica sua sicut fieri solet in die sabbati et egredietur claudeturque porta postquam exierit
EZEK|46|13|et agnum eiusdem anni inmaculatum faciet holocaustum cotidie Domino semper mane faciet illud
EZEK|46|14|et sacrificium faciet super eo cata mane mane sextam partem oephi et de oleo tertiam partem hin ut misceatur similae sacrificium Domino legitimum iuge atque perpetuum
EZEK|46|15|faciet agnum et sacrificium et oleum cata mane mane holocaustum sempiternum
EZEK|46|16|haec dicit Dominus Deus si dederit princeps donum alicui de filiis suis hereditas eius filiorum suorum erit possidebunt ea hereditarie
EZEK|46|17|si autem dederit legatum de hereditate sua uni servorum suorum erit illius usque ad annum remissionis et revertetur ad principem hereditas autem eius filiis eius erit
EZEK|46|18|et non accipiet princeps de hereditate populi per violentiam et de possessione eorum sed de possessione sua hereditatem dabit filiis suis ut non dispergatur populus meus unusquisque a possessione sua
EZEK|46|19|et introduxit me per ingressum qui erat ex latere portae in gazofilacia sanctuarii ad sacerdotes quae respiciebant ad aquilonem et erat ibi locus vergens ad occidentem
EZEK|46|20|et dixit ad me iste est locus ubi coquent sacerdotes pro delicto et pro peccato ubi coquent sacrificium ut non efferant in atrio exteriori et sanctificetur populus
EZEK|46|21|et eduxit me in atrium exterius et circumduxit me per quattuor angulos atrii et ecce atriolum erat in angulo atrii atriola singula per angulos atrii
EZEK|46|22|in quattuor angulos atrii atriola disposita quadraginta cubitorum per longum et triginta per latum mensurae unius quattuor erant
EZEK|46|23|et paries per circuitum ambiens quattuor atriola et culinae fabricatae erant subter porticus per gyrum
EZEK|46|24|et dixit ad me haec est domus culinarum in qua coquent ministri domus Domini victimas populi
EZEK|47|1|et convertit me ad portam domus et ecce aquae egrediebantur subter limen domus ad orientem facies enim domus respiciebat ad orientem aquae autem descendebant in latus templi dextrum ad meridiem altaris
EZEK|47|2|et eduxit me per viam portae aquilonis et convertit me ad viam foras portam exteriorem viam quae respiciebat ad orientem et ecce aquae redundantes a latere dextro
EZEK|47|3|cum egrederetur vir ad orientem qui habebat funiculum in manu sua et mensus est mille cubitos et transduxit me per aquam usque ad talos
EZEK|47|4|rursumque mensus est mille et transduxit me per aquam usque ad genua
EZEK|47|5|et mensus est mille et transduxit me per aquam usque ad renes et mensus est mille torrentem quem non potui pertransire quoniam intumuerant aquae profundae torrentis qui non potest transvadari
EZEK|47|6|et dixit ad me certe vidisti fili hominis et duxit me et convertit ad ripam torrentis
EZEK|47|7|cumque me convertissem ecce in ripa torrentis ligna multa nimis ex utraque parte
EZEK|47|8|et ait ad me aquae istae quae egrediuntur ad tumulos sabuli orientalis et descendunt ad plana deserti intrabunt mare et exibunt et sanabuntur aquae
EZEK|47|9|et omnis anima vivens quae serpit quocumque venerit torrens vivet et erunt pisces multi satis postquam venerint illuc aquae istae et sanabuntur et vivent omnia ad quae venerit torrens
EZEK|47|10|vivent et stabunt super illa piscatores ab Engaddi usque ad Engallim siccatio sagenarum erunt plurimae species erunt piscium eius sicut pisces maris magni multitudinis nimiae
EZEK|47|11|in litoribus autem eius et in palustribus non sanabuntur quia in salinas dabuntur
EZEK|47|12|et super torrentem orietur in ripis eius ex utraque parte omne lignum pomiferum non defluet folium ex eo et non deficiet fructus eius per singulos menses adferet primitiva quia aquae eius de sanctuario egredientur et erunt fructus eius in cibum et folia eius ad medicinam
EZEK|47|13|haec dicit Dominus Deus hic est terminus in quo possidebitis terram in duodecim tribubus Israhel quia Ioseph duplicem funiculum habet
EZEK|47|14|possidebitis autem eam singuli aeque ut frater suus quam levavi manum meam ut darem patribus vestris et cadet terra haec vobis in possessionem
EZEK|47|15|hic est autem terminus terrae ad plagam septentrionalem a mari magno via Bethalon venientibus Sadada
EZEK|47|16|Emath Berotha Sabarim quae est inter terminum Damasci et confinium Emath domus Atticon quae est iuxta terminos Auran
EZEK|47|17|et erit terminus a mari usque ad atrium Aenon terminus Damasci et ab aquilone ad aquilonem et terminus Emath plaga autem septentrionalis
EZEK|47|18|porro plaga orientalis de medio Auran et de medio Damasci et de medio Galaad et de medio terrae Israhel Iordanis disterminans ad mare orientale metiemini etiam plagam orientalem
EZEK|47|19|plaga autem australis meridiana a Thamar usque ad aquas Contradictionis Cades et torrens usque ad mare magnum et plaga ad meridiem australis
EZEK|47|20|et plaga maris mare magnum a confinio per directum donec venias Emath haec est plaga maris
EZEK|47|21|et dividetis terram istam vobis per tribus Israhel
EZEK|47|22|et mittetis eam in hereditatem vobis et advenis qui accesserint ad vos qui genuerint filios in medio vestrum et erunt vobis sicut indigenae inter filios Israhel vobiscum divident possessionem in medio tribuum Israhel
EZEK|47|23|in tribu autem quacumque fuerit advena ibi dabitis possessionem illi ait Dominus Deus
EZEK|48|1|et haec nomina tribuum a finibus aquilonis iuxta viam Aethlon pergentibus Emath atrium Aenon terminus Damasci ad aquilonem iuxta Emath et erit ei plaga orientalis mare Dan una
EZEK|48|2|et ad terminum Dan a plaga orientali usque ad plagam maris Aser una
EZEK|48|3|et super terminum Aser a plaga orientali usque ad plagam maris Nepthalim una
EZEK|48|4|et super terminum Nepthalim a plaga orientali usque ad plagam maris Manasse una
EZEK|48|5|et super terminum Manasse a plaga orientali usque ad plagam maris Ephraim una
EZEK|48|6|et super terminum Ephraim a plaga orientali usque ad plagam maris Ruben una
EZEK|48|7|et super terminum Ruben a plaga orientali usque ad plagam maris Iuda una
EZEK|48|8|et super terminum Iuda a plaga orientali usque ad plagam maris erunt primitiae quas separabitis viginti quinque milibus latitudinis et longitudinis sicuti singulae partes a plaga orientali usque ad plagam maris et erit sanctuarium in medio eius
EZEK|48|9|primitiae quas separastis Domino longitudo viginti quinque milibus et latitudo decem milibus
EZEK|48|10|hae autem erunt primitiae sanctuarii sacerdotum ad aquilonem viginti quinque milia et ad mare latitudinis decem milia sed et ad orientem latitudinis decem milia et ad meridiem longitudinis viginti quinque milia et erit sanctuarium Domini in medio eius
EZEK|48|11|sacerdotibus sanctuarium erit de filiis Sadoc qui custodierunt caerimonias meas et non erraverunt cum errarent filii Israhel sicut erraverunt et Levitae
EZEK|48|12|et erunt eis primitiae de primitiis terrae sanctum sanctorum iuxta terminum Levitarum
EZEK|48|13|sed et Levitis similiter iuxta fines sacerdotum viginti quinque milia longitudinis et latitudinis decem milia omnis longitudo viginti et quinque milium et latitudo decem milium
EZEK|48|14|et non venundabunt ex eo neque mutabunt nec transferentur primitiae terrae quia sanctificatae sunt Domino
EZEK|48|15|quinque milia autem quae supersunt in latitudine per viginti quinque milia profana erunt urbis in habitaculum et in suburbana et erit civitas in medio eius
EZEK|48|16|et heae mensurae eius ad plagam septentrionalem quingenti et quattuor milia et ad plagam meridianam quingenti et quattuor milia et ad plagam orientalem quingenti et quattuor milia et ad plagam occidentalem quingenti et quattuor milia
EZEK|48|17|erunt autem suburbana civitatis ad aquilonem ducenti quinquaginta et in meridie ducenti quinquaginta et ad orientem ducenti quinquaginta et ad mare ducenti quinquaginta
EZEK|48|18|quod autem reliquum fuerit in longitudine secundum primitias sanctuarii decem milia in orientem et decem milia ad occidentem erunt sicut primitiae sanctuarii et erunt fruges eius in panes his qui serviunt civitati
EZEK|48|19|servientes autem civitati operabuntur ex omnibus tribubus Israhel
EZEK|48|20|omnes primitiae viginti quinque milium per viginti quinque milia in quadrum separabuntur in primitias sanctuarii et possessionem civitatis
EZEK|48|21|quod autem reliquum fuerit principis erit ex omni parte primitiarum sanctuarii et possessionis civitatis e regione viginti quinque milium primitiarum usque ad terminum orientalem sed et ad mare e regione viginti quinque milium usque ad terminum maris similiter in partibus principis erit et erunt primitiae sanctuarii et sanctuarium templi in medio eius
EZEK|48|22|de possessione autem Levitarum et de possessione civitatis in medio partium principis erit inter terminum Iuda et inter terminum Beniamin et ad principem pertinebit
EZEK|48|23|et reliquis tribubus a plaga orientali usque ad plagam occidentalem Beniamin una
EZEK|48|24|et contra terminum Beniamin a plaga orientali usque ad plagam occidentalem Symeon una
EZEK|48|25|et super terminum Symeonis a plaga orientali usque ad plagam occidentis Isachar una
EZEK|48|26|et super terminum Isachar a plaga orientali usque ad plagam occidentalem Zabulon una
EZEK|48|27|et super terminum Zabulon a plaga orientali usque ad plagam maris Gad una
EZEK|48|28|et super terminum Gad ad plagam austri in meridiem et erit finis de Thamar usque ad aquas Contradictionis Cades hereditas contra mare magnum
EZEK|48|29|haec est terra quam mittetis in sortem tribubus Israhel et hae partitiones earum ait Dominus Deus
EZEK|48|30|et hii egressus civitatis a plaga septentrionali quingentos et quattuor milia mensurabis
EZEK|48|31|et portae civitatis in nominibus tribuum Israhel portae tres a septentrione porta Ruben una porta Iudae una porta Levi una
EZEK|48|32|et ad plagam orientalem quingentos et quattuor milia et portae tres porta Ioseph una porta Beniamin una porta Dan una
EZEK|48|33|et ad plagam meridianam quingentos et quattuor milia metieris portam Symeonis unam portam Isachar unam portam Zabulon unam
EZEK|48|34|et ad plagam occidentalem quingenti et quattuor milia portae eorum tres porta Gad una porta Aser una porta Nepthalim una
EZEK|48|35|per circuitum decem et octo milia et nomen civitatis ex illa die Dominus ibidem
DAN|1|1|anno tertio regni Ioachim regis Iuda venit Nabuchodonosor rex Babylonis Hierusalem et obsedit eam
DAN|1|2|et tradidit Dominus in manu eius Ioachim regem Iudae et partem vasorum domus Dei et asportavit ea in terram Sennaar in domum dei sui et vasa intulit in domum thesauri dei sui
DAN|1|3|et ait rex Asfanaz praeposito eunuchorum suorum ut introduceret de filiis Israhel et de semine regio et tyrannorum
DAN|1|4|pueros in quibus nulla esset macula decoros forma et eruditos omni sapientia cautos scientia et doctos disciplina et qui possent stare in palatio regis ut doceret eos litteras et linguam Chaldeorum
DAN|1|5|et constituit eis rex annonam per singulos dies de cibis suis et de vino unde bibebat ipse ut enutriti tribus annis postea starent in conspectu regis
DAN|1|6|fuerunt ergo inter eos de filiis Iuda Danihel Ananias Misahel et Azarias
DAN|1|7|et inposuit eis praepositus eunuchorum nomina Daniheli Balthasar et Ananiae Sedrac Misaheli Misac et Azariae Abdenago
DAN|1|8|proposuit autem Danihel in corde suo ne pollueretur de mensa regis neque de vino potus eius et rogavit eunuchorum praepositum ne contaminaretur
DAN|1|9|dedit autem Deus Daniheli gratiam et misericordiam in conspectu principis eunuchorum
DAN|1|10|et ait princeps eunuchorum ad Danihel timeo ego dominum meum regem qui constituit vobis cibum et potum qui si viderit vultus vestros macilentiores prae ceteris adulescentibus coaevis vestris condemnabitis caput meum regi
DAN|1|11|et dixit Danihel ad Malassar quem constituerat princeps eunuchorum super Danihel Ananiam Misahel et Azariam
DAN|1|12|tempta nos obsecro servos tuos diebus decem et dentur nobis legumina ad vescendum et aqua ad bibendum
DAN|1|13|et contemplare vultus nostros et vultus puerorum qui vescuntur cibo regio et sicut videris facies cum servis tuis
DAN|1|14|qui audito sermone huiuscemodi temptavit eos diebus decem
DAN|1|15|post dies autem decem apparuerunt vultus eorum meliores et corpulentiores prae omnibus pueris qui vescebantur cibo regio
DAN|1|16|porro Malassar tollebat cibaria et vinum potus eorum dabatque eis legumina
DAN|1|17|pueris autem his dedit Deus scientiam et disciplinam in omni libro et sapientia Daniheli autem intellegentiam omnium visionum et somniorum
DAN|1|18|conpletis itaque diebus post quos dixerat rex ut introducerentur introduxit eos praepositus eunuchorum in conspectu Nabuchodonosor
DAN|1|19|cumque locutus eis fuisset rex non sunt inventi de universis tales ut Danihel Ananias Misahel et Azarias et steterunt in conspectu regis
DAN|1|20|et omne verbum sapientiae et intellectus quod sciscitatus est ab eis rex invenit in eis decuplum super cunctos ariolos et magos qui erant in universo regno eius
DAN|1|21|fuit autem Danihel usque ad annum primum Cyri regis
DAN|2|1|in anno secundo regni Nabuchodonosor vidit Nabuchodonosor somnium et conterritus est spiritus eius et somnium eius fugit ab eo
DAN|2|2|praecepit ergo rex ut convocarentur arioli et magi et malefici et Chaldei et indicarent regi somnia sua qui cum venissent steterunt coram rege
DAN|2|3|et dixit ad eos rex vidi somnium et mente confusus ignoro quid viderim
DAN|2|4|responderuntque Chaldei regi syriace rex in sempiternum vive dic somnium servis tuis et interpretationem eius indicabimus
DAN|2|5|et respondens rex ait Chaldeis sermo recessit a me nisi indicaveritis mihi somnium et coniecturam eius peribitis vos et domus vestrae publicabuntur
DAN|2|6|si autem somnium et coniecturam eius narraveritis praemia et dona et honorem multum accipietis a me somnium igitur et interpretationem eius indicate mihi
DAN|2|7|responderunt secundo atque dixerunt rex somnium dicat servis suis et interpretationem illius indicabimus
DAN|2|8|respondit rex et ait certo novi quia tempus redimitis scientes quod recesserit a me sermo
DAN|2|9|si ergo somnium non indicaveritis mihi una est de vobis sententia quod interpretationem quoque fallacem et deceptione plenam conposueritis ut loquamini mihi donec tempus pertranseat somnium itaque dicite mihi ut sciam quod interpretationem quoque eius veram loquamini
DAN|2|10|respondentes ergo Chaldei coram rege dixerunt non est homo super terram qui sermonem tuum rex possit implere sed neque regum quisquam magnus et potens verbum huiuscemodi sciscitatur ab omni ariolo et mago et Chaldeo
DAN|2|11|sermo enim quem tu rex quaeris gravis est nec repperietur quisquam qui indicet illum in conspectu regis exceptis diis quorum non est cum hominibus conversatio
DAN|2|12|quo audito rex in furore et in ira magna praecepit ut perirent omnes sapientes Babylonis
DAN|2|13|et egressa sententia sapientes interficiebantur quaerebaturque Danihel et socii eius ut perirent
DAN|2|14|tunc Danihel requisivit de lege atque sententia ab Arioch principe militiae regis qui egressus fuerat ad interficiendos sapientes Babylonis
DAN|2|15|et interrogavit eum qui a rege acceperat potestatem quam ob causam tam crudelis sententia a facie esset regis egressa cum ergo rem indicasset Arioch Daniheli
DAN|2|16|Danihel ingressus rogavit regem ut tempus daret sibi ad solutionem indicandam regi
DAN|2|17|et ingressus est domum suam Ananiaeque Misaheli et Azariae sociis suis indicavit negotium
DAN|2|18|ut quaererent misericordiam a facie Dei caeli super sacramento isto et non perirent Danihel et socii eius cum ceteris sapientibus Babylonis
DAN|2|19|tunc Daniheli per visionem nocte mysterium revelatum est et Danihel benedixit Deo caeli
DAN|2|20|et locutus ait sit nomen Domini benedictum a saeculo et usque in saeculum quia sapientia et fortitudo eius sunt
DAN|2|21|et ipse mutat tempora et aetates transfert regna atque constituit dat sapientiam sapientibus et scientiam intellegentibus disciplinam
DAN|2|22|ipse revelat profunda et abscondita et novit in tenebris constituta et lux cum eo est
DAN|2|23|tibi Deus patrum meorum confiteor teque laudo quia sapientiam et fortitudinem dedisti mihi et nunc ostendisti mihi quae rogavimus te quia sermonem regis aperuisti nobis
DAN|2|24|post haec Danihel ingressus ad Arioch quem constituerat rex ut perderet sapientes Babylonis sic ei locutus est sapientes Babylonis ne perdas introduc me in conspectu regis et solutionem regi enarrabo
DAN|2|25|tunc Arioch festinus introduxit Danihelem ad regem et dixit ei inveni hominem de filiis transmigrationis Iudae qui solutionem regi adnuntiet
DAN|2|26|respondit rex et dixit Daniheli cuius nomen erat Balthasar putasne vere potes indicare mihi somnium quod vidi et interpretationem eius
DAN|2|27|et respondens Danihel coram rege ait mysterium quod rex interrogat sapientes magi et arioli et aruspices non queunt indicare regi
DAN|2|28|sed est Deus in caelo revelans mysteria qui indicavit tibi rex Nabuchodonosor quae ventura sunt novissimis temporibus somnium tuum et visiones capitis tui in cubili tuo huiuscemodi sunt
DAN|2|29|tu rex cogitare coepisti in stratu tuo quid esset futurum post haec et qui revelat mysteria ostendit tibi quae ventura sunt
DAN|2|30|mihi quoque non in sapientia quae est in me plus quam in cunctis viventibus sacramentum hoc revelatum est sed ut interpretatio regi manifesta fieret et cogitationes mentis tuae scires
DAN|2|31|tu rex videbas et ecce quasi statua una grandis statua illa magna et statura sublimis stabat contra te et intuitus eius erat terribilis
DAN|2|32|huius statuae caput ex auro optimo erat pectus autem et brachia de argento porro venter et femora ex aere
DAN|2|33|tibiae autem ferreae pedum quaedam pars erat ferrea quaedam fictilis
DAN|2|34|videbas ita donec abscisus est lapis sine manibus et percussit statuam in pedibus eius ferreis et fictilibus et comminuit eos
DAN|2|35|tunc contrita sunt pariter ferrum testa aes argentum et aurum et redacta quasi in favillam aestivae areae rapta sunt vento nullusque locus inventus est eis lapis autem qui percusserat statuam factus est mons magnus et implevit universam terram
DAN|2|36|hoc est somnium interpretationem quoque eius dicemus coram te rex
DAN|2|37|tu rex regum es et Deus caeli regnum fortitudinem et imperium et gloriam dedit tibi
DAN|2|38|et omnia in quibus habitant filii hominum et bestiae agri volucresque caeli dedit in manu tua et sub dicione tua universa constituit tu es ergo caput aureum
DAN|2|39|et post te consurget regnum aliud minus te et regnum tertium aliud aereum quod imperabit universae terrae
DAN|2|40|et regnum quartum erit velut ferrum quomodo ferrum comminuit et domat omnia sic comminuet omnia haec et conteret
DAN|2|41|porro quia vidisti pedum et digitorum partem testae figuli et partem ferream regnum divisum erit quod tamen de plantario ferri orietur secundum quod vidisti ferrum mixtum testae ex luto
DAN|2|42|et digitos pedum ex parte ferreos et ex parte fictiles ex parte regnum erit solidum et ex parte contritum
DAN|2|43|quia autem vidisti ferrum mixtum testae ex luto commiscebuntur quidem humano semine sed non adherebunt sibi sicuti ferrum misceri non potest testae
DAN|2|44|in diebus autem regnorum illorum suscitabit Deus caeli regnum quod in aeternum non dissipabitur et regnum eius populo alteri non tradetur comminuet et consumet universa regna haec et ipsum stabit in aeternum
DAN|2|45|secundum quod vidisti quod de monte abscisus est lapis sine manibus et comminuit testam et ferrum et aes et argentum et aurum Deus magnus ostendit regi quae futura sunt postea et verum est somnium et fidelis interpretatio eius
DAN|2|46|tunc rex Nabuchodonosor cecidit in faciem suam et Danihelum adoravit et hostias et incensum praecepit ut sacrificarent ei
DAN|2|47|loquens ergo rex ait Daniheli vere Deus vester Deus deorum est et Dominus regum et revelans mysteria quoniam potuisti aperire sacramentum hoc
DAN|2|48|tunc rex Danihelum in sublime extulit et munera multa et magna dedit ei et constituit eum principem super omnes provincias Babylonis et praefectum magistratuum super cunctos sapientes Babylonis
DAN|2|49|Danihel autem postulavit a rege et constituit super opera provinciae Babylonis Sedrac Misac et Abdenago ipse autem Danihel erat in foribus regis
DAN|3|1|Nabuchodonosor rex fecit statuam auream altitudine cubitorum sexaginta latitudine cubitorum sex et statuit eam in campo Duram provinciae Babylonis
DAN|3|2|itaque Nabuchodonosor rex misit ad congregandos satrapas magistratus et iudices duces et tyrannos et praefectos omnesque principes regionum ut convenirent ad dedicationem statuae quam erexerat Nabuchodonosor rex
DAN|3|3|tunc congregati sunt satrapae magistratus et iudices duces et tyranni et optimates qui erant in potestatibus constituti et universi principes regionum ut convenirent ad dedicationem statuae quam erexerat Nabuchodonosor rex stabant autem in conspectu statuae quam posuerat Nabuchodonosor
DAN|3|4|et praeco clamabat valenter vobis dicitur populis tribubus et linguis
DAN|3|5|in hora qua audieritis sonitum tubae et fistulae et citharae sambucae et psalterii et symphoniae et universi generis musicorum cadentes adorate statuam auream quam constituit Nabuchodonosor rex
DAN|3|6|si quis autem non prostratus adoraverit eadem hora mittetur in fornacem ignis ardentis
DAN|3|7|post haec igitur statim ut audierunt omnes populi sonitum tubae fistulae et citharae sambucae et psalterii et symphoniae et omnis generis musicorum cadentes omnes populi et tribus et linguae adoraverunt statuam auream quam constituerat Nabuchodonosor rex
DAN|3|8|statimque et in ipso tempore accedentes viri chaldei accusaverunt Iudaeos
DAN|3|9|dixeruntque Nabuchodonosor regi rex in aeternum vive
DAN|3|10|tu rex posuisti decretum ut omnis homo qui audierit sonitum tubae fistulae et citharae sambucae et psalterii et symphoniae et universi generis musicorum prosternat se et adoret statuam auream
DAN|3|11|si quis autem non procidens adoraverit mittatur in fornacem ignis ardentem
DAN|3|12|sunt ergo viri iudaei quos constituisti super opera regionis Babyloniae Sedrac Misac et Abdenago viri isti contempserunt rex decretum tuum deos tuos non colunt et statuam auream quam erexisti non adorant
DAN|3|13|tunc Nabuchodonosor in furore et in ira praecepit ut adducerentur Sedrac Misac et Abdenago qui confestim adducti sunt in conspectu regis
DAN|3|14|pronuntiansque Nabuchodonosor rex ait eis verene Sedrac Misac et Abdenago deos meos non colitis et statuam auream quam constitui non adoratis
DAN|3|15|nunc ergo si estis parati quacumque hora audieritis sonitum tubae fistulae et citharae sambucae psalterii et symphoniae omnisque generis musicorum prosternite vos et adorate statuam quam feci quod si non adoraveritis eadem hora mittemini in fornacem ignis ardentem et quis est Deus qui eripiat vos de manu mea
DAN|3|16|respondentes Sedrac Misac et Abdenago dixerunt regi Nabuchodonosor non oportet nos de hac re respondere tibi
DAN|3|17|ecce enim Deus noster quem colimus potest eripere nos de camino ignis ardentis et de manibus tuis rex liberare
DAN|3|18|quod si noluerit notum tibi sit rex quia deos tuos non colimus et statuam auream quam erexisti non adoramus
DAN|3|19|tunc Nabuchodonosor repletus est furore et aspectus faciei illius inmutatus est super Sedrac Misac et Abdenago et praecepit ut succenderetur fornax septuplum quam succendi consuerat
DAN|3|20|et viris fortissimis de exercitu suo iussit ut ligatis pedibus Sedrac Misac et Abdenago mitterent eos in fornacem ignis ardentem
DAN|3|21|et confestim viri illi vincti cum bracis suis et tiaris et calciamentis et vestibus missi sunt in medium fornacis ignis ardentis
DAN|3|22|nam iussio regis urguebat fornax autem succensa erat nimis porro viros illos qui miserant Sedrac Misac et Abdenago interfecit flamma ignis
DAN|3|23|viri autem hii id est tres Sedrac Misac et Abdenago ceciderunt in medio camini ignis ardentis conligati
DAN|3|24|et ambulabant in medio flammae laudantes Deum et benedicentes Domino
DAN|3|25|stans autem Azarias oravit sic aperiensque os suum in medio ignis ait
DAN|3|26|benedictus es Domine Deus patrum nostrorum et laudabilis et gloriosum nomen tuum in saecula
DAN|3|27|quia iustus es in omnibus quae fecisti nobis et universa opera tua vera et viae tuae rectae et omnia iudicia tua vera
DAN|3|28|iudicia enim vera fecisti iuxta omnia quae induxisti super nos et super civitatem sanctam patrum nostrorum Hierusalem quia in veritate et in iudicio induxisti omnia haec propter peccata nostra
DAN|3|29|peccavimus enim et inique egimus recedentes a te et deliquimus in omnibus
DAN|3|30|et praecepta tua non audivimus nec observavimus nec fecimus sicut praeceperas nobis ut bene nobis esset
DAN|3|31|omnia ergo quae induxisti super nos et universa quae fecisti nobis vero iudicio fecisti
DAN|3|32|et tradidisti nos in manibus inimicorum iniquorum et pessimorum praevaricatorumque et regi iniusto et pessimo ultra omnem terram
DAN|3|33|et nunc non possumus aperire os confusio et obprobrium facti sumus servis tuis et his qui colunt te
DAN|3|34|ne quaesumus tradas nos in perpetuum propter nomen tuum et ne dissipes testamentum tuum
DAN|3|35|neque auferas misericordiam tuam a nobis propter Abraham dilectum tuum et Isaac servum tuum et Israhel sanctum tuum
DAN|3|36|quibus locutus es pollicens quod multiplicares semen eorum sicut stellas caeli et sicut harenam quae est in litore maris
DAN|3|37|quia Domine inminuti sumus plus quam omnes gentes sumusque humiles in universa terra hodie propter peccata nostra
DAN|3|38|et non est in tempore hoc princeps et propheta et dux neque holocaustum neque sacrificium neque oblatio neque incensum neque locus primitiarum coram te
DAN|3|39|ut possimus invenire misericordiam sed in anima contrita et spiritu humilitatis suscipiamur
DAN|3|40|sicut in holocaustum arietum et taurorum et sicut in milibus agnorum pinguium sic fiat sacrificium nostrum in conspectu tuo hodie ut placeat tibi quoniam non est confusio confidentibus in te
DAN|3|41|et nunc sequimur in toto corde et timemus te et quaerimus faciem tuam
DAN|3|42|ne confundas nos sed fac nobiscum iuxta mansuetudinem tuam et secundum multitudinem misericordiae tuae
DAN|3|43|et erue nos in mirabilibus tuis et da gloriam nomini tuo Domine
DAN|3|44|et confundantur omnes qui ostendunt servis tuis mala confundantur in omni potentia et robur eorum conteratur
DAN|3|45|sciant quia tu Domine Deus solus et gloriosus super orbem terrarum
DAN|3|46|et non cessabant qui inmiserant eos ministri regis succendere fornacem naptha et stuppa et pice et malleolis
DAN|3|47|et effundebatur flamma super fornacem cubitis quadraginta novem
DAN|3|48|et erupit et incendit quos repperit iuxta fornacem de Chaldeis
DAN|3|49|angelus autem descendit cum Azaria et sociis eius in fornacem et excussit flammam ignis de fornace
DAN|3|50|et fecit medium fornacis quasi ventum roris flantem et non tetigit eos omnino ignis neque contristavit nec quicquam molestiae intulit
DAN|3|51|tunc hii tres quasi ex uno ore laudabant et glorificabant et benedicebant Deo in fornace dicentes
DAN|3|52|benedictus es Domine Deus patrum nostrorum et laudabilis et superexaltatus in saecula et benedictum nomen gloriae tuae sanctum et laudabile et superexaltatum in omnibus saeculis
DAN|3|53|benedictus es in templo sancto gloriae tuae et superlaudabilis et supergloriosus in saecula
DAN|3|54|benedictus es in throno regni tui et superlaudabilis et superexaltatus in saecula
DAN|3|55|benedictus es qui intueris abyssos et sedes super cherubin et laudabilis et superexaltatus in saecula
DAN|3|56|benedictus es in firmamento caeli et laudabilis et gloriosus in saecula
DAN|3|57|benedicite omnia opera Domini Domino laudate et superexaltate eum in saecula
DAN|3|58|benedicite angeli Domino laudate et superexaltate eum in saecula
DAN|3|59|benedicite caeli Domino laudate et superexaltate eum in saecula
DAN|3|60|benedicite aquae omnes quae super caelos sunt Domino laudate et superexaltate eum in saecula
DAN|3|61|benedicite omnes virtutes Domini Domino laudate et superexaltate eum in saecula
DAN|3|62|benedicite sol et luna Domino laudate et superexaltate eum in saecula
DAN|3|63|benedicite stellae caeli Domino laudate et superexaltate eum in saecula
DAN|3|64|benedicite omnis imber et ros Domino laudate et superexaltate eum in saecula
DAN|3|65|benedicite omnis spiritus Domino laudate et superexaltate eum in saecula
DAN|3|66|benedicite ignis et aestus Domino laudate et superexaltate eum in saecula
DAN|3|67|benedicite frigus et aestus Domino laudate et superexaltate eum in saecula
DAN|3|68|benedicite rores et pruina Domino laudate et superexaltate eum in saecula
DAN|3|69|benedicite gelu et frigus Domino laudate et superexaltate eum in saecula
DAN|3|70|benedicite glacies et nives Domino laudate et superexaltate eum in saecula
DAN|3|71|benedicite noctes et dies Domino laudate et superexaltate eum in saecula
DAN|3|72|benedicite lux et tenebrae Domino laudate et superexaltate eum in saecula
DAN|3|73|benedicite fulgura et nubes Domino laudate et superexaltate eum in saecula
DAN|3|74|benedicat terra Dominum laudet et superexaltet eum in saecula
DAN|3|75|benedicite montes et colles Domino laudate et superexaltate eum in saecula
DAN|3|76|benedicite universa germinantia in terra Domino laudate et superexaltate eum in saecula
DAN|3|77|benedicite fontes Domino laudate et superexaltate eum in saecula
DAN|3|78|benedicite maria et flumina Domino laudate et superexaltate eum in saecula
DAN|3|79|benedicite cete et omnia quae moventur in aquis Domino laudate et superexaltate eum in saecula
DAN|3|80|benedicite omnes volucres caeli Domino laudate et superexaltate eum in saecula
DAN|3|81|benedicite omnes bestiae et pecora Domino laudate et superexaltate eum in saecula
DAN|3|82|benedicite filii hominum Domino laudate et superexaltate eum in saecula
DAN|3|83|benedic Israhel Domino laudate et superexaltate eum in saecula
DAN|3|84|benedicite sacerdotes Domini Domino laudate et superexaltate eum in saecula
DAN|3|85|benedicite servi Domini Domino laudate et superexaltate eum in saecula
DAN|3|86|benedicite spiritus et animae iustorum Domino laudate et superexaltate eum in saecula
DAN|3|87|benedicite sancti et humiles corde Domino laudate et superexaltate eum in saecula
DAN|3|88|benedicite Anania Azaria et Misahel Domino laudate et superexaltate eum in saecula quia eruit nos de inferno et salvos fecit de manu mortis et liberavit de medio ardentis flammae et de medio ignis eruit nos
DAN|3|89|confitemini Domino quoniam bonus quoniam in saeculum misericordia eius
DAN|3|90|benedicite omnes religiosi Domino Deo deorum laudate et confitemini quia in omnia saecula misericordia eius
DAN|3|91|tunc Nabuchodonosor rex obstipuit et surrexit propere et ait optimatibus suis nonne tres viros misimus in medio ignis conpeditos qui respondentes dixerunt regi vere rex
DAN|3|92|respondit et ait ecce ego video viros quattuor solutos et ambulantes in medio ignis et nihil corruptionis in eis est et species quarti similis filio Dei
DAN|3|93|tunc accessit Nabuchodonosor ad ostium fornacis ignis ardentis et ait Sedrac Misac et Abdenago servi Dei excelsi egredimini et venite statimque egressi sunt Sedrac Misac et Abdenago de medio ignis
DAN|3|94|et congregati satrapae magistratus et iudices et potentes regis contemplabantur viros illos quoniam nihil potestatis habuisset ignis in corporibus eorum et capillus capitis eorum non esset adustus et sarabara eorum non fuissent inmutata et odor ignis non transisset per eos
DAN|3|95|et erumpens Nabuchodonosor ait benedictus Deus eorum Sedrac videlicet Misac et Abdenago qui misit angelum suum et eruit servos suos quia crediderunt in eo et verbum regis inmutaverunt et tradiderunt corpora sua ne servirent et ne adorarent omnem deum excepto Deo suo
DAN|3|96|a me ergo positum est hoc decretum ut omnis populus et tribus et lingua quaecumque locuta fuerit blasphemiam contra Deum Sedrac Misac et Abdenago dispereat et domus eius vastetur neque enim est Deus alius qui possit ita salvare
DAN|3|97|tunc rex promovit Sedrac Misac et Abdenago in provincia Babylonis
DAN|3|98|Nabuchodonosor rex omnibus populis gentibus et linguis quae habitant in universa terra pax vobis multiplicetur
DAN|3|99|signa et mirabilia fecit apud me Deus excelsus placuit ergo mihi praedicare
DAN|3|100|signa eius quia magna sunt et mirabilia eius quia fortia et regnum eius regnum sempiternum et potestas eius in generationem et generationem
DAN|4|1|ego Nabuchodonosor quietus eram in domo mea et florens in palatio meo
DAN|4|2|somnium vidi quod perterruit me et cogitationes meae in stratu meo et visiones capitis mei conturbaverunt me
DAN|4|3|et per me propositum est decretum ut introducerentur in conspectu meo cuncti sapientes Babylonis et ut solutionem somnii indicarent mihi
DAN|4|4|tunc ingrediebantur arioli magi Chaldei et aruspices et somnium narravi in conspectu eorum et solutionem eius non indicaverunt mihi
DAN|4|5|donec collega ingressus est in conspectu meo Danihel cuius nomen Balthasar secundum nomen dei mei qui habet spiritum deorum sanctorum in semet ipso et somnium coram eo locutus sum
DAN|4|6|Balthasar princeps ariolorum quem ego scio quod spiritum deorum sanctorum habeas in te et omne sacramentum non est inpossibile tibi visiones somniorum meorum quas vidi et solutionem eorum narra
DAN|4|7|visio capitis mei in cubili meo videbam et ecce arbor in medio terrae et altitudo eius nimia
DAN|4|8|magna arbor et fortis et proceritas eius contingens caelum aspectus illius erat usque ad terminos universae terrae
DAN|4|9|folia eius pulcherrima et fructus eius nimius et esca universorum in ea subter eam habitabant animalia et bestiae et in ramis eius conversabantur volucres caeli et ex ea vescebatur omnis caro
DAN|4|10|videbam in visione capitis mei super stratum meum et ecce vigil et sanctus de caelo descendit
DAN|4|11|clamavit fortiter et sic ait succidite arborem et praecidite ramos eius excutite folia eius et dispergite fructum eius fugiant bestiae quae subter eam sunt et volucres de ramis eius
DAN|4|12|verumtamen germen radicum eius in terra sinite et alligetur vinculo ferreo et aereo in herbis quae foris sunt et rore caeli tinguatur et cum feris pars eius in herba terrae
DAN|4|13|cor eius ab humano commutetur et cor ferae detur ei et septem tempora mutentur super eum
DAN|4|14|in sententia vigilum decretum est et sermo sanctorum et petitio donec cognoscant viventes quoniam dominatur Excelsus in regno hominum et cuicumque voluerit dabit illud et humillimum hominem constituet super eo
DAN|4|15|hoc somnium vidi ego rex Nabuchodonosor tu ergo Balthasar interpretationem narra festinus quia omnes sapientes regni mei non queunt solutionem edicere mihi tu autem potes quia spiritus deorum sanctorum in te est
DAN|4|16|tunc Danihel cuius nomen Balthasar coepit intra semet ipsum tacitus cogitare quasi hora una et cogitationes eius conturbabant eum respondens autem rex ait Balthasar somnium et interpretatio eius non conturbent te respondit Balthasar et dixit domine mi somnium his qui te oderunt et interpretatio eius hostibus tuis sit
DAN|4|17|arborem quam vidisti sublimem atque robustam cuius altitudo pertingit ad caelum et aspectus illius in omnem terram
DAN|4|18|et rami eius pulcherrimi et fructus eius nimius et esca omnium in ea subter eam habitantes bestiae agri et in ramis eius commorantes aves caeli
DAN|4|19|tu es rex qui magnificatus es et invaluisti et magnitudo tua crevit et pervenit usque ad caelum et potestas tua in terminos universae terrae
DAN|4|20|quod autem vidit rex vigilem et sanctum descendere de caelo et dicere succidite arborem et dissipate illam attamen germen radicum eius in terra dimittite et vinciatur ferro et aere in herbis foris et rore caeli conspergatur et cum feris sit pabulum eius donec septem tempora commutentur super eum
DAN|4|21|haec est interpretatio sententiae Altissimi quae pervenit super dominum meum regem
DAN|4|22|eicient te ab hominibus et cum bestiis feris erit habitatio tua et faenum ut bos comedes et rore caeli infunderis septem quoque tempora mutabuntur super te donec scias quod dominetur Excelsus super regnum hominum et cuicumque voluerit det illud
DAN|4|23|quod autem praecepit ut relinqueretur germen radicum eius id est arboris regnum tuum tibi manebit postquam cognoveris potestatem esse caelestem
DAN|4|24|quam ob rem rex consilium meum placeat tibi et peccata tua elemosynis redime et iniquitates tuas misericordiis pauperum forsitan ignoscat delictis tuis
DAN|4|25|omnia venerunt super Nabuchodonosor regem
DAN|4|26|post finem mensuum duodecim in aula Babylonis deambulabat
DAN|4|27|responditque rex et ait nonne haec est Babylon magna quam ego aedificavi in domum regni in robore fortitudinis meae et in gloria decoris mei
DAN|4|28|cum adhuc sermo esset in ore regis vox de caelo ruit tibi dicitur Nabuchodonosor rex regnum transiit a te
DAN|4|29|et ab hominibus te eicient et cum bestiis feris erit habitatio tua faenum quasi bos comedes et septem tempora mutabuntur super te donec scias quod dominetur Excelsus in regno hominum et cuicumque voluerit det illud
DAN|4|30|eadem hora sermo conpletus est super Nabuchodonosor ex hominibus abiectus est et faenum ut bos comedit et rore caeli corpus eius infectum est donec capilli eius in similitudinem aquilarum crescerent et ungues eius quasi avium
DAN|4|31|igitur post finem dierum ego Nabuchodonosor oculos meos ad caelum levavi et sensus meus redditus est mihi et Altissimo benedixi et viventem in sempiternum laudavi et glorificavi quia potestas eius potestas sempiterna et regnum eius in generationem et generationem
DAN|4|32|et omnes habitatores terrae apud eum in nihilum reputati sunt iuxta voluntatem enim suam facit tam in virtutibus caeli quam in habitatoribus terrae et non est qui resistat manui eius et dicat ei quare fecisti
DAN|4|33|in ipso tempore sensus meus reversus est ad me et ad honorem regni mei decoremque perveni et figura mea reversa est ad me et optimates mei et magistratus mei requisierunt me et in regno meo constitutus sum et magnificentia amplior addita est mihi
DAN|4|34|nunc igitur ego Nabuchodonosor laudo et magnifico et glorifico Regem caeli quia omnia opera eius vera et viae eius iudicia et gradientes in superbia potest humiliare
DAN|5|1|Balthasar rex fecit grande convivium optimatibus suis mille et unusquisque secundum suam bibebat aetatem
DAN|5|2|praecepit ergo iam temulentus ut adferrentur vasa aurea et argentea quae asportaverat Nabuchodonosor pater eius de templo quod fuit in Hierusalem ut biberent in eis rex et optimates eius uxoresque eius et concubinae
DAN|5|3|tunc adlata sunt vasa aurea quae asportaverat de templo quod fuerat in Hierusalem et biberunt in eis rex et optimates eius uxores et concubinae illius
DAN|5|4|bibebant vinum et laudabant deos suos aureos et argenteos et aereos ferreos ligneosque et lapideos
DAN|5|5|in eadem hora apparuerunt digiti quasi manus hominis scribentis contra candelabrum in superficie parietis aulae regiae et rex aspiciebat articulos manus scribentis
DAN|5|6|tunc regis facies commutata est et cogitationes eius conturbabant eum et conpages renum eius solvebantur et genua eius ad se invicem conlidebantur
DAN|5|7|exclamavit itaque rex fortiter ut introducerent magos Chaldeos et aruspices et proloquens rex ait sapientibus Babylonis quicumque legerit scripturam hanc et interpretationem eius manifestam mihi fecerit purpura vestietur et torquem auream habebit in collo et tertius in regno meo erit
DAN|5|8|tunc ingressi omnes sapientes regis non potuerunt nec scripturam legere nec interpretationem indicare regi
DAN|5|9|unde rex Balthasar satis conturbatus est et vultus illius inmutatus est sed et optimates eius turbabantur
DAN|5|10|regina autem pro re quae acciderat regi et optimatibus eius domum convivii ingressa est et proloquens ait rex in aeternum vive non te conturbent cogitationes tuae neque facies tua inmutetur
DAN|5|11|est vir in regno tuo qui spiritum deorum sanctorum habet in se et in diebus patris tui scientia et sapientia inventae sunt in eo nam et rex Nabuchodonosor pater tuus principem magorum incantatorum Chaldeorum et aruspicum constituit eum pater inquam tuus o rex
DAN|5|12|quia spiritus amplior et prudentia intellegentiaque interpretatio somniorum et ostensio secretorum ac solutio ligatorum inventae sunt in eo hoc est in Danihelo cui rex posuit nomen Balthasar nunc itaque Danihel vocetur et interpretationem narrabit
DAN|5|13|igitur introductus est Danihel coram rege ad quem praefatus rex ait tu es Danihel de filiis captivitatis Iudae quam adduxit rex pater meus de Iudaea
DAN|5|14|audivi de te quoniam spiritum deorum habeas et scientia intellegentiaque ac sapientia ampliores inventae sint in te
DAN|5|15|et nunc introgressi sunt in conspectu meo sapientes magi ut scripturam hanc legerent et interpretationem eius indicarent mihi et nequiverunt sensum sermonis huius edicere
DAN|5|16|porro ego audivi de te quod possis obscura interpretari et ligata dissolvere si ergo vales scripturam legere et interpretationem indicare mihi purpura vestieris et torquem auream circa collum tuum habebis et tertius in regno meo princeps eris
DAN|5|17|ad quae respondens Danihel ait coram rege munera tua sint tibi et dona domus tuae alteri da scripturam autem legam tibi rex et interpretationem eius ostendam tibi
DAN|5|18|o rex Deus altissimus regnum et magnificentiam gloriam et honorem dedit Nabuchodonosor patri tuo
DAN|5|19|et propter magnificentiam quam dederat ei universi populi tribus et linguae tremebant et metuebant eum quos volebat interficiebat et quos volebat percutiebat quos volebat exaltabat et quos volebat humiliabat
DAN|5|20|quando autem elevatum est cor eius et spiritus illius obfirmatus est ad superbiam depositus est de solio regni sui et gloria eius ablata est
DAN|5|21|et a filiis hominum eiectus est sed et cor eius cum bestiis positum est et cum onagris erat habitatio eius faenum quoque ut bos comedebat et rore caeli corpus eius infectum est donec cognosceret quod potestatem habeat Altissimus in regno hominum et quemcumque voluerit suscitabit super illud
DAN|5|22|tu quoque filius eius Balthasar non humiliasti cor tuum cum scires haec omnia
DAN|5|23|sed adversum Dominatorem caeli elevatus es et vasa domus eius adlata sunt coram te et tu et optimates tui et uxores tuae et concubinae vinum bibistis in eis deos quoque argenteos et aureos et aereos ferreos ligneosque et lapideos qui non vident neque audiunt neque sentiunt laudasti porro Deum qui habet flatum tuum in manu sua et omnes vias tuas non glorificasti
DAN|5|24|idcirco ab eo missus est articulus manus quae scripsit hoc quod exaratum est
DAN|5|25|haec est autem scriptura quae digesta est mane thecel fares
DAN|5|26|et haec interpretatio sermonis mane numeravit Deus regnum tuum et conplevit illud
DAN|5|27|thecel adpensum est in statera et inventus es minus habens
DAN|5|28|fares divisum est regnum tuum et datum est Medis et Persis
DAN|5|29|tunc iubente rege indutus est Danihel purpura et circumdata est torques aurea collo eius et praedicatum est de eo quod haberet potestatem tertius in regno
DAN|5|30|eadem nocte interfectus est Balthasar rex Chaldeus
DAN|5|31|et Darius Medus successit in regnum annos natus sexaginta duo
DAN|6|1|placuit Dario et constituit supra regnum satrapas centum viginti ut essent in toto regno suo
DAN|6|2|et super eos principes tres ex quibus Danihel unus erat ut satrapae illis redderent rationem et rex non sustineret molestiam
DAN|6|3|igitur Danihel superabat omnes principes et satrapas quia spiritus Dei amplior erat in eo
DAN|6|4|porro rex cogitabat constituere eum super omne regnum unde principes et satrapae quaerebant occasionem ut invenirent Daniheli ex latere regni nullamque causam et suspicionem repperire potuerunt eo quod fidelis esset et omnis culpa et suspicio non inveniretur in eo
DAN|6|5|dixerunt ergo viri illi non inveniemus Daniheli huic aliquam occasionem nisi forte in lege Dei sui
DAN|6|6|tunc principes et satrapae subripuerunt regi et sic locuti sunt ei Darie rex in aeternum vive
DAN|6|7|consilium inierunt cuncti principes regni magistratus et satrapae senatores et iudices ut decretum imperatorium exeat et edictum ut omnis qui petierit aliquam petitionem a quocumque deo et homine usque ad dies triginta nisi a te rex mittatur in lacum leonum
DAN|6|8|nunc itaque rex confirma sententiam et scribe decretum ut non inmutetur quod statutum est a Medis atque Persis nec praevaricari cuiquam liceat
DAN|6|9|porro rex Darius proposuit edictum et statuit
DAN|6|10|quod cum Danihel conperisset id est constitutam legem ingressus est domum suam et fenestris apertis in cenaculo suo contra Hierusalem tribus temporibus in die flectebat genua sua et adorabat confitebaturque coram Deo suo sicut et ante facere consueverat
DAN|6|11|viri igitur illi curiosius inquirentes invenerunt Danihel orantem et obsecrantem Deum suum
DAN|6|12|et accedentes locuti sunt regi super edicto rex numquid non constituisti ut omnis homo qui rogaret quemquam de diis et hominibus usque ad dies triginta nisi a te rex mitteretur in lacum leonum ad quod respondens rex ait verus sermo iuxta decretum Medorum atque Persarum quod praevaricari non licet
DAN|6|13|tunc respondentes dixerunt coram rege Danihel de filiis captivitatis Iudae non curavit de lege tua et de edicto quod constituisti sed tribus temporibus per diem orat obsecratione sua
DAN|6|14|quod verbum cum audisset rex satis contristatus est et pro Danihel posuit cor ut liberaret eum et usque ad occasum solis laborabat ut erueret illum
DAN|6|15|viri autem illi intellegentes regem dixerunt ei scito rex quia lex Medorum est atque Persarum ut omne decretum quod constituit rex non liceat inmutari
DAN|6|16|tunc rex praecepit et adduxerunt Danihelem et miserunt eum in lacum leonum dixitque rex Daniheli Deus tuus quem colis semper ipse liberabit te
DAN|6|17|adlatusque est lapis unus et positus est super os laci quem obsignavit rex anulo suo et anulo optimatum suorum ne quid fieret contra Danihel
DAN|6|18|et abiit rex in domum suam et dormivit incenatus cibique non sunt inlati coram eo insuper et somnus recessit ab eo
DAN|6|19|tunc rex primo diluculo consurgens festinus ad lacum leonum perrexit
DAN|6|20|adpropinquansque lacui Danihelem voce lacrimabili inclamavit et affatus est eum Danihel serve Dei viventis Deus tuus cui tu servis semper putasne valuit liberare te a leonibus
DAN|6|21|et Danihel regi respondens ait rex in aeternum vive
DAN|6|22|Deus meus misit angelum suum et conclusit ora leonum et non nocuerunt mihi quia coram eo iustitia inventa est in me sed et coram te rex delictum non feci
DAN|6|23|tunc rex vehementer gavisus est super eo et Danihelem praecepit educi de lacu eductusque est Danihel de lacu et nulla laesio inventa est in eo quia credidit Deo suo
DAN|6|24|iubente autem rege adducti sunt viri illi qui accusaverant Danihelem et in lacum leonum missi sunt ipsi et filii et uxores eorum et non pervenerunt usque ad pavimentum laci donec arriperent eos leones et omnia ossa eorum comminuerunt
DAN|6|25|tunc Darius rex scripsit universis populis tribubus et linguis habitantibus in universa terra pax vobis multiplicetur
DAN|6|26|a me constitutum est decretum ut in universo imperio et regno meo tremescant et paveant Deum Danihelis ipse est enim Deus vivens et aeternus in saecula et regnum eius non dissipabitur et potestas eius usque in aeternum
DAN|6|27|ipse liberator atque salvator faciens signa et mirabilia in caelo et in terra qui liberavit Danihelem de manu leonum
DAN|6|28|porro Danihel perseveravit usque ad regnum Darii regnumque Cyri Persae
DAN|7|1|anno primo Balthasar regis Babylonis Danihel somnium vidit visio autem capitis eius in cubili suo et somnium scribens brevi sermone conprehendit summatimque perstringens ait
DAN|7|2|videbam in visione mea nocte et ecce quattuor venti caeli pugnabant in mari magno
DAN|7|3|et quattuor bestiae grandes ascendebant de mari diversae inter se
DAN|7|4|prima quasi leaena et alas habebat aquilae aspiciebam donec evulsae sunt alae eius et sublata est de terra et super pedes quasi homo stetit et cor eius datum est ei
DAN|7|5|et ecce bestia alia similis urso in parte stetit et tres ordines erant in ore eius et in dentibus eius et sic dicebant ei surge comede carnes plurimas
DAN|7|6|post hoc aspiciebam et ecce alia quasi pardus et alas habebat avis quattuor super se et quattuor capita erant in bestia et potestas data est ei
DAN|7|7|post hoc aspiciebam in visione noctis et ecce bestia quarta terribilis atque mirabilis et fortis nimis dentes ferreos habebat magnos comedens atque comminuens et reliqua pedibus suis conculcans dissimilis autem erat ceteris bestiis quas videram ante eam et habebat cornua decem
DAN|7|8|considerabam cornua et ecce cornu aliud parvulum ortum est de medio eorum et tria de cornibus primis evulsa sunt a facie eius et ecce oculi quasi oculi hominis erant in cornu isto et os loquens ingentia
DAN|7|9|aspiciebam donec throni positi sunt et antiquus dierum sedit vestimentum eius quasi nix candidum et capilli capitis eius quasi lana munda thronus eius flammae ignis rotae eius ignis accensus
DAN|7|10|fluvius igneus rapidusque egrediebatur a facie eius milia milium ministrabant ei et decies milies centena milia adsistebant ei iudicium sedit et libri aperti sunt
DAN|7|11|aspiciebam propter vocem sermonum grandium quos cornu illud loquebatur et vidi quoniam interfecta esset bestia et perisset corpus eius et traditum esset ad conburendum igni
DAN|7|12|aliarum quoque bestiarum ablata esset potestas et tempora vitae constituta essent eis usque ad tempus et tempus
DAN|7|13|aspiciebam ergo in visione noctis et ecce cum nubibus caeli quasi filius hominis veniebat et usque ad antiquum dierum pervenit et in conspectu eius obtulerunt eum
DAN|7|14|et dedit ei potestatem et honorem et regnum et omnes populi tribus ac linguae ipsi servient potestas eius potestas aeterna quae non auferetur et regnum eius quod non corrumpetur
DAN|7|15|horruit spiritus meus ego Danihel territus sum in his et visiones capitis mei conturbaverunt me
DAN|7|16|accessi ad unum de adsistentibus et veritatem quaerebam ab eo de omnibus his qui dixit mihi interpretationem sermonum et edocuit me
DAN|7|17|hae bestiae magnae quattuor quattuor regna consurgent de terra
DAN|7|18|suscipient autem regnum sancti Dei altissimi et obtinebunt regnum usque in saeculum et saeculum saeculorum
DAN|7|19|post hoc volui diligenter discere de bestia quarta quia erat dissimilis valde ab omnibus et terribilis nimis dentes et ungues eius ferrei comedebat et comminuebat et reliquias pedibus suis conculcabat
DAN|7|20|et de cornibus decem quae habebat in capite et de alio quod ortum fuerat ante quod ceciderant tria cornua de cornu illo quod habebat oculos et os loquens grandia et maius erat ceteris
DAN|7|21|aspiciebam et ecce cornu illud faciebat bellum adversus sanctos et praevalebat eis
DAN|7|22|donec venit antiquus dierum et iudicium dedit sanctis Excelsi et tempus advenit et regnum obtinuerunt sancti
DAN|7|23|et sic ait bestia quarta regnum quartum erit in terra quod maius erit omnibus regnis et devorabit universam terram et conculcabit et comminuet eam
DAN|7|24|porro cornua decem ipsius regni decem reges erunt et alius consurget post eos et ipse potentior erit prioribus et tres reges humiliabit
DAN|7|25|et sermones contra Excelsum loquetur et sanctos Altissimi conteret et putabit quod possit mutare tempora et leges et tradentur in manu eius usque ad tempus et tempora et dimidium temporis
DAN|7|26|et iudicium sedebit ut auferatur potentia et conteratur et dispereat usque in finem
DAN|7|27|regnum autem et potestas et magnitudo regni quae est subter omne caelum detur populo sanctorum Altissimi cuius regnum regnum sempiternum est et omnes reges servient ei et oboedient
DAN|7|28|hucusque finis verbi ego Danihel multum cogitationibus meis conturbabar et facies mea mutata est in me verbum autem in corde meo conservavi
DAN|8|1|anno tertio regni Balthasar regis visio apparuit mihi ego Danihel post id quod videram in principio
DAN|8|2|vidi in visione mea cum essem in Susis castro quod est in Aelam civitate vidi autem in visione esse me super portam Ulai
DAN|8|3|et levavi oculos meos et vidi et ecce aries unus stabat ante paludem habens cornua excelsa et unum excelsius altero atque succrescens postea
DAN|8|4|vidi arietem cornibus ventilantem contra occidentem et contra aquilonem et contra meridiem et omnes bestiae non poterant resistere ei neque liberari de manu eius fecitque secundum voluntatem suam et magnificatus est
DAN|8|5|et ego intellegebam ecce autem hircus caprarum veniebat ab occidente super faciem totius terrae et non tangebat terram porro hircus habebat cornu insigne inter oculos suos
DAN|8|6|et venit usque ad arietem illum cornutum quem videram stantem ante portam et cucurrit ad eum in impetu fortitudinis suae
DAN|8|7|cumque adpropinquasset prope arietem efferatus est in eum et percussit arietem et comminuit duo cornua eius et non poterat aries resistere ei cumque eum misisset in terram conculcavit et nemo quibat liberare arietem de manu eius
DAN|8|8|hircus autem caprarum magnus factus est nimis cumque crevisset fractum est cornu magnum et orta sunt cornua quattuor subter illud per quattuor ventos caeli
DAN|8|9|de uno autem ex eis egressum est cornu unum modicum et factum est grande contra meridiem et contra orientem et contra fortitudinem
DAN|8|10|et magnificatum est usque ad fortitudinem caeli et deiecit de fortitudine et de stellis et conculcavit eas
DAN|8|11|et usque ad principem fortitudinis magnificatus est et ab eo tulit iuge sacrificium et deiecit locum sanctificationis eius
DAN|8|12|robur autem datum est contra iuge sacrificium propter peccata et prosternetur veritas in terra et faciet et prosperabitur
DAN|8|13|et audivi unum de sanctis loquentem et dixit unus sanctus alteri nescio cui loquenti usquequo visio et iuge sacrificium et peccatum desolationis quae facta est et sanctuarium et fortitudo conculcabitur
DAN|8|14|et dixit ei usque ad vesperam et mane duo milia trecenti et mundabitur sanctuarium
DAN|8|15|factum est autem cum viderem ego Danihel visionem et quaererem intellegentiam ecce stetit in conspectu meo quasi species viri
DAN|8|16|et audivi vocem viri inter Ulai et clamavit et ait Gabrihel fac intellegere istum visionem
DAN|8|17|et venit et stetit iuxta ubi ego stabam cumque venisset pavens corrui in faciem meam et ait ad me intellege fili hominis quoniam in tempore finis conplebitur visio
DAN|8|18|cumque loqueretur ad me conlapsus sum pronus in terram et tetigit me et statuit me in gradu meo
DAN|8|19|dixitque mihi ego ostendam tibi quae futura sint in novissimo maledictionis quoniam habet tempus finem suum
DAN|8|20|aries quem vidisti habere cornua rex Medorum est atque Persarum
DAN|8|21|porro hircus caprarum rex Graecorum est et cornu grande quod erat inter oculos eius ipse est rex primus
DAN|8|22|quod autem fracto illo surrexerunt quattuor pro eo quattuor reges de gente eius consurgent sed non in fortitudine eius
DAN|8|23|et post regnum eorum cum creverint iniquitates consurget rex inpudens facie et intellegens propositiones
DAN|8|24|et roborabitur fortitudo eius sed non in viribus suis et supra quam credi potest universa vastabit et prosperabitur et faciet et interficiet robustos et populum sanctorum
DAN|8|25|secundum voluntatem suam et dirigetur dolus in manu eius et cor suum magnificabit et in copia rerum omnium occidet plurimos et contra principem principum consurget et sine manu conteretur
DAN|8|26|et visio vespere et mane quae dicta est vera est tu ergo signa visionem quia post dies multos erit
DAN|8|27|et ego Danihel langui et aegrotavi per dies cumque surrexissem faciebam opera regis et stupebam ad visionem et non erat qui interpretaretur
DAN|9|1|in anno primo Darii filii Asueri de semine Medorum qui imperavit super regnum Chaldeorum
DAN|9|2|anno uno regni eius ego Danihel intellexi in libris numerum annorum de quo factus est sermo Domini ad Hieremiam prophetam ut conplerentur desolationes Hierusalem septuaginta anni
DAN|9|3|et posui faciem meam ad Dominum Deum rogare et deprecari in ieiuniis sacco et cinere
DAN|9|4|et oravi Dominum Deum meum et confessus sum et dixi obsecro Domine Deus magne et terribilis custodiens pactum et misericordiam diligentibus te et custodientibus mandata tua
DAN|9|5|peccavimus inique fecimus impie egimus et recessimus et declinavimus a mandatis tuis ac iudiciis
DAN|9|6|non oboedivimus servis tuis prophetis qui locuti sunt in nomine tuo regibus nostris principibus nostris patribus nostris omnique populo terrae
DAN|9|7|tibi Domine iustitia nobis autem confusio faciei sicut est hodie viro Iuda et habitatoribus Hierusalem et omni Israhel his qui prope sunt et his qui procul in universis terris ad quas eiecisti eos propter iniquitates eorum in quibus peccaverunt in te
DAN|9|8|Domine nobis confusio faciei regibus nostris principibus nostris et patribus nostris qui peccaverunt
DAN|9|9|tibi autem Domino Deo nostro misericordia et propitiatio quia recessimus a te
DAN|9|10|et non audivimus vocem Domini Dei nostri ut ambularemus in lege eius quam posuit nobis per servos suos prophetas
DAN|9|11|et omnis Israhel praevaricati sunt legem tuam et declinaverunt ne audirent vocem tuam et stillavit super nos maledictio et detestatio quae scripta est in libro Mosi servi Dei quia peccavimus ei
DAN|9|12|et statuit sermones suos quos locutus est super nos et super principes nostros qui iudicaverunt nos ut superducerent in nos malum magnum quale numquam fuit sub omni caelo secundum quod factum est in Hierusalem
DAN|9|13|sicut scriptum est in lege Mosi omne malum hoc venit super nos et non rogavimus faciem tuam Domine Deus noster ut reverteremur ab iniquitatibus nostris et cogitaremus veritatem tuam
DAN|9|14|et vigilavit Dominus et adduxit eam super nos iustus Dominus Deus noster in omnibus operibus suis quae fecit non enim audivimus vocem eius
DAN|9|15|et nunc Domine Deus noster qui eduxisti populum tuum de terra Aegypti in manu forti et fecisti tibi nomen secundum diem hanc peccavimus iniquitatem fecimus
DAN|9|16|Domine in omnem iustitiam tuam avertatur obsecro ira tua et furor tuus a civitate tua Hierusalem et monte sancto tuo propter peccata enim nostra et iniquitates patrum nostrorum Hierusalem et populus tuus in obprobrium sunt omnibus per circuitum nostrum
DAN|9|17|nunc ergo exaudi Deus noster orationem servi tui et preces eius et ostende faciem tuam super sanctuarium tuum quod desertum est propter temet ipsum
DAN|9|18|inclina Deus meus aurem tuam et audi aperi oculos tuos et vide desolationem nostram et civitatem super quam invocatum est nomen tuum neque enim in iustificationibus nostris prosternimus preces ante faciem tuam sed in miserationibus tuis multis
DAN|9|19|exaudi Domine placare Domine adtende et fac ne moreris propter temet ipsum Deus meus quia nomen tuum invocatum est super civitatem et super populum tuum
DAN|9|20|cumque adhuc loquerer et orarem et confiterer peccata mea et peccata populi mei Israhel ut prosternerem preces meas in conspectu Dei mei pro monte sancto Dei mei
DAN|9|21|adhuc me loquente in oratione ecce vir Gabrihel quem videram in visione principio cito volans tetigit me in tempore sacrificii vespertini
DAN|9|22|et docuit me et locutus est mihi dixitque Danihel nunc egressus sum ut docerem te et intellegeres
DAN|9|23|ab exordio precum tuarum egressus est sermo ego autem veni ut indicarem tibi quia vir desideriorum es tu ergo animadverte sermonem et intellege visionem
DAN|9|24|septuaginta ebdomades adbreviatae sunt super populum tuum et super urbem sanctam tuam ut consummetur praevaricatio et finem accipiat peccatum et deleatur iniquitas et adducatur iustitia sempiterna et impleatur visio et prophetes et unguatur sanctus sanctorum
DAN|9|25|scito ergo et animadverte ab exitu sermonis ut iterum aedificetur Hierusalem usque ad christum ducem ebdomades septem et ebdomades sexaginta duae erunt et rursum aedificabitur platea et muri in angustia temporum
DAN|9|26|et post ebdomades sexaginta duas occidetur christus et non erit eius et civitatem et sanctuarium dissipabit populus cum duce venturo et finis eius vastitas et post finem belli statuta desolatio
DAN|9|27|confirmabit autem pactum multis ebdomas una et in dimidio ebdomadis deficiet hostia et sacrificium et in templo erit abominatio desolationis et usque ad consummationem et finem perseverabit desolatio
DAN|10|1|anno tertio Cyri regis Persarum verbum revelatum est Daniheli cognomento Balthasar et verum verbum et fortitudo magna intellexitque sermonem intellegentia est enim opus in visione
DAN|10|2|in diebus illis ego Danihel lugebam trium ebdomadarum diebus
DAN|10|3|panem desiderabilem non comedi et caro et vinum non introierunt in os meum sed neque unguento unctus sum donec conplerentur trium ebdomadarum dies
DAN|10|4|die autem vicesima et quarta mensis primi eram iuxta fluvium magnum qui est Tigris
DAN|10|5|et levavi oculos meos et vidi et ecce vir unus vestitus lineis et renes eius accincti auro obrizo
DAN|10|6|et corpus eius quasi chrysolitus et facies eius velut species fulgoris et oculi eius ut lampas ardens et brachia eius et quae deorsum usque ad pedes quasi species aeris candentis et vox sermonum eius ut vox multitudinis
DAN|10|7|vidi autem ego Danihel solus visionem porro viri qui erant mecum non viderunt sed terror nimius inruit super eos et fugerunt in absconditum
DAN|10|8|ego autem relictus solus vidi visionem grandem hanc et non remansit in me fortitudo sed et species mea inmutata est in me et emarcui nec habui quicquam virium
DAN|10|9|et audivi vocem sermonum eius et audiens iacebam consternatus super faciem meam vultusque meus herebat terrae
DAN|10|10|et ecce manus tetigit me et erexit me super genua mea et super articulos manuum mearum
DAN|10|11|et dixit ad me Danihel vir desideriorum intellege verba quae ego loquor ad te et sta in gradu tuo nunc enim sum missus ad te cumque dixisset mihi sermonem istum steti tremens
DAN|10|12|et ait ad me noli metuere Danihel quia ex die primo quo posuisti cor tuum ad intellegendum ut te adfligeres in conspectu Dei tui exaudita sunt verba tua et ego veni propter sermones tuos
DAN|10|13|princeps autem regni Persarum restitit mihi viginti et uno diebus et ecce Michahel unus de principibus primis venit in adiutorium meum et ego remansi ibi iuxta regem Persarum
DAN|10|14|veni autem ut docerem te quae ventura sunt populo tuo in novissimis diebus quoniam adhuc visio in dies
DAN|10|15|cumque loqueretur mihi huiuscemodi verbis deieci vultum meum ad terram et tacui
DAN|10|16|et ecce quasi similitudo filii hominis tetigit labia mea et aperiens os meum locutus sum et dixi ad eum qui stabat contra me domine mi in visione tua dissolutae sunt conpages meae et nihil in me remansit virium
DAN|10|17|et quomodo poterit servus domini mei loqui cum domino meo nihil enim in me remansit virium sed et halitus meus intercluditur
DAN|10|18|rursum ergo tetigit me quasi visio hominis et confortavit me
DAN|10|19|et dixit noli timere vir desideriorum pax tibi confortare et esto robustus cumque loqueretur mecum convalui et dixi loquere domine mi quia confortasti me
DAN|10|20|et ait numquid scis quare venerim ad te et nunc revertar ut proelier adversum principem Persarum cum enim egrederer apparuit princeps Graecorum veniens
DAN|10|21|verumtamen adnuntiabo tibi quod expressum est in scriptura veritatis et nemo est adiutor meus in omnibus his nisi Michahel princeps vester
DAN|11|1|ego autem ab anno primo Darii Medi stabam ut confortaretur et roboraretur
DAN|11|2|et nunc veritatem adnuntiabo tibi ecce adhuc tres reges stabunt in Perside et quartus ditabitur opibus nimiis super omnes et cum invaluerit divitiis suis concitabit omnes adversum regnum Graeciae
DAN|11|3|surget vero rex fortis et dominabitur potestate multa et faciet quod placuerit ei
DAN|11|4|et cum steterit conteretur regnum eius et dividetur in quattuor ventos caeli sed non in posteros eius neque secundum potentiam illius qua dominatus est lacerabitur enim regnum eius etiam in externos exceptis his
DAN|11|5|et confortabitur rex austri et de principibus eius praevalebit super eum et dominabitur dicione multa enim dominatio eius
DAN|11|6|et post finem annorum foederabuntur filiaque regis austri veniet ad regem aquilonis facere amicitiam et non obtinebit fortitudinem brachii nec stabit semen eius et tradetur ipsa et qui adduxerunt eam adulescentes eius et qui confortabant eam in temporibus
DAN|11|7|et stabit de germine radicum eius plantatio et veniet cum exercitu et ingredietur provinciam regis aquilonis et abutetur eis et obtinebit
DAN|11|8|insuper et deos eorum et sculptilia vasa quoque pretiosa argenti et auri captiva ducet in Aegyptum ipse praevalebit adversum regem aquilonis
DAN|11|9|et intrabit in regnum rex austri et revertetur ad terram suam
DAN|11|10|filii autem eius provocabuntur et congregabunt multitudinem exercituum plurimorum et veniet properans et inundans et revertetur et concitabitur et congredietur cum robore eius
DAN|11|11|et provocatus rex austri egredietur et pugnabit adversum regem aquilonis et praeparabit multitudinem nimiam et dabitur multitudo in manu eius
DAN|11|12|et capiet multitudinem et exaltabitur cor eius et deiciet multa milia sed non praevalebit
DAN|11|13|convertetur enim rex aquilonis et praeparabit multitudinem multo maiorem quam prius et in fine temporum annorumque veniet properans cum exercitu magno et opibus nimiis
DAN|11|14|et in temporibus illis multi consurgent adversum regem austri filii quoque praevaricatorum populi tui extollentur ut impleant visionem et corruent
DAN|11|15|et veniet rex aquilonis et conportabit aggerem et capiet urbes munitissimas et brachia austri non sustinebunt et consurgent electi eius ad resistendum et non erit fortitudo
DAN|11|16|et faciet veniens super eum iuxta placitum suum et non erit qui stet contra faciem eius et stabit in terra inclita et consumetur in manu eius
DAN|11|17|et ponet faciem suam ut veniat ad tenendum universum regnum eius et recta faciet cum eo et filiam feminarum dabit ei ut evertat illud et non stabit nec illius erit
DAN|11|18|et convertet faciem suam ad insulas et capiet multas et cessare faciet principem obprobrii sui et obprobrium eius convertetur in eum
DAN|11|19|et convertet faciem suam ad imperium terrae suae et inpinget et corruet et non invenietur
DAN|11|20|et stabit in loco eius vilissimus et indignus decore regio et in paucis diebus conteretur non in furore nec in proelio
DAN|11|21|et stabit in loco eius despectus et non tribuetur ei honor regius et veniet clam et obtinebit regnum in fraudulentia
DAN|11|22|et brachia pugnantis expugnabuntur a facie eius et conterentur insuper et dux foederis
DAN|11|23|et post amicitias cum eo faciet dolum et ascendet et superabit in modico populo
DAN|11|24|abundantes et uberes urbes ingredietur et faciet quae non fecerunt patres eius et patres patrum eius rapinas et praedam et divitias eorum dissipabit et contra firmissimas cogitationes iniet et hoc usque ad tempus
DAN|11|25|et concitabitur fortitudo eius et cor eius adversum regem austri in exercitu magno et rex austri provocabitur ad bellum multis auxiliis et fortibus nimis et non stabunt quia inibunt adversum eum consilia
DAN|11|26|et comedentes panem cum eo conterent illum exercitusque eius opprimetur et cadent interfecti plurimi
DAN|11|27|duorum quoque regum cor erit ut malefaciant et ad mensam unam mendacium loquentur et non proficient quia adhuc finis in aliud tempus
DAN|11|28|et revertetur in terram suam cum opibus multis et cor eius adversus testamentum sanctum et faciet et revertetur in terram suam
DAN|11|29|statuto tempore revertetur et veniet ad austrum et non erit priori simile novissimum
DAN|11|30|et venient super eum trieres et Romani et percutietur et revertetur et indignabitur contra testamentum sanctuarii et faciet reverteturque et cogitabit adversum eos qui dereliquerunt testamentum sanctuarii
DAN|11|31|et brachia ex eo stabunt et polluent sanctuarium fortitudinis et auferent iuge sacrificium et dabunt abominationem in desolationem
DAN|11|32|et impii in testamentum simulabunt fraudulenter populus autem sciens Deum suum obtinebit et faciet
DAN|11|33|et docti in populo docebunt plurimos et ruent in gladio et in flamma in captivitate et rapina dierum
DAN|11|34|cumque corruerint sublevabuntur auxilio parvulo et adplicabuntur eis plurimi fraudulenter
DAN|11|35|et de eruditis ruent ut conflentur et eligantur et dealbentur usque ad tempus praefinitum quia adhuc aliud tempus erit
DAN|11|36|et faciet iuxta voluntatem suam rex et elevabitur et magnificabitur adversum omnem deum et adversum Deum deorum loquetur magnifica et diriget donec conpleatur iracundia perpetrata est quippe definitio
DAN|11|37|et Deum patrum suorum non reputabit et erit in concupiscentiis feminarum nec quemquam deorum curabit quia adversum universa consurget
DAN|11|38|deum autem Maozim in loco suo venerabitur et deum quem ignoraverunt patres eius colet auro et argento et lapide pretioso rebusque pretiosis
DAN|11|39|et faciet ut muniat Maozim cum deo alieno quem cognovit et multiplicabit gloriam et dabit eis potestatem in multis et terram dividet gratuito
DAN|11|40|et in tempore praefinito proeliabitur adversum eum rex austri et quasi tempestas veniet contra illum rex aquilonis in curribus et in equitibus et in classe magna et ingredietur terras et conteret et pertransiet
DAN|11|41|et introibit in terram gloriosam et multae corruent hae autem solae salvabuntur de manu eius Edom et Moab et principium filiorum Ammon
DAN|11|42|et mittet manum suam in terras et terra Aegypti non effugiet
DAN|11|43|et dominabitur thesaurorum auri et argenti et in omnibus pretiosis Aegypti per Lybias quoque et Aethiopias transibit
DAN|11|44|et fama turbabit eum ab oriente et ab aquilone et veniet in multitudine magna ut conterat et interficiat plurimos
DAN|11|45|et figet tabernaculum suum Apedno inter maria super montem inclitum et sanctum et veniet usque ad summitatem eius et nemo auxiliabitur ei
DAN|12|1|in tempore autem illo consurget Michahel princeps magnus qui stat pro filiis populi tui et veniet tempus quale non fuit ab eo quo gentes esse coeperunt usque ad tempus illud et in tempore illo salvabitur populus tuus omnis qui inventus fuerit scriptus in libro
DAN|12|2|et multi de his qui dormiunt in terrae pulvere evigilabunt alii in vitam aeternam et alii in obprobrium ut videant semper
DAN|12|3|qui autem docti fuerint fulgebunt quasi splendor firmamenti et qui ad iustitiam erudiunt multos quasi stellae in perpetuas aeternitates
DAN|12|4|tu autem Danihel clude sermones et signa librum usque ad tempus statutum pertransibunt plurimi et multiplex erit scientia
DAN|12|5|et vidi ego Danihel et ecce quasi duo alii stabant unus hinc super ripam fluminis et alius inde ex altera ripa fluminis
DAN|12|6|et dixi viro qui indutus erat lineis qui stabat super aquas fluminis usquequo finis horum mirabilium
DAN|12|7|et audivi virum qui indutus erat lineis qui stabat super aquas fluminis cum levasset dexteram et sinistram suam in caelum et iurasset per viventem in aeternum quia in tempus temporum et dimidium temporis et cum conpleta fuerit dispersio manus populi sancti conplebuntur universa haec
DAN|12|8|et ego audivi et non intellexi et dixi domine mi quid erit post haec
DAN|12|9|et ait vade Danihel quia clausi sunt signatique sermones usque ad tempus praefinitum
DAN|12|10|eligentur et dealbabuntur et quasi ignis probabuntur multi et impie agent impii neque intellegent omnes impii porro docti intellegent
DAN|12|11|et a tempore cum ablatum fuerit iuge sacrificium et posita fuerit abominatio in desolatione dies mille ducenti nonaginta
DAN|12|12|beatus qui expectat et pervenit ad dies mille trecentos triginta quinque
DAN|12|13|tu autem vade ad praefinitum et requiesce et stabis in sorte tua in fine dierum
HOS|1|1|verbum Domini quod factum est ad Osee filium Beeri in diebus Oziae Ioatham Ahaz Ezechiae regum Iuda et in diebus Hieroboam filii Ioas regis Israhel
HOS|1|2|principium loquendi Dominum in Osee et dixit Dominus ad Osee vade sume tibi uxorem fornicationum et filios fornicationum quia fornicans fornicabitur terra a Domino
HOS|1|3|et abiit et accepit Gomer filiam Debelaim et concepit et peperit filium
HOS|1|4|et dixit Dominus ad eum voca nomen eius Hiezrahel quoniam adhuc modicum et visitabo sanguinem Hiezrahel super domum Hieu et quiescere faciam regnum domus Israhel
HOS|1|5|et in illa die conteram arcum Israhel in valle Hiezrahel
HOS|1|6|et concepit adhuc et peperit filiam et dixit ei voca nomen eius Absque misericordia quia non addam ultra misereri domui Israhel sed oblivione obliviscar eorum
HOS|1|7|et domui Iuda miserebor et salvabo eos in Domino Deo suo et non salvabo eos in arcu et gladio et in bello et in equis et in equitibus
HOS|1|8|et ablactavit eam quae erat absque misericordia et concepit et peperit filium
HOS|1|9|et dixit voca nomen eius Non populus meus quia vos non populus meus et ego non ero vester
HOS|1|10|et erit numerus filiorum Israhel quasi harena maris quae sine mensura est et non numerabitur et erit in loco ubi dicetur eis non populus meus vos dicetur eis filii Dei viventis
HOS|1|11|et congregabuntur filii Iuda et filii Israhel pariter et ponent sibimet caput unum et ascendent de terra quia magnus dies Hiezrahel
HOS|2|1|dicite fratribus vestris Populus meus et sorori vestrae Misericordiam consecuta
HOS|2|2|iudicate matrem vestram iudicate quoniam ipsa non uxor mea et ego non vir eius auferat fornicationes suas a facie sua et adulteria sua de medio uberum suorum
HOS|2|3|ne forte expoliem eam nudam et statuam eam secundum diem nativitatis suae et ponam eam quasi solitudinem et statuam eam velut terram inviam et interficiam eam siti
HOS|2|4|et filiorum illius non miserebor quoniam filii fornicationum sunt
HOS|2|5|quia fornicata est mater eorum confusa est quae concepit eos quia dixit vadam post amatores meos qui dant panes mihi et aquas meas lanam meam et linum meum oleum meum et potum meum
HOS|2|6|propter hoc ecce ego sepiam viam tuam spinis et sepiam eam maceria et semitas suas non inveniet
HOS|2|7|et sequetur amatores suos et non adprehendet eos et quaeret eos et non inveniet et dicet vadam et revertar ad virum meum priorem quia bene mihi erat tunc magis quam nunc
HOS|2|8|et haec nescivit quia ego dedi ei frumentum et vinum et oleum et argentum multiplicavi ei et aurum quae fecerunt Baal
HOS|2|9|idcirco convertar et sumam frumentum meum in tempore suo et vinum meum in tempore suo et liberabo lanam meam et linum meum quae operiebant ignominiam eius
HOS|2|10|et nunc revelabo stultitiam eius in oculis amatorum eius et vir non eruet eam de manu mea
HOS|2|11|et cessare faciam omne gaudium eius sollemnitatem eius neomeniam eius sabbatum eius et omnia festa tempora eius
HOS|2|12|et corrumpam vineam eius et ficum eius de quibus dixit mercedes hae meae sunt quas dederunt mihi amatores mei et ponam eam in saltu et comedet illam bestia agri
HOS|2|13|et visitabo super eam dies Baalim quibus accendebat incensum et ornabatur inaure sua et monili suo et ibat post amatores suos et mei obliviscebatur dicit Dominus
HOS|2|14|propter hoc ecce ego lactabo eam et ducam eam in solitudinem et loquar ad cor eius
HOS|2|15|et dabo ei vinitores eius ex eodem loco et vallem Achor ad aperiendam spem et canet ibi iuxta dies iuventutis suae et iuxta dies ascensionis suae de terra Aegypti
HOS|2|16|et erit in die illo ait Dominus vocabit me Vir meus et non vocabit me ultra Baali
HOS|2|17|et auferam nomina Baalim de ore eius et non recordabitur ultra nominis eorum
HOS|2|18|et percutiam eis foedus in die illa cum bestia agri et cum volucre caeli et cum reptili terrae et arcum et gladium et bellum conteram de terra et dormire eos faciam fiducialiter
HOS|2|19|et sponsabo te mihi in sempiternum et sponsabo te mihi in iustitia et iudicio et in misericordia et miserationibus
HOS|2|20|et sponsabo te mihi in fide et scies quia ego Dominus
HOS|2|21|et erit in illa die exaudiam dicit Dominus exaudiam caelos et illi exaudient terram
HOS|2|22|et terra exaudiet triticum et vinum et oleum et haec exaudient Hiezrahel
HOS|2|23|et seminabo eam mihi in terram et miserebor eius quae fuit absque misericordia
HOS|2|24|et dicam non populo meo populus meus tu et ipse dicet Dominus meus es tu
HOS|3|1|et dixit Dominus ad me adhuc vade dilige mulierem dilectam amico et adulteram sicut diligit Dominus filios Israhel et ipsi respectant ad deos alienos et diligunt vinacea uvarum
HOS|3|2|et fodi eam mihi quindecim argenteis et choro hordei et dimidio choro hordei
HOS|3|3|et dixi ad eam dies multos expectabis me non fornicaberis et non eris viro sed et ego expectabo te
HOS|3|4|quia dies multos sedebunt filii Israhel sine rege et sine principe et sine sacrificio et sine altari et sine ephod et sine therafin
HOS|3|5|et post haec revertentur filii Israhel et quaerent Dominum Deum suum et David regem suum et pavebunt ad Dominum et ad bonum eius in novissimo dierum
HOS|4|1|audite verbum Domini filii Israhel quia iudicium Domino cum habitatoribus terrae non est enim veritas et non est misericordia et non est scientia Dei in terra
HOS|4|2|maledictum et mendacium et homicidium et furtum et adulterium inundaverunt et sanguis sanguinem tetigit
HOS|4|3|propter hoc lugebit terra et infirmabitur omnis qui habitat in ea in bestia agri et in volucre caeli sed et pisces maris congregabuntur
HOS|4|4|verumtamen unusquisque non iudicet et non arguatur vir populus enim tuus sicut hii qui contradicunt sacerdoti
HOS|4|5|et corrues hodie et corruet etiam propheta tecum nocte tacere feci matrem tuam
HOS|4|6|conticuit populus meus eo quod non habuerit scientiam quia tu scientiam reppulisti repellam te ne sacerdotio fungaris mihi et oblita es legis Dei tui obliviscar filiorum tuorum et ego
HOS|4|7|secundum multitudinem eorum sic peccaverunt mihi gloriam eorum in ignominiam commutabo
HOS|4|8|peccata populi mei comedent et ad iniquitatem eorum sublevabunt animas eorum
HOS|4|9|et erit sicut populus sic sacerdos et visitabo super eum vias eius et cogitationes eius reddam ei
HOS|4|10|et comedent et non saturabuntur fornicati sunt et non cessaverunt quoniam Dominum reliquerunt in non custodiendo
HOS|4|11|fornicatio et vinum et ebrietas aufert cor
HOS|4|12|populus meus in ligno suo interrogavit et baculus eius adnuntiavit ei spiritus enim fornicationum decepit eos et fornicati sunt a Deo suo
HOS|4|13|super capita montium sacrificabant et super colles accendebant thymiama subtus quercum et populum et terebinthum quia bona erat umbra eius ideo fornicabuntur filiae vestrae et sponsae vestrae adulterae erunt
HOS|4|14|non visitabo super filias vestras cum fuerint fornicatae et super sponsas vestras cum adulteraverint quoniam ipsi cum meretricibus versabantur et cum effeminatis sacrificabant et populus non intellegens vapulabit
HOS|4|15|si fornicaris tu Israhel non delinquat saltim Iuda et nolite ingredi in Galgala et ne ascenderitis in Bethaven neque iuraveritis vivit Dominus
HOS|4|16|quoniam sicut vacca lasciviens declinavit Israhel nunc pascet eos Dominus quasi agnum in latitudine
HOS|4|17|particeps idolorum Ephraim dimitte eum
HOS|4|18|separatum est convivium eorum fornicatione fornicati sunt dilexerunt adferre ignominiam protectores eius
HOS|4|19|ligavit spiritus eam in alis suis et confundentur a sacrificiis suis
HOS|5|1|audite hoc sacerdotes et adtendite domus Israhel et domus regis auscultate quia vobis iudicium est quoniam laqueus facti estis speculationi et rete expansum super Thabor
HOS|5|2|et victimas declinastis in profundum et ego eruditor omnium eorum
HOS|5|3|ego scio Ephraim et Israhel non est absconditus a me quia nunc fornicatus est Ephraim contaminatus est Israhel
HOS|5|4|non dabunt cogitationes suas ut revertantur ad Dominum suum quia spiritus fornicationis in medio eorum et Dominum non cognoverunt
HOS|5|5|et respondebit arrogantia Israhel in facie eius et Israhel et Ephraim ruent in iniquitate sua ruet etiam Iudas cum eis
HOS|5|6|in gregibus suis et in armentis suis vadent ad quaerendum Dominum et non invenient ablatus est ab eis
HOS|5|7|in Domino praevaricati sunt quia filios alienos genuerunt nunc devorabit eos mensis cum partibus suis
HOS|5|8|clangite bucina in Gabaa tuba in Rama ululate in Bethaven post tergum tuum Beniamin
HOS|5|9|Ephraim in desolatione erit in die correptionis in tribubus Israhel ostendi fidem
HOS|5|10|facti sunt principes Iuda quasi adsumentes terminum super eos effundam quasi aquam iram meam
HOS|5|11|calumniam patiens Ephraim fractus iudicio quoniam coepit abire post sordem
HOS|5|12|et ego quasi tinea Ephraim et quasi putredo domui Iuda
HOS|5|13|et vidit Ephraim languorem suum et Iudas vinculum suum et abiit Ephraim ad Assur et misit ad regem ultorem et ipse non poterit sanare vos nec solvere poterit a vobis vinculum
HOS|5|14|quoniam ego quasi leaena Ephraim et quasi catulus leonis domui Iuda ego ego capiam et vadam tollam et non est qui eruat
HOS|5|15|vadens revertar ad locum meum donec deficiatis et quaeratis faciem meam
HOS|6|1|in tribulatione sua mane consurgunt ad me venite et revertamur ad Dominum
HOS|6|2|quia ipse cepit et sanabit nos percutiet et curabit nos
HOS|6|3|vivificabit nos post duos dies in die tertia suscitabit nos et vivemus in conspectu eius sciemus sequemurque ut cognoscamus Dominum quasi diluculum praeparatus est egressus eius et veniet quasi imber nobis temporaneus et serotinus terrae
HOS|6|4|quid faciam tibi Ephraim quid faciam tibi Iuda misericordia vestra quasi nubes matutina et quasi ros mane pertransiens
HOS|6|5|propter hoc dolavi in prophetis occidi eos in verbis oris mei et iudicia tua quasi lux egredientur
HOS|6|6|quia misericordiam volui et non sacrificium et scientiam Dei plus quam holocausta
HOS|6|7|ipsi autem sicut Adam transgressi sunt pactum ibi praevaricati sunt in me
HOS|6|8|Galaad civitas operantium idolum subplantata sanguine
HOS|6|9|et quasi fauces virorum latronum particeps sacerdotum in via interficientium pergentes de Sychem quia scelus operati sunt
HOS|6|10|in domo Israhel vidi horrendum ibi fornicationes Ephraim contaminatus est Israhel
HOS|6|11|sed et Iuda pone messem tibi cum convertero captivitatem populi mei
HOS|7|1|cum sanare vellem Israhel revelata est iniquitas Ephraim et malitia Samariae quia operati sunt mendacium et fur ingressus est spolians latrunculus foris
HOS|7|2|et ne forte dicant in cordibus suis omnem malitiam eorum me recordatum nunc circumdederunt eos adinventiones suae coram facie mea factae sunt
HOS|7|3|in malitia sua laetificaverunt regem et in mendaciis suis principes
HOS|7|4|omnes adulterantes quasi clibanus succensus a coquente quievit paululum civitas a commixtione fermenti donec fermentaretur totum
HOS|7|5|dies regis nostri coeperunt principes furere a vino extendit manum suam cum inlusoribus
HOS|7|6|quia adplicuerunt quasi clibanum cor suum cum insidiaretur eis tota nocte dormivit coquens eos mane ipse succensus quasi ignis flammae
HOS|7|7|omnes calefacti sunt quasi clibanus et devoraverunt iudices suos omnes reges eorum ceciderunt non est qui clamet in eis ad me
HOS|7|8|Ephraim in populis ipse commiscebatur Ephraim factus est subcinericius qui non reversatur
HOS|7|9|comederunt alieni robur eius et ipse nescivit sed et cani effusi sunt in eo et ipse ignoravit
HOS|7|10|et humiliabitur superbia Israhel in facie eius nec reversi sunt ad Dominum Deum suum et non quaesierunt eum in omnibus his
HOS|7|11|et factus est Ephraim quasi columba seducta non habens cor Aegyptum invocabant ad Assyrios abierunt
HOS|7|12|et cum profecti fuerint expandam super eos rete meum quasi volucrem caeli detraham eos caedam eos secundum auditionem coetus eorum
HOS|7|13|vae eis quoniam recesserunt a me vastabuntur quia praevaricati sunt in me et ego redemi eos et ipsi locuti sunt contra me mendacia
HOS|7|14|et non clamaverunt ad me in corde suo sed ululabant in cubilibus suis super triticum et vinum ruminabant recesserunt a me
HOS|7|15|et ego erudivi et confortavi brachia eorum et in me cogitaverunt malitiam
HOS|7|16|reversi sunt ut essent absque iugo facti sunt quasi arcus dolosus cadent in gladio principes eorum a furore linguae suae ista subsannatio eorum in terra Aegypti
HOS|8|1|in gutture tuo sit tuba quasi aquila super domum Domini pro eo quod transgressi sunt foedus meum et legem meam praevaricati sunt
HOS|8|2|me invocabunt Deus meus cognovimus te Israhel
HOS|8|3|proiecit Israhel bonum inimicus persequetur eum
HOS|8|4|ipsi regnaverunt et non ex me principes extiterunt et non cognovi argentum suum et aurum suum fecerunt sibi idola ut interirent
HOS|8|5|proiectus est vitulus tuus Samaria iratus est furor meus in eis usquequo non poterunt emundari
HOS|8|6|quia ex Israhel et ipse est artifex fecit illum et non est Deus quoniam in aranearum telas erit vitulus Samariae
HOS|8|7|quia ventum seminabunt et turbinem metent culmus stans non est in eis germen non faciet farinam quod si et fecerit alieni comedent eam
HOS|8|8|devoratus est Israhel nunc factus est in nationibus quasi vas inmundum
HOS|8|9|quia ipsi ascenderunt ad Assur onager solitarius sibi Ephraim munera dederunt amatoribus
HOS|8|10|sed et cum mercede conduxerint nationes nunc congregabo eos et quiescent paulisper ab onere regis et principum
HOS|8|11|quia multiplicavit Ephraim altaria ad peccandum factae sunt ei arae in delictum
HOS|8|12|scribam ei multiplices leges meas quae velut alienae conputatae sunt
HOS|8|13|hostias adfer adfer immolabunt carnes et comedent Dominus non suscipiet eas nunc recordabitur iniquitatis eorum et visitabit peccata eorum ipsi in Aegyptum convertentur
HOS|8|14|et oblitus est Israhel factoris sui et aedificavit delubra et Iudas multiplicavit urbes munitas et mittam ignem in civitates eius et devorabit aedes illius
HOS|9|1|noli laetari Israhel noli exultare sicut populi quia fornicatus es a Deo tuo dilexisti mercedem super omnes areas tritici
HOS|9|2|area et torcular non pascet eos et vinum mentietur eis
HOS|9|3|non habitabunt in terra Domini reversus est Ephraim Aegyptum et in Assyriis pollutum comedit
HOS|9|4|non libabunt Domino vinum et non placebunt ei sacrificia eorum quasi panis lugentium omnes qui comedunt eum contaminabuntur quia panis eorum animae ipsorum non intrabit in domum Domini
HOS|9|5|quid facietis in die sollemni in die festivitatis Domini
HOS|9|6|ecce enim profecti sunt a vastitate Aegyptus congregavit eos Memphis sepeliet eos desiderabile argenti eorum urtica hereditabit lappa in tabernaculis eorum
HOS|9|7|venerunt dies visitationis venerunt dies retributionis scitote Israhel stultum prophetam insanum virum spiritalem propter multitudinem iniquitatis tuae et multitudo amentiae
HOS|9|8|speculator Ephraim cum Deo meo propheta laqueus ruinae super omnes vias eius insania in domo Dei eius
HOS|9|9|profunde peccaverunt sicut in diebus Gabaa recordabitur iniquitatis eorum et visitabit peccata eorum
HOS|9|10|quasi uvas in deserto inveni Israhel quasi prima poma ficulneae in cacumine eius vidi patres eorum ipsi autem intraverunt ad Beelphegor et abalienati sunt in confusione et facti sunt abominabiles sicut ea quae dilexerunt
HOS|9|11|Ephraim quasi avis avolavit gloria eorum a partu et ab utero et a conceptu
HOS|9|12|quod si et enutrierint filios suos absque liberis eos faciam in hominibus sed et vae eis cum recessero ab eis
HOS|9|13|Ephraim ut vidi Tyrus erat fundata in pulchritudine et Ephraim educit ad interfectorem filios suos
HOS|9|14|da eis Domine quid dabis eis da eis vulvam sine liberis et ubera arentia
HOS|9|15|omnes nequitiae eorum in Galgal quia ibi exosos habui eos propter malitiam adinventionum eorum de domo mea eiciam eos non addam ut diligam eos omnes principes eorum recedentes
HOS|9|16|percussus est Ephraim radix eorum exsiccata est fructum nequaquam facient quod si et genuerint interficiam amantissima uteri eorum
HOS|9|17|abiciet eos Deus meus quia non audierunt eum et erunt vagi in nationibus
HOS|10|1|vitis frondosa Israhel fructus adaequatus est ei secundum multitudinem fructus sui multiplicavit altaria iuxta ubertatem terrae suae exuberavit simulacris
HOS|10|2|divisum est cor eorum nunc interibunt ipse confringet simulacra eorum depopulabitur aras eorum
HOS|10|3|quia nunc dicent non est rex nobis non enim timemus Dominum et rex quid faciet nobis
HOS|10|4|loquimini verba visionis inutilis et ferietis foedus et germinabit quasi amaritudo iudicium super sulcos agri
HOS|10|5|vaccas Bethaven coluerunt habitatores Samariae quia luxit super eum populus eius et aeditui eius super eum exultaverunt in gloria eius quia migravit ab eo
HOS|10|6|siquidem et ipse in Assur delatus est munus regi ultori confusio Ephraim capiet et confundetur Israhel in voluntate sua
HOS|10|7|transire fecit Samaria regem suum quasi spumam super faciem aquae
HOS|10|8|et disperdentur excelsa idoli peccatum Israhel lappa et tribulus ascendet super aras eorum et dicent montibus operite nos et collibus cadite super nos
HOS|10|9|ex diebus Gabaa peccavit Israhel ibi steterunt non conprehendet eos in Gabaa proelium super filios iniquitatis
HOS|10|10|iuxta desiderium meum corripiam eos congregabuntur super eos populi cum corripientur propter duas iniquitates suas
HOS|10|11|Ephraim vitula docta diligere trituram et ego transivi super pulchritudinem colli eius ascendam super Ephraim arabit Iudas confringet sibi sulcos Iacob
HOS|10|12|seminate vobis in iustitia metite in ore misericordiae innovate vobis novale tempus autem requirendi Dominum cum venerit qui docebit vos iustitiam
HOS|10|13|arastis impietatem iniquitatem messuistis comedistis frugem mendacii quia confisus es in viis tuis in multitudine fortium tuorum
HOS|10|14|consurget tumultus in populo tuo et omnes munitiones tuae vastabuntur sicut vastatus est Salman a domo eius qui iudicavit Baal in die proelii matre super filios adlisa
HOS|10|15|sic fecit vobis Bethel a facie malitiae nequitiarum vestrarum
HOS|11|1|sicuti mane transit pertransiit rex Israhel quia puer Israhel et dilexi eum et ex Aegypto vocavi filium meum
HOS|11|2|vocaverunt eos sic abierunt a facie eorum Baalim immolabant et simulacris sacrificabant
HOS|11|3|et ego quasi nutricius Ephraim portabam eos in brachiis meis et nescierunt quod curarem eos
HOS|11|4|in funiculis Adam traham eos in vinculis caritatis et ero eis quasi exaltans iugum super maxillas eorum et declinavi ad eum ut vesceretur
HOS|11|5|non revertetur in terram Aegypti et Assur ipse rex eius quoniam noluerunt converti
HOS|11|6|coepit gladius in civitatibus eius et consumet electos eius et comedet capita eorum
HOS|11|7|et populus meus pendebit ad reditum meum iugum autem inponetur ei simul quod non auferetur
HOS|11|8|quomodo dabo te Ephraim protegam te Israhel quomodo dabo te sicut Adama ponam te ut Seboim conversum est in me cor meum pariter conturbata est paenitudo mea
HOS|11|9|non faciam furorem irae meae non convertar ut disperdam Ephraim quoniam Deus ego et non homo in medio tui Sanctus et non ingrediar civitatem
HOS|11|10|post Dominum ambulabunt quasi leo rugiet quia ipse rugiet et formidabunt filii maris
HOS|11|11|et avolabunt quasi avis ex Aegypto et quasi columba de terra Assyriorum et conlocabo eos in domibus suis dicit Dominus
HOS|11|12|circumdedit me in negatione Ephraim et in dolo domus Israhel Iudas autem testis descendit cum Deo et cum sanctis fidelis
HOS|12|1|Ephraim pascit ventum et sequitur aestum tota die mendacium et vastitatem multiplicat et foedus cum Assyriis iniit et oleum in Aegyptum ferebat
HOS|12|2|iudicium ergo Domini cum Iuda et visitatio super Iacob iuxta vias eius et iuxta adinventiones eius reddet ei
HOS|12|3|in utero subplantavit fratrem suum et in fortitudine sua directus est cum angelo
HOS|12|4|et invaluit ad angelum et confortatus est flevit et rogavit eum in Bethel invenit eum et ibi locutus est nobiscum
HOS|12|5|et Dominus Deus exercituum Dominus memoriale eius
HOS|12|6|et tu ad Deum tuum converteris misericordiam et iudicium custodi et spera in Deo tuo semper
HOS|12|7|Chanaan in manu eius statera dolosa calumniam dilexit
HOS|12|8|et dixit Ephraim verumtamen dives effectus sum inveni idolum mihi omnes labores mei non invenient mihi iniquitatem quam peccavi
HOS|12|9|et ego Dominus Deus tuus ex terra Aegypti adhuc sedere te faciam in tabernaculis sicut in diebus festivitatis
HOS|12|10|et locutus sum super prophetas et ego visionem multiplicavi et in manu prophetarum adsimilatus sum
HOS|12|11|si Galaad idolum tamen frustra erant in Galgal bubus immolantes nam et altaria eorum quasi acervi super sulcos agri
HOS|12|12|fugit Iacob in regionem Syriae et servivit Israhel in uxore et in uxore servavit
HOS|12|13|in propheta autem eduxit Dominus Israhel de Aegypto et in propheta servatus est
HOS|12|14|ad iracundiam me provocavit Ephraim in amaritudinibus suis et sanguis eius super eum veniet et obprobrium eius restituet ei Dominus suus
HOS|13|1|loquente Ephraim horror invasit Israhel et deliquit in Baal et mortuus est
HOS|13|2|et nunc addiderunt ad peccandum feceruntque sibi conflatile de argento suo quasi similitudinem idolorum factura artificum totum est his ipsi dicunt immolate homines vitulos adorantes
HOS|13|3|idcirco erunt quasi nubes matutina et sicut ros matutinus praeteriens sicut pulvis turbine raptus ex area et sicut fumus de fumario
HOS|13|4|ego autem Dominus Deus tuus ex terra Aegypti et Deum absque me nescies et salvator non est praeter me
HOS|13|5|ego cognovi te in deserto in terra solitudinis
HOS|13|6|iuxta pascua sua et adimpleti sunt et saturati elevaverunt cor suum et obliti sunt mei
HOS|13|7|et ero eis quasi leaena sicut pardus in via Assyriorum
HOS|13|8|occurram eis quasi ursa raptis catulis et disrumpam interiora iecoris eorum et consumam eos ibi quasi leo bestia agri scindet eos
HOS|13|9|perditio tua Israhel tantummodo in me auxilium tuum
HOS|13|10|ubi est rex tuus maxime nunc salvet te in omnibus urbibus tuis et iudices tui de quibus dixisti da mihi regem et principes
HOS|13|11|dabo tibi regem in furore meo et auferam in indignatione mea
HOS|13|12|conligata est iniquitas Ephraim absconditum peccatum eius
HOS|13|13|dolores parturientis venient ei ipse filius non sapiens nunc enim non stabit in contritione filiorum
HOS|13|14|de manu mortis liberabo eos de morte redimam eos ero mors tua o mors ero morsus tuus inferne consolatio abscondita est ab oculis meis
HOS|13|15|quia ipse inter fratres dividet adducet urentem ventum Dominus de deserto ascendentem et siccabit venas eius et desolabit fontem eius et ipse diripiet thesaurum omnis vasis desiderabilis
HOS|14|1|pereat Samaria quoniam ad amaritudinem concitavit Dominum suum in gladio pereat parvuli eorum elidantur et fetae eius discindantur
HOS|14|2|convertere Israhel ad Dominum Deum tuum quoniam corruisti in iniquitate tua
HOS|14|3|tollite vobiscum verba et convertimini ad Dominum dicite ei omnem aufer iniquitatem et accipe bonum et reddemus vitulos labiorum nostrorum
HOS|14|4|Assur non salvabit nos super equum non ascendemus nec dicemus ultra dii nostri opera manuum nostrarum quia eius qui in te est misereberis pupilli
HOS|14|5|sanabo contritiones eorum diligam eos spontanee quia aversus est furor meus ab eo
HOS|14|6|ero quasi ros Israhel germinabit quasi lilium et erumpet radix eius ut Libani
HOS|14|7|ibunt rami eius et erit quasi oliva gloria eius et odor eius ut Libani
HOS|14|8|convertentur sedentes in umbra eius vivent tritico et germinabunt quasi vinea memoriale eius sicut vinum Libani
HOS|14|9|Ephraim quid mihi ultra idola ego exaudiam et dirigam eum ego ut abietem virentem ex me fructus tuus inventus est
HOS|14|10|quis sapiens et intelleget ista intellegens et sciet haec quia rectae viae Domini et iusti ambulabunt in eis praevaricatores vero corruent in eis
JOEL|1|1|verbum Domini quod factum est ad Iohel filium Fatuhel
JOEL|1|2|audite hoc senes et auribus percipite omnes habitatores terrae si factum est istud in diebus vestris aut in diebus patrum vestrorum
JOEL|1|3|super hoc filiis vestris narrate et filii vestri filiis suis et filii eorum generationi alterae
JOEL|1|4|residuum erucae comedit lucusta et residuum lucustae comedit bruchus et residuum bruchi comedit rubigo
JOEL|1|5|expergescimini ebrii et flete et ululate omnes qui bibitis vinum in dulcedine quoniam periit ab ore vestro
JOEL|1|6|gens enim ascendit super terram meam fortis et innumerabilis dentes eius ut dentes leonis et molares eius ut catuli leonis
JOEL|1|7|posuit vineam meam in desertum et ficum meam decorticavit nudans spoliavit eam et proiecit albi facti sunt rami eius
JOEL|1|8|plange quasi virgo accincta sacco super virum pubertatis suae
JOEL|1|9|periit sacrificium et libatio de domo Domini luxerunt sacerdotes ministri Domini
JOEL|1|10|depopulata est regio luxit humus quoniam devastatum est triticum confusum est vinum elanguit oleum
JOEL|1|11|confusi sunt agricolae ululaverunt vinitores super frumento et hordeo quia periit messis agri
JOEL|1|12|vinea confusa est et ficus elanguit malogranatum et palma et malum et omnia ligna agri aruerunt quia confusum est gaudium a filiis hominum
JOEL|1|13|accingite vos et plangite sacerdotes ululate ministri altaris ingredimini cubate in sacco ministri Dei mei quoniam interiit de domo Dei vestri sacrificium et libatio
JOEL|1|14|sanctificate ieiunium vocate coetum congregate senes omnes habitatores terrae in domum Dei vestri et clamate ad Dominum
JOEL|1|15|a a a diei quia prope est dies Domini et quasi vastitas a potente veniet
JOEL|1|16|numquid non coram oculis vestris alimenta perierunt de domo Dei nostri laetitia et exultatio
JOEL|1|17|conputruerunt iumenta in stercore suo demolita sunt horrea dissipatae sunt apothecae quoniam confusum est triticum
JOEL|1|18|quid ingemuit animal mugierunt greges armenti quia non est pascua eis sed et greges pecorum disperierunt
JOEL|1|19|ad te Domine clamabo quia ignis comedit speciosa deserti et flamma succendit omnia ligna regionis
JOEL|1|20|sed et bestiae agri quasi area sitiens imbrem suspexerunt ad te quoniam exsiccati sunt fontes aquarum et ignis devoravit speciosa deserti
JOEL|2|1|canite tuba in Sion ululate in monte sancto meo conturbentur omnes habitatores terrae quia venit dies Domini quia prope est
JOEL|2|2|dies tenebrarum et caliginis dies nubis et turbinis quasi mane expansum super montes populus multus et fortis similis ei non fuit a principio et post eum non erit usque in annos generationis et generationis
JOEL|2|3|ante faciem eius ignis vorans et post eum exurens flamma quasi hortus voluptatis terra coram eo et post eum solitudo deserti neque est qui effugiat eum
JOEL|2|4|quasi aspectus equorum aspectus eorum et quasi equites sic current
JOEL|2|5|sicut sonitus quadrigarum super capita montium exilient sicut sonitus flammae ignis devorantis stipulam velut populus fortis praeparatus ad proelium
JOEL|2|6|a facie eius cruciabuntur populi omnes vultus redigentur in ollam
JOEL|2|7|sicut fortes current quasi viri bellatores ascendent murum vir in viis suis gradietur et non declinabunt a semitis suis
JOEL|2|8|unusquisque fratrem suum non coartabit singuli in calle suo ambulabunt sed et per fenestras cadent et non demolientur
JOEL|2|9|urbem ingredientur in muro current domos conscendent per fenestras intrabunt quasi fur
JOEL|2|10|a facie eius contremuit terra moti sunt caeli sol et luna obtenebrati sunt et stellae retraxerunt splendorem suum
JOEL|2|11|et Dominus dedit vocem suam ante faciem exercitus sui quia multa sunt nimis castra eius quia fortia et facientia verbum eius magnus enim dies Domini et terribilis valde et quis sustinebit eum
JOEL|2|12|nunc ergo dicit Dominus convertimini ad me in toto corde vestro in ieiunio et in fletu et in planctu
JOEL|2|13|et scindite corda vestra et non vestimenta vestra et convertimini ad Dominum Deum vestrum quia benignus et misericors est patiens et multae misericordiae et praestabilis super malitia
JOEL|2|14|quis scit si convertatur et ignoscat et relinquat post se benedictionem sacrificium et libamen Domino Deo nostro
JOEL|2|15|canite tuba in Sion sanctificate ieiunium vocate coetum
JOEL|2|16|congregate populum sanctificate ecclesiam coadunate senes congregate parvulos et sugentes ubera egrediatur sponsus de cubili suo et sponsa de thalamo suo
JOEL|2|17|inter vestibulum et altare plorabunt sacerdotes ministri Domini et dicent parce Domine populo tuo et ne des hereditatem tuam in obprobrium ut dominentur eis nationes quare dicunt in populis ubi est Deus eorum
JOEL|2|18|zelatus est Dominus terram suam et pepercit populo suo
JOEL|2|19|et respondit Dominus et dixit populo suo ecce ego mittam vobis frumentum et vinum et oleum et replebimini eo et non dabo vos ultra obprobrium in gentibus
JOEL|2|20|et eum qui ab aquilone est procul faciam a vobis et expellam eum in terram inviam et desertam faciem eius contra mare orientale et extremum eius ad mare novissimum et ascendet fetor eius et ascendet putredo eius quia superbe egit
JOEL|2|21|noli timere terra exulta et laetare quoniam magnificavit Dominus ut faceret
JOEL|2|22|nolite timere animalia regionis quia germinaverunt speciosa deserti quia lignum adtulit fructum suum ficus et vinea dederunt virtutem suam
JOEL|2|23|et filii Sion exultate et laetamini in Domino Deo vestro quia dedit vobis doctorem iustitiae et descendere faciet ad vos imbrem matutinum et serotinum in principio
JOEL|2|24|et implebuntur areae frumento et redundabunt torcularia vino et oleo
JOEL|2|25|et reddam vobis annos quos comedit lucusta bruchus et rubigo et eruca fortitudo mea magna quam misi in vos
JOEL|2|26|et comedetis vescentes et saturabimini et laudabitis nomen Domini Dei vestri qui fecit vobiscum mirabilia et non confundetur populus meus in sempiternum
JOEL|2|27|et scietis quia in medio Israhel ego sum et ego Dominus Deus vester et non est amplius et non confundetur populus meus in aeternum
JOEL|2|28|et erit post haec effundam spiritum meum super omnem carnem et prophetabunt filii vestri et filiae vestrae senes vestri somnia somniabunt et iuvenes vestri visiones videbunt
JOEL|2|29|sed et super servos et ancillas in diebus illis effundam spiritum meum
JOEL|2|30|et dabo prodigia in caelo et in terra sanguinem et ignem et vaporem fumi
JOEL|2|31|sol vertetur in tenebras et luna in sanguinem antequam veniat dies Domini magnus et horribilis
JOEL|2|32|et erit omnis qui invocaverit nomen Domini salvus erit quia in monte Sion et in Hierusalem erit salvatio sicut dixit Dominus et in residuis quos Dominus vocaverit
JOEL|3|1|quia ecce in diebus illis et in tempore illo cum convertero captivitatem Iuda et Hierusalem
JOEL|3|2|congregabo omnes gentes et deducam eas in valle Iosaphat et disceptabo cum eis ibi super populo meo et hereditate mea Israhel quos disperserunt in nationibus et terram meam diviserunt
JOEL|3|3|et super populum meum miserunt sortem et posuerunt puerum in prostibulum et puellam vendiderunt pro vino ut biberent
JOEL|3|4|verum quid vobis et mihi Tyrus et Sidon et omnis terminus Palestinorum numquid ultionem vos redditis mihi et si ulciscimini vos contra me cito velociter reddam vicissitudinem vobis super caput vestrum
JOEL|3|5|argentum enim meum et aurum tulistis et desiderabilia mea et pulcherrima intulistis in delubra vestra
JOEL|3|6|et filios Iuda et filios Hierusalem vendidistis filiis Graecorum ut longe faceretis eos de finibus suis
JOEL|3|7|ecce ego suscitabo eos de loco in quo vendidistis eos et convertam retributionem vestram in caput vestrum
JOEL|3|8|et vendam filios vestros et filias vestras in manibus filiorum Iuda et venundabunt eos Sabeis genti longinquae quia Dominus locutus est
JOEL|3|9|clamate hoc in gentibus sanctificate bellum suscitate robustos accedant ascendant omnes viri bellatores
JOEL|3|10|concidite aratra vestra in gladios et ligones vestros in lanceas infirmus dicat quia fortis ego sum
JOEL|3|11|erumpite et venite omnes gentes de circuitu et congregamini ibi occumbere faciet Dominus robustos tuos
JOEL|3|12|consurgant et ascendant gentes in vallem Iosaphat quia ibi sedebo ut iudicem omnes gentes in circuitu
JOEL|3|13|mittite falces quoniam maturavit messis venite et descendite quia plenum est torcular exuberant torcularia quia multiplicata est malitia eorum
JOEL|3|14|populi populi in valle concisionis quia iuxta est dies Domini in valle concisionis
JOEL|3|15|sol et luna obtenebricata sunt et stellae retraxerunt splendorem suum
JOEL|3|16|et Dominus de Sion rugiet et de Hierusalem dabit vocem suam et movebuntur caeli et terra et Dominus spes populi sui et fortitudo filiorum Israhel
JOEL|3|17|et scietis quia ego Dominus Deus vester habitans in Sion in monte sancto meo et erit Hierusalem sancta et alieni non transibunt per eam amplius
JOEL|3|18|et erit in die illa stillabunt montes dulcedinem et colles fluent lacte et per omnes rivos Iuda ibunt aquae et fons de domo Domini egredietur et inrigabit torrentem Spinarum
JOEL|3|19|Aegyptus in desolatione erit et Idumea in desertum perditionis pro eo quod inique egerint in filios Iuda et effuderint sanguinem innocentem in terra sua
JOEL|3|20|et Iudaea in aeternum habitabitur et Hierusalem in generatione et generationem
JOEL|3|21|et mundabo sanguinem eorum quem non mundaveram et Dominus commorabitur in Sion
AMOS|1|1|verba Amos qui fuit in pastoralibus de Thecuae quae vidit super Israhel in diebus Oziae regis Iuda et in diebus Hieroboam filii Ioas regis Israhel ante duos annos terraemotus
AMOS|1|2|et dixit Dominus de Sion rugiet et de Hierusalem dabit vocem suam et luxerunt speciosa pastorum et exsiccatus est vertex Carmeli
AMOS|1|3|haec dicit Dominus super tribus sceleribus Damasci et super quattuor non convertam eum eo quod trituraverint in plaustris ferreis Galaad
AMOS|1|4|et mittam ignem in domum Azahel et devorabit domos Benadad
AMOS|1|5|et conteram vectem Damasci et disperdam habitatorem de campo Idoli et tenentem sceptrum de domo Voluptatis et transferetur populus Syriae Cyrenen dicit Dominus
AMOS|1|6|haec dicit Dominus super tribus sceleribus Gazae et super quattuor non convertam eum eo quod transtulerit captivitatem perfectam ut concluderet eam in Idumea
AMOS|1|7|et mittam ignem in murum Gazae et devorabit aedes eius
AMOS|1|8|et disperdam habitatorem de Azoto et tenentem sceptrum de Ascalone et convertam manum meam super Accaron et peribunt reliqui Philisthinorum dicit Dominus Deus
AMOS|1|9|haec dicit Dominus super tribus sceleribus Tyri et super quattuor non convertam eum eo quod concluserint captivitatem perfectam in Idumea et non sint recordati foederis fratrum
AMOS|1|10|et emittam ignem in murum Tyri et devorabit aedes eius
AMOS|1|11|haec dicit Dominus super tribus sceleribus Edom et super quattuor non convertam eum eo quod persecutus sit in gladio fratrem suum et violaverit misericordiam eius et tenuerit ultra furorem suum et indignationem suam servaverit usque in finem
AMOS|1|12|mittam ignem in Theman et devorabit aedes Bosrae
AMOS|1|13|haec dicit Dominus super tribus sceleribus filiorum Ammon et super quattuor non convertam eum eo quod dissecuerit praegnantes Galaad ad dilatandum terminum suum
AMOS|1|14|et succendam ignem in muro Rabbae et devorabit aedes eius in ululatu in die belli et in turbine in die commotionis
AMOS|1|15|et ibit Melchom in captivitatem ipse et principes eius simul dicit Dominus
AMOS|2|1|haec dicit Dominus super tribus sceleribus Moab et super quattuor non convertam eum eo quod incenderit ossa regis Idumeae usque ad cinerem
AMOS|2|2|et mittam ignem in Moab et devorabit aedes Carioth et morietur in sonitu Moab in clangore tubae
AMOS|2|3|et disperdam iudicem de medio eius et omnes principes eius interficiam cum eo dicit Dominus
AMOS|2|4|haec dicit Dominus super tribus sceleribus Iuda et super quattuor non convertam eum eo quod abiecerint legem Domini et mandata eius non custodierint deceperunt enim eos idola sua post quae abierant patres eorum
AMOS|2|5|et mittam ignem in Iuda et devorabit aedes Hierusalem
AMOS|2|6|haec dicit Dominus super tribus sceleribus Israhel et super quattuor non convertam eum pro eo quod vendiderit argento iustum et pauperem pro calciamentis
AMOS|2|7|qui conterunt super pulverem terrae capita pauperum et viam humilium declinant et filius ac pater eius ierunt ad puellam ut violarent nomen sanctum meum
AMOS|2|8|et super vestimentis pigneratis accubuerunt iuxta omne altare et vinum damnatorum bibebant in domo Dei sui
AMOS|2|9|ego autem exterminavi Amorreum a facie eorum cuius altitudo cedrorum altitudo eius et fortis ipse quasi quercus et contrivi fructum eius desuper et radices eius subter
AMOS|2|10|ego sum qui ascendere vos feci de terra Aegypti et eduxi vos in deserto quadraginta annis ut possideretis terram Amorrei
AMOS|2|11|et suscitavi de filiis vestris in prophetas et de iuvenibus vestris nazarenos numquid non ita est filii Israhel dicit Dominus
AMOS|2|12|et propinabatis nazarenis vino et prophetis mandabatis dicentes ne prophetetis
AMOS|2|13|ecce ego stridebo super vos sicut stridet plaustrum onustum faeno
AMOS|2|14|et peribit fuga a veloce et fortis non obtinebit virtutem suam et robustus non salvabit animam suam
AMOS|2|15|et tenens arcum non stabit et velox pedibus suis non salvabitur et ascensor equi non salvabit animam suam
AMOS|2|16|et robustus corde inter fortes nudus fugiet in die illa dicit Dominus
AMOS|3|1|audite verbum quod locutus est Dominus super vos filii Israhel super omni cognatione quam eduxi de terra Aegypti dicens
AMOS|3|2|tantummodo vos cognovi ex omnibus cognationibus terrae idcirco visitabo super vos omnes iniquitates vestras
AMOS|3|3|numquid ambulabunt duo pariter nisi convenerit eis
AMOS|3|4|numquid rugiet leo in saltu nisi habuerit praedam numquid dabit catulus leonis vocem de cubili suo nisi aliquid adprehenderit
AMOS|3|5|numquid cadet avis in laqueum terrae absque aucupe numquid auferetur laqueus de terra antequam quid ceperit
AMOS|3|6|si clanget tuba in civitate et populus non expavescet si erit malum in civitate quod Dominus non fecit
AMOS|3|7|quia non faciet Dominus Deus verbum nisi revelaverit secretum suum ad servos suos prophetas
AMOS|3|8|leo rugiet quis non timebit Dominus Deus locutus est quis non prophetabit
AMOS|3|9|auditum facite in aedibus Azoti et in aedibus terrae Aegypti et dicite congregamini super montes Samariae et videte insanias multas in medio eius et calumniam patientes in penetrabilibus eius
AMOS|3|10|et nescierunt facere rectum dicit Dominus thesaurizantes iniquitatem et rapinas in aedibus suis
AMOS|3|11|propterea haec dicit Dominus Deus tribulabitur et circumietur terra et detrahetur ex te fortitudo tua et diripientur aedes tuae
AMOS|3|12|haec dicit Dominus quomodo si eruat pastor de ore leonis duo crura aut extremum auriculae sic eruentur filii Israhel qui habitant in Samaria in plaga lectuli et in Damasco grabatti
AMOS|3|13|audite et contestamini in domo Iacob dicit Dominus Deus exercituum
AMOS|3|14|quia in die cum visitare coepero praevaricationes Israhel super eum visitabo et super altaria Bethel et amputabuntur cornua altaris et cadent in terram
AMOS|3|15|et percutiam domum hiemalem cum domo aestiva et peribunt domus eburneae et dissipabuntur aedes multae dicit Dominus
AMOS|4|1|audite verbum hoc vaccae pingues quae estis in monte Samariae quae calumniam facitis egenis et confringitis pauperes quae dicitis dominis vestris adferte et bibemus
AMOS|4|2|iuravit Dominus Deus in sancto suo quia ecce dies venient super vos et levabunt vos in contis et reliquias vestras in ollis ferventibus
AMOS|4|3|et per aperturas exibitis altera contra alteram et proiciemini in Armon dicit Dominus
AMOS|4|4|venite ad Bethel et impie agite ad Galgalam et multiplicate praevaricationem et offerte mane victimas vestras tribus diebus decimas vestras
AMOS|4|5|et sacrificate de fermentato laudem et vocate voluntarias oblationes et adnuntiate sic enim voluistis filii Israhel dicit Dominus Deus
AMOS|4|6|unde et ego dedi vobis stuporem dentium in cunctis urbibus vestris et indigentiam panum in omnibus locis vestris et non estis reversi ad me dicit Dominus
AMOS|4|7|ego quoque prohibui a vobis imbrem cum adhuc tres menses superessent usque ad messem et plui super civitatem unam et super civitatem alteram non plui pars una conpluta est et pars super quam non plui aruit
AMOS|4|8|et venerunt duae et tres civitates ad civitatem unam ut biberent aquam et non sunt satiatae et non redistis ad me dicit Dominus
AMOS|4|9|percussi vos in vento urente et in aurugine multitudinem hortorum vestrorum et vinearum vestrarum oliveta vestra et ficeta vestra comedit eruca et non redistis ad me dicit Dominus
AMOS|4|10|misi in vos mortem in via Aegypti percussi in gladio iuvenes vestros usque ad captivitatem equorum vestrorum et ascendere feci putredinem castrorum vestrorum in nares vestras et non redistis ad me dicit Dominus
AMOS|4|11|subverti vos sicut subvertit Deus Sodomam et Gomorram et facti estis quasi torris raptus de incendio et non redistis ad me dicit Dominus
AMOS|4|12|quapropter haec faciam tibi Israhel postquam autem haec fecero tibi praeparare in occursum Dei tui Israhel
AMOS|4|13|quia ecce formans montes et creans ventum et adnuntians homini eloquium suum faciens matutinam nebulam et gradiens super excelsa terrae Dominus Deus exercituum nomen eius
AMOS|5|1|audite verbum istud quod ego levo super vos planctum domus Israhel cecidit non adiciet ut resurgat
AMOS|5|2|virgo Israhel proiecta est in terram suam non est qui suscitet eam
AMOS|5|3|quia haec dicit Dominus Deus urbs de qua egrediebantur mille relinquentur in ea centum et de qua egrediebantur centum relinquentur in ea decem in domo Israhel
AMOS|5|4|quia haec dicit Dominus domui Israhel quaerite me et vivetis
AMOS|5|5|et nolite quaerere Bethel et in Galgala nolite intrare et in Bersabee non transibitis quia Galgala captiva ducetur et Bethel erit inutilis
AMOS|5|6|quaerite Dominum et vivite ne forte conburatur ut ignis domus Ioseph et devorabit et non erit qui extinguat Bethel
AMOS|5|7|qui convertitis in absinthium iudicium et iustitiam in terra relinquitis
AMOS|5|8|facientem Arcturum et Orionem et convertentem in mane tenebras et diem nocte mutantem qui vocat aquas maris et effundit eas super faciem terrae Dominus nomen eius
AMOS|5|9|qui subridet vastitatem super robustum et depopulationem super potentem adfert
AMOS|5|10|odio habuerunt in porta corripientem et loquentem perfecte abominati sunt
AMOS|5|11|idcirco pro eo quod diripiebatis pauperem et praedam electam tollebatis ab eo domos quadro lapide aedificabitis et non habitabitis in eis vineas amantissimas plantabitis et non bibetis vinum earum
AMOS|5|12|quia cognovi multa scelera vestra et fortia peccata vestra hostes iusti accipientes munus et pauperes in porta deprimentes
AMOS|5|13|ideo prudens in tempore illo tacebit quia tempus malum est
AMOS|5|14|quaerite bonum et non malum ut vivatis et erit Dominus Deus exercituum vobiscum sicut dixistis
AMOS|5|15|odite malum et diligite bonum et constituite in porta iudicium si forte misereatur Dominus Deus exercituum reliquiis Ioseph
AMOS|5|16|propterea haec dicit Dominus Deus exercituum Dominator in omnibus plateis planctus et in cunctis quae foris sunt dicetur vae vae et vocabunt agricolam ad luctum et ad planctum eos qui sciunt plangere
AMOS|5|17|et in omnibus vineis erit planctus quia pertransibo in medio tui dicit Dominus
AMOS|5|18|vae desiderantibus diem Domini ad quid eam vobis dies Domini ista tenebrae et non lux
AMOS|5|19|quomodo si fugiat vir a facie leonis et occurrat ei ursus et ingrediatur domum et innitatur manu sua super parietem et mordeat eum coluber
AMOS|5|20|numquid non tenebrae dies Domini et non lux et caligo et non splendor in ea
AMOS|5|21|odi et proieci festivitates vestras et non capiam odorem coetuum vestrorum
AMOS|5|22|quod si adtuleritis mihi holocaustomata et munera vestra non suscipiam et vota pinguium vestrorum non respiciam
AMOS|5|23|aufer a me tumultum carminum tuorum et cantica lyrae tuae non audiam
AMOS|5|24|et revelabitur quasi aqua iudicium et iustitia quasi torrens fortis
AMOS|5|25|numquid hostias et sacrificium obtulistis mihi in deserto quadraginta annis domus Israhel
AMOS|5|26|et portastis tabernaculum Moloch vestro et imaginem idolorum vestrorum sidus dei vestri quae fecistis vobis
AMOS|5|27|et migrare vos faciam trans Damascum dixit Dominus Deus exercituum nomen eius
AMOS|6|1|vae qui opulenti estis in Sion et confiditis in monte Samariae optimates capita populorum ingredientes pompatice domum Israhel
AMOS|6|2|transite in Chalanne et videte et ite inde in Emath magnam et descendite in Geth Palestinorum et ad optima quaeque regna horum si latior terminus eorum termino vestro est
AMOS|6|3|qui separati estis in diem malum et adpropinquatis solio iniquitatis
AMOS|6|4|qui dormitis in lectis eburneis et lascivitis in stratis vestris qui comeditis agnum de grege et vitulos de medio armenti
AMOS|6|5|qui canitis ad vocem psalterii sicut David putaverunt se habere vasa cantici
AMOS|6|6|bibentes in fialis vinum et optimo unguento delibuti et nihil patiebantur super contritione Ioseph
AMOS|6|7|quapropter nunc migrabunt in capite transmigrantium et auferetur factio lascivientium
AMOS|6|8|iuravit Dominus Deus in anima sua dicit Dominus Deus exercituum detestor ego superbiam Iacob et domos eius odi et tradam civitatem cum habitatoribus suis
AMOS|6|9|quod si reliqui fuerint decem viri in domo una et ipsi morientur
AMOS|6|10|et tollet eum propinquus suus et conburet eum ut efferat ossa de domo et dicet ei qui in penetrabilibus domus est numquid adhuc est apud te
AMOS|6|11|et respondebit finis est et dicet ei tace et non recorderis nominis Domini
AMOS|6|12|quia ecce Dominus mandabit et percutiet domum maiorem ruinis et domum minorem scissionibus
AMOS|6|13|numquid currere queunt in petris equi aut arari potest in bubalis quoniam convertistis in amaritudinem iudicium et fructum iustitiae in absinthium
AMOS|6|14|qui laetamini in nihili qui dicitis numquid non in fortitudine nostra adsumpsimus nobis cornua
AMOS|6|15|ecce enim suscitabo super vos domus Israhel dicit Dominus Deus exercituum gentem et conterent vos ab introitu Emath usque ad torrentem Deserti
AMOS|7|1|haec ostendit mihi Dominus Deus et ecce fictor lucustae in principio germinantium serotini imbris et ecce serotinus post tonsorem regis
AMOS|7|2|et factum est cum consummasset comedere herbam terrae et dixi Domine Deus propitius esto obsecro quis suscitabit Iacob quia parvulus est
AMOS|7|3|misertus est Dominus super hoc non erit dixit Dominus
AMOS|7|4|haec ostendit mihi Dominus Deus et ecce vocabat iudicium ad ignem Dominus Deus et devoravit abyssum multam et comedit simul partem
AMOS|7|5|et dixi Domine Deus quiesce obsecro quis suscitabit Iacob quia parvulus est
AMOS|7|6|misertus est Dominus super hoc sed et istud non erit dixit Dominus Deus
AMOS|7|7|haec ostendit mihi et ecce Dominus stans super murum litum et in manu eius trulla cementarii
AMOS|7|8|et dixit Dominus ad me quid tu vides Amos et dixi trullam cementarii et dixit Dominus ecce ego ponam trullam in medio populi mei Israhel non adiciam ultra superinducere eum
AMOS|7|9|et demolientur excelsa idoli et sanctificationes Israhel desolabuntur et consurgam super domum Hieroboam in gladio
AMOS|7|10|et misit Amasias sacerdos Bethel ad Hieroboam regem Israhel dicens rebellavit contra te Amos in medio domus Israhel non poterit terra sustinere universos sermones eius
AMOS|7|11|haec enim dicit Amos in gladio morietur Hieroboam et Israhel captivus migrabit de terra sua
AMOS|7|12|et dixit Amasias ad Amos qui vides gradere fuge in terram Iuda et comede ibi panem et ibi prophetabis
AMOS|7|13|et in Bethel non adicies ultra ut prophetes quia sanctificatio regis est et domus regni est
AMOS|7|14|et respondit Amos et dixit ad Amasiam non sum propheta et non sum filius prophetae sed armentarius ego sum vellicans sycomoros
AMOS|7|15|et tulit me Dominus cum sequerer gregem et dixit ad me Dominus vade propheta ad populum meum Israhel
AMOS|7|16|et nunc audi verbum Domini tu dicis non prophetabis super Israhel et non stillabis super domum idoli
AMOS|7|17|propter hoc haec dicit Dominus uxor tua in civitate fornicabitur et filii tui et filiae tuae in gladio cadent et humus tua funiculo metietur et tu in terra polluta morieris et Israhel captivus migrabit de terra sua
AMOS|8|1|haec ostendit mihi Dominus Deus et ecce uncinus pomorum
AMOS|8|2|et dixit quid tu vides Amos et dixi uncinum pomorum et dixit Dominus ad me venit finis super populum meum Israhel non adiciam ultra ut pertranseam eum
AMOS|8|3|et stridebunt cardines templi in die illa dicit Dominus Deus multi morientur in omni loco proicietur silentium
AMOS|8|4|audite hoc qui conteritis pauperem et deficere facitis egenos terrae
AMOS|8|5|dicentes quando transibit mensis et venundabimus merces et sabbatum et aperiemus frumentum ut inminuamus mensuram et augeamus siclum et subponamus stateras dolosas
AMOS|8|6|ut possideamus in argento egenos et pauperes pro calciamentis et quisquilias frumenti vendamus
AMOS|8|7|iuravit Dominus in superbia Iacob si oblitus fuero usque ad finem omnia opera eorum
AMOS|8|8|numquid super isto non commovebitur terra et lugebit omnis habitator eius et ascendet quasi fluvius universus et eicietur et defluet quasi rivus Aegypti
AMOS|8|9|et erit in die illa dicit Dominus occidet sol meridie et tenebrescere faciam terram in die luminis
AMOS|8|10|et convertam festivitates vestras in luctum et omnia cantica vestra in planctum et inducam super omne dorsum vestrum saccum et super omne caput calvitium et ponam eam quasi luctum unigeniti et novissima eius quasi diem amarum
AMOS|8|11|ecce dies veniunt dicit Dominus et mittam famem in terram non famem panis neque sitim aquae sed audiendi verbum Domini
AMOS|8|12|et commovebuntur a mari usque ad mare et ab aquilone usque ad orientem circumibunt quaerentes verbum Domini et non invenient
AMOS|8|13|in die illa deficient virgines pulchrae et adulescentes in siti
AMOS|8|14|qui iurant in delicto Samariae et dicunt vivit deus tuus Dan et vivit via Bersabee et cadent et non resurgent ultra
AMOS|9|1|vidi Dominum stantem super altare et dixit percute cardinem et commoveantur superliminaria avaritia enim in capite omnium et novissimum eorum in gladio interficiam non erit fuga eis fugiet et non salvabitur ex eis qui fugerit
AMOS|9|2|si descenderint usque ad infernum inde manus mea educet eos et si ascenderint usque ad caelum inde detraham eos
AMOS|9|3|et si absconditi fuerint in vertice Carmeli inde scrutans auferam eos et si celaverint se ab oculis meis in fundo maris ibi mandabo serpenti et mordebit eos
AMOS|9|4|et si abierint in captivitatem coram inimicis suis ibi mandabo gladio et occidet eos et ponam oculos meos super eos in malum et non in bonum
AMOS|9|5|et Dominus Deus exercituum qui tangit terram et tabescet et lugebunt omnes habitantes in ea et ascendet sicut rivus omnis et defluet sicut fluvius Aegypti
AMOS|9|6|qui aedificat in caelo ascensionem suam et fasciculum suum super terram fundavit qui vocat aquas maris et effundit eas super faciem terrae Dominus nomen eius
AMOS|9|7|numquid non ut filii Aethiopum vos estis mihi filii Israhel ait Dominus numquid non Israhel ascendere feci de terra Aegypti et Palestinos de Cappadocia et Syros de Cyrene
AMOS|9|8|ecce oculi Domini Dei super regnum peccans et conteram illud a facie terrae verumtamen conterens non conteram domum Iacob dicit Dominus
AMOS|9|9|ecce enim ego mandabo et concutiam in omnibus gentibus domum Israhel sicut concutitur in cribro et non cadet lapillus super terram
AMOS|9|10|in gladio morientur omnes peccatores populi mei qui dicunt non adpropinquabit et non veniet super nos malum
AMOS|9|11|in die illo suscitabo tabernaculum David quod cecidit et reaedificabo aperturas murorum eius et ea quae corruerant instaurabo et reaedificabo eum sicut diebus antiquis
AMOS|9|12|ut possideant reliquias Idumeae et omnes nationes eo quod invocatum sit nomen meum super eos dicit Dominus faciens haec
AMOS|9|13|ecce dies veniunt dicit Dominus et conprehendet arator messorem et calcator uvae mittentem semen et stillabunt montes dulcedinem et omnes colles culti erunt
AMOS|9|14|et convertam captivitatem populi mei Israhel et aedificabunt civitates desertas et habitabunt et plantabunt vineas et bibent vinum earum et facient hortos et comedent fructus eorum
OBAD|1|1|visio Abdiae haec dicit Dominus Deus ad Edom auditum audivimus a Domino et legatum ad gentes misit surgite et consurgamus adversum eum in proelium
OBAD|1|2|ecce parvulum te dedi in gentibus contemptibilis tu es valde
OBAD|1|3|superbia cordis tui extulit te habitantem in scissuris petrae exaltantem solium suum qui dicit in corde suo quis detrahet me in terram
OBAD|1|4|si exaltatus fueris ut aquila et si inter sidera posueris nidum tuum inde detraham te dicit Dominus
OBAD|1|5|si fures introissent ad te si latrones per noctem quomodo conticuisses nonne furati essent sufficientia sibi si vindemiatores introissent ad te numquid saltim racemos reliquissent tibi
OBAD|1|6|quomodo scrutati sunt Esau investigaverunt abscondita eius
OBAD|1|7|usque ad terminum emiserunt te omnes viri foederis tui inluserunt tibi invaluerunt adversum te viri pacis tuae qui comedunt tecum ponent insidias subter te non est prudentia in eo
OBAD|1|8|numquid non in die illa dicit Dominus perdam sapientes de Idumea et prudentiam de monte Esau
OBAD|1|9|et timebunt fortes tui a meridie ut intereat vir de monte Esau
OBAD|1|10|propter interfectionem et propter iniquitatem in fratrem tuum Iacob operiet te confusio et peribis in aeternum
OBAD|1|11|in die cum stares adversus quando capiebant alieni exercitum eius et extranei ingrediebantur portas eius et super Hierusalem mittebant sortem tu quoque eras quasi unus ex eis
OBAD|1|12|et non despicies in die fratris tui in die peregrinationis eius et non laetaberis super filios Iuda in die perditionis eorum et non magnificabis os tuum in die angustiae
OBAD|1|13|neque ingredieris portam populi mei in die ruinae eorum neque despicies et tu in malis eius in die vastitatis illius et non emitteris adversum exercitum eius in die vastitatis illius
OBAD|1|14|neque stabis in exitibus ut interficias eos qui fugerint et non concludes reliquos eius in die tribulationis
OBAD|1|15|quoniam iuxta est dies Domini super omnes gentes sicut fecisti fiet tibi retributionem tuam convertet in caput tuum
OBAD|1|16|quomodo enim bibisti super montem sanctum meum bibent omnes gentes iugiter et bibent et absorbent et erunt quasi non sint
OBAD|1|17|et in monte Sion erit salvatio et erit sanctus et possidebit domus Iacob eos qui se possederant
OBAD|1|18|et erit domus Iacob ignis et domus Ioseph flamma et domus Esau stipula et succendentur in eis et devorabunt eos et non erunt reliquiae domus Esau quia Dominus locutus est
OBAD|1|19|et hereditabunt hii qui ad austrum montem Esau et qui in campestribus Philisthim et possidebunt regionem Ephraim et regionem Samariae et Beniamin possidebit Galaad
OBAD|1|20|et transmigratio exercitus huius filiorum Israhel omnia Chananeorum usque ad Saraptham et transmigratio Hierusalem quae in Bosforo est possidebit civitates austri
OBAD|1|21|et ascendent salvatores in montem Sion iudicare montem Esau et erit Domino regnum
JONAH|1|1|et factum est verbum Domini ad Ionam filium Amathi dicens
JONAH|1|2|surge vade in Nineven civitatem grandem et praedica in ea quia ascendit malitia eius coram me
JONAH|1|3|et surrexit Iona ut fugeret in Tharsis a facie Domini et descendit Ioppen et invenit navem euntem in Tharsis et dedit naulum eius et descendit in eam ut iret cum eis in Tharsis a facie Domini
JONAH|1|4|Dominus autem misit ventum magnum in mari et facta est tempestas magna in mari et navis periclitabatur conteri
JONAH|1|5|et timuerunt nautae et clamaverunt viri ad deum suum et miserunt vasa quae erant in navi in mare ut adleviaretur ab eis et Iona descendit ad interiora navis et dormiebat sopore gravi
JONAH|1|6|et accessit ad eum gubernator et dixit ei quid tu sopore deprimeris surge invoca Deum tuum si forte recogitet Deus de nobis et non pereamus
JONAH|1|7|et dixit vir ad collegam suum venite et mittamus sortes et sciamus quare hoc malum sit nobis et miserunt sortes et cecidit sors super Ionam
JONAH|1|8|et dixerunt ad eum indica nobis cuius causa malum istud sit nobis quod est opus tuum quae terra tua et quo vel ex quo populo es tu
JONAH|1|9|et dixit ad eos Hebraeus ego sum et Dominum Deum caeli ego timeo qui fecit mare et aridam
JONAH|1|10|et timuerunt viri timore magno et dixerunt ad eum quid hoc fecisti cognoverunt enim viri quod a facie Domini fugeret quia indicaverat eis
JONAH|1|11|et dixerunt ad eum quid faciemus tibi et cessabit mare a nobis quia mare ibat et intumescebat
JONAH|1|12|et dixit ad eos tollite me et mittite in mare et cessabit mare a vobis scio enim ego quoniam propter me tempestas grandis haec super vos
JONAH|1|13|et remigabant viri ut reverterentur ad aridam et non valebant quia mare ibat et intumescebat super eos
JONAH|1|14|et clamaverunt ad Dominum et dixerunt quaesumus Domine ne pereamus in anima viri istius et ne des super nos sanguinem innocentem quia tu Domine sicut voluisti fecisti
JONAH|1|15|et tulerunt Ionam et miserunt in mare et stetit mare a fervore suo
JONAH|1|16|et timuerunt viri timore magno Dominum et immolaverunt hostias Domino et voverunt vota
JONAH|2|1|et praeparavit Dominus piscem grandem ut degluttiret Ionam et erat Iona in ventre piscis tribus diebus et tribus noctibus
JONAH|2|2|et oravit Iona ad Dominum Deum suum de utero piscis
JONAH|2|3|et dixit clamavi de tribulatione mea ad Dominum et exaudivit me de ventre inferni clamavi et exaudisti vocem meam
JONAH|2|4|et proiecisti me in profundum in corde maris et flumen circumdedit me omnes gurgites tui et fluctus tui super me transierunt
JONAH|2|5|et ego dixi abiectus sum a conspectu oculorum tuorum verumtamen rursus videbo templum sanctum tuum
JONAH|2|6|circumdederunt me aquae usque ad animam abyssus vallavit me pelagus operuit caput meum
JONAH|2|7|ad extrema montium descendi terrae vectes concluserunt me in aeternum et sublevabis de corruptione vitam meam Domine Deus meus
JONAH|2|8|cum angustiaretur in me anima mea Domini recordatus sum ut veniat ad te oratio mea ad templum sanctum tuum
JONAH|2|9|qui custodiunt vanitates frustra misericordiam suam derelinquunt
JONAH|2|10|ego autem in voce laudis immolabo tibi quaecumque vovi reddam pro salute Domino
JONAH|2|11|et dixit Dominus pisci et evomuit Ionam in aridam
JONAH|3|1|et factum est verbum Domini ad Ionam secundo dicens
JONAH|3|2|surge vade ad Nineven civitatem magnam et praedica in ea praedicationem quam ego loquor ad te
JONAH|3|3|et surrexit Iona et abiit in Nineven iuxta verbum Domini et Nineve erat civitas magna Dei itinere dierum trium
JONAH|3|4|et coepit Iona introire in civitatem itinere diei unius et clamavit et dixit adhuc quadraginta dies et Nineve subvertetur
JONAH|3|5|et crediderunt viri ninevitae in Deo et praedicaverunt ieiunium et vestiti sunt saccis a maiore usque ad minorem
JONAH|3|6|et pervenit verbum ad regem Nineve et surrexit de solio suo et abiecit vestimentum suum a se et indutus est sacco et sedit in cinere
JONAH|3|7|et clamavit et dixit in Nineve ex ore regis et principum eius dicens homines et iumenta et boves et pecora non gustent quicquam nec pascantur et aquam non bibant
JONAH|3|8|et operiantur saccis homines et iumenta et clament ad Dominum in fortitudine et convertatur vir a via sua mala et ab iniquitate quae est in manibus eorum
JONAH|3|9|quis scit si convertatur et ignoscat Deus et revertatur a furore irae suae et non peribimus
JONAH|3|10|et vidit Deus opera eorum quia conversi sunt a via sua mala et misertus est Deus super malitiam quam locutus fuerat ut faceret eis et non fecit
JONAH|4|1|et adflictus est Iona adflictione magna et iratus est
JONAH|4|2|et oravit ad Dominum et dixit obsecro Domine numquid non hoc est verbum meum cum adhuc essem in terra mea propter hoc praeoccupavi ut fugerem in Tharsis scio enim quia tu Deus clemens et misericors es patiens et multae miserationis et ignoscens super malitia
JONAH|4|3|et nunc Domine tolle quaeso animam meam a me quia melior est mihi mors quam vita
JONAH|4|4|et dixit Dominus putasne bene irasceris tu
JONAH|4|5|et egressus est Iona de civitate et sedit contra orientem civitatis et fecit sibimet ibi umbraculum et sedebat subter eum in umbra donec videret quid accideret civitati
JONAH|4|6|et praeparavit Dominus Deus hederam et ascendit super caput Ionae ut esset umbra super caput eius et protegeret eum laboraverat enim et laetatus est Iona super hedera laetitia magna
JONAH|4|7|et paravit Deus vermem ascensu diluculo in crastinum et percussit hederam et exaruit
JONAH|4|8|et cum ortus fuisset sol praecepit Dominus vento calido et urenti et percussit sol super caput Ionae et aestuabat et petivit animae suae ut moreretur et dixit melius est mihi mori quam vivere
JONAH|4|9|et dixit Dominus ad Ionam putasne bene irasceris tu super hederam et dixit bene irascor ego usque ad mortem
JONAH|4|10|et dixit Dominus tu doles super hederam in qua non laborasti neque fecisti ut cresceret quae sub una nocte nata est et una nocte periit
JONAH|4|11|et ego non parcam Nineve civitati magnae in qua sunt plus quam centum viginti milia hominum qui nesciunt quid sit inter dexteram et sinistram suam et iumenta multa
MIC|1|1|verbum Domini quod factum est ad Micham Morasthiten in diebus Ioatham Ahaz Ezechiae regum Iuda quod vidit super Samariam et Hierusalem
MIC|1|2|audite populi omnes et adtendat terra et plenitudo eius et sit Dominus Deus vobis in testem Dominus de templo sancto suo
MIC|1|3|quia ecce Dominus egreditur de loco suo et descendet et calcabit super excelsa terrae
MIC|1|4|et consumentur montes subtus eum et valles scindentur sicut cera a facie ignis sicut aquae quae decurrunt in praeceps
MIC|1|5|in scelere Iacob omne istud et in peccatis domus Israhel quod scelus Iacob nonne Samaria et quae excelsa Iudae nonne Hierusalem
MIC|1|6|et ponam Samariam quasi acervum lapidum in agro cum plantatur vinea et detraham in vallem lapides eius et fundamenta eius revelabo
MIC|1|7|et omnia sculptilia eius concidentur et omnes mercedes eius conburentur igni et omnia idola eius ponam in perditionem quia de mercedibus meretricis congregata sunt et usque ad mercedem meretricis revertentur
MIC|1|8|super hoc plangam et ululabo vadam spoliatus et nudus faciam planctum velut draconum et luctum quasi strutionum
MIC|1|9|quia desperata est plaga eius quia venit usque ad Iudam tetigit portam populi mei usque ad Hierusalem
MIC|1|10|in Geth nolite adnuntiare lacrimis ne ploretis in domo Pulveris pulvere vos conspergite
MIC|1|11|et transite vobis habitatio Pulchra confusa ignominia non est egressa quae habitat in Exitu planctum domus Vicinae accipiet ex vobis quae stetit sibimet
MIC|1|12|quia infirmata est in bonum quae habitat in Amaritudinibus quia descendit malum a Domino in portam Hierusalem
MIC|1|13|tumultus quadrigae stuporis habitanti Lachis principium peccati est filiae Sion quia in te inventa sunt scelera Israhel
MIC|1|14|propterea dabit emissarios super hereditatem Geth domus Mendacii in deceptionem regibus Israhel
MIC|1|15|adhuc heredem adducam tibi quae habitas in Maresa usque Adollam veniet gloria Israhel
MIC|1|16|decalvare et tondere super filios deliciarum tuarum dilata calvitium tuum sicut aquila quoniam captivi ducti sunt ex te
MIC|2|1|vae qui cogitatis inutile et operamini malum in cubilibus vestris in luce matutina faciunt illud quoniam contra Deum est manus eorum
MIC|2|2|et concupierunt agros et violenter tulerunt et domos rapuerunt et calumniabantur virum et domum eius virum et hereditatem eius
MIC|2|3|idcirco haec dicit Dominus ecce ego cogito super familiam istam malum unde non auferetis colla vestra et non ambulabitis superbi quoniam tempus pessimum est
MIC|2|4|in die illa sumetur super vos parabola et cantabitur canticum cum suavitate dicentium depopulatione vastati sumus pars populi mei commutata est quomodo recedet a me cum revertatur qui regiones nostras dividat
MIC|2|5|propter hoc non erit tibi mittens funiculum sortis in coetu Domini
MIC|2|6|ne loquamini loquentes non stillabit super istos non conprehendet confusio
MIC|2|7|dicit domus Iacob numquid adbreviatus est spiritus Domini aut tales sunt cogitationes eius nonne verba mea bona sunt cum eo qui recte graditur
MIC|2|8|et e contrario populus meus in adversarium consurrexit desuper tunica pallium sustulistis eos qui transiebant simpliciter convertistis in bellum
MIC|2|9|mulieres populi mei eiecistis de domo deliciarum suarum a parvulis earum tulistis laudem meam in perpetuum
MIC|2|10|surgite et ite quia non habetis hic requiem propter inmunditiam eius corrumpetur putredine pessima
MIC|2|11|utinam non essem vir habens spiritum et mendacium potius loquerer stillabo tibi in vinum et in ebrietatem et erit super quem stillatur populus iste
MIC|2|12|congregatione congregabo Iacob totum te in unum conducam reliquias Israhel pariter ponam illum quasi gregem in ovili quasi pecus in medio caularum tumultuabuntur a multitudine hominum
MIC|2|13|ascendet enim pandens iter ante eos divident et transibunt portam et egredientur per eam et transibit rex eorum coram eis et Dominus in capite eorum
MIC|3|1|et dixi audite principes Iacob et duces domus Israhel numquid non vestrum est scire iudicium
MIC|3|2|qui odio habetis bonum et diligitis malum qui violenter tollitis pelles eorum desuper eos et carnem eorum desuper ossibus eorum
MIC|3|3|qui comederunt carnem populi mei et pellem eorum desuper excoriaverunt et ossa eorum confregerunt et conciderunt sicut in lebete et quasi carnem in medio ollae
MIC|3|4|tunc clamabunt ad Dominum et non exaudiet eos et abscondet faciem suam ab eis in tempore illo sicut nequiter egerunt in adinventionibus suis
MIC|3|5|haec dicit Dominus super prophetas qui seducunt populum meum qui mordent dentibus suis et praedicant pacem et si quis non dederit in ore eorum quippiam sanctificant super eum proelium
MIC|3|6|propterea nox vobis pro visione erit et tenebrae vobis pro divinatione et occumbet sol super prophetas et obtenebrabitur super eos dies
MIC|3|7|et confundentur qui vident visiones et confundentur divini et operient vultus suos omnes quia non est responsum Dei
MIC|3|8|verumtamen ego repletus sum fortitudine spiritus Domini iudicio et virtute ut adnuntiem Iacob scelus suum et Israhel peccatum suum
MIC|3|9|audite haec principes domus Iacob et iudices domus Israhel qui abominamini iudicium et omnia recta pervertitis
MIC|3|10|qui aedificatis Sion in sanguinibus et Hierusalem in iniquitate
MIC|3|11|principes eius in muneribus iudicabant et sacerdotes eius in mercede docebant et prophetae eius in pecunia divinabant et super Dominum requiescebant dicentes numquid non Dominus in medio nostrum non venient super nos mala
MIC|3|12|propter hoc causa vestri Sion quasi ager arabitur et Hierusalem quasi acervus lapidum erit et mons templi in excelsa silvarum
MIC|4|1|et in novissimo dierum erit mons domus Domini praeparatus in vertice montium et sublimis super colles et fluent ad eum populi
MIC|4|2|et properabunt gentes multae et dicent venite ascendamus ad montem Domini et ad domum Dei Iacob et docebit nos de viis suis et ibimus in semitis eius quia de Sion egredietur lex et verbum Domini de Hierusalem
MIC|4|3|et iudicabit inter populos multos et corripiet gentes fortes usque in longinquum et concident gladios suos in vomeres et hastas suas in ligones non sumet gens adversus gentem gladium et non discent ultra belligerare
MIC|4|4|et sedebit vir subtus vineam suam et subtus ficum suam et non erit qui deterreat quia os Domini exercituum locutum est
MIC|4|5|quia omnes populi ambulabunt unusquisque in nomine dei sui nos autem ambulabimus in nomine Domini Dei nostri in aeternum et ultra
MIC|4|6|in die illa dicit Dominus congregabo claudicantem et eam quam eieceram colligam et quam adflixeram
MIC|4|7|et ponam claudicantem in reliquias et eam quae laboraverat in gentem robustam et regnabit Dominus super eos in monte Sion ex hoc nunc et usque in aeternum
MIC|4|8|et tu turris Gregis nebulosa filiae Sion usque ad te veniet et veniet potestas prima regnum filiae Hierusalem
MIC|4|9|nunc quare maerore contraheris numquid rex non est tibi aut consiliarius tuus periit quia conprehendit te dolor sicut parturientem
MIC|4|10|dole et satage filia Sion quasi parturiens quia nunc egredieris de civitate et habitabis in regione et venies usque ad Babylonem ibi liberaberis ibi redimet te Dominus de manu inimicorum tuorum
MIC|4|11|et nunc congregatae sunt super te gentes multae quae dicunt lapidetur et aspiciat in Sion oculus noster
MIC|4|12|ipsi autem non cognoverunt cogitationes Domini et non intellexerunt consilium eius quia congregavit eos quasi faenum areae
MIC|4|13|surge et tritura filia Sion quia cornu tuum ponam ferreum et ungulas tuas ponam aereas et comminues populos multos et interficiam Domino rapinas eorum et fortitudinem eorum Domino universae terrae
MIC|5|1|nunc vastaberis filia latronis obsidionem posuerunt super nos in virga percutient maxillam iudicis Israhel
MIC|5|2|et tu Bethleem Ephrata parvulus es in milibus Iuda ex te mihi egredietur qui sit dominator in Israhel et egressus eius ab initio a diebus aeternitatis
MIC|5|3|propter hoc dabit eos usque ad tempus in quo parturiens pariet reliquiae fratrum eius convertentur ad filios Israhel
MIC|5|4|et stabit et pascet in fortitudine Domini in sublimitate nominis Domini Dei sui et convertentur quia nunc magnificabitur usque ad terminos terrae
MIC|5|5|et erit iste pax Assyrius cum venerit in terram nostram et quando calcaverit in domibus nostris et suscitabimus super eum septem pastores et octo primates homines
MIC|5|6|et pascent terram Assur in gladio et terram Nemrod in lanceis eius et liberabit ab Assur cum venerit in terram nostram et cum calcaverit in finibus nostris
MIC|5|7|et erunt reliquiae Iacob in medio populorum multorum quasi ros a Domino et quasi stillae super herbam quae non expectat virum et non praestolatur filios hominum
MIC|5|8|et erunt reliquiae Iacob in gentibus in medio populorum multorum quasi leo in iumentis silvarum et quasi catulus leonis in gregibus pecorum qui cum transierit et conculcaverit et ceperit non est qui eruat
MIC|5|9|exaltabitur manus tua super hostes tuos et omnes inimici tui interibunt
MIC|5|10|et erit in die illa dicit Dominus auferam equos tuos de medio tui et disperdam quadrigas tuas
MIC|5|11|et perdam civitates terrae tuae et destruam omnes munitiones tuas et auferam maleficia de manu tua et divinationes non erunt in te
MIC|5|12|et perire faciam sculptilia tua et statuas tuas de medio tui et non adorabis ultra opera manuum tuarum
MIC|5|13|et evellam lucos tuos de medio tui et conteram civitates tuas
MIC|5|14|et faciam in furore et in indignatione ultionem in omnibus gentibus quae non audierunt
MIC|6|1|audite quae Dominus loquitur surge contende iudicio adversum montes et audiant colles vocem tuam
MIC|6|2|audiant montes iudicium Domini et fortia fundamenta terrae quia iudicium Domini cum populo suo et cum Israhel diiudicabitur
MIC|6|3|populus meus quid feci tibi et quid molestus fui tibi responde mihi
MIC|6|4|quia eduxi te de terra Aegypti et de domo servientium liberavi te et misi ante faciem tuam Mosen et Aaron et Mariam
MIC|6|5|populus meus memento quaeso quid cogitaverit Balac rex Moab et quid responderit ei Balaam filius Beor de Setthim usque ad Galgalam ut cognosceret iustitias Domini
MIC|6|6|quid dignum offeram Domino curvem genu Deo excelso numquid offeram ei holocaustomata et vitulos anniculos
MIC|6|7|numquid placari potest Dominus in milibus arietum aut in multis milibus hircorum pinguium numquid dabo primogenitum meum pro scelere meo fructum ventris mei pro peccato animae meae
MIC|6|8|indicabo tibi o homo quid sit bonum et quid Dominus quaerat a te utique facere iudicium et diligere misericordiam et sollicitum ambulare cum Deo tuo
MIC|6|9|vox Domini ad civitatem clamat et salus erit timentibus nomen tuum audite tribus et quis adprobabit illud
MIC|6|10|adhuc ignis in domo impii thesauri iniquitatis et mensura minor irae plena
MIC|6|11|numquid iustificabo stateram impiam et saccelli pondera dolosa
MIC|6|12|in quibus divites eius repleti sunt iniquitate et habitantes in ea loquebantur mendacium et lingua eorum fraudulenta in ore eorum
MIC|6|13|et ego ergo coepi percutere te perditione super peccatis tuis
MIC|6|14|tu comedes et non saturaberis et humiliatio tua in medio tui et adprehendes et non salvabis et quos salvaveris in gladium dabo
MIC|6|15|tu seminabis et non metes tu calcabis olivam et non ungueris oleo et mustum et non bibes vinum
MIC|6|16|et custodisti praecepta Omri et omne opus domus Achab et ambulasti in voluntatibus eorum ut darem te in perditionem et habitantes in ea in sibilum et obprobrium populi mei portabitis
MIC|7|1|vae mihi quia factus sum sicut qui colligit in autumno racemos vindemiae non est botrus ad comedendum praecoquas ficus desideravit anima mea
MIC|7|2|periit sanctus de terra et rectus in hominibus non est omnes in sanguine insidiantur vir fratrem suum venatur ad mortem
MIC|7|3|malum manuum suarum dicunt bonum princeps postulat et iudex in reddendo est et magnus locutus est desiderium animae suae et conturbaverunt eam
MIC|7|4|qui optimus in eis est quasi paliurus et qui rectus quasi spina de sepe dies speculationis tuae visitatio tua venit nunc erit vastitas eorum
MIC|7|5|nolite credere amico et nolite confidere in duce ab ea quae dormit in sinu tuo custodi claustra oris tui
MIC|7|6|quia filius contumeliam facit patri filia consurgit adversus matrem suam nurus contra socrum suam inimici hominis domestici eius
MIC|7|7|ego autem ad Dominum aspiciam expectabo Deum salvatorem meum audiet me Deus meus
MIC|7|8|ne laeteris inimica mea super me quia cecidi consurgam cum sedero in tenebris Dominus lux mea est
MIC|7|9|iram Domini portabo quoniam peccavi ei donec iudicet causam meam et faciat iudicium meum educet me in lucem videbo in iustitiam eius
MIC|7|10|et aspiciet inimica mea et operietur confusione quae dicit ad me ubi est Dominus Deus tuus oculi mei videbunt in eam nunc erit in conculcationem ut lutum platearum
MIC|7|11|dies ut aedificentur maceriae tuae in die illa longe fiet lex
MIC|7|12|in die illa et usque ad te veniet Assur et usque ad civitates munitas et a civitatibus munitis usque ad flumen et ad mare de mari et ad montem de monte
MIC|7|13|et erit terra in desolationem propter habitatores suos et propter fructum cogitationum eorum
MIC|7|14|pasce populum tuum in virga tua gregem hereditatis tuae habitantes solos in saltu in medio Carmeli pascentur Basan et Galaad iuxta dies antiquos
MIC|7|15|secundum dies egressionis tuae de terra Aegypti ostendam ei mirabilia
MIC|7|16|videbunt gentes et confundentur super omni fortitudine sua ponent manus super os aures eorum surdae erunt
MIC|7|17|lingent pulverem sicut serpens velut reptilia terrae proturbabuntur de aedibus suis Dominum Deum nostrum desiderabunt et timebunt te
MIC|7|18|quis Deus similis tui qui aufers iniquitatem et transis peccatum reliquiarum hereditatis tuae non inmittet ultra furorem suum quoniam volens misericordiam est
MIC|7|19|revertetur et miserebitur nostri deponet iniquitates nostras et proiciet in profundum maris omnia peccata nostra
MIC|7|20|dabis veritatem Iacob misericordiam Abraham quae iurasti patribus nostris a diebus antiquis
NAH|1|1|onus Nineve liber visionis Naum Helcesei
NAH|1|2|Deus aemulator et ulciscens Dominus ulciscens Dominus et habens furorem ulciscens Dominus in hostes suos et irascens ipse inimicis suis
NAH|1|3|Dominus patiens et magnus fortitudine et mundans non faciet innocentem Dominus in tempestate et turbine viae eius et nebulae pulvis pedum eius
NAH|1|4|increpans mare et exsiccans illud et omnia flumina ad desertum deducens infirmatus est Basan et Carmelus et flos Libani elanguit
NAH|1|5|montes commoti sunt ab eo et colles adsolati sunt et contremuit terra a facie eius et orbis et omnes habitantes in eo
NAH|1|6|ante faciem indignationis eius quis stabit et quis resistet in ira furoris eius indignatio eius effusa est ut ignis et petrae dissolutae sunt ab eo
NAH|1|7|bonus Dominus et confortans in die tribulationis et sciens sperantes in se
NAH|1|8|et in diluvio praetereunte consummationem faciet loci eius et inimicos eius persequentur tenebrae
NAH|1|9|quid cogitatis contra Dominum consummationem ipse faciet non consurget duplex tribulatio
NAH|1|10|quia sicut spinae se invicem conplectuntur sic convivium eorum pariter potantium consumentur quasi stipula ariditate plena
NAH|1|11|ex te exivit cogitans contra Dominum malitiam mente pertractans praevaricationem
NAH|1|12|haec dicit Dominus si perfecti fuerint et ita plures sic quoque adtondentur et pertransibit adflixi te et non adfligam te ultra
NAH|1|13|et nunc conteram virgam eius de dorso tuo et vincula tua disrumpam
NAH|1|14|et praecipiet super te Dominus non seminabitur ex nomine tuo amplius de domo Dei tui interficiam sculptile et conflatile ponam sepulchrum tuum quia inhonoratus es
NAH|1|15|ecce super montes pedes evangelizantis et adnuntiantis pacem celebra Iuda festivitates tuas et redde vota tua quia non adiciet ultra ut pertranseat in te Belial universus interiit
NAH|2|1|ascendit qui dispergat coram te qui custodit obsidionem contemplare viam conforta lumbos robora virtutem valde
NAH|2|2|quia reddidit Dominus superbiam Iacob sicut superbiam Israhel quia vastatores dissipaverunt eos et propagines eorum corruperunt
NAH|2|3|clypeus fortium eius ignitus viri exercitus in coccineis igneae habenae currus in die praeparationis eius et agitatores consopiti sunt
NAH|2|4|in itineribus conturbati sunt quadrigae conlisae sunt in plateis aspectus eorum quasi lampades quasi fulgura discurrentia
NAH|2|5|recordabitur fortium suorum ruent in itineribus suis velociter ascendent muros eius et praeparabitur umbraculum
NAH|2|6|portae fluviorum apertae sunt et templum ad solum dirutum
NAH|2|7|et miles captivus abductus est et ancillae eius minabantur gementes ut columbae murmurantes in cordibus suis
NAH|2|8|et Nineve quasi piscina aquarum aquae eius ipsi vero fugerunt state state et non est qui revertatur
NAH|2|9|diripite argentum diripite aurum et non est finis divitiarum ex omnibus vasis desiderabilibus
NAH|2|10|dissipata et scissa et dilacerata et cor tabescens et dissolutio geniculorum et defectio in cunctis renibus et facies omnium sicut nigredo ollae
NAH|2|11|ubi est habitaculum leonum et pascua catulorum leonum ad quam ivit leo ut ingrederetur illuc catulus leonis et non est qui exterreat
NAH|2|12|leo cepit sufficienter catulis suis et necavit leaenis suis et implevit praeda speluncas suas et cubile suum rapina
NAH|2|13|ecce ego ad te dicit Dominus exercituum et succendam usque ad fumum quadrigas eius et leunculos tuos comedet gladius et exterminabo de terra praedam tuam et non audietur ultra vox nuntiorum tuorum
NAH|3|1|vae civitas sanguinum universa mendacii dilaceratione plena non recedet a te rapina
NAH|3|2|vox flagelli et vox impetus rotae et equi frementis et quadrigae ferventis equitis ascendentis
NAH|3|3|et micantis gladii et fulgurantis hastae et multitudinis interfectae et gravis ruinae nec est finis cadaverum et corruent in corporibus suis
NAH|3|4|propter multitudinem fornicationum meretricis speciosae et gratae et habentis maleficia quae vendidit gentes in fornicationibus suis et familias in maleficiis suis
NAH|3|5|ecce ego ad te dicit Dominus exercituum et revelabo pudenda tua in facie tua et ostendam gentibus nuditatem tuam et regnis ignominiam tuam
NAH|3|6|et proiciam super te abominationes et contumeliis te adficiam et ponam te in exemplum
NAH|3|7|et erit omnis qui viderit te resiliet a te et dicet vastata est Nineve quis commovebit super te caput unde quaeram consolatorem tibi
NAH|3|8|numquid melior es ab Alexandria populorum quae habitat in fluminibus aqua in circuitu eius cuius divitiae mare aquae muri eius
NAH|3|9|Aethiopia fortitudo et Aegyptus et non est finis Africa et Lybies fuerunt in auxilio tuo
NAH|3|10|sed et ipsa in transmigrationem ducta est in captivitatem parvuli eius elisi sunt in capite omnium viarum et super inclitos eius miserunt sortem et omnes optimates eius confixi sunt in conpedibus
NAH|3|11|et tu ergo inebriaberis eris despecta et tu quaeres auxilium ab inimico
NAH|3|12|omnes munitiones tuae sicuti ficus cum grossis suis si concussae fuerint cadent in os comedentis
NAH|3|13|ecce populus tuus mulieres in medio tui inimicis tuis adapertione pandentur portae terrae tuae devorabit ignis vectes tuos
NAH|3|14|aquam propter obsidionem hauri tibi extrue munitiones tuas intra in lutum et calca subigens tene laterem
NAH|3|15|ibi comedet te ignis peribis gladio devorabit te ut bruchus congregare ut bruchus multiplicare ut lucusta
NAH|3|16|plures fecisti negotiationes tuas quam stellae sunt caeli bruchus expansus est et avolavit
NAH|3|17|custodes tui quasi lucustae et parvuli tui quasi lucustae lucustarum quae considunt in sepibus in die frigoris sol ortus est et avolaverunt et non est cognitus locus earum ubi fuerint
NAH|3|18|dormitaverunt pastores tui rex Assur sepelientur principes tui latitavit populus tuus in montibus et non est qui congreget
NAH|3|19|non est obscura contritio tua pessima est plaga tua omnes qui audierunt auditionem tuam conpresserunt manum super te quia super quem non transiit malitia tua semper
HAB|1|1|onus quod vidit Abacuc propheta
HAB|1|2|usquequo Domine clamabo et non exaudies vociferabor ad te vim patiens et non salvabis
HAB|1|3|quare ostendisti mihi iniquitatem et laborem videre praeda et iniustitia contra me et factum est iudicium et contradictio potentior
HAB|1|4|propter hoc lacerata est lex et non pervenit usque ad finem iudicium quia impius praevalet adversus iustum propterea egreditur iudicium perversum
HAB|1|5|aspicite in gentibus et videte et admiramini et obstupescite quia opus factum est in diebus vestris quod nemo credet cum narrabitur
HAB|1|6|quia ecce ego suscitabo Chaldeos gentem amaram et velocem ambulantem super latitudinem terrae ut possideat tabernacula non sua
HAB|1|7|horribilis et terribilis est ex semet ipsa iudicium et onus eius egredietur
HAB|1|8|leviores pardis equi eius et velociores lupis vespertinis et diffundentur equites eius equites namque eius de longe venient volabunt quasi aquila festinans ad comedendum
HAB|1|9|omnes ad praedam venient facies eorum ventus urens et congregabit quasi harenam captivitatem
HAB|1|10|et ipse de regibus triumphabit et tyranni ridiculi eius erunt ipse super omnem munitionem ridebit et conportabit aggerem et capiet eam
HAB|1|11|tunc mutabitur spiritus et pertransibit et corruet haec est fortitudo eius dei sui
HAB|1|12|numquid non tu a principio Domine Deus meus Sancte meus et non moriemur Domine in iudicium posuisti eum et fortem ut corriperes fundasti eum
HAB|1|13|mundi sunt oculi tui ne videas malum et respicere ad iniquitatem non poteris quare non respicis super inique agentes et taces devorante impio iustiorem se
HAB|1|14|et facies homines quasi pisces maris et quasi reptile non habens principem
HAB|1|15|totum in hamo sublevavit traxit illud in sagena sua et congregavit in rete suo super hoc laetabitur et exultabit
HAB|1|16|propterea immolabit sagenae suae et sacrificabit reti suo quia in ipsis incrassata est pars eius et cibus eius electus
HAB|1|17|propter hoc ergo expandit sagenam suam et semper interficere gentes non parcet
HAB|2|1|super custodiam meam stabo et figam gradum super munitionem et contemplabor ut videam quid dicatur mihi et quid respondeam ad arguentem me
HAB|2|2|et respondit mihi Dominus et dixit scribe visum et explana eum super tabulas ut percurrat qui legerit eum
HAB|2|3|quia adhuc visus procul et apparebit in finem et non mentietur si moram fecerit expecta illum quia veniens veniet et non tardabit
HAB|2|4|ecce qui incredulus est non erit recta anima eius in semet ipso iustus autem in fide sua vivet
HAB|2|5|et quomodo vinum potantem decipit sic erit vir superbus et non decorabitur qui dilatavit quasi infernus animam suam et ipse quasi mors et non adimpletur et congregabit ad se omnes gentes et coacervabit ad se omnes populos
HAB|2|6|numquid non omnes isti super eum parabolam sument et loquellam enigmatum eius et dicetur vae ei qui multiplicat non sua usquequo et adgravat contra se densum lutum
HAB|2|7|numquid non repente consurgent qui mordeant te et suscitabuntur lacerantes te et eris in rapinam eis
HAB|2|8|quia tu spoliasti gentes multas spoliabunt te omnes qui reliqui fuerint de populis propter sanguinem hominis et iniquitatem terrae civitatis et omnium habitantium in ea
HAB|2|9|vae qui congregat avaritiam malam domui suae ut sit in excelso nidus eius et liberari se putat de manu mali
HAB|2|10|cogitasti confusionem domui tuae concidisti populos multos et peccavit anima tua
HAB|2|11|quia lapis de pariete clamabit et lignum quod inter iuncturas aedificiorum est respondebit
HAB|2|12|vae qui aedificat civitatem in sanguinibus et praeparat urbem in iniquitate
HAB|2|13|numquid non haec a Domino sunt exercituum laborabunt enim populi in multo igni et gentes in vacuum et deficient
HAB|2|14|quia replebitur terra ut cognoscat gloriam Domini quasi aquae operientes mare
HAB|2|15|vae qui potum dat amico suo mittens fel suum et inebrians ut aspiciat nuditatem eius
HAB|2|16|repletus est ignominia pro gloria bibe tu quoque et consopire circumdabit te calix dexterae Domini et vomitus ignominiae super gloriam tuam
HAB|2|17|quia iniquitas Libani operiet te et vastitas animalium deterrebit eos de sanguinibus hominis et iniquitate terrae et civitatis et omnium habitantium in ea
HAB|2|18|quid prodest sculptile quia sculpsit illud fictor suus conflatile et imaginem falsam quia speravit in figmento fictor eius ut faceret simulacra muta
HAB|2|19|vae qui dicit ligno expergiscere surge lapidi tacenti numquid ipse docere poterit ecce iste coopertus est auro et argento et omnis spiritus non est in visceribus eius
HAB|2|20|Dominus autem in templo sancto suo sileat a facie eius omnis terra
HAB|3|1|oratio Abacuc prophetae pro ignorationibus
HAB|3|2|Domine audivi auditionem tuam et timui Domine opus tuum in medio annorum vivifica illud in medio annorum notum facies cum iratus fueris misericordiae recordaberis
HAB|3|3|Deus ab austro veniet et Sanctus de monte Pharan semper operuit caelos gloria eius et laudis eius plena est terra
HAB|3|4|splendor eius ut lux erit cornua in manibus eius ibi abscondita est fortitudo eius
HAB|3|5|ante faciem eius ibit mors et egredietur diabolus ante pedes eius
HAB|3|6|stetit et mensus est terram aspexit et dissolvit gentes et contriti sunt montes saeculi incurvati sunt colles mundi ab itineribus aeternitatis eius
HAB|3|7|pro iniquitate vidi tentoria Aethiopiae turbabuntur pelles terrae Madian
HAB|3|8|numquid in fluminibus iratus es Domine aut in fluminibus furor tuus vel in mari indignatio tua quia ascendes super equos tuos et quadrigae tuae salvatio
HAB|3|9|suscitans suscitabis arcum tuum iuramenta tribubus quae locutus es semper fluvios scindes terrae
HAB|3|10|viderunt te et doluerunt montes gurges aquarum transiit dedit abyssus vocem suam altitudo manus suas levavit
HAB|3|11|sol et luna steterunt in habitaculo suo in luce sagittarum tuarum ibunt in splendore fulgurantis hastae tuae
HAB|3|12|in fremitu conculcabis terram in furore obstupefacies gentes
HAB|3|13|egressus es in salutem populi tui in salutem cum christo tuo percussisti caput de domo impii denudasti fundamentum usque ad collum semper
HAB|3|14|maledixisti sceptris eius capiti bellatorum eius venientibus ut turbo ad dispergendum me exultatio eorum sicut eius qui devorat pauperem in abscondito
HAB|3|15|viam fecisti in mari equis tuis in luto aquarum multarum
HAB|3|16|audivi et conturbatus est venter meus ad vocem contremuerunt labia mea ingrediatur putredo in ossibus meis et subter me scateat ut requiescam in die tribulationis ut ascendam ad populum accinctum nostrum
HAB|3|17|ficus enim non florebit et non erit germen in vineis mentietur opus olivae et arva non adferent cibum abscidetur de ovili pecus et non erit armentum in praesepibus
HAB|3|18|ego autem in Domino gaudebo exultabo in Deo Iesu meo
HAB|3|19|Dominus Deus fortitudo mea et ponet pedes meos quasi cervorum et super excelsa mea deducet me victori in psalmis canentem
ZEPH|1|1|verbum Domini quod factum est ad Sofoniam filium Chusi filium Godoliae filii Amariae filii Ezechiae in diebus Iosiae filii Amon regis Iuda
ZEPH|1|2|congregans congregabo omnia a facie terrae dicit Dominus
ZEPH|1|3|congregans hominem et pecus congregans volatile caeli et pisces maris et ruinae impiorum erunt et disperdam homines a facie terrae dicit Dominus
ZEPH|1|4|et extendam manum meam super Iudam et super omnes habitantes Hierusalem et disperdam de loco hoc reliquias Baal et nomina aedituorum cum sacerdotibus
ZEPH|1|5|et eos qui adorant super tecta militiam caeli et adorant et iurant in Domino et iurant in Melchom
ZEPH|1|6|et qui avertuntur de post tergum Domini et qui non quaesierunt Dominum nec investigaverunt eum
ZEPH|1|7|silete a facie Domini Dei quia iuxta est dies Domini quia praeparavit Dominus hostiam sanctificavit vocatos suos
ZEPH|1|8|et erit in die hostiae Domini visitabo super principes et super filios regis et super omnes qui induti sunt veste peregrina
ZEPH|1|9|et visitabo omnem qui arroganter ingreditur super limen in die illa qui conplent domum Domini Dei sui iniquitate et dolo
ZEPH|1|10|et erit in die illa dicit Dominus vox clamoris a porta Piscium et ululatus a secunda et contritio magna a collibus
ZEPH|1|11|ululate habitatores pilae conticuit omnis populus Chanaan disperierunt omnes involuti argento
ZEPH|1|12|et erit in tempore illo scrutabor Hierusalem in lucernis et visitabo super viros defixos in fecibus suis qui dicunt in cordibus suis non faciet bene Dominus et non faciet male
ZEPH|1|13|et erit fortitudo eorum in direptionem et domus eorum in desertum et aedificabunt domos et non habitabunt et plantabunt vineas et non bibent vinum earum
ZEPH|1|14|iuxta est dies Domini magnus iuxta et velox nimis vox diei Domini amara tribulabitur ibi fortis
ZEPH|1|15|dies irae dies illa dies tribulationis et angustiae dies calamitatis et miseriae dies tenebrarum et caliginis dies nebulae et turbinis
ZEPH|1|16|dies tubae et clangoris super civitates munitas et super angulos excelsos
ZEPH|1|17|et tribulabo homines et ambulabunt ut caeci quia Domino peccaverunt et effundetur sanguis eorum sicut humus et corpus eorum sicut stercora
ZEPH|1|18|sed et argentum eorum et aurum eorum non poterit liberare eos in die irae Domini in igne zeli eius devorabitur omnis terra quia consummationem cum festinatione faciet cunctis habitantibus terram
ZEPH|2|1|convenite congregamini gens non amabilis
ZEPH|2|2|priusquam pariat iussio quasi pulverem transeuntem diem antequam veniat super vos ira furoris Domini antequam veniat super vos dies furoris Domini
ZEPH|2|3|quaerite Dominum omnes mansueti terrae qui iudicium eius estis operati quaerite iustum quaerite mansuetum si quo modo abscondamini in die furoris Domini
ZEPH|2|4|quia Gaza destructa erit et Ascalon in desertum Azotum in meridie eicient et Accaron eradicabitur
ZEPH|2|5|vae qui habitatis funiculum maris gens perditorum verbum Domini super vos Chanaan terra Philisthinorum et disperdam te ita ut non sit inhabitator
ZEPH|2|6|et erit funiculus maris requies pastorum et caulae pecorum
ZEPH|2|7|et erit funiculus eius qui remanserit de domo Iuda ibi pascentur in domibus Ascalonis ad vesperam requiescent quia visitabit eos Dominus Deus eorum et avertet captivitatem eorum
ZEPH|2|8|audivi obprobrium Moab et blasphemias filiorum Ammon quae exprobraverunt populo meo et magnificati sunt super terminos eorum
ZEPH|2|9|propterea vivo ego dicit Dominus exercituum Deus Israhel quia Moab ut Sodoma erit et filii Ammon quasi Gomorra siccitas spinarum et acervi salis et desertum usque in aeternum reliquiae populi mei diripient illos residui gentis meae possidebunt eos
ZEPH|2|10|hoc eis eveniet pro superbia sua quia blasphemaverunt et magnificati sunt super populum Domini exercituum
ZEPH|2|11|horribilis Dominus super eos et adtenuabit omnes deos terrae et adorabunt eum vir de loco suo omnes insulae gentium
ZEPH|2|12|sed et vos Aethiopes interfecti gladio meo eritis
ZEPH|2|13|et extendet manum suam super aquilonem et perdet Assur et ponet speciosam in solitudinem et in invium et quasi desertum
ZEPH|2|14|et accubabunt in medio eius greges omnes bestiae gentium et onocrotalus et ericius in liminibus eius morabuntur vox cantantis in fenestra corvus in superliminari quoniam adtenuabo robur eius
ZEPH|2|15|haec est civitas gloriosa habitans in confidentia quae dicebat in corde suo ego sum et extra me non est alia amplius quomodo facta est in desertum cubile bestiae omnis qui transit per eam sibilabit et movebit manum suam
ZEPH|3|1|vae provocatrix et redempta civitas columba
ZEPH|3|2|non audivit vocem et non suscepit disciplinam in Domino non est confisa ad Deum suum non adpropiavit
ZEPH|3|3|principes eius in medio eius quasi leones rugientes iudices eius lupi vespere non relinquebant in mane
ZEPH|3|4|prophetae eius vesani viri infideles sacerdotes eius polluerunt sanctum iniuste egerunt contra legem
ZEPH|3|5|Dominus iustus in medio eius non faciet iniquitatem mane mane iudicium suum dabit in luce et non abscondetur nescivit autem iniquus confusionem
ZEPH|3|6|disperdi gentes et dissipati sunt anguli earum desertas feci vias eorum dum non est qui transeat desolatae sunt civitates eorum non remanente viro nec ullo habitatore
ZEPH|3|7|dixi attamen timebis me suscipies disciplinam et non peribit habitaculum eius propter omnia in quibus visitavi eam verumtamen diluculo surgentes corruperunt omnes cogitationes suas
ZEPH|3|8|quapropter expecta me dicit Dominus in die resurrectionis meae in futurum quia iudicium meum ut congregem gentes et colligam regna ut effundam super eas indignationem meam omnem iram furoris mei in igne enim zeli mei devorabitur omnis terra
ZEPH|3|9|quia tunc reddam populis labium electum ut vocent omnes in nomine Domini et serviant ei umero uno
ZEPH|3|10|ultra flumina Aethiopiae inde supplices mei filii dispersorum meorum deferent munus mihi
ZEPH|3|11|in die illa non confunderis super cunctis adinventionibus tuis quibus praevaricata es in me quia tunc auferam de medio tui magniloquos superbiae tuae et non adicies exaltari amplius in monte sancto meo
ZEPH|3|12|et derelinquam in medio tui populum pauperem et egenum et sperabunt in nomine Domini
ZEPH|3|13|reliquiae Israhel non facient iniquitatem nec loquentur mendacium et non invenietur in ore eorum lingua dolosa quoniam ipsi pascentur et accubabunt et non erit qui exterreat
ZEPH|3|14|lauda filia Sion iubilate Israhel laetare et exulta in omni corde filia Hierusalem
ZEPH|3|15|abstulit Dominus iudicium tuum avertit inimicos tuos rex Israhel Dominus in medio tui non timebis malum ultra
ZEPH|3|16|in die illa dicetur Hierusalem noli timere Sion non dissolvantur manus tuae
ZEPH|3|17|Dominus Deus tuus in medio tui Fortis ipse salvabit gaudebit super te in laetitia silebit in dilectione tua exultabit super te in laude
ZEPH|3|18|nugas qui a lege recesserant congregabo quia ex te erant ut non ultra habeas super eis obprobrium
ZEPH|3|19|ecce ego interficiam omnes qui adflixerunt te in tempore illo et salvabo claudicantem et eam quae eiecta fuerat congregabo et ponam eos in laudem et in nomen in omni terra confusionis eorum
ZEPH|3|20|in tempore illo quo adducam vos et in tempore quo congregabo vos dabo enim vos in nomen et in laudem omnibus populis terrae cum convertero captivitatem vestram coram oculis vestris dicit Dominus
HAG|1|1|in anno secundo Darii regis in mense sexto in die una mensis factum est verbum Domini in manu Aggei prophetae ad Zorobabel filium Salathihel ducem Iuda et ad Iesum filium Iosedech sacerdotem magnum dicens
HAG|1|2|haec ait Dominus exercituum dicens populus iste dicit nondum venit tempus domus Domini aedificandae
HAG|1|3|et factum est verbum Domini in manu Aggei prophetae dicens
HAG|1|4|numquid tempus vobis est ut habitetis in domibus laqueatis et domus ista deserta
HAG|1|5|et nunc haec dicit Dominus exercituum ponite corda vestra super vias vestras
HAG|1|6|seminastis multum et intulistis parum comedistis et non estis satiati bibistis et non estis inebriati operuistis vos et non estis calefacti et qui mercedes congregavit misit eas in sacculum pertusum
HAG|1|7|haec dicit Dominus exercituum ponite corda vestra super vias vestras
HAG|1|8|ascendite in montem portate lignum et aedificate domum et acceptabilis mihi erit et glorificabor dicit Dominus
HAG|1|9|respexistis ad amplius et ecce factum est minus et intulistis in domum et exsuflavi illud quam ob causam dicit Dominus exercituum quia domus mea deserta est et vos festinatis unusquisque in domum suam
HAG|1|10|propter hoc super vos prohibiti sunt caeli ne darent rorem et terra prohibita est ne daret germen suum
HAG|1|11|et vocavi siccitatem super terram et super montes et super triticum et super vinum et super oleum et quaecumque profert humus et super homines et super iumenta et super omnem laborem manuum
HAG|1|12|et audivit Zorobabel filius Salathihel et Iesus filius Iosedech sacerdos magnus et omnes reliquiae populi vocem Dei sui et verba Aggei prophetae sicut misit eum Dominus Deus eorum ad ipsos et timuit populus a facie Domini
HAG|1|13|et dixit Aggeus nuntius Domini de nuntiis Domini populo dicens ego vobiscum dicit Dominus
HAG|1|14|et suscitavit Dominus spiritum Zorobabel filii Salathihel ducis Iuda et spiritum Iesu filii Iosedech sacerdotis magni et spiritum reliquorum de omni populo et ingressi sunt et faciebant opus in domo Domini exercituum Dei sui
HAG|2|1|in die vicesima et quarta mensis in sexto mense in anno secundo Darii regis
HAG|2|2|in septimo mense vicesima et prima mensis factum est verbum Domini in manu Aggei prophetae dicens
HAG|2|3|loquere ad Zorobabel filium Salathihel ducem Iuda et ad Iesum filium Iosedech sacerdotem magnum et ad reliquos populi dicens
HAG|2|4|quis in vobis est derelictus qui vidit domum istam in gloria sua prima et quid vos videtis hanc nunc numquid non ita est quasi non sit in oculis vestris
HAG|2|5|et nunc confortare Zorobabel dicit Dominus et confortare Iesu fili Iosedech sacerdos magne et confortare omnis popule terrae dicit Dominus exercituum et facite quoniam ego vobiscum sum dicit Dominus exercituum
HAG|2|6|verbum quod placui vobiscum cum egrederemini de terra Aegypti et spiritus meus erit in medio vestrum nolite timere
HAG|2|7|quia haec dicit Dominus exercituum adhuc unum modicum est et ego commovebo caelum et terram et mare et aridam
HAG|2|8|et movebo omnes gentes et veniet desideratus cunctis gentibus et implebo domum istam gloria dicit Dominus exercituum
HAG|2|9|meum est argentum et meum est aurum dicit Dominus exercituum
HAG|2|10|magna erit gloria domus istius novissimae plus quam primae dicit Dominus exercituum et in loco isto dabo pacem dicit Dominus exercituum
HAG|2|11|in vicesima et quarta noni mensis in anno secundo Darii factum est verbum Domini ad Aggeum prophetam dicens
HAG|2|12|haec dicit Dominus exercituum interroga sacerdotes legem dicens
HAG|2|13|si tulerit homo carnem sanctificatam in ora vestimenti sui et tetigerit de summitate eius panem aut pulmentum aut vinum aut oleum aut omnem cibum numquid sanctificabitur respondentes autem sacerdotes dixerunt non
HAG|2|14|et dixit Aggeus si tetigerit pollutus in anima ex omnibus his numquid contaminabitur et responderunt sacerdotes et dixerunt contaminabitur
HAG|2|15|et respondit Aggeus et dixit sic populus iste et sic gens ista ante faciem meam dicit Dominus et sic omne opus manuum eorum et omnia quae obtulerint ibi contaminata erunt
HAG|2|16|et nunc ponite corda vestra a die hac et supra antequam poneretur lapis super lapidem in templo Domini
HAG|2|17|cum accederetis ad acervum viginti modiorum et fierent decem intraretis ad torcular ut exprimeretis quinquaginta lagoenas et fiebant viginti
HAG|2|18|percussi vos vento urente et aurugine et grandine omnia opera manuum vestrarum et non fuit in vobis qui reverteretur ad me dicit Dominus
HAG|2|19|ponite corda vestra ex die ista et in futurum a die vicesima et quarta noni mensis a die qua fundamenta iacta sunt templi Domini ponite super cor vestrum
HAG|2|20|numquid iam semen in germine est et adhuc vinea et ficus et malogranatum et lignum olivae non floruit ex die ista benedicam
HAG|2|21|et factum est verbum Domini secundo ad Aggeum in vicesima et quarta mensis dicens
HAG|2|22|loquere ad Zorobabel ducem Iuda dicens ego movebo caelum pariter et terram
HAG|2|23|et subvertam solium regnorum et conteram fortitudinem regni gentium et subvertam quadrigam et ascensorem eius et descendent equi et ascensores eorum vir in gladio fratris sui
HAG|2|24|in die illo dicit Dominus exercituum adsumam te Zorobabel fili Salathihel serve meus dicit Dominus et ponam te quasi signaculum quia te elegi dicit Dominus exercituum
ZECH|1|1|in mense octavo in anno secundo Darii factum est verbum Domini ad Zacchariam filium Barachiae filium Addo prophetam dicens
ZECH|1|2|iratus est Dominus super patres vestros iracundia
ZECH|1|3|et dices ad eos haec dicit Dominus exercituum convertimini ad me ait Dominus exercituum et convertar ad vos dicit Dominus exercituum
ZECH|1|4|ne sitis sicut patres vestri ad quos clamabant prophetae priores dicentes haec dicit Dominus exercituum convertimini de viis vestris malis et cogitationibus vestris pessimis et non audierunt neque adtenderunt ad me dicit Dominus
ZECH|1|5|patres vestri ubi sunt et prophetae numquid in sempiternum vivent
ZECH|1|6|verumtamen verba mea et legitima mea quae mandavi servis meis prophetis numquid non conprehenderunt patres vestros et conversi sunt et dixerunt sicut cogitavit Dominus exercituum facere nobis secundum vias nostras et secundum adinventiones nostras fecit nobis
ZECH|1|7|in die vicesima et quarta undecimo mense sabath in anno secundo Darii factum est verbum Domini ad Zacchariam filium Barachiae filium Addo prophetam dicens
ZECH|1|8|vidi per noctem et ecce vir ascendens super equum rufum et ipse stabat inter myrteta quae erant in profundo et post eum equi rufi varii et albi
ZECH|1|9|et dixi quid sunt isti domine mi et dixit ad me angelus qui loquebatur in me ego ostendam tibi quid sint haec
ZECH|1|10|et respondit vir qui stabat inter myrteta et dixit isti sunt quos misit Dominus ut perambularent terram
ZECH|1|11|et responderunt angelo Domini qui stabat inter myrteta et dixerunt perambulavimus terram et ecce omnis terra habitatur et quiescit
ZECH|1|12|et respondit angelus Domini et dixit Domine exercituum usquequo tu non misereberis Hierusalem et urbium Iuda quibus iratus es iste septuagesimus annus est
ZECH|1|13|et respondit Dominus angelo qui loquebatur in me verba bona verba consolatoria
ZECH|1|14|et dixit ad me angelus qui loquebatur in me clama dicens haec dicit Dominus exercituum zelatus sum Hierusalem et Sion zelo magno
ZECH|1|15|et ira magna ego irascor super gentes opulentas quia ego iratus sum parum ipsi vero adiuverunt in malum
ZECH|1|16|propterea haec dicit Dominus revertar ad Hierusalem in misericordiis domus mea aedificabitur in ea ait Dominus exercituum et perpendiculum extendetur super Hierusalem
ZECH|1|17|adhuc clama dicens haec dicit Dominus exercituum adhuc affluent civitates meae bonis et consolabitur Dominus adhuc Sion et eliget adhuc Hierusalem
ZECH|1|18|et levavi oculos meos et vidi et ecce quattuor cornua
ZECH|1|19|et dixi ad angelum qui loquebatur in me quid sunt haec et dixit ad me haec sunt cornua quae ventilaverunt Iudam et Israhel et Hierusalem
ZECH|1|20|et ostendit mihi Dominus quattuor fabros
ZECH|1|21|et dixi quid isti veniunt facere qui ait dicens haec sunt cornua quae ventilaverunt Iudam per singulos viros et nemo eorum levavit caput suum et venerunt isti deterrere ea ut deiciant cornua gentium quae levaverunt cornu super terram Iuda ut dispergerent eam
ZECH|2|1|et levavi oculos meos et vidi et ecce vir et in manu eius funiculus mensorum
ZECH|2|2|et dixi quo tu vadis et dixit ad me ut metiar Hierusalem et videam quanta sit latitudo eius et quanta longitudo eius
ZECH|2|3|et ecce angelus qui loquebatur in me egrediebatur et angelus alius egrediebatur in occursum eius
ZECH|2|4|et dixit ad eum curre loquere ad puerum istum dicens absque muro habitabitur Hierusalem prae multitudine hominum et iumentorum in medio eius
ZECH|2|5|et ego ero ei ait Dominus murus ignis in circuitu et in gloria ero in medio eius
ZECH|2|6|o o fugite de terra aquilonis dicit Dominus quoniam in quattuor ventos caeli dispersi vos dicit Dominus
ZECH|2|7|o Sion fuge quae habitas apud filiam Babylonis
ZECH|2|8|quia haec dicit Dominus exercituum post gloriam misit me ad gentes quae spoliaverunt vos qui enim tetigerit vos tangit pupillam oculi eius
ZECH|2|9|quia ecce ego levo manum meam super eos et erunt praedae his qui serviebant sibi et cognoscetis quia Dominus exercituum misit me
ZECH|2|10|lauda et laetare filia Sion quia ecce ego venio et habitabo in medio tui ait Dominus
ZECH|2|11|et adplicabuntur gentes multae ad Dominum in die illa et erunt mihi in populum et habitabo in medio tui et scies quia Dominus exercituum misit me ad te
ZECH|2|12|et possidebit Dominus Iudam partem suam in terra sanctificata et eliget adhuc Hierusalem
ZECH|2|13|sileat omnis caro a facie Domini quia consurrexit de habitaculo sancto suo
ZECH|3|1|et ostendit mihi Iesum sacerdotem magnum stantem coram angelo Domini et Satan stabat a dextris eius ut adversaretur ei
ZECH|3|2|et dixit Dominus ad Satan increpet Dominus in te Satan et increpet Dominus in te qui elegit Hierusalem numquid non iste torris est erutus de igne
ZECH|3|3|et Iesus erat indutus vestibus sordidis et stabat ante faciem angeli
ZECH|3|4|qui respondit et ait ad eos qui stabant coram se dicens auferte vestimenta sordida ab eo et dixit ad eum ecce abstuli a te iniquitatem tuam et indui te mutatoriis
ZECH|3|5|et dixit ponite cidarim mundam super caput eius et posuerunt cidarim mundam super caput eius et induerunt eum vestibus et angelus Domini stabat
ZECH|3|6|et contestabatur angelus Domini Iesum dicens
ZECH|3|7|haec dicit Dominus exercituum si in viis meis ambulaveris et custodiam meam custodieris tu quoque iudicabis domum meam et custodies atria mea et dabo tibi ambulantes de his qui nunc hic adsistunt
ZECH|3|8|audi Iesu sacerdos magne tu et amici tui qui habitant coram te quia viri portendentes sunt ecce enim ego adducam servum meum orientem
ZECH|3|9|quia ecce lapis quem dedi coram Iesu super lapidem unum septem oculi sunt ecce ego celabo sculpturam eius ait Dominus exercituum et auferam iniquitatem terrae illius in die una
ZECH|3|10|in die illa dicit Dominus exercituum vocabit vir amicum suum subter vineam et subter ficum
ZECH|4|1|et reversus est angelus qui loquebatur in me et suscitavit me quasi virum qui suscitatur de somno suo
ZECH|4|2|et dixit ad me quid tu vides et dixi vidi et ecce candelabrum aureum totum et lampas eius super caput ipsius et septem lucernae eius super illud septem et septem infusoria lucernis quae erant super caput illius
ZECH|4|3|et duae olivae super illud una a dextris lampadis et una a sinistris eius
ZECH|4|4|et respondi et aio ad angelum qui loquebatur in me dicens quid sunt haec domine mi
ZECH|4|5|et respondit angelus qui loquebatur in me et dixit ad me numquid nescis quid sunt haec et dixi non domine mi
ZECH|4|6|et respondit et ait ad me dicens hoc est verbum Domini ad Zorobabel dicens non in exercitu nec in robore sed in spiritu meo dicit Dominus exercituum
ZECH|4|7|quis tu mons magne coram Zorobabel in planum et educet lapidem primarium et exaequabit gratiam gratiae eius
ZECH|4|8|et factum est verbum Domini ad me dicens
ZECH|4|9|manus Zorobabel fundaverunt domum istam et manus eius perficient eam et scietis quia Dominus exercituum misit me ad vos
ZECH|4|10|quis enim despexit dies parvos et laetabuntur et videbunt lapidem stagneum in manu Zorobabel septem isti oculi Domini qui discurrunt in universa terra
ZECH|4|11|et respondi et dixi ad eum quid sunt duae olivae istae ad dextram candelabri et ad sinistram eius
ZECH|4|12|et respondi secundo et dixi ad eum quid sunt duae spicae olivarum quae sunt iuxta duo rostra aurea in quibus sunt suffusoria ex auro
ZECH|4|13|et ait ad me dicens numquid nescis quid sunt haec et dixi non domine
ZECH|4|14|et dixit isti duo filii olei qui adsistunt Dominatori universae terrae
ZECH|5|1|et conversus sum et levavi oculos meos et vidi et ecce volumen volans
ZECH|5|2|et dixit ad me quid tu vides et dixi ego video volumen volans longitudo eius viginti cubitorum et latitudo eius decem cubitorum
ZECH|5|3|et dixit ad me haec est maledictio quae egreditur super faciem omnis terrae quia omnis fur sicut ibi scriptum est iudicabitur et omnis iurans ex hoc similiter iudicabitur
ZECH|5|4|educam illud dicit Dominus exercituum et veniet ad domum furis et ad domum iurantis in nomine meo mendaciter et commorabitur in medio domus eius et consumet eam et ligna eius et lapides eius
ZECH|5|5|et egressus est angelus qui loquebatur in me et dixit ad me leva oculos tuos et vide quid est hoc quod egreditur
ZECH|5|6|et dixi quidnam est et ait haec est amphora egrediens et dixit haec est oculus eorum in universa terra
ZECH|5|7|et ecce talentum plumbi portabatur et ecce mulier una sedens in medio amphorae
ZECH|5|8|et dixit haec est impietas et proiecit eam in medio amphorae et misit massam plumbeam in os eius
ZECH|5|9|et levavi oculos meos et vidi et ecce duae mulieres egredientes et spiritus in alis earum et habebant alas quasi alas milvi et levaverunt amphoram inter terram et caelum
ZECH|5|10|et dixi ad angelum qui loquebatur in me quo istae deferunt amphoram
ZECH|5|11|et dixit ad me ut aedificetur ei domus in terra Sennaar et stabiliatur et ponatur ibi super basem suam
ZECH|6|1|et conversus sum et levavi oculos meos et vidi et ecce quattuor quadrigae egredientes de medio duorum montium et montes montes aerei
ZECH|6|2|in quadriga prima equi rufi et in quadriga secunda equi nigri
ZECH|6|3|et in quadriga tertia equi albi et in quadriga quarta equi varii fortes
ZECH|6|4|et respondi et dixi ad angelum qui loquebatur in me quid sunt haec domine mi
ZECH|6|5|et respondit angelus et ait ad me isti sunt quattuor venti caeli qui egrediuntur ut stent coram Dominatore omnis terrae
ZECH|6|6|in quo erant equi nigri egrediebantur in terra aquilonis et albi egressi sunt post eos et varii egressi sunt ad terram austri
ZECH|6|7|qui autem erant robustissimi exierunt et quaerebant ire et discurrere per omnem terram et dixit ite perambulate terram et perambulaverunt terram
ZECH|6|8|et vocavit me et locutus est ad me dicens ecce qui egrediuntur in terram aquilonis requiescere fecerunt spiritum meum in terra aquilonis
ZECH|6|9|et factum est verbum Domini ad me dicens
ZECH|6|10|sume a transmigratione ab Oldai et a Tobia et ab Idaia et venies tu in die illa et intrabis domum Iosiae filii Sofoniae qui venerunt de Babylone
ZECH|6|11|et sumes argentum et aurum et facies coronas et pones in capite Iesu filii Iosedech sacerdotis magni
ZECH|6|12|et loqueris ad eum dicens haec ait Dominus exercituum dicens ecce vir Oriens nomen eius et subter eum orietur et aedificabit templum Domino
ZECH|6|13|et ipse extruet templum Domino et ipse portabit gloriam et sedebit et dominabitur super solio suo et erit sacerdos super solio suo et consilium pacis erit inter duos illos
ZECH|6|14|et coronae erunt Helem et Tobiae et Idaiae et Hen filio Sofoniae memoriale in templo Domini
ZECH|6|15|et qui procul sunt venient et aedificabunt in templo Domini et scietis quia Dominus exercituum misit me ad vos erit autem hoc si auditu audieritis vocem Domini Dei vestri
ZECH|7|1|et factum est in anno quarto Darii regis factum est verbum Domini ad Zacchariam in quarta mensis noni qui est casleu
ZECH|7|2|et miserunt ad domum Dei Sarasar et Rogomelech et viri qui erant cum eo ad deprecandam faciem Domini
ZECH|7|3|ut dicerent sacerdotibus domus Domini exercituum et prophetis loquentes numquid flendum mihi est in mense quinto vel sanctificare me debeo sicuti feci iam multis annis
ZECH|7|4|et factum est verbum Domini exercituum ad me dicens
ZECH|7|5|loquere ad omnem populum terrae et ad sacerdotes dicens cum ieiunaretis et plangeretis in quinto et septimo per hos septuaginta annos numquid ieiunium ieiunastis mihi
ZECH|7|6|et cum comedistis et cum bibistis numquid non vobis comedistis et vobismet ipsis bibistis
ZECH|7|7|numquid non sunt verba quae locutus est Dominus in manu prophetarum priorum cum adhuc Hierusalem habitaretur et esset opulenta ipsa et urbes in circuitu eius et ad austrum et in campestribus habitaretur
ZECH|7|8|et factum est verbum Domini ad Zacchariam dicens
ZECH|7|9|haec ait Dominus exercituum dicens iudicium verum iudicate et misericordiam et miserationes facite unusquisque cum fratre suo
ZECH|7|10|et viduam et pupillum et advenam et pauperem nolite calumniari et malum vir fratri suo non cogitet in corde suo
ZECH|7|11|et noluerunt adtendere et verterunt scapulam recedentem et aures suas adgravaverunt ne audirent
ZECH|7|12|et cor suum posuerunt adamantem ne audirent legem et verba quae misit Dominus exercituum in spiritu suo per manum prophetarum priorum et facta est indignatio magna a Domino exercituum
ZECH|7|13|et factum est sicut locutus est et non audierunt sic clamabunt et non exaudiam dicit Dominus exercituum
ZECH|7|14|et dispersi eos per omnia regna quae nesciunt et terra desolata est ab eis eo quod non esset transiens et revertens et posuerunt terram desiderabilem in desertum
ZECH|8|1|et factum est verbum Domini exercituum dicens
ZECH|8|2|haec dicit Dominus exercituum zelatus sum Sion zelo magno et indignatione magna zelatus sum eam
ZECH|8|3|haec dicit Dominus exercituum reversus sum ad Sion et habitabo in medio Hierusalem et vocabitur Hierusalem civitas veritatis et mons Domini exercituum mons sanctificatus
ZECH|8|4|haec dicit Dominus exercituum adhuc habitabunt senes et anus in plateis Hierusalem et viri baculus in manu eius prae multitudine dierum
ZECH|8|5|et plateae civitatis conplebuntur infantibus et puellis ludentibus in plateis eius
ZECH|8|6|haec dicit Dominus exercituum si difficile videbitur in oculis reliquiarum populi huius in diebus illis numquid in oculis meis difficile erit dicit Dominus exercituum
ZECH|8|7|haec dicit Dominus exercituum ecce ego salvabo populum meum de terra orientis et de terra occasus solis
ZECH|8|8|et adducam eos et habitabunt in medio Hierusalem et erunt mihi in populum et ego ero eis in Deum in veritate et iustitia
ZECH|8|9|haec dicit Dominus exercituum confortentur manus vestrae qui auditis in diebus his sermones istos per os prophetarum in die qua fundata est domus Domini exercituum ut templum aedificaretur
ZECH|8|10|siquidem ante dies illos merces hominum non erat nec merces iumentorum erat neque introeunti et exeunti erat pax prae tribulatione et dimisi omnes homines unumquemque contra proximum suum
ZECH|8|11|nunc autem non iuxta dies priores ego faciam reliquiis populi huius dicit Dominus exercituum
ZECH|8|12|sed semen pacis erit vinea dabit fructum suum et terra dabit germen suum et caeli dabunt rorem suum et possidere faciam reliquias populi huius universa haec
ZECH|8|13|et erit sicut eratis maledictio in gentibus domus Iuda et domus Israhel sic salvabo vos et eritis benedictio nolite timere confortentur manus vestrae
ZECH|8|14|quia haec dicit Dominus exercituum sicut cogitavi ut adfligerem vos cum ad iracundiam provocassent patres vestri me dicit Dominus
ZECH|8|15|et non sum misertus sic conversus cogitavi in diebus istis ut benefaciam Hierusalem et domui Iuda nolite timere
ZECH|8|16|haec sunt ergo verba quae facietis loquimini veritatem unusquisque cum proximo suo veritatem et iudicium pacis iudicate in portis vestris
ZECH|8|17|et unusquisque malum contra amicum suum ne cogitetis in cordibus vestris et iuramentum mendax ne diligatis omnia enim haec sunt quae odi dicit Dominus
ZECH|8|18|et factum est verbum Domini exercituum ad me dicens
ZECH|8|19|haec dicit Dominus exercituum ieiunium quarti et ieiunium quinti et ieiunium septimi et ieiunium decimi erit domui Iuda in gaudium et in laetitiam et in sollemnitates praeclaras veritatem tantum et pacem diligite
ZECH|8|20|haec dicit Dominus exercituum usquequo veniant populi et habitent in civitatibus multis
ZECH|8|21|et vadant habitatores unus ad alterum dicentes eamus et deprecemur faciem Domini et quaeramus Dominum exercituum vadam etiam ego
ZECH|8|22|et venient populi multi et gentes robustae ad quaerendum Dominum exercituum in Hierusalem et deprecandam faciem Domini
ZECH|8|23|haec dicit Dominus exercituum in diebus illis in quibus adprehendent decem homines ex omnibus linguis gentium et adprehendent fimbriam viri iudaei dicentes ibimus vobiscum audivimus enim quoniam Deus vobiscum est
ZECH|9|1|onus verbi Domini in terra Adrach et Damasci requiei eius quia Domini est oculus hominis et omnium tribuum Israhel
ZECH|9|2|Emath quoque in terminis eius et Tyrus et Sidon adsumpserunt quippe sibi sapientiam valde
ZECH|9|3|et aedificavit Tyrus munitionem suam et coacervavit argentum quasi humum et aurum ut lutum platearum
ZECH|9|4|ecce Dominus possidebit eam et percutiet in mari fortitudinem eius et haec igni devorabitur
ZECH|9|5|videbit Ascalon et timebit et Gaza et dolebit nimis et Accaron quoniam confusa est spes eius et peribit rex de Gaza et Ascalon non habitabitur
ZECH|9|6|et sedebit separator in Azoto et disperdam superbiam Philisthinorum
ZECH|9|7|et auferam sanguinem eius de ore eius et abominationes eius de medio dentium eius et relinquetur etiam ipse Deo nostro et erit quasi dux in Iuda et Accaron quasi Iebuseus
ZECH|9|8|et circumdabo domum meam ex his qui militant mihi euntes et revertentes et non transibit super eos ultra exactor quia nunc vidi in oculis meis
ZECH|9|9|exulta satis filia Sion iubila filia Hierusalem ecce rex tuus veniet tibi iustus et salvator ipse pauper et ascendens super asinum et super pullum filium asinae
ZECH|9|10|et disperdam quadrigam ex Ephraim et equum de Hierusalem et dissipabitur arcus belli et loquetur pacem gentibus et potestas eius a mari usque ad mare et a fluminibus usque ad fines terrae
ZECH|9|11|tu quoque in sanguine testamenti tui emisisti vinctos tuos de lacu in quo non est aqua
ZECH|9|12|convertimini ad munitionem vincti spei hodie quoque adnuntians duplicia reddam tibi
ZECH|9|13|quoniam extendi mihi Iudam quasi arcum implevi Ephraim et suscitabo filios tuos Sion super filios tuos Graecia et ponam te quasi gladium fortium
ZECH|9|14|et Dominus Deus super eos videbitur et exibit ut fulgur iaculum eius et Dominus Deus in tuba canet et vadet in turbine austri
ZECH|9|15|Dominus exercituum proteget eos et devorabunt et subicient lapidibus fundae et bibentes inebriabuntur quasi vino et replebuntur ut fialae et quasi cornua altaris
ZECH|9|16|et salvabit eos Dominus Deus eorum in die illa ut gregem populi sui quia lapides sancti elevantur super terram eius
ZECH|9|17|quid enim bonum eius est et quid pulchrum eius nisi frumentum electorum et vinum germinans virgines
ZECH|10|1|petite a Domino pluviam in tempore serotino et Dominus faciet nives et pluviam imbris dabit eis singulis herbam in agro
ZECH|10|2|quia simulacra locuta sunt inutile et divini viderunt mendacium et somniatores frustra locuti sunt vane consolabantur idcirco abducti sunt quasi grex adfligentur quia non est eis pastor
ZECH|10|3|super pastores iratus est furor meus et super hircos visitabo quia visitavit Dominus exercituum gregem suum domum Iuda et posuit eos quasi equum gloriae suae in bello
ZECH|10|4|ex ipso angulus ex ipso paxillus ex ipso arcus proelii ex ipso egredietur omnis exactor simul
ZECH|10|5|et erunt quasi fortes conculcantes lutum viarum in proelio et bellabunt quia Dominus cum eis et confundentur ascensores equorum
ZECH|10|6|et confortabo domum Iuda et domum Ioseph salvabo et convertam eos quia miserebor eorum et erunt sicut fuerunt quando non proieceram eos ego enim Dominus Deus eorum et exaudiam eos
ZECH|10|7|et erunt quasi fortes Ephraim et laetabitur cor eorum quasi a vino et filii eorum videbunt et laetabuntur et exultabit cor eorum in Domino
ZECH|10|8|sibilabo eis et congregabo illos quia redemi eos et multiplicabo eos sicut ante fuerant multiplicati
ZECH|10|9|et seminabo eos in populis et de longe recordabuntur mei et vivent cum filiis suis et revertentur
ZECH|10|10|et reducam eos de terra Aegypti et de Assyriis congregabo eos et ad terram Galaad et Libani adducam eos et non invenietur eis locus
ZECH|10|11|et transibit in maris freto et percutiet in mari fluctus et confundentur omnia profunda Fluminis et humiliabitur superbia Assur et sceptrum Aegypti recedet
ZECH|10|12|confortabo eos in Domino et in nomine eius ambulabunt dicit Dominus
ZECH|11|1|aperi Libane portas tuas et comedat ignis cedros tuas
ZECH|11|2|ulula abies quia cecidit cedrus quoniam magnifici vastati sunt ululate quercus Basan quoniam succisus est saltus munitus
ZECH|11|3|vox ululatus pastorum quia vastata est magnificentia eorum vox rugitus leonum quoniam vastata est superbia Iordanis
ZECH|11|4|haec dicit Dominus Deus meus pasce pecora occisionis
ZECH|11|5|quae qui possederant occidebant et non dolebant et vendebant ea dicentes benedictus Dominus divites facti sumus et pastores eorum non parcebant eis
ZECH|11|6|et ego non parcam ultra super habitantes terram dicit Dominus ecce ego tradam homines unumquemque in manu proximi sui et in manu regis sui et concident terram et non eruam de manu eorum
ZECH|11|7|et pascam pecus occisionis propter hoc o pauperes gregis et adsumpsi mihi duas virgas unam vocavi Decorem et alteram vocavi Funiculos et pavi gregem
ZECH|11|8|et succidi tres pastores in mense uno et contracta est anima mea in eis siquidem anima eorum variavit in me
ZECH|11|9|et dixi non pascam vos quod moritur moriatur et quod succiditur succidatur et reliqui vorent unusquisque carnem proximi sui
ZECH|11|10|et tuli virgam meam quae vocabatur Decus et abscidi eam ut irritum facerem foedus meum quod percussi cum omnibus populis
ZECH|11|11|et in irritum deductum est in die illa et cognoverunt sic pauperes gregis qui custodiunt mihi quia verbum Domini est
ZECH|11|12|et dixi ad eos si bonum est in oculis vestris adferte mercedem meam et si non quiescite et adpenderunt mercedem meam triginta argenteos
ZECH|11|13|et dixit Dominus ad me proice illud ad statuarium decorum pretium quod adpretiatus sum ab eis et tuli triginta argenteos et proieci illos in domo Domini ad statuarium
ZECH|11|14|et praecidi virgam meam secundam quae appellabatur Funiculus ut dissolverem germanitatem inter Iudam et inter Israhel
ZECH|11|15|et dixit Dominus ad me adhuc sume tibi vasa pastoris stulti
ZECH|11|16|quia ecce ego suscitabo pastorem in terra qui derelicta non visitabit dispersum non quaeret et contritum non sanabit et id quod stat non enutriet et carnes pinguium comedet et ungulas eorum dissolvet
ZECH|11|17|o pastor et idolum derelinquens gregem gladius super brachium eius et super oculum dextrum eius brachium eius ariditate siccabitur et oculus dexter eius tenebrescens obscurabitur
ZECH|12|1|onus verbi Domini super Israhel dixit Dominus extendens caelum et fundans terram et fingens spiritum hominis in eo
ZECH|12|2|ecce ego ponam Hierusalem superliminare crapulae omnibus populis in circuitu sed et Iuda erit in obsidione contra Hierusalem
ZECH|12|3|et erit in die illa ponam Hierusalem lapidem oneris cunctis populis omnes qui levabunt eam concisione lacerabuntur et colligentur adversum eam omnia regna terrae
ZECH|12|4|in die illa dicit Dominus percutiam omnem equum in stuporem et ascensorem eius in amentiam et super domum Iuda aperiam oculos meos et omnem equum populorum percutiam in caecitate
ZECH|12|5|et dicent duces Iuda in corde suo confortentur mihi habitatores Hierusalem in Domino exercituum Deo eorum
ZECH|12|6|in die illo ponam duces Iuda sicut caminum ignis in lignis et sicut facem ignis in faeno et devorabunt ad dextram et ad sinistram omnes populos in circuitu et habitabitur Hierusalem rursum in loco suo in Hierusalem
ZECH|12|7|et salvabit Dominus tabernacula Iuda sicut in principio ut non magnifice glorietur domus David et gloria habitantium Hierusalem contra Iudam
ZECH|12|8|in die illo proteget Dominus habitatores Hierusalem et erit qui offenderit ex eis in die illa quasi David et domus David quasi Dei sicut angelus Domini in conspectu eius
ZECH|12|9|et erit in die illa quaeram conterere omnes gentes quae veniunt contra Hierusalem
ZECH|12|10|et effundam super domum David et super habitatores Hierusalem spiritum gratiae et precum et aspicient ad me quem confixerunt et plangent eum planctu quasi super unigenitum et dolebunt super eum ut doleri solet in morte primogeniti
ZECH|12|11|in die illa magnus erit planctus in Hierusalem sicut planctus Adadremmon in campo Mageddon
ZECH|12|12|et planget terra familiae et familiae seorsum familiae domus David seorsum et mulieres eorum seorsum
ZECH|12|13|familiae domus Nathan seorsum et mulieres eorum seorsum familiae domus Levi seorsum et mulieres eorum seorsum familiae Semei seorsum et mulieres eorum seorsum
ZECH|12|14|omnes familiae reliquae familiae et familiae seorsum et mulieres eorum seorsum
ZECH|13|1|in die illa erit fons patens domus David et habitantibus Hierusalem in ablutionem peccatoris et menstruatae
ZECH|13|2|et erit in die illa dicit Dominus exercituum disperdam nomina idolorum de terra et non memorabuntur ultra et prophetas et spiritum inmundum auferam de terra
ZECH|13|3|et erit cum prophetaverit quispiam ultra dicent ei pater eius et mater eius qui genuerunt eum non vives quia mendacium locutus es in nomine Domini et configent eum pater eius et mater eius genitores eius cum prophetaverit
ZECH|13|4|et erit in die illa confundentur prophetae unusquisque ex visione sua cum prophetaverit nec operientur pallio saccino ut mentiantur
ZECH|13|5|sed dicet non sum propheta homo agricola ego sum quoniam Adam exemplum meum ab adulescentia mea
ZECH|13|6|et dicetur ei quid sunt plagae istae in medio manuum tuarum et dicet his plagatus sum in domo eorum qui diligebant me
ZECH|13|7|framea suscitare super pastorem meum et super virum coherentem mihi dicit Dominus exercituum percute pastorem et dispergantur oves et convertam manum meam ad parvulos
ZECH|13|8|et erunt in omni terra dicit Dominus partes duae in ea disperdentur et deficient et tertia pars relinquetur in ea
ZECH|13|9|et ducam tertiam partem per ignem et uram eas sicut uritur argentum et probabo eos sicut probatur aurum ipse vocabit nomen meum et ego exaudiam eum dicam populus meus es et ipse dicet Dominus Deus meus
ZECH|14|1|ecce dies veniunt Domini et dividentur spolia tua in medio tui
ZECH|14|2|et congregabo omnes gentes ad Hierusalem in proelium et capietur civitas et vastabuntur domus et mulieres violabuntur et egredietur media pars civitatis in captivitatem et reliquum populi non auferetur ex urbe
ZECH|14|3|et egredietur Dominus et proeliabitur contra gentes illas sicut proeliatus est in die certaminis
ZECH|14|4|et stabunt pedes eius in die illa super montem Olivarum qui est contra Hierusalem ad orientem et scindetur mons Olivarum ex media parte sui ad orientem et occidentem praerupto grandi valde et separabitur medium montis ad aquilonem et medium eius ad meridiem
ZECH|14|5|et fugietis ad vallem montium meorum quoniam coniungetur vallis montium usque ad proximum et fugietis sicut fugistis a facie terraemotus in diebus Oziae regis Iuda et veniet Dominus Deus meus omnesque sancti cum eo
ZECH|14|6|et erit in die illa non erit lux sed frigus et gelu
ZECH|14|7|et erit dies una quae nota est Domino non dies neque nox et in tempore vesperae erit lux
ZECH|14|8|et erit in die illa exibunt aquae vivae de Hierusalem medium earum ad mare orientale et medium earum ad mare novissimum in aestate et in hieme erunt
ZECH|14|9|et erit Dominus rex super omnem terram in die illa erit Dominus unus et erit nomen eius unum
ZECH|14|10|et revertetur omnis terra usque ad desertum de colle Remmon ad austrum Hierusalem et exaltabitur et habitabit in loco suo a porta Beniamin usque ad locum portae Prioris usque ad portam Angulorum et a turre Ananehel usque ad torcularia regis
ZECH|14|11|et habitabunt in ea et anathema non erit amplius sed sedebit Hierusalem secura
ZECH|14|12|et haec erit plaga qua percutiet Dominus omnes gentes quae pugnaverunt adversus Hierusalem tabescet caro uniuscuiusque stantis super pedes suos et oculi eius contabescent in foraminibus suis et lingua eorum contabescet in ore suo
ZECH|14|13|in die illo erit tumultus Domini magnus in eis et adprehendet vir manum proximi sui et conseretur manus eius super manum proximi sui
ZECH|14|14|sed et Iudas pugnabit adversus Hierusalem et congregabuntur divitiae omnium gentium in circuitu aurum et argentum et vestes multae satis
ZECH|14|15|et sic erit ruina equi et muli cameli et asini et omnium iumentorum quae fuerint in castris illis sicut ruina haec
ZECH|14|16|et omnes qui reliqui fuerint de universis gentibus quae venerint contra Hierusalem ascendent ab anno in annum ut adorent regem Dominum exercituum et celebrent festivitatem tabernaculorum
ZECH|14|17|et erit qui non ascenderit de familiis terrae ad Hierusalem ut adoret regem Dominum exercituum non erit super eos imber
ZECH|14|18|quod si et familia Aegypti non ascenderit et non venerit nec super eos erit sed erit ruina qua percutiet Dominus omnes gentes quae non ascenderint ad celebrandam festivitatem tabernaculorum
ZECH|14|19|hoc erit peccatum Aegypti et hoc peccatum omnium gentium quae non ascenderint ad celebrandam festivitatem tabernaculorum
ZECH|14|20|in die illo erit quod super frenum equi est sanctum Domino et erunt lebetes in domo Domini quasi fialae coram altari
ZECH|14|21|et erit omnis lebes in Hierusalem et in Iuda sanctificatus Domino exercituum et venient omnes immolantes et sument ex eis et coquent in eis et non erit mercator ultra in domo Domini exercituum in die illo
MAL|1|1|onus verbi Domini ad Israhel in manu Malachi
MAL|1|2|dilexi vos dicit Dominus et dixistis in quo dilexisti nos nonne frater erat Esau Iacob dicit Dominus et dilexi Iacob
MAL|1|3|Esau autem odio habui et posui montes eius in solitudinem et hereditatem eius in dracones deserti
MAL|1|4|quod si dixerit Idumea destructi sumus sed revertentes aedificabimus quae deserta sunt haec dicit Dominus exercituum isti aedificabunt et ego destruam et vocabuntur Termini impietatis et Populus cui iratus est Dominus usque in aeternum
MAL|1|5|et oculi vestri videbunt et vos dicetis magnificetur Dominus super terminum Israhel
MAL|1|6|filius honorat patrem et servus dominum suum si ergo pater ego sum ubi est honor meus et si dominus ego sum ubi est timor meus dicit Dominus exercituum ad vos o sacerdotes qui despicitis nomen meum et dixistis in quo despeximus nomen tuum
MAL|1|7|offertis super altare meum panem pollutum et dicitis in quo polluimus te in eo quod dicitis mensa Domini despecta est
MAL|1|8|si offeratis caecum ad immolandum nonne malum est et si offeratis claudum et languidum nonne malum est offer illud duci tuo si placuerit ei aut si susceperit faciem tuam dicit Dominus exercituum
MAL|1|9|et nunc deprecamini vultum Dei ut misereatur vestri de manu enim vestra factum est hoc si quo modo suscipiat facies vestras dicit Dominus exercituum
MAL|1|10|quis est in vobis qui claudat ostia et incendat altare meum gratuito non est mihi voluntas in vobis dicit Dominus exercituum et munus non suscipiam de manu vestra
MAL|1|11|ab ortu enim solis usque ad occasum magnum est nomen meum in gentibus et in omni loco sacrificatur et offertur nomini meo oblatio munda quia magnum nomen meum in gentibus dicit Dominus exercituum
MAL|1|12|et vos polluistis illud in eo quod dicitis mensa Domini contaminata est et quod superponitur contemptibile est cum igni qui illud devorat
MAL|1|13|et dixistis ecce de labore et exsuflastis illud dicit Dominus exercituum et intulistis de rapinis claudum et languidum et intulistis munus numquid suscipiam illud de manu vestra dicit Dominus
MAL|1|14|maledictus dolosus qui habet in grege suo masculum et votum faciens immolat debile Domino quia rex magnus ego dicit Dominus exercituum et nomen meum horribile in gentibus
MAL|2|1|et nunc ad vos mandatum hoc o sacerdotes
MAL|2|2|si nolueritis audire et si nolueritis ponere super cor ut detis gloriam nomini meo ait Dominus exercituum mittam in vos egestatem et maledicam benedictionibus vestris et maledicam illis quoniam non posuistis super cor
MAL|2|3|ecce ego proiciam vobis brachium et dispergam super vultum vestrum stercus sollemnitatum vestrarum et adsumet vos secum
MAL|2|4|et scietis quia misi ad vos mandatum istud ut esset pactum meum cum Levi dicit Dominus exercituum
MAL|2|5|pactum meum fuit cum eo vitae et pacis et dedi ei timorem et timuit me et a facie nominis mei pavebat
MAL|2|6|lex veritatis fuit in ore eius et iniquitas non est inventa in labiis eius in pace et in aequitate ambulavit mecum et multos avertit ab iniquitate
MAL|2|7|labia enim sacerdotis custodient scientiam et legem requirent ex ore eius quia angelus Domini exercituum est
MAL|2|8|vos autem recessistis de via et scandalizastis plurimos in lege irritum fecistis pactum Levi dicit Dominus exercituum
MAL|2|9|propter quod et ego dedi vos contemptibiles et humiles omnibus populis sicut non servastis vias meas et accepistis faciem in lege
MAL|2|10|numquid non pater unus omnium nostrum numquid non Deus unus creavit nos quare ergo despicit unusquisque nostrum fratrem suum violans pactum patrum nostrorum
MAL|2|11|transgressus est Iuda et abominatio facta est in Israhel et in Hierusalem quia contaminavit Iudas sanctificationem Domini quam dilexit et habuit filiam dei alieni
MAL|2|12|disperdat Dominus virum qui fecerit hoc magistrum et discipulum de tabernaculis Iacob et offerentem munus Domino exercituum
MAL|2|13|et hoc rursum fecistis operiebatis lacrimis altare Domini fletu et mugitu ita ut ultra non respiciam ad sacrificium nec accipiam placabile quid de manu vestra
MAL|2|14|et dixistis quam ob causam quia Dominus testificatus est inter te et uxorem pubertatis tuae quam tu despexisti et haec particeps tua et uxor foederis tui
MAL|2|15|nonne unus fecit et residuum spiritus eius est et quid unus quaerit nisi semen Dei custodite ergo spiritum vestrum et uxorem adulescentiae tuae noli despicere
MAL|2|16|cum odio habueris dimitte dicit Dominus Deus Israhel operiet autem iniquitas vestimentum eius dicit Dominus exercituum custodite spiritum vestrum et nolite despicere
MAL|2|17|laborare fecistis Dominum in sermonibus vestris et dixistis in quo eum fecimus laborare in eo cum diceretis omnis qui facit malum bonus est in conspectu Domini et tales ei placent aut certe ubi est Deus iudicii
MAL|3|1|ecce ego mittam angelum meum et praeparabit viam ante faciem meam et statim veniet ad templum suum dominator quem vos quaeritis et angelus testamenti quem vos vultis ecce venit dicit Dominus exercituum
MAL|3|2|et quis poterit cogitare diem adventus eius et quis stabit ad videndum eum ipse enim quasi ignis conflans et quasi herba fullonum
MAL|3|3|et sedebit conflans et emundans argentum et purgabit filios Levi et colabit eos quasi aurum et quasi argentum et erunt Domino offerentes sacrificia in iustitia
MAL|3|4|et placebit Domino sacrificium Iuda et Hierusalem sicut dies saeculi et sicut anni antiqui
MAL|3|5|et accedam ad vos in iudicio et ero testis velox maleficis et adulteris et periuris et qui calumniantur mercedem mercennarii viduas et pupillos et opprimunt peregrinum nec timuerunt me dicit Dominus exercituum
MAL|3|6|ego enim Dominus et non mutor et vos filii Iacob non estis consumpti
MAL|3|7|a diebus enim patrum vestrorum recessistis a legitimis meis et non custodistis revertimini ad me et revertar ad vos dicit Dominus exercituum et dixistis in quo revertemur
MAL|3|8|si adfiget homo Deum quia vos configitis me et dixistis in quo confiximus te in decimis et in primitivis
MAL|3|9|et in penuria vos maledicti estis et me vos configitis gens tota
MAL|3|10|inferte omnem decimam in horreum et sit cibus in domo mea et probate me super hoc dicit Dominus si non aperuero vobis cataractas caeli et effudero vobis benedictionem usque ad abundantiam
MAL|3|11|et increpabo pro vobis devorantem et non corrumpet fructum terrae vestrae nec erit sterilis vinea in agro dicit Dominus exercituum
MAL|3|12|et beatos vos dicent omnes gentes eritis enim vos terra desiderabilis dicit Dominus exercituum
MAL|3|13|invaluerunt super me verba vestra dicit Dominus
MAL|3|14|et dixistis quid locuti sumus contra te dixistis vanus est qui servit Deo et quod emolumentum quia custodivimus praecepta eius et quia ambulavimus tristes coram Domino exercituum
MAL|3|15|ergo nunc beatos dicimus arrogantes siquidem aedificati sunt facientes impietatem et temptaverunt Deum et salvi facti sunt
MAL|3|16|tunc locuti sunt timentes Deum unusquisque cum proximo suo et adtendit Dominus et audivit et scriptus est liber monumenti coram eo timentibus Dominum et cogitantibus nomen eius
MAL|3|17|et erunt mihi ait Dominus exercituum in die qua ego facio in peculium et parcam eis sicut parcit vir filio suo servienti sibi
MAL|3|18|et convertemini et videbitis quid sit inter iustum et impium et inter servientem Deo et non servientem ei
MAL|4|1|ecce enim dies veniet succensa quasi caminus et erunt omnes superbi et omnes facientes impietatem stipula et inflammabit eos dies veniens dicit Dominus exercituum quae non relinquet eis radicem et germen
MAL|4|2|et orietur vobis timentibus nomen meum sol iustitiae et sanitas in pinnis eius et egrediemini et salietis sicut vituli de armento
MAL|4|3|et calcabitis impios cum fuerint cinis sub planta pedum vestrorum in die qua ego facio dicit Dominus exercituum
MAL|4|4|mementote legis Mosi servi mei quam mandavi ei in Choreb ad omnem Israhel praecepta et iudicia
MAL|4|5|ecce ego mittam vobis Heliam prophetam antequam veniat dies Domini magnus et horribilis
MAL|4|6|et convertet cor patrum ad filios et cor filiorum ad patres eorum ne forte veniam et percutiam terram anathemate
MATT|1|1|liber generationis Iesu Christi filii David filii Abraham
MATT|1|2|Abraham genuit Isaac Isaac autem genuit Iacob Iacob autem genuit Iudam et fratres eius
MATT|1|3|Iudas autem genuit Phares et Zara de Thamar Phares autem genuit Esrom Esrom autem genuit Aram
MATT|1|4|Aram autem genuit Aminadab Aminadab autem genuit Naasson Naasson autem genuit Salmon
MATT|1|5|Salmon autem genuit Booz de Rachab Booz autem genuit Obed ex Ruth Obed autem genuit Iesse Iesse autem genuit David regem
MATT|1|6|David autem rex genuit Salomonem ex ea quae fuit Uriae
MATT|1|7|Salomon autem genuit Roboam Roboam autem genuit Abiam Abia autem genuit Asa
MATT|1|8|Asa autem genuit Iosaphat Iosaphat autem genuit Ioram Ioram autem genuit Oziam
MATT|1|9|Ozias autem genuit Ioatham Ioatham autem genuit Achaz Achaz autem genuit Ezechiam
MATT|1|10|Ezechias autem genuit Manassen Manasses autem genuit Amon Amon autem genuit Iosiam
MATT|1|11|Iosias autem genuit Iechoniam et fratres eius in transmigratione Babylonis
MATT|1|12|et post transmigrationem Babylonis Iechonias genuit Salathihel Salathihel autem genuit Zorobabel
MATT|1|13|Zorobabel autem genuit Abiud Abiud autem genuit Eliachim Eliachim autem genuit Azor
MATT|1|14|Azor autem genuit Saddoc Saddoc autem genuit Achim Achim autem genuit Eliud
MATT|1|15|Eliud autem genuit Eleazar Eleazar autem genuit Matthan Matthan autem genuit Iacob
MATT|1|16|Iacob autem genuit Ioseph virum Mariae de qua natus est Iesus qui vocatur Christus
MATT|1|17|omnes ergo generationes ab Abraham usque ad David generationes quattuordecim et a David usque ad transmigrationem Babylonis generationes quattuordecim et a transmigratione Babylonis usque ad Christum generationes quattuordecim
MATT|1|18|Christi autem generatio sic erat cum esset desponsata mater eius Maria Ioseph antequam convenirent inventa est in utero habens de Spiritu Sancto
MATT|1|19|Ioseph autem vir eius cum esset iustus et nollet eam traducere voluit occulte dimittere eam
MATT|1|20|haec autem eo cogitante ecce angelus Domini in somnis apparuit ei dicens Ioseph fili David noli timere accipere Mariam coniugem tuam quod enim in ea natum est de Spiritu Sancto est
MATT|1|21|pariet autem filium et vocabis nomen eius Iesum ipse enim salvum faciet populum suum a peccatis eorum
MATT|1|22|hoc autem totum factum est ut adimpleretur id quod dictum est a Domino per prophetam dicentem
MATT|1|23|ecce virgo in utero habebit et pariet filium et vocabunt nomen eius Emmanuhel quod est interpretatum Nobiscum Deus
MATT|1|24|exsurgens autem Ioseph a somno fecit sicut praecepit ei angelus Domini et accepit coniugem suam
MATT|1|25|et non cognoscebat eam donec peperit filium suum primogenitum et vocavit nomen eius Iesum
MATT|2|1|cum ergo natus esset Iesus in Bethleem Iudaeae in diebus Herodis regis ecce magi ab oriente venerunt Hierosolymam
MATT|2|2|dicentes ubi est qui natus est rex Iudaeorum vidimus enim stellam eius in oriente et venimus adorare eum
MATT|2|3|audiens autem Herodes rex turbatus est et omnis Hierosolyma cum illo
MATT|2|4|et congregans omnes principes sacerdotum et scribas populi sciscitabatur ab eis ubi Christus nasceretur
MATT|2|5|at illi dixerunt ei in Bethleem Iudaeae sic enim scriptum est per prophetam
MATT|2|6|et tu Bethleem terra Iuda nequaquam minima es in principibus Iuda ex te enim exiet dux qui reget populum meum Israhel
MATT|2|7|tunc Herodes clam vocatis magis diligenter didicit ab eis tempus stellae quae apparuit eis
MATT|2|8|et mittens illos in Bethleem dixit ite et interrogate diligenter de puero et cum inveneritis renuntiate mihi ut et ego veniens adorem eum
MATT|2|9|qui cum audissent regem abierunt et ecce stella quam viderant in oriente antecedebat eos usque dum veniens staret supra ubi erat puer
MATT|2|10|videntes autem stellam gavisi sunt gaudio magno valde
MATT|2|11|et intrantes domum invenerunt puerum cum Maria matre eius et procidentes adoraverunt eum et apertis thesauris suis obtulerunt ei munera aurum tus et murram
MATT|2|12|et responso accepto in somnis ne redirent ad Herodem per aliam viam reversi sunt in regionem suam
MATT|2|13|qui cum recessissent ecce angelus Domini apparuit in somnis Ioseph dicens surge et accipe puerum et matrem eius et fuge in Aegyptum et esto ibi usque dum dicam tibi futurum est enim ut Herodes quaerat puerum ad perdendum eum
MATT|2|14|qui consurgens accepit puerum et matrem eius nocte et recessit in Aegyptum
MATT|2|15|et erat ibi usque ad obitum Herodis ut adimpleretur quod dictum est a Domino per prophetam dicentem ex Aegypto vocavi filium meum
MATT|2|16|tunc Herodes videns quoniam inlusus esset a magis iratus est valde et mittens occidit omnes pueros qui erant in Bethleem et in omnibus finibus eius a bimatu et infra secundum tempus quod exquisierat a magis
MATT|2|17|tunc adimpletum est quod dictum est per Hieremiam prophetam dicentem
MATT|2|18|vox in Rama audita est ploratus et ululatus multus Rachel plorans filios suos et noluit consolari quia non sunt
MATT|2|19|defuncto autem Herode ecce apparuit angelus Domini in somnis Ioseph in Aegypto
MATT|2|20|dicens surge et accipe puerum et matrem eius et vade in terram Israhel defuncti sunt enim qui quaerebant animam pueri
MATT|2|21|qui surgens accepit puerum et matrem eius et venit in terram Israhel
MATT|2|22|audiens autem quod Archelaus regnaret in Iudaea pro Herode patre suo timuit illo ire et admonitus in somnis secessit in partes Galilaeae
MATT|2|23|et veniens habitavit in civitate quae vocatur Nazareth ut adimpleretur quod dictum est per prophetas quoniam Nazareus vocabitur
MATT|3|1|in diebus autem illis venit Iohannes Baptista praedicans in deserto Iudaeae
MATT|3|2|et dicens paenitentiam agite adpropinquavit enim regnum caelorum
MATT|3|3|hic est enim qui dictus est per Esaiam prophetam dicentem vox clamantis in deserto parate viam Domini rectas facite semitas eius
MATT|3|4|ipse autem Iohannes habebat vestimentum de pilis camelorum et zonam pelliciam circa lumbos suos esca autem eius erat lucustae et mel silvestre
MATT|3|5|tunc exiebat ad eum Hierosolyma et omnis Iudaea et omnis regio circa Iordanen
MATT|3|6|et baptizabantur in Iordane ab eo confitentes peccata sua
MATT|3|7|videns autem multos Pharisaeorum et Sadducaeorum venientes ad baptismum suum dixit eis progenies viperarum quis demonstravit vobis fugere a futura ira
MATT|3|8|facite ergo fructum dignum paenitentiae
MATT|3|9|et ne velitis dicere intra vos patrem habemus Abraham dico enim vobis quoniam potest Deus de lapidibus istis suscitare filios Abrahae
MATT|3|10|iam enim securis ad radicem arborum posita est omnis ergo arbor quae non facit fructum bonum exciditur et in ignem mittitur
MATT|3|11|ego quidem vos baptizo in aqua in paenitentiam qui autem post me venturus est fortior me est cuius non sum dignus calciamenta portare ipse vos baptizabit in Spiritu Sancto et igni
MATT|3|12|cuius ventilabrum in manu sua et permundabit aream suam et congregabit triticum suum in horreum paleas autem conburet igni inextinguibili
MATT|3|13|tunc venit Iesus a Galilaea in Iordanen ad Iohannem ut baptizaretur ab eo
MATT|3|14|Iohannes autem prohibebat eum dicens ego a te debeo baptizari et tu venis ad me
MATT|3|15|respondens autem Iesus dixit ei sine modo sic enim decet nos implere omnem iustitiam tunc dimisit eum
MATT|3|16|baptizatus autem confestim ascendit de aqua et ecce aperti sunt ei caeli et vidit Spiritum Dei descendentem sicut columbam venientem super se
MATT|3|17|et ecce vox de caelis dicens hic est Filius meus dilectus in quo mihi conplacui
MATT|4|1|tunc Iesus ductus est in desertum ab Spiritu ut temptaretur a diabolo
MATT|4|2|et cum ieiunasset quadraginta diebus et quadraginta noctibus postea esuriit
MATT|4|3|et accedens temptator dixit ei si Filius Dei es dic ut lapides isti panes fiant
MATT|4|4|qui respondens dixit scriptum est non in pane solo vivet homo sed in omni verbo quod procedit de ore Dei
MATT|4|5|tunc adsumit eum diabolus in sanctam civitatem et statuit eum supra pinnaculum templi
MATT|4|6|et dixit ei si Filius Dei es mitte te deorsum scriptum est enim quia angelis suis mandabit de te et in manibus tollent te ne forte offendas ad lapidem pedem tuum
MATT|4|7|ait illi Iesus rursum scriptum est non temptabis Dominum Deum tuum
MATT|4|8|iterum adsumit eum diabolus in montem excelsum valde et ostendit ei omnia regna mundi et gloriam eorum
MATT|4|9|et dixit illi haec tibi omnia dabo si cadens adoraveris me
MATT|4|10|tunc dicit ei Iesus vade Satanas scriptum est Dominum Deum tuum adorabis et illi soli servies
MATT|4|11|tunc reliquit eum diabolus et ecce angeli accesserunt et ministrabant ei
MATT|4|12|cum autem audisset quod Iohannes traditus esset secessit in Galilaeam
MATT|4|13|et relicta civitate Nazareth venit et habitavit in Capharnaum maritimam in finibus Zabulon et Nepthalim
MATT|4|14|ut adimpleretur quod dictum est per Esaiam prophetam
MATT|4|15|terra Zabulon et terra Nepthalim via maris trans Iordanen Galilaeae gentium
MATT|4|16|populus qui sedebat in tenebris lucem vidit magnam et sedentibus in regione et umbra mortis lux orta est eis
MATT|4|17|exinde coepit Iesus praedicare et dicere paenitentiam agite adpropinquavit enim regnum caelorum
MATT|4|18|ambulans autem iuxta mare Galilaeae vidit duos fratres Simonem qui vocatur Petrus et Andream fratrem eius mittentes rete in mare erant enim piscatores
MATT|4|19|et ait illis venite post me et faciam vos fieri piscatores hominum
MATT|4|20|at illi continuo relictis retibus secuti sunt eum
MATT|4|21|et procedens inde vidit alios duos fratres Iacobum Zebedaei et Iohannem fratrem eius in navi cum Zebedaeo patre eorum reficientes retia sua et vocavit eos
MATT|4|22|illi autem statim relictis retibus et patre secuti sunt eum
MATT|4|23|et circumibat Iesus totam Galilaeam docens in synagogis eorum et praedicans evangelium regni et sanans omnem languorem et omnem infirmitatem in populo
MATT|4|24|et abiit opinio eius in totam Syriam et obtulerunt ei omnes male habentes variis languoribus et tormentis conprehensos et qui daemonia habebant et lunaticos et paralyticos et curavit eos
MATT|4|25|et secutae sunt eum turbae multae de Galilaea et Decapoli et Hierosolymis et Iudaea et de trans Iordanen
MATT|5|1|videns autem turbas ascendit in montem et cum sedisset accesserunt ad eum discipuli eius
MATT|5|2|et aperiens os suum docebat eos dicens
MATT|5|3|beati pauperes spiritu quoniam ipsorum est regnum caelorum
MATT|5|4|beati mites quoniam ipsi possidebunt terram
MATT|5|5|beati qui lugent quoniam ipsi consolabuntur
MATT|5|6|beati qui esuriunt et sitiunt iustitiam quoniam ipsi saturabuntur
MATT|5|7|beati misericordes quia ipsi misericordiam consequentur
MATT|5|8|beati mundo corde quoniam ipsi Deum videbunt
MATT|5|9|beati pacifici quoniam filii Dei vocabuntur
MATT|5|10|beati qui persecutionem patiuntur propter iustitiam quoniam ipsorum est regnum caelorum
MATT|5|11|beati estis cum maledixerint vobis et persecuti vos fuerint et dixerint omne malum adversum vos mentientes propter me
MATT|5|12|gaudete et exultate quoniam merces vestra copiosa est in caelis sic enim persecuti sunt prophetas qui fuerunt ante vos
MATT|5|13|vos estis sal terrae quod si sal evanuerit in quo sallietur ad nihilum valet ultra nisi ut mittatur foras et conculcetur ab hominibus
MATT|5|14|vos estis lux mundi non potest civitas abscondi supra montem posita
MATT|5|15|neque accendunt lucernam et ponunt eam sub modio sed super candelabrum ut luceat omnibus qui in domo sunt
MATT|5|16|sic luceat lux vestra coram hominibus ut videant vestra bona opera et glorificent Patrem vestrum qui in caelis est
MATT|5|17|nolite putare quoniam veni solvere legem aut prophetas non veni solvere sed adimplere
MATT|5|18|amen quippe dico vobis donec transeat caelum et terra iota unum aut unus apex non praeteribit a lege donec omnia fiant
MATT|5|19|qui ergo solverit unum de mandatis istis minimis et docuerit sic homines minimus vocabitur in regno caelorum qui autem fecerit et docuerit hic magnus vocabitur in regno caelorum
MATT|5|20|dico enim vobis quia nisi abundaverit iustitia vestra plus quam scribarum et Pharisaeorum non intrabitis in regnum caelorum
MATT|5|21|audistis quia dictum est antiquis non occides qui autem occiderit reus erit iudicio
MATT|5|22|ego autem dico vobis quia omnis qui irascitur fratri suo reus erit iudicio qui autem dixerit fratri suo racha reus erit concilio qui autem dixerit fatue reus erit gehennae ignis
MATT|5|23|si ergo offeres munus tuum ad altare et ibi recordatus fueris quia frater tuus habet aliquid adversum te
MATT|5|24|relinque ibi munus tuum ante altare et vade prius reconciliare fratri tuo et tunc veniens offers munus tuum
MATT|5|25|esto consentiens adversario tuo cito dum es in via cum eo ne forte tradat te adversarius iudici et iudex tradat te ministro et in carcerem mittaris
MATT|5|26|amen dico tibi non exies inde donec reddas novissimum quadrantem
MATT|5|27|audistis quia dictum est antiquis non moechaberis
MATT|5|28|ego autem dico vobis quoniam omnis qui viderit mulierem ad concupiscendum eam iam moechatus est eam in corde suo
MATT|5|29|quod si oculus tuus dexter scandalizat te erue eum et proice abs te expedit enim tibi ut pereat unum membrorum tuorum quam totum corpus tuum mittatur in gehennam
MATT|5|30|et si dextera manus tua scandalizat te abscide eam et proice abs te expedit tibi ut pereat unum membrorum tuorum quam totum corpus tuum eat in gehennam
MATT|5|31|dictum est autem quicumque dimiserit uxorem suam det illi libellum repudii
MATT|5|32|ego autem dico vobis quia omnis qui dimiserit uxorem suam excepta fornicationis causa facit eam moechari et qui dimissam duxerit adulterat
MATT|5|33|iterum audistis quia dictum est antiquis non peierabis reddes autem Domino iuramenta tua
MATT|5|34|ego autem dico vobis non iurare omnino neque per caelum quia thronus Dei est
MATT|5|35|neque per terram quia scabillum est pedum eius neque per Hierosolymam quia civitas est magni Regis
MATT|5|36|neque per caput tuum iuraveris quia non potes unum capillum album facere aut nigrum
MATT|5|37|sit autem sermo vester est est non non quod autem his abundantius est a malo est
MATT|5|38|audistis quia dictum est oculum pro oculo et dentem pro dente
MATT|5|39|ego autem dico vobis non resistere malo sed si quis te percusserit in dextera maxilla tua praebe illi et alteram
MATT|5|40|et ei qui vult tecum iudicio contendere et tunicam tuam tollere remitte ei et pallium
MATT|5|41|et quicumque te angariaverit mille passus vade cum illo alia duo
MATT|5|42|qui petit a te da ei et volenti mutuari a te ne avertaris
MATT|5|43|audistis quia dictum est diliges proximum tuum et odio habebis inimicum tuum
MATT|5|44|ego autem dico vobis diligite inimicos vestros benefacite his qui oderunt vos et orate pro persequentibus et calumniantibus vos
MATT|5|45|ut sitis filii Patris vestri qui in caelis est qui solem suum oriri facit super bonos et malos et pluit super iustos et iniustos
MATT|5|46|si enim diligatis eos qui vos diligunt quam mercedem habebitis nonne et publicani hoc faciunt
MATT|5|47|et si salutaveritis fratres vestros tantum quid amplius facitis nonne et ethnici hoc faciunt
MATT|5|48|estote ergo vos perfecti sicut et Pater vester caelestis perfectus est
MATT|6|1|adtendite ne iustitiam vestram faciatis coram hominibus ut videamini ab eis alioquin mercedem non habebitis apud Patrem vestrum qui in caelis est
MATT|6|2|cum ergo facies elemosynam noli tuba canere ante te sicut hypocritae faciunt in synagogis et in vicis ut honorificentur ab hominibus amen dico vobis receperunt mercedem suam
MATT|6|3|te autem faciente elemosynam nesciat sinistra tua quid faciat dextera tua
MATT|6|4|ut sit elemosyna tua in abscondito et Pater tuus qui videt in abscondito reddet tibi
MATT|6|5|et cum oratis non eritis sicut hypocritae qui amant in synagogis et in angulis platearum stantes orare ut videantur ab hominibus amen dico vobis receperunt mercedem suam
MATT|6|6|tu autem cum orabis intra in cubiculum tuum et cluso ostio tuo ora Patrem tuum in abscondito et Pater tuus qui videt in abscondito reddet tibi
MATT|6|7|orantes autem nolite multum loqui sicut ethnici putant enim quia in multiloquio suo exaudiantur
MATT|6|8|nolite ergo adsimilari eis scit enim Pater vester quibus opus sit vobis antequam petatis eum
MATT|6|9|sic ergo vos orabitis Pater noster qui in caelis es sanctificetur nomen tuum
MATT|6|10|veniat regnum tuum fiat voluntas tua sicut in caelo et in terra
MATT|6|11|panem nostrum supersubstantialem da nobis hodie
MATT|6|12|et dimitte nobis debita nostra sicut et nos dimisimus debitoribus nostris
MATT|6|13|et ne inducas nos in temptationem sed libera nos a malo
MATT|6|14|si enim dimiseritis hominibus peccata eorum dimittet et vobis Pater vester caelestis delicta vestra
MATT|6|15|si autem non dimiseritis hominibus nec Pater vester dimittet peccata vestra
MATT|6|16|cum autem ieiunatis nolite fieri sicut hypocritae tristes demoliuntur enim facies suas ut pareant hominibus ieiunantes amen dico vobis quia receperunt mercedem suam
MATT|6|17|tu autem cum ieiunas ungue caput tuum et faciem tuam lava
MATT|6|18|ne videaris hominibus ieiunans sed Patri tuo qui est in abscondito et Pater tuus qui videt in abscondito reddet tibi
MATT|6|19|nolite thesaurizare vobis thesauros in terra ubi erugo et tinea demolitur ubi fures effodiunt et furantur
MATT|6|20|thesaurizate autem vobis thesauros in caelo ubi neque erugo neque tinea demolitur et ubi fures non effodiunt nec furantur
MATT|6|21|ubi enim est thesaurus tuus ibi est et cor tuum
MATT|6|22|lucerna corporis est oculus si fuerit oculus tuus simplex totum corpus tuum lucidum erit
MATT|6|23|si autem oculus tuus nequam fuerit totum corpus tuum tenebrosum erit si ergo lumen quod in te est tenebrae sunt tenebrae quantae erunt
MATT|6|24|nemo potest duobus dominis servire aut enim unum odio habebit et alterum diliget aut unum sustinebit et alterum contemnet non potestis Deo servire et mamonae
MATT|6|25|ideo dico vobis ne solliciti sitis animae vestrae quid manducetis neque corpori vestro quid induamini nonne anima plus est quam esca et corpus plus est quam vestimentum
MATT|6|26|respicite volatilia caeli quoniam non serunt neque metunt neque congregant in horrea et Pater vester caelestis pascit illa nonne vos magis pluris estis illis
MATT|6|27|quis autem vestrum cogitans potest adicere ad staturam suam cubitum unum
MATT|6|28|et de vestimento quid solliciti estis considerate lilia agri quomodo crescunt non laborant nec nent
MATT|6|29|dico autem vobis quoniam nec Salomon in omni gloria sua coopertus est sicut unum ex istis
MATT|6|30|si autem faenum agri quod hodie est et cras in clibanum mittitur Deus sic vestit quanto magis vos minimae fidei
MATT|6|31|nolite ergo solliciti esse dicentes quid manducabimus aut quid bibemus aut quo operiemur
MATT|6|32|haec enim omnia gentes inquirunt scit enim Pater vester quia his omnibus indigetis
MATT|6|33|quaerite autem primum regnum et iustitiam eius et omnia haec adicientur vobis
MATT|6|34|nolite ergo esse solliciti in crastinum crastinus enim dies sollicitus erit sibi ipse sufficit diei malitia sua
MATT|7|1|nolite iudicare ut non iudicemini
MATT|7|2|in quo enim iudicio iudicaveritis iudicabimini et in qua mensura mensi fueritis metietur vobis
MATT|7|3|quid autem vides festucam in oculo fratris tui et trabem in oculo tuo non vides
MATT|7|4|aut quomodo dicis fratri tuo sine eiciam festucam de oculo tuo et ecce trabis est in oculo tuo
MATT|7|5|hypocrita eice primum trabem de oculo tuo et tunc videbis eicere festucam de oculo fratris tui
MATT|7|6|nolite dare sanctum canibus neque mittatis margaritas vestras ante porcos ne forte conculcent eas pedibus suis et conversi disrumpant vos
MATT|7|7|petite et dabitur vobis quaerite et invenietis pulsate et aperietur vobis
MATT|7|8|omnis enim qui petit accipit et qui quaerit invenit et pulsanti aperietur
MATT|7|9|aut quis est ex vobis homo quem si petierit filius suus panem numquid lapidem porriget ei
MATT|7|10|aut si piscem petet numquid serpentem porriget ei
MATT|7|11|si ergo vos cum sitis mali nostis bona dare filiis vestris quanto magis Pater vester qui in caelis est dabit bona petentibus se
MATT|7|12|omnia ergo quaecumque vultis ut faciant vobis homines et vos facite eis haec est enim lex et prophetae
MATT|7|13|intrate per angustam portam quia lata porta et spatiosa via quae ducit ad perditionem et multi sunt qui intrant per eam
MATT|7|14|quam angusta porta et arta via quae ducit ad vitam et pauci sunt qui inveniunt eam
MATT|7|15|adtendite a falsis prophetis qui veniunt ad vos in vestimentis ovium intrinsecus autem sunt lupi rapaces
MATT|7|16|a fructibus eorum cognoscetis eos numquid colligunt de spinis uvas aut de tribulis ficus
MATT|7|17|sic omnis arbor bona fructus bonos facit mala autem arbor fructus malos facit
MATT|7|18|non potest arbor bona fructus malos facere neque arbor mala fructus bonos facere
MATT|7|19|omnis arbor quae non facit fructum bonum exciditur et in ignem mittitur
MATT|7|20|igitur ex fructibus eorum cognoscetis eos
MATT|7|21|non omnis qui dicit mihi Domine Domine intrabit in regnum caelorum sed qui facit voluntatem Patris mei qui in caelis est ipse intrabit in regnum caelorum
MATT|7|22|multi dicent mihi in illa die Domine Domine nonne in nomine tuo prophetavimus et in tuo nomine daemonia eiecimus et in tuo nomine virtutes multas fecimus
MATT|7|23|et tunc confitebor illis quia numquam novi vos discedite a me qui operamini iniquitatem
MATT|7|24|omnis ergo qui audit verba mea haec et facit ea adsimilabitur viro sapienti qui aedificavit domum suam supra petram
MATT|7|25|et descendit pluvia et venerunt flumina et flaverunt venti et inruerunt in domum illam et non cecidit fundata enim erat super petram
MATT|7|26|et omnis qui audit verba mea haec et non facit ea similis erit viro stulto qui aedificavit domum suam supra harenam
MATT|7|27|et descendit pluvia et venerunt flumina et flaverunt venti et inruerunt in domum illam et cecidit et fuit ruina eius magna
MATT|7|28|et factum est cum consummasset Iesus verba haec admirabantur turbae super doctrinam eius
MATT|7|29|erat enim docens eos sicut potestatem habens non sicut scribae eorum et Pharisaei
MATT|8|1|cum autem descendisset de monte secutae sunt eum turbae multae
MATT|8|2|et ecce leprosus veniens adorabat eum dicens Domine si vis potes me mundare
MATT|8|3|et extendens manum tetigit eum Iesus dicens volo mundare et confestim mundata est lepra eius
MATT|8|4|et ait illi Iesus vide nemini dixeris sed vade ostende te sacerdoti et offer munus quod praecepit Moses in testimonium illis
MATT|8|5|cum autem introisset Capharnaum accessit ad eum centurio rogans eum
MATT|8|6|et dicens Domine puer meus iacet in domo paralyticus et male torquetur
MATT|8|7|et ait illi Iesus ego veniam et curabo eum
MATT|8|8|et respondens centurio ait Domine non sum dignus ut intres sub tectum meum sed tantum dic verbo et sanabitur puer meus
MATT|8|9|nam et ego homo sum sub potestate habens sub me milites et dico huic vade et vadit et alio veni et venit et servo meo fac hoc et facit
MATT|8|10|audiens autem Iesus miratus est et sequentibus se dixit amen dico vobis non inveni tantam fidem in Israhel
MATT|8|11|dico autem vobis quod multi ab oriente et occidente venient et recumbent cum Abraham et Isaac et Iacob in regno caelorum
MATT|8|12|filii autem regni eicientur in tenebras exteriores ibi erit fletus et stridor dentium
MATT|8|13|et dixit Iesus centurioni vade et sicut credidisti fiat tibi et sanatus est puer in hora illa
MATT|8|14|et cum venisset Iesus in domum Petri vidit socrum eius iacentem et febricitantem
MATT|8|15|et tetigit manum eius et dimisit eam febris et surrexit et ministrabat eis
MATT|8|16|vespere autem facto obtulerunt ei multos daemonia habentes et eiciebat spiritus verbo et omnes male habentes curavit
MATT|8|17|ut adimpleretur quod dictum est per Esaiam prophetam dicentem ipse infirmitates nostras accepit et aegrotationes portavit
MATT|8|18|videns autem Iesus turbas multas circum se iussit ire trans fretum
MATT|8|19|et accedens unus scriba ait illi magister sequar te quocumque ieris
MATT|8|20|et dicit ei Iesus vulpes foveas habent et volucres caeli tabernacula Filius autem hominis non habet ubi caput reclinet
MATT|8|21|alius autem de discipulis eius ait illi Domine permitte me primum ire et sepelire patrem meum
MATT|8|22|Iesus autem ait illi sequere me et dimitte mortuos sepelire mortuos suos
MATT|8|23|et ascendente eo in navicula secuti sunt eum discipuli eius
MATT|8|24|et ecce motus magnus factus est in mari ita ut navicula operiretur fluctibus ipse vero dormiebat
MATT|8|25|et accesserunt et suscitaverunt eum dicentes Domine salva nos perimus
MATT|8|26|et dicit eis quid timidi estis modicae fidei tunc surgens imperavit ventis et mari et facta est tranquillitas magna
MATT|8|27|porro homines mirati sunt dicentes qualis est hic quia et venti et mare oboediunt ei
MATT|8|28|et cum venisset trans fretum in regionem Gerasenorum occurrerunt ei duo habentes daemonia de monumentis exeuntes saevi nimis ita ut nemo posset transire per viam illam
MATT|8|29|et ecce clamaverunt dicentes quid nobis et tibi Fili Dei venisti huc ante tempus torquere nos
MATT|8|30|erat autem non longe ab illis grex porcorum multorum pascens
MATT|8|31|daemones autem rogabant eum dicentes si eicis nos mitte nos in gregem porcorum
MATT|8|32|et ait illis ite at illi exeuntes abierunt in porcos et ecce impetu abiit totus grex per praeceps in mare et mortui sunt in aquis
MATT|8|33|pastores autem fugerunt et venientes in civitatem nuntiaverunt omnia et de his qui daemonia habuerant
MATT|8|34|et ecce tota civitas exiit obviam Iesu et viso eo rogabant ut transiret a finibus eorum
MATT|9|1|et ascendens in naviculam transfretavit et venit in civitatem suam
MATT|9|2|et ecce offerebant ei paralyticum iacentem in lecto et videns Iesus fidem illorum dixit paralytico confide fili remittuntur tibi peccata tua
MATT|9|3|et ecce quidam de scribis dixerunt intra se hic blasphemat
MATT|9|4|et cum vidisset Iesus cogitationes eorum dixit ut quid cogitatis mala in cordibus vestris
MATT|9|5|quid est facilius dicere dimittuntur tibi peccata aut dicere surge et ambula
MATT|9|6|ut sciatis autem quoniam Filius hominis habet potestatem in terra dimittendi peccata tunc ait paralytico surge tolle lectum tuum et vade in domum tuam
MATT|9|7|et surrexit et abiit in domum suam
MATT|9|8|videntes autem turbae timuerunt et glorificaverunt Deum qui dedit potestatem talem hominibus
MATT|9|9|et cum transiret inde Iesus vidit hominem sedentem in teloneo Mattheum nomine et ait illi sequere me et surgens secutus est eum
MATT|9|10|et factum est discumbente eo in domo ecce multi publicani et peccatores venientes discumbebant cum Iesu et discipulis eius
MATT|9|11|et videntes Pharisaei dicebant discipulis eius quare cum publicanis et peccatoribus manducat magister vester
MATT|9|12|at Iesus audiens ait non est opus valentibus medico sed male habentibus
MATT|9|13|euntes autem discite quid est misericordiam volo et non sacrificium non enim veni vocare iustos sed peccatores
MATT|9|14|tunc accesserunt ad eum discipuli Iohannis dicentes quare nos et Pharisaei ieiunamus frequenter discipuli autem tui non ieiunant
MATT|9|15|et ait illis Iesus numquid possunt filii sponsi lugere quamdiu cum illis est sponsus venient autem dies cum auferetur ab eis sponsus et tunc ieiunabunt
MATT|9|16|nemo autem inmittit commissuram panni rudis in vestimentum vetus tollit enim plenitudinem eius a vestimento et peior scissura fit
MATT|9|17|neque mittunt vinum novum in utres veteres alioquin rumpuntur utres et vinum effunditur et utres pereunt sed vinum novum in utres novos mittunt et ambo conservantur
MATT|9|18|haec illo loquente ad eos ecce princeps unus accessit et adorabat eum dicens filia mea modo defuncta est sed veni inpone manum super eam et vivet
MATT|9|19|et surgens Iesus sequebatur eum et discipuli eius
MATT|9|20|et ecce mulier quae sanguinis fluxum patiebatur duodecim annis accessit retro et tetigit fimbriam vestimenti eius
MATT|9|21|dicebat enim intra se si tetigero tantum vestimentum eius salva ero
MATT|9|22|at Iesus conversus et videns eam dixit confide filia fides tua te salvam fecit et salva facta est mulier ex illa hora
MATT|9|23|et cum venisset Iesus in domum principis et vidisset tibicines et turbam tumultuantem
MATT|9|24|dicebat recedite non est enim mortua puella sed dormit et deridebant eum
MATT|9|25|et cum eiecta esset turba intravit et tenuit manum eius et surrexit puella
MATT|9|26|et exiit fama haec in universam terram illam
MATT|9|27|et transeunte inde Iesu secuti sunt eum duo caeci clamantes et dicentes miserere nostri Fili David
MATT|9|28|cum autem venisset domum accesserunt ad eum caeci et dicit eis Iesus creditis quia possum hoc facere vobis dicunt ei utique Domine
MATT|9|29|tunc tetigit oculos eorum dicens secundum fidem vestram fiat vobis
MATT|9|30|et aperti sunt oculi illorum et comminatus est illis Iesus dicens videte ne quis sciat
MATT|9|31|illi autem exeuntes diffamaverunt eum in tota terra illa
MATT|9|32|egressis autem illis ecce obtulerunt ei hominem mutum daemonium habentem
MATT|9|33|et eiecto daemone locutus est mutus et miratae sunt turbae dicentes numquam paruit sic in Israhel
MATT|9|34|Pharisaei autem dicebant in principe daemoniorum eicit daemones
MATT|9|35|et circumibat Iesus civitates omnes et castella docens in synagogis eorum et praedicans evangelium regni et curans omnem languorem et omnem infirmitatem
MATT|9|36|videns autem turbas misertus est eis quia erant vexati et iacentes sicut oves non habentes pastorem
MATT|9|37|tunc dicit discipulis suis messis quidem multa operarii autem pauci
MATT|9|38|rogate ergo dominum messis ut eiciat operarios in messem suam
MATT|10|1|et convocatis duodecim discipulis suis dedit illis potestatem spirituum inmundorum ut eicerent eos et curarent omnem languorem et omnem infirmitatem
MATT|10|2|duodecim autem apostolorum nomina sunt haec primus Simon qui dicitur Petrus et Andreas frater eius
MATT|10|3|Iacobus Zebedaei et Iohannes frater eius Philippus et Bartholomeus Thomas et Mattheus publicanus et Iacobus Alphei et Thaddeus
MATT|10|4|Simon Cananeus et Iudas Scariotes qui et tradidit eum
MATT|10|5|hos duodecim misit Iesus praecipiens eis et dicens in viam gentium ne abieritis et in civitates Samaritanorum ne intraveritis
MATT|10|6|sed potius ite ad oves quae perierunt domus Israhel
MATT|10|7|euntes autem praedicate dicentes quia adpropinquavit regnum caelorum
MATT|10|8|infirmos curate mortuos suscitate leprosos mundate daemones eicite gratis accepistis gratis date
MATT|10|9|nolite possidere aurum neque argentum neque pecuniam in zonis vestris
MATT|10|10|non peram in via neque duas tunicas neque calciamenta neque virgam dignus enim est operarius cibo suo
MATT|10|11|in quamcumque civitatem aut castellum intraveritis interrogate quis in ea dignus sit et ibi manete donec exeatis
MATT|10|12|intrantes autem in domum salutate eam
MATT|10|13|et siquidem fuerit domus digna veniat pax vestra super eam si autem non fuerit digna pax vestra ad vos revertatur
MATT|10|14|et quicumque non receperit vos neque audierit sermones vestros exeuntes foras de domo vel de civitate excutite pulverem de pedibus vestris
MATT|10|15|amen dico vobis tolerabilius erit terrae Sodomorum et Gomorraeorum in die iudicii quam illi civitati
MATT|10|16|ecce ego mitto vos sicut oves in medio luporum estote ergo prudentes sicut serpentes et simplices sicut columbae
MATT|10|17|cavete autem ab hominibus tradent enim vos in conciliis et in synagogis suis flagellabunt vos
MATT|10|18|et ad praesides et ad reges ducemini propter me in testimonium illis et gentibus
MATT|10|19|cum autem tradent vos nolite cogitare quomodo aut quid loquamini dabitur enim vobis in illa hora quid loquamini
MATT|10|20|non enim vos estis qui loquimini sed Spiritus Patris vestri qui loquitur in vobis
MATT|10|21|tradet autem frater fratrem in mortem et pater filium et insurgent filii in parentes et morte eos adficient
MATT|10|22|et eritis odio omnibus propter nomen meum qui autem perseveraverit in finem hic salvus erit
MATT|10|23|cum autem persequentur vos in civitate ista fugite in aliam amen enim dico vobis non consummabitis civitates Israhel donec veniat Filius hominis
MATT|10|24|non est discipulus super magistrum nec servus super dominum suum
MATT|10|25|sufficit discipulo ut sit sicut magister eius et servus sicut dominus eius si patrem familias Beelzebub vocaverunt quanto magis domesticos eius
MATT|10|26|ne ergo timueritis eos nihil enim opertum quod non revelabitur et occultum quod non scietur
MATT|10|27|quod dico vobis in tenebris dicite in lumine et quod in aure auditis praedicate super tecta
MATT|10|28|et nolite timere eos qui occidunt corpus animam autem non possunt occidere sed potius eum timete qui potest et animam et corpus perdere in gehennam
MATT|10|29|nonne duo passeres asse veneunt et unus ex illis non cadet super terram sine Patre vestro
MATT|10|30|vestri autem et capilli capitis omnes numerati sunt
MATT|10|31|nolite ergo timere multis passeribus meliores estis vos
MATT|10|32|omnis ergo qui confitebitur me coram hominibus confitebor et ego eum coram Patre meo qui est in caelis
MATT|10|33|qui autem negaverit me coram hominibus negabo et ego eum coram Patre meo qui est in caelis
MATT|10|34|nolite arbitrari quia venerim mittere pacem in terram non veni pacem mittere sed gladium
MATT|10|35|veni enim separare hominem adversus patrem suum et filiam adversus matrem suam et nurum adversus socrum suam
MATT|10|36|et inimici hominis domestici eius
MATT|10|37|qui amat patrem aut matrem plus quam me non est me dignus et qui amat filium aut filiam super me non est me dignus
MATT|10|38|et qui non accipit crucem suam et sequitur me non est me dignus
MATT|10|39|qui invenit animam suam perdet illam et qui perdiderit animam suam propter me inveniet eam
MATT|10|40|qui recipit vos me recipit et qui me recipit recipit eum qui me misit
MATT|10|41|qui recipit prophetam in nomine prophetae mercedem prophetae accipiet et qui recipit iustum in nomine iusti mercedem iusti accipiet
MATT|10|42|et quicumque potum dederit uni ex minimis istis calicem aquae frigidae tantum in nomine discipuli amen dico vobis non perdet mercedem suam
MATT|11|1|et factum est cum consummasset Iesus praecipiens duodecim discipulis suis transiit inde ut doceret et praedicaret in civitatibus eorum
MATT|11|2|Iohannes autem cum audisset in vinculis opera Christi mittens duos de discipulis suis
MATT|11|3|ait illi tu es qui venturus es an alium expectamus
MATT|11|4|et respondens Iesus ait illis euntes renuntiate Iohanni quae auditis et videtis
MATT|11|5|caeci vident claudi ambulant leprosi mundantur surdi audiunt mortui resurgunt pauperes evangelizantur
MATT|11|6|et beatus est qui non fuerit scandalizatus in me
MATT|11|7|illis autem abeuntibus coepit Iesus dicere ad turbas de Iohanne quid existis in desertum videre harundinem vento agitatam
MATT|11|8|sed quid existis videre hominem mollibus vestitum ecce qui mollibus vestiuntur in domibus regum sunt
MATT|11|9|sed quid existis videre prophetam etiam dico vobis et plus quam prophetam
MATT|11|10|hic enim est de quo scriptum est ecce ego mitto angelum meum ante faciem tuam qui praeparabit viam tuam ante te
MATT|11|11|amen dico vobis non surrexit inter natos mulierum maior Iohanne Baptista qui autem minor est in regno caelorum maior est illo
MATT|11|12|a diebus autem Iohannis Baptistae usque nunc regnum caelorum vim patitur et violenti rapiunt illud
MATT|11|13|omnes enim prophetae et lex usque ad Iohannem prophetaverunt
MATT|11|14|et si vultis recipere ipse est Helias qui venturus est
MATT|11|15|qui habet aures audiendi audiat
MATT|11|16|cui autem similem aestimabo generationem istam similis est pueris sedentibus in foro qui clamantes coaequalibus
MATT|11|17|dicunt cecinimus vobis et non saltastis lamentavimus et non planxistis
MATT|11|18|venit enim Iohannes neque manducans neque bibens et dicunt daemonium habet
MATT|11|19|venit Filius hominis manducans et bibens et dicunt ecce homo vorax et potator vini publicanorum et peccatorum amicus et iustificata est sapientia a filiis suis
MATT|11|20|tunc coepit exprobrare civitatibus in quibus factae sunt plurimae virtutes eius quia non egissent paenitentiam
MATT|11|21|vae tibi Corazain vae tibi Bethsaida quia si in Tyro et Sidone factae essent virtutes quae factae sunt in vobis olim in cilicio et cinere paenitentiam egissent
MATT|11|22|verumtamen dico vobis Tyro et Sidoni remissius erit in die iudicii quam vobis
MATT|11|23|et tu Capharnaum numquid usque in caelum exaltaberis usque in infernum descendes quia si in Sodomis factae fuissent virtutes quae factae sunt in te forte mansissent usque in hunc diem
MATT|11|24|verumtamen dico vobis quia terrae Sodomorum remissius erit in die iudicii quam tibi
MATT|11|25|in illo tempore respondens Iesus dixit confiteor tibi Pater Domine caeli et terrae quia abscondisti haec a sapientibus et prudentibus et revelasti ea parvulis
MATT|11|26|ita Pater quoniam sic fuit placitum ante te
MATT|11|27|omnia mihi tradita sunt a Patre meo et nemo novit Filium nisi Pater neque Patrem quis novit nisi Filius et cui voluerit Filius revelare
MATT|11|28|venite ad me omnes qui laboratis et onerati estis et ego reficiam vos
MATT|11|29|tollite iugum meum super vos et discite a me quia mitis sum et humilis corde et invenietis requiem animabus vestris
MATT|11|30|iugum enim meum suave est et onus meum leve est
MATT|12|1|in illo tempore abiit Iesus sabbato per sata discipuli autem eius esurientes coeperunt vellere spicas et manducare
MATT|12|2|Pharisaei autem videntes dixerunt ei ecce discipuli tui faciunt quod non licet eis facere sabbatis
MATT|12|3|at ille dixit eis non legistis quid fecerit David quando esuriit et qui cum eo erant
MATT|12|4|quomodo intravit in domum Dei et panes propositionis comedit quos non licebat ei edere neque his qui cum eo erant nisi solis sacerdotibus
MATT|12|5|aut non legistis in lege quia sabbatis sacerdotes in templo sabbatum violant et sine crimine sunt
MATT|12|6|dico autem vobis quia templo maior est hic
MATT|12|7|si autem sciretis quid est misericordiam volo et non sacrificium numquam condemnassetis innocentes
MATT|12|8|dominus est enim Filius hominis etiam sabbati
MATT|12|9|et cum inde transisset venit in synagogam eorum
MATT|12|10|et ecce homo manum habens aridam et interrogabant eum dicentes si licet sabbatis curare ut accusarent eum
MATT|12|11|ipse autem dixit illis quis erit ex vobis homo qui habeat ovem unam et si ceciderit haec sabbatis in foveam nonne tenebit et levabit eam
MATT|12|12|quanto magis melior est homo ove itaque licet sabbatis benefacere
MATT|12|13|tunc ait homini extende manum tuam et extendit et restituta est sanitati sicut altera
MATT|12|14|exeuntes autem Pharisaei consilium faciebant adversus eum quomodo eum perderent
MATT|12|15|Iesus autem sciens recessit inde et secuti sunt eum multi et curavit eos omnes
MATT|12|16|et praecepit eis ne manifestum eum facerent
MATT|12|17|ut adimpleretur quod dictum est per Esaiam prophetam dicentem
MATT|12|18|ecce puer meus quem elegi dilectus meus in quo bene placuit animae meae ponam spiritum meum super eum et iudicium gentibus nuntiabit
MATT|12|19|non contendet neque clamabit neque audiet aliquis in plateis vocem eius
MATT|12|20|harundinem quassatam non confringet et linum fumigans non extinguet donec eiciat ad victoriam iudicium
MATT|12|21|et in nomine eius gentes sperabunt
MATT|12|22|tunc oblatus est ei daemonium habens caecus et mutus et curavit eum ita ut loqueretur et videret
MATT|12|23|et stupebant omnes turbae et dicebant numquid hic est Filius David
MATT|12|24|Pharisaei autem audientes dixerunt hic non eicit daemones nisi in Beelzebub principe daemoniorum
MATT|12|25|Iesus autem sciens cogitationes eorum dixit eis omne regnum divisum contra se desolatur et omnis civitas vel domus divisa contra se non stabit
MATT|12|26|et si Satanas Satanan eicit adversus se divisus est quomodo ergo stabit regnum eius
MATT|12|27|et si ego in Beelzebub eicio daemones filii vestri in quo eiciunt ideo ipsi iudices erunt vestri
MATT|12|28|si autem ego in Spiritu Dei eicio daemones igitur pervenit in vos regnum Dei
MATT|12|29|aut quomodo potest quisquam intrare in domum fortis et vasa eius diripere nisi prius alligaverit fortem et tunc domum illius diripiat
MATT|12|30|qui non est mecum contra me est et qui non congregat mecum spargit
MATT|12|31|ideo dico vobis omne peccatum et blasphemia remittetur hominibus Spiritus autem blasphemia non remittetur
MATT|12|32|et quicumque dixerit verbum contra Filium hominis remittetur ei qui autem dixerit contra Spiritum Sanctum non remittetur ei neque in hoc saeculo neque in futuro
MATT|12|33|aut facite arborem bonam et fructum eius bonum aut facite arborem malam et fructum eius malum siquidem ex fructu arbor agnoscitur
MATT|12|34|progenies viperarum quomodo potestis bona loqui cum sitis mali ex abundantia enim cordis os loquitur
MATT|12|35|bonus homo de bono thesauro profert bona et malus homo de malo thesauro profert mala
MATT|12|36|dico autem vobis quoniam omne verbum otiosum quod locuti fuerint homines reddent rationem de eo in die iudicii
MATT|12|37|ex verbis enim tuis iustificaberis et ex verbis tuis condemnaberis
MATT|12|38|tunc responderunt ei quidam de scribis et Pharisaeis dicentes magister volumus a te signum videre
MATT|12|39|qui respondens ait illis generatio mala et adultera signum quaerit et signum non dabitur ei nisi signum Ionae prophetae
MATT|12|40|sicut enim fuit Ionas in ventre ceti tribus diebus et tribus noctibus sic erit Filius hominis in corde terrae tribus diebus et tribus noctibus
MATT|12|41|viri ninevitae surgent in iudicio cum generatione ista et condemnabunt eam quia paenitentiam egerunt in praedicatione Ionae et ecce plus quam Iona hic
MATT|12|42|regina austri surget in iudicio cum generatione ista et condemnabit eam quia venit a finibus terrae audire sapientiam Salomonis et ecce plus quam Salomon hic
MATT|12|43|cum autem inmundus spiritus exierit ab homine ambulat per loca arida quaerens requiem et non invenit
MATT|12|44|tunc dicit revertar in domum meam unde exivi et veniens invenit vacantem scopis mundatam et ornatam
MATT|12|45|tunc vadit et adsumit septem alios spiritus secum nequiores se et intrantes habitant ibi et fiunt novissima hominis illius peiora prioribus sic erit et generationi huic pessimae
MATT|12|46|adhuc eo loquente ad turbas ecce mater eius et fratres stabant foris quaerentes loqui ei
MATT|12|47|dixit autem ei quidam ecce mater tua et fratres tui foris stant quaerentes te
MATT|12|48|at ipse respondens dicenti sibi ait quae est mater mea et qui sunt fratres mei
MATT|12|49|et extendens manum in discipulos suos dixit ecce mater mea et fratres mei
MATT|12|50|quicumque enim fecerit voluntatem Patris mei qui in caelis est ipse meus et frater et soror et mater est
MATT|13|1|in illo die exiens Iesus de domo sedebat secus mare
MATT|13|2|et congregatae sunt ad eum turbae multae ita ut in naviculam ascendens sederet et omnis turba stabat in litore
MATT|13|3|et locutus est eis multa in parabolis dicens ecce exiit qui seminat seminare
MATT|13|4|et dum seminat quaedam ceciderunt secus viam et venerunt volucres et comederunt ea
MATT|13|5|alia autem ceciderunt in petrosa ubi non habebat terram multam et continuo exorta sunt quia non habebant altitudinem terrae
MATT|13|6|sole autem orto aestuaverunt et quia non habebant radicem aruerunt
MATT|13|7|alia autem ceciderunt in spinas et creverunt spinae et suffocaverunt ea
MATT|13|8|alia vero ceciderunt in terram bonam et dabant fructum aliud centesimum aliud sexagesimum aliud tricesimum
MATT|13|9|qui habet aures audiendi audiat
MATT|13|10|et accedentes discipuli dixerunt ei quare in parabolis loqueris eis
MATT|13|11|qui respondens ait illis quia vobis datum est nosse mysteria regni caelorum illis autem non est datum
MATT|13|12|qui enim habet dabitur ei et abundabit qui autem non habet et quod habet auferetur ab eo
MATT|13|13|ideo in parabolis loquor eis quia videntes non vident et audientes non audiunt neque intellegunt
MATT|13|14|et adimpletur eis prophetia Esaiae dicens auditu audietis et non intellegetis et videntes videbitis et non videbitis
MATT|13|15|incrassatum est enim cor populi huius et auribus graviter audierunt et oculos suos cluserunt nequando oculis videant et auribus audiant et corde intellegant et convertantur et sanem eos
MATT|13|16|vestri autem beati oculi quia vident et aures vestrae quia audiunt
MATT|13|17|amen quippe dico vobis quia multi prophetae et iusti cupierunt videre quae videtis et non viderunt et audire quae auditis et non audierunt
MATT|13|18|vos ergo audite parabolam seminantis
MATT|13|19|omnis qui audit verbum regni et non intellegit venit malus et rapit quod seminatum est in corde eius hic est qui secus viam seminatus est
MATT|13|20|qui autem supra petrosa seminatus est hic est qui verbum audit et continuo cum gaudio accipit illud
MATT|13|21|non habet autem in se radicem sed est temporalis facta autem tribulatione et persecutione propter verbum continuo scandalizatur
MATT|13|22|qui autem est seminatus in spinis hic est qui verbum audit et sollicitudo saeculi istius et fallacia divitiarum suffocat verbum et sine fructu efficitur
MATT|13|23|qui vero in terra bona seminatus est hic est qui audit verbum et intellegit et fructum adfert et facit aliud quidem centum aliud autem sexaginta porro aliud triginta
MATT|13|24|aliam parabolam proposuit illis dicens simile factum est regnum caelorum homini qui seminavit bonum semen in agro suo
MATT|13|25|cum autem dormirent homines venit inimicus eius et superseminavit zizania in medio tritici et abiit
MATT|13|26|cum autem crevisset herba et fructum fecisset tunc apparuerunt et zizania
MATT|13|27|accedentes autem servi patris familias dixerunt ei domine nonne bonum semen seminasti in agro tuo unde ergo habet zizania
MATT|13|28|et ait illis inimicus homo hoc fecit servi autem dixerunt ei vis imus et colligimus ea
MATT|13|29|et ait non ne forte colligentes zizania eradicetis simul cum eis et triticum
MATT|13|30|sinite utraque crescere usque ad messem et in tempore messis dicam messoribus colligite primum zizania et alligate ea fasciculos ad conburendum triticum autem congregate in horreum meum
MATT|13|31|aliam parabolam proposuit eis dicens simile est regnum caelorum grano sinapis quod accipiens homo seminavit in agro suo
MATT|13|32|quod minimum quidem est omnibus seminibus cum autem creverit maius est omnibus holeribus et fit arbor ita ut volucres caeli veniant et habitent in ramis eius
MATT|13|33|aliam parabolam locutus est eis simile est regnum caelorum fermento quod acceptum mulier abscondit in farinae satis tribus donec fermentatum est totum
MATT|13|34|haec omnia locutus est Iesus in parabolis ad turbas et sine parabolis non loquebatur eis
MATT|13|35|ut impleretur quod dictum erat per prophetam dicentem aperiam in parabolis os meum eructabo abscondita a constitutione mundi
MATT|13|36|tunc dimissis turbis venit in domum et accesserunt ad eum discipuli eius dicentes dissere nobis parabolam zizaniorum agri
MATT|13|37|qui respondens ait qui seminat bonum semen est Filius hominis
MATT|13|38|ager autem est mundus bonum vero semen hii sunt filii regni zizania autem filii sunt nequam
MATT|13|39|inimicus autem qui seminavit ea est diabolus messis vero consummatio saeculi est messores autem angeli sunt
MATT|13|40|sicut ergo colliguntur zizania et igni conburuntur sic erit in consummatione saeculi
MATT|13|41|mittet Filius hominis angelos suos et colligent de regno eius omnia scandala et eos qui faciunt iniquitatem
MATT|13|42|et mittent eos in caminum ignis ibi erit fletus et stridor dentium
MATT|13|43|tunc iusti fulgebunt sicut sol in regno Patris eorum qui habet aures audiat
MATT|13|44|simile est regnum caelorum thesauro abscondito in agro quem qui invenit homo abscondit et prae gaudio illius vadit et vendit universa quae habet et emit agrum illum
MATT|13|45|iterum simile est regnum caelorum homini negotiatori quaerenti bonas margaritas
MATT|13|46|inventa autem una pretiosa margarita abiit et vendidit omnia quae habuit et emit eam
MATT|13|47|iterum simile est regnum caelorum sagenae missae in mare et ex omni genere congreganti
MATT|13|48|quam cum impleta esset educentes et secus litus sedentes elegerunt bonos in vasa malos autem foras miserunt
MATT|13|49|sic erit in consummatione saeculi exibunt angeli et separabunt malos de medio iustorum
MATT|13|50|et mittent eos in caminum ignis ibi erit fletus et stridor dentium
MATT|13|51|intellexistis haec omnia dicunt ei etiam
MATT|13|52|ait illis ideo omnis scriba doctus in regno caelorum similis est homini patri familias qui profert de thesauro suo nova et vetera
MATT|13|53|et factum est cum consummasset Iesus parabolas istas transiit inde
MATT|13|54|et veniens in patriam suam docebat eos in synagogis eorum ita ut mirarentur et dicerent unde huic sapientia haec et virtutes
MATT|13|55|nonne hic est fabri filius nonne mater eius dicitur Maria et fratres eius Iacobus et Ioseph et Simon et Iudas
MATT|13|56|et sorores eius nonne omnes apud nos sunt unde ergo huic omnia ista
MATT|13|57|et scandalizabantur in eo Iesus autem dixit eis non est propheta sine honore nisi in patria sua et in domo sua
MATT|13|58|et non fecit ibi virtutes multas propter incredulitatem illorum
MATT|14|1|in illo tempore audiit Herodes tetrarcha famam Iesu
MATT|14|2|et ait pueris suis hic est Iohannes Baptista ipse surrexit a mortuis et ideo virtutes inoperantur in eo
MATT|14|3|Herodes enim tenuit Iohannem et alligavit eum et posuit in carcere propter Herodiadem uxorem fratris sui
MATT|14|4|dicebat enim illi Iohannes non licet tibi habere eam
MATT|14|5|et volens illum occidere timuit populum quia sicut prophetam eum habebant
MATT|14|6|die autem natalis Herodis saltavit filia Herodiadis in medio et placuit Herodi
MATT|14|7|unde cum iuramento pollicitus est ei dare quodcumque postulasset ab eo
MATT|14|8|at illa praemonita a matre sua da mihi inquit hic in disco caput Iohannis Baptistae
MATT|14|9|et contristatus est rex propter iuramentum autem et eos qui pariter recumbebant iussit dari
MATT|14|10|misitque et decollavit Iohannem in carcere
MATT|14|11|et adlatum est caput eius in disco et datum est puellae et tulit matri suae
MATT|14|12|et accedentes discipuli eius tulerunt corpus et sepelierunt illud et venientes nuntiaverunt Iesu
MATT|14|13|quod cum audisset Iesus secessit inde in navicula in locum desertum seorsum et cum audissent turbae secutae sunt eum pedestres de civitatibus
MATT|14|14|et exiens vidit turbam multam et misertus est eius et curavit languidos eorum
MATT|14|15|vespere autem facto accesserunt ad eum discipuli eius dicentes desertus est locus et hora iam praeteriit dimitte turbas ut euntes in castella emant sibi escas
MATT|14|16|Iesus autem dixit eis non habent necesse ire date illis vos manducare
MATT|14|17|responderunt ei non habemus hic nisi quinque panes et duos pisces
MATT|14|18|qui ait eis adferte illos mihi huc
MATT|14|19|et cum iussisset turbam discumbere supra faenum acceptis quinque panibus et duobus piscibus aspiciens in caelum benedixit et fregit et dedit discipulis panes discipuli autem turbis
MATT|14|20|et manducaverunt omnes et saturati sunt et tulerunt reliquias duodecim cofinos fragmentorum plenos
MATT|14|21|manducantium autem fuit numerus quinque milia virorum exceptis mulieribus et parvulis
MATT|14|22|et statim iussit discipulos ascendere in navicula et praecedere eum trans fretum donec dimitteret turbas
MATT|14|23|et dimissa turba ascendit in montem solus orare vespere autem facto solus erat ibi
MATT|14|24|navicula autem in medio mari iactabatur fluctibus erat enim contrarius ventus
MATT|14|25|quarta autem vigilia noctis venit ad eos ambulans supra mare
MATT|14|26|et videntes eum supra mare ambulantem turbati sunt dicentes quia fantasma est et prae timore clamaverunt
MATT|14|27|statimque Iesus locutus est eis dicens habete fiduciam ego sum nolite timere
MATT|14|28|respondens autem Petrus dixit Domine si tu es iube me venire ad te super aquas
MATT|14|29|at ipse ait veni et descendens Petrus de navicula ambulabat super aquam ut veniret ad Iesum
MATT|14|30|videns vero ventum validum timuit et cum coepisset mergi clamavit dicens Domine salvum me fac
MATT|14|31|et continuo Iesus extendens manum adprehendit eum et ait illi modicae fidei quare dubitasti
MATT|14|32|et cum ascendissent in naviculam cessavit ventus
MATT|14|33|qui autem in navicula erant venerunt et adoraverunt eum dicentes vere Filius Dei es
MATT|14|34|et cum transfretassent venerunt in terram Gennesar
MATT|14|35|et cum cognovissent eum viri loci illius miserunt in universam regionem illam et obtulerunt ei omnes male habentes
MATT|14|36|et rogabant eum ut vel fimbriam vestimenti eius tangerent et quicumque tetigerunt salvi facti sunt
MATT|15|1|tunc accesserunt ad eum ab Hierosolymis scribae et Pharisaei dicentes
MATT|15|2|quare discipuli tui transgrediuntur traditionem seniorum non enim lavant manus suas cum panem manducant
MATT|15|3|ipse autem respondens ait illis quare et vos transgredimini mandatum Dei propter traditionem vestram
MATT|15|4|nam Deus dixit honora patrem et matrem et qui maledixerit patri vel matri morte moriatur
MATT|15|5|vos autem dicitis quicumque dixerit patri vel matri munus quodcumque est ex me tibi proderit
MATT|15|6|et non honorificabit patrem suum aut matrem et irritum fecistis mandatum Dei propter traditionem vestram
MATT|15|7|hypocritae bene prophetavit de vobis Esaias dicens
MATT|15|8|populus hic labiis me honorat cor autem eorum longe est a me
MATT|15|9|sine causa autem colunt me docentes doctrinas mandata hominum
MATT|15|10|et convocatis ad se turbis dixit eis audite et intellegite
MATT|15|11|non quod intrat in os coinquinat hominem sed quod procedit ex ore hoc coinquinat hominem
MATT|15|12|tunc accedentes discipuli eius dixerunt ei scis quia Pharisaei audito verbo scandalizati sunt
MATT|15|13|at ille respondens ait omnis plantatio quam non plantavit Pater meus caelestis eradicabitur
MATT|15|14|sinite illos caeci sunt duces caecorum caecus autem si caeco ducatum praestet ambo in foveam cadunt
MATT|15|15|respondens autem Petrus dixit ei edissere nobis parabolam istam
MATT|15|16|at ille dixit adhuc et vos sine intellectu estis
MATT|15|17|non intellegitis quia omne quod in os intrat in ventrem vadit et in secessum emittitur
MATT|15|18|quae autem procedunt de ore de corde exeunt et ea coinquinant hominem
MATT|15|19|de corde enim exeunt cogitationes malae homicidia adulteria fornicationes furta falsa testimonia blasphemiae
MATT|15|20|haec sunt quae coinquinant hominem non lotis autem manibus manducare non coinquinat hominem
MATT|15|21|et egressus inde Iesus secessit in partes Tyri et Sidonis
MATT|15|22|et ecce mulier chananea a finibus illis egressa clamavit dicens ei miserere mei Domine Fili David filia mea male a daemonio vexatur
MATT|15|23|qui non respondit ei verbum et accedentes discipuli eius rogabant eum dicentes dimitte eam quia clamat post nos
MATT|15|24|ipse autem respondens ait non sum missus nisi ad oves quae perierunt domus Israhel
MATT|15|25|at illa venit et adoravit eum dicens Domine adiuva me
MATT|15|26|qui respondens ait non est bonum sumere panem filiorum et mittere canibus
MATT|15|27|at illa dixit etiam Domine nam et catelli edunt de micis quae cadunt de mensa dominorum suorum
MATT|15|28|tunc respondens Iesus ait illi o mulier magna est fides tua fiat tibi sicut vis et sanata est filia illius ex illa hora
MATT|15|29|et cum transisset inde Iesus venit secus mare Galilaeae et ascendens in montem sedebat ibi
MATT|15|30|et accesserunt ad eum turbae multae habentes secum mutos clodos caecos debiles et alios multos et proiecerunt eos ad pedes eius et curavit eos
MATT|15|31|ita ut turbae mirarentur videntes mutos loquentes clodos ambulantes caecos videntes et magnificabant Deum Israhel
MATT|15|32|Iesus autem convocatis discipulis suis dixit misereor turbae quia triduo iam perseverant mecum et non habent quod manducent et dimittere eos ieiunos nolo ne deficiant in via
MATT|15|33|et dicunt ei discipuli unde ergo nobis in deserto panes tantos ut saturemus turbam tantam
MATT|15|34|et ait illis Iesus quot panes habetis at illi dixerunt septem et paucos pisciculos
MATT|15|35|et praecepit turbae ut discumberet super terram
MATT|15|36|et accipiens septem panes et pisces et gratias agens fregit et dedit discipulis suis et discipuli dederunt populo
MATT|15|37|et comederunt omnes et saturati sunt et quod superfuit de fragmentis tulerunt septem sportas plenas
MATT|15|38|erant autem qui manducaverant quattuor milia hominum extra parvulos et mulieres
MATT|15|39|et dimissa turba ascendit in naviculam et venit in fines Magedan
MATT|16|1|et accesserunt ad eum Pharisaei et Sadducaei temptantes et rogaverunt eum ut signum de caelo ostenderet eis
MATT|16|2|at ille respondens ait eis facto vespere dicitis serenum erit rubicundum est enim caelum
MATT|16|3|et mane hodie tempestas rutilat enim triste caelum
MATT|16|4|faciem ergo caeli diiudicare nostis signa autem temporum non potestis generatio mala et adultera signum quaerit et signum non dabitur ei nisi signum Ionae et relictis illis abiit
MATT|16|5|et cum venissent discipuli eius trans fretum obliti sunt panes accipere
MATT|16|6|qui dixit illis intuemini et cavete a fermento Pharisaeorum et Sadducaeorum
MATT|16|7|at illi cogitabant inter se dicentes quia panes non accepimus
MATT|16|8|sciens autem Iesus dixit quid cogitatis inter vos modicae fidei quia panes non habetis
MATT|16|9|nondum intellegitis neque recordamini quinque panum quinque milium hominum et quot cofinos sumpsistis
MATT|16|10|neque septem panum quattuor milium hominum et quot sportas sumpsistis
MATT|16|11|quare non intellegitis quia non de pane dixi vobis cavete a fermento Pharisaeorum et Sadducaeorum
MATT|16|12|tunc intellexerunt quia non dixerit cavendum a fermento panum sed a doctrina Pharisaeorum et Sadducaeorum
MATT|16|13|venit autem Iesus in partes Caesareae Philippi et interrogabat discipulos suos dicens quem dicunt homines esse Filium hominis
MATT|16|14|at illi dixerunt alii Iohannem Baptistam alii autem Heliam alii vero Hieremiam aut unum ex prophetis
MATT|16|15|dicit illis vos autem quem me esse dicitis
MATT|16|16|respondens Simon Petrus dixit tu es Christus Filius Dei vivi
MATT|16|17|respondens autem Iesus dixit ei beatus es Simon Bar Iona quia caro et sanguis non revelavit tibi sed Pater meus qui in caelis est
MATT|16|18|et ego dico tibi quia tu es Petrus et super hanc petram aedificabo ecclesiam meam et portae inferi non praevalebunt adversum eam
MATT|16|19|et tibi dabo claves regni caelorum et quodcumque ligaveris super terram erit ligatum in caelis et quodcumque solveris super terram erit solutum in caelis
MATT|16|20|tunc praecepit discipulis suis ut nemini dicerent quia ipse esset Iesus Christus
MATT|16|21|exinde coepit Iesus ostendere discipulis suis quia oporteret eum ire Hierosolymam et multa pati a senioribus et scribis et principibus sacerdotum et occidi et tertia die resurgere
MATT|16|22|et adsumens eum Petrus coepit increpare illum dicens absit a te Domine non erit tibi hoc
MATT|16|23|qui conversus dixit Petro vade post me Satana scandalum es mihi quia non sapis ea quae Dei sunt sed ea quae hominum
MATT|16|24|tunc Iesus dixit discipulis suis si quis vult post me venire abneget semet ipsum et tollat crucem suam et sequatur me
MATT|16|25|qui enim voluerit animam suam salvam facere perdet eam qui autem perdiderit animam suam propter me inveniet eam
MATT|16|26|quid enim prodest homini si mundum universum lucretur animae vero suae detrimentum patiatur aut quam dabit homo commutationem pro anima sua
MATT|16|27|Filius enim hominis venturus est in gloria Patris sui cum angelis suis et tunc reddet unicuique secundum opus eius
MATT|16|28|amen dico vobis sunt quidam de hic stantibus qui non gustabunt mortem donec videant Filium hominis venientem in regno suo
MATT|17|1|et post dies sex adsumpsit Iesus Petrum et Iacobum et Iohannem fratrem eius et ducit illos in montem excelsum seorsum
MATT|17|2|et transfiguratus est ante eos et resplenduit facies eius sicut sol vestimenta autem eius facta sunt alba sicut nix
MATT|17|3|et ecce apparuit illis Moses et Helias cum eo loquentes
MATT|17|4|respondens autem Petrus dixit ad Iesum Domine bonum est nos hic esse si vis faciamus hic tria tabernacula tibi unum et Mosi unum et Heliae unum
MATT|17|5|adhuc eo loquente ecce nubes lucida obumbravit eos et ecce vox de nube dicens hic est Filius meus dilectus in quo mihi bene conplacuit ipsum audite
MATT|17|6|et audientes discipuli ceciderunt in faciem suam et timuerunt valde
MATT|17|7|et accessit Iesus et tetigit eos dixitque eis surgite et nolite timere
MATT|17|8|levantes autem oculos suos neminem viderunt nisi solum Iesum
MATT|17|9|et descendentibus illis de monte praecepit Iesus dicens nemini dixeritis visionem donec Filius hominis a mortuis resurgat
MATT|17|10|et interrogaverunt eum discipuli dicentes quid ergo scribae dicunt quod Heliam oporteat primum venire
MATT|17|11|at ille respondens ait eis Helias quidem venturus est et restituet omnia
MATT|17|12|dico autem vobis quia Helias iam venit et non cognoverunt eum sed fecerunt in eo quaecumque voluerunt sic et Filius hominis passurus est ab eis
MATT|17|13|tunc intellexerunt discipuli quia de Iohanne Baptista dixisset eis
MATT|17|14|et cum venisset ad turbam accessit ad eum homo genibus provolutus ante eum dicens Domine miserere filii mei quia lunaticus est et male patitur nam saepe cadit in ignem et crebro in aquam
MATT|17|15|et obtuli eum discipulis tuis et non potuerunt curare eum
MATT|17|16|respondens Iesus ait o generatio incredula et perversa quousque ero vobiscum usquequo patiar vos adferte huc illum ad me
MATT|17|17|et increpavit ei Iesus et exiit ab eo daemonium et curatus est puer ex illa hora
MATT|17|18|tunc accesserunt discipuli ad Iesum secreto et dixerunt quare nos non potuimus eicere illum
MATT|17|19|dicit illis propter incredulitatem vestram amen quippe dico vobis si habueritis fidem sicut granum sinapis dicetis monti huic transi hinc et transibit et nihil inpossibile erit vobis
MATT|17|20|hoc autem genus non eicitur nisi per orationem et ieiunium
MATT|17|21|conversantibus autem eis in Galilaea dixit illis Iesus Filius hominis tradendus est in manus hominum
MATT|17|22|et occident eum et tertio die resurget et contristati sunt vehementer
MATT|17|23|et cum venissent Capharnaum accesserunt qui didragma accipiebant ad Petrum et dixerunt magister vester non solvit didragma
MATT|17|24|ait etiam et cum intrasset domum praevenit eum Iesus dicens quid tibi videtur Simon reges terrae a quibus accipiunt tributum vel censum a filiis suis an ab alienis
MATT|17|25|et ille dixit ab alienis dixit illi Iesus ergo liberi sunt filii
MATT|17|26|ut autem non scandalizemus eos vade ad mare et mitte hamum et eum piscem qui primus ascenderit tolle et aperto ore eius invenies staterem illum sumens da eis pro me et te
MATT|17|27|
MATT|18|1|in illa hora accesserunt discipuli ad Iesum dicentes quis putas maior est in regno caelorum
MATT|18|2|et advocans Iesus parvulum statuit eum in medio eorum
MATT|18|3|et dixit amen dico vobis nisi conversi fueritis et efficiamini sicut parvuli non intrabitis in regnum caelorum
MATT|18|4|quicumque ergo humiliaverit se sicut parvulus iste hic est maior in regno caelorum
MATT|18|5|et qui susceperit unum parvulum talem in nomine meo me suscipit
MATT|18|6|qui autem scandalizaverit unum de pusillis istis qui in me credunt expedit ei ut suspendatur mola asinaria in collo eius et demergatur in profundum maris
MATT|18|7|vae mundo ab scandalis necesse est enim ut veniant scandala verumtamen vae homini per quem scandalum venit
MATT|18|8|si autem manus tua vel pes tuus scandalizat te abscide eum et proice abs te bonum tibi est ad vitam ingredi debilem vel clodum quam duas manus vel duos pedes habentem mitti in ignem aeternum
MATT|18|9|et si oculus tuus scandalizat te erue eum et proice abs te bonum tibi est unoculum in vitam intrare quam duos oculos habentem mitti in gehennam ignis
MATT|18|10|videte ne contemnatis unum ex his pusillis dico enim vobis quia angeli eorum in caelis semper vident faciem Patris mei qui in caelis est
MATT|18|11|venit enim Filius hominis salvare quod perierat
MATT|18|12|quid vobis videtur si fuerint alicui centum oves et erraverit una ex eis nonne relinquet nonaginta novem in montibus et vadit quaerere eam quae erravit
MATT|18|13|et si contigerit ut inveniat eam amen dico vobis quia gaudebit super eam magis quam super nonaginta novem quae non erraverunt
MATT|18|14|sic non est voluntas ante Patrem vestrum qui in caelis est ut pereat unus de pusillis istis
MATT|18|15|si autem peccaverit in te frater tuus vade et corripe eum inter te et ipsum solum si te audierit lucratus es fratrem tuum
MATT|18|16|si autem non te audierit adhibe tecum adhuc unum vel duos ut in ore duorum testium vel trium stet omne verbum
MATT|18|17|quod si non audierit eos dic ecclesiae si autem et ecclesiam non audierit sit tibi sicut ethnicus et publicanus
MATT|18|18|amen dico vobis quaecumque alligaveritis super terram erunt ligata et in caelo et quaecumque solveritis super terram erunt soluta et in caelo
MATT|18|19|iterum dico vobis quia si duo ex vobis consenserint super terram de omni re quacumque petierint fiet illis a Patre meo qui in caelis est
MATT|18|20|ubi enim sunt duo vel tres congregati in nomine meo ibi sum in medio eorum
MATT|18|21|tunc accedens Petrus ad eum dixit Domine quotiens peccabit in me frater meus et dimittam ei usque septies
MATT|18|22|dicit illi Iesus non dico tibi usque septies sed usque septuagies septies
MATT|18|23|ideo adsimilatum est regnum caelorum homini regi qui voluit rationem ponere cum servis suis
MATT|18|24|et cum coepisset rationem ponere oblatus est ei unus qui debebat decem milia talenta
MATT|18|25|cum autem non haberet unde redderet iussit eum dominus venundari et uxorem eius et filios et omnia quae habebat et reddi
MATT|18|26|procidens autem servus ille orabat eum dicens patientiam habe in me et omnia reddam tibi
MATT|18|27|misertus autem dominus servi illius dimisit eum et debitum dimisit ei
MATT|18|28|egressus autem servus ille invenit unum de conservis suis qui debebat ei centum denarios et tenens suffocabat eum dicens redde quod debes
MATT|18|29|et procidens conservus eius rogabat eum dicens patientiam habe in me et omnia reddam tibi
MATT|18|30|ille autem noluit sed abiit et misit eum in carcerem donec redderet debitum
MATT|18|31|videntes autem conservi eius quae fiebant contristati sunt valde et venerunt et narraverunt domino suo omnia quae facta erant
MATT|18|32|tunc vocavit illum dominus suus et ait illi serve nequam omne debitum dimisi tibi quoniam rogasti me
MATT|18|33|non ergo oportuit et te misereri conservi tui sicut et ego tui misertus sum
MATT|18|34|et iratus dominus eius tradidit eum tortoribus quoadusque redderet universum debitum
MATT|18|35|sic et Pater meus caelestis faciet vobis si non remiseritis unusquisque fratri suo de cordibus vestris
MATT|19|1|et factum est cum consummasset Iesus sermones istos migravit a Galilaea et venit in fines Iudaeae trans Iordanen
MATT|19|2|et secutae sunt eum turbae multae et curavit eos ibi
MATT|19|3|et accesserunt ad eum Pharisaei temptantes eum et dicentes si licet homini dimittere uxorem suam quacumque ex causa
MATT|19|4|qui respondens ait eis non legistis quia qui fecit ab initio masculum et feminam fecit eos
MATT|19|5|et dixit propter hoc dimittet homo patrem et matrem et adherebit uxori suae et erunt duo in carne una
MATT|19|6|itaque iam non sunt duo sed una caro quod ergo Deus coniunxit homo non separet
MATT|19|7|dicunt illi quid ergo Moses mandavit dari libellum repudii et dimittere
MATT|19|8|ait illis quoniam Moses ad duritiam cordis vestri permisit vobis dimittere uxores vestras ab initio autem non sic fuit
MATT|19|9|dico autem vobis quia quicumque dimiserit uxorem suam nisi ob fornicationem et aliam duxerit moechatur et qui dimissam duxerit moechatur
MATT|19|10|dicunt ei discipuli eius si ita est causa homini cum uxore non expedit nubere
MATT|19|11|qui dixit non omnes capiunt verbum istud sed quibus datum est
MATT|19|12|sunt enim eunuchi qui de matris utero sic nati sunt et sunt eunuchi qui facti sunt ab hominibus et sunt eunuchi qui se ipsos castraverunt propter regnum caelorum qui potest capere capiat
MATT|19|13|tunc oblati sunt ei parvuli ut manus eis inponeret et oraret discipuli autem increpabant eis
MATT|19|14|Iesus vero ait eis sinite parvulos et nolite eos prohibere ad me venire talium est enim regnum caelorum
MATT|19|15|et cum inposuisset eis manus abiit inde
MATT|19|16|et ecce unus accedens ait illi magister bone quid boni faciam ut habeam vitam aeternam
MATT|19|17|qui dixit ei quid me interrogas de bono unus est bonus Deus si autem vis ad vitam ingredi serva mandata
MATT|19|18|dicit illi quae Iesus autem dixit non homicidium facies non adulterabis non facies furtum non falsum testimonium dices
MATT|19|19|honora patrem et matrem et diliges proximum tuum sicut te ipsum
MATT|19|20|dicit illi adulescens omnia haec custodivi quid adhuc mihi deest
MATT|19|21|ait illi Iesus si vis perfectus esse vade vende quae habes et da pauperibus et habebis thesaurum in caelo et veni sequere me
MATT|19|22|cum audisset autem adulescens verbum abiit tristis erat enim habens multas possessiones
MATT|19|23|Iesus autem dixit discipulis suis amen dico vobis quia dives difficile intrabit in regnum caelorum
MATT|19|24|et iterum dico vobis facilius est camelum per foramen acus transire quam divitem intrare in regnum caelorum
MATT|19|25|auditis autem his discipuli mirabantur valde dicentes quis ergo poterit salvus esse
MATT|19|26|aspiciens autem Iesus dixit illis apud homines hoc inpossibile est apud Deum autem omnia possibilia sunt
MATT|19|27|tunc respondens Petrus dixit ei ecce nos reliquimus omnia et secuti sumus te quid ergo erit nobis
MATT|19|28|Iesus autem dixit illis amen dico vobis quod vos qui secuti estis me in regeneratione cum sederit Filius hominis in sede maiestatis suae sedebitis et vos super sedes duodecim iudicantes duodecim tribus Israhel
MATT|19|29|et omnis qui reliquit domum vel fratres aut sorores aut patrem aut matrem aut uxorem aut filios aut agros propter nomen meum centuplum accipiet et vitam aeternam possidebit
MATT|19|30|multi autem erunt primi novissimi et novissimi primi
MATT|20|1|simile est enim regnum caelorum homini patri familias qui exiit primo mane conducere operarios in vineam suam
MATT|20|2|conventione autem facta cum operariis ex denario diurno misit eos in vineam suam
MATT|20|3|et egressus circa horam tertiam vidit alios stantes in foro otiosos
MATT|20|4|et illis dixit ite et vos in vineam et quod iustum fuerit dabo vobis
MATT|20|5|illi autem abierunt iterum autem exiit circa sextam et nonam horam et fecit similiter
MATT|20|6|circa undecimam vero exiit et invenit alios stantes et dicit illis quid hic statis tota die otiosi
MATT|20|7|dicunt ei quia nemo nos conduxit dicit illis ite et vos in vineam
MATT|20|8|cum sero autem factum esset dicit dominus vineae procuratori suo voca operarios et redde illis mercedem incipiens a novissimis usque ad primos
MATT|20|9|cum venissent ergo qui circa undecimam horam venerant acceperunt singulos denarios
MATT|20|10|venientes autem et primi arbitrati sunt quod plus essent accepturi acceperunt autem et ipsi singulos denarios
MATT|20|11|et accipientes murmurabant adversus patrem familias
MATT|20|12|dicentes hii novissimi una hora fecerunt et pares illos nobis fecisti qui portavimus pondus diei et aestus
MATT|20|13|at ille respondens uni eorum dixit amice non facio tibi iniuriam nonne ex denario convenisti mecum
MATT|20|14|tolle quod tuum est et vade volo autem et huic novissimo dare sicut et tibi
MATT|20|15|aut non licet mihi quod volo facere an oculus tuus nequam est quia ego bonus sum
MATT|20|16|sic erunt novissimi primi et primi novissimi multi sunt enim vocati pauci autem electi
MATT|20|17|et ascendens Iesus Hierosolymam adsumpsit duodecim discipulos secreto et ait illis
MATT|20|18|ecce ascendimus Hierosolymam et Filius hominis tradetur principibus sacerdotum et scribis et condemnabunt eum morte
MATT|20|19|et tradent eum gentibus ad deludendum et flagellandum et crucifigendum et tertia die resurget
MATT|20|20|tunc accessit ad eum mater filiorum Zebedaei cum filiis suis adorans et petens aliquid ab eo
MATT|20|21|qui dixit ei quid vis ait illi dic ut sedeant hii duo filii mei unus ad dexteram tuam et unus ad sinistram in regno tuo
MATT|20|22|respondens autem Iesus dixit nescitis quid petatis potestis bibere calicem quem ego bibiturus sum dicunt ei possumus
MATT|20|23|ait illis calicem quidem meum bibetis sedere autem ad dexteram meam et sinistram non est meum dare vobis sed quibus paratum est a Patre meo
MATT|20|24|et audientes decem indignati sunt de duobus fratribus
MATT|20|25|Iesus autem vocavit eos ad se et ait scitis quia principes gentium dominantur eorum et qui maiores sunt potestatem exercent in eos
MATT|20|26|non ita erit inter vos sed quicumque voluerit inter vos maior fieri sit vester minister
MATT|20|27|et qui voluerit inter vos primus esse erit vester servus
MATT|20|28|sicut Filius hominis non venit ministrari sed ministrare et dare animam suam redemptionem pro multis
MATT|20|29|et egredientibus eis ab Hiericho secuta est eum turba multa
MATT|20|30|et ecce duo caeci sedentes secus viam audierunt quia Iesus transiret et clamaverunt dicentes Domine miserere nostri Fili David
MATT|20|31|turba autem increpabat eos ut tacerent at illi magis clamabant dicentes Domine miserere nostri Fili David
MATT|20|32|et stetit Iesus et vocavit eos et ait quid vultis ut faciam vobis
MATT|20|33|dicunt illi Domine ut aperiantur oculi nostri
MATT|20|34|misertus autem eorum Iesus tetigit oculos eorum et confestim viderunt et secuti sunt eum
MATT|21|1|et cum adpropinquassent Hierosolymis et venissent Bethfage ad montem Oliveti tunc Iesus misit duos discipulos
MATT|21|2|dicens eis ite in castellum quod contra vos est et statim invenietis asinam alligatam et pullum cum ea solvite et adducite mihi
MATT|21|3|et si quis vobis aliquid dixerit dicite quia Dominus his opus habet et confestim dimittet eos
MATT|21|4|hoc autem factum est ut impleretur quod dictum est per prophetam dicentem
MATT|21|5|dicite filiae Sion ecce rex tuus venit tibi mansuetus et sedens super asinam et pullum filium subiugalis
MATT|21|6|euntes autem discipuli fecerunt sicut praecepit illis Iesus
MATT|21|7|et adduxerunt asinam et pullum et inposuerunt super eis vestimenta sua et eum desuper sedere fecerunt
MATT|21|8|plurima autem turba straverunt vestimenta sua in via alii autem caedebant ramos de arboribus et sternebant in via
MATT|21|9|turbae autem quae praecedebant et quae sequebantur clamabant dicentes osanna Filio David benedictus qui venturus est in nomine Domini osanna in altissimis
MATT|21|10|et cum intrasset Hierosolymam commota est universa civitas dicens quis est hic
MATT|21|11|populi autem dicebant hic est Iesus propheta a Nazareth Galilaeae
MATT|21|12|et intravit Iesus in templum Dei et eiciebat omnes vendentes et ementes in templo et mensas nummulariorum et cathedras vendentium columbas evertit
MATT|21|13|et dicit eis scriptum est domus mea domus orationis vocabitur vos autem fecistis eam speluncam latronum
MATT|21|14|et accesserunt ad eum caeci et claudi in templo et sanavit eos
MATT|21|15|videntes autem principes sacerdotum et scribae mirabilia quae fecit et pueros clamantes in templo et dicentes osanna Filio David indignati sunt
MATT|21|16|et dixerunt ei audis quid isti dicant Iesus autem dicit eis utique numquam legistis quia ex ore infantium et lactantium perfecisti laudem
MATT|21|17|et relictis illis abiit foras extra civitatem in Bethaniam ibique mansit
MATT|21|18|mane autem revertens in civitatem esuriit
MATT|21|19|et videns fici arborem unam secus viam venit ad eam et nihil invenit in ea nisi folia tantum et ait illi numquam ex te fructus nascatur in sempiternum et arefacta est continuo ficulnea
MATT|21|20|et videntes discipuli mirati sunt dicentes quomodo continuo aruit
MATT|21|21|respondens autem Iesus ait eis amen dico vobis si habueritis fidem et non haesitaveritis non solum de ficulnea facietis sed et si monti huic dixeritis tolle et iacta te in mare fiet
MATT|21|22|et omnia quaecumque petieritis in oratione credentes accipietis
MATT|21|23|et cum venisset in templum accesserunt ad eum docentem principes sacerdotum et seniores populi dicentes in qua potestate haec facis et quis tibi dedit hanc potestatem
MATT|21|24|respondens Iesus dixit illis interrogabo vos et ego unum sermonem quem si dixeritis mihi et ego vobis dicam in qua potestate haec facio
MATT|21|25|baptismum Iohannis unde erat e caelo an ex hominibus at illi cogitabant inter se dicentes si dixerimus e caelo dicet nobis quare ergo non credidistis illi
MATT|21|26|si autem dixerimus ex hominibus timemus turbam omnes enim habent Iohannem sicut prophetam
MATT|21|27|et respondentes Iesu dixerunt nescimus ait illis et ipse nec ego dico vobis in qua potestate haec facio
MATT|21|28|quid autem vobis videtur homo habebat duos filios et accedens ad primum dixit fili vade hodie operare in vinea mea
MATT|21|29|ille autem respondens ait nolo postea autem paenitentia motus abiit
MATT|21|30|accedens autem ad alterum dixit similiter at ille respondens ait eo domine et non ivit
MATT|21|31|quis ex duobus fecit voluntatem patris dicunt novissimus dicit illis Iesus amen dico vobis quia publicani et meretrices praecedunt vos in regno Dei
MATT|21|32|venit enim ad vos Iohannes in via iustitiae et non credidistis ei publicani autem et meretrices crediderunt ei vos autem videntes nec paenitentiam habuistis postea ut crederetis ei
MATT|21|33|aliam parabolam audite homo erat pater familias qui plantavit vineam et sepem circumdedit ei et fodit in ea torcular et aedificavit turrem et locavit eam agricolis et peregre profectus est
MATT|21|34|cum autem tempus fructuum adpropinquasset misit servos suos ad agricolas ut acciperent fructus eius
MATT|21|35|et agricolae adprehensis servis eius alium ceciderunt alium occiderunt alium vero lapidaverunt
MATT|21|36|iterum misit alios servos plures prioribus et fecerunt illis similiter
MATT|21|37|novissime autem misit ad eos filium suum dicens verebuntur filium meum
MATT|21|38|agricolae autem videntes filium dixerunt intra se hic est heres venite occidamus eum et habebimus hereditatem eius
MATT|21|39|et adprehensum eum eiecerunt extra vineam et occiderunt
MATT|21|40|cum ergo venerit dominus vineae quid faciet agricolis illis
MATT|21|41|aiunt illi malos male perdet et vineam locabit aliis agricolis qui reddant ei fructum temporibus suis
MATT|21|42|dicit illis Iesus numquam legistis in scripturis lapidem quem reprobaverunt aedificantes hic factus est in caput anguli a Domino factum est istud et est mirabile in oculis nostris
MATT|21|43|ideo dico vobis quia auferetur a vobis regnum Dei et dabitur genti facienti fructus eius
MATT|21|44|et qui ceciderit super lapidem istum confringetur super quem vero ceciderit conteret eum
MATT|21|45|et cum audissent principes sacerdotum et Pharisaei parabolas eius cognoverunt quod de ipsis diceret
MATT|21|46|et quaerentes eum tenere timuerunt turbas quoniam sicut prophetam eum habebant
MATT|22|1|et respondens Iesus dixit iterum in parabolis eis dicens
MATT|22|2|simile factum est regnum caelorum homini regi qui fecit nuptias filio suo
MATT|22|3|et misit servos suos vocare invitatos ad nuptias et nolebant venire
MATT|22|4|iterum misit alios servos dicens dicite invitatis ecce prandium meum paravi tauri mei et altilia occisa et omnia parata venite ad nuptias
MATT|22|5|illi autem neglexerunt et abierunt alius in villam suam alius vero ad negotiationem suam
MATT|22|6|reliqui vero tenuerunt servos eius et contumelia adfectos occiderunt
MATT|22|7|rex autem cum audisset iratus est et missis exercitibus suis perdidit homicidas illos et civitatem illorum succendit
MATT|22|8|tunc ait servis suis nuptiae quidem paratae sunt sed qui invitati erant non fuerunt digni
MATT|22|9|ite ergo ad exitus viarum et quoscumque inveneritis vocate ad nuptias
MATT|22|10|et egressi servi eius in vias congregaverunt omnes quos invenerunt malos et bonos et impletae sunt nuptiae discumbentium
MATT|22|11|intravit autem rex ut videret discumbentes et vidit ibi hominem non vestitum veste nuptiali
MATT|22|12|et ait illi amice quomodo huc intrasti non habens vestem nuptialem at ille obmutuit
MATT|22|13|tunc dixit rex ministris ligatis pedibus eius et manibus mittite eum in tenebras exteriores ibi erit fletus et stridor dentium
MATT|22|14|multi autem sunt vocati pauci vero electi
MATT|22|15|tunc abeuntes Pharisaei consilium inierunt ut caperent eum in sermone
MATT|22|16|et mittunt ei discipulos suos cum Herodianis dicentes magister scimus quia verax es et viam Dei in veritate doces et non est tibi cura de aliquo non enim respicis personam hominum
MATT|22|17|dic ergo nobis quid tibi videatur licet censum dare Caesari an non
MATT|22|18|cognita autem Iesus nequitia eorum ait quid me temptatis hypocritae
MATT|22|19|ostendite mihi nomisma census at illi obtulerunt ei denarium
MATT|22|20|et ait illis Iesus cuius est imago haec et suprascriptio
MATT|22|21|dicunt ei Caesaris tunc ait illis reddite ergo quae sunt Caesaris Caesari et quae sunt Dei Deo
MATT|22|22|et audientes mirati sunt et relicto eo abierunt
MATT|22|23|in illo die accesserunt ad eum Sadducaei qui dicunt non esse resurrectionem et interrogaverunt eum
MATT|22|24|dicentes magister Moses dixit si quis mortuus fuerit non habens filium ut ducat frater eius uxorem illius et suscitet semen fratri suo
MATT|22|25|erant autem apud nos septem fratres et primus uxore ducta defunctus est et non habens semen reliquit uxorem suam fratri suo
MATT|22|26|similiter secundus et tertius usque ad septimum
MATT|22|27|novissime autem omnium et mulier defuncta est
MATT|22|28|in resurrectione ergo cuius erit de septem uxor omnes enim habuerunt eam
MATT|22|29|respondens autem Iesus ait illis erratis nescientes scripturas neque virtutem Dei
MATT|22|30|in resurrectione enim neque nubent neque nubentur sed sunt sicut angeli Dei in caelo
MATT|22|31|de resurrectione autem mortuorum non legistis quod dictum est a Deo dicente vobis
MATT|22|32|ego sum Deus Abraham et Deus Isaac et Deus Iacob non est Deus mortuorum sed viventium
MATT|22|33|et audientes turbae mirabantur in doctrina eius
MATT|22|34|Pharisaei autem audientes quod silentium inposuisset Sadducaeis convenerunt in unum
MATT|22|35|et interrogavit eum unus ex eis legis doctor temptans eum
MATT|22|36|magister quod est mandatum magnum in lege
MATT|22|37|ait illi Iesus diliges Dominum Deum tuum ex toto corde tuo et in tota anima tua et in tota mente tua
MATT|22|38|hoc est maximum et primum mandatum
MATT|22|39|secundum autem simile est huic diliges proximum tuum sicut te ipsum
MATT|22|40|in his duobus mandatis universa lex pendet et prophetae
MATT|22|41|congregatis autem Pharisaeis interrogavit eos Iesus
MATT|22|42|dicens quid vobis videtur de Christo cuius filius est dicunt ei David
MATT|22|43|ait illis quomodo ergo David in spiritu vocat eum Dominum dicens
MATT|22|44|dixit Dominus Domino meo sede a dextris meis donec ponam inimicos tuos scabillum pedum tuorum
MATT|22|45|si ergo David vocat eum Dominum quomodo filius eius est
MATT|22|46|et nemo poterat respondere ei verbum neque ausus fuit quisquam ex illa die eum amplius interrogare
MATT|23|1|tunc Iesus locutus est ad turbas et discipulos suos
MATT|23|2|dicens super cathedram Mosi sederunt scribae et Pharisaei
MATT|23|3|omnia ergo quaecumque dixerint vobis servate et facite secundum opera vero eorum nolite facere dicunt enim et non faciunt
MATT|23|4|alligant autem onera gravia et inportabilia et inponunt in umeros hominum digito autem suo nolunt ea movere
MATT|23|5|omnia vero opera sua faciunt ut videantur ab hominibus dilatant enim phylacteria sua et magnificant fimbrias
MATT|23|6|amant autem primos recubitus in cenis et primas cathedras in synagogis
MATT|23|7|et salutationes in foro et vocari ab hominibus rabbi
MATT|23|8|vos autem nolite vocari rabbi unus enim est magister vester omnes autem vos fratres estis
MATT|23|9|et patrem nolite vocare vobis super terram unus enim est Pater vester qui in caelis est
MATT|23|10|nec vocemini magistri quia magister vester unus est Christus
MATT|23|11|qui maior est vestrum erit minister vester
MATT|23|12|qui autem se exaltaverit humiliabitur et qui se humiliaverit exaltabitur
MATT|23|13|vae autem vobis scribae et Pharisaei hypocritae quia clauditis regnum caelorum ante homines vos enim non intratis nec introeuntes sinitis intrare
MATT|23|14|
MATT|23|15|vae vobis scribae et Pharisaei hypocritae quia circuitis mare et aridam ut faciatis unum proselytum et cum fuerit factus facitis eum filium gehennae duplo quam vos
MATT|23|16|vae vobis duces caeci qui dicitis quicumque iuraverit per templum nihil est qui autem iuraverit in aurum templi debet
MATT|23|17|stulti et caeci quid enim maius est aurum an templum quod sanctificat aurum
MATT|23|18|et quicumque iuraverit in altari nihil est quicumque autem iuraverit in dono quod est super illud debet
MATT|23|19|caeci quid enim maius est donum an altare quod sanctificat donum
MATT|23|20|qui ergo iurat in altare iurat in eo et in omnibus quae super illud sunt
MATT|23|21|et qui iuraverit in templo iurat in illo et in eo qui inhabitat in ipso
MATT|23|22|et qui iurat in caelo iurat in throno Dei et in eo qui sedet super eum
MATT|23|23|vae vobis scribae et Pharisaei hypocritae quia decimatis mentam et anethum et cyminum et reliquistis quae graviora sunt legis iudicium et misericordiam et fidem haec oportuit facere et illa non omittere
MATT|23|24|duces caeci excolantes culicem camelum autem gluttientes
MATT|23|25|vae vobis scribae et Pharisaei hypocritae quia mundatis quod de foris est calicis et parapsidis intus autem pleni sunt rapina et inmunditia
MATT|23|26|Pharisaee caece munda prius quod intus est calicis et parapsidis ut fiat et id quod de foris est mundum
MATT|23|27|vae vobis scribae et Pharisaei hypocritae quia similes estis sepulchris dealbatis quae a foris parent hominibus speciosa intus vero plena sunt ossibus mortuorum et omni spurcitia
MATT|23|28|sic et vos a foris quidem paretis hominibus iusti intus autem pleni estis hypocrisi et iniquitate
MATT|23|29|vae vobis scribae et Pharisaei hypocritae quia aedificatis sepulchra prophetarum et ornatis monumenta iustorum
MATT|23|30|et dicitis si fuissemus in diebus patrum nostrorum non essemus socii eorum in sanguine prophetarum
MATT|23|31|itaque testimonio estis vobismet ipsis quia filii estis eorum qui prophetas occiderunt
MATT|23|32|et vos implete mensuram patrum vestrorum
MATT|23|33|serpentes genimina viperarum quomodo fugietis a iudicio gehennae
MATT|23|34|ideo ecce ego mitto ad vos prophetas et sapientes et scribas ex illis occidetis et crucifigetis et ex eis flagellabitis in synagogis vestris et persequemini de civitate in civitatem
MATT|23|35|ut veniat super vos omnis sanguis iustus qui effusus est super terram a sanguine Abel iusti usque ad sanguinem Zacchariae filii Barachiae quem occidistis inter templum et altare
MATT|23|36|amen dico vobis venient haec omnia super generationem istam
MATT|23|37|Hierusalem Hierusalem quae occidis prophetas et lapidas eos qui ad te missi sunt quotiens volui congregare filios tuos quemadmodum gallina congregat pullos suos sub alas et noluisti
MATT|23|38|ecce relinquitur vobis domus vestra deserta
MATT|23|39|dico enim vobis non me videbitis amodo donec dicatis benedictus qui venit in nomine Domini
MATT|24|1|et egressus Iesus de templo ibat et accesserunt discipuli eius ut ostenderent ei aedificationes templi
MATT|24|2|ipse autem respondens dixit eis videtis haec omnia amen dico vobis non relinquetur hic lapis super lapidem qui non destruatur
MATT|24|3|sedente autem eo super montem Oliveti accesserunt ad eum discipuli secreto dicentes dic nobis quando haec erunt et quod signum adventus tui et consummationis saeculi
MATT|24|4|et respondens Iesus dixit eis videte ne quis vos seducat
MATT|24|5|multi enim venient in nomine meo dicentes ego sum Christus et multos seducent
MATT|24|6|audituri autem estis proelia et opiniones proeliorum videte ne turbemini oportet enim haec fieri sed nondum est finis
MATT|24|7|consurget enim gens in gentem et regnum in regnum et erunt pestilentiae et fames et terraemotus per loca
MATT|24|8|haec autem omnia initia sunt dolorum
MATT|24|9|tunc tradent vos in tribulationem et occident vos et eritis odio omnibus gentibus propter nomen meum
MATT|24|10|et tunc scandalizabuntur multi et invicem tradent et odio habebunt invicem
MATT|24|11|et multi pseudoprophetae surgent et seducent multos
MATT|24|12|et quoniam abundabit iniquitas refrigescet caritas multorum
MATT|24|13|qui autem permanserit usque in finem hic salvus erit
MATT|24|14|et praedicabitur hoc evangelium regni in universo orbe in testimonium omnibus gentibus et tunc veniet consummatio
MATT|24|15|cum ergo videritis abominationem desolationis quae dicta est a Danihelo propheta stantem in loco sancto qui legit intellegat
MATT|24|16|tunc qui in Iudaea sunt fugiant ad montes
MATT|24|17|et qui in tecto non descendat tollere aliquid de domo sua
MATT|24|18|et qui in agro non revertatur tollere tunicam suam
MATT|24|19|vae autem praegnatibus et nutrientibus in illis diebus
MATT|24|20|orate autem ut non fiat fuga vestra hieme vel sabbato
MATT|24|21|erit enim tunc tribulatio magna qualis non fuit ab initio mundi usque modo neque fiet
MATT|24|22|et nisi breviati fuissent dies illi non fieret salva omnis caro sed propter electos breviabuntur dies illi
MATT|24|23|tunc si quis vobis dixerit ecce hic Christus aut illic nolite credere
MATT|24|24|surgent enim pseudochristi et pseudoprophetae et dabunt signa magna et prodigia ita ut in errorem inducantur si fieri potest etiam electi
MATT|24|25|ecce praedixi vobis
MATT|24|26|si ergo dixerint vobis ecce in deserto est nolite exire ecce in penetrabilibus nolite credere
MATT|24|27|sicut enim fulgur exit ab oriente et paret usque in occidente ita erit et adventus Filii hominis
MATT|24|28|ubicumque fuerit corpus illuc congregabuntur aquilae
MATT|24|29|statim autem post tribulationem dierum illorum sol obscurabitur et luna non dabit lumen suum et stellae cadent de caelo et virtutes caelorum commovebuntur
MATT|24|30|et tunc parebit signum Filii hominis in caelo et tunc plangent omnes tribus terrae et videbunt Filium hominis venientem in nubibus caeli cum virtute multa et maiestate
MATT|24|31|et mittet angelos suos cum tuba et voce magna et congregabunt electos eius a quattuor ventis a summis caelorum usque ad terminos eorum
MATT|24|32|ab arbore autem fici discite parabolam cum iam ramus eius tener fuerit et folia nata scitis quia prope est aestas
MATT|24|33|ita et vos cum videritis haec omnia scitote quia prope est in ianuis
MATT|24|34|amen dico vobis quia non praeteribit haec generatio donec omnia haec fiant
MATT|24|35|caelum et terra transibunt verba vero mea non praeteribunt
MATT|24|36|de die autem illa et hora nemo scit neque angeli caelorum nisi Pater solus
MATT|24|37|sicut autem in diebus Noe ita erit et adventus Filii hominis
MATT|24|38|sicut enim erant in diebus ante diluvium comedentes et bibentes nubentes et nuptum tradentes usque ad eum diem quo introivit in arcam Noe
MATT|24|39|et non cognoverunt donec venit diluvium et tulit omnes ita erit et adventus Filii hominis
MATT|24|40|tunc duo erunt in agro unus adsumetur et unus relinquetur
MATT|24|41|duae molentes in mola una adsumetur et una relinquetur
MATT|24|42|vigilate ergo quia nescitis qua hora Dominus vester venturus sit
MATT|24|43|illud autem scitote quoniam si sciret pater familias qua hora fur venturus esset vigilaret utique et non sineret perfodiri domum suam
MATT|24|44|ideoque et vos estote parati quia qua nescitis hora Filius hominis venturus est
MATT|24|45|quis putas est fidelis servus et prudens quem constituit dominus suus supra familiam suam ut det illis cibum in tempore
MATT|24|46|beatus ille servus quem cum venerit dominus eius invenerit sic facientem
MATT|24|47|amen dico vobis quoniam super omnia bona sua constituet eum
MATT|24|48|si autem dixerit malus servus ille in corde suo moram facit dominus meus venire
MATT|24|49|et coeperit percutere conservos suos manducet autem et bibat cum ebriis
MATT|24|50|veniet dominus servi illius in die qua non sperat et hora qua ignorat
MATT|24|51|et dividet eum partemque eius ponet cum hypocritis illic erit fletus et stridor dentium
MATT|25|1|tunc simile erit regnum caelorum decem virginibus quae accipientes lampadas suas exierunt obviam sponso et sponsae
MATT|25|2|quinque autem ex eis erant fatuae et quinque prudentes
MATT|25|3|sed quinque fatuae acceptis lampadibus non sumpserunt oleum secum
MATT|25|4|prudentes vero acceperunt oleum in vasis suis cum lampadibus
MATT|25|5|moram autem faciente sponso dormitaverunt omnes et dormierunt
MATT|25|6|media autem nocte clamor factus est ecce sponsus venit exite obviam ei
MATT|25|7|tunc surrexerunt omnes virgines illae et ornaverunt lampades suas
MATT|25|8|fatuae autem sapientibus dixerunt date nobis de oleo vestro quia lampades nostrae extinguntur
MATT|25|9|responderunt prudentes dicentes ne forte non sufficiat nobis et vobis ite potius ad vendentes et emite vobis
MATT|25|10|dum autem irent emere venit sponsus et quae paratae erant intraverunt cum eo ad nuptias et clausa est ianua
MATT|25|11|novissime veniunt et reliquae virgines dicentes domine domine aperi nobis
MATT|25|12|at ille respondens ait amen dico vobis nescio vos
MATT|25|13|vigilate itaque quia nescitis diem neque horam
MATT|25|14|sicut enim homo proficiscens vocavit servos suos et tradidit illis bona sua
MATT|25|15|et uni dedit quinque talenta alii autem duo alii vero unum unicuique secundum propriam virtutem et profectus est statim
MATT|25|16|abiit autem qui quinque talenta acceperat et operatus est in eis et lucratus est alia quinque
MATT|25|17|similiter qui duo acceperat lucratus est alia duo
MATT|25|18|qui autem unum acceperat abiens fodit in terra et abscondit pecuniam domini sui
MATT|25|19|post multum vero temporis venit dominus servorum illorum et posuit rationem cum eis
MATT|25|20|et accedens qui quinque talenta acceperat obtulit alia quinque talenta dicens domine quinque talenta mihi tradidisti ecce alia quinque superlucratus sum
MATT|25|21|ait illi dominus eius euge bone serve et fidelis quia super pauca fuisti fidelis super multa te constituam intra in gaudium domini tui
MATT|25|22|accessit autem et qui duo talenta acceperat et ait domine duo talenta tradidisti mihi ecce alia duo lucratus sum
MATT|25|23|ait illi dominus eius euge serve bone et fidelis quia super pauca fuisti fidelis supra multa te constituam intra in gaudium domini tui
MATT|25|24|accedens autem et qui unum talentum acceperat ait domine scio quia homo durus es metis ubi non seminasti et congregas ubi non sparsisti
MATT|25|25|et timens abii et abscondi talentum tuum in terra ecce habes quod tuum est
MATT|25|26|respondens autem dominus eius dixit ei serve male et piger sciebas quia meto ubi non semino et congrego ubi non sparsi
MATT|25|27|oportuit ergo te mittere pecuniam meam nummulariis et veniens ego recepissem utique quod meum est cum usura
MATT|25|28|tollite itaque ab eo talentum et date ei qui habet decem talenta
MATT|25|29|omni enim habenti dabitur et abundabit ei autem qui non habet et quod videtur habere auferetur ab eo
MATT|25|30|et inutilem servum eicite in tenebras exteriores illic erit fletus et stridor dentium
MATT|25|31|cum autem venerit Filius hominis in maiestate sua et omnes angeli cum eo tunc sedebit super sedem maiestatis suae
MATT|25|32|et congregabuntur ante eum omnes gentes et separabit eos ab invicem sicut pastor segregat oves ab hedis
MATT|25|33|et statuet oves quidem a dextris suis hedos autem a sinistris
MATT|25|34|tunc dicet rex his qui a dextris eius erunt venite benedicti Patris mei possidete paratum vobis regnum a constitutione mundi
MATT|25|35|esurivi enim et dedistis mihi manducare sitivi et dedistis mihi bibere hospes eram et collexistis me
MATT|25|36|nudus et operuistis me infirmus et visitastis me in carcere eram et venistis ad me
MATT|25|37|tunc respondebunt ei iusti dicentes Domine quando te vidimus esurientem et pavimus sitientem et dedimus tibi potum
MATT|25|38|quando autem te vidimus hospitem et colleximus te aut nudum et cooperuimus
MATT|25|39|aut quando te vidimus infirmum aut in carcere et venimus ad te
MATT|25|40|et respondens rex dicet illis amen dico vobis quamdiu fecistis uni de his fratribus meis minimis mihi fecistis
MATT|25|41|tunc dicet et his qui a sinistris erunt discedite a me maledicti in ignem aeternum qui paratus est diabolo et angelis eius
MATT|25|42|esurivi enim et non dedistis mihi manducare sitivi et non dedistis mihi potum
MATT|25|43|hospes eram et non collexistis me nudus et non operuistis me infirmus et in carcere et non visitastis me
MATT|25|44|tunc respondebunt et ipsi dicentes Domine quando te vidimus esurientem aut sitientem aut hospitem aut nudum aut infirmum vel in carcere et non ministravimus tibi
MATT|25|45|tunc respondebit illis dicens amen dico vobis quamdiu non fecistis uni de minoribus his nec mihi fecistis
MATT|25|46|et ibunt hii in supplicium aeternum iusti autem in vitam aeternam
MATT|26|1|et factum est cum consummasset Iesus sermones hos omnes dixit discipulis suis
MATT|26|2|scitis quia post biduum pascha fiet et Filius hominis tradetur ut crucifigatur
MATT|26|3|tunc congregati sunt principes sacerdotum et seniores populi in atrium principis sacerdotum qui dicebatur Caiaphas
MATT|26|4|et consilium fecerunt ut Iesum dolo tenerent et occiderent
MATT|26|5|dicebant autem non in die festo ne forte tumultus fieret in populo
MATT|26|6|cum autem esset Iesus in Bethania in domo Simonis leprosi
MATT|26|7|accessit ad eum mulier habens alabastrum unguenti pretiosi et effudit super caput ipsius recumbentis
MATT|26|8|videntes autem discipuli indignati sunt dicentes ut quid perditio haec
MATT|26|9|potuit enim istud venundari multo et dari pauperibus
MATT|26|10|sciens autem Iesus ait illis quid molesti estis mulieri opus bonum operata est in me
MATT|26|11|nam semper pauperes habetis vobiscum me autem non semper habetis
MATT|26|12|mittens enim haec unguentum hoc in corpus meum ad sepeliendum me fecit
MATT|26|13|amen dico vobis ubicumque praedicatum fuerit hoc evangelium in toto mundo dicetur et quod haec fecit in memoriam eius
MATT|26|14|tunc abiit unus de duodecim qui dicitur Iudas Scarioth ad principes sacerdotum
MATT|26|15|et ait illis quid vultis mihi dare et ego vobis eum tradam at illi constituerunt ei triginta argenteos
MATT|26|16|et exinde quaerebat oportunitatem ut eum traderet
MATT|26|17|prima autem azymorum accesserunt discipuli ad Iesum dicentes ubi vis paremus tibi comedere pascha
MATT|26|18|at Iesus dixit ite in civitatem ad quendam et dicite ei magister dicit tempus meum prope est apud te facio pascha cum discipulis meis
MATT|26|19|et fecerunt discipuli sicut constituit illis Iesus et paraverunt pascha
MATT|26|20|vespere autem facto discumbebat cum duodecim discipulis
MATT|26|21|et edentibus illis dixit amen dico vobis quia unus vestrum me traditurus est
MATT|26|22|et contristati valde coeperunt singuli dicere numquid ego sum Domine
MATT|26|23|at ipse respondens ait qui intinguit mecum manum in parapside hic me tradet
MATT|26|24|Filius quidem hominis vadit sicut scriptum est de illo vae autem homini illi per quem Filius hominis traditur bonum erat ei si natus non fuisset homo ille
MATT|26|25|respondens autem Iudas qui tradidit eum dixit numquid ego sum rabbi ait illi tu dixisti
MATT|26|26|cenantibus autem eis accepit Iesus panem et benedixit ac fregit deditque discipulis suis et ait accipite et comedite hoc est corpus meum
MATT|26|27|et accipiens calicem gratias egit et dedit illis dicens bibite ex hoc omnes
MATT|26|28|hic est enim sanguis meus novi testamenti qui pro multis effunditur in remissionem peccatorum
MATT|26|29|dico autem vobis non bibam amodo de hoc genimine vitis usque in diem illum cum illud bibam vobiscum novum in regno Patris mei
MATT|26|30|et hymno dicto exierunt in montem Oliveti
MATT|26|31|tunc dicit illis Iesus omnes vos scandalum patiemini in me in ista nocte scriptum est enim percutiam pastorem et dispergentur oves gregis
MATT|26|32|postquam autem resurrexero praecedam vos in Galilaeam
MATT|26|33|respondens autem Petrus ait illi et si omnes scandalizati fuerint in te ego numquam scandalizabor
MATT|26|34|ait illi Iesus amen dico tibi quia in hac nocte antequam gallus cantet ter me negabis
MATT|26|35|ait illi Petrus etiam si oportuerit me mori tecum non te negabo similiter et omnes discipuli dixerunt
MATT|26|36|tunc venit Iesus cum illis in villam quae dicitur Gethsemani et dixit discipulis suis sedete hic donec vadam illuc et orem
MATT|26|37|et adsumpto Petro et duobus filiis Zebedaei coepit contristari et maestus esse
MATT|26|38|tunc ait illis tristis est anima mea usque ad mortem sustinete hic et vigilate mecum
MATT|26|39|et progressus pusillum procidit in faciem suam orans et dicens mi Pater si possibile est transeat a me calix iste verumtamen non sicut ego volo sed sicut tu
MATT|26|40|et venit ad discipulos et invenit eos dormientes et dicit Petro sic non potuistis una hora vigilare mecum
MATT|26|41|vigilate et orate ut non intretis in temptationem spiritus quidem promptus est caro autem infirma
MATT|26|42|iterum secundo abiit et oravit dicens Pater mi si non potest hic calix transire nisi bibam illum fiat voluntas tua
MATT|26|43|et venit iterum et invenit eos dormientes erant enim oculi eorum gravati
MATT|26|44|et relictis illis iterum abiit et oravit tertio eundem sermonem dicens
MATT|26|45|tunc venit ad discipulos suos et dicit illis dormite iam et requiescite ecce adpropinquavit hora et Filius hominis traditur in manus peccatorum
MATT|26|46|surgite eamus ecce adpropinquavit qui me tradit
MATT|26|47|adhuc ipso loquente ecce Iudas unus de duodecim venit et cum eo turba multa cum gladiis et fustibus a principibus sacerdotum et senioribus populi
MATT|26|48|qui autem tradidit eum dedit illis signum dicens quemcumque osculatus fuero ipse est tenete eum
MATT|26|49|et confestim accedens ad Iesum dixit have rabbi et osculatus est eum
MATT|26|50|dixitque illi Iesus amice ad quod venisti tunc accesserunt et manus iniecerunt in Iesum et tenuerunt eum
MATT|26|51|et ecce unus ex his qui erant cum Iesu extendens manum exemit gladium suum et percutiens servum principis sacerdotum amputavit auriculam eius
MATT|26|52|tunc ait illi Iesus converte gladium tuum in locum suum omnes enim qui acceperint gladium gladio peribunt
MATT|26|53|an putas quia non possum rogare Patrem meum et exhibebit mihi modo plus quam duodecim legiones angelorum
MATT|26|54|quomodo ergo implebuntur scripturae quia sic oportet fieri
MATT|26|55|in illa hora dixit Iesus turbis tamquam ad latronem existis cum gladiis et fustibus conprehendere me cotidie apud vos sedebam docens in templo et non me tenuistis
MATT|26|56|hoc autem totum factum est ut implerentur scripturae prophetarum tunc discipuli omnes relicto eo fugerunt
MATT|26|57|at illi tenentes Iesum duxerunt ad Caiaphan principem sacerdotum ubi scribae et seniores convenerant
MATT|26|58|Petrus autem sequebatur eum a longe usque in atrium principis sacerdotum et ingressus intro sedebat cum ministris ut videret finem
MATT|26|59|principes autem sacerdotum et omne concilium quaerebant falsum testimonium contra Iesum ut eum morti traderent
MATT|26|60|et non invenerunt cum multi falsi testes accessissent novissime autem venerunt duo falsi testes
MATT|26|61|et dixerunt hic dixit possum destruere templum Dei et post triduum aedificare illud
MATT|26|62|et surgens princeps sacerdotum ait illi nihil respondes ad ea quae isti adversum te testificantur
MATT|26|63|Iesus autem tacebat et princeps sacerdotum ait illi adiuro te per Deum vivum ut dicas nobis si tu es Christus Filius Dei
MATT|26|64|dicit illi Iesus tu dixisti verumtamen dico vobis amodo videbitis Filium hominis sedentem a dextris virtutis et venientem in nubibus caeli
MATT|26|65|tunc princeps sacerdotum scidit vestimenta sua dicens blasphemavit quid adhuc egemus testibus ecce nunc audistis blasphemiam
MATT|26|66|quid vobis videtur at illi respondentes dixerunt reus est mortis
MATT|26|67|tunc expuerunt in faciem eius et colaphis eum ceciderunt alii autem palmas in faciem ei dederunt
MATT|26|68|dicentes prophetiza nobis Christe quis est qui te percussit
MATT|26|69|Petrus vero sedebat foris in atrio et accessit ad eum una ancilla dicens et tu cum Iesu Galilaeo eras
MATT|26|70|at ille negavit coram omnibus dicens nescio quid dicis
MATT|26|71|exeunte autem illo ianuam vidit eum alia et ait his qui erant ibi et hic erat cum Iesu Nazareno
MATT|26|72|et iterum negavit cum iuramento quia non novi hominem
MATT|26|73|et post pusillum accesserunt qui stabant et dixerunt Petro vere et tu ex illis es nam et loquella tua manifestum te facit
MATT|26|74|tunc coepit detestari et iurare quia non novisset hominem et continuo gallus cantavit
MATT|26|75|et recordatus est Petrus verbi Iesu quod dixerat priusquam gallus cantet ter me negabis et egressus foras ploravit amare
MATT|27|1|mane autem facto consilium inierunt omnes principes sacerdotum et seniores populi adversus Iesum ut eum morti traderent
MATT|27|2|et vinctum adduxerunt eum et tradiderunt Pontio Pilato praesidi
MATT|27|3|tunc videns Iudas qui eum tradidit quod damnatus esset paenitentia ductus rettulit triginta argenteos principibus sacerdotum et senioribus
MATT|27|4|dicens peccavi tradens sanguinem iustum at illi dixerunt quid ad nos tu videris
MATT|27|5|et proiectis argenteis in templo recessit et abiens laqueo se suspendit
MATT|27|6|principes autem sacerdotum acceptis argenteis dixerunt non licet mittere eos in corbanan quia pretium sanguinis est
MATT|27|7|consilio autem inito emerunt ex illis agrum figuli in sepulturam peregrinorum
MATT|27|8|propter hoc vocatus est ager ille Acheldemach ager sanguinis usque in hodiernum diem
MATT|27|9|tunc impletum est quod dictum est per Hieremiam prophetam dicentem et acceperunt triginta argenteos pretium adpretiati quem adpretiaverunt a filiis Israhel
MATT|27|10|et dederunt eos in agrum figuli sicut constituit mihi Dominus
MATT|27|11|Iesus autem stetit ante praesidem et interrogavit eum praeses dicens tu es rex Iudaeorum dicit ei Iesus tu dicis
MATT|27|12|et cum accusaretur a principibus sacerdotum et senioribus nihil respondit
MATT|27|13|tunc dicit illi Pilatus non audis quanta adversum te dicant testimonia
MATT|27|14|et non respondit ei ad ullum verbum ita ut miraretur praeses vehementer
MATT|27|15|per diem autem sollemnem consueverat praeses dimittere populo unum vinctum quem voluissent
MATT|27|16|habebat autem tunc vinctum insignem qui dicebatur Barabbas
MATT|27|17|congregatis ergo illis dixit Pilatus quem vultis dimittam vobis Barabban an Iesum qui dicitur Christus
MATT|27|18|sciebat enim quod per invidiam tradidissent eum
MATT|27|19|sedente autem illo pro tribunali misit ad illum uxor eius dicens nihil tibi et iusto illi multa enim passa sum hodie per visum propter eum
MATT|27|20|princeps autem sacerdotum et seniores persuaserunt populis ut peterent Barabban Iesum vero perderent
MATT|27|21|respondens autem praeses ait illis quem vultis vobis de duobus dimitti at illi dixerunt Barabban
MATT|27|22|dicit illis Pilatus quid igitur faciam de Iesu qui dicitur Christus
MATT|27|23|dicunt omnes crucifigatur ait illis praeses quid enim mali fecit at illi magis clamabant dicentes crucifigatur
MATT|27|24|videns autem Pilatus quia nihil proficeret sed magis tumultus fieret accepta aqua lavit manus coram populo dicens innocens ego sum a sanguine iusti huius vos videritis
MATT|27|25|et respondens universus populus dixit sanguis eius super nos et super filios nostros
MATT|27|26|tunc dimisit illis Barabban Iesum autem flagellatum tradidit eis ut crucifigeretur
MATT|27|27|tunc milites praesidis suscipientes Iesum in praetorio congregaverunt ad eum universam cohortem
MATT|27|28|et exuentes eum clamydem coccineam circumdederunt ei
MATT|27|29|et plectentes coronam de spinis posuerunt super caput eius et harundinem in dextera eius et genu flexo ante eum inludebant dicentes have rex Iudaeorum
MATT|27|30|et expuentes in eum acceperunt harundinem et percutiebant caput eius
MATT|27|31|et postquam inluserunt ei exuerunt eum clamydem et induerunt eum vestimentis eius et duxerunt eum ut crucifigerent
MATT|27|32|exeuntes autem invenerunt hominem cyreneum nomine Simonem hunc angariaverunt ut tolleret crucem eius
MATT|27|33|et venerunt in locum qui dicitur Golgotha quod est Calvariae locus
MATT|27|34|et dederunt ei vinum bibere cum felle mixtum et cum gustasset noluit bibere
MATT|27|35|postquam autem crucifixerunt eum diviserunt vestimenta eius sortem mittentes
MATT|27|36|et sedentes servabant eum
MATT|27|37|et inposuerunt super caput eius causam ipsius scriptam hic est Iesus rex Iudaeorum
MATT|27|38|tunc crucifixi sunt cum eo duo latrones unus a dextris et unus a sinistris
MATT|27|39|praetereuntes autem blasphemabant eum moventes capita sua
MATT|27|40|et dicentes qui destruit templum et in triduo illud reaedificat salva temet ipsum si Filius Dei es descende de cruce
MATT|27|41|similiter et principes sacerdotum inludentes cum scribis et senioribus dicentes
MATT|27|42|alios salvos fecit se ipsum non potest salvum facere si rex Israhel est descendat nunc de cruce et credemus ei
MATT|27|43|confidet in Deo liberet nunc eum si vult dixit enim quia Dei Filius sum
MATT|27|44|id ipsum autem et latrones qui fixi erant cum eo inproperabant ei
MATT|27|45|a sexta autem hora tenebrae factae sunt super universam terram usque ad horam nonam
MATT|27|46|et circa horam nonam clamavit Iesus voce magna dicens Heli Heli lema sabacthani hoc est Deus meus Deus meus ut quid dereliquisti me
MATT|27|47|quidam autem illic stantes et audientes dicebant Heliam vocat iste
MATT|27|48|et continuo currens unus ex eis acceptam spongiam implevit aceto et inposuit harundini et dabat ei bibere
MATT|27|49|ceteri vero dicebant sine videamus an veniat Helias liberans eum
MATT|27|50|Iesus autem iterum clamans voce magna emisit spiritum
MATT|27|51|et ecce velum templi scissum est in duas partes a summo usque deorsum et terra mota est et petrae scissae sunt
MATT|27|52|et monumenta aperta sunt et multa corpora sanctorum qui dormierant surrexerunt
MATT|27|53|et exeuntes de monumentis post resurrectionem eius venerunt in sanctam civitatem et apparuerunt multis
MATT|27|54|centurio autem et qui cum eo erant custodientes Iesum viso terraemotu et his quae fiebant timuerunt valde dicentes vere Dei Filius erat iste
MATT|27|55|erant autem ibi mulieres multae a longe quae secutae erant Iesum a Galilaea ministrantes ei
MATT|27|56|inter quas erat Maria Magdalene et Maria Iacobi et Ioseph mater et mater filiorum Zebedaei
MATT|27|57|cum sero autem factum esset venit quidam homo dives ab Arimathia nomine Ioseph qui et ipse discipulus erat Iesu
MATT|27|58|hic accessit ad Pilatum et petiit corpus Iesu tunc Pilatus iussit reddi corpus
MATT|27|59|et accepto corpore Ioseph involvit illud sindone munda
MATT|27|60|et posuit illud in monumento suo novo quod exciderat in petra et advolvit saxum magnum ad ostium monumenti et abiit
MATT|27|61|erat autem ibi Maria Magdalene et altera Maria sedentes contra sepulchrum
MATT|27|62|altera autem die quae est post parasceven convenerunt principes sacerdotum et Pharisaei ad Pilatum
MATT|27|63|dicentes domine recordati sumus quia seductor ille dixit adhuc vivens post tres dies resurgam
MATT|27|64|iube ergo custodiri sepulchrum usque in diem tertium ne forte veniant discipuli eius et furentur eum et dicant plebi surrexit a mortuis et erit novissimus error peior priore
MATT|27|65|ait illis Pilatus habetis custodiam ite custodite sicut scitis
MATT|27|66|illi autem abeuntes munierunt sepulchrum signantes lapidem cum custodibus
MATT|28|1|vespere autem sabbati quae lucescit in primam sabbati venit Maria Magdalene et altera Maria videre sepulchrum
MATT|28|2|et ecce terraemotus factus est magnus angelus enim Domini descendit de caelo et accedens revolvit lapidem et sedebat super eum
MATT|28|3|erat autem aspectus eius sicut fulgur et vestimentum eius sicut nix
MATT|28|4|prae timore autem eius exterriti sunt custodes et facti sunt velut mortui
MATT|28|5|respondens autem angelus dixit mulieribus nolite timere vos scio enim quod Iesum qui crucifixus est quaeritis
MATT|28|6|non est hic surrexit enim sicut dixit venite videte locum ubi positus erat Dominus
MATT|28|7|et cito euntes dicite discipulis eius quia surrexit et ecce praecedit vos in Galilaeam ibi eum videbitis ecce praedixi vobis
MATT|28|8|et exierunt cito de monumento cum timore et magno gaudio currentes nuntiare discipulis eius
MATT|28|9|et ecce Iesus occurrit illis dicens havete illae autem accesserunt et tenuerunt pedes eius et adoraverunt eum
MATT|28|10|tunc ait illis Iesus nolite timere ite nuntiate fratribus meis ut eant in Galilaeam ibi me videbunt
MATT|28|11|quae cum abissent ecce quidam de custodibus venerunt in civitatem et nuntiaverunt principibus sacerdotum omnia quae facta fuerant
MATT|28|12|et congregati cum senioribus consilio accepto pecuniam copiosam dederunt militibus
MATT|28|13|dicentes dicite quia discipuli eius nocte venerunt et furati sunt eum nobis dormientibus
MATT|28|14|et si hoc auditum fuerit a praeside nos suadebimus ei et securos vos faciemus
MATT|28|15|at illi accepta pecunia fecerunt sicut erant docti et divulgatum est verbum istud apud Iudaeos usque in hodiernum diem
MATT|28|16|undecim autem discipuli abierunt in Galilaeam in montem ubi constituerat illis Iesus
MATT|28|17|et videntes eum adoraverunt quidam autem dubitaverunt
MATT|28|18|et accedens Iesus locutus est eis dicens data est mihi omnis potestas in caelo et in terra
MATT|28|19|euntes ergo docete omnes gentes baptizantes eos in nomine Patris et Filii et Spiritus Sancti
MATT|28|20|docentes eos servare omnia quaecumque mandavi vobis et ecce ego vobiscum sum omnibus diebus usque ad consummationem saeculi
MARK|1|1|initium evangelii Iesu Christi Filii Dei
MARK|1|2|sicut scriptum est in Esaia propheta ecce mitto angelum meum ante faciem tuam qui praeparabit viam tuam
MARK|1|3|vox clamantis in deserto parate viam Domini rectas facite semitas eius
MARK|1|4|fuit Iohannes in deserto baptizans et praedicans baptismum paenitentiae in remissionem peccatorum
MARK|1|5|et egrediebatur ad illum omnis Iudaeae regio et Hierosolymitae universi et baptizabantur ab illo in Iordane flumine confitentes peccata sua
MARK|1|6|et erat Iohannes vestitus pilis cameli et zona pellicia circa lumbos eius et lucustas et mel silvestre edebat
MARK|1|7|et praedicabat dicens venit fortior me post me cuius non sum dignus procumbens solvere corrigiam calciamentorum eius
MARK|1|8|ego baptizavi vos aqua ille vero baptizabit vos Spiritu Sancto
MARK|1|9|et factum est in diebus illis venit Iesus a Nazareth Galilaeae et baptizatus est in Iordane ab Iohanne
MARK|1|10|et statim ascendens de aqua vidit apertos caelos et Spiritum tamquam columbam descendentem et manentem in ipso
MARK|1|11|et vox facta est de caelis tu es Filius meus dilectus in te conplacui
MARK|1|12|et statim Spiritus expellit eum in desertum
MARK|1|13|et erat in deserto quadraginta diebus et quadraginta noctibus et temptabatur a Satana eratque cum bestiis et angeli ministrabant illi
MARK|1|14|postquam autem traditus est Iohannes venit Iesus in Galilaeam praedicans evangelium regni Dei
MARK|1|15|et dicens quoniam impletum est tempus et adpropinquavit regnum Dei paenitemini et credite evangelio
MARK|1|16|et praeteriens secus mare Galilaeae vidit Simonem et Andream fratrem eius mittentes retia in mare erant enim piscatores
MARK|1|17|et dixit eis Iesus venite post me et faciam vos fieri piscatores hominum
MARK|1|18|et protinus relictis retibus secuti sunt eum
MARK|1|19|et progressus inde pusillum vidit Iacobum Zebedaei et Iohannem fratrem eius et ipsos in navi conponentes retia
MARK|1|20|et statim vocavit illos et relicto patre suo Zebedaeo in navi cum mercennariis secuti sunt eum
MARK|1|21|et ingrediuntur Capharnaum et statim sabbatis ingressus synagogam docebat eos
MARK|1|22|et stupebant super doctrina eius erat enim docens eos quasi potestatem habens et non sicut scribae
MARK|1|23|et erat in synagoga eorum homo in spiritu inmundo et exclamavit
MARK|1|24|dicens quid nobis et tibi Iesu Nazarene venisti perdere nos scio qui sis Sanctus Dei
MARK|1|25|et comminatus est ei Iesus dicens obmutesce et exi de homine
MARK|1|26|et discerpens eum spiritus inmundus et exclamans voce magna exivit ab eo
MARK|1|27|et mirati sunt omnes ita ut conquirerent inter se dicentes quidnam est hoc quae doctrina haec nova quia in potestate et spiritibus inmundis imperat et oboediunt ei
MARK|1|28|et processit rumor eius statim in omnem regionem Galilaeae
MARK|1|29|et protinus egredientes de synagoga venerunt in domum Simonis et Andreae cum Iacobo et Iohanne
MARK|1|30|decumbebat autem socrus Simonis febricitans et statim dicunt ei de illa
MARK|1|31|et accedens elevavit eam adprehensa manu eius et continuo dimisit eam febris et ministrabat eis
MARK|1|32|vespere autem facto cum occidisset sol adferebant ad eum omnes male habentes et daemonia habentes
MARK|1|33|et erat omnis civitas congregata ad ianuam
MARK|1|34|et curavit multos qui vexabantur variis languoribus et daemonia multa eiciebat et non sinebat loqui ea quoniam sciebant eum
MARK|1|35|et diluculo valde surgens egressus abiit in desertum locum ibique orabat
MARK|1|36|et persecutus est eum Simon et qui cum illo erant
MARK|1|37|et cum invenissent eum dixerunt ei quia omnes quaerunt te
MARK|1|38|et ait illis eamus in proximos vicos et civitates ut et ibi praedicem ad hoc enim veni
MARK|1|39|et erat praedicans in synagogis eorum et omni Galilaea et daemonia eiciens
MARK|1|40|et venit ad eum leprosus deprecans eum et genu flexo dixit si vis potes me mundare
MARK|1|41|Iesus autem misertus eius extendit manum suam et tangens eum ait illi volo mundare
MARK|1|42|et cum dixisset statim discessit ab eo lepra et mundatus est
MARK|1|43|et comminatus ei statim eiecit illum
MARK|1|44|et dicit ei vide nemini dixeris sed vade ostende te principi sacerdotum et offer pro emundatione tua quae praecepit Moses in testimonium illis
MARK|1|45|at ille egressus coepit praedicare et diffamare sermonem ita ut iam non posset manifeste in civitatem introire sed foris in desertis locis esse et conveniebant ad eum undique
MARK|2|1|et iterum intravit Capharnaum post dies
MARK|2|2|et auditum est quod in domo esset et convenerunt multi ita ut non caperet neque ad ianuam et loquebatur eis verbum
MARK|2|3|et venerunt ferentes ad eum paralyticum qui a quattuor portabatur
MARK|2|4|et cum non possent offerre eum illi prae turba nudaverunt tectum ubi erat et patefacientes submiserunt grabattum in quo paralyticus iacebat
MARK|2|5|cum vidisset autem Iesus fidem illorum ait paralytico fili dimittuntur tibi peccata
MARK|2|6|erant autem illic quidam de scribis sedentes et cogitantes in cordibus suis
MARK|2|7|quid hic sic loquitur blasphemat quis potest dimittere peccata nisi solus Deus
MARK|2|8|quo statim cognito Iesus spiritu suo quia sic cogitarent intra se dicit illis quid ista cogitatis in cordibus vestris
MARK|2|9|quid est facilius dicere paralytico dimittuntur tibi peccata an dicere surge et tolle grabattum tuum et ambula
MARK|2|10|ut autem sciatis quia potestatem habet Filius hominis in terra dimittendi peccata ait paralytico
MARK|2|11|tibi dico surge tolle grabattum tuum et vade in domum tuam
MARK|2|12|et statim ille surrexit et sublato grabatto abiit coram omnibus ita ut admirarentur omnes et honorificarent Deum dicentes quia numquam sic vidimus
MARK|2|13|et egressus est rursus ad mare omnisque turba veniebat ad eum et docebat eos
MARK|2|14|et cum praeteriret vidit Levin Alphei sedentem ad teloneum et ait illi sequere me et surgens secutus est eum
MARK|2|15|et factum est cum accumberet in domo illius multi publicani et peccatores simul discumbebant cum Iesu et discipulis eius erant enim multi qui et sequebantur eum
MARK|2|16|et scribae et Pharisaei videntes quia manducaret cum peccatoribus et publicanis dicebant discipulis eius quare cum publicanis et peccatoribus manducat et bibit magister vester
MARK|2|17|hoc audito Iesus ait illis non necesse habent sani medicum sed qui male habent non enim veni vocare iustos sed peccatores
MARK|2|18|et erant discipuli Iohannis et Pharisaei ieiunantes et veniunt et dicunt illi cur discipuli Iohannis et Pharisaeorum ieiunant tui autem discipuli non ieiunant
MARK|2|19|et ait illis Iesus numquid possunt filii nuptiarum quamdiu sponsus cum illis est ieiunare quanto tempore habent secum sponsum non possunt ieiunare
MARK|2|20|venient autem dies cum auferetur ab eis sponsus et tunc ieiunabunt in illa die
MARK|2|21|nemo adsumentum panni rudis adsuit vestimento veteri alioquin aufert supplementum novum a veteri et maior scissura fit
MARK|2|22|et nemo mittit vinum novellum in utres veteres alioquin disrumpet vinum utres et vinum effunditur et utres peribunt sed vinum novum in utres novos mitti debet
MARK|2|23|et factum est iterum cum sabbatis ambularet per sata et discipuli eius coeperunt praegredi et vellere spicas
MARK|2|24|Pharisaei autem dicebant ei ecce quid faciunt sabbatis quod non licet
MARK|2|25|et ait illis numquam legistis quid fecerit David quando necessitatem habuit et esuriit ipse et qui cum eo erant
MARK|2|26|quomodo introiit in domum Dei sub Abiathar principe sacerdotum et panes propositionis manducavit quos non licet manducare nisi sacerdotibus et dedit eis qui cum eo erant
MARK|2|27|et dicebat eis sabbatum propter hominem factum est et non homo propter sabbatum
MARK|2|28|itaque dominus est Filius hominis etiam sabbati
MARK|3|1|et introivit iterum synagogam et erat ibi homo habens manum aridam
MARK|3|2|et observabant eum si sabbatis curaret ut accusarent illum
MARK|3|3|et ait homini habenti manum aridam surge in medium
MARK|3|4|et dicit eis licet sabbatis bene facere an male animam salvam facere an perdere at illi tacebant
MARK|3|5|et circumspiciens eos cum ira contristatus super caecitatem cordis eorum dicit homini extende manum tuam et extendit et restituta est manus illi
MARK|3|6|exeuntes autem statim Pharisaei cum Herodianis consilium faciebant adversus eum quomodo eum perderent
MARK|3|7|et Iesus cum discipulis suis secessit ad mare et multa turba a Galilaea et Iudaea secuta est eum
MARK|3|8|et ab Hierosolymis et ab Idumea et trans Iordanen et qui circa Tyrum et Sidonem multitudo magna audientes quae faciebat venerunt ad eum
MARK|3|9|et dixit discipulis suis ut navicula sibi deserviret propter turbam ne conprimerent eum
MARK|3|10|multos enim sanabat ita ut inruerent in eum ut illum tangerent quotquot habebant plagas
MARK|3|11|et spiritus inmundi cum illum videbant procidebant ei et clamabant dicentes
MARK|3|12|tu es Filius Dei et vehementer comminabatur eis ne manifestarent illum
MARK|3|13|et ascendens in montem vocavit ad se quos voluit ipse et venerunt ad eum
MARK|3|14|et fecit ut essent duodecim cum illo et ut mitteret eos praedicare
MARK|3|15|et dedit illis potestatem curandi infirmitates et eiciendi daemonia
MARK|3|16|et inposuit Simoni nomen Petrus
MARK|3|17|et Iacobum Zebedaei et Iohannem fratrem Iacobi et inposuit eis nomina Boanerges quod est Filii tonitrui
MARK|3|18|et Andream et Philippum et Bartholomeum et Mattheum et Thomam et Iacobum Alphei et Thaddeum et Simonem Cananeum
MARK|3|19|et Iudam Scarioth qui et tradidit illum
MARK|3|20|et veniunt ad domum et convenit iterum turba ita ut non possent neque panem manducare
MARK|3|21|et cum audissent sui exierunt tenere eum dicebant enim quoniam in furorem versus est
MARK|3|22|et scribae qui ab Hierosolymis descenderant dicebant quoniam Beelzebub habet et quia in principe daemonum eicit daemonia
MARK|3|23|et convocatis eis in parabolis dicebat illis quomodo potest Satanas Satanan eicere
MARK|3|24|et si regnum in se dividatur non potest stare regnum illud
MARK|3|25|et si domus super semet ipsam dispertiatur non poterit domus illa stare
MARK|3|26|et si Satanas consurrexit in semet ipsum dispertitus est et non potest stare sed finem habet
MARK|3|27|nemo potest vasa fortis ingressus in domum diripere nisi prius fortem alliget et tunc domum eius diripiet
MARK|3|28|amen dico vobis quoniam omnia dimittentur filiis hominum peccata et blasphemiae quibus blasphemaverint
MARK|3|29|qui autem blasphemaverit in Spiritum Sanctum non habet remissionem in aeternum sed reus erit aeterni delicti
MARK|3|30|quoniam dicebant spiritum inmundum habet
MARK|3|31|et veniunt mater eius et fratres et foris stantes miserunt ad eum vocantes eum
MARK|3|32|et sedebat circa eum turba et dicunt ei ecce mater tua et fratres tui foris quaerunt te
MARK|3|33|et respondens eis ait quae est mater mea et fratres mei
MARK|3|34|et circumspiciens eos qui in circuitu eius sedebant ait ecce mater mea et fratres mei
MARK|3|35|qui enim fecerit voluntatem Dei hic frater meus et soror mea et mater est
MARK|4|1|et iterum coepit docere ad mare et congregata est ad eum turba multa ita ut in navem ascendens sederet in mari et omnis turba circa mare super terram erat
MARK|4|2|et docebat eos in parabolis multa et dicebat illis in doctrina sua
MARK|4|3|audite ecce exiit seminans ad seminandum
MARK|4|4|et dum seminat aliud cecidit circa viam et venerunt volucres et comederunt illud
MARK|4|5|aliud vero cecidit super petrosa ubi non habuit terram multam et statim exortum est quoniam non habebat altitudinem terrae
MARK|4|6|et quando exortus est sol exaestuavit et eo quod non haberet radicem exaruit
MARK|4|7|et aliud cecidit in spinas et ascenderunt spinae et offocaverunt illud et fructum non dedit
MARK|4|8|et aliud cecidit in terram bonam et dabat fructum ascendentem et crescentem et adferebat unum triginta et unum sexaginta et unum centum
MARK|4|9|et dicebat qui habet aures audiendi audiat
MARK|4|10|et cum esset singularis interrogaverunt eum hii qui cum eo erant cum duodecim parabolas
MARK|4|11|et dicebat eis vobis datum est mysterium regni Dei illis autem qui foris sunt in parabolis omnia fiunt
MARK|4|12|ut videntes videant et non videant et audientes audiant et non intellegant nequando convertantur et dimittantur eis peccata
MARK|4|13|et ait illis nescitis parabolam hanc et quomodo omnes parabolas cognoscetis
MARK|4|14|qui seminat verbum seminat
MARK|4|15|hii autem sunt qui circa viam ubi seminatur verbum et cum audierint confestim venit Satanas et aufert verbum quod seminatum est in corda eorum
MARK|4|16|et hii sunt similiter qui super petrosa seminantur qui cum audierint verbum statim cum gaudio accipiunt illud
MARK|4|17|et non habent radicem in se sed temporales sunt deinde orta tribulatione et persecutione propter verbum confestim scandalizantur
MARK|4|18|et alii sunt qui in spinis seminantur hii sunt qui verbum audiunt
MARK|4|19|et aerumnae saeculi et deceptio divitiarum et circa reliqua concupiscentiae introeuntes suffocant verbum et sine fructu efficitur
MARK|4|20|et hii sunt qui super terram bonam seminati sunt qui audiunt verbum et suscipiunt et fructificant unum triginta et unum sexaginta et unum centum
MARK|4|21|et dicebat illis numquid venit lucerna ut sub modio ponatur aut sub lecto nonne ut super candelabrum ponatur
MARK|4|22|non enim est aliquid absconditum quod non manifestetur nec factum est occultum sed ut in palam veniat
MARK|4|23|si quis habet aures audiendi audiat
MARK|4|24|et dicebat illis videte quid audiatis in qua mensura mensi fueritis remetietur vobis et adicietur vobis
MARK|4|25|qui enim habet dabitur illi et qui non habet etiam quod habet auferetur ab illo
MARK|4|26|et dicebat sic est regnum Dei quemadmodum si homo iaciat sementem in terram
MARK|4|27|et dormiat et exsurgat nocte ac die et semen germinet et increscat dum nescit ille
MARK|4|28|ultro enim terra fructificat primum herbam deinde spicam deinde plenum frumentum in spica
MARK|4|29|et cum se produxerit fructus statim mittit falcem quoniam adest messis
MARK|4|30|et dicebat cui adsimilabimus regnum Dei aut cui parabolae conparabimus illud
MARK|4|31|sicut granum sinapis quod cum seminatum fuerit in terra minus est omnibus seminibus quae sunt in terra
MARK|4|32|et cum seminatum fuerit ascendit et fit maius omnibus holeribus et facit ramos magnos ita ut possint sub umbra eius aves caeli habitare
MARK|4|33|et talibus multis parabolis loquebatur eis verbum prout poterant audire
MARK|4|34|sine parabola autem non loquebatur eis seorsum autem discipulis suis disserebat omnia
MARK|4|35|et ait illis illa die cum sero esset factum transeamus contra
MARK|4|36|et dimittentes turbam adsumunt eum ita ut erat in navi et aliae naves erant cum illo
MARK|4|37|et facta est procella magna venti et fluctus mittebat in navem ita ut impleretur navis
MARK|4|38|et erat ipse in puppi supra cervical dormiens et excitant eum et dicunt ei magister non ad te pertinet quia perimus
MARK|4|39|et exsurgens comminatus est vento et dixit mari tace obmutesce et cessavit ventus et facta est tranquillitas magna
MARK|4|40|et ait illis quid timidi estis necdum habetis fidem et timuerunt magno timore et dicebant ad alterutrum quis putas est iste quia et ventus et mare oboediunt ei
MARK|5|1|et venerunt trans fretum maris in regionem Gerasenorum
MARK|5|2|et exeunti ei de navi statim occurrit ei de monumentis homo in spiritu inmundo
MARK|5|3|qui domicilium habebat in monumentis et neque catenis iam quisquam eum poterat ligare
MARK|5|4|quoniam saepe conpedibus et catenis vinctus disrupisset catenas et conpedes comminuisset et nemo poterat eum domare
MARK|5|5|et semper nocte ac die in monumentis et in montibus erat clamans et concidens se lapidibus
MARK|5|6|videns autem Iesum a longe cucurrit et adoravit eum
MARK|5|7|et clamans voce magna dicit quid mihi et tibi Iesu Fili Dei summi adiuro te per Deum ne me torqueas
MARK|5|8|dicebat enim illi exi spiritus inmunde ab homine
MARK|5|9|et interrogabat eum quod tibi nomen est et dicit ei Legio nomen mihi est quia multi sumus
MARK|5|10|et deprecabatur eum multum ne se expelleret extra regionem
MARK|5|11|erat autem ibi circa montem grex porcorum magnus pascens
MARK|5|12|et deprecabantur eum spiritus dicentes mitte nos in porcos ut in eos introeamus
MARK|5|13|et concessit eis statim Iesus et exeuntes spiritus inmundi introierunt in porcos et magno impetu grex praecipitatus est in mare ad duo milia et suffocati sunt in mare
MARK|5|14|qui autem pascebant eos fugerunt et nuntiaverunt in civitatem et in agros et egressi sunt videre quid esset facti
MARK|5|15|et veniunt ad Iesum et vident illum qui a daemonio vexabatur sedentem vestitum et sanae mentis et timuerunt
MARK|5|16|et narraverunt illis qui viderant qualiter factum esset ei qui daemonium habuerat et de porcis
MARK|5|17|et rogare eum coeperunt ut discederet de finibus eorum
MARK|5|18|cumque ascenderet navem coepit illum deprecari qui daemonio vexatus fuerat ut esset cum illo
MARK|5|19|et non admisit eum sed ait illi vade in domum tuam ad tuos et adnuntia illis quanta tibi Dominus fecerit et misertus sit tui
MARK|5|20|et abiit et coepit praedicare in Decapoli quanta sibi fecisset Iesus et omnes mirabantur
MARK|5|21|et cum transcendisset Iesus in navi rursus trans fretum convenit turba multa ad illum et erat circa mare
MARK|5|22|et venit quidam de archisynagogis nomine Iairus et videns eum procidit ad pedes eius
MARK|5|23|et deprecabatur eum multum dicens quoniam filia mea in extremis est veni inpone manus super eam ut salva sit et vivat
MARK|5|24|et abiit cum illo et sequebatur eum turba multa et conprimebant illum
MARK|5|25|et mulier quae erat in profluvio sanguinis annis duodecim
MARK|5|26|et fuerat multa perpessa a conpluribus medicis et erogaverat omnia sua nec quicquam profecerat sed magis deterius habebat
MARK|5|27|cum audisset de Iesu venit in turba retro et tetigit vestimentum eius
MARK|5|28|dicebat enim quia si vel vestimentum eius tetigero salva ero
MARK|5|29|et confestim siccatus est fons sanguinis eius et sensit corpore quod sanata esset a plaga
MARK|5|30|et statim Iesus cognoscens in semet ipso virtutem quae exierat de eo conversus ad turbam aiebat quis tetigit vestimenta mea
MARK|5|31|et dicebant ei discipuli sui vides turbam conprimentem te et dicis quis me tetigit
MARK|5|32|et circumspiciebat videre eam quae hoc fecerat
MARK|5|33|mulier autem timens et tremens sciens quod factum esset in se venit et procidit ante eum et dixit ei omnem veritatem
MARK|5|34|ille autem dixit ei filia fides tua te salvam fecit vade in pace et esto sana a plaga tua
MARK|5|35|adhuc eo loquente veniunt ab archisynagogo dicentes quia filia tua mortua est quid ultra vexas magistrum
MARK|5|36|Iesus autem verbo quod dicebatur audito ait archisynagogo noli timere tantummodo crede
MARK|5|37|et non admisit quemquam sequi se nisi Petrum et Iacobum et Iohannem fratrem Iacobi
MARK|5|38|et veniunt in domum archisynagogi et videt tumultum et flentes et heiulantes multum
MARK|5|39|et ingressus ait eis quid turbamini et ploratis puella non est mortua sed dormit
MARK|5|40|et inridebant eum ipse vero eiectis omnibus adsumit patrem et matrem puellae et qui secum erant et ingreditur ubi erat puella iacens
MARK|5|41|et tenens manum puellae ait illi talitha cumi quod est interpretatum puella tibi dico surge
MARK|5|42|et confestim surrexit puella et ambulabat erat autem annorum duodecim et obstipuerunt stupore maximo
MARK|5|43|et praecepit illis vehementer ut nemo id sciret et dixit dari illi manducare
MARK|6|1|et egressus inde abiit in patriam suam et sequebantur illum discipuli sui
MARK|6|2|et facto sabbato coepit in synagoga docere et multi audientes admirabantur in doctrina eius dicentes unde huic haec omnia et quae est sapientia quae data est illi et virtutes tales quae per manus eius efficiuntur
MARK|6|3|nonne iste est faber filius Mariae frater Iacobi et Ioseph et Iudae et Simonis nonne et sorores eius hic nobiscum sunt et scandalizabantur in illo
MARK|6|4|et dicebat eis Iesus quia non est propheta sine honore nisi in patria sua et in cognatione sua et in domo sua
MARK|6|5|et non poterat ibi virtutem ullam facere nisi paucos infirmos inpositis manibus curavit
MARK|6|6|et mirabatur propter incredulitatem eorum
MARK|6|7|et circumibat castella in circuitu docens et convocavit duodecim et coepit eos mittere binos et dabat illis potestatem spirituum inmundorum
MARK|6|8|et praecepit eis ne quid tollerent in via nisi virgam tantum non peram non panem neque in zona aes
MARK|6|9|sed calciatos sandaliis et ne induerentur duabus tunicis
MARK|6|10|et dicebat eis quocumque introieritis in domum illic manete donec exeatis inde
MARK|6|11|et quicumque non receperint vos nec audierint vos exeuntes inde excutite pulverem de pedibus vestris in testimonium illis
MARK|6|12|et exeuntes praedicabant ut paenitentiam agerent
MARK|6|13|et daemonia multa eiciebant et unguebant oleo multos aegrotos et sanabant
MARK|6|14|et audivit Herodes rex manifestum enim factum est nomen eius et dicebat quia Iohannes Baptista resurrexit a mortuis et propterea inoperantur virtutes in illo
MARK|6|15|alii autem dicebant quia Helias est alii vero dicebant propheta est quasi unus ex prophetis
MARK|6|16|quo audito Herodes ait quem ego decollavi Iohannem hic a mortuis resurrexit
MARK|6|17|ipse enim Herodes misit ac tenuit Iohannem et vinxit eum in carcere propter Herodiadem uxorem Philippi fratris sui quia duxerat eam
MARK|6|18|dicebat enim Iohannes Herodi non licet tibi habere uxorem fratris tui
MARK|6|19|Herodias autem insidiabatur illi et volebat occidere eum nec poterat
MARK|6|20|Herodes enim metuebat Iohannem sciens eum virum iustum et sanctum et custodiebat eum et audito eo multa faciebat et libenter eum audiebat
MARK|6|21|et cum dies oportunus accidisset Herodes natalis sui cenam fecit principibus et tribunis et primis Galilaeae
MARK|6|22|cumque introisset filia ipsius Herodiadis et saltasset et placuisset Herodi simulque recumbentibus rex ait puellae pete a me quod vis et dabo tibi
MARK|6|23|et iuravit illi quia quicquid petieris dabo tibi licet dimidium regni mei
MARK|6|24|quae cum exisset dixit matri suae quid petam et illa dixit caput Iohannis Baptistae
MARK|6|25|cumque introisset statim cum festinatione ad regem petivit dicens volo ut protinus des mihi in disco caput Iohannis Baptistae
MARK|6|26|et contristatus rex propter iusiurandum et propter simul recumbentes noluit eam contristare
MARK|6|27|sed misso speculatore praecepit adferri caput eius in disco et decollavit eum in carcere
MARK|6|28|et adtulit caput eius in disco et dedit illud puellae et puella dedit matri suae
MARK|6|29|quo audito discipuli eius venerunt et tulerunt corpus eius et posuerunt illud in monumento
MARK|6|30|et convenientes apostoli ad Iesum renuntiaverunt illi omnia quae egerant et docuerant
MARK|6|31|et ait illis venite seorsum in desertum locum et requiescite pusillum erant enim qui veniebant et rediebant multi et nec manducandi spatium habebant
MARK|6|32|et ascendentes in navi abierunt in desertum locum seorsum
MARK|6|33|et viderunt eos abeuntes et cognoverunt multi et pedestre et de omnibus civitatibus concurrerunt illuc et praevenerunt eos
MARK|6|34|et exiens vidit multam turbam Iesus et misertus est super eos quia erant sicut oves non habentes pastorem et coepit docere illos multa
MARK|6|35|et cum iam hora multa fieret accesserunt discipuli eius dicentes desertus est locus hic et iam hora praeterivit
MARK|6|36|dimitte illos ut euntes in proximas villas et vicos emant sibi cibos quos manducent
MARK|6|37|et respondens ait illis date illis manducare et dixerunt ei euntes emamus denariis ducentis panes et dabimus eis manducare
MARK|6|38|et dicit eis quot panes habetis ite et videte et cum cognovissent dicunt quinque et duos pisces
MARK|6|39|et praecepit illis ut accumbere facerent omnes secundum contubernia super viride faenum
MARK|6|40|et discubuerunt in partes per centenos et per quinquagenos
MARK|6|41|et acceptis quinque panibus et duobus piscibus intuens in caelum benedixit et fregit panes et dedit discipulis suis ut ponerent ante eos et duos pisces divisit omnibus
MARK|6|42|et manducaverunt omnes et saturati sunt
MARK|6|43|et sustulerunt reliquias fragmentorum duodecim cofinos plenos et de piscibus
MARK|6|44|erant autem qui manducaverunt quinque milia virorum
MARK|6|45|et statim coegit discipulos suos ascendere navem ut praecederent eum trans fretum ad Bethsaidam dum ipse dimitteret populum
MARK|6|46|et cum dimisisset eos abiit in montem orare
MARK|6|47|et cum sero esset erat navis in medio mari et ipse solus in terra
MARK|6|48|et videns eos laborantes in remigando erat enim ventus contrarius eis et circa quartam vigiliam noctis venit ad eos ambulans super mare et volebat praeterire eos
MARK|6|49|at illi ut viderunt eum ambulantem super mare putaverunt fantasma esse et exclamaverunt
MARK|6|50|omnes enim eum viderunt et conturbati sunt et statim locutus est cum eis et dixit illis confidite ego sum nolite timere
MARK|6|51|et ascendit ad illos in navem et cessavit ventus et plus magis intra se stupebant
MARK|6|52|non enim intellexerant de panibus erat enim cor illorum obcaecatum
MARK|6|53|et cum transfretassent pervenerunt in terram Gennesareth et adplicuerunt
MARK|6|54|cumque egressi essent de navi continuo cognoverunt eum
MARK|6|55|et percurrentes universam regionem illam coeperunt in grabattis eos qui se male habebant circumferre ubi audiebant eum esse
MARK|6|56|et quocumque introibat in vicos vel in villas aut civitates in plateis ponebant infirmos et deprecabantur eum ut vel fimbriam vestimenti eius tangerent et quotquot tangebant eum salvi fiebant
MARK|7|1|et conveniunt ad eum Pharisaei et quidam de scribis venientes ab Hierosolymis
MARK|7|2|et cum vidissent quosdam ex discipulis eius communibus manibus id est non lotis manducare panes vituperaverunt
MARK|7|3|Pharisaei enim et omnes Iudaei nisi crebro lavent manus non manducant tenentes traditionem seniorum
MARK|7|4|et a foro nisi baptizentur non comedunt et alia multa sunt quae tradita sunt illis servare baptismata calicum et urceorum et aeramentorum et lectorum
MARK|7|5|et interrogant eum Pharisaei et scribae quare discipuli tui non ambulant iuxta traditionem seniorum sed communibus manibus manducant panem
MARK|7|6|at ille respondens dixit eis bene prophetavit Esaias de vobis hypocritis sicut scriptum est populus hic labiis me honorat cor autem eorum longe est a me
MARK|7|7|in vanum autem me colunt docentes doctrinas praecepta hominum
MARK|7|8|relinquentes enim mandatum Dei tenetis traditionem hominum baptismata urceorum et calicum et alia similia his facitis multa
MARK|7|9|et dicebat illis bene irritum facitis praeceptum Dei ut traditionem vestram servetis
MARK|7|10|Moses enim dixit honora patrem tuum et matrem tuam et qui maledixerit patri aut matri morte moriatur
MARK|7|11|vos autem dicitis si dixerit homo patri aut matri corban quod est donum quodcumque ex me tibi profuerit
MARK|7|12|et ultra non dimittitis eum quicquam facere patri suo aut matri
MARK|7|13|rescindentes verbum Dei per traditionem vestram quam tradidistis et similia huiusmodi multa facitis
MARK|7|14|et advocans iterum turbam dicebat illis audite me omnes et intellegite
MARK|7|15|nihil est extra hominem introiens in eum quod possit eum coinquinare sed quae de homine procedunt illa sunt quae communicant hominem
MARK|7|16|si quis habet aures audiendi audiat
MARK|7|17|et cum introisset in domum a turba interrogabant eum discipuli eius parabolam
MARK|7|18|et ait illis sic et vos inprudentes estis non intellegitis quia omne extrinsecus introiens in hominem non potest eum communicare
MARK|7|19|quia non introit in cor eius sed in ventrem et in secessum exit purgans omnes escas
MARK|7|20|dicebat autem quoniam quae de homine exeunt illa communicant hominem
MARK|7|21|ab intus enim de corde hominum cogitationes malae procedunt adulteria fornicationes homicidia
MARK|7|22|furta avaritiae nequitiae dolus inpudicitia oculus malus blasphemia superbia stultitia
MARK|7|23|omnia haec mala ab intus procedunt et communicant hominem
MARK|7|24|et inde surgens abiit in fines Tyri et Sidonis et ingressus domum neminem voluit scire et non potuit latere
MARK|7|25|mulier enim statim ut audivit de eo cuius habebat filia spiritum inmundum intravit et procidit ad pedes eius
MARK|7|26|erat autem mulier gentilis Syrophoenissa genere et rogabat eum ut daemonium eiceret de filia eius
MARK|7|27|qui dixit illi sine prius saturari filios non est enim bonum sumere panem filiorum et mittere canibus
MARK|7|28|at illa respondit et dicit ei utique Domine nam et catelli sub mensa comedunt de micis puerorum
MARK|7|29|et ait illi propter hunc sermonem vade exiit daemonium de filia tua
MARK|7|30|et cum abisset domum suam invenit puellam iacentem supra lectum et daemonium exisse
MARK|7|31|et iterum exiens de finibus Tyri venit per Sidonem ad mare Galilaeae inter medios fines Decapoleos
MARK|7|32|et adducunt ei surdum et mutum et deprecantur eum ut inponat illi manum
MARK|7|33|et adprehendens eum de turba seorsum misit digitos suos in auriculas et expuens tetigit linguam eius
MARK|7|34|et suspiciens in caelum ingemuit et ait illi eppheta quod est adaperire
MARK|7|35|et statim apertae sunt aures eius et solutum est vinculum linguae eius et loquebatur recte
MARK|7|36|et praecepit illis ne cui dicerent quanto autem eis praecipiebat tanto magis plus praedicabant
MARK|7|37|et eo amplius admirabantur dicentes bene omnia fecit et surdos facit audire et mutos loqui
MARK|8|1|in illis diebus iterum cum turba multa esset nec haberent quod manducarent convocatis discipulis ait illis
MARK|8|2|misereor super turba quia ecce iam triduo sustinent me nec habent quod manducent
MARK|8|3|et si dimisero eos ieiunos in domum suam deficient in via quidam enim ex eis de longe venerunt
MARK|8|4|et responderunt ei discipuli sui unde istos poterit quis hic saturare panibus in solitudine
MARK|8|5|et interrogavit eos quot panes habetis qui dixerunt septem
MARK|8|6|et praecepit turbae discumbere supra terram et accipiens septem panes gratias agens fregit et dabat discipulis suis ut adponerent et adposuerunt turbae
MARK|8|7|et habebant pisciculos paucos et ipsos benedixit et iussit adponi
MARK|8|8|et manducaverunt et saturati sunt et sustulerunt quod superaverat de fragmentis septem sportas
MARK|8|9|erant autem qui manducaverunt quasi quattuor milia et dimisit eos
MARK|8|10|et statim ascendens navem cum discipulis suis venit in partes Dalmanutha
MARK|8|11|et exierunt Pharisaei et coeperunt conquirere cum eo quaerentes ab illo signum de caelo temptantes eum
MARK|8|12|et ingemescens spiritu ait quid generatio ista quaerit signum amen dico vobis si dabitur generationi isti signum
MARK|8|13|et dimittens eos ascendens iterum abiit trans fretum
MARK|8|14|et obliti sunt sumere panes et nisi unum panem non habebant secum in navi
MARK|8|15|et praecipiebat eis dicens videte cavete a fermento Pharisaeorum et fermento Herodis
MARK|8|16|et cogitabant ad alterutrum dicentes quia panes non habemus
MARK|8|17|quo cognito Iesus ait illis quid cogitatis quia panes non habetis nondum cognoscitis nec intellegitis adhuc caecatum habetis cor vestrum
MARK|8|18|oculos habentes non videtis et aures habentes non auditis nec recordamini
MARK|8|19|quando quinque panes fregi in quinque milia et quot cofinos fragmentorum plenos sustulistis dicunt ei duodecim
MARK|8|20|quando et septem panes in quattuor milia quot sportas fragmentorum tulistis et dicunt ei septem
MARK|8|21|et dicebat eis quomodo nondum intellegitis
MARK|8|22|et veniunt Bethsaida et adducunt ei caecum et rogabant eum ut illum tangeret
MARK|8|23|et adprehendens manum caeci eduxit eum extra vicum et expuens in oculos eius inpositis manibus suis interrogavit eum si aliquid videret
MARK|8|24|et aspiciens ait video homines velut arbores ambulantes
MARK|8|25|deinde iterum inposuit manus super oculos eius et coepit videre et restitutus est ita ut videret clare omnia
MARK|8|26|et misit illum in domum suam dicens vade in domum tuam et si in vicum introieris nemini dixeris
MARK|8|27|et egressus est Iesus et discipuli eius in castella Caesareae Philippi et in via interrogabat discipulos suos dicens eis quem me dicunt esse homines
MARK|8|28|qui responderunt illi dicentes Iohannem Baptistam alii Heliam alii vero quasi unum de prophetis
MARK|8|29|tunc dicit illis vos vero quem me dicitis esse respondens Petrus ait ei tu es Christus
MARK|8|30|et comminatus est eis ne cui dicerent de illo
MARK|8|31|et coepit docere illos quoniam oportet Filium hominis multa pati et reprobari a senioribus et a summis sacerdotibus et scribis et occidi et post tres dies resurgere
MARK|8|32|et palam verbum loquebatur et adprehendens eum Petrus coepit increpare eum
MARK|8|33|qui conversus et videns discipulos suos comminatus est Petro dicens vade retro me Satana quoniam non sapis quae Dei sunt sed quae sunt hominum
MARK|8|34|et convocata turba cum discipulis suis dixit eis si quis vult post me sequi deneget se ipsum et tollat crucem suam et sequatur me
MARK|8|35|qui enim voluerit animam suam salvam facere perdet eam qui autem perdiderit animam suam propter me et evangelium salvam eam faciet
MARK|8|36|quid enim proderit homini si lucretur mundum totum et detrimentum faciat animae suae
MARK|8|37|aut quid dabit homo commutationem pro anima sua
MARK|8|38|qui enim me confusus fuerit et mea verba in generatione ista adultera et peccatrice et Filius hominis confundetur eum cum venerit in gloria Patris sui cum angelis sanctis
MARK|8|39|et dicebat illis amen dico vobis quia sunt quidam de hic stantibus qui non gustabunt mortem donec videant regnum Dei veniens in virtute
MARK|9|1|et post dies sex adsumit Iesus Petrum et Iacobum et Iohannem et ducit illos in montem excelsum seorsum solos et transfiguratus est coram ipsis
MARK|9|2|et vestimenta eius facta sunt splendentia candida nimis velut nix qualia fullo super terram non potest candida facere
MARK|9|3|et apparuit illis Helias cum Mose et erant loquentes cum Iesu
MARK|9|4|et respondens Petrus ait Iesu rabbi bonum est hic nos esse et faciamus tria tabernacula tibi unum et Mosi unum et Heliae unum
MARK|9|5|non enim sciebat quid diceret erant enim timore exterriti
MARK|9|6|et facta est nubes obumbrans eos et venit vox de nube dicens hic est Filius meus carissimus audite illum
MARK|9|7|et statim circumspicientes neminem amplius viderunt nisi Iesum tantum secum
MARK|9|8|et descendentibus illis de monte praecepit illis ne cui quae vidissent narrarent nisi cum Filius hominis a mortuis resurrexerit
MARK|9|9|et verbum continuerunt apud se conquirentes quid esset cum a mortuis resurrexerit
MARK|9|10|et interrogabant eum dicentes quid ergo dicunt Pharisaei et scribae quia Heliam oporteat venire primum
MARK|9|11|qui respondens ait illis Helias cum venerit primo restituet omnia et quomodo scriptum est in Filium hominis ut multa patiatur et contemnatur
MARK|9|12|sed dico vobis quia et Helias venit et fecerunt illi quaecumque voluerunt sicut scriptum est de eo
MARK|9|13|et veniens ad discipulos suos vidit turbam magnam circa eos et scribas conquirentes cum illis
MARK|9|14|et confestim omnis populus videns eum stupefactus est et adcurrentes salutabant eum
MARK|9|15|et interrogavit eos quid inter vos conquiritis
MARK|9|16|et respondens unus de turba dixit magister adtuli filium meum ad te habentem spiritum mutum
MARK|9|17|qui ubicumque eum adprehenderit adlidit eum et spumat et stridet dentibus et arescit et dixi discipulis tuis ut eicerent illum et non potuerunt
MARK|9|18|qui respondens eis dicit o generatio incredula quamdiu apud vos ero quamdiu vos patiar adferte illum ad me
MARK|9|19|et adtulerunt eum et cum vidisset illum statim spiritus conturbavit eum et elisus in terram volutabatur spumans
MARK|9|20|et interrogavit patrem eius quantum temporis est ex quo hoc ei accidit at ille ait ab infantia
MARK|9|21|et frequenter eum et in ignem et in aquas misit ut eum perderet sed si quid potes adiuva nos misertus nostri
MARK|9|22|Iesus autem ait illi si potes credere omnia possibilia credenti
MARK|9|23|et continuo exclamans pater pueri cum lacrimis aiebat credo adiuva incredulitatem meam
MARK|9|24|et cum videret Iesus concurrentem turbam comminatus est spiritui inmundo dicens illi surde et mute spiritus ego tibi praecipio exi ab eo et amplius ne introeas in eum
MARK|9|25|et clamans et multum discerpens eum exiit ab eo et factus est sicut mortuus ita ut multi dicerent quia mortuus est
MARK|9|26|Iesus autem tenens manum eius elevavit illum et surrexit
MARK|9|27|et cum introisset in domum discipuli eius secreto interrogabant eum quare nos non potuimus eicere eum
MARK|9|28|et dixit illis hoc genus in nullo potest exire nisi in oratione et ieiunio
MARK|9|29|et inde profecti praetergrediebantur Galilaeam nec volebat quemquam scire
MARK|9|30|docebat autem discipulos suos et dicebat illis quoniam Filius hominis tradetur in manus hominum et occident eum et occisus tertia die resurget
MARK|9|31|at illi ignorabant verbum et timebant eum interrogare
MARK|9|32|et venerunt Capharnaum qui cum domi esset interrogabat eos quid in via tractabatis
MARK|9|33|at illi tacebant siquidem inter se in via disputaverant quis esset illorum maior
MARK|9|34|et residens vocavit duodecim et ait illis si quis vult primus esse erit omnium novissimus et omnium minister
MARK|9|35|et accipiens puerum statuit eum in medio eorum quem cum conplexus esset ait illis
MARK|9|36|quisquis unum ex huiusmodi pueris receperit in nomine meo me recipit et quicumque me susceperit non me suscipit sed eum qui me misit
MARK|9|37|respondit illi Iohannes dicens magister vidimus quendam in nomine tuo eicientem daemonia qui non sequitur nos et prohibuimus eum
MARK|9|38|Iesus autem ait nolite prohibere eum nemo est enim qui faciat virtutem in nomine meo et possit cito male loqui de me
MARK|9|39|qui enim non est adversum vos pro vobis est
MARK|9|40|quisquis enim potum dederit vobis calicem aquae in nomine meo quia Christi estis amen dico vobis non perdet mercedem suam
MARK|9|41|et quisquis scandalizaverit unum ex his pusillis credentibus in me bonum est ei magis si circumdaretur mola asinaria collo eius et in mare mitteretur
MARK|9|42|et si scandalizaverit te manus tua abscide illam bonum est tibi debilem introire in vitam quam duas manus habentem ire in gehennam in ignem inextinguibilem
MARK|9|43|ubi vermis eorum non moritur et ignis non extinguitur
MARK|9|44|et si pes tuus te scandalizat amputa illum bonum est tibi claudum introire in vitam aeternam quam duos pedes habentem mitti in gehennam ignis inextinguibilis
MARK|9|45|ubi vermis eorum non moritur et ignis non extinguitur
MARK|9|46|quod si oculus tuus scandalizat te eice eum bonum est tibi luscum introire in regnum Dei quam duos oculos habentem mitti in gehennam ignis
MARK|9|47|ubi vermis eorum non moritur et ignis non extinguitur
MARK|9|48|omnis enim igne sallietur et omnis victima sallietur
MARK|9|49|bonum est sal quod si sal insulsum fuerit in quo illud condietis habete in vobis sal et pacem habete inter vos
MARK|9|50|
MARK|10|1|et inde exsurgens venit in fines Iudaeae ultra Iordanen et conveniunt iterum turbae ad eum et sicut consueverat iterum docebat illos
MARK|10|2|et accedentes Pharisaei interrogabant eum si licet viro uxorem dimittere temptantes eum
MARK|10|3|at ille respondens dixit eis quid vobis praecepit Moses
MARK|10|4|qui dixerunt Moses permisit libellum repudii scribere et dimittere
MARK|10|5|quibus respondens Iesus ait ad duritiam cordis vestri scripsit vobis praeceptum istud
MARK|10|6|ab initio autem creaturae masculum et feminam fecit eos Deus
MARK|10|7|propter hoc relinquet homo patrem suum et matrem et adherebit ad uxorem suam
MARK|10|8|et erunt duo in carne una itaque iam non sunt duo sed una caro
MARK|10|9|quod ergo Deus iunxit homo non separet
MARK|10|10|et in domo iterum discipuli eius de eodem interrogaverunt eum
MARK|10|11|et dicit illis quicumque dimiserit uxorem suam et aliam duxerit adulterium committit super eam
MARK|10|12|et si uxor dimiserit virum suum et alii nupserit moechatur
MARK|10|13|et offerebant illi parvulos ut tangeret illos discipuli autem comminabantur offerentibus
MARK|10|14|quos cum videret Iesus indigne tulit et ait illis sinite parvulos venire ad me et ne prohibueritis eos talium est enim regnum Dei
MARK|10|15|amen dico vobis quisque non receperit regnum Dei velut parvulus non intrabit in illud
MARK|10|16|et conplexans eos et inponens manus super illos benedicebat eos
MARK|10|17|et cum egressus esset in viam procurrens quidam genu flexo ante eum rogabat eum magister bone quid faciam ut vitam aeternam percipiam
MARK|10|18|Iesus autem dixit ei quid me dicis bonum nemo bonus nisi unus Deus
MARK|10|19|praecepta nosti ne adulteres ne occidas ne fureris ne falsum testimonium dixeris ne fraudem feceris honora patrem tuum et matrem
MARK|10|20|et ille respondens ait illi magister omnia haec conservavi a iuventute mea
MARK|10|21|Iesus autem intuitus eum dilexit eum et dixit illi unum tibi deest vade quaecumque habes vende et da pauperibus et habebis thesaurum in caelo et veni sequere me
MARK|10|22|qui contristatus in verbo abiit maerens erat enim habens possessiones multas
MARK|10|23|et circumspiciens Iesus ait discipulis suis quam difficile qui pecunias habent in regnum Dei introibunt
MARK|10|24|discipuli autem obstupescebant in verbis eius at Iesus rursus respondens ait illis filioli quam difficile est confidentes in pecuniis regnum Dei introire
MARK|10|25|facilius est camelum per foramen acus transire quam divitem intrare in regnum Dei
MARK|10|26|qui magis admirabantur dicentes ad semet ipsos et quis potest salvus fieri
MARK|10|27|et intuens illos Iesus ait apud homines inpossibile est sed non apud Deum omnia enim possibilia sunt apud Deum
MARK|10|28|coepit Petrus ei dicere ecce nos dimisimus omnia et secuti sumus te
MARK|10|29|respondens Iesus ait amen dico vobis nemo est qui reliquerit domum aut fratres aut sorores aut matrem aut patrem aut filios aut agros propter me et propter evangelium
MARK|10|30|qui non accipiat centies tantum nunc in tempore hoc domos et fratres et sorores et matres et filios et agros cum persecutionibus et in saeculo futuro vitam aeternam
MARK|10|31|multi autem erunt primi novissimi et novissimi primi
MARK|10|32|erant autem in via ascendentes in Hierosolyma et praecedebat illos Iesus et stupebant et sequentes timebant et adsumens iterum duodecim coepit illis dicere quae essent ei ventura
MARK|10|33|quia ecce ascendimus in Hierosolyma et Filius hominis tradetur principibus sacerdotum et scribis et senioribus et damnabunt eum morti et tradent eum gentibus
MARK|10|34|et inludent ei et conspuent eum et flagellabunt eum et interficient eum et tertia die resurget
MARK|10|35|et accedunt ad illum Iacobus et Iohannes filii Zebedaei dicentes magister volumus ut quodcumque petierimus facias nobis
MARK|10|36|at ille dixit eis quid vultis ut faciam vobis
MARK|10|37|et dixerunt da nobis ut unus ad dexteram tuam et alius ad sinistram tuam sedeamus in gloria tua
MARK|10|38|Iesus autem ait eis nescitis quid petatis potestis bibere calicem quem ego bibo aut baptismum quo ego baptizor baptizari
MARK|10|39|at illi dixerunt ei possumus Iesus autem ait eis calicem quidem quem ego bibo bibetis et baptismum quo ego baptizor baptizabimini
MARK|10|40|sedere autem ad dexteram meam vel ad sinistram non est meum dare sed quibus paratum est
MARK|10|41|et audientes decem coeperunt indignari de Iacobo et Iohanne
MARK|10|42|Iesus autem vocans eos ait illis scitis quia hii qui videntur principari gentibus dominantur eis et principes eorum potestatem habent ipsorum
MARK|10|43|non ita est autem in vobis sed quicumque voluerit fieri maior erit vester minister
MARK|10|44|et quicumque voluerit in vobis primus esse erit omnium servus
MARK|10|45|nam et Filius hominis non venit ut ministraretur ei sed ut ministraret et daret animam suam redemptionem pro multis
MARK|10|46|et veniunt Hierichum et proficiscente eo de Hiericho et discipulis eius et plurima multitudine filius Timei Bartimeus caecus sedebat iuxta viam mendicans
MARK|10|47|qui cum audisset quia Iesus Nazarenus est coepit clamare et dicere Fili David Iesu miserere mei
MARK|10|48|et comminabantur illi multi ut taceret at ille multo magis clamabat Fili David miserere mei
MARK|10|49|et stans Iesus praecepit illum vocari et vocant caecum dicentes ei animaequior esto surge vocat te
MARK|10|50|qui proiecto vestimento suo exiliens venit ad eum
MARK|10|51|et respondens illi Iesus dixit quid vis tibi faciam caecus autem dixit ei rabboni ut videam
MARK|10|52|Iesus autem ait illi vade fides tua te salvum fecit et confestim vidit et sequebatur eum in via
MARK|11|1|et cum adpropinquarent Hierosolymae et Bethaniae ad montem Olivarum mittit duos ex discipulis suis
MARK|11|2|et ait illis ite in castellum quod est contra vos et statim introeuntes illuc invenietis pullum ligatum super quem nemo adhuc hominum sedit solvite illum et adducite
MARK|11|3|et si quis vobis dixerit quid facitis dicite quia Domino necessarius est et continuo illum dimittet huc
MARK|11|4|et abeuntes invenerunt pullum ligatum ante ianuam foris in bivio et solvunt eum
MARK|11|5|et quidam de illic stantibus dicebant illis quid facitis solventes pullum
MARK|11|6|qui dixerunt eis sicut praeceperat illis Iesus et dimiserunt eis
MARK|11|7|et duxerunt pullum ad Iesum et inponunt illi vestimenta sua et sedit super eo
MARK|11|8|multi autem vestimenta sua straverunt in via alii autem frondes caedebant de arboribus et sternebant in via
MARK|11|9|et qui praeibant et qui sequebantur clamabant dicentes osanna benedictus qui venit in nomine Domini
MARK|11|10|benedictum quod venit regnum patris nostri David osanna in excelsis
MARK|11|11|et introivit Hierosolyma in templum et circumspectis omnibus cum iam vespera esset hora exivit in Bethania cum duodecim
MARK|11|12|et alia die cum exirent a Bethania esuriit
MARK|11|13|cumque vidisset a longe ficum habentem folia venit si quid forte inveniret in ea et cum venisset ad eam nihil invenit praeter folia non enim erat tempus ficorum
MARK|11|14|et respondens dixit ei iam non amplius in aeternum quisquam fructum ex te manducet et audiebant discipuli eius
MARK|11|15|et veniunt Hierosolymam et cum introisset templum coepit eicere vendentes et ementes in templo et mensas nummulariorum et cathedras vendentium columbas evertit
MARK|11|16|et non sinebat ut quisquam vas transferret per templum
MARK|11|17|et docebat dicens eis non scriptum est quia domus mea domus orationis vocabitur omnibus gentibus vos autem fecistis eam speluncam latronum
MARK|11|18|quo audito principes sacerdotum et scribae quaerebant quomodo eum perderent timebant enim eum quoniam universa turba admirabatur super doctrina eius
MARK|11|19|et cum vespera facta esset egrediebatur de civitate
MARK|11|20|et cum mane transirent viderunt ficum aridam factam a radicibus
MARK|11|21|et recordatus Petrus dicit ei rabbi ecce ficus cui maledixisti aruit
MARK|11|22|et respondens Iesus ait illis habete fidem Dei
MARK|11|23|amen dico vobis quicumque dixerit huic monti tollere et mittere in mare et non haesitaverit in corde suo sed crediderit quia quodcumque dixerit fiat fiet ei
MARK|11|24|propterea dico vobis omnia quaecumque orantes petitis credite quia accipietis et veniet vobis
MARK|11|25|et cum stabitis ad orandum dimittite si quid habetis adversus aliquem ut et Pater vester qui in caelis est dimittat vobis peccata vestra
MARK|11|26|quod si vos non dimiseritis nec Pater vester qui in caelis est dimittet vobis peccata vestra
MARK|11|27|et veniunt rursus Hierosolymam et cum ambularet in templo accedunt ad eum summi sacerdotes et scribae et seniores
MARK|11|28|et dicunt illi in qua potestate haec facis et quis tibi dedit hanc potestatem ut ista facias
MARK|11|29|Iesus autem respondens ait illis interrogabo vos et ego unum verbum et respondete mihi et dicam vobis in qua potestate haec faciam
MARK|11|30|baptismum Iohannis de caelo erat an ex hominibus respondete mihi
MARK|11|31|at illi cogitabant secum dicentes si dixerimus de caelo dicet quare ergo non credidistis ei
MARK|11|32|sed dicemus ex hominibus timebant populum omnes enim habebant Iohannem quia vere propheta esset
MARK|11|33|et respondentes dicunt Iesu nescimus respondens Iesus ait illis neque ego dico vobis in qua potestate haec faciam
MARK|12|1|et coepit illis in parabolis loqui vineam pastinavit homo et circumdedit sepem et fodit lacum et aedificavit turrem et locavit eam agricolis et peregre profectus est
MARK|12|2|et misit ad agricolas in tempore servum ut ab agricolis acciperet de fructu vineae
MARK|12|3|qui adprehensum eum ceciderunt et dimiserunt vacuum
MARK|12|4|et iterum misit ad illos alium servum et illum capite vulneraverunt et contumeliis adfecerunt
MARK|12|5|et rursum alium misit et illum occiderunt et plures alios quosdam caedentes alios vero occidentes
MARK|12|6|adhuc ergo unum habens filium carissimum et illum misit ad eos novissimum dicens quia reverebuntur filium meum
MARK|12|7|coloni autem dixerunt ad invicem hic est heres venite occidamus eum et nostra erit hereditas
MARK|12|8|et adprehendentes eum occiderunt et eiecerunt extra vineam
MARK|12|9|quid ergo faciet dominus vineae veniet et perdet colonos et dabit vineam aliis
MARK|12|10|nec scripturam hanc legistis lapidem quem reprobaverunt aedificantes hic factus est in caput anguli
MARK|12|11|a Domino factum est istud et est mirabile in oculis nostris
MARK|12|12|et quaerebant eum tenere et timuerunt turbam cognoverunt enim quoniam ad eos parabolam hanc dixerit et relicto eo abierunt
MARK|12|13|et mittunt ad eum quosdam ex Pharisaeis et Herodianis ut eum caperent in verbo
MARK|12|14|qui venientes dicunt ei magister scimus quoniam verax es et non curas quemquam nec enim vides in faciem hominis sed in veritate viam Dei doces licet dari tributum Caesari an non dabimus
MARK|12|15|qui sciens versutiam eorum ait illis quid me temptatis adferte mihi denarium ut videam
MARK|12|16|at illi adtulerunt et ait illis cuius est imago haec et inscriptio dicunt illi Caesaris
MARK|12|17|respondens autem Iesus dixit illis reddite igitur quae sunt Caesaris Caesari et quae sunt Dei Deo et mirabantur super eo
MARK|12|18|et venerunt ad eum Sadducaei qui dicunt resurrectionem non esse et interrogabant eum dicentes
MARK|12|19|magister Moses nobis scripsit ut si cuius frater mortuus fuerit et dimiserit uxorem et filios non reliquerit accipiat frater eius uxorem ipsius et resuscitet semen fratri suo
MARK|12|20|septem ergo fratres erant et primus accepit uxorem et mortuus est non relicto semine
MARK|12|21|et secundus accepit eam et mortuus est et nec iste reliquit semen et tertius similiter
MARK|12|22|et acceperunt eam similiter septem et non reliquerunt semen novissima omnium defuncta est et mulier
MARK|12|23|in resurrectione ergo cum resurrexerint cuius de his erit uxor septem enim habuerunt eam uxorem
MARK|12|24|et respondens Iesus ait illis non ideo erratis non scientes scripturas neque virtutem Dei
MARK|12|25|cum enim a mortuis resurrexerint neque nubent neque nubentur sed sunt sicut angeli in caelis
MARK|12|26|de mortuis autem quod resurgant non legistis in libro Mosi super rubum quomodo dixerit illi Deus inquiens ego sum Deus Abraham et Deus Isaac et Deus Iacob
MARK|12|27|non est Deus mortuorum sed vivorum vos ergo multum erratis
MARK|12|28|et accessit unus de scribis qui audierat illos conquirentes et videns quoniam bene illis responderit interrogavit eum quod esset primum omnium mandatum
MARK|12|29|Iesus autem respondit ei quia primum omnium mandatum est audi Israhel Dominus Deus noster Deus unus est
MARK|12|30|et diliges Dominum Deum tuum ex toto corde tuo et ex tota anima tua et ex tota mente tua et ex tota virtute tua hoc est primum mandatum
MARK|12|31|secundum autem simile illi diliges proximum tuum tamquam te ipsum maius horum aliud mandatum non est
MARK|12|32|et ait illi scriba bene magister in veritate dixisti quia unus est et non est alius praeter eum
MARK|12|33|et ut diligatur ex toto corde et ex toto intellectu et ex tota anima et ex tota fortitudine et diligere proximum tamquam se ipsum maius est omnibus holocaustomatibus et sacrificiis
MARK|12|34|Iesus autem videns quod sapienter respondisset dixit illi non es longe a regno Dei et nemo iam audebat eum interrogare
MARK|12|35|et respondens Iesus dicebat docens in templo quomodo dicunt scribae Christum Filium esse David
MARK|12|36|ipse enim David dicit in Spiritu Sancto dixit Dominus Domino meo sede a dextris meis donec ponam inimicos tuos scabillum pedum tuorum
MARK|12|37|ipse ergo David dicit eum Dominum et unde est filius eius et multa turba eum libenter audivit
MARK|12|38|et dicebat eis in doctrina sua cavete a scribis qui volunt in stolis ambulare et salutari in foro
MARK|12|39|et in primis cathedris sedere in synagogis et primos discubitus in cenis
MARK|12|40|qui devorant domos viduarum sub obtentu prolixae orationis hii accipient prolixius iudicium
MARK|12|41|et sedens Iesus contra gazofilacium aspiciebat quomodo turba iactaret aes in gazofilacium et multi divites iactabant multa
MARK|12|42|cum venisset autem una vidua pauper misit duo minuta quod est quadrans
MARK|12|43|et convocans discipulos suos ait illis amen dico vobis quoniam vidua haec pauper plus omnibus misit qui miserunt in gazofilacium
MARK|12|44|omnes enim ex eo quod abundabat illis miserunt haec vero de penuria sua omnia quae habuit misit totum victum suum
MARK|13|1|et cum egrederetur de templo ait illi unus ex discipulis suis magister aspice quales lapides et quales structurae
MARK|13|2|et respondens Iesus ait illi vides has omnes magnas aedificationes non relinquetur lapis super lapidem qui non destruatur
MARK|13|3|et cum sederet in montem Olivarum contra templum interrogabant eum separatim Petrus et Iacobus et Iohannes et Andreas
MARK|13|4|dic nobis quando ista fient et quod signum erit quando haec omnia incipient consummari
MARK|13|5|et respondens Iesus coepit dicere illis videte ne quis vos seducat
MARK|13|6|multi enim venient in nomine meo dicentes quia ego sum et multos seducent
MARK|13|7|cum audieritis autem bella et opiniones bellorum ne timueritis oportet enim fieri sed nondum finis
MARK|13|8|exsurget autem gens super gentem et regnum super regnum et erunt terraemotus per loca et fames initium dolorum haec
MARK|13|9|videte autem vosmet ipsos tradent enim vos conciliis et in synagogis vapulabitis et ante praesides et reges stabitis propter me in testimonium illis
MARK|13|10|et in omnes gentes primum oportet praedicari evangelium
MARK|13|11|et cum duxerint vos tradentes nolite praecogitare quid loquamini sed quod datum vobis fuerit in illa hora id loquimini non enim estis vos loquentes sed Spiritus Sanctus
MARK|13|12|tradet autem frater fratrem in mortem et pater filium et consurgent filii in parentes et morte adficient eos
MARK|13|13|et eritis odio omnibus propter nomen meum qui autem sustinuerit in finem hic salvus erit
MARK|13|14|cum autem videritis abominationem desolationis stantem ubi non debet qui legit intellegat tunc qui in Iudaea sunt fugiant in montes
MARK|13|15|et qui super tectum ne descendat in domum nec introeat ut tollat quid de domo sua
MARK|13|16|et qui in agro erit non revertatur retro tollere vestimentum suum
MARK|13|17|vae autem praegnatibus et nutrientibus in illis diebus
MARK|13|18|orate vero ut hieme non fiant
MARK|13|19|erunt enim dies illi tribulationes tales quales non fuerunt ab initio creaturae quam condidit Deus usque nunc neque fient
MARK|13|20|et nisi breviasset Dominus dies non fuisset salva omnis caro sed propter electos quos elegit breviavit dies
MARK|13|21|et tunc si quis vobis dixerit ecce hic est Christus ecce illic ne credideritis
MARK|13|22|exsurgent enim pseudochristi et pseudoprophetae et dabunt signa et portenta ad seducendos si potest fieri etiam electos
MARK|13|23|vos ergo videte ecce praedixi vobis omnia
MARK|13|24|sed in illis diebus post tribulationem illam sol contenebrabitur et luna non dabit splendorem suum
MARK|13|25|et erunt stellae caeli decidentes et virtutes quae sunt in caelis movebuntur
MARK|13|26|et tunc videbunt Filium hominis venientem in nubibus cum virtute multa et gloria
MARK|13|27|et tunc mittet angelos suos et congregabit electos suos a quattuor ventis a summo terrae usque ad summum caeli
MARK|13|28|a ficu autem discite parabolam cum iam ramus eius tener fuerit et nata fuerint folia cognoscitis quia in proximo sit aestas
MARK|13|29|sic et vos cum videritis haec fieri scitote quod in proximo sit in ostiis
MARK|13|30|amen dico vobis quoniam non transiet generatio haec donec omnia ista fiant
MARK|13|31|caelum et terra transibunt verba autem mea non transibunt
MARK|13|32|de die autem illo vel hora nemo scit neque angeli in caelo neque Filius nisi Pater
MARK|13|33|videte vigilate et orate nescitis enim quando tempus sit
MARK|13|34|sicut homo qui peregre profectus reliquit domum suam et dedit servis suis potestatem cuiusque operis et ianitori praecipiat ut vigilet
MARK|13|35|vigilate ergo nescitis enim quando dominus domus veniat sero an media nocte an galli cantu an mane
MARK|13|36|ne cum venerit repente inveniat vos dormientes
MARK|13|37|quod autem vobis dico omnibus dico vigilate
MARK|14|1|erat autem pascha et azyma post biduum et quaerebant summi sacerdotes et scribae quomodo eum dolo tenerent et occiderent
MARK|14|2|dicebant enim non in die festo ne forte tumultus fieret populi
MARK|14|3|et cum esset Bethaniae in domo Simonis leprosi et recumberet venit mulier habens alabastrum unguenti nardi spicati pretiosi et fracto alabastro effudit super caput eius
MARK|14|4|erant autem quidam indigne ferentes intra semet ipsos et dicentes ut quid perditio ista unguenti facta est
MARK|14|5|poterat enim unguentum istud veniri plus quam trecentis denariis et dari pauperibus et fremebant in eam
MARK|14|6|Iesus autem dixit sinite eam quid illi molesti estis bonum opus operata est in me
MARK|14|7|semper enim pauperes habetis vobiscum et cum volueritis potestis illis benefacere me autem non semper habetis
MARK|14|8|quod habuit haec fecit praevenit unguere corpus meum in sepulturam
MARK|14|9|amen dico vobis ubicumque praedicatum fuerit evangelium istud in universum mundum et quod fecit haec narrabitur in memoriam eius
MARK|14|10|et Iudas Scariotis unus de duodecim abiit ad summos sacerdotes ut proderet eum illis
MARK|14|11|qui audientes gavisi sunt et promiserunt ei pecuniam se daturos et quaerebat quomodo illum oportune traderet
MARK|14|12|et primo die azymorum quando pascha immolabant dicunt ei discipuli quo vis eamus et paremus tibi ut manduces pascha
MARK|14|13|et mittit duos ex discipulis suis et dicit eis ite in civitatem et occurret vobis homo laguenam aquae baiulans sequimini eum
MARK|14|14|et quocumque introierit dicite domino domus quia magister dicit ubi est refectio mea ubi pascha cum discipulis meis manducem
MARK|14|15|et ipse vobis demonstrabit cenaculum grande stratum et illic parate nobis
MARK|14|16|et abierunt discipuli eius et venerunt in civitatem et invenerunt sicut dixerat illis et praeparaverunt pascha
MARK|14|17|vespere autem facto venit cum duodecim
MARK|14|18|et discumbentibus eis et manducantibus ait Iesus amen dico vobis quia unus ex vobis me tradet qui manducat mecum
MARK|14|19|at illi coeperunt contristari et dicere ei singillatim numquid ego
MARK|14|20|qui ait illis unus ex duodecim qui intinguit mecum in catino
MARK|14|21|et Filius quidem hominis vadit sicut scriptum est de eo vae autem homini illi per quem Filius hominis traditur bonum ei si non esset natus homo ille
MARK|14|22|et manducantibus illis accepit Iesus panem et benedicens fregit et dedit eis et ait sumite hoc est corpus meum
MARK|14|23|et accepto calice gratias agens dedit eis et biberunt ex illo omnes
MARK|14|24|et ait illis hic est sanguis meus novi testamenti qui pro multis effunditur
MARK|14|25|amen dico vobis quod iam non bibam de genimine vitis usque in diem illum cum illud bibam novum in regno Dei
MARK|14|26|et hymno dicto exierunt in montem Olivarum
MARK|14|27|et ait eis Iesus omnes scandalizabimini in nocte ista quia scriptum est percutiam pastorem et dispergentur oves
MARK|14|28|sed posteaquam resurrexero praecedam vos in Galilaeam
MARK|14|29|Petrus autem ait ei et si omnes scandalizati fuerint sed non ego
MARK|14|30|et ait illi Iesus amen dico tibi quia tu hodie in nocte hac priusquam bis gallus vocem dederit ter me es negaturus
MARK|14|31|at ille amplius loquebatur et si oportuerit me simul conmori tibi non te negabo similiter autem et omnes dicebant
MARK|14|32|et veniunt in praedium cui nomen Gethsemani et ait discipulis suis sedete hic donec orem
MARK|14|33|et adsumit Petrum et Iacobum et Iohannem secum et coepit pavere et taedere
MARK|14|34|et ait illis tristis est anima mea usque ad mortem sustinete hic et vigilate
MARK|14|35|et cum processisset paululum procidit super terram et orabat ut si fieri posset transiret ab eo hora
MARK|14|36|et dixit Abba Pater omnia possibilia tibi sunt transfer calicem hunc a me sed non quod ego volo sed quod tu
MARK|14|37|et venit et invenit eos dormientes et ait Petro Simon dormis non potuisti una hora vigilare
MARK|14|38|vigilate et orate ut non intretis in temptationem spiritus quidem promptus caro vero infirma
MARK|14|39|et iterum abiens oravit eundem sermonem dicens
MARK|14|40|et reversus denuo invenit eos dormientes erant enim oculi illorum ingravati et ignorabant quid responderent ei
MARK|14|41|et venit tertio et ait illis dormite iam et requiescite sufficit venit hora ecce traditur Filius hominis in manus peccatorum
MARK|14|42|surgite eamus ecce qui me tradit prope est
MARK|14|43|et adhuc eo loquente venit Iudas Scarioth unus ex duodecim et cum illo turba cum gladiis et lignis a summis sacerdotibus et a scribis et a senioribus
MARK|14|44|dederat autem traditor eius signum eis dicens quemcumque osculatus fuero ipse est tenete eum et ducite
MARK|14|45|et cum venisset statim accedens ad eum ait rabbi et osculatus est eum
MARK|14|46|at illi manus iniecerunt in eum et tenuerunt eum
MARK|14|47|unus autem quidam de circumstantibus educens gladium percussit servum summi sacerdotis et amputavit illi auriculam
MARK|14|48|et respondens Iesus ait illis tamquam ad latronem existis cum gladiis et lignis conprehendere me
MARK|14|49|cotidie eram apud vos in templo docens et non me tenuistis sed ut adimpleantur scripturae
MARK|14|50|tunc discipuli eius relinquentes eum omnes fugerunt
MARK|14|51|adulescens autem quidam sequebatur illum amictus sindone super nudo et tenuerunt eum
MARK|14|52|at ille reiecta sindone nudus profugit ab eis
MARK|14|53|et adduxerunt Iesum ad summum sacerdotem et conveniunt omnes sacerdotes et scribae et seniores
MARK|14|54|Petrus autem a longe secutus est eum usque intro in atrium summi sacerdotis et sedebat cum ministris et calefaciebat se ad ignem
MARK|14|55|summi vero sacerdotes et omne concilium quaerebant adversum Iesum testimonium ut eum morti traderent nec inveniebant
MARK|14|56|multi enim testimonium falsum dicebant adversus eum et convenientia testimonia non erant
MARK|14|57|et quidam surgentes falsum testimonium ferebant adversus eum dicentes
MARK|14|58|quoniam nos audivimus eum dicentem ego dissolvam templum hoc manufactum et per triduum aliud non manufactum aedificabo
MARK|14|59|et non erat conveniens testimonium illorum
MARK|14|60|et exsurgens summus sacerdos in medium interrogavit Iesum dicens non respondes quicquam ad ea quae tibi obiciuntur ab his
MARK|14|61|ille autem tacebat et nihil respondit rursum summus sacerdos interrogabat eum et dicit ei tu es Christus Filius Benedicti
MARK|14|62|Iesus autem dixit illi ego sum et videbitis Filium hominis a dextris sedentem Virtutis et venientem cum nubibus caeli
MARK|14|63|summus autem sacerdos scindens vestimenta sua ait quid adhuc desideramus testes
MARK|14|64|audistis blasphemiam quid vobis videtur qui omnes condemnaverunt eum esse reum mortis
MARK|14|65|et coeperunt quidam conspuere eum et velare faciem eius et colaphis eum caedere et dicere ei prophetiza et ministri alapis eum caedebant
MARK|14|66|et cum esset Petrus in atrio deorsum venit una ex ancillis summi sacerdotis
MARK|14|67|et cum vidisset Petrum calefacientem se aspiciens illum ait et tu cum Iesu Nazareno eras
MARK|14|68|at ille negavit dicens neque scio neque novi quid dicas et exiit foras ante atrium et gallus cantavit
MARK|14|69|rursus autem cum vidisset illum ancilla coepit dicere circumstantibus quia hic ex illis est
MARK|14|70|at ille iterum negavit et post pusillum rursus qui adstabant dicebant Petro vere ex illis es nam et Galilaeus es
MARK|14|71|ille autem coepit anathematizare et iurare quia nescio hominem istum quem dicitis
MARK|14|72|et statim iterum gallus cantavit et recordatus est Petrus verbi quod dixerat ei Iesus priusquam gallus cantet bis ter me negabis et coepit flere
MARK|15|1|et confestim mane consilium facientes summi sacerdotes cum senioribus et scribis et universo concilio vincientes Iesum duxerunt et tradiderunt Pilato
MARK|15|2|et interrogavit eum Pilatus tu es rex Iudaeorum at ille respondens ait illi tu dicis
MARK|15|3|et accusabant eum summi sacerdotes in multis
MARK|15|4|Pilatus autem rursum interrogavit eum dicens non respondes quicquam vide in quantis te accusant
MARK|15|5|Iesus autem amplius nihil respondit ita ut miraretur Pilatus
MARK|15|6|per diem autem festum dimittere solebat illis unum ex vinctis quemcumque petissent
MARK|15|7|erat autem qui dicebatur Barabbas qui cum seditiosis erat vinctus qui in seditione fecerant homicidium
MARK|15|8|et cum ascendisset turba coepit rogare sicut semper faciebat illis
MARK|15|9|Pilatus autem respondit eis et dixit vultis dimittam vobis regem Iudaeorum
MARK|15|10|sciebat enim quod per invidiam tradidissent eum summi sacerdotes
MARK|15|11|pontifices autem concitaverunt turbam ut magis Barabban dimitteret eis
MARK|15|12|Pilatus autem iterum respondens ait illis quid ergo vultis faciam regi Iudaeorum
MARK|15|13|at illi iterum clamaverunt crucifige eum
MARK|15|14|Pilatus vero dicebat eis quid enim mali fecit at illi magis clamabant crucifige eum
MARK|15|15|Pilatus autem volens populo satisfacere dimisit illis Barabban et tradidit Iesum flagellis caesum ut crucifigeretur
MARK|15|16|milites autem duxerunt eum intro in atrium praetorii et convocant totam cohortem
MARK|15|17|et induunt eum purpuram et inponunt ei plectentes spineam coronam
MARK|15|18|et coeperunt salutare eum have rex Iudaeorum
MARK|15|19|et percutiebant caput eius harundine et conspuebant eum et ponentes genua adorabant eum
MARK|15|20|et postquam inluserunt ei exuerunt illum purpuram et induerunt eum vestimentis suis et educunt illum ut crucifigerent eum
MARK|15|21|et angariaverunt praetereuntem quempiam Simonem Cyreneum venientem de villa patrem Alexandri et Rufi ut tolleret crucem eius
MARK|15|22|et perducunt illum in Golgotha locum quod est interpretatum Calvariae locus
MARK|15|23|et dabant ei bibere murratum vinum et non accepit
MARK|15|24|et crucifigentes eum diviserunt vestimenta eius mittentes sortem super eis quis quid tolleret
MARK|15|25|erat autem hora tertia et crucifixerunt eum
MARK|15|26|et erat titulus causae eius inscriptus rex Iudaeorum
MARK|15|27|et cum eo crucifigunt duos latrones unum a dextris et alium a sinistris eius
MARK|15|28|et adimpleta est scriptura quae dicit et cum iniquis reputatus est
MARK|15|29|et praetereuntes blasphemabant eum moventes capita sua et dicentes va qui destruit templum et in tribus diebus aedificat
MARK|15|30|salvum fac temet ipsum descendens de cruce
MARK|15|31|similiter et summi sacerdotes ludentes ad alterutrum cum scribis dicebant alios salvos fecit se ipsum non potest salvum facere
MARK|15|32|Christus rex Israhel descendat nunc de cruce ut videamus et credamus et qui cum eo crucifixi erant conviciabantur ei
MARK|15|33|et facta hora sexta tenebrae factae sunt per totam terram usque in horam nonam
MARK|15|34|et hora nona exclamavit Iesus voce magna dicens Heloi Heloi lama sabacthani quod est interpretatum Deus meus Deus meus ut quid dereliquisti me
MARK|15|35|et quidam de circumstantibus audientes dicebant ecce Heliam vocat
MARK|15|36|currens autem unus et implens spongiam aceto circumponensque calamo potum dabat ei dicens sinite videamus si veniat Helias ad deponendum eum
MARK|15|37|Iesus autem emissa voce magna exspiravit
MARK|15|38|et velum templi scissum est in duo a sursum usque deorsum
MARK|15|39|videns autem centurio qui ex adverso stabat quia sic clamans exspirasset ait vere homo hic Filius Dei erat
MARK|15|40|erant autem et mulieres de longe aspicientes inter quas et Maria Magdalene et Maria Iacobi minoris et Ioseph mater et Salome
MARK|15|41|et cum esset in Galilaea sequebantur eum et ministrabant ei et aliae multae quae simul cum eo ascenderant Hierosolyma
MARK|15|42|et cum iam sero esset factum quia erat parasceve quod est ante sabbatum
MARK|15|43|venit Ioseph ab Arimathia nobilis decurio qui et ipse erat expectans regnum Dei et audacter introiit ad Pilatum et petiit corpus Iesu
MARK|15|44|Pilatus autem mirabatur si iam obisset et accersito centurione interrogavit eum si iam mortuus esset
MARK|15|45|et cum cognovisset a centurione donavit corpus Ioseph
MARK|15|46|Ioseph autem mercatus sindonem et deponens eum involvit sindone et posuit eum in monumento quod erat excisum de petra et advolvit lapidem ad ostium monumenti
MARK|15|47|Maria autem Magdalene et Maria Ioseph aspiciebant ubi poneretur
MARK|16|1|et cum transisset sabbatum Maria Magdalene et Maria Iacobi et Salome emerunt aromata ut venientes unguerent eum
MARK|16|2|et valde mane una sabbatorum veniunt ad monumentum orto iam sole
MARK|16|3|et dicebant ad invicem quis revolvet nobis lapidem ab ostio monumenti
MARK|16|4|et respicientes vident revolutum lapidem erat quippe magnus valde
MARK|16|5|et introeuntes in monumento viderunt iuvenem sedentem in dextris coopertum stola candida et obstipuerunt
MARK|16|6|qui dicit illis nolite expavescere Iesum quaeritis Nazarenum crucifixum surrexit non est hic ecce locus ubi posuerunt eum
MARK|16|7|sed ite et dicite discipulis eius et Petro quia praecedit vos in Galilaeam ibi eum videbitis sicut dixit vobis
MARK|16|8|at illae exeuntes fugerunt de monumento invaserat enim eas tremor et pavor et nemini quicquam dixerunt timebant enim
MARK|16|9|surgens autem mane prima sabbati apparuit primo Mariae Magdalenae de qua eiecerat septem daemonia
MARK|16|10|illa vadens nuntiavit his qui cum eo fuerant lugentibus et flentibus
MARK|16|11|et illi audientes quia viveret et visus esset ab ea non crediderunt
MARK|16|12|post haec autem duobus ex eis ambulantibus ostensus est in alia effigie euntibus in villam
MARK|16|13|et illi euntes nuntiaverunt ceteris nec illis crediderunt
MARK|16|14|novissime recumbentibus illis undecim apparuit et exprobravit incredulitatem illorum et duritiam cordis quia his qui viderant eum resurrexisse non crediderant
MARK|16|15|et dixit eis euntes in mundum universum praedicate evangelium omni creaturae
MARK|16|16|qui crediderit et baptizatus fuerit salvus erit qui vero non crediderit condemnabitur
MARK|16|17|signa autem eos qui crediderint haec sequentur in nomine meo daemonia eicient linguis loquentur novis
MARK|16|18|serpentes tollent et si mortiferum quid biberint non eos nocebit super aegrotos manus inponent et bene habebunt
MARK|16|19|et Dominus quidem postquam locutus est eis adsumptus est in caelum et sedit a dextris Dei
MARK|16|20|illi autem profecti praedicaverunt ubique Domino cooperante et sermonem confirmante sequentibus signis
LUKE|1|1|quoniam quidem multi conati sunt ordinare narrationem quae in nobis conpletae sunt rerum
LUKE|1|2|sicut tradiderunt nobis qui ab initio ipsi viderunt et ministri fuerunt sermonis
LUKE|1|3|visum est et mihi adsecuto a principio omnibus diligenter ex ordine tibi scribere optime Theophile
LUKE|1|4|ut cognoscas eorum verborum de quibus eruditus es veritatem
LUKE|1|5|fuit in diebus Herodis regis Iudaeae sacerdos quidam nomine Zaccharias de vice Abia et uxor illi de filiabus Aaron et nomen eius Elisabeth
LUKE|1|6|erant autem iusti ambo ante Deum incedentes in omnibus mandatis et iustificationibus Domini sine querella
LUKE|1|7|et non erat illis filius eo quod esset Elisabeth sterilis et ambo processissent in diebus suis
LUKE|1|8|factum est autem cum sacerdotio fungeretur in ordine vicis suae ante Deum
LUKE|1|9|secundum consuetudinem sacerdotii sorte exiit ut incensum poneret ingressus in templum Domini
LUKE|1|10|et omnis multitudo erat populi orans foris hora incensi
LUKE|1|11|apparuit autem illi angelus Domini stans a dextris altaris incensi
LUKE|1|12|et Zaccharias turbatus est videns et timor inruit super eum
LUKE|1|13|ait autem ad illum angelus ne timeas Zaccharia quoniam exaudita est deprecatio tua et uxor tua Elisabeth pariet tibi filium et vocabis nomen eius Iohannem
LUKE|1|14|et erit gaudium tibi et exultatio et multi in nativitate eius gaudebunt
LUKE|1|15|erit enim magnus coram Domino et vinum et sicera non bibet et Spiritu Sancto replebitur adhuc ex utero matris suae
LUKE|1|16|et multos filiorum Israhel convertet ad Dominum Deum ipsorum
LUKE|1|17|et ipse praecedet ante illum in spiritu et virtute Heliae ut convertat corda patrum in filios et incredibiles ad prudentiam iustorum parare Domino plebem perfectam
LUKE|1|18|et dixit Zaccharias ad angelum unde hoc sciam ego enim sum senex et uxor mea processit in diebus suis
LUKE|1|19|et respondens angelus dixit ei ego sum Gabrihel qui adsto ante Deum et missus sum loqui ad te et haec tibi evangelizare
LUKE|1|20|et ecce eris tacens et non poteris loqui usque in diem quo haec fiant pro eo quod non credidisti verbis meis quae implebuntur in tempore suo
LUKE|1|21|et erat plebs expectans Zacchariam et mirabantur quod tardaret ipse in templo
LUKE|1|22|egressus autem non poterat loqui ad illos et cognoverunt quod visionem vidisset in templo et ipse erat innuens illis et permansit mutus
LUKE|1|23|et factum est ut impleti sunt dies officii eius abiit in domum suam
LUKE|1|24|post hos autem dies concepit Elisabeth uxor eius et occultabat se mensibus quinque dicens
LUKE|1|25|quia sic mihi fecit Dominus in diebus quibus respexit auferre obprobrium meum inter homines
LUKE|1|26|in mense autem sexto missus est angelus Gabrihel a Deo in civitatem Galilaeae cui nomen Nazareth
LUKE|1|27|ad virginem desponsatam viro cui nomen erat Ioseph de domo David et nomen virginis Maria
LUKE|1|28|et ingressus angelus ad eam dixit have gratia plena Dominus tecum benedicta tu in mulieribus
LUKE|1|29|quae cum vidisset turbata est in sermone eius et cogitabat qualis esset ista salutatio
LUKE|1|30|et ait angelus ei ne timeas Maria invenisti enim gratiam apud Deum
LUKE|1|31|ecce concipies in utero et paries filium et vocabis nomen eius Iesum
LUKE|1|32|hic erit magnus et Filius Altissimi vocabitur et dabit illi Dominus Deus sedem David patris eius
LUKE|1|33|et regnabit in domo Iacob in aeternum et regni eius non erit finis
LUKE|1|34|dixit autem Maria ad angelum quomodo fiet istud quoniam virum non cognosco
LUKE|1|35|et respondens angelus dixit ei Spiritus Sanctus superveniet in te et virtus Altissimi obumbrabit tibi ideoque et quod nascetur sanctum vocabitur Filius Dei
LUKE|1|36|et ecce Elisabeth cognata tua et ipsa concepit filium in senecta sua et hic mensis est sextus illi quae vocatur sterilis
LUKE|1|37|quia non erit inpossibile apud Deum omne verbum
LUKE|1|38|dixit autem Maria ecce ancilla Domini fiat mihi secundum verbum tuum et discessit ab illa angelus
LUKE|1|39|exsurgens autem Maria in diebus illis abiit in montana cum festinatione in civitatem Iuda
LUKE|1|40|et intravit in domum Zacchariae et salutavit Elisabeth
LUKE|1|41|et factum est ut audivit salutationem Mariae Elisabeth exultavit infans in utero eius et repleta est Spiritu Sancto Elisabeth
LUKE|1|42|et exclamavit voce magna et dixit benedicta tu inter mulieres et benedictus fructus ventris tui
LUKE|1|43|et unde hoc mihi ut veniat mater Domini mei ad me
LUKE|1|44|ecce enim ut facta est vox salutationis tuae in auribus meis exultavit in gaudio infans in utero meo
LUKE|1|45|et beata quae credidit quoniam perficientur ea quae dicta sunt ei a Domino
LUKE|1|46|et ait Maria magnificat anima mea Dominum
LUKE|1|47|et exultavit spiritus meus in Deo salutari meo
LUKE|1|48|quia respexit humilitatem ancillae suae ecce enim ex hoc beatam me dicent omnes generationes
LUKE|1|49|quia fecit mihi magna qui potens est et sanctum nomen eius
LUKE|1|50|et misericordia eius in progenies et progenies timentibus eum
LUKE|1|51|fecit potentiam in brachio suo dispersit superbos mente cordis sui
LUKE|1|52|deposuit potentes de sede et exaltavit humiles
LUKE|1|53|esurientes implevit bonis et divites dimisit inanes
LUKE|1|54|suscepit Israhel puerum suum memorari misericordiae
LUKE|1|55|sicut locutus est ad patres nostros Abraham et semini eius in saecula
LUKE|1|56|mansit autem Maria cum illa quasi mensibus tribus et reversa est in domum suam
LUKE|1|57|Elisabeth autem impletum est tempus pariendi et peperit filium
LUKE|1|58|et audierunt vicini et cognati eius quia magnificavit Dominus misericordiam suam cum illa et congratulabantur ei
LUKE|1|59|et factum est in die octavo venerunt circumcidere puerum et vocabant eum nomine patris eius Zacchariam
LUKE|1|60|et respondens mater eius dixit nequaquam sed vocabitur Iohannes
LUKE|1|61|et dixerunt ad illam quia nemo est in cognatione tua qui vocetur hoc nomine
LUKE|1|62|innuebant autem patri eius quem vellet vocari eum
LUKE|1|63|et postulans pugillarem scripsit dicens Iohannes est nomen eius et mirati sunt universi
LUKE|1|64|apertum est autem ilico os eius et lingua eius et loquebatur benedicens Deum
LUKE|1|65|et factus est timor super omnes vicinos eorum et super omnia montana Iudaeae divulgabantur omnia verba haec
LUKE|1|66|et posuerunt omnes qui audierant in corde suo dicentes quid putas puer iste erit etenim manus Domini erat cum illo
LUKE|1|67|et Zaccharias pater eius impletus est Spiritu Sancto et prophetavit dicens
LUKE|1|68|benedictus Deus Israhel quia visitavit et fecit redemptionem plebi suae
LUKE|1|69|et erexit cornu salutis nobis in domo David pueri sui
LUKE|1|70|sicut locutus est per os sanctorum qui a saeculo sunt prophetarum eius
LUKE|1|71|salutem ex inimicis nostris et de manu omnium qui oderunt nos
LUKE|1|72|ad faciendam misericordiam cum patribus nostris et memorari testamenti sui sancti
LUKE|1|73|iusiurandum quod iuravit ad Abraham patrem nostrum
LUKE|1|74|daturum se nobis ut sine timore de manu inimicorum nostrorum liberati serviamus illi
LUKE|1|75|in sanctitate et iustitia coram ipso omnibus diebus nostris
LUKE|1|76|et tu puer propheta Altissimi vocaberis praeibis enim ante faciem Domini parare vias eius
LUKE|1|77|ad dandam scientiam salutis plebi eius in remissionem peccatorum eorum
LUKE|1|78|per viscera misericordiae Dei nostri in quibus visitavit nos oriens ex alto
LUKE|1|79|inluminare his qui in tenebris et in umbra mortis sedent ad dirigendos pedes nostros in viam pacis
LUKE|1|80|puer autem crescebat et confortabatur spiritu et erat in deserto usque in diem ostensionis suae ad Israhel
LUKE|2|1|factum est autem in diebus illis exiit edictum a Caesare Augusto ut describeretur universus orbis
LUKE|2|2|haec descriptio prima facta est praeside Syriae Cyrino
LUKE|2|3|et ibant omnes ut profiterentur singuli in suam civitatem
LUKE|2|4|ascendit autem et Ioseph a Galilaea de civitate Nazareth in Iudaeam civitatem David quae vocatur Bethleem eo quod esset de domo et familia David
LUKE|2|5|ut profiteretur cum Maria desponsata sibi uxore praegnate
LUKE|2|6|factum est autem cum essent ibi impleti sunt dies ut pareret
LUKE|2|7|et peperit filium suum primogenitum et pannis eum involvit et reclinavit eum in praesepio quia non erat eis locus in diversorio
LUKE|2|8|et pastores erant in regione eadem vigilantes et custodientes vigilias noctis supra gregem suum
LUKE|2|9|et ecce angelus Domini stetit iuxta illos et claritas Dei circumfulsit illos et timuerunt timore magno
LUKE|2|10|et dixit illis angelus nolite timere ecce enim evangelizo vobis gaudium magnum quod erit omni populo
LUKE|2|11|quia natus est vobis hodie salvator qui est Christus Dominus in civitate David
LUKE|2|12|et hoc vobis signum invenietis infantem pannis involutum et positum in praesepio
LUKE|2|13|et subito facta est cum angelo multitudo militiae caelestis laudantium Deum et dicentium
LUKE|2|14|gloria in altissimis Deo et in terra pax in hominibus bonae voluntatis
LUKE|2|15|et factum est ut discesserunt ab eis angeli in caelum pastores loquebantur ad invicem transeamus usque Bethleem et videamus hoc verbum quod factum est quod fecit Dominus et ostendit nobis
LUKE|2|16|et venerunt festinantes et invenerunt Mariam et Ioseph et infantem positum in praesepio
LUKE|2|17|videntes autem cognoverunt de verbo quod dictum erat illis de puero hoc
LUKE|2|18|et omnes qui audierunt mirati sunt et de his quae dicta erant a pastoribus ad ipsos
LUKE|2|19|Maria autem conservabat omnia verba haec conferens in corde suo
LUKE|2|20|et reversi sunt pastores glorificantes et laudantes Deum in omnibus quae audierant et viderant sicut dictum est ad illos
LUKE|2|21|et postquam consummati sunt dies octo ut circumcideretur vocatum est nomen eius Iesus quod vocatum est ab angelo priusquam in utero conciperetur
LUKE|2|22|et postquam impleti sunt dies purgationis eius secundum legem Mosi tulerunt illum in Hierusalem ut sisterent eum Domino
LUKE|2|23|sicut scriptum est in lege Domini quia omne masculinum adaperiens vulvam sanctum Domino vocabitur
LUKE|2|24|et ut darent hostiam secundum quod dictum est in lege Domini par turturum aut duos pullos columbarum
LUKE|2|25|et ecce homo erat in Hierusalem cui nomen Symeon et homo iste iustus et timoratus expectans consolationem Israhel et Spiritus Sanctus erat in eo
LUKE|2|26|et responsum acceperat ab Spiritu Sancto non visurum se mortem nisi prius videret Christum Domini
LUKE|2|27|et venit in Spiritu in templum et cum inducerent puerum Iesum parentes eius ut facerent secundum consuetudinem legis pro eo
LUKE|2|28|et ipse accepit eum in ulnas suas et benedixit Deum et dixit
LUKE|2|29|nunc dimittis servum tuum Domine secundum verbum tuum in pace
LUKE|2|30|quia viderunt oculi mei salutare tuum
LUKE|2|31|quod parasti ante faciem omnium populorum
LUKE|2|32|lumen ad revelationem gentium et gloriam plebis tuae Israhel
LUKE|2|33|et erat pater eius et mater mirantes super his quae dicebantur de illo
LUKE|2|34|et benedixit illis Symeon et dixit ad Mariam matrem eius ecce positus est hic in ruinam et resurrectionem multorum in Israhel et in signum cui contradicetur
LUKE|2|35|et tuam ipsius animam pertransiet gladius ut revelentur ex multis cordibus cogitationes
LUKE|2|36|et erat Anna prophetissa filia Phanuhel de tribu Aser haec processerat in diebus multis et vixerat cum viro suo annis septem a virginitate sua
LUKE|2|37|et haec vidua usque ad annos octoginta quattuor quae non discedebat de templo ieiuniis et obsecrationibus serviens nocte ac die
LUKE|2|38|et haec ipsa hora superveniens confitebatur Domino et loquebatur de illo omnibus qui expectabant redemptionem Hierusalem
LUKE|2|39|et ut perfecerunt omnia secundum legem Domini reversi sunt in Galilaeam in civitatem suam Nazareth
LUKE|2|40|puer autem crescebat et confortabatur plenus sapientia et gratia Dei erat in illo
LUKE|2|41|et ibant parentes eius per omnes annos in Hierusalem in die sollemni paschae
LUKE|2|42|et cum factus esset annorum duodecim ascendentibus illis in Hierosolymam secundum consuetudinem diei festi
LUKE|2|43|consummatisque diebus cum redirent remansit puer Iesus in Hierusalem et non cognoverunt parentes eius
LUKE|2|44|existimantes autem illum esse in comitatu venerunt iter diei et requirebant eum inter cognatos et notos
LUKE|2|45|et non invenientes regressi sunt in Hierusalem requirentes eum
LUKE|2|46|et factum est post triduum invenerunt illum in templo sedentem in medio doctorum audientem illos et interrogantem
LUKE|2|47|stupebant autem omnes qui eum audiebant super prudentia et responsis eius
LUKE|2|48|et videntes admirati sunt et dixit mater eius ad illum fili quid fecisti nobis sic ecce pater tuus et ego dolentes quaerebamus te
LUKE|2|49|et ait ad illos quid est quod me quaerebatis nesciebatis quia in his quae Patris mei sunt oportet me esse
LUKE|2|50|et ipsi non intellexerunt verbum quod locutus est ad illos
LUKE|2|51|et descendit cum eis et venit Nazareth et erat subditus illis et mater eius conservabat omnia verba haec in corde suo
LUKE|2|52|et Iesus proficiebat sapientia aetate et gratia apud Deum et homines
LUKE|3|1|anno autem quintodecimo imperii Tiberii Caesaris procurante Pontio Pilato Iudaeam tetrarcha autem Galilaeae Herode Philippo autem fratre eius tetrarcha Itureae et Trachonitidis regionis et Lysania Abilinae tetrarcha
LUKE|3|2|sub principibus sacerdotum Anna et Caiapha factum est verbum Dei super Iohannem Zacchariae filium in deserto
LUKE|3|3|et venit in omnem regionem Iordanis praedicans baptismum paenitentiae in remissionem peccatorum
LUKE|3|4|sicut scriptum est in libro sermonum Esaiae prophetae vox clamantis in deserto parate viam Domini rectas facite semitas eius
LUKE|3|5|omnis vallis implebitur et omnis mons et collis humiliabitur et erunt prava in directa et aspera in vias planas
LUKE|3|6|et videbit omnis caro salutare Dei
LUKE|3|7|dicebat ergo ad turbas quae exiebant ut baptizarentur ab ipso genimina viperarum quis ostendit vobis fugere a ventura ira
LUKE|3|8|facite ergo fructus dignos paenitentiae et ne coeperitis dicere patrem habemus Abraham dico enim vobis quia potest Deus de lapidibus istis suscitare filios Abrahae
LUKE|3|9|iam enim securis ad radicem arborum posita est omnis ergo arbor non faciens fructum exciditur et in ignem mittitur
LUKE|3|10|et interrogabant eum turbae dicentes quid ergo faciemus
LUKE|3|11|respondens autem dicebat illis qui habet duas tunicas det non habenti et qui habet escas similiter faciat
LUKE|3|12|venerunt autem et publicani ut baptizarentur et dixerunt ad illum magister quid faciemus
LUKE|3|13|at ille dixit ad eos nihil amplius quam quod constitutum est vobis faciatis
LUKE|3|14|interrogabant autem eum et milites dicentes quid faciemus et nos et ait illis neminem concutiatis neque calumniam faciatis et contenti estote stipendiis vestris
LUKE|3|15|existimante autem populo et cogitantibus omnibus in cordibus suis de Iohanne ne forte ipse esset Christus
LUKE|3|16|respondit Iohannes dicens omnibus ego quidem aqua baptizo vos venit autem fortior me cuius non sum dignus solvere corrigiam calciamentorum eius ipse vos baptizabit in Spiritu Sancto et igni
LUKE|3|17|cuius ventilabrum in manu eius et purgabit aream suam et congregabit triticum in horreum suum paleas autem conburet igni inextinguibili
LUKE|3|18|multa quidem et alia exhortans evangelizabat populum
LUKE|3|19|Herodes autem tetrarcha cum corriperetur ab illo de Herodiade uxore fratris sui et de omnibus malis quae fecit Herodes
LUKE|3|20|adiecit et hoc supra omnia et inclusit Iohannem in carcere
LUKE|3|21|factum est autem cum baptizaretur omnis populus et Iesu baptizato et orante apertum est caelum
LUKE|3|22|et descendit Spiritus Sanctus corporali specie sicut columba in ipsum et vox de caelo facta est tu es Filius meus dilectus in te conplacuit mihi
LUKE|3|23|et ipse Iesus erat incipiens quasi annorum triginta ut putabatur filius Ioseph qui fuit Heli
LUKE|3|24|qui fuit Matthat qui fuit Levi qui fuit Melchi qui fuit Iannae qui fuit Ioseph
LUKE|3|25|qui fuit Matthathiae qui fuit Amos qui fuit Naum qui fuit Esli qui fuit Naggae
LUKE|3|26|qui fuit Maath qui fuit Matthathiae qui fuit Semei qui fuit Iosech qui fuit Ioda
LUKE|3|27|qui fuit Iohanna qui fuit Resa qui fuit Zorobabel qui fuit Salathihel qui fuit Neri
LUKE|3|28|qui fuit Melchi qui fuit Addi qui fuit Cosam qui fuit Helmadam qui fuit Her
LUKE|3|29|qui fuit Iesu qui fuit Eliezer qui fuit Iorim qui fuit Matthat qui fuit Levi
LUKE|3|30|qui fuit Symeon qui fuit Iuda qui fuit Ioseph qui fuit Iona qui fuit Eliachim
LUKE|3|31|qui fuit Melea qui fuit Menna qui fuit Matthata qui fuit Nathan qui fuit David
LUKE|3|32|qui fuit Iesse qui fuit Obed qui fuit Booz qui fuit Salmon qui fuit Naasson
LUKE|3|33|qui fuit Aminadab qui fuit Aram qui fuit Esrom qui fuit Phares qui fuit Iudae
LUKE|3|34|qui fuit Iacob qui fuit Isaac qui fuit Abraham qui fuit Thare qui fuit Nachor
LUKE|3|35|qui fuit Seruch qui fuit Ragau qui fuit Phalec qui fuit Eber qui fuit Sale
LUKE|3|36|qui fuit Cainan qui fuit Arfaxat qui fuit Sem qui fuit Noe qui fuit Lamech
LUKE|3|37|qui fuit Mathusalae qui fuit Enoch qui fuit Iared qui fuit Malelehel qui fuit Cainan
LUKE|3|38|qui fuit Enos qui fuit Seth qui fuit Adam qui fuit Dei
LUKE|4|1|Iesus autem plenus Spiritu Sancto regressus est ab Iordane et agebatur in Spiritu in desertum
LUKE|4|2|diebus quadraginta et temptabatur a diabolo et nihil manducavit in diebus illis et consummatis illis esuriit
LUKE|4|3|dixit autem illi diabolus si Filius Dei es dic lapidi huic ut panis fiat
LUKE|4|4|et respondit ad illum Iesus scriptum est quia non in pane solo vivet homo sed in omni verbo Dei
LUKE|4|5|et duxit illum diabolus et ostendit illi omnia regna orbis terrae in momento temporis
LUKE|4|6|et ait ei tibi dabo potestatem hanc universam et gloriam illorum quia mihi tradita sunt et cui volo do illa
LUKE|4|7|tu ergo si adoraveris coram me erunt tua omnia
LUKE|4|8|et respondens Iesus dixit illi scriptum est Dominum Deum tuum adorabis et illi soli servies
LUKE|4|9|et duxit illum in Hierusalem et statuit eum supra pinnam templi et dixit illi si Filius Dei es mitte te hinc deorsum
LUKE|4|10|scriptum est enim quod angelis suis mandabit de te ut conservent te
LUKE|4|11|et quia in manibus tollent te ne forte offendas ad lapidem pedem tuum
LUKE|4|12|et respondens Iesus ait illi dictum est non temptabis Dominum Deum tuum
LUKE|4|13|et consummata omni temptatione diabolus recessit ab illo usque ad tempus
LUKE|4|14|et regressus est Iesus in virtute Spiritus in Galilaeam et fama exiit per universam regionem de illo
LUKE|4|15|et ipse docebat in synagogis eorum et magnificabatur ab omnibus
LUKE|4|16|et venit Nazareth ubi erat nutritus et intravit secundum consuetudinem suam die sabbati in synagogam et surrexit legere
LUKE|4|17|et traditus est illi liber prophetae Esaiae et ut revolvit librum invenit locum ubi scriptum erat
LUKE|4|18|Spiritus Domini super me propter quod unxit me evangelizare pauperibus misit me
LUKE|4|19|praedicare captivis remissionem et caecis visum dimittere confractos in remissionem praedicare annum Domini acceptum et diem retributionis
LUKE|4|20|et cum plicuisset librum reddidit ministro et sedit et omnium in synagoga oculi erant intendentes in eum
LUKE|4|21|coepit autem dicere ad illos quia hodie impleta est haec scriptura in auribus vestris
LUKE|4|22|et omnes testimonium illi dabant et mirabantur in verbis gratiae quae procedebant de ore ipsius et dicebant nonne hic filius est Ioseph
LUKE|4|23|et ait illis utique dicetis mihi hanc similitudinem medice cura te ipsum quanta audivimus facta in Capharnaum fac et hic in patria tua
LUKE|4|24|ait autem amen dico vobis quia nemo propheta acceptus est in patria sua
LUKE|4|25|in veritate dico vobis multae viduae erant in diebus Heliae in Israhel quando clusum est caelum annis tribus et mensibus sex cum facta est fames magna in omni terra
LUKE|4|26|et ad nullam illarum missus est Helias nisi in Sareptha Sidoniae ad mulierem viduam
LUKE|4|27|et multi leprosi erant in Israhel sub Heliseo propheta et nemo eorum mundatus est nisi Neman Syrus
LUKE|4|28|et repleti sunt omnes in synagoga ira haec audientes
LUKE|4|29|et surrexerunt et eiecerunt illum extra civitatem et duxerunt illum usque ad supercilium montis supra quem civitas illorum erat aedificata ut praecipitarent eum
LUKE|4|30|ipse autem transiens per medium illorum ibat
LUKE|4|31|et descendit in Capharnaum civitatem Galilaeae ibique docebat illos sabbatis
LUKE|4|32|et stupebant in doctrina eius quia in potestate erat sermo ipsius
LUKE|4|33|et in synagoga erat homo habens daemonium inmundum et exclamavit voce magna
LUKE|4|34|dicens sine quid nobis et tibi Iesu Nazarene venisti perdere nos scio te qui sis Sanctus Dei
LUKE|4|35|et increpavit illi Iesus dicens obmutesce et exi ab illo et cum proiecisset illum daemonium in medium exiit ab illo nihilque illum nocuit
LUKE|4|36|et factus est pavor in omnibus et conloquebantur ad invicem dicentes quod est hoc verbum quia in potestate et virtute imperat inmundis spiritibus et exeunt
LUKE|4|37|et divulgabatur fama de illo in omnem locum regionis
LUKE|4|38|surgens autem de synagoga introivit in domum Simonis socrus autem Simonis tenebatur magnis febribus et rogaverunt illum pro ea
LUKE|4|39|et stans super illam imperavit febri et dimisit illam et continuo surgens ministrabat illis
LUKE|4|40|cum sol autem occidisset omnes qui habebant infirmos variis languoribus ducebant illos ad eum at ille singulis manus inponens curabat eos
LUKE|4|41|exiebant autem etiam daemonia a multis clamantia et dicentia quia tu es Filius Dei et increpans non sinebat ea loqui quia sciebant ipsum esse Christum
LUKE|4|42|facta autem die egressus ibat in desertum locum et turbae requirebant eum et venerunt usque ad ipsum et detinebant illum ne discederet ab eis
LUKE|4|43|quibus ille ait quia et aliis civitatibus oportet me evangelizare regnum Dei quia ideo missus sum
LUKE|4|44|et erat praedicans in synagogis Galilaeae
LUKE|5|1|factum est autem cum turbae inruerent in eum ut audirent verbum Dei et ipse stabat secus stagnum Gennesareth
LUKE|5|2|et vidit duas naves stantes secus stagnum piscatores autem descenderant et lavabant retia
LUKE|5|3|ascendens autem in unam navem quae erat Simonis rogavit eum a terra reducere pusillum et sedens docebat de navicula turbas
LUKE|5|4|ut cessavit autem loqui dixit ad Simonem duc in altum et laxate retia vestra in capturam
LUKE|5|5|et respondens Simon dixit illi praeceptor per totam noctem laborantes nihil cepimus in verbo autem tuo laxabo rete
LUKE|5|6|et cum hoc fecissent concluserunt piscium multitudinem copiosam rumpebatur autem rete eorum
LUKE|5|7|et annuerunt sociis qui erant in alia navi ut venirent et adiuvarent eos et venerunt et impleverunt ambas naviculas ita ut mergerentur
LUKE|5|8|quod cum videret Simon Petrus procidit ad genua Iesu dicens exi a me quia homo peccator sum Domine
LUKE|5|9|stupor enim circumdederat eum et omnes qui cum illo erant in captura piscium quam ceperant
LUKE|5|10|similiter autem Iacobum et Iohannem filios Zebedaei qui erant socii Simonis et ait ad Simonem Iesus noli timere ex hoc iam homines eris capiens
LUKE|5|11|et subductis ad terram navibus relictis omnibus secuti sunt illum
LUKE|5|12|et factum est cum esset in una civitatum et ecce vir plenus lepra et videns Iesum et procidens in faciem rogavit eum dicens Domine si vis potes me mundare
LUKE|5|13|et extendens manum tetigit illum dicens volo mundare et confestim lepra discessit ab illo
LUKE|5|14|et ipse praecepit illi ut nemini diceret sed vade ostende te sacerdoti et offer pro emundatione tua sicut praecepit Moses in testimonium illis
LUKE|5|15|perambulabat autem magis sermo de illo et conveniebant turbae multae ut audirent et curarentur ab infirmitatibus suis
LUKE|5|16|ipse autem secedebat in deserto et orabat
LUKE|5|17|et factum est in una dierum et ipse sedebat docens et erant Pharisaei sedentes et legis doctores qui venerant ex omni castello Galilaeae et Iudaeae et Hierusalem et virtus erat Domini ad sanandum eos
LUKE|5|18|et ecce viri portantes in lecto hominem qui erat paralyticus et quaerebant eum inferre et ponere ante eum
LUKE|5|19|et non invenientes qua parte illum inferrent prae turba ascenderunt supra tectum per tegulas submiserunt illum cum lecto in medium ante Iesum
LUKE|5|20|quorum fidem ut vidit dixit homo remittuntur tibi peccata tua
LUKE|5|21|et coeperunt cogitare scribae et Pharisaei dicentes quis est hic qui loquitur blasphemias quis potest dimittere peccata nisi solus Deus
LUKE|5|22|ut cognovit autem Iesus cogitationes eorum respondens dixit ad illos quid cogitatis in cordibus vestris
LUKE|5|23|quid est facilius dicere dimittuntur tibi peccata an dicere surge et ambula
LUKE|5|24|ut autem sciatis quia Filius hominis potestatem habet in terra dimittere peccata ait paralytico tibi dico surge tolle lectum tuum et vade in domum tuam
LUKE|5|25|et confestim surgens coram illis tulit in quo iacebat et abiit in domum suam magnificans Deum
LUKE|5|26|et stupor adprehendit omnes et magnificabant Deum et repleti sunt timore dicentes quia vidimus mirabilia hodie
LUKE|5|27|et post haec exiit et vidit publicanum nomine Levi sedentem ad teloneum et ait illi sequere me
LUKE|5|28|et relictis omnibus surgens secutus est eum
LUKE|5|29|et fecit ei convivium magnum Levi in domo sua et erat turba multa publicanorum et aliorum qui cum illis erant discumbentes
LUKE|5|30|et murmurabant Pharisaei et scribae eorum dicentes ad discipulos eius quare cum publicanis et peccatoribus manducatis et bibitis
LUKE|5|31|et respondens Iesus dixit ad illos non egent qui sani sunt medico sed qui male habent
LUKE|5|32|non veni vocare iustos sed peccatores in paenitentiam
LUKE|5|33|at illi dixerunt ad eum quare discipuli Iohannis ieiunant frequenter et obsecrationes faciunt similiter et Pharisaeorum tui autem edunt et bibunt
LUKE|5|34|quibus ipse ait numquid potestis filios sponsi dum cum illis est sponsus facere ieiunare
LUKE|5|35|venient autem dies et cum ablatus fuerit ab illis sponsus tunc ieiunabunt in illis diebus
LUKE|5|36|dicebat autem et similitudinem ad illos quia nemo commissuram a vestimento novo inmittit in vestimentum vetus alioquin et novum rumpit et veteri non convenit commissura a novo
LUKE|5|37|et nemo mittit vinum novum in utres veteres alioquin rumpet vinum novum utres et ipsum effundetur et utres peribunt
LUKE|5|38|sed vinum novum in utres novos mittendum est et utraque conservantur
LUKE|5|39|et nemo bibens vetus statim vult novum dicit enim vetus melius est
LUKE|6|1|factum est autem in sabbato secundoprimo cum transiret per sata vellebant discipuli eius spicas et manducabant confricantes manibus
LUKE|6|2|quidam autem Pharisaeorum dicebant illis quid facitis quod non licet in sabbatis
LUKE|6|3|et respondens Iesus ad eos dixit nec hoc legistis quod fecit David cum esurisset ipse et qui cum eo erant
LUKE|6|4|quomodo intravit in domum Dei et panes propositionis sumpsit et manducavit et dedit his qui cum ipso erant quos non licet manducare nisi tantum sacerdotibus
LUKE|6|5|et dicebat illis quia dominus est Filius hominis etiam sabbati
LUKE|6|6|factum est autem et in alio sabbato ut intraret in synagogam et doceret et erat ibi homo et manus eius dextra erat arida
LUKE|6|7|observabant autem scribae et Pharisaei si in sabbato curaret ut invenirent accusare illum
LUKE|6|8|ipse vero sciebat cogitationes eorum et ait homini qui habebat manum aridam surge et sta in medium et surgens stetit
LUKE|6|9|ait autem ad illos Iesus interrogo vos si licet sabbato bene facere an male animam salvam facere an perdere
LUKE|6|10|et circumspectis omnibus dixit homini extende manum tuam et extendit et restituta est manus eius
LUKE|6|11|ipsi autem repleti sunt insipientia et conloquebantur ad invicem quidnam facerent Iesu
LUKE|6|12|factum est autem in illis diebus exiit in montem orare et erat pernoctans in oratione Dei
LUKE|6|13|et cum dies factus esset vocavit discipulos suos et elegit duodecim ex ipsis quos et apostolos nominavit
LUKE|6|14|Simonem quem cognominavit Petrum et Andream fratrem eius Iacobum et Iohannem Philippum et Bartholomeum
LUKE|6|15|Mattheum et Thomam Iacobum Alphei et Simonem qui vocatur Zelotes
LUKE|6|16|Iudam Iacobi et Iudam Scarioth qui fuit proditor
LUKE|6|17|et descendens cum illis stetit in loco campestri et turba discipulorum eius et multitudo copiosa plebis ab omni Iudaea et Hierusalem et maritimae Tyri et Sidonis
LUKE|6|18|qui venerunt ut audirent eum et sanarentur a languoribus suis et qui vexabantur ab spiritibus inmundis curabantur
LUKE|6|19|et omnis turba quaerebant eum tangere quia virtus de illo exiebat et sanabat omnes
LUKE|6|20|et ipse elevatis oculis in discipulos suos dicebat beati pauperes quia vestrum est regnum Dei
LUKE|6|21|beati qui nunc esuritis quia saturabimini beati qui nunc fletis quia ridebitis
LUKE|6|22|beati eritis cum vos oderint homines et cum separaverint vos et exprobraverint et eiecerint nomen vestrum tamquam malum propter Filium hominis
LUKE|6|23|gaudete in illa die et exultate ecce enim merces vestra multa in caelo secundum haec enim faciebant prophetis patres eorum
LUKE|6|24|verumtamen vae vobis divitibus quia habetis consolationem vestram
LUKE|6|25|vae vobis qui saturati estis quia esurietis vae vobis qui ridetis nunc quia lugebitis et flebitis
LUKE|6|26|vae cum bene vobis dixerint omnes homines secundum haec faciebant prophetis patres eorum
LUKE|6|27|sed vobis dico qui auditis diligite inimicos vestros benefacite his qui vos oderunt
LUKE|6|28|benedicite maledicentibus vobis orate pro calumniantibus vos
LUKE|6|29|ei qui te percutit in maxillam praebe et alteram et ab eo qui aufert tibi vestimentum etiam tunicam noli prohibere
LUKE|6|30|omni autem petenti te tribue et qui aufert quae tua sunt ne repetas
LUKE|6|31|et prout vultis ut faciant vobis homines et vos facite illis similiter
LUKE|6|32|et si diligitis eos qui vos diligunt quae vobis est gratia nam et peccatores diligentes se diligunt
LUKE|6|33|et si benefeceritis his qui vobis benefaciunt quae vobis est gratia siquidem et peccatores hoc faciunt
LUKE|6|34|et si mutuum dederitis his a quibus speratis recipere quae gratia est vobis nam et peccatores peccatoribus fenerantur ut recipiant aequalia
LUKE|6|35|verumtamen diligite inimicos vestros et benefacite et mutuum date nihil desperantes et erit merces vestra multa et eritis filii Altissimi quia ipse benignus est super ingratos et malos
LUKE|6|36|estote ergo misericordes sicut et Pater vester misericors est
LUKE|6|37|nolite iudicare et non iudicabimini nolite condemnare et non condemnabimini dimittite et dimittemini
LUKE|6|38|date et dabitur vobis mensuram bonam confersam et coagitatam et supereffluentem dabunt in sinum vestrum eadem quippe mensura qua mensi fueritis remetietur vobis
LUKE|6|39|dicebat autem illis et similitudinem numquid potest caecus caecum ducere nonne ambo in foveam cadent
LUKE|6|40|non est discipulus super magistrum perfectus autem omnis erit sicut magister eius
LUKE|6|41|quid autem vides festucam in oculo fratris tui trabem autem quae in oculo tuo est non consideras
LUKE|6|42|et quomodo potes dicere fratri tuo frater sine eiciam festucam de oculo tuo ipse in oculo tuo trabem non videns hypocrita eice primum trabem de oculo tuo et tunc perspicies ut educas festucam de oculo fratris tui
LUKE|6|43|non est enim arbor bona quae facit fructus malos neque arbor mala faciens fructum bonum
LUKE|6|44|unaquaeque enim arbor de fructu suo cognoscitur neque enim de spinis colligunt ficus neque de rubo vindemiant uvam
LUKE|6|45|bonus homo de bono thesauro cordis sui profert bonum et malus homo de malo profert malum ex abundantia enim cordis os loquitur
LUKE|6|46|quid autem vocatis me Domine Domine et non facitis quae dico
LUKE|6|47|omnis qui venit ad me et audit sermones meos et facit eos ostendam vobis cui similis est
LUKE|6|48|similis est homini aedificanti domum qui fodit in altum et posuit fundamenta supra petram inundatione autem facta inlisum est flumen domui illi et non potuit eam movere fundata enim erat supra petram
LUKE|6|49|qui autem audivit et non fecit similis est homini aedificanti domum suam supra terram sine fundamento in quam inlisus est fluvius et continuo concidit et facta est ruina domus illius magna
LUKE|7|1|cum autem implesset omnia verba sua in aures plebis intravit Capharnaum
LUKE|7|2|centurionis autem cuiusdam servus male habens erat moriturus qui illi erat pretiosus
LUKE|7|3|et cum audisset de Iesu misit ad eum seniores Iudaeorum rogans eum ut veniret et salvaret servum eius
LUKE|7|4|at illi cum venissent ad Iesum rogabant eum sollicite dicentes ei quia dignus est ut hoc illi praestes
LUKE|7|5|diligit enim gentem nostram et synagogam ipse aedificavit nobis
LUKE|7|6|Iesus autem ibat cum illis et cum iam non longe esset a domo misit ad eum centurio amicos dicens Domine noli vexari non enim dignus sum ut sub tectum meum intres
LUKE|7|7|propter quod et me ipsum non sum dignum arbitratus ut venirem ad te sed dic verbo et sanabitur puer meus
LUKE|7|8|nam et ego homo sum sub potestate constitutus habens sub me milites et dico huic vade et vadit et alio veni et venit et servo meo fac hoc et facit
LUKE|7|9|quo audito Iesus miratus est et conversus sequentibus se turbis dixit amen dico vobis nec in Israhel tantam fidem inveni
LUKE|7|10|et reversi qui missi fuerant domum invenerunt servum qui languerat sanum
LUKE|7|11|et factum est deinceps ibat in civitatem quae vocatur Naim et ibant cum illo discipuli eius et turba copiosa
LUKE|7|12|cum autem adpropinquaret portae civitatis et ecce defunctus efferebatur filius unicus matri suae et haec vidua erat et turba civitatis multa cum illa
LUKE|7|13|quam cum vidisset Dominus misericordia motus super ea dixit illi noli flere
LUKE|7|14|et accessit et tetigit loculum hii autem qui portabant steterunt et ait adulescens tibi dico surge
LUKE|7|15|et resedit qui erat mortuus et coepit loqui et dedit illum matri suae
LUKE|7|16|accepit autem omnes timor et magnificabant Deum dicentes quia propheta magnus surrexit in nobis et quia Deus visitavit plebem suam
LUKE|7|17|et exiit hic sermo in universam Iudaeam de eo et omnem circa regionem
LUKE|7|18|et nuntiaverunt Iohanni discipuli eius de omnibus his
LUKE|7|19|et convocavit duos de discipulis suis Iohannes et misit ad Dominum dicens tu es qui venturus es an alium expectamus
LUKE|7|20|cum autem venissent ad eum viri dixerunt Iohannes Baptista misit nos ad te dicens tu es qui venturus es an alium expectamus
LUKE|7|21|in ipsa autem hora curavit multos a languoribus et plagis et spiritibus malis et caecis multis donavit visum
LUKE|7|22|et respondens dixit illis euntes nuntiate Iohanni quae vidistis et audistis quia caeci vident claudi ambulant leprosi mundantur surdi audiunt mortui resurgunt pauperes evangelizantur
LUKE|7|23|et beatus est quicumque non fuerit scandalizatus in me
LUKE|7|24|et cum discessissent nuntii Iohannis coepit dicere de Iohanne ad turbas quid existis in desertum videre harundinem vento moveri
LUKE|7|25|sed quid existis videre hominem mollibus vestimentis indutum ecce qui in veste pretiosa sunt et deliciis in domibus regum sunt
LUKE|7|26|sed quid existis videre prophetam utique dico vobis et plus quam prophetam
LUKE|7|27|hic est de quo scriptum est ecce mitto angelum meum ante faciem tuam qui praeparabit viam tuam ante te
LUKE|7|28|dico enim vobis maior inter natos mulierum propheta Iohanne Baptista nemo est qui autem minor est in regno Dei maior est illo
LUKE|7|29|et omnis populus audiens et publicani iustificaverunt Deum baptizati baptismo Iohannis
LUKE|7|30|Pharisaei autem et legis periti consilium Dei spreverunt in semet ipsos non baptizati ab eo
LUKE|7|31|cui ergo similes dicam homines generationis huius et cui similes sunt
LUKE|7|32|similes sunt pueris sedentibus in foro et loquentibus ad invicem et dicentibus cantavimus vobis tibiis et non saltastis lamentavimus et non plorastis
LUKE|7|33|venit enim Iohannes Baptista neque manducans panem neque bibens vinum et dicitis daemonium habet
LUKE|7|34|venit Filius hominis manducans et bibens et dicitis ecce homo devorator et bibens vinum amicus publicanorum et peccatorum
LUKE|7|35|et iustificata est sapientia ab omnibus filiis suis
LUKE|7|36|rogabat autem illum quidam de Pharisaeis ut manducaret cum illo et ingressus domum Pharisaei discubuit
LUKE|7|37|et ecce mulier quae erat in civitate peccatrix ut cognovit quod accubuit in domo Pharisaei adtulit alabastrum unguenti
LUKE|7|38|et stans retro secus pedes eius lacrimis coepit rigare pedes eius et capillis capitis sui tergebat et osculabatur pedes eius et unguento unguebat
LUKE|7|39|videns autem Pharisaeus qui vocaverat eum ait intra se dicens hic si esset propheta sciret utique quae et qualis mulier quae tangit eum quia peccatrix est
LUKE|7|40|et respondens Iesus dixit ad illum Simon habeo tibi aliquid dicere at ille ait magister dic
LUKE|7|41|duo debitores erant cuidam feneratori unus debebat denarios quingentos alius quinquaginta
LUKE|7|42|non habentibus illis unde redderent donavit utrisque quis ergo eum plus diliget
LUKE|7|43|respondens Simon dixit aestimo quia is cui plus donavit at ille dixit ei recte iudicasti
LUKE|7|44|et conversus ad mulierem dixit Simoni vides hanc mulierem intravi in domum tuam aquam pedibus meis non dedisti haec autem lacrimis rigavit pedes meos et capillis suis tersit
LUKE|7|45|osculum mihi non dedisti haec autem ex quo intravit non cessavit osculari pedes meos
LUKE|7|46|oleo caput meum non unxisti haec autem unguento unxit pedes meos
LUKE|7|47|propter quod dico tibi remittentur ei peccata multa quoniam dilexit multum cui autem minus dimittitur minus diligit
LUKE|7|48|dixit autem ad illam remittuntur tibi peccata
LUKE|7|49|et coeperunt qui simul accumbebant dicere intra se quis est hic qui etiam peccata dimittit
LUKE|7|50|dixit autem ad mulierem fides tua te salvam fecit vade in pace
LUKE|8|1|et factum est deinceps et ipse iter faciebat per civitatem et castellum praedicans et evangelizans regnum Dei et duodecim cum illo
LUKE|8|2|et mulieres aliquae quae erant curatae ab spiritibus malignis et infirmitatibus Maria quae vocatur Magdalene de qua daemonia septem exierant
LUKE|8|3|et Iohanna uxor Chuza procuratoris Herodis et Susanna et aliae multae quae ministrabant eis de facultatibus suis
LUKE|8|4|cum autem turba plurima conveniret et de civitatibus properarent ad eum dixit per similitudinem
LUKE|8|5|exiit qui seminat seminare semen suum et dum seminat aliud cecidit secus viam et conculcatum est et volucres caeli comederunt illud
LUKE|8|6|et aliud cecidit supra petram et natum aruit quia non habebat humorem
LUKE|8|7|et aliud cecidit inter spinas et simul exortae spinae suffocaverunt illud
LUKE|8|8|et aliud cecidit in terram bonam et ortum fecit fructum centuplum haec dicens clamabat qui habet aures audiendi audiat
LUKE|8|9|interrogabant autem eum discipuli eius quae esset haec parabola
LUKE|8|10|quibus ipse dixit vobis datum est nosse mysterium regni Dei ceteris autem in parabolis ut videntes non videant et audientes non intellegant
LUKE|8|11|est autem haec parabola semen est verbum Dei
LUKE|8|12|qui autem secus viam sunt qui audiunt deinde venit diabolus et tollit verbum de corde eorum ne credentes salvi fiant
LUKE|8|13|nam qui supra petram qui cum audierint cum gaudio suscipiunt verbum et hii radices non habent qui ad tempus credunt et in tempore temptationis recedunt
LUKE|8|14|quod autem in spinis cecidit hii sunt qui audierunt et a sollicitudinibus et divitiis et voluptatibus vitae euntes suffocantur et non referunt fructum
LUKE|8|15|quod autem in bonam terram hii sunt qui in corde bono et optimo audientes verbum retinent et fructum adferunt in patientia
LUKE|8|16|nemo autem lucernam accendens operit eam vaso aut subtus lectum ponit sed supra candelabrum ponit ut intrantes videant lumen
LUKE|8|17|non enim est occultum quod non manifestetur nec absconditum quod non cognoscatur et in palam veniat
LUKE|8|18|videte ergo quomodo auditis qui enim habet dabitur illi et quicumque non habet etiam quod putat se habere auferetur ab illo
LUKE|8|19|venerunt autem ad illum mater et fratres eius et non poterant adire ad eum prae turba
LUKE|8|20|et nuntiatum est illi mater tua et fratres tui stant foris volentes te videre
LUKE|8|21|qui respondens dixit ad eos mater mea et fratres mei hii sunt qui verbum Dei audiunt et faciunt
LUKE|8|22|factum est autem in una dierum et ipse ascendit in naviculam et discipuli eius et ait ad illos transfretemus trans stagnum et ascenderunt
LUKE|8|23|navigantibus autem illis obdormiit et descendit procella venti in stagnum et conplebantur et periclitabantur
LUKE|8|24|accedentes autem suscitaverunt eum dicentes praeceptor perimus at ille surgens increpavit ventum et tempestatem aquae et cessavit et facta est tranquillitas
LUKE|8|25|dixit autem illis ubi est fides vestra qui timentes mirati sunt dicentes ad invicem quis putas hic est quia et ventis imperat et mari et oboediunt ei
LUKE|8|26|enavigaverunt autem ad regionem Gerasenorum quae est contra Galilaeam
LUKE|8|27|et cum egressus esset ad terram occurrit illi vir quidam qui habebat daemonium iam temporibus multis et vestimento non induebatur neque in domo manebat sed in monumentis
LUKE|8|28|is ut vidit Iesum procidit ante illum et exclamans voce magna dixit quid mihi et tibi est Iesu Fili Dei altissimi obsecro te ne me torqueas
LUKE|8|29|praecipiebat enim spiritui inmundo ut exiret ab homine multis enim temporibus arripiebat illum et vinciebatur catenis et conpedibus custoditus et ruptis vinculis agebatur a daemonio in deserta
LUKE|8|30|interrogavit autem illum Iesus dicens quod tibi nomen est at ille dixit Legio quia intraverunt daemonia multa in eum
LUKE|8|31|et rogabant illum ne imperaret illis ut in abyssum irent
LUKE|8|32|erat autem ibi grex porcorum multorum pascentium in monte et rogabant eum ut permitteret eos in illos ingredi et permisit illos
LUKE|8|33|exierunt ergo daemonia ab homine et intraverunt in porcos et impetu abiit grex per praeceps in stagnum et suffocatus est
LUKE|8|34|quod ut viderunt factum qui pascebant fugerunt et nuntiaverunt in civitatem et in villas
LUKE|8|35|exierunt autem videre quod factum est et venerunt ad Iesum et invenerunt hominem sedentem a quo daemonia exierant vestitum ac sana mente ad pedes eius et timuerunt
LUKE|8|36|nuntiaverunt autem illis et qui viderant quomodo sanus factus esset a Legione
LUKE|8|37|et rogaverunt illum omnis multitudo regionis Gerasenorum ut discederet ab ipsis quia timore magno tenebantur ipse autem ascendens navem reversus est
LUKE|8|38|et rogabat illum vir a quo daemonia exierant ut cum eo esset dimisit autem eum Iesus dicens
LUKE|8|39|redi domum tuam et narra quanta tibi fecit Deus et abiit per universam civitatem praedicans quanta illi fecisset Iesus
LUKE|8|40|factum est autem cum redisset Iesus excepit illum turba erant enim omnes expectantes eum
LUKE|8|41|et ecce venit vir cui nomen Iairus et ipse princeps synagogae erat et cecidit ad pedes Iesu rogans eum ut intraret in domum eius
LUKE|8|42|quia filia unica erat illi fere annorum duodecim et haec moriebatur et contigit dum iret a turbis conprimebatur
LUKE|8|43|et mulier quaedam erat in fluxu sanguinis ab annis duodecim quae in medicos erogaverat omnem substantiam suam nec ab ullo potuit curari
LUKE|8|44|accessit retro et tetigit fimbriam vestimenti eius et confestim stetit fluxus sanguinis eius
LUKE|8|45|et ait Iesus quis est qui me tetigit negantibus autem omnibus dixit Petrus et qui cum illo erant praeceptor turbae te conprimunt et adfligunt et dicis quis me tetigit
LUKE|8|46|et dixit Iesus tetigit me aliquis nam ego novi virtutem de me exisse
LUKE|8|47|videns autem mulier quia non latuit tremens venit et procidit ante pedes illius et ob quam causam tetigerit eum indicavit coram omni populo et quemadmodum confestim sanata sit
LUKE|8|48|at ipse dixit illi filia fides tua te salvam fecit vade in pace
LUKE|8|49|adhuc illo loquente venit a principe synagogae dicens ei quia mortua est filia tua noli vexare illum
LUKE|8|50|Iesus autem audito hoc verbo respondit patri puellae noli timere crede tantum et salva erit
LUKE|8|51|et cum venisset domum non permisit intrare secum quemquam nisi Petrum et Iohannem et Iacobum et patrem et matrem puellae
LUKE|8|52|flebant autem omnes et plangebant illam at ille dixit nolite flere non est mortua sed dormit
LUKE|8|53|et deridebant eum scientes quia mortua esset
LUKE|8|54|ipse autem tenens manum eius clamavit dicens puella surge
LUKE|8|55|et reversus est spiritus eius et surrexit continuo et iussit illi dari manducare
LUKE|8|56|et stupuerunt parentes eius quibus praecepit ne alicui dicerent quod factum erat
LUKE|9|1|convocatis autem duodecim apostolis dedit illis virtutem et potestatem super omnia daemonia et ut languores curarent
LUKE|9|2|et misit illos praedicare regnum Dei et sanare infirmos
LUKE|9|3|et ait ad illos nihil tuleritis in via neque virgam neque peram neque panem neque pecuniam neque duas tunicas habeatis
LUKE|9|4|et in quamcumque domum intraveritis ibi manete et inde ne exeatis
LUKE|9|5|et quicumque non receperint vos exeuntes de civitate illa etiam pulverem pedum vestrorum excutite in testimonium supra illos
LUKE|9|6|egressi autem circumibant per castella evangelizantes et curantes ubique
LUKE|9|7|audivit autem Herodes tetrarcha omnia quae fiebant ab eo et haesitabat eo quod diceretur
LUKE|9|8|a quibusdam quia Iohannes surrexit a mortuis a quibusdam vero quia Helias apparuit ab aliis autem quia propheta unus de antiquis surrexit
LUKE|9|9|et ait Herodes Iohannem ego decollavi quis autem est iste de quo audio ego talia et quaerebat videre eum
LUKE|9|10|et reversi apostoli narraverunt illi quaecumque fecerunt et adsumptis illis secessit seorsum in locum desertum qui est Bethsaida
LUKE|9|11|quod cum cognovissent turbae secutae sunt illum et excepit illos et loquebatur illis de regno Dei et eos qui cura indigebant sanabat
LUKE|9|12|dies autem coeperat declinare et accedentes duodecim dixerunt illi dimitte turbas ut euntes in castella villasque quae circa sunt devertant et inveniant escas quia hic in loco deserto sumus
LUKE|9|13|ait autem ad illos vos date illis manducare at illi dixerunt non sunt nobis plus quam quinque panes et duo pisces nisi forte nos eamus et emamus in omnem hanc turbam escas
LUKE|9|14|erant autem fere viri quinque milia ait autem ad discipulos suos facite illos discumbere per convivia quinquagenos
LUKE|9|15|et ita fecerunt et discumbere fecerunt omnes
LUKE|9|16|acceptis autem quinque panibus et duobus piscibus respexit in caelum et benedixit illis et fregit et distribuit discipulis suis ut ponerent ante turbas
LUKE|9|17|et manducaverunt omnes et saturati sunt et sublatum est quod superfuit illis fragmentorum cofini duodecim
LUKE|9|18|et factum est cum solus esset orans erant cum illo et discipuli et interrogavit illos dicens quem me dicunt esse turbae
LUKE|9|19|at illi responderunt et dixerunt Iohannem Baptistam alii autem Heliam alii quia propheta unus de prioribus surrexit
LUKE|9|20|dixit autem illis vos autem quem me esse dicitis respondens Simon Petrus dixit Christum Dei
LUKE|9|21|at ille increpans illos praecepit ne cui dicerent hoc
LUKE|9|22|dicens quia oportet Filium hominis multa pati et reprobari a senioribus et principibus sacerdotum et scribis et occidi et tertia die resurgere
LUKE|9|23|dicebat autem ad omnes si quis vult post me venire abneget se ipsum et tollat crucem suam cotidie et sequatur me
LUKE|9|24|qui enim voluerit animam suam salvam facere perdet illam nam qui perdiderit animam suam propter me salvam faciet illam
LUKE|9|25|quid enim proficit homo si lucretur universum mundum se autem ipsum perdat et detrimentum sui faciat
LUKE|9|26|nam qui me erubuerit et meos sermones hunc Filius hominis erubescet cum venerit in maiestate sua et Patris et sanctorum angelorum
LUKE|9|27|dico autem vobis vere sunt aliqui hic stantes qui non gustabunt mortem donec videant regnum Dei
LUKE|9|28|factum est autem post haec verba fere dies octo et adsumpsit Petrum et Iohannem et Iacobum et ascendit in montem ut oraret
LUKE|9|29|et factum est dum oraret species vultus eius altera et vestitus eius albus refulgens
LUKE|9|30|et ecce duo viri loquebantur cum illo erant autem Moses et Helias
LUKE|9|31|visi in maiestate et dicebant excessum eius quem conpleturus erat in Hierusalem
LUKE|9|32|Petrus vero et qui cum illo gravati erant somno et evigilantes viderunt maiestatem eius et duos viros qui stabant cum illo
LUKE|9|33|et factum est cum discederent ab illo ait Petrus ad Iesum praeceptor bonum est nos hic esse et faciamus tria tabernacula unum tibi et unum Mosi et unum Heliae nesciens quid diceret
LUKE|9|34|haec autem illo loquente facta est nubes et obumbravit eos et timuerunt intrantibus illis in nubem
LUKE|9|35|et vox facta est de nube dicens hic est Filius meus electus ipsum audite
LUKE|9|36|et dum fieret vox inventus est Iesus solus et ipsi tacuerunt et nemini dixerunt in illis diebus quicquam ex his quae viderant
LUKE|9|37|factum est autem in sequenti die descendentibus illis de monte occurrit illi turba multa
LUKE|9|38|et ecce vir de turba exclamavit dicens magister obsecro te respice in filium meum quia unicus est mihi
LUKE|9|39|et ecce spiritus adprehendit illum et subito clamat et elidit et dissipat eum cum spuma et vix discedit dilanians eum
LUKE|9|40|et rogavi discipulos tuos ut eicerent illum et non potuerunt
LUKE|9|41|respondens autem Iesus dixit o generatio infidelis et perversa usquequo ero apud vos et patiar vos adduc huc filium tuum
LUKE|9|42|et cum accederet elisit illum daemonium et dissipavit
LUKE|9|43|et increpavit Iesus spiritum inmundum et sanavit puerum et reddidit illum patri eius
LUKE|9|44|stupebant autem omnes in magnitudine Dei omnibusque mirantibus in omnibus quae faciebat dixit ad discipulos suos ponite vos in cordibus vestris sermones istos Filius enim hominis futurum est ut tradatur in manus hominum
LUKE|9|45|at illi ignorabant verbum istud et erat velatum ante eos ut non sentirent illud et timebant interrogare eum de hoc verbo
LUKE|9|46|intravit autem cogitatio in eos quis eorum maior esset
LUKE|9|47|at Iesus videns cogitationes cordis illorum adprehendens puerum statuit eum secus se
LUKE|9|48|et ait illis quicumque susceperit puerum istum in nomine meo me recipit et quicumque me recipit recipit eum qui me misit nam qui minor est inter omnes vos hic maior est
LUKE|9|49|respondens autem Iohannes dixit praeceptor vidimus quendam in nomine tuo eicientem daemonia et prohibuimus eum quia non sequitur nobiscum
LUKE|9|50|et ait ad illum Iesus nolite prohibere qui enim non est adversum vos pro vobis est
LUKE|9|51|factum est autem dum conplerentur dies adsumptionis eius et ipse faciem suam firmavit ut iret Hierusalem
LUKE|9|52|et misit nuntios ante conspectum suum et euntes intraverunt in civitatem Samaritanorum ut pararent illi
LUKE|9|53|et non receperunt eum quia facies eius erat euntis Hierusalem
LUKE|9|54|cum vidissent autem discipuli eius Iacobus et Iohannes dixerunt Domine vis dicimus ut ignis descendat de caelo et consumat illos
LUKE|9|55|et conversus increpavit illos
LUKE|9|56|et abierunt in aliud castellum
LUKE|9|57|factum est autem ambulantibus illis in via dixit quidam ad illum sequar te quocumque ieris
LUKE|9|58|et ait illi Iesus vulpes foveas habent et volucres caeli nidos Filius autem hominis non habet ubi caput reclinet
LUKE|9|59|ait autem ad alterum sequere me ille autem dixit Domine permitte mihi primum ire sepelire patrem meum
LUKE|9|60|dixitque ei Iesus sine ut mortui sepeliant mortuos suos tu autem vade adnuntia regnum Dei
LUKE|9|61|et ait alter sequar te Domine sed primum permitte mihi renuntiare his qui domi sunt
LUKE|9|62|ait ad illum Iesus nemo mittens manum suam in aratrum et aspiciens retro aptus est regno Dei
LUKE|10|1|post haec autem designavit Dominus et alios septuaginta duos et misit illos binos ante faciem suam in omnem civitatem et locum quo erat ipse venturus
LUKE|10|2|et dicebat illis messis quidem multa operarii autem pauci rogate ergo Dominum messis ut mittat operarios in messem
LUKE|10|3|ite ecce ego mitto vos sicut agnos inter lupos
LUKE|10|4|nolite portare sacculum neque peram neque calciamenta et neminem per viam salutaveritis
LUKE|10|5|in quamcumque domum intraveritis primum dicite pax huic domui
LUKE|10|6|et si ibi fuerit filius pacis requiescet super illam pax vestra sin autem ad vos revertetur
LUKE|10|7|in eadem autem domo manete edentes et bibentes quae apud illos sunt dignus enim est operarius mercede sua nolite transire de domo in domum
LUKE|10|8|et in quamcumque civitatem intraveritis et susceperint vos manducate quae adponuntur vobis
LUKE|10|9|et curate infirmos qui in illa sunt et dicite illis adpropinquavit in vos regnum Dei
LUKE|10|10|in quamcumque civitatem intraveritis et non receperint vos exeuntes in plateas eius dicite
LUKE|10|11|etiam pulverem qui adhesit nobis de civitate vestra extergimus in vos tamen hoc scitote quia adpropinquavit regnum Dei
LUKE|10|12|dico vobis quia Sodomis in die illa remissius erit quam illi civitati
LUKE|10|13|vae tibi Corazain vae tibi Bethsaida quia si in Tyro et Sidone factae fuissent virtutes quae in vobis factae sunt olim in cilicio et cinere sedentes paeniterent
LUKE|10|14|verumtamen Tyro et Sidoni remissius erit in iudicio quam vobis
LUKE|10|15|et tu Capharnaum usque in caelum exaltata usque ad infernum demergeris
LUKE|10|16|qui vos audit me audit et qui vos spernit me spernit qui autem me spernit spernit eum qui me misit
LUKE|10|17|reversi sunt autem septuaginta duo cum gaudio dicentes Domine etiam daemonia subiciuntur nobis in nomine tuo
LUKE|10|18|et ait illis videbam Satanan sicut fulgur de caelo cadentem
LUKE|10|19|ecce dedi vobis potestatem calcandi supra serpentes et scorpiones et supra omnem virtutem inimici et nihil vobis nocebit
LUKE|10|20|verumtamen in hoc nolite gaudere quia spiritus vobis subiciuntur gaudete autem quod nomina vestra scripta sunt in caelis
LUKE|10|21|in ipsa hora exultavit Spiritu Sancto et dixit confiteor tibi Pater Domine caeli et terrae quod abscondisti haec a sapientibus et prudentibus et revelasti ea parvulis etiam Pater quia sic placuit ante te
LUKE|10|22|omnia mihi tradita sunt a Patre meo et nemo scit qui sit Filius nisi Pater et qui sit Pater nisi Filius et cui voluerit Filius revelare
LUKE|10|23|et conversus ad discipulos suos dixit beati oculi qui vident quae videtis
LUKE|10|24|dico enim vobis quod multi prophetae et reges voluerunt videre quae vos videtis et non viderunt et audire quae auditis et non audierunt
LUKE|10|25|et ecce quidam legis peritus surrexit temptans illum et dicens magister quid faciendo vitam aeternam possidebo
LUKE|10|26|at ille dixit ad eum in lege quid scriptum est quomodo legis
LUKE|10|27|ille respondens dixit diliges Dominum Deum tuum ex toto corde tuo et ex tota anima tua et ex omnibus viribus tuis et ex omni mente tua et proximum tuum sicut te ipsum
LUKE|10|28|dixitque illi recte respondisti hoc fac et vives
LUKE|10|29|ille autem volens iustificare se ipsum dixit ad Iesum et quis est meus proximus
LUKE|10|30|suscipiens autem Iesus dixit homo quidam descendebat ab Hierusalem in Hiericho et incidit in latrones qui etiam despoliaverunt eum et plagis inpositis abierunt semivivo relicto
LUKE|10|31|accidit autem ut sacerdos quidam descenderet eadem via et viso illo praeterivit
LUKE|10|32|similiter et Levita cum esset secus locum et videret eum pertransiit
LUKE|10|33|Samaritanus autem quidam iter faciens venit secus eum et videns eum misericordia motus est
LUKE|10|34|et adpropians alligavit vulnera eius infundens oleum et vinum et inponens illum in iumentum suum duxit in stabulum et curam eius egit
LUKE|10|35|et altera die protulit duos denarios et dedit stabulario et ait curam illius habe et quodcumque supererogaveris ego cum rediero reddam tibi
LUKE|10|36|quis horum trium videtur tibi proximus fuisse illi qui incidit in latrones
LUKE|10|37|at ille dixit qui fecit misericordiam in illum et ait illi Iesus vade et tu fac similiter
LUKE|10|38|factum est autem dum irent et ipse intravit in quoddam castellum et mulier quaedam Martha nomine excepit illum in domum suam
LUKE|10|39|et huic erat soror nomine Maria quae etiam sedens secus pedes Domini audiebat verbum illius
LUKE|10|40|Martha autem satagebat circa frequens ministerium quae stetit et ait Domine non est tibi curae quod soror mea reliquit me solam ministrare dic ergo illi ut me adiuvet
LUKE|10|41|et respondens dixit illi Dominus Martha Martha sollicita es et turbaris erga plurima
LUKE|10|42|porro unum est necessarium Maria optimam partem elegit quae non auferetur ab ea
LUKE|11|1|et factum est cum esset in loco quodam orans ut cessavit dixit unus ex discipulis eius ad eum Domine doce nos orare sicut et Iohannes docuit discipulos suos
LUKE|11|2|et ait illis cum oratis dicite Pater sanctificetur nomen tuum adveniat regnum tuum
LUKE|11|3|panem nostrum cotidianum da nobis cotidie
LUKE|11|4|et dimitte nobis peccata nostra siquidem et ipsi dimittimus omni debenti nobis et ne nos inducas in temptationem
LUKE|11|5|et ait ad illos quis vestrum habebit amicum et ibit ad illum media nocte et dicit illi amice commoda mihi tres panes
LUKE|11|6|quoniam amicus meus venit de via ad me et non habeo quod ponam ante illum
LUKE|11|7|et ille de intus respondens dicat noli mihi molestus esse iam ostium clausum est et pueri mei mecum sunt in cubili non possum surgere et dare tibi
LUKE|11|8|dico vobis et si non dabit illi surgens eo quod amicus eius sit propter inprobitatem tamen eius surget et dabit illi quotquot habet necessarios
LUKE|11|9|et ego vobis dico petite et dabitur vobis quaerite et invenietis pulsate et aperietur vobis
LUKE|11|10|omnis enim qui petit accipit et qui quaerit invenit et pulsanti aperietur
LUKE|11|11|quis autem ex vobis patrem petet panem numquid lapidem dabit illi aut piscem numquid pro pisce serpentem dabit illi
LUKE|11|12|aut si petierit ovum numquid porriget illi scorpionem
LUKE|11|13|si ergo vos cum sitis mali nostis bona data dare filiis vestris quanto magis Pater vester de caelo dabit spiritum bonum petentibus se
LUKE|11|14|et erat eiciens daemonium et illud erat mutum et cum eiecisset daemonium locutus est mutus et admiratae sunt turbae
LUKE|11|15|quidam autem ex eis dixerunt in Beelzebub principe daemoniorum eicit daemonia
LUKE|11|16|et alii temptantes signum de caelo quaerebant ab eo
LUKE|11|17|ipse autem ut vidit cogitationes eorum dixit eis omne regnum in se ipsum divisum desolatur et domus supra domum cadet
LUKE|11|18|si autem et Satanas in se ipsum divisus est quomodo stabit regnum ipsius quia dicitis in Beelzebub eicere me daemonia
LUKE|11|19|si autem ego in Beelzebub eicio daemonia filii vestri in quo eiciunt ideo ipsi iudices vestri erunt
LUKE|11|20|porro si in digito Dei eicio daemonia profecto praevenit in vos regnum Dei
LUKE|11|21|cum fortis armatus custodit atrium suum in pace sunt ea quae possidet
LUKE|11|22|si autem fortior illo superveniens vicerit eum universa arma eius aufert in quibus confidebat et spolia eius distribuit
LUKE|11|23|qui non est mecum adversum me est et qui non colligit mecum dispergit
LUKE|11|24|cum inmundus spiritus exierit de homine perambulat per loca inaquosa quaerens requiem et non inveniens dicit revertar in domum meam unde exivi
LUKE|11|25|et cum venerit invenit scopis mundatam
LUKE|11|26|et tunc vadit et adsumit septem alios spiritus nequiores se et ingressi habitant ibi et sunt novissima hominis illius peiora prioribus
LUKE|11|27|factum est autem cum haec diceret extollens vocem quaedam mulier de turba dixit illi beatus venter qui te portavit et ubera quae suxisti
LUKE|11|28|at ille dixit quippini beati qui audiunt verbum Dei et custodiunt
LUKE|11|29|turbis autem concurrentibus coepit dicere generatio haec generatio nequam est signum quaerit et signum non dabitur illi nisi signum Ionae
LUKE|11|30|nam sicut Ionas fuit signum Ninevitis ita erit et Filius hominis generationi isti
LUKE|11|31|regina austri surget in iudicio cum viris generationis huius et condemnabit illos quia venit a finibus terrae audire sapientiam Salomonis et ecce plus Salomone hic
LUKE|11|32|viri ninevitae surgent in iudicio cum generatione hac et condemnabunt illam quia paenitentiam egerunt ad praedicationem Ionae et ecce plus Iona hic
LUKE|11|33|nemo lucernam accendit et in abscondito ponit neque sub modio sed supra candelabrum ut qui ingrediuntur lumen videant
LUKE|11|34|lucerna corporis tui est oculus tuus si oculus tuus fuerit simplex totum corpus tuum lucidum erit si autem nequam fuerit etiam corpus tuum tenebrosum erit
LUKE|11|35|vide ergo ne lumen quod in te est tenebrae sint
LUKE|11|36|si ergo corpus tuum totum lucidum fuerit non habens aliquam partem tenebrarum erit lucidum totum et sicut lucerna fulgoris inluminabit te
LUKE|11|37|et cum loqueretur rogavit illum quidam Pharisaeus ut pranderet apud se et ingressus recubuit
LUKE|11|38|Pharisaeus autem coepit intra se reputans dicere quare non baptizatus esset ante prandium
LUKE|11|39|et ait Dominus ad illum nunc vos Pharisaei quod de foris est calicis et catini mundatis quod autem intus est vestrum plenum est rapina et iniquitate
LUKE|11|40|stulti nonne qui fecit quod de foris est etiam id quod de intus est fecit
LUKE|11|41|verumtamen quod superest date elemosynam et ecce omnia munda sunt vobis
LUKE|11|42|sed vae vobis Pharisaeis quia decimatis mentam et rutam et omne holus et praeteritis iudicium et caritatem Dei haec autem oportuit facere et illa non omittere
LUKE|11|43|vae vobis Pharisaeis quia diligitis primas cathedras in synagogis et salutationes in foro
LUKE|11|44|vae vobis quia estis ut monumenta quae non parent et homines ambulantes supra nesciunt
LUKE|11|45|respondens autem quidam ex legis peritis ait illi magister haec dicens etiam nobis contumeliam facis
LUKE|11|46|at ille ait et vobis legis peritis vae quia oneratis homines oneribus quae portari non possunt et ipsi uno digito vestro non tangitis sarcinas
LUKE|11|47|vae vobis quia aedificatis monumenta prophetarum patres autem vestri occiderunt illos
LUKE|11|48|profecto testificamini quod consentitis operibus patrum vestrorum quoniam quidem ipsi eos occiderunt vos autem aedificatis eorum sepulchra
LUKE|11|49|propterea et sapientia Dei dixit mittam ad illos prophetas et apostolos et ex illis occident et persequentur
LUKE|11|50|ut inquiratur sanguis omnium prophetarum qui effusus est a constitutione mundi a generatione ista
LUKE|11|51|a sanguine Abel usque ad sanguinem Zacchariae qui periit inter altare et aedem ita dico vobis requiretur ab hac generatione
LUKE|11|52|vae vobis legis peritis quia tulistis clavem scientiae ipsi non introistis et eos qui introibant prohibuistis
LUKE|11|53|cum haec ad illos diceret coeperunt Pharisaei et legis periti graviter insistere et os eius opprimere de multis
LUKE|11|54|insidiantes et quaerentes capere aliquid ex ore eius ut accusarent eum
LUKE|12|1|multis autem turbis circumstantibus ita ut se invicem conculcarent coepit dicere ad discipulos suos adtendite a fermento Pharisaeorum quae est hypocrisis
LUKE|12|2|nihil autem opertum est quod non reveletur neque absconditum quod non sciatur
LUKE|12|3|quoniam quae in tenebris dixistis in lumine dicentur et quod in aurem locuti estis in cubiculis praedicabitur in tectis
LUKE|12|4|dico autem vobis amicis meis ne terreamini ab his qui occidunt corpus et post haec non habent amplius quod faciant
LUKE|12|5|ostendam autem vobis quem timeatis timete eum qui postquam occiderit habet potestatem mittere in gehennam ita dico vobis hunc timete
LUKE|12|6|nonne quinque passeres veneunt dipundio et unus ex illis non est in oblivione coram Deo
LUKE|12|7|sed et capilli capitis vestri omnes numerati sunt nolite ergo timere multis passeribus pluris estis
LUKE|12|8|dico autem vobis omnis quicumque confessus fuerit in me coram hominibus et Filius hominis confitebitur in illo coram angelis Dei
LUKE|12|9|qui autem negaverit me coram hominibus denegabitur coram angelis Dei
LUKE|12|10|et omnis qui dicit verbum in Filium hominis remittetur illi ei autem qui in Spiritum Sanctum blasphemaverit non remittetur
LUKE|12|11|cum autem inducent vos in synagogas et ad magistratus et potestates nolite solliciti esse qualiter aut quid respondeatis aut quid dicatis
LUKE|12|12|Spiritus enim Sanctus docebit vos in ipsa hora quae oporteat dicere
LUKE|12|13|ait autem quidam ei de turba magister dic fratri meo ut dividat mecum hereditatem
LUKE|12|14|at ille dixit ei homo quis me constituit iudicem aut divisorem super vos
LUKE|12|15|dixitque ad illos videte et cavete ab omni avaritia quia non in abundantia cuiusquam vita eius est ex his quae possidet
LUKE|12|16|dixit autem similitudinem ad illos dicens hominis cuiusdam divitis uberes fructus ager adtulit
LUKE|12|17|et cogitabat intra se dicens quid faciam quod non habeo quo congregem fructus meos
LUKE|12|18|et dixit hoc faciam destruam horrea mea et maiora faciam et illuc congregabo omnia quae nata sunt mihi et bona mea
LUKE|12|19|et dicam animae meae anima habes multa bona posita in annos plurimos requiesce comede bibe epulare
LUKE|12|20|dixit autem illi Deus stulte hac nocte animam tuam repetunt a te quae autem parasti cuius erunt
LUKE|12|21|sic est qui sibi thesaurizat et non est in Deum dives
LUKE|12|22|dixitque ad discipulos suos ideo dico vobis nolite solliciti esse animae quid manducetis neque corpori quid vestiamini
LUKE|12|23|anima plus est quam esca et corpus quam vestimentum
LUKE|12|24|considerate corvos quia non seminant neque metunt quibus non est cellarium neque horreum et Deus pascit illos quanto magis vos pluris estis illis
LUKE|12|25|quis autem vestrum cogitando potest adicere ad staturam suam cubitum unum
LUKE|12|26|si ergo neque quod minimum est potestis quid de ceteris solliciti estis
LUKE|12|27|considerate lilia quomodo crescunt non laborant non nent dico autem vobis nec Salomon in omni gloria sua vestiebatur sicut unum ex istis
LUKE|12|28|si autem faenum quod hodie in agro est et cras in clibanum mittitur Deus sic vestit quanto magis vos pusillae fidei
LUKE|12|29|et vos nolite quaerere quid manducetis aut quid bibatis et nolite in sublime tolli
LUKE|12|30|haec enim omnia gentes mundi quaerunt Pater autem vester scit quoniam his indigetis
LUKE|12|31|verumtamen quaerite regnum Dei et haec omnia adicientur vobis
LUKE|12|32|nolite timere pusillus grex quia conplacuit Patri vestro dare vobis regnum
LUKE|12|33|vendite quae possidetis et date elemosynam facite vobis sacculos qui non veterescunt thesaurum non deficientem in caelis quo fur non adpropiat neque tinea corrumpit
LUKE|12|34|ubi enim thesaurus vester est ibi et cor vestrum erit
LUKE|12|35|sint lumbi vestri praecincti et lucernae ardentes
LUKE|12|36|et vos similes hominibus expectantibus dominum suum quando revertatur a nuptiis ut cum venerit et pulsaverit confestim aperiant ei
LUKE|12|37|beati servi illi quos cum venerit dominus invenerit vigilantes amen dico vobis quod praecinget se et faciet illos discumbere et transiens ministrabit illis
LUKE|12|38|et si venerit in secunda vigilia et si in tertia vigilia venerit et ita invenerit beati sunt servi illi
LUKE|12|39|hoc autem scitote quia si sciret pater familias qua hora fur veniret vigilaret utique et non sineret perfodiri domum suam
LUKE|12|40|et vos estote parati quia qua hora non putatis Filius hominis venit
LUKE|12|41|ait autem ei Petrus Domine ad nos dicis hanc parabolam an et ad omnes
LUKE|12|42|dixit autem Dominus quis putas est fidelis dispensator et prudens quem constituet dominus super familiam suam ut det illis in tempore tritici mensuram
LUKE|12|43|beatus ille servus quem cum venerit dominus invenerit ita facientem
LUKE|12|44|vere dico vobis quia supra omnia quae possidet constituet illum
LUKE|12|45|quod si dixerit servus ille in corde suo moram facit dominus meus venire et coeperit percutere pueros et ancillas et edere et bibere et inebriari
LUKE|12|46|veniet dominus servi illius in die qua non sperat et hora qua nescit et dividet eum partemque eius cum infidelibus ponet
LUKE|12|47|ille autem servus qui cognovit voluntatem domini sui et non praeparavit et non fecit secundum voluntatem eius vapulabit multas
LUKE|12|48|qui autem non cognovit et fecit digna plagis vapulabit paucis omni autem cui multum datum est multum quaeretur ab eo et cui commendaverunt multum plus petent ab eo
LUKE|12|49|ignem veni mittere in terram et quid volo si accendatur
LUKE|12|50|baptisma autem habeo baptizari et quomodo coartor usque dum perficiatur
LUKE|12|51|putatis quia pacem veni dare in terram non dico vobis sed separationem
LUKE|12|52|erunt enim ex hoc quinque in domo una divisi tres in duo et duo in tres
LUKE|12|53|dividentur pater in filium et filius in patrem suum mater in filiam et filia in matrem socrus in nurum suam et nurus in socrum suam
LUKE|12|54|dicebat autem et ad turbas cum videritis nubem orientem ab occasu statim dicitis nimbus venit et ita fit
LUKE|12|55|et cum austrum flantem dicitis quia aestus erit et fit
LUKE|12|56|hypocritae faciem terrae et caeli nostis probare hoc autem tempus quomodo non probatis
LUKE|12|57|quid autem et a vobis ipsis non iudicatis quod iustum est
LUKE|12|58|cum autem vadis cum adversario tuo ad principem in via da operam liberari ab illo ne forte trahat te apud iudicem et iudex tradat te exactori et exactor mittat te in carcerem
LUKE|12|59|dico tibi non exies inde donec etiam novissimum minutum reddas
LUKE|13|1|aderant autem quidam ipso in tempore nuntiantes illi de Galilaeis quorum sanguinem Pilatus miscuit cum sacrificiis eorum
LUKE|13|2|et respondens dixit illis putatis quod hii Galilaei prae omnibus Galilaeis peccatores fuerunt quia talia passi sunt
LUKE|13|3|non dico vobis sed nisi paenitentiam habueritis omnes similiter peribitis
LUKE|13|4|sicut illi decem et octo supra quos cecidit turris in Siloam et occidit eos putatis quia et ipsi debitores fuerunt praeter omnes homines habitantes in Hierusalem
LUKE|13|5|non dico vobis sed si non paenitentiam egeritis omnes similiter peribitis
LUKE|13|6|dicebat autem hanc similitudinem arborem fici habebat quidam plantatam in vinea sua et venit quaerens fructum in illa et non invenit
LUKE|13|7|dixit autem ad cultorem vineae ecce anni tres sunt ex quo venio quaerens fructum in ficulnea hac et non invenio succide ergo illam ut quid etiam terram occupat
LUKE|13|8|at ille respondens dixit illi domine dimitte illam et hoc anno usque dum fodiam circa illam et mittam stercora
LUKE|13|9|et si quidem fecerit fructum sin autem in futurum succides eam
LUKE|13|10|erat autem docens in synagoga eorum sabbatis
LUKE|13|11|et ecce mulier quae habebat spiritum infirmitatis annis decem et octo et erat inclinata nec omnino poterat sursum respicere
LUKE|13|12|quam cum videret Iesus vocavit ad se et ait illi mulier dimissa es ab infirmitate tua
LUKE|13|13|et inposuit illi manus et confestim erecta est et glorificabat Deum
LUKE|13|14|respondens autem archisynagogus indignans quia sabbato curasset Iesus dicebat turbae sex dies sunt in quibus oportet operari in his ergo venite et curamini et non in die sabbati
LUKE|13|15|respondit autem ad illum Dominus et dixit hypocritae unusquisque vestrum sabbato non solvit bovem suum aut asinum a praesepio et ducit adaquare
LUKE|13|16|hanc autem filiam Abrahae quam alligavit Satanas ecce decem et octo annis non oportuit solvi a vinculo isto die sabbati
LUKE|13|17|et cum haec diceret erubescebant omnes adversarii eius et omnis populus gaudebat in universis quae gloriose fiebant ab eo
LUKE|13|18|dicebat ergo cui simile est regnum Dei et cui simile esse existimabo illud
LUKE|13|19|simile est grano sinapis quod acceptum homo misit in hortum suum et crevit et factum est in arborem magnam et volucres caeli requieverunt in ramis eius
LUKE|13|20|et iterum dixit cui simile aestimabo regnum Dei
LUKE|13|21|simile est fermento quod acceptum mulier abscondit in farinae sata tria donec fermentaretur totum
LUKE|13|22|et ibat per civitates et castella docens et iter faciens in Hierusalem
LUKE|13|23|ait autem illi quidam Domine si pauci sunt qui salvantur ipse autem dixit ad illos
LUKE|13|24|contendite intrare per angustam portam quia multi dico vobis quaerunt intrare et non poterunt
LUKE|13|25|cum autem intraverit pater familias et cluserit ostium et incipietis foris stare et pulsare ostium dicentes Domine aperi nobis et respondens dicet vobis nescio vos unde sitis
LUKE|13|26|tunc incipietis dicere manducavimus coram te et bibimus et in plateis nostris docuisti
LUKE|13|27|et dicet vobis nescio vos unde sitis discedite a me omnes operarii iniquitatis
LUKE|13|28|ibi erit fletus et stridor dentium cum videritis Abraham et Isaac et Iacob et omnes prophetas in regno Dei vos autem expelli foras
LUKE|13|29|et venient ab oriente et occidente et aquilone et austro et accumbent in regno Dei
LUKE|13|30|et ecce sunt novissimi qui erunt primi et sunt primi qui erunt novissimi
LUKE|13|31|in ipsa die accesserunt quidam Pharisaeorum dicentes illi exi et vade hinc quia Herodes vult te occidere
LUKE|13|32|et ait illis ite dicite vulpi illi ecce eicio daemonia et sanitates perficio hodie et cras et tertia consummor
LUKE|13|33|verumtamen oportet me hodie et cras et sequenti ambulare quia non capit prophetam perire extra Hierusalem
LUKE|13|34|Hierusalem Hierusalem quae occidis prophetas et lapidas eos qui mittuntur ad te quotiens volui congregare filios tuos quemadmodum avis nidum suum sub pinnis et noluisti
LUKE|13|35|ecce relinquitur vobis domus vestra dico autem vobis quia non videbitis me donec veniat cum dicetis benedictus qui venit in nomine Domini
LUKE|14|1|et factum est cum intraret in domum cuiusdam principis Pharisaeorum sabbato manducare panem et ipsi observabant eum
LUKE|14|2|et ecce homo quidam hydropicus erat ante illum
LUKE|14|3|et respondens Iesus dixit ad legis peritos et Pharisaeos dicens si licet sabbato curare
LUKE|14|4|at illi tacuerunt ipse vero adprehensum sanavit eum ac dimisit
LUKE|14|5|et respondens ad illos dixit cuius vestrum asinus aut bos in puteum cadet et non continuo extrahet illum die sabbati
LUKE|14|6|et non poterant ad haec respondere illi
LUKE|14|7|dicebat autem et ad invitatos parabolam intendens quomodo primos accubitus eligerent dicens ad illos
LUKE|14|8|cum invitatus fueris ad nuptias non discumbas in primo loco ne forte honoratior te sit invitatus ab eo
LUKE|14|9|et veniens is qui te et illum vocavit dicat tibi da huic locum et tunc incipias cum rubore novissimum locum tenere
LUKE|14|10|sed cum vocatus fueris vade recumbe in novissimo loco ut cum venerit qui te invitavit dicat tibi amice ascende superius tunc erit tibi gloria coram simul discumbentibus
LUKE|14|11|quia omnis qui se exaltat humiliabitur et qui se humiliat exaltabitur
LUKE|14|12|dicebat autem et ei qui se invitaverat cum facis prandium aut cenam noli vocare amicos tuos neque fratres tuos neque cognatos neque vicinos divites ne forte et ipsi te reinvitent et fiat tibi retributio
LUKE|14|13|sed cum facis convivium voca pauperes debiles claudos caecos
LUKE|14|14|et beatus eris quia non habent retribuere tibi retribuetur enim tibi in resurrectione iustorum
LUKE|14|15|haec cum audisset quidam de simul discumbentibus dixit illi beatus qui manducabit panem in regno Dei
LUKE|14|16|at ipse dixit ei homo quidam fecit cenam magnam et vocavit multos
LUKE|14|17|et misit servum suum hora cenae dicere invitatis ut venirent quia iam parata sunt omnia
LUKE|14|18|et coeperunt simul omnes excusare primus dixit ei villam emi et necesse habeo exire et videre illam rogo te habe me excusatum
LUKE|14|19|et alter dixit iuga boum emi quinque et eo probare illa rogo te habe me excusatum
LUKE|14|20|et alius dixit uxorem duxi et ideo non possum venire
LUKE|14|21|et reversus servus nuntiavit haec domino suo tunc iratus pater familias dixit servo suo exi cito in plateas et vicos civitatis et pauperes ac debiles et caecos et claudos introduc huc
LUKE|14|22|et ait servus domine factum est ut imperasti et adhuc locus est
LUKE|14|23|et ait dominus servo exi in vias et sepes et conpelle intrare ut impleatur domus mea
LUKE|14|24|dico autem vobis quod nemo virorum illorum qui vocati sunt gustabit cenam meam
LUKE|14|25|ibant autem turbae multae cum eo et conversus dixit ad illos
LUKE|14|26|si quis venit ad me et non odit patrem suum et matrem et uxorem et filios et fratres et sorores adhuc autem et animam suam non potest esse meus discipulus
LUKE|14|27|et qui non baiulat crucem suam et venit post me non potest esse meus discipulus
LUKE|14|28|quis enim ex vobis volens turrem aedificare non prius sedens conputat sumptus qui necessarii sunt si habet ad perficiendum
LUKE|14|29|ne posteaquam posuerit fundamentum et non potuerit perficere omnes qui vident incipiant inludere ei
LUKE|14|30|dicentes quia hic homo coepit aedificare et non potuit consummare
LUKE|14|31|aut qui rex iturus committere bellum adversus alium regem non sedens prius cogitat si possit cum decem milibus occurrere ei qui cum viginti milibus venit ad se
LUKE|14|32|alioquin adhuc illo longe agente legationem mittens rogat ea quae pacis sunt
LUKE|14|33|sic ergo omnis ex vobis qui non renuntiat omnibus quae possidet non potest meus esse discipulus
LUKE|14|34|bonum est sal si autem sal quoque evanuerit in quo condietur
LUKE|14|35|neque in terram neque in sterquilinium utile est sed foras mittetur qui habet aures audiendi audiat
LUKE|15|1|erant autem adpropinquantes ei publicani et peccatores ut audirent illum
LUKE|15|2|et murmurabant Pharisaei et scribae dicentes quia hic peccatores recipit et manducat cum illis
LUKE|15|3|et ait ad illos parabolam istam dicens
LUKE|15|4|quis ex vobis homo qui habet centum oves et si perdiderit unam ex illis nonne dimittit nonaginta novem in deserto et vadit ad illam quae perierat donec inveniat illam
LUKE|15|5|et cum invenerit eam inponit in umeros suos gaudens
LUKE|15|6|et veniens domum convocat amicos et vicinos dicens illis congratulamini mihi quia inveni ovem meam quae perierat
LUKE|15|7|dico vobis quod ita gaudium erit in caelo super uno peccatore paenitentiam habente quam super nonaginta novem iustis qui non indigent paenitentia
LUKE|15|8|aut quae mulier habens dragmas decem si perdiderit dragmam unam nonne accendit lucernam et everrit domum et quaerit diligenter donec inveniat
LUKE|15|9|et cum invenerit convocat amicas et vicinas dicens congratulamini mihi quia inveni dragmam quam perdideram
LUKE|15|10|ita dico vobis gaudium erit coram angelis Dei super uno peccatore paenitentiam agente
LUKE|15|11|ait autem homo quidam habuit duos filios
LUKE|15|12|et dixit adulescentior ex illis patri pater da mihi portionem substantiae quae me contingit et divisit illis substantiam
LUKE|15|13|et non post multos dies congregatis omnibus adulescentior filius peregre profectus est in regionem longinquam et ibi dissipavit substantiam suam vivendo luxuriose
LUKE|15|14|et postquam omnia consummasset facta est fames valida in regione illa et ipse coepit egere
LUKE|15|15|et abiit et adhesit uni civium regionis illius et misit illum in villam suam ut pasceret porcos
LUKE|15|16|et cupiebat implere ventrem suum de siliquis quas porci manducabant et nemo illi dabat
LUKE|15|17|in se autem reversus dixit quanti mercennarii patris mei abundant panibus ego autem hic fame pereo
LUKE|15|18|surgam et ibo ad patrem meum et dicam illi pater peccavi in caelum et coram te
LUKE|15|19|et iam non sum dignus vocari filius tuus fac me sicut unum de mercennariis tuis
LUKE|15|20|et surgens venit ad patrem suum cum autem adhuc longe esset vidit illum pater ipsius et misericordia motus est et adcurrens cecidit supra collum eius et osculatus est illum
LUKE|15|21|dixitque ei filius pater peccavi in caelum et coram te iam non sum dignus vocari filius tuus
LUKE|15|22|dixit autem pater ad servos suos cito proferte stolam primam et induite illum et date anulum in manum eius et calciamenta in pedes
LUKE|15|23|et adducite vitulum saginatum et occidite et manducemus et epulemur
LUKE|15|24|quia hic filius meus mortuus erat et revixit perierat et inventus est et coeperunt epulari
LUKE|15|25|erat autem filius eius senior in agro et cum veniret et adpropinquaret domui audivit symphoniam et chorum
LUKE|15|26|et vocavit unum de servis et interrogavit quae haec essent
LUKE|15|27|isque dixit illi frater tuus venit et occidit pater tuus vitulum saginatum quia salvum illum recepit
LUKE|15|28|indignatus est autem et nolebat introire pater ergo illius egressus coepit rogare illum
LUKE|15|29|at ille respondens dixit patri suo ecce tot annis servio tibi et numquam mandatum tuum praeterii et numquam dedisti mihi hedum ut cum amicis meis epularer
LUKE|15|30|sed postquam filius tuus hic qui devoravit substantiam suam cum meretricibus venit occidisti illi vitulum saginatum
LUKE|15|31|at ipse dixit illi fili tu semper mecum es et omnia mea tua sunt
LUKE|15|32|epulari autem et gaudere oportebat quia frater tuus hic mortuus erat et revixit perierat et inventus est
LUKE|16|1|dicebat autem et ad discipulos suos homo quidam erat dives qui habebat vilicum et hic diffamatus est apud illum quasi dissipasset bona ipsius
LUKE|16|2|et vocavit illum et ait illi quid hoc audio de te redde rationem vilicationis tuae iam enim non poteris vilicare
LUKE|16|3|ait autem vilicus intra se quid faciam quia dominus meus aufert a me vilicationem fodere non valeo mendicare erubesco
LUKE|16|4|scio quid faciam ut cum amotus fuero a vilicatione recipiant me in domos suas
LUKE|16|5|convocatis itaque singulis debitoribus domini sui dicebat primo quantum debes domino meo
LUKE|16|6|at ille dixit centum cados olei dixitque illi accipe cautionem tuam et sede cito scribe quinquaginta
LUKE|16|7|deinde alio dixit tu vero quantum debes qui ait centum choros tritici ait illi accipe litteras tuas et scribe octoginta
LUKE|16|8|et laudavit dominus vilicum iniquitatis quia prudenter fecisset quia filii huius saeculi prudentiores filiis lucis in generatione sua sunt
LUKE|16|9|et ego vobis dico facite vobis amicos de mamona iniquitatis ut cum defeceritis recipiant vos in aeterna tabernacula
LUKE|16|10|qui fidelis est in minimo et in maiori fidelis est et qui in modico iniquus est et in maiori iniquus est
LUKE|16|11|si ergo in iniquo mamona fideles non fuistis quod verum est quis credet vobis
LUKE|16|12|et si in alieno fideles non fuistis quod vestrum est quis dabit vobis
LUKE|16|13|nemo servus potest duobus dominis servire aut enim unum odiet et alterum diliget aut uni adherebit et alterum contemnet non potestis Deo servire et mamonae
LUKE|16|14|audiebant autem omnia haec Pharisaei qui erant avari et deridebant illum
LUKE|16|15|et ait illis vos estis qui iustificatis vos coram hominibus Deus autem novit corda vestra quia quod hominibus altum est abominatio est ante Deum
LUKE|16|16|lex et prophetae usque ad Iohannem ex eo regnum Dei evangelizatur et omnis in illud vim facit
LUKE|16|17|facilius est autem caelum et terram praeterire quam de lege unum apicem cadere
LUKE|16|18|omnis qui dimittit uxorem suam et ducit alteram moechatur et qui dimissam a viro ducit moechatur
LUKE|16|19|homo quidam erat dives et induebatur purpura et bysso et epulabatur cotidie splendide
LUKE|16|20|et erat quidam mendicus nomine Lazarus qui iacebat ad ianuam eius ulceribus plenus
LUKE|16|21|cupiens saturari de micis quae cadebant de mensa divitis sed et canes veniebant et lingebant ulcera eius
LUKE|16|22|factum est autem ut moreretur mendicus et portaretur ab angelis in sinum Abrahae mortuus est autem et dives et sepultus est in inferno
LUKE|16|23|elevans oculos suos cum esset in tormentis videbat Abraham a longe et Lazarum in sinu eius
LUKE|16|24|et ipse clamans dixit pater Abraham miserere mei et mitte Lazarum ut intinguat extremum digiti sui in aqua ut refrigeret linguam meam quia crucior in hac flamma
LUKE|16|25|et dixit illi Abraham fili recordare quia recepisti bona in vita tua et Lazarus similiter mala nunc autem hic consolatur tu vero cruciaris
LUKE|16|26|et in his omnibus inter nos et vos chasma magnum firmatum est ut hii qui volunt hinc transire ad vos non possint neque inde huc transmeare
LUKE|16|27|et ait rogo ergo te pater ut mittas eum in domum patris mei
LUKE|16|28|habeo enim quinque fratres ut testetur illis ne et ipsi veniant in locum hunc tormentorum
LUKE|16|29|et ait illi Abraham habent Mosen et prophetas audiant illos
LUKE|16|30|at ille dixit non pater Abraham sed si quis ex mortuis ierit ad eos paenitentiam agent
LUKE|16|31|ait autem illi si Mosen et prophetas non audiunt neque si quis ex mortuis resurrexerit credent
LUKE|17|1|et ad discipulos suos ait inpossibile est ut non veniant scandala vae autem illi per quem veniunt
LUKE|17|2|utilius est illi si lapis molaris inponatur circa collum eius et proiciatur in mare quam ut scandalizet unum de pusillis istis
LUKE|17|3|adtendite vobis si peccaverit frater tuus increpa illum et si paenitentiam egerit dimitte illi
LUKE|17|4|et si septies in die peccaverit in te et septies in die conversus fuerit ad te dicens paenitet me dimitte illi
LUKE|17|5|et dixerunt apostoli Domino adauge nobis fidem
LUKE|17|6|dixit autem Dominus si haberetis fidem sicut granum sinapis diceretis huic arbori moro eradicare et transplantare in mare et oboediret vobis
LUKE|17|7|quis autem vestrum habens servum arantem aut pascentem qui regresso de agro dicet illi statim transi recumbe
LUKE|17|8|et non dicet ei para quod cenem et praecinge te et ministra mihi donec manducem et bibam et post haec tu manducabis et bibes
LUKE|17|9|numquid gratiam habet servo illi quia fecit quae sibi imperaverat non puto
LUKE|17|10|sic et vos cum feceritis omnia quae praecepta sunt vobis dicite servi inutiles sumus quod debuimus facere fecimus
LUKE|17|11|et factum est dum iret in Hierusalem transiebat per mediam Samariam et Galilaeam
LUKE|17|12|et cum ingrederetur quoddam castellum occurrerunt ei decem viri leprosi qui steterunt a longe
LUKE|17|13|et levaverunt vocem dicentes Iesu praeceptor miserere nostri
LUKE|17|14|quos ut vidit dixit ite ostendite vos sacerdotibus et factum est dum irent mundati sunt
LUKE|17|15|unus autem ex illis ut vidit quia mundatus est regressus est cum magna voce magnificans Deum
LUKE|17|16|et cecidit in faciem ante pedes eius gratias agens et hic erat Samaritanus
LUKE|17|17|respondens autem Iesus dixit nonne decem mundati sunt et novem ubi sunt
LUKE|17|18|non est inventus qui rediret et daret gloriam Deo nisi hic alienigena
LUKE|17|19|et ait illi surge vade quia fides tua te salvum fecit
LUKE|17|20|interrogatus autem a Pharisaeis quando venit regnum Dei respondit eis et dixit non venit regnum Dei cum observatione
LUKE|17|21|neque dicent ecce hic aut ecce illic ecce enim regnum Dei intra vos est
LUKE|17|22|et ait ad discipulos venient dies quando desideretis videre unum diem Filii hominis et non videbitis
LUKE|17|23|et dicent vobis ecce hic ecce illic nolite ire neque sectemini
LUKE|17|24|nam sicut fulgur coruscans de sub caelo in ea quae sub caelo sunt fulget ita erit Filius hominis in die sua
LUKE|17|25|primum autem oportet illum multa pati et reprobari a generatione hac
LUKE|17|26|et sicut factum est in diebus Noe ita erit et in diebus Filii hominis
LUKE|17|27|edebant et bibebant uxores ducebant et dabantur ad nuptias usque in diem qua intravit Noe in arcam et venit diluvium et perdidit omnes
LUKE|17|28|similiter sicut factum est in diebus Loth edebant et bibebant emebant et vendebant plantabant aedificabant
LUKE|17|29|qua die autem exiit Loth a Sodomis pluit ignem et sulphur de caelo et omnes perdidit
LUKE|17|30|secundum haec erit qua die Filius hominis revelabitur
LUKE|17|31|in illa hora qui fuerit in tecto et vasa eius in domo ne descendat tollere illa et qui in agro similiter non redeat retro
LUKE|17|32|memores estote uxoris Loth
LUKE|17|33|quicumque quaesierit animam suam salvare perdet illam et qui perdiderit illam vivificabit eam
LUKE|17|34|dico vobis illa nocte erunt duo in lecto uno unus adsumetur et alter relinquetur
LUKE|17|35|duae erunt molentes in unum una adsumetur et altera relinquetur duo in agro unus adsumetur et alter relinquetur
LUKE|17|36|respondentes dicunt illi ubi Domine
LUKE|17|37|qui dixit eis ubicumque fuerit corpus illuc congregabuntur aquilae
LUKE|18|1|dicebat autem et parabolam ad illos quoniam oportet semper orare et non deficere
LUKE|18|2|dicens iudex quidam erat in quadam civitate qui Deum non timebat et hominem non verebatur
LUKE|18|3|vidua autem quaedam erat in civitate illa et veniebat ad eum dicens vindica me de adversario meo
LUKE|18|4|et nolebat per multum tempus post haec autem dixit intra se et si Deum non timeo nec hominem revereor
LUKE|18|5|tamen quia molesta est mihi haec vidua vindicabo illam ne in novissimo veniens suggillet me
LUKE|18|6|ait autem Dominus audite quid iudex iniquitatis dicit
LUKE|18|7|Deus autem non faciet vindictam electorum suorum clamantium ad se die ac nocte et patientiam habebit in illis
LUKE|18|8|dico vobis quia cito faciet vindictam illorum verumtamen Filius hominis veniens putas inveniet fidem in terra
LUKE|18|9|dixit autem et ad quosdam qui in se confidebant tamquam iusti et aspernabantur ceteros parabolam istam
LUKE|18|10|duo homines ascenderunt in templum ut orarent unus Pharisaeus et alter publicanus
LUKE|18|11|Pharisaeus stans haec apud se orabat Deus gratias ago tibi quia non sum sicut ceteri hominum raptores iniusti adulteri vel ut etiam hic publicanus
LUKE|18|12|ieiuno bis in sabbato decimas do omnium quae possideo
LUKE|18|13|et publicanus a longe stans nolebat nec oculos ad caelum levare sed percutiebat pectus suum dicens Deus propitius esto mihi peccatori
LUKE|18|14|dico vobis descendit hic iustificatus in domum suam ab illo quia omnis qui se exaltat humiliabitur et qui se humiliat exaltabitur
LUKE|18|15|adferebant autem ad illum et infantes ut eos tangeret quod cum viderent discipuli increpabant illos
LUKE|18|16|Iesus autem convocans illos dixit sinite pueros venire ad me et nolite eos vetare talium est enim regnum Dei
LUKE|18|17|amen dico vobis quicumque non acceperit regnum Dei sicut puer non intrabit in illud
LUKE|18|18|et interrogavit eum quidam princeps dicens magister bone quid faciens vitam aeternam possidebo
LUKE|18|19|dixit autem ei Iesus quid me dicis bonum nemo bonus nisi solus Deus
LUKE|18|20|mandata nosti non occides non moechaberis non furtum facies non falsum testimonium dices honora patrem tuum et matrem
LUKE|18|21|qui ait haec omnia custodivi a iuventute mea
LUKE|18|22|quo audito Iesus ait ei adhuc unum tibi deest omnia quaecumque habes vende et da pauperibus et habebis thesaurum in caelo et veni sequere me
LUKE|18|23|his ille auditis contristatus est quia dives erat valde
LUKE|18|24|videns autem illum Iesus tristem factum dixit quam difficile qui pecunias habent in regnum Dei intrabunt
LUKE|18|25|facilius est enim camelum per foramen acus transire quam divitem intrare in regnum Dei
LUKE|18|26|et dixerunt qui audiebant et quis potest salvus fieri
LUKE|18|27|ait illis quae inpossibilia sunt apud homines possibilia sunt apud Deum
LUKE|18|28|ait autem Petrus ecce nos dimisimus omnia et secuti sumus te
LUKE|18|29|qui dixit eis amen dico vobis nemo est qui reliquit domum aut parentes aut fratres aut uxorem aut filios propter regnum Dei
LUKE|18|30|et non recipiat multo plura in hoc tempore et in saeculo venturo vitam aeternam
LUKE|18|31|adsumpsit autem Iesus duodecim et ait illis ecce ascendimus Hierosolyma et consummabuntur omnia quae scripta sunt per prophetas de Filio hominis
LUKE|18|32|tradetur enim gentibus et inludetur et flagellabitur et conspuetur
LUKE|18|33|et postquam flagellaverint occident eum et die tertia resurget
LUKE|18|34|et ipsi nihil horum intellexerunt et erat verbum istud absconditum ab eis et non intellegebant quae dicebantur
LUKE|18|35|factum est autem cum adpropinquaret Hiericho caecus quidam sedebat secus viam mendicans
LUKE|18|36|et cum audiret turbam praetereuntem interrogabat quid hoc esset
LUKE|18|37|dixerunt autem ei quod Iesus Nazarenus transiret
LUKE|18|38|et clamavit dicens Iesu Fili David miserere mei
LUKE|18|39|et qui praeibant increpabant eum ut taceret ipse vero multo magis clamabat Fili David miserere mei
LUKE|18|40|stans autem Iesus iussit illum adduci ad se et cum adpropinquasset interrogavit illum
LUKE|18|41|dicens quid tibi vis faciam at ille dixit Domine ut videam
LUKE|18|42|et Iesus dixit illi respice fides tua te salvum fecit
LUKE|18|43|et confestim vidit et sequebatur illum magnificans Deum et omnis plebs ut vidit dedit laudem Deo
LUKE|19|1|et ingressus perambulabat Hiericho
LUKE|19|2|et ecce vir nomine Zaccheus et hic erat princeps publicanorum et ipse dives
LUKE|19|3|et quaerebat videre Iesum quis esset et non poterat prae turba quia statura pusillus erat
LUKE|19|4|et praecurrens ascendit in arborem sycomorum ut videret illum quia inde erat transiturus
LUKE|19|5|et cum venisset ad locum suspiciens Iesus vidit illum et dixit ad eum Zacchee festinans descende quia hodie in domo tua oportet me manere
LUKE|19|6|et festinans descendit et excepit illum gaudens
LUKE|19|7|et cum viderent omnes murmurabant dicentes quod ad hominem peccatorem devertisset
LUKE|19|8|stans autem Zaccheus dixit ad Dominum ecce dimidium bonorum meorum Domine do pauperibus et si quid aliquem defraudavi reddo quadruplum
LUKE|19|9|ait Iesus ad eum quia hodie salus domui huic facta est eo quod et ipse filius sit Abrahae
LUKE|19|10|venit enim Filius hominis quaerere et salvum facere quod perierat
LUKE|19|11|haec illis audientibus adiciens dixit parabolam eo quod esset prope Hierusalem et quia existimarent quod confestim regnum Dei manifestaretur
LUKE|19|12|dixit ergo homo quidam nobilis abiit in regionem longinquam accipere sibi regnum et reverti
LUKE|19|13|vocatis autem decem servis suis dedit illis decem mnas et ait ad illos negotiamini dum venio
LUKE|19|14|cives autem eius oderant illum et miserunt legationem post illum dicentes nolumus hunc regnare super nos
LUKE|19|15|et factum est ut rediret accepto regno et iussit vocari servos quibus dedit pecuniam ut sciret quantum quisque negotiatus esset
LUKE|19|16|venit autem primus dicens domine mna tua decem mnas adquisivit
LUKE|19|17|et ait illi euge bone serve quia in modico fidelis fuisti eris potestatem habens supra decem civitates
LUKE|19|18|et alter venit dicens domine mna tua fecit quinque mnas
LUKE|19|19|et huic ait et tu esto supra quinque civitates
LUKE|19|20|et alter venit dicens domine ecce mna tua quam habui repositam in sudario
LUKE|19|21|timui enim te quia homo austeris es tollis quod non posuisti et metis quod non seminasti
LUKE|19|22|dicit ei de ore tuo te iudico serve nequam sciebas quod ego austeris homo sum tollens quod non posui et metens quod non seminavi
LUKE|19|23|et quare non dedisti pecuniam meam ad mensam et ego veniens cum usuris utique exegissem illud
LUKE|19|24|et adstantibus dixit auferte ab illo mnam et date illi qui decem mnas habet
LUKE|19|25|et dixerunt ei domine habet decem mnas
LUKE|19|26|dico autem vobis quia omni habenti dabitur ab eo autem qui non habet et quod habet auferetur ab eo
LUKE|19|27|verumtamen inimicos meos illos qui noluerunt me regnare super se adducite huc et interficite ante me
LUKE|19|28|et his dictis praecedebat ascendens in Hierosolyma
LUKE|19|29|et factum est cum adpropinquasset ad Bethfage et Bethania ad montem qui vocatur Oliveti misit duos discipulos suos
LUKE|19|30|dicens ite in castellum quod contra est in quod introeuntes invenietis pullum asinae alligatum cui nemo umquam hominum sedit solvite illum et adducite
LUKE|19|31|et si quis vos interrogaverit quare solvitis sic dicetis ei quia Dominus operam eius desiderat
LUKE|19|32|abierunt autem qui missi erant et invenerunt sicut dixit illis stantem pullum
LUKE|19|33|solventibus autem illis pullum dixerunt domini eius ad illos quid solvitis pullum
LUKE|19|34|at illi dixerunt quia Dominus eum necessarium habet
LUKE|19|35|et duxerunt illum ad Iesum et iactantes vestimenta sua supra pullum inposuerunt Iesum
LUKE|19|36|eunte autem illo substernebant vestimenta sua in via
LUKE|19|37|et cum adpropinquaret iam ad descensum montis Oliveti coeperunt omnes turbae discentium gaudentes laudare Deum voce magna super omnibus quas viderant virtutibus
LUKE|19|38|dicentes benedictus qui venit rex in nomine Domini pax in caelo et gloria in excelsis
LUKE|19|39|et quidam Pharisaeorum de turbis dixerunt ad illum magister increpa discipulos tuos
LUKE|19|40|quibus ipse ait dico vobis quia si hii tacuerint lapides clamabunt
LUKE|19|41|et ut adpropinquavit videns civitatem flevit super illam dicens
LUKE|19|42|quia si cognovisses et tu et quidem in hac die tua quae ad pacem tibi nunc autem abscondita sunt ab oculis tuis
LUKE|19|43|quia venient dies in te et circumdabunt te inimici tui vallo et circumdabunt te et coangustabunt te undique
LUKE|19|44|ad terram prosternent te et filios qui in te sunt et non relinquent in te lapidem super lapidem eo quod non cognoveris tempus visitationis tuae
LUKE|19|45|et ingressus in templum coepit eicere vendentes in illo et ementes
LUKE|19|46|dicens illis scriptum est quia domus mea domus orationis est vos autem fecistis illam speluncam latronum
LUKE|19|47|et erat docens cotidie in templo principes autem sacerdotum et scribae et principes plebis quaerebant illum perdere
LUKE|19|48|et non inveniebant quid facerent illi omnis enim populus suspensus erat audiens illum
LUKE|20|1|et factum est in una dierum docente illo populum in templo et evangelizante convenerunt principes sacerdotum et scribae cum senioribus
LUKE|20|2|et aiunt dicentes ad illum dic nobis in qua potestate haec facis aut quis est qui dedit tibi hanc potestatem
LUKE|20|3|respondens autem dixit ad illos interrogabo vos et ego verbum respondete mihi
LUKE|20|4|baptismum Iohannis de caelo erat an ex hominibus
LUKE|20|5|at illi cogitabant inter se dicentes quia si dixerimus de caelo dicet quare ergo non credidistis illi
LUKE|20|6|si autem dixerimus ex hominibus plebs universa lapidabit nos certi sunt enim Iohannem prophetam esse
LUKE|20|7|et responderunt se nescire unde esset
LUKE|20|8|et Iesus ait illis neque ego dico vobis in qua potestate haec facio
LUKE|20|9|coepit autem dicere ad plebem parabolam hanc homo plantavit vineam et locavit eam colonis et ipse peregre fuit multis temporibus
LUKE|20|10|et in tempore misit ad cultores servum ut de fructu vineae darent illi qui caesum dimiserunt eum inanem
LUKE|20|11|et addidit alterum servum mittere illi autem hunc quoque caedentes et adficientes contumelia dimiserunt inanem
LUKE|20|12|et addidit tertium mittere qui et illum vulnerantes eiecerunt
LUKE|20|13|dixit autem dominus vineae quid faciam mittam filium meum dilectum forsitan cum hunc viderint verebuntur
LUKE|20|14|quem cum vidissent coloni cogitaverunt inter se dicentes hic est heres occidamus illum ut nostra fiat hereditas
LUKE|20|15|et eiectum illum extra vineam occiderunt quid ergo faciet illis dominus vineae
LUKE|20|16|veniet et perdet colonos istos et dabit vineam aliis quo audito dixerunt illi absit
LUKE|20|17|ille autem aspiciens eos ait quid est ergo hoc quod scriptum est lapidem quem reprobaverunt aedificantes hic factus est in caput anguli
LUKE|20|18|omnis qui ceciderit supra illum lapidem conquassabitur supra quem autem ceciderit comminuet illum
LUKE|20|19|et quaerebant principes sacerdotum et scribae mittere in illum manus illa hora et timuerunt populum cognoverunt enim quod ad ipsos dixerit similitudinem istam
LUKE|20|20|et observantes miserunt insidiatores qui se iustos simularent ut caperent eum in sermone et traderent illum principatui et potestati praesidis
LUKE|20|21|et interrogaverunt illum dicentes magister scimus quia recte dicis et doces et non accipis personam sed in veritate viam Dei doces
LUKE|20|22|licet nobis dare tributum Caesari an non
LUKE|20|23|considerans autem dolum illorum dixit ad eos quid me temptatis
LUKE|20|24|ostendite mihi denarium cuius habet imaginem et inscriptionem respondentes dixerunt Caesaris
LUKE|20|25|et ait illis reddite ergo quae Caesaris sunt Caesari et quae Dei sunt Deo
LUKE|20|26|et non potuerunt verbum eius reprehendere coram plebe et mirati in responso eius tacuerunt
LUKE|20|27|accesserunt autem quidam Sadducaeorum qui negant esse resurrectionem et interrogaverunt eum
LUKE|20|28|dicentes magister Moses scripsit nobis si frater alicuius mortuus fuerit habens uxorem et hic sine filiis fuerit ut accipiat eam frater eius uxorem et suscitet semen fratri suo
LUKE|20|29|septem ergo fratres erant et primus accepit uxorem et mortuus est sine filiis
LUKE|20|30|et sequens accepit illam et ipse mortuus est sine filio
LUKE|20|31|et tertius accepit illam similiter et omnes septem et non reliquerunt semen et mortui sunt
LUKE|20|32|novissima omnium mortua est et mulier
LUKE|20|33|in resurrectione ergo cuius eorum erit uxor siquidem septem habuerunt eam uxorem
LUKE|20|34|et ait illis Iesus filii saeculi huius nubunt et traduntur ad nuptias
LUKE|20|35|illi autem qui digni habebuntur saeculo illo et resurrectione ex mortuis neque nubunt neque ducunt uxores
LUKE|20|36|neque enim ultra mori poterunt aequales enim angelis sunt et filii sunt Dei cum sint filii resurrectionis
LUKE|20|37|quia vero resurgant mortui et Moses ostendit secus rubum sicut dicit Dominum Deum Abraham et Deum Isaac et Deum Iacob
LUKE|20|38|Deus autem non est mortuorum sed vivorum omnes enim vivunt ei
LUKE|20|39|respondentes autem quidam scribarum dixerunt magister bene dixisti
LUKE|20|40|et amplius non audebant eum quicquam interrogare
LUKE|20|41|dixit autem ad illos quomodo dicunt Christum Filium David esse
LUKE|20|42|et ipse David dicit in libro Psalmorum dixit Dominus Domino meo sede a dextris meis
LUKE|20|43|donec ponam inimicos tuos scabillum pedum tuorum
LUKE|20|44|David ergo Dominum illum vocat et quomodo filius eius est
LUKE|20|45|audiente autem omni populo dixit discipulis suis
LUKE|20|46|adtendite a scribis qui volunt ambulare in stolis et amant salutationes in foro et primas cathedras in synagogis et primos discubitus in conviviis
LUKE|20|47|qui devorant domos viduarum simulantes longam orationem hii accipient damnationem maiorem
LUKE|21|1|respiciens autem vidit eos qui mittebant munera sua in gazofilacium divites
LUKE|21|2|vidit autem et quandam viduam pauperculam mittentem aera minuta duo
LUKE|21|3|et dixit vere dico vobis quia vidua haec pauper plus quam omnes misit
LUKE|21|4|nam omnes hii ex abundanti sibi miserunt in munera Dei haec autem ex eo quod deest illi omnem victum suum quem habuit misit
LUKE|21|5|et quibusdam dicentibus de templo quod lapidibus bonis et donis ornatum esset dixit
LUKE|21|6|haec quae videtis venient dies in quibus non relinquetur lapis super lapidem qui non destruatur
LUKE|21|7|interrogaverunt autem illum dicentes praeceptor quando haec erunt et quod signum cum fieri incipient
LUKE|21|8|qui dixit videte ne seducamini multi enim venient in nomine meo dicentes quia ego sum et tempus adpropinquavit nolite ergo ire post illos
LUKE|21|9|cum autem audieritis proelia et seditiones nolite terreri oportet primum haec fieri sed non statim finis
LUKE|21|10|tunc dicebat illis surget gens contra gentem et regnum adversus regnum
LUKE|21|11|terraemotus magni erunt per loca et pestilentiae et fames terroresque de caelo et signa magna erunt
LUKE|21|12|sed ante haec omnia inicient vobis manus suas et persequentur tradentes in synagogas et custodias trahentes ad reges et praesides propter nomen meum
LUKE|21|13|continget autem vobis in testimonium
LUKE|21|14|ponite ergo in cordibus vestris non praemeditari quemadmodum respondeatis
LUKE|21|15|ego enim dabo vobis os et sapientiam cui non poterunt resistere et contradicere omnes adversarii vestri
LUKE|21|16|trademini autem a parentibus et fratribus et cognatis et amicis et morte adficient ex vobis
LUKE|21|17|et eritis odio omnibus propter nomen meum
LUKE|21|18|et capillus de capite vestro non peribit
LUKE|21|19|in patientia vestra possidebitis animas vestras
LUKE|21|20|cum autem videritis circumdari ab exercitu Hierusalem tunc scitote quia adpropinquavit desolatio eius
LUKE|21|21|tunc qui in Iudaea sunt fugiant in montes et qui in medio eius discedant et qui in regionibus non intrent in eam
LUKE|21|22|quia dies ultionis hii sunt ut impleantur omnia quae scripta sunt
LUKE|21|23|vae autem praegnatibus et nutrientibus in illis diebus erit enim pressura magna supra terram et ira populo huic
LUKE|21|24|et cadent in ore gladii et captivi ducentur in omnes gentes et Hierusalem calcabitur a gentibus donec impleantur tempora nationum
LUKE|21|25|et erunt signa in sole et luna et stellis et in terris pressura gentium prae confusione sonitus maris et fluctuum
LUKE|21|26|arescentibus hominibus prae timore et expectatione quae supervenient universo orbi nam virtutes caelorum movebuntur
LUKE|21|27|et tunc videbunt Filium hominis venientem in nube cum potestate magna et maiestate
LUKE|21|28|his autem fieri incipientibus respicite et levate capita vestra quoniam adpropinquat redemptio vestra
LUKE|21|29|et dixit illis similitudinem videte ficulneam et omnes arbores
LUKE|21|30|cum producunt iam ex se fructum scitis quoniam prope est aestas
LUKE|21|31|ita et vos cum videritis haec fieri scitote quoniam prope est regnum Dei
LUKE|21|32|amen dico vobis quia non praeteribit generatio haec donec omnia fiant
LUKE|21|33|caelum et terra transibunt verba autem mea non transient
LUKE|21|34|adtendite autem vobis ne forte graventur corda vestra in crapula et ebrietate et curis huius vitae et superveniat in vos repentina dies illa
LUKE|21|35|tamquam laqueus enim superveniet in omnes qui sedent super faciem omnis terrae
LUKE|21|36|vigilate itaque omni tempore orantes ut digni habeamini fugere ista omnia quae futura sunt et stare ante Filium hominis
LUKE|21|37|erat autem diebus docens in templo noctibus vero exiens morabatur in monte qui vocatur Oliveti
LUKE|21|38|et omnis populus manicabat ad eum in templo audire eum
LUKE|22|1|adpropinquabat autem dies festus azymorum qui dicitur pascha
LUKE|22|2|et quaerebant principes sacerdotum et scribae quomodo eum interficerent timebant vero plebem
LUKE|22|3|intravit autem Satanas in Iudam qui cognominatur Scarioth unum de duodecim
LUKE|22|4|et abiit et locutus est cum principibus sacerdotum et magistratibus quemadmodum illum traderet eis
LUKE|22|5|et gavisi sunt et pacti sunt pecuniam illi dare
LUKE|22|6|et spopondit et quaerebat oportunitatem ut traderet illum sine turbis
LUKE|22|7|venit autem dies azymorum in qua necesse erat occidi pascha
LUKE|22|8|et misit Petrum et Iohannem dicens euntes parate nobis pascha ut manducemus
LUKE|22|9|at illi dixerunt ubi vis paremus
LUKE|22|10|et dixit ad eos ecce introeuntibus vobis in civitatem occurret vobis homo amphoram aquae portans sequimini eum in domum in qua intrat
LUKE|22|11|et dicetis patri familias domus dicit tibi magister ubi est diversorium ubi pascha cum discipulis meis manducem
LUKE|22|12|et ipse vobis ostendet cenaculum magnum stratum et ibi parate
LUKE|22|13|euntes autem invenerunt sicut dixit illis et paraverunt pascha
LUKE|22|14|et cum facta esset hora discubuit et duodecim apostoli cum eo
LUKE|22|15|et ait illis desiderio desideravi hoc pascha manducare vobiscum antequam patiar
LUKE|22|16|dico enim vobis quia ex hoc non manducabo illud donec impleatur in regno Dei
LUKE|22|17|et accepto calice gratias egit et dixit accipite et dividite inter vos
LUKE|22|18|dico enim vobis quod non bibam de generatione vitis donec regnum Dei veniat
LUKE|22|19|et accepto pane gratias egit et fregit et dedit eis dicens hoc est corpus meum quod pro vobis datur hoc facite in meam commemorationem
LUKE|22|20|similiter et calicem postquam cenavit dicens hic est calix novum testamentum in sanguine meo quod pro vobis funditur
LUKE|22|21|verumtamen ecce manus tradentis me mecum est in mensa
LUKE|22|22|et quidem Filius hominis secundum quod definitum est vadit verumtamen vae illi homini per quem traditur
LUKE|22|23|et ipsi coeperunt quaerere inter se quis esset ex eis qui hoc facturus esset
LUKE|22|24|facta est autem et contentio inter eos quis eorum videretur esse maior
LUKE|22|25|dixit autem eis reges gentium dominantur eorum et qui potestatem habent super eos benefici vocantur
LUKE|22|26|vos autem non sic sed qui maior est in vobis fiat sicut iunior et qui praecessor est sicut ministrator
LUKE|22|27|nam quis maior est qui recumbit an qui ministrat nonne qui recumbit ego autem in medio vestrum sum sicut qui ministrat
LUKE|22|28|vos autem estis qui permansistis mecum in temptationibus meis
LUKE|22|29|et ego dispono vobis sicut disposuit mihi Pater meus regnum
LUKE|22|30|ut edatis et bibatis super mensam meam in regno et sedeatis super thronos iudicantes duodecim tribus Israhel
LUKE|22|31|ait autem Dominus Simon Simon ecce Satanas expetivit vos ut cribraret sicut triticum
LUKE|22|32|ego autem rogavi pro te ut non deficiat fides tua et tu aliquando conversus confirma fratres tuos
LUKE|22|33|qui dixit ei Domine tecum paratus sum et in carcerem et in mortem ire
LUKE|22|34|et ille dixit dico tibi Petre non cantabit hodie gallus donec ter abneges nosse me
LUKE|22|35|et dixit eis quando misi vos sine sacculo et pera et calciamentis numquid aliquid defuit vobis at illi dixerunt nihil
LUKE|22|36|dixit ergo eis sed nunc qui habet sacculum tollat similiter et peram et qui non habet vendat tunicam suam et emat gladium
LUKE|22|37|dico enim vobis quoniam adhuc hoc quod scriptum est oportet impleri in me et quod cum iniustis deputatus est etenim ea quae sunt de me finem habent
LUKE|22|38|at illi dixerunt Domine ecce gladii duo hic at ille dixit eis satis est
LUKE|22|39|et egressus ibat secundum consuetudinem in montem Olivarum secuti sunt autem illum et discipuli
LUKE|22|40|et cum pervenisset ad locum dixit illis orate ne intretis in temptationem
LUKE|22|41|et ipse avulsus est ab eis quantum iactus est lapidis et positis genibus orabat
LUKE|22|42|dicens Pater si vis transfer calicem istum a me verumtamen non mea voluntas sed tua fiat
LUKE|22|43|apparuit autem illi angelus de caelo confortans eum et factus in agonia prolixius orabat
LUKE|22|44|et factus est sudor eius sicut guttae sanguinis decurrentis in terram
LUKE|22|45|et cum surrexisset ab oratione et venisset ad discipulos suos invenit eos dormientes prae tristitia
LUKE|22|46|et ait illis quid dormitis surgite orate ne intretis in temptationem
LUKE|22|47|adhuc eo loquente ecce turba et qui vocabatur Iudas unus de duodecim antecedebat eos et adpropinquavit Iesu ut oscularetur eum
LUKE|22|48|Iesus autem dixit ei Iuda osculo Filium hominis tradis
LUKE|22|49|videntes autem hii qui circa ipsum erant quod futurum erat dixerunt ei Domine si percutimus in gladio
LUKE|22|50|et percussit unus ex illis servum principis sacerdotum et amputavit auriculam eius dextram
LUKE|22|51|respondens autem Iesus ait sinite usque huc et cum tetigisset auriculam eius sanavit eum
LUKE|22|52|dixit autem Iesus ad eos qui venerant ad se principes sacerdotum et magistratus templi et seniores quasi ad latronem existis cum gladiis et fustibus
LUKE|22|53|cum cotidie vobiscum fuerim in templo non extendistis manus in me sed haec est hora vestra et potestas tenebrarum
LUKE|22|54|conprehendentes autem eum duxerunt ad domum principis sacerdotum Petrus vero sequebatur a longe
LUKE|22|55|accenso autem igni in medio atrio et circumsedentibus illis erat Petrus in medio eorum
LUKE|22|56|quem cum vidisset ancilla quaedam sedentem ad lumen et eum fuisset intuita dixit et hic cum illo erat
LUKE|22|57|at ille negavit eum dicens mulier non novi illum
LUKE|22|58|et post pusillum alius videns eum dixit et tu de illis es Petrus vero ait o homo non sum
LUKE|22|59|et intervallo facto quasi horae unius alius quidam adfirmabat dicens vere et hic cum illo erat nam et Galilaeus est
LUKE|22|60|et ait Petrus homo nescio quod dicis et continuo adhuc illo loquente cantavit gallus
LUKE|22|61|et conversus Dominus respexit Petrum et recordatus est Petrus verbi Domini sicut dixit quia priusquam gallus cantet ter me negabis
LUKE|22|62|et egressus foras Petrus flevit amare
LUKE|22|63|et viri qui tenebant illum inludebant ei caedentes
LUKE|22|64|et velaverunt eum et percutiebant faciem eius et interrogabant eum dicentes prophetiza quis est qui te percussit
LUKE|22|65|et alia multa blasphemantes dicebant in eum
LUKE|22|66|et ut factus est dies convenerunt seniores plebis et principes sacerdotum et scribae et duxerunt illum in concilium suum dicentes si tu es Christus dic nobis
LUKE|22|67|et ait illis si vobis dixero non creditis mihi
LUKE|22|68|si autem et interrogavero non respondebitis mihi neque dimittetis
LUKE|22|69|ex hoc autem erit Filius hominis sedens a dextris virtutis Dei
LUKE|22|70|dixerunt autem omnes tu ergo es Filius Dei qui ait vos dicitis quia ego sum
LUKE|22|71|at illi dixerunt quid adhuc desideramus testimonium ipsi enim audivimus de ore eius
LUKE|23|1|et surgens omnis multitudo eorum duxerunt illum ad Pilatum
LUKE|23|2|coeperunt autem accusare illum dicentes hunc invenimus subvertentem gentem nostram et prohibentem tributa dari Caesari et dicentem se Christum regem esse
LUKE|23|3|Pilatus autem interrogavit eum dicens tu es rex Iudaeorum at ille respondens ait tu dicis
LUKE|23|4|ait autem Pilatus ad principes sacerdotum et turbas nihil invenio causae in hoc homine
LUKE|23|5|at illi invalescebant dicentes commovet populum docens per universam Iudaeam et incipiens a Galilaea usque huc
LUKE|23|6|Pilatus autem audiens Galilaeam interrogavit si homo Galilaeus esset
LUKE|23|7|et ut cognovit quod de Herodis potestate esset remisit eum ad Herodem qui et ipse Hierosolymis erat illis diebus
LUKE|23|8|Herodes autem viso Iesu gavisus est valde erat enim cupiens ex multo tempore videre eum eo quod audiret multa de illo et sperabat signum aliquod videre ab eo fieri
LUKE|23|9|interrogabat autem illum multis sermonibus at ipse nihil illi respondebat
LUKE|23|10|stabant etiam principes sacerdotum et scribae constanter accusantes eum
LUKE|23|11|sprevit autem illum Herodes cum exercitu suo et inlusit indutum veste alba et remisit ad Pilatum
LUKE|23|12|et facti sunt amici Herodes et Pilatus in ipsa die nam antea inimici erant ad invicem
LUKE|23|13|Pilatus autem convocatis principibus sacerdotum et magistratibus et plebe
LUKE|23|14|dixit ad illos obtulistis mihi hunc hominem quasi avertentem populum et ecce ego coram vobis interrogans nullam causam inveni in homine isto ex his in quibus eum accusatis
LUKE|23|15|sed neque Herodes nam remisi vos ad illum et ecce nihil dignum morte actum est ei
LUKE|23|16|emendatum ergo illum dimittam
LUKE|23|17|necesse autem habebat dimittere eis per diem festum unum
LUKE|23|18|exclamavit autem simul universa turba dicens tolle hunc et dimitte nobis Barabban
LUKE|23|19|qui erat propter seditionem quandam factam in civitate et homicidium missus in carcerem
LUKE|23|20|iterum autem Pilatus locutus est ad illos volens dimittere Iesum
LUKE|23|21|at illi succlamabant dicentes crucifige crucifige illum
LUKE|23|22|ille autem tertio dixit ad illos quid enim mali fecit iste nullam causam mortis invenio in eo corripiam ergo illum et dimittam
LUKE|23|23|at illi instabant vocibus magnis postulantes ut crucifigeretur et invalescebant voces eorum
LUKE|23|24|et Pilatus adiudicavit fieri petitionem eorum
LUKE|23|25|dimisit autem illis eum qui propter homicidium et seditionem missus fuerat in carcerem quem petebant Iesum vero tradidit voluntati eorum
LUKE|23|26|et cum ducerent eum adprehenderunt Simonem quendam Cyrenensem venientem de villa et inposuerunt illi crucem portare post Iesum
LUKE|23|27|sequebatur autem illum multa turba populi et mulierum quae plangebant et lamentabant eum
LUKE|23|28|conversus autem ad illas Iesus dixit filiae Hierusalem nolite flere super me sed super vos ipsas flete et super filios vestros
LUKE|23|29|quoniam ecce venient dies in quibus dicent beatae steriles et ventres qui non genuerunt et ubera quae non lactaverunt
LUKE|23|30|tunc incipient dicere montibus cadite super nos et collibus operite nos
LUKE|23|31|quia si in viridi ligno haec faciunt in arido quid fiet
LUKE|23|32|ducebantur autem et alii duo nequam cum eo ut interficerentur
LUKE|23|33|et postquam venerunt in locum qui vocatur Calvariae ibi crucifixerunt eum et latrones unum a dextris et alterum a sinistris
LUKE|23|34|Iesus autem dicebat Pater dimitte illis non enim sciunt quid faciunt dividentes vero vestimenta eius miserunt sortes
LUKE|23|35|et stabat populus expectans et deridebant illum principes cum eis dicentes alios salvos fecit se salvum faciat si hic est Christus Dei electus
LUKE|23|36|inludebant autem ei et milites accedentes et acetum offerentes illi
LUKE|23|37|dicentes si tu es rex Iudaeorum salvum te fac
LUKE|23|38|erat autem et superscriptio inscripta super illum litteris graecis et latinis et hebraicis hic est rex Iudaeorum
LUKE|23|39|unus autem de his qui pendebant latronibus blasphemabat eum dicens si tu es Christus salvum fac temet ipsum et nos
LUKE|23|40|respondens autem alter increpabat illum dicens neque tu times Deum quod in eadem damnatione es
LUKE|23|41|et nos quidem iuste nam digna factis recipimus hic vero nihil mali gessit
LUKE|23|42|et dicebat ad Iesum Domine memento mei cum veneris in regnum tuum
LUKE|23|43|et dixit illi Iesus amen dico tibi hodie mecum eris in paradiso
LUKE|23|44|erat autem fere hora sexta et tenebrae factae sunt in universa terra usque in nonam horam
LUKE|23|45|et obscuratus est sol et velum templi scissum est medium
LUKE|23|46|et clamans voce magna Iesus ait Pater in manus tuas commendo spiritum meum et haec dicens exspiravit
LUKE|23|47|videns autem centurio quod factum fuerat glorificavit Deum dicens vere hic homo iustus erat
LUKE|23|48|et omnis turba eorum qui simul aderant ad spectaculum istud et videbant quae fiebant percutientes pectora sua revertebantur
LUKE|23|49|stabant autem omnes noti eius a longe et mulieres quae secutae erant eum a Galilaea haec videntes
LUKE|23|50|et ecce vir nomine Ioseph qui erat decurio vir bonus et iustus
LUKE|23|51|hic non consenserat consilio et actibus eorum ab Arimathia civitate Iudaeae qui expectabat et ipse regnum Dei
LUKE|23|52|hic accessit ad Pilatum et petiit corpus Iesu
LUKE|23|53|et depositum involvit sindone et posuit eum in monumento exciso in quo nondum quisquam positus fuerat
LUKE|23|54|et dies erat parasceves et sabbatum inlucescebat
LUKE|23|55|subsecutae autem mulieres quae cum ipso venerant de Galilaea viderunt monumentum et quemadmodum positum erat corpus eius
LUKE|23|56|et revertentes paraverunt aromata et unguenta et sabbato quidem siluerunt secundum mandatum
LUKE|24|1|una autem sabbati valde diluculo venerunt ad monumentum portantes quae paraverant aromata
LUKE|24|2|et invenerunt lapidem revolutum a monumento
LUKE|24|3|et ingressae non invenerunt corpus Domini Iesu
LUKE|24|4|et factum est dum mente consternatae essent de isto ecce duo viri steterunt secus illas in veste fulgenti
LUKE|24|5|cum timerent autem et declinarent vultum in terram dixerunt ad illas quid quaeritis viventem cum mortuis
LUKE|24|6|non est hic sed surrexit recordamini qualiter locutus est vobis cum adhuc in Galilaea esset
LUKE|24|7|dicens quia oportet Filium hominis tradi in manus hominum peccatorum et crucifigi et die tertia resurgere
LUKE|24|8|et recordatae sunt verborum eius
LUKE|24|9|et regressae a monumento nuntiaverunt haec omnia illis undecim et ceteris omnibus
LUKE|24|10|erat autem Maria Magdalene et Iohanna et Maria Iacobi et ceterae quae cum eis erant quae dicebant ad apostolos haec
LUKE|24|11|et visa sunt ante illos sicut deliramentum verba ista et non credebant illis
LUKE|24|12|Petrus autem surgens cucurrit ad monumentum et procumbens videt linteamina sola posita et abiit secum mirans quod factum fuerat
LUKE|24|13|et ecce duo ex illis ibant ipsa die in castellum quod erat in spatio stadiorum sexaginta ab Hierusalem nomine Emmaus
LUKE|24|14|et ipsi loquebantur ad invicem de his omnibus quae acciderant
LUKE|24|15|et factum est dum fabularentur et secum quaererent et ipse Iesus adpropinquans ibat cum illis
LUKE|24|16|oculi autem illorum tenebantur ne eum agnoscerent
LUKE|24|17|et ait ad illos qui sunt hii sermones quos confertis ad invicem ambulantes et estis tristes
LUKE|24|18|et respondens unus cui nomen Cleopas dixit ei tu solus peregrinus es in Hierusalem et non cognovisti quae facta sunt in illa his diebus
LUKE|24|19|quibus ille dixit quae et dixerunt de Iesu Nazareno qui fuit vir propheta potens in opere et sermone coram Deo et omni populo
LUKE|24|20|et quomodo eum tradiderunt summi sacerdotum et principes nostri in damnationem mortis et crucifixerunt eum
LUKE|24|21|nos autem sperabamus quia ipse esset redempturus Israhel et nunc super haec omnia tertia dies hodie quod haec facta sunt
LUKE|24|22|sed et mulieres quaedam ex nostris terruerunt nos quae ante lucem fuerunt ad monumentum
LUKE|24|23|et non invento corpore eius venerunt dicentes se etiam visionem angelorum vidisse qui dicunt eum vivere
LUKE|24|24|et abierunt quidam ex nostris ad monumentum et ita invenerunt sicut mulieres dixerunt ipsum vero non viderunt
LUKE|24|25|et ipse dixit ad eos o stulti et tardi corde ad credendum in omnibus quae locuti sunt prophetae
LUKE|24|26|nonne haec oportuit pati Christum et ita intrare in gloriam suam
LUKE|24|27|et incipiens a Mose et omnibus prophetis interpretabatur illis in omnibus scripturis quae de ipso erant
LUKE|24|28|et adpropinquaverunt castello quo ibant et ipse se finxit longius ire
LUKE|24|29|et coegerunt illum dicentes mane nobiscum quoniam advesperascit et inclinata est iam dies et intravit cum illis
LUKE|24|30|et factum est dum recumberet cum illis accepit panem et benedixit ac fregit et porrigebat illis
LUKE|24|31|et aperti sunt oculi eorum et cognoverunt eum et ipse evanuit ex oculis eorum
LUKE|24|32|et dixerunt ad invicem nonne cor nostrum ardens erat in nobis dum loqueretur in via et aperiret nobis scripturas
LUKE|24|33|et surgentes eadem hora regressi sunt in Hierusalem et invenerunt congregatos undecim et eos qui cum ipsis erant
LUKE|24|34|dicentes quod surrexit Dominus vere et apparuit Simoni
LUKE|24|35|et ipsi narrabant quae gesta erant in via et quomodo cognoverunt eum in fractione panis
LUKE|24|36|dum haec autem loquuntur Iesus stetit in medio eorum et dicit eis pax vobis ego sum nolite timere
LUKE|24|37|conturbati vero et conterriti existimabant se spiritum videre
LUKE|24|38|et dixit eis quid turbati estis et cogitationes ascendunt in corda vestra
LUKE|24|39|videte manus meas et pedes quia ipse ego sum palpate et videte quia spiritus carnem et ossa non habet sicut me videtis habere
LUKE|24|40|et cum hoc dixisset ostendit eis manus et pedes
LUKE|24|41|adhuc autem illis non credentibus et mirantibus prae gaudio dixit habetis hic aliquid quod manducetur
LUKE|24|42|at illi obtulerunt ei partem piscis assi et favum mellis
LUKE|24|43|et cum manducasset coram eis sumens reliquias dedit eis
LUKE|24|44|et dixit ad eos haec sunt verba quae locutus sum ad vos cum adhuc essem vobiscum quoniam necesse est impleri omnia quae scripta sunt in lege Mosi et prophetis et psalmis de me
LUKE|24|45|tunc aperuit illis sensum ut intellegerent scripturas
LUKE|24|46|et dixit eis quoniam sic scriptum est et sic oportebat Christum pati et resurgere a mortuis die tertia
LUKE|24|47|et praedicari in nomine eius paenitentiam et remissionem peccatorum in omnes gentes incipientibus ab Hierosolyma
LUKE|24|48|vos autem estis testes horum
LUKE|24|49|et ego mitto promissum Patris mei in vos vos autem sedete in civitate quoadusque induamini virtutem ex alto
LUKE|24|50|eduxit autem eos foras in Bethaniam et elevatis manibus suis benedixit eis
LUKE|24|51|et factum est dum benediceret illis recessit ab eis et ferebatur in caelum
LUKE|24|52|et ipsi adorantes regressi sunt in Hierusalem cum gaudio magno
LUKE|24|53|et erant semper in templo laudantes et benedicentes Deum amen
JOHN|1|1|in principio erat Verbum et Verbum erat apud Deum et Deus erat Verbum
JOHN|1|2|hoc erat in principio apud Deum
JOHN|1|3|omnia per ipsum facta sunt et sine ipso factum est nihil quod factum est
JOHN|1|4|in ipso vita erat et vita erat lux hominum
JOHN|1|5|et lux in tenebris lucet et tenebrae eam non conprehenderunt
JOHN|1|6|fuit homo missus a Deo cui nomen erat Iohannes
JOHN|1|7|hic venit in testimonium ut testimonium perhiberet de lumine ut omnes crederent per illum
JOHN|1|8|non erat ille lux sed ut testimonium perhiberet de lumine
JOHN|1|9|erat lux vera quae inluminat omnem hominem venientem in mundum
JOHN|1|10|in mundo erat et mundus per ipsum factus est et mundus eum non cognovit
JOHN|1|11|in propria venit et sui eum non receperunt
JOHN|1|12|quotquot autem receperunt eum dedit eis potestatem filios Dei fieri his qui credunt in nomine eius
JOHN|1|13|qui non ex sanguinibus neque ex voluntate carnis neque ex voluntate viri sed ex Deo nati sunt
JOHN|1|14|et Verbum caro factum est et habitavit in nobis et vidimus gloriam eius gloriam quasi unigeniti a Patre plenum gratiae et veritatis
JOHN|1|15|Iohannes testimonium perhibet de ipso et clamat dicens hic erat quem dixi vobis qui post me venturus est ante me factus est quia prior me erat
JOHN|1|16|et de plenitudine eius nos omnes accepimus et gratiam pro gratia
JOHN|1|17|quia lex per Mosen data est gratia et veritas per Iesum Christum facta est
JOHN|1|18|Deum nemo vidit umquam unigenitus Filius qui est in sinu Patris ipse enarravit
JOHN|1|19|et hoc est testimonium Iohannis quando miserunt Iudaei ab Hierosolymis sacerdotes et Levitas ad eum ut interrogarent eum tu quis es
JOHN|1|20|et confessus est et non negavit et confessus est quia non sum ego Christus
JOHN|1|21|et interrogaverunt eum quid ergo Helias es tu et dicit non sum propheta es tu et respondit non
JOHN|1|22|dixerunt ergo ei quis es ut responsum demus his qui miserunt nos quid dicis de te ipso
JOHN|1|23|ait ego vox clamantis in deserto dirigite viam Domini sicut dixit Esaias propheta
JOHN|1|24|et qui missi fuerant erant ex Pharisaeis
JOHN|1|25|et interrogaverunt eum et dixerunt ei quid ergo baptizas si tu non es Christus neque Helias neque propheta
JOHN|1|26|respondit eis Iohannes dicens ego baptizo in aqua medius autem vestrum stetit quem vos non scitis
JOHN|1|27|ipse est qui post me venturus est qui ante me factus est cuius ego non sum dignus ut solvam eius corrigiam calciamenti
JOHN|1|28|haec in Bethania facta sunt trans Iordanen ubi erat Iohannes baptizans
JOHN|1|29|altera die videt Iohannes Iesum venientem ad se et ait ecce agnus Dei qui tollit peccatum mundi
JOHN|1|30|hic est de quo dixi post me venit vir qui ante me factus est quia prior me erat
JOHN|1|31|et ego nesciebam eum sed ut manifestaretur Israhel propterea veni ego in aqua baptizans
JOHN|1|32|et testimonium perhibuit Iohannes dicens quia vidi Spiritum descendentem quasi columbam de caelo et mansit super eum
JOHN|1|33|et ego nesciebam eum sed qui misit me baptizare in aqua ille mihi dixit super quem videris Spiritum descendentem et manentem super eum hic est qui baptizat in Spiritu Sancto
JOHN|1|34|et ego vidi et testimonium perhibui quia hic est Filius Dei
JOHN|1|35|altera die iterum stabat Iohannes et ex discipulis eius duo
JOHN|1|36|et respiciens Iesum ambulantem dicit ecce agnus Dei
JOHN|1|37|et audierunt eum duo discipuli loquentem et secuti sunt Iesum
JOHN|1|38|conversus autem Iesus et videns eos sequentes dicit eis quid quaeritis qui dixerunt ei rabbi quod dicitur interpretatum magister ubi habitas
JOHN|1|39|dicit eis venite et videte venerunt et viderunt ubi maneret et apud eum manserunt die illo hora autem erat quasi decima
JOHN|1|40|erat autem Andreas frater Simonis Petri unus ex duobus qui audierant ab Iohanne et secuti fuerant eum
JOHN|1|41|invenit hic primum fratrem suum Simonem et dicit ei invenimus Messiam quod est interpretatum Christus
JOHN|1|42|et adduxit eum ad Iesum intuitus autem eum Iesus dixit tu es Simon filius Iohanna tu vocaberis Cephas quod interpretatur Petrus
JOHN|1|43|in crastinum voluit exire in Galilaeam et invenit Philippum et dicit ei Iesus sequere me
JOHN|1|44|erat autem Philippus a Bethsaida civitate Andreae et Petri
JOHN|1|45|invenit Philippus Nathanahel et dicit ei quem scripsit Moses in lege et prophetae invenimus Iesum filium Ioseph a Nazareth
JOHN|1|46|et dixit ei Nathanahel a Nazareth potest aliquid boni esse dicit ei Philippus veni et vide
JOHN|1|47|vidit Iesus Nathanahel venientem ad se et dicit de eo ecce vere Israhelita in quo dolus non est
JOHN|1|48|dicit ei Nathanahel unde me nosti respondit Iesus et dixit ei priusquam te Philippus vocaret cum esses sub ficu vidi te
JOHN|1|49|respondit ei Nathanahel et ait rabbi tu es Filius Dei tu es rex Israhel
JOHN|1|50|respondit Iesus et dixit ei quia dixi tibi vidi te sub ficu credis maius his videbis
JOHN|1|51|et dicit ei amen amen dico vobis videbitis caelum apertum et angelos Dei ascendentes et descendentes supra Filium hominis
JOHN|2|1|et die tertio nuptiae factae sunt in Cana Galilaeae et erat mater Iesu ibi
JOHN|2|2|vocatus est autem ibi et Iesus et discipuli eius ad nuptias
JOHN|2|3|et deficiente vino dicit mater Iesu ad eum vinum non habent
JOHN|2|4|et dicit ei Iesus quid mihi et tibi est mulier nondum venit hora mea
JOHN|2|5|dicit mater eius ministris quodcumque dixerit vobis facite
JOHN|2|6|erant autem ibi lapideae hydriae sex positae secundum purificationem Iudaeorum capientes singulae metretas binas vel ternas
JOHN|2|7|dicit eis Iesus implete hydrias aqua et impleverunt eas usque ad summum
JOHN|2|8|et dicit eis Iesus haurite nunc et ferte architriclino et tulerunt
JOHN|2|9|ut autem gustavit architriclinus aquam vinum factam et non sciebat unde esset ministri autem sciebant qui haurierant aquam vocat sponsum architriclinus
JOHN|2|10|et dicit ei omnis homo primum bonum vinum ponit et cum inebriati fuerint tunc id quod deterius est tu servasti bonum vinum usque adhuc
JOHN|2|11|hoc fecit initium signorum Iesus in Cana Galilaeae et manifestavit gloriam suam et crediderunt in eum discipuli eius
JOHN|2|12|post hoc descendit Capharnaum ipse et mater eius et fratres eius et discipuli eius et ibi manserunt non multis diebus
JOHN|2|13|et prope erat pascha Iudaeorum et ascendit Hierosolyma Iesus
JOHN|2|14|et invenit in templo vendentes boves et oves et columbas et nummularios sedentes
JOHN|2|15|et cum fecisset quasi flagellum de funiculis omnes eiecit de templo oves quoque et boves et nummulariorum effudit aes et mensas subvertit
JOHN|2|16|et his qui columbas vendebant dixit auferte ista hinc nolite facere domum Patris mei domum negotiationis
JOHN|2|17|recordati vero sunt discipuli eius quia scriptum est zelus domus tuae comedit me
JOHN|2|18|responderunt ergo Iudaei et dixerunt ei quod signum ostendis nobis quia haec facis
JOHN|2|19|respondit Iesus et dixit eis solvite templum hoc et in tribus diebus excitabo illud
JOHN|2|20|dixerunt ergo Iudaei quadraginta et sex annis aedificatum est templum hoc et tu tribus diebus excitabis illud
JOHN|2|21|ille autem dicebat de templo corporis sui
JOHN|2|22|cum ergo resurrexisset a mortuis recordati sunt discipuli eius quia hoc dicebat et crediderunt scripturae et sermoni quem dixit Iesus
JOHN|2|23|cum autem esset Hierosolymis in pascha in die festo multi crediderunt in nomine eius videntes signa eius quae faciebat
JOHN|2|24|ipse autem Iesus non credebat semet ipsum eis eo quod ipse nosset omnes
JOHN|2|25|et quia opus ei non erat ut quis testimonium perhiberet de homine ipse enim sciebat quid esset in homine
JOHN|3|1|erat autem homo ex Pharisaeis Nicodemus nomine princeps Iudaeorum
JOHN|3|2|hic venit ad eum nocte et dixit ei rabbi scimus quia a Deo venisti magister nemo enim potest haec signa facere quae tu facis nisi fuerit Deus cum eo
JOHN|3|3|respondit Iesus et dixit ei amen amen dico tibi nisi quis natus fuerit denuo non potest videre regnum Dei
JOHN|3|4|dicit ad eum Nicodemus quomodo potest homo nasci cum senex sit numquid potest in ventrem matris suae iterato introire et nasci
JOHN|3|5|respondit Iesus amen amen dico tibi nisi quis renatus fuerit ex aqua et Spiritu non potest introire in regnum Dei
JOHN|3|6|quod natum est ex carne caro est et quod natum est ex Spiritu spiritus est
JOHN|3|7|non mireris quia dixi tibi oportet vos nasci denuo
JOHN|3|8|Spiritus ubi vult spirat et vocem eius audis sed non scis unde veniat et quo vadat sic est omnis qui natus est ex Spiritu
JOHN|3|9|respondit Nicodemus et dixit ei quomodo possunt haec fieri
JOHN|3|10|respondit Iesus et dixit ei tu es magister Israhel et haec ignoras
JOHN|3|11|amen amen dico tibi quia quod scimus loquimur et quod vidimus testamur et testimonium nostrum non accipitis
JOHN|3|12|si terrena dixi vobis et non creditis quomodo si dixero vobis caelestia credetis
JOHN|3|13|et nemo ascendit in caelum nisi qui descendit de caelo Filius hominis qui est in caelo
JOHN|3|14|et sicut Moses exaltavit serpentem in deserto ita exaltari oportet Filium hominis
JOHN|3|15|ut omnis qui credit in ipso non pereat sed habeat vitam aeternam
JOHN|3|16|sic enim dilexit Deus mundum ut Filium suum unigenitum daret ut omnis qui credit in eum non pereat sed habeat vitam aeternam
JOHN|3|17|non enim misit Deus Filium suum in mundum ut iudicet mundum sed ut salvetur mundus per ipsum
JOHN|3|18|qui credit in eum non iudicatur qui autem non credit iam iudicatus est quia non credidit in nomine unigeniti Filii Dei
JOHN|3|19|hoc est autem iudicium quia lux venit in mundum et dilexerunt homines magis tenebras quam lucem erant enim eorum mala opera
JOHN|3|20|omnis enim qui mala agit odit lucem et non venit ad lucem ut non arguantur opera eius
JOHN|3|21|qui autem facit veritatem venit ad lucem ut manifestentur eius opera quia in Deo sunt facta
JOHN|3|22|post haec venit Iesus et discipuli eius in iudaeam terram et illic demorabatur cum eis et baptizabat
JOHN|3|23|erat autem et Iohannes baptizans in Aenon iuxta Salim quia aquae multae erant illic et adveniebant et baptizabantur
JOHN|3|24|nondum enim missus fuerat in carcerem Iohannes
JOHN|3|25|facta est ergo quaestio ex discipulis Iohannis cum Iudaeis de purificatione
JOHN|3|26|et venerunt ad Iohannem et dixerunt ei rabbi qui erat tecum trans Iordanen cui tu testimonium perhibuisti ecce hic baptizat et omnes veniunt ad eum
JOHN|3|27|respondit Iohannes et dixit non potest homo accipere quicquam nisi fuerit ei datum de caelo
JOHN|3|28|ipsi vos mihi testimonium perhibetis quod dixerim ego non sum Christus sed quia missus sum ante illum
JOHN|3|29|qui habet sponsam sponsus est amicus autem sponsi qui stat et audit eum gaudio gaudet propter vocem sponsi hoc ergo gaudium meum impletum est
JOHN|3|30|illum oportet crescere me autem minui
JOHN|3|31|qui desursum venit supra omnes est qui est de terra de terra est et de terra loquitur qui de caelo venit supra omnes est
JOHN|3|32|et quod vidit et audivit hoc testatur et testimonium eius nemo accipit
JOHN|3|33|qui accipit eius testimonium signavit quia Deus verax est
JOHN|3|34|quem enim misit Deus verba Dei loquitur non enim ad mensuram dat Deus Spiritum
JOHN|3|35|Pater diligit Filium et omnia dedit in manu eius
JOHN|3|36|qui credit in Filium habet vitam aeternam qui autem incredulus est Filio non videbit vitam sed ira Dei manet super eum
JOHN|4|1|ut ergo cognovit Iesus quia audierunt Pharisaei quia Iesus plures discipulos facit et baptizat quam Iohannes
JOHN|4|2|quamquam Iesus non baptizaret sed discipuli eius
JOHN|4|3|reliquit Iudaeam et abiit iterum in Galilaeam
JOHN|4|4|oportebat autem eum transire per Samariam
JOHN|4|5|venit ergo in civitatem Samariae quae dicitur Sychar iuxta praedium quod dedit Iacob Ioseph filio suo
JOHN|4|6|erat autem ibi fons Iacob Iesus ergo fatigatus ex itinere sedebat sic super fontem hora erat quasi sexta
JOHN|4|7|venit mulier de Samaria haurire aquam dicit ei Iesus da mihi bibere
JOHN|4|8|discipuli enim eius abierant in civitatem ut cibos emerent
JOHN|4|9|dicit ergo ei mulier illa samaritana quomodo tu Iudaeus cum sis bibere a me poscis quae sum mulier samaritana non enim coutuntur Iudaei Samaritanis
JOHN|4|10|respondit Iesus et dixit ei si scires donum Dei et quis est qui dicit tibi da mihi bibere tu forsitan petisses ab eo et dedisset tibi aquam vivam
JOHN|4|11|dicit ei mulier Domine neque in quo haurias habes et puteus altus est unde ergo habes aquam vivam
JOHN|4|12|numquid tu maior es patre nostro Iacob qui dedit nobis puteum et ipse ex eo bibit et filii eius et pecora eius
JOHN|4|13|respondit Iesus et dixit ei omnis qui bibit ex aqua hac sitiet iterum qui autem biberit ex aqua quam ego dabo ei non sitiet in aeternum
JOHN|4|14|sed aqua quam dabo ei fiet in eo fons aquae salientis in vitam aeternam
JOHN|4|15|dicit ad eum mulier Domine da mihi hanc aquam ut non sitiam neque veniam huc haurire
JOHN|4|16|dicit ei Iesus vade voca virum tuum et veni huc
JOHN|4|17|respondit mulier et dixit non habeo virum dicit ei Iesus bene dixisti quia non habeo virum
JOHN|4|18|quinque enim viros habuisti et nunc quem habes non est tuus vir hoc vere dixisti
JOHN|4|19|dicit ei mulier Domine video quia propheta es tu
JOHN|4|20|patres nostri in monte hoc adoraverunt et vos dicitis quia Hierosolymis est locus ubi adorare oportet
JOHN|4|21|dicit ei Iesus mulier crede mihi quia veniet hora quando neque in monte hoc neque in Hierosolymis adorabitis Patrem
JOHN|4|22|vos adoratis quod nescitis nos adoramus quod scimus quia salus ex Iudaeis est
JOHN|4|23|sed venit hora et nunc est quando veri adoratores adorabunt Patrem in spiritu et veritate nam et Pater tales quaerit qui adorent eum
JOHN|4|24|spiritus est Deus et eos qui adorant eum in spiritu et veritate oportet adorare
JOHN|4|25|dicit ei mulier scio quia Messias venit qui dicitur Christus cum ergo venerit ille nobis adnuntiabit omnia
JOHN|4|26|dicit ei Iesus ego sum qui loquor tecum
JOHN|4|27|et continuo venerunt discipuli eius et mirabantur quia cum muliere loquebatur nemo tamen dixit quid quaeris aut quid loqueris cum ea
JOHN|4|28|reliquit ergo hydriam suam mulier et abiit in civitatem et dicit illis hominibus
JOHN|4|29|venite videte hominem qui dixit mihi omnia quaecumque feci numquid ipse est Christus
JOHN|4|30|exierunt de civitate et veniebant ad eum
JOHN|4|31|interea rogabant eum discipuli dicentes rabbi manduca
JOHN|4|32|ille autem dixit eis ego cibum habeo manducare quem vos nescitis
JOHN|4|33|dicebant ergo discipuli ad invicem numquid aliquis adtulit ei manducare
JOHN|4|34|dicit eis Iesus meus cibus est ut faciam voluntatem eius qui misit me ut perficiam opus eius
JOHN|4|35|nonne vos dicitis quod adhuc quattuor menses sunt et messis venit ecce dico vobis levate oculos vestros et videte regiones quia albae sunt iam ad messem
JOHN|4|36|et qui metit mercedem accipit et congregat fructum in vitam aeternam ut et qui seminat simul gaudeat et qui metit
JOHN|4|37|in hoc enim est verbum verum quia alius est qui seminat et alius est qui metit
JOHN|4|38|ego misi vos metere quod vos non laborastis alii laboraverunt et vos in laborem eorum introistis
JOHN|4|39|ex civitate autem illa multi crediderunt in eum Samaritanorum propter verbum mulieris testimonium perhibentis quia dixit mihi omnia quaecumque feci
JOHN|4|40|cum venissent ergo ad illum Samaritani rogaverunt eum ut ibi maneret et mansit ibi duos dies
JOHN|4|41|et multo plures crediderunt propter sermonem eius
JOHN|4|42|et mulieri dicebant quia iam non propter tuam loquellam credimus ipsi enim audivimus et scimus quia hic est vere salvator mundi
JOHN|4|43|post duos autem dies exiit inde et abiit in Galilaeam
JOHN|4|44|ipse enim Iesus testimonium perhibuit quia propheta in sua patria honorem non habet
JOHN|4|45|cum ergo venisset in Galilaeam exceperunt eum Galilaei cum omnia vidissent quae fecerat Hierosolymis in die festo et ipsi enim venerant in diem festum
JOHN|4|46|venit ergo iterum in Cana Galilaeae ubi fecit aquam vinum et erat quidam regulus cuius filius infirmabatur Capharnaum
JOHN|4|47|hic cum audisset quia Iesus adveniret a Iudaea in Galilaeam abiit ad eum et rogabat eum ut descenderet et sanaret filium eius incipiebat enim mori
JOHN|4|48|dixit ergo Iesus ad eum nisi signa et prodigia videritis non creditis
JOHN|4|49|dicit ad eum regulus Domine descende priusquam moriatur filius meus
JOHN|4|50|dicit ei Iesus vade filius tuus vivit credidit homo sermoni quem dixit ei Iesus et ibat
JOHN|4|51|iam autem eo descendente servi occurrerunt ei et nuntiaverunt dicentes quia filius eius viveret
JOHN|4|52|interrogabat ergo horam ab eis in qua melius habuerit et dixerunt ei quia heri hora septima reliquit eum febris
JOHN|4|53|cognovit ergo pater quia illa hora erat in qua dixit ei Iesus filius tuus vivit et credidit ipse et domus eius tota
JOHN|4|54|hoc iterum secundum signum fecit Iesus cum venisset a Iudaea in Galilaeam
JOHN|5|1|post haec erat dies festus Iudaeorum et ascendit Iesus Hierosolymis
JOHN|5|2|est autem Hierosolymis super Probatica piscina quae cognominatur hebraice Bethsaida quinque porticus habens
JOHN|5|3|in his iacebat multitudo magna languentium caecorum claudorum aridorum expectantium aquae motum
JOHN|5|4|
JOHN|5|5|erat autem quidam homo ibi triginta et octo annos habens in infirmitate sua
JOHN|5|6|hunc cum vidisset Iesus iacentem et cognovisset quia multum iam tempus habet dicit ei vis sanus fieri
JOHN|5|7|respondit ei languidus Domine hominem non habeo ut cum turbata fuerit aqua mittat me in piscinam dum venio enim ego alius ante me descendit
JOHN|5|8|dicit ei Iesus surge tolle grabattum tuum et ambula
JOHN|5|9|et statim sanus factus est homo et sustulit grabattum suum et ambulabat erat autem sabbatum in illo die
JOHN|5|10|dicebant Iudaei illi qui sanatus fuerat sabbatum est non licet tibi tollere grabattum tuum
JOHN|5|11|respondit eis qui me fecit sanum ille mihi dixit tolle grabattum tuum et ambula
JOHN|5|12|interrogaverunt ergo eum quis est ille homo qui dixit tibi tolle grabattum tuum et ambula
JOHN|5|13|is autem qui sanus fuerat effectus nesciebat quis esset Iesus enim declinavit turba constituta in loco
JOHN|5|14|postea invenit eum Iesus in templo et dixit illi ecce sanus factus es iam noli peccare ne deterius tibi aliquid contingat
JOHN|5|15|abiit ille homo et nuntiavit Iudaeis quia Iesus esset qui fecit eum sanum
JOHN|5|16|propterea persequebantur Iudaei Iesum quia haec faciebat in sabbato
JOHN|5|17|Iesus autem respondit eis Pater meus usque modo operatur et ego operor
JOHN|5|18|propterea ergo magis quaerebant eum Iudaei interficere quia non solum solvebat sabbatum sed et Patrem suum dicebat Deum aequalem se faciens Deo respondit itaque Iesus et dixit eis
JOHN|5|19|amen amen dico vobis non potest Filius a se facere quicquam nisi quod viderit Patrem facientem quaecumque enim ille fecerit haec et Filius similiter facit
JOHN|5|20|Pater enim diligit Filium et omnia demonstrat ei quae ipse facit et maiora his demonstrabit ei opera ut vos miremini
JOHN|5|21|sicut enim Pater suscitat mortuos et vivificat sic et Filius quos vult vivificat
JOHN|5|22|neque enim Pater iudicat quemquam sed iudicium omne dedit Filio
JOHN|5|23|ut omnes honorificent Filium sicut honorificant Patrem qui non honorificat Filium non honorificat Patrem qui misit illum
JOHN|5|24|amen amen dico vobis quia qui verbum meum audit et credit ei qui misit me habet vitam aeternam et in iudicium non venit sed transit a morte in vitam
JOHN|5|25|amen amen dico vobis quia venit hora et nunc est quando mortui audient vocem Filii Dei et qui audierint vivent
JOHN|5|26|sicut enim Pater habet vitam in semet ipso sic dedit et Filio vitam habere in semet ipso
JOHN|5|27|et potestatem dedit ei et iudicium facere quia Filius hominis est
JOHN|5|28|nolite mirari hoc quia venit hora in qua omnes qui in monumentis sunt audient vocem eius
JOHN|5|29|et procedent qui bona fecerunt in resurrectionem vitae qui vero mala egerunt in resurrectionem iudicii
JOHN|5|30|non possum ego a me ipso facere quicquam sicut audio iudico et iudicium meum iustum est quia non quaero voluntatem meam sed voluntatem eius qui misit me
JOHN|5|31|si ego testimonium perhibeo de me testimonium meum non est verum
JOHN|5|32|alius est qui testimonium perhibet de me et scio quia verum est testimonium quod perhibet de me
JOHN|5|33|vos misistis ad Iohannem et testimonium perhibuit veritati
JOHN|5|34|ego autem non ab homine testimonium accipio sed haec dico ut vos salvi sitis
JOHN|5|35|ille erat lucerna ardens et lucens vos autem voluistis exultare ad horam in luce eius
JOHN|5|36|ego autem habeo testimonium maius Iohanne opera enim quae dedit mihi Pater ut perficiam ea ipsa opera quae ego facio testimonium perhibent de me quia Pater me misit
JOHN|5|37|et qui misit me Pater ipse testimonium perhibuit de me neque vocem eius umquam audistis neque speciem eius vidistis
JOHN|5|38|et verbum eius non habetis in vobis manens quia quem misit ille huic vos non creditis
JOHN|5|39|scrutamini scripturas quia vos putatis in ipsis vitam aeternam habere et illae sunt quae testimonium perhibent de me
JOHN|5|40|et non vultis venire ad me ut vitam habeatis
JOHN|5|41|claritatem ab hominibus non accipio
JOHN|5|42|sed cognovi vos quia dilectionem Dei non habetis in vobis
JOHN|5|43|ego veni in nomine Patris mei et non accipitis me si alius venerit in nomine suo illum accipietis
JOHN|5|44|quomodo potestis vos credere qui gloriam ab invicem accipitis et gloriam quae a solo est Deo non quaeritis
JOHN|5|45|nolite putare quia ego accusaturus sim vos apud Patrem est qui accuset vos Moses in quo vos speratis
JOHN|5|46|si enim crederetis Mosi crederetis forsitan et mihi de me enim ille scripsit
JOHN|5|47|si autem illius litteris non creditis quomodo meis verbis credetis
JOHN|6|1|post haec abiit Iesus trans mare Galilaeae quod est Tiberiadis
JOHN|6|2|et sequebatur eum multitudo magna quia videbant signa quae faciebat super his qui infirmabantur
JOHN|6|3|subiit ergo in montem Iesus et ibi sedebat cum discipulis suis
JOHN|6|4|erat autem proximum pascha dies festus Iudaeorum
JOHN|6|5|cum sublevasset ergo oculos Iesus et vidisset quia multitudo maxima venit ad eum dicit ad Philippum unde ememus panes ut manducent hii
JOHN|6|6|hoc autem dicebat temptans eum ipse enim sciebat quid esset facturus
JOHN|6|7|respondit ei Philippus ducentorum denariorum panes non sufficiunt eis ut unusquisque modicum quid accipiat
JOHN|6|8|dicit ei unus ex discipulis eius Andreas frater Simonis Petri
JOHN|6|9|est puer unus hic qui habet quinque panes hordiacios et duos pisces sed haec quid sunt inter tantos
JOHN|6|10|dixit ergo Iesus facite homines discumbere erat autem faenum multum in loco discubuerunt ergo viri numero quasi quinque milia
JOHN|6|11|accepit ergo panes Iesus et cum gratias egisset distribuit discumbentibus similiter et ex piscibus quantum volebant
JOHN|6|12|ut autem impleti sunt dixit discipulis suis colligite quae superaverunt fragmenta ne pereant
JOHN|6|13|collegerunt ergo et impleverunt duodecim cofinos fragmentorum ex quinque panibus hordiaciis quae superfuerunt his qui manducaverunt
JOHN|6|14|illi ergo homines cum vidissent quod fecerat signum dicebant quia hic est vere propheta qui venturus est in mundum
JOHN|6|15|Iesus ergo cum cognovisset quia venturi essent ut raperent eum et facerent eum regem fugit iterum in montem ipse solus
JOHN|6|16|ut autem sero factum est descenderunt discipuli eius ad mare
JOHN|6|17|et cum ascendissent navem venerunt trans mare in Capharnaum et tenebrae iam factae erant et non venerat ad eos Iesus
JOHN|6|18|mare autem vento magno flante exsurgebat
JOHN|6|19|cum remigassent ergo quasi stadia viginti quinque aut triginta vident Iesum ambulantem super mare et proximum navi fieri et timuerunt
JOHN|6|20|ille autem dicit eis ego sum nolite timere
JOHN|6|21|voluerunt ergo accipere eum in navi et statim fuit navis ad terram quam ibant
JOHN|6|22|altera die turba quae stabat trans mare vidit quia navicula alia non erat ibi nisi una et quia non introisset cum discipulis suis Iesus in navem sed soli discipuli eius abissent
JOHN|6|23|aliae vero supervenerunt naves a Tiberiade iuxta locum ubi manducaverant panem gratias agente Domino
JOHN|6|24|cum ergo vidisset turba quia Iesus non esset ibi neque discipuli eius ascenderunt naviculas et venerunt Capharnaum quaerentes Iesum
JOHN|6|25|et cum invenissent eum trans mare dixerunt ei rabbi quando huc venisti
JOHN|6|26|respondit eis Iesus et dixit amen amen dico vobis quaeritis me non quia vidistis signa sed quia manducastis ex panibus et saturati estis
JOHN|6|27|operamini non cibum qui perit sed qui permanet in vitam aeternam quem Filius hominis vobis dabit hunc enim Pater signavit Deus
JOHN|6|28|dixerunt ergo ad eum quid faciemus ut operemur opera Dei
JOHN|6|29|respondit Iesus et dixit eis hoc est opus Dei ut credatis in eum quem misit ille
JOHN|6|30|dixerunt ergo ei quod ergo tu facis signum ut videamus et credamus tibi quid operaris
JOHN|6|31|patres nostri manna manducaverunt in deserto sicut scriptum est panem de caelo dedit eis manducare
JOHN|6|32|dixit ergo eis Iesus amen amen dico vobis non Moses dedit vobis panem de caelo sed Pater meus dat vobis panem de caelo verum
JOHN|6|33|panis enim Dei est qui descendit de caelo et dat vitam mundo
JOHN|6|34|dixerunt ergo ad eum Domine semper da nobis panem hunc
JOHN|6|35|dixit autem eis Iesus ego sum panis vitae qui veniet ad me non esuriet et qui credit in me non sitiet umquam
JOHN|6|36|sed dixi vobis quia et vidistis me et non creditis
JOHN|6|37|omne quod dat mihi Pater ad me veniet et eum qui venit ad me non eiciam foras
JOHN|6|38|quia descendi de caelo non ut faciam voluntatem meam sed voluntatem eius qui misit me
JOHN|6|39|haec est autem voluntas eius qui misit me Patris ut omne quod dedit mihi non perdam ex eo sed resuscitem illum novissimo die
JOHN|6|40|haec est enim voluntas Patris mei qui misit me ut omnis qui videt Filium et credit in eum habeat vitam aeternam et resuscitabo ego eum in novissimo die
JOHN|6|41|murmurabant ergo Iudaei de illo quia dixisset ego sum panis qui de caelo descendi
JOHN|6|42|et dicebant nonne hic est Iesus filius Ioseph cuius nos novimus patrem et matrem quomodo ergo dicit hic quia de caelo descendi
JOHN|6|43|respondit ergo Iesus et dixit eis nolite murmurare in invicem
JOHN|6|44|nemo potest venire ad me nisi Pater qui misit me traxerit eum et ego resuscitabo eum novissimo die
JOHN|6|45|est scriptum in prophetis et erunt omnes docibiles Dei omnis qui audivit a Patre et didicit venit ad me
JOHN|6|46|non quia Patrem vidit quisquam nisi is qui est a Deo hic vidit Patrem
JOHN|6|47|amen amen dico vobis qui credit in me habet vitam aeternam
JOHN|6|48|ego sum panis vitae
JOHN|6|49|patres vestri manducaverunt in deserto manna et mortui sunt
JOHN|6|50|hic est panis de caelo descendens ut si quis ex ipso manducaverit non moriatur
JOHN|6|51|ego sum panis vivus qui de caelo descendi
JOHN|6|52|si quis manducaverit ex hoc pane vivet in aeternum et panis quem ego dabo caro mea est pro mundi vita
JOHN|6|53|litigabant ergo Iudaei ad invicem dicentes quomodo potest hic nobis carnem suam dare ad manducandum
JOHN|6|54|dixit ergo eis Iesus amen amen dico vobis nisi manducaveritis carnem Filii hominis et biberitis eius sanguinem non habetis vitam in vobis
JOHN|6|55|qui manducat meam carnem et bibit meum sanguinem habet vitam aeternam et ego resuscitabo eum in novissimo die
JOHN|6|56|caro enim mea vere est cibus et sanguis meus vere est potus
JOHN|6|57|qui manducat meam carnem et bibit meum sanguinem in me manet et ego in illo
JOHN|6|58|sicut misit me vivens Pater et ego vivo propter Patrem et qui manducat me et ipse vivet propter me
JOHN|6|59|hic est panis qui de caelo descendit non sicut manducaverunt patres vestri manna et mortui sunt qui manducat hunc panem vivet in aeternum
JOHN|6|60|haec dixit in synagoga docens in Capharnaum
JOHN|6|61|multi ergo audientes ex discipulis eius dixerunt durus est hic sermo quis potest eum audire
JOHN|6|62|sciens autem Iesus apud semet ipsum quia murmurarent de hoc discipuli eius dixit eis hoc vos scandalizat
JOHN|6|63|si ergo videritis Filium hominis ascendentem ubi erat prius
JOHN|6|64|spiritus est qui vivificat caro non prodest quicquam verba quae ego locutus sum vobis spiritus et vita sunt
JOHN|6|65|sed sunt quidam ex vobis qui non credunt sciebat enim ab initio Iesus qui essent credentes et quis traditurus esset eum
JOHN|6|66|et dicebat propterea dixi vobis quia nemo potest venire ad me nisi fuerit ei datum a Patre meo
JOHN|6|67|ex hoc multi discipulorum eius abierunt retro et iam non cum illo ambulabant
JOHN|6|68|dixit ergo Iesus ad duodecim numquid et vos vultis abire
JOHN|6|69|respondit ergo ei Simon Petrus Domine ad quem ibimus verba vitae aeternae habes
JOHN|6|70|et nos credidimus et cognovimus quia tu es Christus Filius Dei
JOHN|6|71|respondit eis Iesus nonne ego vos duodecim elegi et ex vobis unus diabolus est
JOHN|6|72|dicebat autem Iudam Simonis Scariotis hic enim erat traditurus eum cum esset unus ex duodecim
JOHN|7|1|post haec ambulabat Iesus in Galilaeam non enim volebat in Iudaeam ambulare quia quaerebant eum Iudaei interficere
JOHN|7|2|erat autem in proximo dies festus Iudaeorum scenopegia
JOHN|7|3|dixerunt autem ad eum fratres eius transi hinc et vade in Iudaeam ut et discipuli tui videant opera tua quae facis
JOHN|7|4|nemo quippe in occulto quid facit et quaerit ipse in palam esse si haec facis manifesta te ipsum mundo
JOHN|7|5|neque enim fratres eius credebant in eum
JOHN|7|6|dicit ergo eis Iesus tempus meum nondum advenit tempus autem vestrum semper est paratum
JOHN|7|7|non potest mundus odisse vos me autem odit quia ego testimonium perhibeo de illo quia opera eius mala sunt
JOHN|7|8|vos ascendite ad diem festum hunc ego non ascendo ad diem festum istum quia meum tempus nondum impletum est
JOHN|7|9|haec cum dixisset ipse mansit in Galilaea
JOHN|7|10|ut autem ascenderunt fratres eius tunc et ipse ascendit ad diem festum non manifeste sed quasi in occulto
JOHN|7|11|Iudaei ergo quaerebant eum in die festo et dicebant ubi est ille
JOHN|7|12|et murmur multus de eo erat in turba; quidam enim dicebant quia bonus est alii autem dicebant non sed seducit turbas
JOHN|7|13|nemo tamen palam loquebatur de illo propter metum Iudaeorum
JOHN|7|14|iam autem die festo mediante ascendit Iesus in templum et docebat
JOHN|7|15|et mirabantur Iudaei dicentes quomodo hic litteras scit cum non didicerit
JOHN|7|16|respondit eis Iesus et dixit mea doctrina non est mea sed eius qui misit me
JOHN|7|17|si quis voluerit voluntatem eius facere cognoscet de doctrina utrum ex Deo sit an ego a me ipso loquar
JOHN|7|18|qui a semet ipso loquitur gloriam propriam quaerit qui autem quaerit gloriam eius qui misit illum hic verax est et iniustitia in illo non est
JOHN|7|19|nonne Moses dedit vobis legem et nemo ex vobis facit legem
JOHN|7|20|quid me quaeritis interficere respondit turba et dixit daemonium habes quis te quaerit interficere
JOHN|7|21|respondit Iesus et dixit eis unum opus feci et omnes miramini
JOHN|7|22|propterea Moses dedit vobis circumcisionem non quia ex Mose est sed ex patribus et in sabbato circumciditis hominem
JOHN|7|23|si circumcisionem accipit homo in sabbato ut non solvatur lex Mosi mihi indignamini quia totum hominem sanum feci in sabbato
JOHN|7|24|nolite iudicare secundum faciem sed iustum iudicium iudicate
JOHN|7|25|dicebant ergo quidam ex Hierosolymis nonne hic est quem quaerunt interficere
JOHN|7|26|et ecce palam loquitur et nihil ei dicunt numquid vere cognoverunt principes quia hic est Christus
JOHN|7|27|sed hunc scimus unde sit Christus autem cum venerit nemo scit unde sit
JOHN|7|28|clamabat ergo docens in templo Iesus et dicens et me scitis et unde sim scitis et a me ipso non veni sed est verus qui misit me quem vos non scitis
JOHN|7|29|ego scio eum quia ab ipso sum et ipse me misit
JOHN|7|30|quaerebant ergo eum adprehendere et nemo misit in illum manus quia nondum venerat hora eius
JOHN|7|31|de turba autem multi crediderunt in eum et dicebant Christus cum venerit numquid plura signa faciet quam quae hic facit
JOHN|7|32|audierunt Pharisaei turbam murmurantem de illo haec et miserunt principes et Pharisaei ministros ut adprehenderent eum
JOHN|7|33|dixit ergo Iesus adhuc modicum tempus vobiscum sum et vado ad eum qui misit me
JOHN|7|34|quaeretis me et non invenietis et ubi sum ego vos non potestis venire
JOHN|7|35|dixerunt ergo Iudaei ad se ipsos quo hic iturus est quia non inveniemus eum numquid in dispersionem gentium iturus est et docturus gentes
JOHN|7|36|quis est hic sermo quem dixit quaeretis me et non invenietis et ubi sum ego non potestis venire
JOHN|7|37|in novissimo autem die magno festivitatis stabat Iesus et clamabat dicens si quis sitit veniat ad me et bibat
JOHN|7|38|qui credit in me sicut dixit scriptura flumina de ventre eius fluent aquae vivae
JOHN|7|39|hoc autem dixit de Spiritu quem accepturi erant credentes in eum non enim erat Spiritus quia Iesus nondum fuerat glorificatus
JOHN|7|40|ex illa ergo turba cum audissent hos sermones eius dicebant hic est vere propheta
JOHN|7|41|alii dicebant hic est Christus quidam autem dicebant numquid a Galilaea Christus venit
JOHN|7|42|nonne scriptura dicit quia ex semine David et Bethleem castello ubi erat David venit Christus
JOHN|7|43|dissensio itaque facta est in turba propter eum
JOHN|7|44|quidam autem ex ipsis volebant adprehendere eum sed nemo misit super illum manus
JOHN|7|45|venerunt ergo ministri ad pontifices et Pharisaeos et dixerunt eis illi quare non adduxistis eum
JOHN|7|46|responderunt ministri numquam sic locutus est homo sicut hic homo
JOHN|7|47|responderunt ergo eis Pharisaei numquid et vos seducti estis
JOHN|7|48|numquid aliquis ex principibus credidit in eum aut ex Pharisaeis
JOHN|7|49|sed turba haec quae non novit legem maledicti sunt
JOHN|7|50|dicit Nicodemus ad eos ille qui venit ad eum nocte qui unus erat ex ipsis
JOHN|7|51|numquid lex nostra iudicat hominem nisi audierit ab ipso prius et cognoverit quid faciat
JOHN|7|52|responderunt et dixerunt ei numquid et tu Galilaeus es scrutare et vide quia propheta a Galilaea non surgit
JOHN|7|53|et reversi sunt unusquisque in domum suam
JOHN|8|1|Iesus autem perrexit in montem Oliveti
JOHN|8|2|et diluculo iterum venit in templum et omnis populus venit ad eum et sedens docebat eos
JOHN|8|3|adducunt autem scribae et Pharisaei mulierem in adulterio deprehensam et statuerunt eam in medio
JOHN|8|4|et dixerunt ei magister haec mulier modo deprehensa est in adulterio
JOHN|8|5|in lege autem Moses mandavit nobis huiusmodi lapidare tu ergo quid dicis
JOHN|8|6|haec autem dicebant temptantes eum ut possent accusare eum Iesus autem inclinans se deorsum digito scribebat in terra
JOHN|8|7|cum autem perseverarent interrogantes eum erexit se et dixit eis qui sine peccato est vestrum primus in illam lapidem mittat
JOHN|8|8|et iterum se inclinans scribebat in terra
JOHN|8|9|audientes autem unus post unum exiebant incipientes a senioribus et remansit solus et mulier in medio stans
JOHN|8|10|erigens autem se Iesus dixit ei mulier ubi sunt nemo te condemnavit
JOHN|8|11|quae dixit nemo Domine dixit autem Iesus nec ego te condemnabo vade et amplius iam noli peccare
JOHN|8|12|iterum ergo locutus est eis Iesus dicens ego sum lux mundi qui sequitur me non ambulabit in tenebris sed habebit lucem vitae
JOHN|8|13|dixerunt ergo ei Pharisaei tu de te ipso testimonium perhibes testimonium tuum non est verum
JOHN|8|14|respondit Iesus et dixit eis et si ego testimonium perhibeo de me ipso verum est testimonium meum quia scio unde veni et quo vado vos autem nescitis unde venio aut quo vado
JOHN|8|15|vos secundum carnem iudicatis ego non iudico quemquam
JOHN|8|16|et si iudico ego iudicium meum verum est quia solus non sum sed ego et qui me misit Pater
JOHN|8|17|et in lege vestra scriptum est quia duorum hominum testimonium verum est
JOHN|8|18|ego sum qui testimonium perhibeo de me ipso et testimonium perhibet de me qui misit me Pater
JOHN|8|19|dicebant ergo ei ubi est Pater tuus respondit Iesus neque me scitis neque Patrem meum si me sciretis forsitan et Patrem meum sciretis
JOHN|8|20|haec verba locutus est in gazofilacio docens in templo et nemo adprehendit eum quia necdum venerat hora eius
JOHN|8|21|dixit ergo iterum eis Iesus ego vado et quaeretis me et in peccato vestro moriemini quo ego vado vos non potestis venire
JOHN|8|22|dicebant ergo Iudaei numquid interficiet semet ipsum quia dicit quo ego vado vos non potestis venire
JOHN|8|23|et dicebat eis vos de deorsum estis ego de supernis sum vos de mundo hoc estis ego non sum de hoc mundo
JOHN|8|24|dixi ergo vobis quia moriemini in peccatis vestris si enim non credideritis quia ego sum moriemini in peccato vestro
JOHN|8|25|dicebant ergo ei tu quis es dixit eis Iesus principium quia et loquor vobis
JOHN|8|26|multa habeo de vobis loqui et iudicare sed qui misit me verax est et ego quae audivi ab eo haec loquor in mundo
JOHN|8|27|et non cognoverunt quia Patrem eis dicebat
JOHN|8|28|dixit ergo eis Iesus cum exaltaveritis Filium hominis tunc cognoscetis quia ego sum et a me ipso facio nihil sed sicut docuit me Pater haec loquor
JOHN|8|29|et qui me misit mecum est non reliquit me solum quia ego quae placita sunt ei facio semper
JOHN|8|30|haec illo loquente multi crediderunt in eum
JOHN|8|31|dicebat ergo Iesus ad eos qui crediderunt ei Iudaeos si vos manseritis in sermone meo vere discipuli mei eritis
JOHN|8|32|et cognoscetis veritatem et veritas liberabit vos
JOHN|8|33|responderunt ei semen Abrahae sumus et nemini servivimus umquam quomodo tu dicis liberi eritis
JOHN|8|34|respondit eis Iesus amen amen dico vobis quia omnis qui facit peccatum servus est peccati
JOHN|8|35|servus autem non manet in domo in aeternum filius manet in aeternum
JOHN|8|36|si ergo Filius vos liberaverit vere liberi eritis
JOHN|8|37|scio quia filii Abrahae estis sed quaeritis me interficere quia sermo meus non capit in vobis
JOHN|8|38|ego quod vidi apud Patrem loquor et vos quae vidistis apud patrem vestrum facitis
JOHN|8|39|responderunt et dixerunt ei pater noster Abraham est dicit eis Iesus si filii Abrahae estis opera Abrahae facite
JOHN|8|40|nunc autem quaeritis me interficere hominem qui veritatem vobis locutus sum quam audivi a Deo hoc Abraham non fecit
JOHN|8|41|vos facitis opera patris vestri dixerunt itaque ei nos ex fornicatione non sumus nati unum patrem habemus Deum
JOHN|8|42|dixit ergo eis Iesus si Deus pater vester esset diligeretis utique me ego enim ex Deo processi et veni neque enim a me ipso veni sed ille me misit
JOHN|8|43|quare loquellam meam non cognoscitis quia non potestis audire sermonem meum
JOHN|8|44|vos ex patre diabolo estis et desideria patris vestri vultis facere ille homicida erat ab initio et in veritate non stetit quia non est veritas in eo cum loquitur mendacium ex propriis loquitur quia mendax est et pater eius
JOHN|8|45|ego autem quia veritatem dico non creditis mihi
JOHN|8|46|quis ex vobis arguit me de peccato si veritatem dico quare vos non creditis mihi
JOHN|8|47|qui est ex Deo verba Dei audit propterea vos non auditis quia ex Deo non estis
JOHN|8|48|responderunt igitur Iudaei et dixerunt ei nonne bene dicimus nos quia Samaritanus es tu et daemonium habes
JOHN|8|49|respondit Iesus ego daemonium non habeo sed honorifico Patrem meum et vos inhonoratis me
JOHN|8|50|ego autem non quaero gloriam meam est qui quaerit et iudicat
JOHN|8|51|amen amen dico vobis si quis sermonem meum servaverit mortem non videbit in aeternum
JOHN|8|52|dixerunt ergo Iudaei nunc cognovimus quia daemonium habes Abraham mortuus est et prophetae et tu dicis si quis sermonem meum servaverit non gustabit mortem in aeternum
JOHN|8|53|numquid tu maior es patre nostro Abraham qui mortuus est et prophetae mortui sunt quem te ipsum facis
JOHN|8|54|respondit Iesus si ego glorifico me ipsum gloria mea nihil est est Pater meus qui glorificat me quem vos dicitis quia Deus noster est
JOHN|8|55|et non cognovistis eum ego autem novi eum et si dixero quia non scio eum ero similis vobis mendax sed scio eum et sermonem eius servo
JOHN|8|56|Abraham pater vester exultavit ut videret diem meum et vidit et gavisus est
JOHN|8|57|dixerunt ergo Iudaei ad eum quinquaginta annos nondum habes et Abraham vidisti
JOHN|8|58|dixit eis Iesus amen amen dico vobis antequam Abraham fieret ego sum
JOHN|8|59|tulerunt ergo lapides ut iacerent in eum Iesus autem abscondit se et exivit de templo
JOHN|9|1|et praeteriens vidit hominem caecum a nativitate
JOHN|9|2|et interrogaverunt eum discipuli sui rabbi quis peccavit hic aut parentes eius ut caecus nasceretur
JOHN|9|3|respondit Iesus neque hic peccavit neque parentes eius sed ut manifestetur opera Dei in illo
JOHN|9|4|me oportet operari opera eius qui misit me donec dies est venit nox quando nemo potest operari
JOHN|9|5|quamdiu in mundo sum lux sum mundi
JOHN|9|6|haec cum dixisset expuit in terram et fecit lutum ex sputo et linuit lutum super oculos eius
JOHN|9|7|et dixit ei vade lava in natatoria Siloae quod interpretatur Missus abiit ergo et lavit et venit videns
JOHN|9|8|itaque vicini et qui videbant eum prius quia mendicus erat dicebant nonne hic est qui sedebat et mendicabat alii dicebant quia hic est
JOHN|9|9|alii autem nequaquam sed similis est eius ille dicebat quia ego sum
JOHN|9|10|dicebant ergo ei quomodo aperti sunt oculi tibi
JOHN|9|11|respondit ille homo qui dicitur Iesus lutum fecit et unxit oculos meos et dixit mihi vade ad natatoriam Siloae et lava et abii et lavi et vidi
JOHN|9|12|dixerunt ei ubi est ille ait nescio
JOHN|9|13|adducunt eum ad Pharisaeos qui caecus fuerat
JOHN|9|14|erat autem sabbatum quando lutum fecit Iesus et aperuit oculos eius
JOHN|9|15|iterum ergo interrogabant eum Pharisaei quomodo vidisset ille autem dixit eis lutum posuit mihi super oculos et lavi et video
JOHN|9|16|dicebant ergo ex Pharisaeis quidam non est hic homo a Deo quia sabbatum non custodit alii dicebant quomodo potest homo peccator haec signa facere et scisma erat in eis
JOHN|9|17|dicunt ergo caeco iterum tu quid dicis de eo qui aperuit oculos tuos ille autem dixit quia propheta est
JOHN|9|18|non crediderunt ergo Iudaei de illo quia caecus fuisset et vidisset donec vocaverunt parentes eius qui viderat
JOHN|9|19|et interrogaverunt eos dicentes hic est filius vester quem vos dicitis quia caecus natus est quomodo ergo nunc videt
JOHN|9|20|responderunt eis parentes eius et dixerunt scimus quia hic est filius noster et quia caecus natus est
JOHN|9|21|quomodo autem nunc videat nescimus aut quis eius aperuit oculos nos nescimus ipsum interrogate aetatem habet ipse de se loquatur
JOHN|9|22|haec dixerunt parentes eius quia timebant Iudaeos iam enim conspiraverant Iudaei ut si quis eum confiteretur Christum extra synagogam fieret
JOHN|9|23|propterea parentes eius dixerunt quia aetatem habet ipsum interrogate
JOHN|9|24|vocaverunt ergo rursum hominem qui fuerat caecus et dixerunt ei da gloriam Deo nos scimus quia hic homo peccator est
JOHN|9|25|dixit ergo ille si peccator est nescio unum scio quia caecus cum essem modo video
JOHN|9|26|dixerunt ergo illi quid fecit tibi quomodo aperuit tibi oculos
JOHN|9|27|respondit eis dixi vobis iam et audistis quid iterum vultis audire numquid et vos vultis discipuli eius fieri
JOHN|9|28|maledixerunt ei et dixerunt tu discipulus illius es nos autem Mosi discipuli sumus
JOHN|9|29|nos scimus quia Mosi locutus est Deus hunc autem nescimus unde sit
JOHN|9|30|respondit ille homo et dixit eis in hoc enim mirabile est quia vos nescitis unde sit et aperuit meos oculos
JOHN|9|31|scimus autem quia peccatores Deus non audit sed si quis Dei cultor est et voluntatem eius facit hunc exaudit
JOHN|9|32|a saeculo non est auditum quia aperuit quis oculos caeci nati
JOHN|9|33|nisi esset hic a Deo non poterat facere quicquam
JOHN|9|34|responderunt et dixerunt ei in peccatis natus es totus et tu doces nos et eiecerunt eum foras
JOHN|9|35|audivit Iesus quia eiecerunt eum foras et cum invenisset eum dixit ei tu credis in Filium Dei
JOHN|9|36|respondit ille et dixit quis est Domine ut credam in eum
JOHN|9|37|et dixit ei Iesus et vidisti eum et qui loquitur tecum ipse est
JOHN|9|38|at ille ait credo Domine et procidens adoravit eum
JOHN|9|39|dixit ei Iesus in iudicium ego in hunc mundum veni ut qui non vident videant et qui vident caeci fiant
JOHN|9|40|et audierunt ex Pharisaeis qui cum ipso erant et dixerunt ei numquid et nos caeci sumus
JOHN|9|41|dixit eis Iesus si caeci essetis non haberetis peccatum nunc vero dicitis quia videmus peccatum vestrum manet
JOHN|10|1|amen amen dico vobis qui non intrat per ostium in ovile ovium sed ascendit aliunde ille fur est et latro
JOHN|10|2|qui autem intrat per ostium pastor est ovium
JOHN|10|3|huic ostiarius aperit et oves vocem eius audiunt et proprias oves vocat nominatim et educit eas
JOHN|10|4|et cum proprias oves emiserit ante eas vadit et oves illum sequuntur quia sciunt vocem eius
JOHN|10|5|alienum autem non sequuntur sed fugient ab eo quia non noverunt vocem alienorum
JOHN|10|6|hoc proverbium dixit eis Iesus illi autem non cognoverunt quid loqueretur eis
JOHN|10|7|dixit ergo eis iterum Iesus amen amen dico vobis quia ego sum ostium ovium
JOHN|10|8|omnes quotquot venerunt fures sunt et latrones sed non audierunt eos oves
JOHN|10|9|ego sum ostium per me si quis introierit salvabitur et ingredietur et egredietur et pascua inveniet
JOHN|10|10|fur non venit nisi ut furetur et mactet et perdat ego veni ut vitam habeant et abundantius habeant
JOHN|10|11|ego sum pastor bonus bonus pastor animam suam dat pro ovibus
JOHN|10|12|mercennarius et qui non est pastor cuius non sunt oves propriae videt lupum venientem et dimittit oves et fugit et lupus rapit et dispergit oves
JOHN|10|13|mercennarius autem fugit quia mercennarius est et non pertinet ad eum de ovibus
JOHN|10|14|ego sum pastor bonus et cognosco meas et cognoscunt me meae
JOHN|10|15|sicut novit me Pater et ego agnosco Patrem et animam meam pono pro ovibus
JOHN|10|16|et alias oves habeo quae non sunt ex hoc ovili et illas oportet me adducere et vocem meam audient et fiet unum ovile unus pastor
JOHN|10|17|propterea me Pater diligit quia ego pono animam meam ut iterum sumam eam
JOHN|10|18|nemo tollit eam a me sed ego pono eam a me ipso potestatem habeo ponendi eam et potestatem habeo iterum sumendi eam hoc mandatum accepi a Patre meo
JOHN|10|19|dissensio iterum facta est inter Iudaeos propter sermones hos
JOHN|10|20|dicebant autem multi ex ipsis daemonium habet et insanit quid eum auditis
JOHN|10|21|alii dicebant haec verba non sunt daemonium habentis numquid daemonium potest caecorum oculos aperire
JOHN|10|22|facta sunt autem encenia in Hierosolymis et hiemps erat
JOHN|10|23|et ambulabat Iesus in templo in porticu Salomonis
JOHN|10|24|circumdederunt ergo eum Iudaei et dicebant ei quousque animam nostram tollis si tu es Christus dic nobis palam
JOHN|10|25|respondit eis Iesus loquor vobis et non creditis opera quae ego facio in nomine Patris mei haec testimonium perhibent de me
JOHN|10|26|sed vos non creditis quia non estis ex ovibus meis
JOHN|10|27|oves meae vocem meam audiunt et ego cognosco eas et sequuntur me
JOHN|10|28|et ego vitam aeternam do eis et non peribunt in aeternum et non rapiet eas quisquam de manu mea
JOHN|10|29|Pater meus quod dedit mihi maius omnibus est et nemo potest rapere de manu Patris mei
JOHN|10|30|ego et Pater unum sumus
JOHN|10|31|sustulerunt lapides Iudaei ut lapidarent eum
JOHN|10|32|respondit eis Iesus multa opera bona ostendi vobis ex Patre meo propter quod eorum opus me lapidatis
JOHN|10|33|responderunt ei Iudaei de bono opere non lapidamus te sed de blasphemia et quia tu homo cum sis facis te ipsum Deum
JOHN|10|34|respondit eis Iesus nonne scriptum est in lege vestra quia ego dixi dii estis
JOHN|10|35|si illos dixit deos ad quos sermo Dei factus est et non potest solvi scriptura
JOHN|10|36|quem Pater sanctificavit et misit in mundum vos dicitis quia blasphemas quia dixi Filius Dei sum
JOHN|10|37|si non facio opera Patris mei nolite credere mihi
JOHN|10|38|si autem facio et si mihi non vultis credere operibus credite ut cognoscatis et credatis quia in me est Pater et ego in Patre
JOHN|10|39|quaerebant ergo eum prendere et exivit de manibus eorum
JOHN|10|40|et abiit iterum trans Iordanen in eum locum ubi erat Iohannes baptizans primum et mansit illic
JOHN|10|41|et multi venerunt ad eum et dicebant quia Iohannes quidem signum fecit nullum
JOHN|10|42|omnia autem quaecumque dixit Iohannes de hoc vera erant et multi crediderunt in eum
JOHN|11|1|erat autem quidam languens Lazarus a Bethania de castello Mariae et Marthae sororis eius
JOHN|11|2|Maria autem erat quae unxit Dominum unguento et extersit pedes eius capillis suis cuius frater Lazarus infirmabatur
JOHN|11|3|miserunt ergo sorores ad eum dicentes Domine ecce quem amas infirmatur
JOHN|11|4|audiens autem Iesus dixit eis infirmitas haec non est ad mortem sed pro gloria Dei ut glorificetur Filius Dei per eam
JOHN|11|5|diligebat autem Iesus Martham et sororem eius Mariam et Lazarum
JOHN|11|6|ut ergo audivit quia infirmabatur tunc quidem mansit in eodem loco duobus diebus
JOHN|11|7|deinde post haec dicit discipulis suis eamus in Iudaeam iterum
JOHN|11|8|dicunt ei discipuli rabbi nunc quaerebant te Iudaei lapidare et iterum vadis illuc
JOHN|11|9|respondit Iesus nonne duodecim horae sunt diei si quis ambulaverit in die non offendit quia lucem huius mundi videt
JOHN|11|10|si autem ambulaverit nocte offendit quia lux non est in eo
JOHN|11|11|haec ait et post hoc dicit eis Lazarus amicus noster dormit sed vado ut a somno exsuscitem eum
JOHN|11|12|dixerunt ergo discipuli eius Domine si dormit salvus erit
JOHN|11|13|dixerat autem Iesus de morte eius illi autem putaverunt quia de dormitione somni diceret
JOHN|11|14|tunc ergo dixit eis Iesus manifeste Lazarus mortuus est
JOHN|11|15|et gaudeo propter vos ut credatis quoniam non eram ibi sed eamus ad eum
JOHN|11|16|dixit ergo Thomas qui dicitur Didymus ad condiscipulos eamus et nos ut moriamur cum eo
JOHN|11|17|venit itaque Iesus et invenit eum quattuor dies iam in monumento habentem
JOHN|11|18|erat autem Bethania iuxta Hierosolyma quasi stadiis quindecim
JOHN|11|19|multi autem ex Iudaeis venerant ad Martham et Mariam ut consolarentur eas de fratre suo
JOHN|11|20|Martha ergo ut audivit quia Iesus venit occurrit illi Maria autem domi sedebat
JOHN|11|21|dixit ergo Martha ad Iesum Domine si fuisses hic frater meus non fuisset mortuus
JOHN|11|22|sed et nunc scio quia quaecumque poposceris a Deo dabit tibi Deus
JOHN|11|23|dicit illi Iesus resurget frater tuus
JOHN|11|24|dicit ei Martha scio quia resurget in resurrectione in novissima die
JOHN|11|25|dixit ei Iesus ego sum resurrectio et vita qui credit in me et si mortuus fuerit vivet
JOHN|11|26|et omnis qui vivit et credit in me non morietur in aeternum credis hoc
JOHN|11|27|ait illi utique Domine ego credidi quia tu es Christus Filius Dei qui in mundum venisti
JOHN|11|28|et cum haec dixisset abiit et vocavit Mariam sororem suam silentio dicens magister adest et vocat te
JOHN|11|29|illa ut audivit surgit cito et venit ad eum
JOHN|11|30|nondum enim venerat Iesus in castellum sed erat adhuc in illo loco ubi occurrerat ei Martha
JOHN|11|31|Iudaei igitur qui erant cum ea in domo et consolabantur eam cum vidissent Mariam quia cito surrexit et exiit secuti sunt eam dicentes quia vadit ad monumentum ut ploret ibi
JOHN|11|32|Maria ergo cum venisset ubi erat Iesus videns eum cecidit ad pedes eius et dixit ei Domine si fuisses hic non esset mortuus frater meus
JOHN|11|33|Iesus ergo ut vidit eam plorantem et Iudaeos qui venerant cum ea plorantes fremuit spiritu et turbavit se ipsum
JOHN|11|34|et dixit ubi posuistis eum dicunt ei Domine veni et vide
JOHN|11|35|et lacrimatus est Iesus
JOHN|11|36|dixerunt ergo Iudaei ecce quomodo amabat eum
JOHN|11|37|quidam autem dixerunt ex ipsis non poterat hic qui aperuit oculos caeci facere ut et hic non moreretur
JOHN|11|38|Iesus ergo rursum fremens in semet ipso venit ad monumentum erat autem spelunca et lapis superpositus erat ei
JOHN|11|39|ait Iesus tollite lapidem dicit ei Martha soror eius qui mortuus fuerat Domine iam fetet quadriduanus enim est
JOHN|11|40|dicit ei Iesus nonne dixi tibi quoniam si credideris videbis gloriam Dei
JOHN|11|41|tulerunt ergo lapidem Iesus autem elevatis sursum oculis dixit Pater gratias ago tibi quoniam audisti me
JOHN|11|42|ego autem sciebam quia semper me audis sed propter populum qui circumstat dixi ut credant quia tu me misisti
JOHN|11|43|haec cum dixisset voce magna clamavit Lazare veni foras
JOHN|11|44|et statim prodiit qui fuerat mortuus ligatus pedes et manus institis et facies illius sudario erat ligata dicit Iesus eis solvite eum et sinite abire
JOHN|11|45|multi ergo ex Iudaeis qui venerant ad Mariam et viderant quae fecit crediderunt in eum
JOHN|11|46|quidam autem ex ipsis abierunt ad Pharisaeos et dixerunt eis quae fecit Iesus
JOHN|11|47|collegerunt ergo pontifices et Pharisaei concilium et dicebant quid facimus quia hic homo multa signa facit
JOHN|11|48|si dimittimus eum sic omnes credent in eum et venient Romani et tollent nostrum et locum et gentem
JOHN|11|49|unus autem ex ipsis Caiaphas cum esset pontifex anni illius dixit eis vos nescitis quicquam
JOHN|11|50|nec cogitatis quia expedit nobis ut unus moriatur homo pro populo et non tota gens pereat
JOHN|11|51|hoc autem a semet ipso non dixit sed cum esset pontifex anni illius prophetavit quia Iesus moriturus erat pro gente
JOHN|11|52|et non tantum pro gente sed et ut filios Dei qui erant dispersi congregaret in unum
JOHN|11|53|ab illo ergo die cogitaverunt ut interficerent eum
JOHN|11|54|Iesus ergo iam non in palam ambulabat apud Iudaeos sed abiit in regionem iuxta desertum in civitatem quae dicitur Efrem et ibi morabatur cum discipulis
JOHN|11|55|proximum autem erat pascha Iudaeorum et ascenderunt multi Hierosolyma de regione ante pascha ut sanctificarent se ipsos
JOHN|11|56|quaerebant ergo Iesum et conloquebantur ad invicem in templo stantes quid putatis quia non veniat ad diem festum
JOHN|11|57|dederant autem pontifices et Pharisaei mandatum ut si quis cognoverit ubi sit indicet ut adprehendant eum
JOHN|12|1|Iesus ergo ante sex dies paschae venit Bethaniam ubi fuerat Lazarus mortuus quem suscitavit Iesus
JOHN|12|2|fecerunt autem ei cenam ibi et Martha ministrabat Lazarus vero unus erat ex discumbentibus cum eo
JOHN|12|3|Maria ergo accepit libram unguenti nardi pistici pretiosi unxit pedes Iesu et extersit capillis suis pedes eius et domus impleta est ex odore unguenti
JOHN|12|4|dicit ergo unus ex discipulis eius Iudas Scariotis qui erat eum traditurus
JOHN|12|5|quare hoc unguentum non veniit trecentis denariis et datum est egenis
JOHN|12|6|dixit autem hoc non quia de egenis pertinebat ad eum sed quia fur erat et loculos habens ea quae mittebantur portabat
JOHN|12|7|dixit ergo Iesus sine illam ut in die sepulturae meae servet illud
JOHN|12|8|pauperes enim semper habetis vobiscum me autem non semper habetis
JOHN|12|9|cognovit ergo turba multa ex Iudaeis quia illic est et venerunt non propter Iesum tantum sed ut Lazarum viderent quem suscitavit a mortuis
JOHN|12|10|cogitaverunt autem principes sacerdotum ut et Lazarum interficerent
JOHN|12|11|quia multi propter illum abibant ex Iudaeis et credebant in Iesum
JOHN|12|12|in crastinum autem turba multa quae venerat ad diem festum cum audissent quia venit Iesus Hierosolyma
JOHN|12|13|acceperunt ramos palmarum et processerunt obviam ei et clamabant osanna benedictus qui venit in nomine Domini rex Israhel
JOHN|12|14|et invenit Iesus asellum et sedit super eum sicut scriptum est
JOHN|12|15|noli timere filia Sion ecce rex tuus venit sedens super pullum asinae
JOHN|12|16|haec non cognoverunt discipuli eius primum sed quando glorificatus est Iesus tunc recordati sunt quia haec erant scripta de eo et haec fecerunt ei
JOHN|12|17|testimonium ergo perhibebat turba quae erat cum eo quando Lazarum vocavit de monumento et suscitavit eum a mortuis
JOHN|12|18|propterea et obviam venit ei turba quia audierunt eum fecisse hoc signum
JOHN|12|19|Pharisaei ergo dixerunt ad semet ipsos videtis quia nihil proficimus ecce mundus totus post eum abiit
JOHN|12|20|erant autem gentiles quidam ex his qui ascenderant ut adorarent in die festo
JOHN|12|21|hii ergo accesserunt ad Philippum qui erat a Bethsaida Galilaeae et rogabant eum dicentes domine volumus Iesum videre
JOHN|12|22|venit Philippus et dicit Andreae Andreas rursum et Philippus dixerunt Iesu
JOHN|12|23|Iesus autem respondit eis dicens venit hora ut clarificetur Filius hominis
JOHN|12|24|amen amen dico vobis nisi granum frumenti cadens in terram mortuum fuerit
JOHN|12|25|ipsum solum manet si autem mortuum fuerit multum fructum adfert qui amat animam suam perdet eam et qui odit animam suam in hoc mundo in vitam aeternam custodit eam
JOHN|12|26|si quis mihi ministrat me sequatur et ubi sum ego illic et minister meus erit si quis mihi ministraverit honorificabit eum Pater meus
JOHN|12|27|nunc anima mea turbata est et quid dicam Pater salvifica me ex hora hac sed propterea veni in horam hanc
JOHN|12|28|Pater clarifica tuum nomen venit ergo vox de caelo et clarificavi et iterum clarificabo
JOHN|12|29|turba ergo quae stabat et audierat dicebant tonitruum factum esse alii dicebant angelus ei locutus est
JOHN|12|30|respondit Iesus et dixit non propter me vox haec venit sed propter vos
JOHN|12|31|nunc iudicium est mundi nunc princeps huius mundi eicietur foras
JOHN|12|32|et ego si exaltatus fuero a terra omnia traham ad me ipsum
JOHN|12|33|hoc autem dicebat significans qua morte esset moriturus
JOHN|12|34|respondit ei turba nos audivimus ex lege quia Christus manet in aeternum et quomodo tu dicis oportet exaltari Filium hominis quis est iste Filius hominis
JOHN|12|35|dixit ergo eis Iesus adhuc modicum lumen in vobis est ambulate dum lucem habetis ut non tenebrae vos conprehendant et qui ambulat in tenebris nescit quo vadat
JOHN|12|36|dum lucem habetis credite in lucem ut filii lucis sitis haec locutus est Iesus et abiit et abscondit se ab eis
JOHN|12|37|cum autem tanta signa fecisset coram eis non credebant in eum
JOHN|12|38|ut sermo Esaiae prophetae impleretur quem dixit Domine quis credidit auditui nostro et brachium Domini cui revelatum est
JOHN|12|39|propterea non poterant credere quia iterum dixit Esaias
JOHN|12|40|excaecavit oculos eorum et induravit eorum cor ut non videant oculis et intellegant corde et convertantur et sanem eos
JOHN|12|41|haec dixit Esaias quando vidit gloriam eius et locutus est de eo
JOHN|12|42|verumtamen et ex principibus multi crediderunt in eum sed propter Pharisaeos non confitebantur ut de synagoga non eicerentur
JOHN|12|43|dilexerunt enim gloriam hominum magis quam gloriam Dei
JOHN|12|44|Iesus autem clamavit et dixit qui credit in me non credit in me sed in eum qui misit me
JOHN|12|45|et qui videt me videt eum qui misit me
JOHN|12|46|ego lux in mundum veni ut omnis qui credit in me in tenebris non maneat
JOHN|12|47|et si quis audierit verba mea et non custodierit ego non iudico eum non enim veni ut iudicem mundum sed ut salvificem mundum
JOHN|12|48|qui spernit me et non accipit verba mea habet qui iudicet eum sermo quem locutus sum ille iudicabit eum in novissimo die
JOHN|12|49|quia ego ex me ipso non sum locutus sed qui misit me Pater ipse mihi mandatum dedit quid dicam et quid loquar
JOHN|12|50|et scio quia mandatum eius vita aeterna est quae ergo ego loquor sicut dixit mihi Pater sic loquor
JOHN|13|1|ante diem autem festum paschae sciens Iesus quia venit eius hora ut transeat ex hoc mundo ad Patrem cum dilexisset suos qui erant in mundo in finem dilexit eos
JOHN|13|2|et cena facta cum diabolus iam misisset in corde ut traderet eum Iudas Simonis Scariotis
JOHN|13|3|sciens quia omnia dedit ei Pater in manus et quia a Deo exivit et ad Deum vadit
JOHN|13|4|surgit a cena et ponit vestimenta sua et cum accepisset linteum praecinxit se
JOHN|13|5|deinde mittit aquam in pelvem et coepit lavare pedes discipulorum et extergere linteo quo erat praecinctus
JOHN|13|6|venit ergo ad Simonem Petrum et dicit ei Petrus Domine tu mihi lavas pedes
JOHN|13|7|respondit Iesus et dicit ei quod ego facio tu nescis modo scies autem postea
JOHN|13|8|dicit ei Petrus non lavabis mihi pedes in aeternum respondit Iesus ei si non lavero te non habes partem mecum
JOHN|13|9|dicit ei Simon Petrus Domine non tantum pedes meos sed et manus et caput
JOHN|13|10|dicit ei Iesus qui lotus est non indiget ut lavet sed est mundus totus et vos mundi estis sed non omnes
JOHN|13|11|sciebat enim quisnam esset qui traderet eum propterea dixit non estis mundi omnes
JOHN|13|12|postquam ergo lavit pedes eorum et accepit vestimenta sua cum recubuisset iterum dixit eis scitis quid fecerim vobis
JOHN|13|13|vos vocatis me magister et Domine et bene dicitis sum etenim
JOHN|13|14|si ergo ego lavi vestros pedes Dominus et magister et vos debetis alter alterius lavare pedes
JOHN|13|15|exemplum enim dedi vobis ut quemadmodum ego feci vobis ita et vos faciatis
JOHN|13|16|amen amen dico vobis non est servus maior domino suo neque apostolus maior eo qui misit illum
JOHN|13|17|si haec scitis beati eritis si feceritis ea
JOHN|13|18|non de omnibus vobis dico ego scio quos elegerim sed ut impleatur scriptura qui manducat mecum panem levavit contra me calcaneum suum
JOHN|13|19|amodo dico vobis priusquam fiat ut credatis cum factum fuerit quia ego sum
JOHN|13|20|amen amen dico vobis qui accipit si quem misero me accipit qui autem me accipit accipit eum qui me misit
JOHN|13|21|cum haec dixisset Iesus turbatus est spiritu et protestatus est et dixit amen amen dico vobis quia unus ex vobis tradet me
JOHN|13|22|aspiciebant ergo ad invicem discipuli haesitantes de quo diceret
JOHN|13|23|erat ergo recumbens unus ex discipulis eius in sinu Iesu quem diligebat Iesus
JOHN|13|24|innuit ergo huic Simon Petrus et dicit ei quis est de quo dicit
JOHN|13|25|itaque cum recubuisset ille supra pectus Iesu dicit ei Domine quis est
JOHN|13|26|respondit Iesus ille est cui ego intinctum panem porrexero et cum intinxisset panem dedit Iudae Simonis Scariotis
JOHN|13|27|et post buccellam tunc introivit in illum Satanas dicit ei Iesus quod facis fac citius
JOHN|13|28|hoc autem nemo scivit discumbentium ad quid dixerit ei
JOHN|13|29|quidam enim putabant quia loculos habebat Iudas quia dicit ei Iesus eme ea quae opus sunt nobis ad diem festum aut egenis ut aliquid daret
JOHN|13|30|cum ergo accepisset ille buccellam exivit continuo erat autem nox
JOHN|13|31|cum ergo exisset dicit Iesus nunc clarificatus est Filius hominis et Deus clarificatus est in eo
JOHN|13|32|si Deus clarificatus est in eo et Deus clarificabit eum in semet ipso et continuo clarificabit eum
JOHN|13|33|filioli adhuc modicum vobiscum sum quaeretis me et sicut dixi Iudaeis quo ego vado vos non potestis venire et vobis dico modo
JOHN|13|34|mandatum novum do vobis ut diligatis invicem sicut dilexi vos ut et vos diligatis invicem
JOHN|13|35|in hoc cognoscent omnes quia mei discipuli estis si dilectionem habueritis ad invicem
JOHN|13|36|dicit ei Simon Petrus Domine quo vadis respondit Iesus quo ego vado non potes me modo sequi sequeris autem postea
JOHN|13|37|dicit ei Petrus quare non possum sequi te modo animam meam pro te ponam
JOHN|13|38|respondit Iesus animam tuam pro me ponis amen amen dico tibi non cantabit gallus donec me ter neges
JOHN|14|1|non turbetur cor vestrum creditis in Deum et in me credite
JOHN|14|2|in domo Patris mei mansiones multae sunt si quo minus dixissem vobis quia vado parare vobis locum
JOHN|14|3|et si abiero et praeparavero vobis locum iterum venio et accipiam vos ad me ipsum ut ubi sum ego et vos sitis
JOHN|14|4|et quo ego vado scitis et viam scitis
JOHN|14|5|dicit ei Thomas Domine nescimus quo vadis et quomodo possumus viam scire
JOHN|14|6|dicit ei Iesus ego sum via et veritas et vita nemo venit ad Patrem nisi per me
JOHN|14|7|si cognovissetis me et Patrem meum utique cognovissetis et amodo cognoscitis eum et vidistis eum
JOHN|14|8|dicit ei Philippus Domine ostende nobis Patrem et sufficit nobis
JOHN|14|9|dicit ei Iesus tanto tempore vobiscum sum et non cognovistis me Philippe qui vidit me vidit et Patrem quomodo tu dicis ostende nobis Patrem
JOHN|14|10|non credis quia ego in Patre et Pater in me est verba quae ego loquor vobis a me ipso non loquor Pater autem in me manens ipse facit opera
JOHN|14|11|non creditis quia ego in Patre et Pater in me est
JOHN|14|12|alioquin propter opera ipsa credite amen amen dico vobis qui credit in me opera quae ego facio et ipse faciet et maiora horum faciet quia ego ad Patrem vado
JOHN|14|13|et quodcumque petieritis in nomine meo hoc faciam ut glorificetur Pater in Filio
JOHN|14|14|si quid petieritis me in nomine meo hoc faciam
JOHN|14|15|si diligitis me mandata mea servate
JOHN|14|16|et ego rogabo Patrem et alium paracletum dabit vobis ut maneat vobiscum in aeternum
JOHN|14|17|Spiritum veritatis quem mundus non potest accipere quia non videt eum nec scit eum vos autem cognoscitis eum quia apud vos manebit et in vobis erit
JOHN|14|18|non relinquam vos orfanos veniam ad vos
JOHN|14|19|adhuc modicum et mundus me iam non videt vos autem videtis me quia ego vivo et vos vivetis
JOHN|14|20|in illo die vos cognoscetis quia ego sum in Patre meo et vos in me et ego in vobis
JOHN|14|21|qui habet mandata mea et servat ea ille est qui diligit me qui autem diligit me diligetur a Patre meo et ego diligam eum et manifestabo ei me ipsum
JOHN|14|22|dicit ei Iudas non ille Scariotis Domine quid factum est quia nobis manifestaturus es te ipsum et non mundo
JOHN|14|23|respondit Iesus et dixit ei si quis diligit me sermonem meum servabit et Pater meus diliget eum et ad eum veniemus et mansiones apud eum faciemus
JOHN|14|24|qui non diligit me sermones meos non servat et sermonem quem audistis non est meus sed eius qui misit me Patris
JOHN|14|25|haec locutus sum vobis apud vos manens
JOHN|14|26|paracletus autem Spiritus Sanctus quem mittet Pater in nomine meo ille vos docebit omnia et suggeret vobis omnia quaecumque dixero vobis
JOHN|14|27|pacem relinquo vobis pacem meam do vobis non quomodo mundus dat ego do vobis non turbetur cor vestrum neque formidet
JOHN|14|28|audistis quia ego dixi vobis vado et venio ad vos si diligeretis me gauderetis utique quia vado ad Patrem quia Pater maior me est
JOHN|14|29|et nunc dixi vobis priusquam fiat ut cum factum fuerit credatis
JOHN|14|30|iam non multa loquar vobiscum venit enim princeps mundi huius et in me non habet quicquam
JOHN|14|31|sed ut cognoscat mundus quia diligo Patrem et sicut mandatum dedit mihi Pater sic facio surgite eamus hinc
JOHN|15|1|ego sum vitis vera et Pater meus agricola est
JOHN|15|2|omnem palmitem in me non ferentem fructum tollet eum et omnem qui fert fructum purgabit eum ut fructum plus adferat
JOHN|15|3|iam vos mundi estis propter sermonem quem locutus sum vobis
JOHN|15|4|manete in me et ego in vobis sicut palmes non potest ferre fructum a semet ipso nisi manserit in vite sic nec vos nisi in me manseritis
JOHN|15|5|ego sum vitis vos palmites qui manet in me et ego in eo hic fert fructum multum quia sine me nihil potestis facere
JOHN|15|6|si quis in me non manserit mittetur foras sicut palmes et aruit et colligent eos et in ignem mittunt et ardent
JOHN|15|7|si manseritis in me et verba mea in vobis manserint quodcumque volueritis petetis et fiet vobis
JOHN|15|8|in hoc clarificatus est Pater meus ut fructum plurimum adferatis et efficiamini mei discipuli
JOHN|15|9|sicut dilexit me Pater et ego dilexi vos manete in dilectione mea
JOHN|15|10|si praecepta mea servaveritis manebitis in dilectione mea sicut et ego Patris mei praecepta servavi et maneo in eius dilectione
JOHN|15|11|haec locutus sum vobis ut gaudium meum in vobis sit et gaudium vestrum impleatur
JOHN|15|12|hoc est praeceptum meum ut diligatis invicem sicut dilexi vos
JOHN|15|13|maiorem hac dilectionem nemo habet ut animam suam quis ponat pro amicis suis
JOHN|15|14|vos amici mei estis si feceritis quae ego praecipio vobis
JOHN|15|15|iam non dico vos servos quia servus nescit quid facit dominus eius vos autem dixi amicos quia omnia quaecumque audivi a Patre meo nota feci vobis
JOHN|15|16|non vos me elegistis sed ego elegi vos et posui vos ut eatis et fructum adferatis et fructus vester maneat ut quodcumque petieritis Patrem in nomine meo det vobis
JOHN|15|17|haec mando vobis ut diligatis invicem
JOHN|15|18|si mundus vos odit scitote quia me priorem vobis odio habuit
JOHN|15|19|si de mundo fuissetis mundus quod suum erat diligeret quia vero de mundo non estis sed ego elegi vos de mundo propterea odit vos mundus
JOHN|15|20|mementote sermonis mei quem ego dixi vobis non est servus maior domino suo si me persecuti sunt et vos persequentur si sermonem meum servaverunt et vestrum servabunt
JOHN|15|21|sed haec omnia facient vobis propter nomen meum quia nesciunt eum qui misit me
JOHN|15|22|si non venissem et locutus fuissem eis peccatum non haberent nunc autem excusationem non habent de peccato suo
JOHN|15|23|qui me odit et Patrem meum odit
JOHN|15|24|si opera non fecissem in eis quae nemo alius fecit peccatum non haberent nunc autem et viderunt et oderunt et me et Patrem meum
JOHN|15|25|sed ut impleatur sermo qui in lege eorum scriptus est quia odio me habuerunt gratis
JOHN|15|26|cum autem venerit paracletus quem ego mittam vobis a Patre Spiritum veritatis qui a Patre procedit ille testimonium perhibebit de me
JOHN|15|27|et vos testimonium perhibetis quia ab initio mecum estis
JOHN|16|1|haec locutus sum vobis ut non scandalizemini
JOHN|16|2|absque synagogis facient vos sed venit hora ut omnis qui interficit vos arbitretur obsequium se praestare Deo
JOHN|16|3|et haec facient quia non noverunt Patrem neque me
JOHN|16|4|sed haec locutus sum vobis ut cum venerit hora eorum reminiscamini quia ego dixi vobis
JOHN|16|5|haec autem vobis ab initio non dixi quia vobiscum eram at nunc vado ad eum qui me misit et nemo ex vobis interrogat me quo vadis
JOHN|16|6|sed quia haec locutus sum vobis tristitia implevit cor vestrum
JOHN|16|7|sed ego veritatem dico vobis expedit vobis ut ego vadam si enim non abiero paracletus non veniet ad vos si autem abiero mittam eum ad vos
JOHN|16|8|et cum venerit ille arguet mundum de peccato et de iustitia et de iudicio
JOHN|16|9|de peccato quidem quia non credunt in me
JOHN|16|10|de iustitia vero quia ad Patrem vado et iam non videbitis me
JOHN|16|11|de iudicio autem quia princeps mundi huius iudicatus est
JOHN|16|12|adhuc multa habeo vobis dicere sed non potestis portare modo
JOHN|16|13|cum autem venerit ille Spiritus veritatis docebit vos in omnem veritatem non enim loquetur a semet ipso sed quaecumque audiet loquetur et quae ventura sunt adnuntiabit vobis
JOHN|16|14|ille me clarificabit quia de meo accipiet et adnuntiabit vobis
JOHN|16|15|omnia quaecumque habet Pater mea sunt propterea dixi quia de meo accipit et adnuntiabit vobis
JOHN|16|16|modicum et iam non videbitis me et iterum modicum et videbitis me quia vado ad Patrem
JOHN|16|17|dixerunt ergo ex discipulis eius ad invicem quid est hoc quod dicit nobis modicum et non videbitis me et iterum modicum et videbitis me et quia vado ad Patrem
JOHN|16|18|dicebant ergo quid est hoc quod dicit modicum nescimus quid loquitur
JOHN|16|19|cognovit autem Iesus quia volebant eum interrogare et dixit eis de hoc quaeritis inter vos quia dixi modicum et non videbitis me et iterum modicum et videbitis me
JOHN|16|20|amen amen dico vobis quia plorabitis et flebitis vos mundus autem gaudebit vos autem contristabimini sed tristitia vestra vertetur in gaudium
JOHN|16|21|mulier cum parit tristitiam habet quia venit hora eius cum autem pepererit puerum iam non meminit pressurae propter gaudium quia natus est homo in mundum
JOHN|16|22|et vos igitur nunc quidem tristitiam habetis iterum autem videbo vos et gaudebit cor vestrum et gaudium vestrum nemo tollit a vobis
JOHN|16|23|et in illo die me non rogabitis quicquam amen amen dico vobis si quid petieritis Patrem in nomine meo dabit vobis
JOHN|16|24|usque modo non petistis quicquam in nomine meo petite et accipietis ut gaudium vestrum sit plenum
JOHN|16|25|haec in proverbiis locutus sum vobis venit hora cum iam non in proverbiis loquar vobis sed palam de Patre adnuntiabo vobis
JOHN|16|26|illo die in nomine meo petetis et non dico vobis quia ego rogabo Patrem de vobis
JOHN|16|27|ipse enim Pater amat vos quia vos me amastis et credidistis quia ego a Deo exivi
JOHN|16|28|exivi a Patre et veni in mundum iterum relinquo mundum et vado ad Patrem
JOHN|16|29|dicunt ei discipuli eius ecce nunc palam loqueris et proverbium nullum dicis
JOHN|16|30|nunc scimus quia scis omnia et non opus est tibi ut quis te interroget in hoc credimus quia a Deo existi
JOHN|16|31|respondit eis Iesus modo creditis
JOHN|16|32|ecce venit hora et iam venit ut dispergamini unusquisque in propria et me solum relinquatis et non sum solus quia Pater mecum est
JOHN|16|33|haec locutus sum vobis ut in me pacem habeatis in mundo pressuram habetis sed confidite ego vici mundum
JOHN|17|1|haec locutus est Iesus et sublevatis oculis in caelum dixit Pater venit hora clarifica Filium tuum ut Filius tuus clarificet te
JOHN|17|2|sicut dedisti ei potestatem omnis carnis ut omne quod dedisti ei det eis vitam aeternam
JOHN|17|3|haec est autem vita aeterna ut cognoscant te solum verum Deum et quem misisti Iesum Christum
JOHN|17|4|ego te clarificavi super terram opus consummavi quod dedisti mihi ut faciam
JOHN|17|5|et nunc clarifica me tu Pater apud temet ipsum claritatem quam habui priusquam mundus esset apud te
JOHN|17|6|manifestavi nomen tuum hominibus quos dedisti mihi de mundo tui erant et mihi eos dedisti et sermonem tuum servaverunt
JOHN|17|7|nunc cognoverunt quia omnia quae dedisti mihi abs te sunt
JOHN|17|8|quia verba quae dedisti mihi dedi eis et ipsi acceperunt et cognoverunt vere quia a te exivi et crediderunt quia tu me misisti
JOHN|17|9|ego pro eis rogo non pro mundo rogo sed pro his quos dedisti mihi quia tui sunt
JOHN|17|10|et mea omnia tua sunt et tua mea sunt et clarificatus sum in eis
JOHN|17|11|et iam non sum in mundo et hii in mundo sunt et ego ad te venio Pater sancte serva eos in nomine tuo quos dedisti mihi ut sint unum sicut et nos
JOHN|17|12|cum essem cum eis ego servabam eos in nomine tuo quos dedisti mihi custodivi et nemo ex his perivit nisi filius perditionis ut scriptura impleatur
JOHN|17|13|nunc autem ad te venio et haec loquor in mundo ut habeant gaudium meum impletum in semet ipsis
JOHN|17|14|ego dedi eis sermonem tuum et mundus odio eos habuit quia non sunt de mundo sicut et ego non sum de mundo
JOHN|17|15|non rogo ut tollas eos de mundo sed ut serves eos ex malo
JOHN|17|16|de mundo non sunt sicut et ego non sum de mundo
JOHN|17|17|sanctifica eos in veritate sermo tuus veritas est
JOHN|17|18|sicut me misisti in mundum et ego misi eos in mundum
JOHN|17|19|et pro eis ego sanctifico me ipsum ut sint et ipsi sanctificati in veritate
JOHN|17|20|non pro his autem rogo tantum sed et pro eis qui credituri sunt per verbum eorum in me
JOHN|17|21|ut omnes unum sint sicut tu Pater in me et ego in te ut et ipsi in nobis unum sint ut mundus credat quia tu me misisti
JOHN|17|22|et ego claritatem quam dedisti mihi dedi eis ut sint unum sicut nos unum sumus
JOHN|17|23|ego in eis et tu in me ut sint consummati in unum et cognoscat mundus quia tu me misisti et dilexisti eos sicut me dilexisti
JOHN|17|24|Pater quos dedisti mihi volo ut ubi ego sum et illi sint mecum ut videant claritatem meam quam dedisti mihi quia dilexisti me ante constitutionem mundi
JOHN|17|25|Pater iuste et mundus te non cognovit ego autem te cognovi et hii cognoverunt quia tu me misisti
JOHN|17|26|et notum feci eis nomen tuum et notum faciam ut dilectio qua dilexisti me in ipsis sit et ego in ipsis
JOHN|18|1|haec cum dixisset Iesus egressus est cum discipulis suis trans torrentem Cedron ubi erat hortus in quem introivit ipse et discipuli eius
JOHN|18|2|sciebat autem et Iudas qui tradebat eum ipsum locum quia frequenter Iesus convenerat illuc cum discipulis suis
JOHN|18|3|Iudas ergo cum accepisset cohortem et a pontificibus et Pharisaeis ministros venit illuc cum lanternis et facibus et armis
JOHN|18|4|Iesus itaque sciens omnia quae ventura erant super eum processit et dicit eis quem quaeritis
JOHN|18|5|responderunt ei Iesum Nazarenum dicit eis Iesus ego sum stabat autem et Iudas qui tradebat eum cum ipsis
JOHN|18|6|ut ergo dixit eis ego sum abierunt retrorsum et ceciderunt in terram
JOHN|18|7|iterum ergo eos interrogavit quem quaeritis illi autem dixerunt Iesum Nazarenum
JOHN|18|8|respondit Iesus dixi vobis quia ego sum si ergo me quaeritis sinite hos abire
JOHN|18|9|ut impleretur sermo quem dixit quia quos dedisti mihi non perdidi ex ipsis quemquam
JOHN|18|10|Simon ergo Petrus habens gladium eduxit eum et percussit pontificis servum et abscidit eius auriculam dextram erat autem nomen servo Malchus
JOHN|18|11|dixit ergo Iesus Petro mitte gladium in vaginam calicem quem dedit mihi Pater non bibam illum
JOHN|18|12|cohors ergo et tribunus et ministri Iudaeorum conprehenderunt Iesum et ligaverunt eum
JOHN|18|13|et adduxerunt eum ad Annam primum erat enim socer Caiaphae qui erat pontifex anni illius
JOHN|18|14|erat autem Caiaphas qui consilium dederat Iudaeis quia expedit unum hominem mori pro populo
JOHN|18|15|sequebatur autem Iesum Simon Petrus et alius discipulus discipulus autem ille erat notus pontifici et introivit cum Iesu in atrium pontificis
JOHN|18|16|Petrus autem stabat ad ostium foris exivit ergo discipulus alius qui erat notus pontifici et dixit ostiariae et introduxit Petrum
JOHN|18|17|dicit ergo Petro ancilla ostiaria numquid et tu ex discipulis es hominis istius dicit ille non sum
JOHN|18|18|stabant autem servi et ministri ad prunas quia frigus erat et calefiebant erat autem cum eis et Petrus stans et calefaciens se
JOHN|18|19|pontifex ergo interrogavit Iesum de discipulis suis et de doctrina eius
JOHN|18|20|respondit ei Iesus ego palam locutus sum mundo ego semper docui in synagoga et in templo quo omnes Iudaei conveniunt et in occulto locutus sum nihil
JOHN|18|21|quid me interrogas interroga eos qui audierunt quid locutus sum ipsis ecce hii sciunt quae dixerim ego
JOHN|18|22|haec autem cum dixisset unus adsistens ministrorum dedit alapam Iesu dicens sic respondes pontifici
JOHN|18|23|respondit ei Iesus si male locutus sum testimonium perhibe de malo si autem bene quid me caedis
JOHN|18|24|et misit eum Annas ligatum ad Caiaphan pontificem
JOHN|18|25|erat autem Simon Petrus stans et calefaciens se dixerunt ergo ei numquid et tu ex discipulis eius es negavit ille et dixit non sum
JOHN|18|26|dicit unus ex servis pontificis cognatus eius cuius abscidit Petrus auriculam nonne ego te vidi in horto cum illo
JOHN|18|27|iterum ergo negavit Petrus et statim gallus cantavit
JOHN|18|28|adducunt ergo Iesum a Caiapha in praetorium erat autem mane et ipsi non introierunt in praetorium ut non contaminarentur sed manducarent pascha
JOHN|18|29|exivit ergo Pilatus ad eos foras et dixit quam accusationem adfertis adversus hominem hunc
JOHN|18|30|responderunt et dixerunt ei si non esset hic malefactor non tibi tradidissemus eum
JOHN|18|31|dixit ergo eis Pilatus accipite eum vos et secundum legem vestram iudicate eum dixerunt ergo ei Iudaei nobis non licet interficere quemquam
JOHN|18|32|ut sermo Iesu impleretur quem dixit significans qua esset morte moriturus
JOHN|18|33|introivit ergo iterum in praetorium Pilatus et vocavit Iesum et dixit ei tu es rex Iudaeorum
JOHN|18|34|et respondit Iesus a temet ipso hoc dicis an alii tibi dixerunt de me
JOHN|18|35|respondit Pilatus numquid ego Iudaeus sum gens tua et pontifices tradiderunt te mihi quid fecisti
JOHN|18|36|respondit Iesus regnum meum non est de mundo hoc si ex hoc mundo esset regnum meum ministri mei decertarent ut non traderer Iudaeis nunc autem meum regnum non est hinc
JOHN|18|37|dixit itaque ei Pilatus ergo rex es tu respondit Iesus tu dicis quia rex sum ego ego in hoc natus sum et ad hoc veni in mundum ut testimonium perhibeam veritati omnis qui est ex veritate audit meam vocem
JOHN|18|38|dicit ei Pilatus quid est veritas et cum hoc dixisset iterum exivit ad Iudaeos et dicit eis ego nullam invenio in eo causam
JOHN|18|39|est autem consuetudo vobis ut unum dimittam vobis in pascha vultis ergo dimittam vobis regem Iudaeorum
JOHN|18|40|clamaverunt rursum omnes dicentes non hunc sed Barabban erat autem Barabbas latro
JOHN|19|1|tunc ergo adprehendit Pilatus Iesum et flagellavit
JOHN|19|2|et milites plectentes coronam de spinis inposuerunt capiti eius et veste purpurea circumdederunt eum
JOHN|19|3|et veniebant ad eum et dicebant have rex Iudaeorum et dabant ei alapas
JOHN|19|4|exiit iterum Pilatus foras et dicit eis ecce adduco vobis eum foras
JOHN|19|5|ut cognoscatis quia in eo nullam causam invenio et purpureum vestimentum et dicit eis ecce homo
JOHN|19|6|cum ergo vidissent eum pontifices et ministri clamabant dicentes crucifige crucifige dicit eis Pilatus accipite eum vos et crucifigite ego enim non invenio in eo causam
JOHN|19|7|responderunt ei Iudaei nos legem habemus et secundum legem debet mori quia Filium Dei se fecit
JOHN|19|8|cum ergo audisset Pilatus hunc sermonem magis timuit
JOHN|19|9|et ingressus est praetorium iterum et dicit ad Iesum unde es tu Iesus autem responsum non dedit ei
JOHN|19|10|dicit ergo ei Pilatus mihi non loqueris nescis quia potestatem habeo crucifigere te et potestatem habeo dimittere te
JOHN|19|11|respondit Iesus non haberes potestatem adversum me ullam nisi tibi esset datum desuper propterea qui tradidit me tibi maius peccatum habet
JOHN|19|12|exinde quaerebat Pilatus dimittere eum Iudaei autem clamabant dicentes si hunc dimittis non es amicus Caesaris omnis qui se regem facit contradicit Caesari
JOHN|19|13|Pilatus ergo cum audisset hos sermones adduxit foras Iesum et sedit pro tribunali in locum qui dicitur Lithostrotus hebraice autem Gabbatha
JOHN|19|14|erat autem parasceve paschae hora quasi sexta et dicit Iudaeis ecce rex vester
JOHN|19|15|illi autem clamabant tolle tolle crucifige eum dixit eis Pilatus regem vestrum crucifigam responderunt pontifices non habemus regem nisi Caesarem
JOHN|19|16|tunc ergo tradidit eis illum ut crucifigeretur susceperunt autem Iesum et eduxerunt
JOHN|19|17|et baiulans sibi crucem exivit in eum qui dicitur Calvariae locum hebraice Golgotha
JOHN|19|18|ubi eum crucifixerunt et cum eo alios duos hinc et hinc medium autem Iesum
JOHN|19|19|scripsit autem et titulum Pilatus et posuit super crucem erat autem scriptum Iesus Nazarenus rex Iudaeorum
JOHN|19|20|hunc ergo titulum multi legerunt Iudaeorum quia prope civitatem erat locus ubi crucifixus est Iesus et erat scriptum hebraice graece et latine
JOHN|19|21|dicebant ergo Pilato pontifices Iudaeorum noli scribere rex Iudaeorum sed quia ipse dixit rex sum Iudaeorum
JOHN|19|22|respondit Pilatus quod scripsi scripsi
JOHN|19|23|milites ergo cum crucifixissent eum acceperunt vestimenta eius et fecerunt quattuor partes unicuique militi partem et tunicam erat autem tunica inconsutilis desuper contexta per totum
JOHN|19|24|dixerunt ergo ad invicem non scindamus eam sed sortiamur de illa cuius sit ut scriptura impleatur dicens partiti sunt vestimenta mea sibi et in vestem meam miserunt sortem et milites quidem haec fecerunt
JOHN|19|25|stabant autem iuxta crucem Iesu mater eius et soror matris eius Maria Cleopae et Maria Magdalene
JOHN|19|26|cum vidisset ergo Iesus matrem et discipulum stantem quem diligebat dicit matri suae mulier ecce filius tuus
JOHN|19|27|deinde dicit discipulo ecce mater tua et ex illa hora accepit eam discipulus in sua
JOHN|19|28|postea sciens Iesus quia iam omnia consummata sunt ut consummaretur scriptura dicit sitio
JOHN|19|29|vas ergo positum erat aceto plenum illi autem spongiam plenam aceto hysopo circumponentes obtulerunt ori eius
JOHN|19|30|cum ergo accepisset Iesus acetum dixit consummatum est et inclinato capite tradidit spiritum
JOHN|19|31|Iudaei ergo quoniam parasceve erat ut non remanerent in cruce corpora sabbato erat enim magnus dies ille sabbati rogaverunt Pilatum ut frangerentur eorum crura et tollerentur
JOHN|19|32|venerunt ergo milites et primi quidem fregerunt crura et alterius qui crucifixus est cum eo
JOHN|19|33|ad Iesum autem cum venissent ut viderunt eum iam mortuum non fregerunt eius crura
JOHN|19|34|sed unus militum lancea latus eius aperuit et continuo exivit sanguis et aqua
JOHN|19|35|et qui vidit testimonium perhibuit et verum est eius testimonium et ille scit quia vera dicit ut et vos credatis
JOHN|19|36|facta sunt enim haec ut scriptura impleatur os non comminuetis ex eo
JOHN|19|37|et iterum alia scriptura dicit videbunt in quem transfixerunt
JOHN|19|38|post haec autem rogavit Pilatum Ioseph ab Arimathia eo quod esset discipulus Iesu occultus autem propter metum Iudaeorum ut tolleret corpus Iesu et permisit Pilatus venit ergo et tulit corpus Iesu
JOHN|19|39|venit autem et Nicodemus qui venerat ad Iesum nocte primum ferens mixturam murrae et aloes quasi libras centum
JOHN|19|40|acceperunt ergo corpus Iesu et ligaverunt eum linteis cum aromatibus sicut mos Iudaeis est sepelire
JOHN|19|41|erat autem in loco ubi crucifixus est hortus et in horto monumentum novum in quo nondum quisquam positus erat
JOHN|19|42|ibi ergo propter parasceven Iudaeorum quia iuxta erat monumentum posuerunt Iesum
JOHN|20|1|una autem sabbati Maria Magdalene venit mane cum adhuc tenebrae essent ad monumentum et videt lapidem sublatum a monumento
JOHN|20|2|cucurrit ergo et venit ad Simonem Petrum et ad alium discipulum quem amabat Iesus et dicit eis tulerunt Dominum de monumento et nescimus ubi posuerunt eum
JOHN|20|3|exiit ergo Petrus et ille alius discipulus et venerunt ad monumentum
JOHN|20|4|currebant autem duo simul et ille alius discipulus praecucurrit citius Petro et venit primus ad monumentum
JOHN|20|5|et cum se inclinasset videt posita linteamina non tamen introivit
JOHN|20|6|venit ergo Simon Petrus sequens eum et introivit in monumentum et videt linteamina posita
JOHN|20|7|et sudarium quod fuerat super caput eius non cum linteaminibus positum sed separatim involutum in unum locum
JOHN|20|8|tunc ergo introivit et ille discipulus qui venerat primus ad monumentum et vidit et credidit
JOHN|20|9|nondum enim sciebant scripturam quia oportet eum a mortuis resurgere
JOHN|20|10|abierunt ergo iterum ad semet ipsos discipuli
JOHN|20|11|Maria autem stabat ad monumentum foris plorans dum ergo fleret inclinavit se et prospexit in monumentum
JOHN|20|12|et vidit duos angelos in albis sedentes unum ad caput et unum ad pedes ubi positum fuerat corpus Iesu
JOHN|20|13|dicunt ei illi mulier quid ploras dicit eis quia tulerunt Dominum meum et nescio ubi posuerunt eum
JOHN|20|14|haec cum dixisset conversa est retrorsum et videt Iesum stantem et non sciebat quia Iesus est
JOHN|20|15|dicit ei Iesus mulier quid ploras quem quaeris illa existimans quia hortulanus esset dicit ei domine si tu sustulisti eum dicito mihi ubi posuisti eum et ego eum tollam
JOHN|20|16|dicit ei Iesus Maria conversa illa dicit ei rabboni quod dicitur magister
JOHN|20|17|dicit ei Iesus noli me tangere nondum enim ascendi ad Patrem meum vade autem ad fratres meos et dic eis ascendo ad Patrem meum et Patrem vestrum et Deum meum et Deum vestrum
JOHN|20|18|venit Maria Magdalene adnuntians discipulis quia vidi Dominum et haec dixit mihi
JOHN|20|19|cum esset ergo sero die illo una sabbatorum et fores essent clausae ubi erant discipuli propter metum Iudaeorum venit Iesus et stetit in medio et dicit eis pax vobis
JOHN|20|20|et hoc cum dixisset ostendit eis manus et latus gavisi sunt ergo discipuli viso Domino
JOHN|20|21|dixit ergo eis iterum pax vobis sicut misit me Pater et ego mitto vos
JOHN|20|22|hoc cum dixisset insuflavit et dicit eis accipite Spiritum Sanctum
JOHN|20|23|quorum remiseritis peccata remittuntur eis quorum retinueritis detenta sunt
JOHN|20|24|Thomas autem unus ex duodecim qui dicitur Didymus non erat cum eis quando venit Iesus
JOHN|20|25|dixerunt ergo ei alii discipuli vidimus Dominum ille autem dixit eis nisi videro in manibus eius figuram clavorum et mittam digitum meum in locum clavorum et mittam manum meam in latus eius non credam
JOHN|20|26|et post dies octo iterum erant discipuli eius intus et Thomas cum eis venit Iesus ianuis clausis et stetit in medio et dixit pax vobis
JOHN|20|27|deinde dicit Thomae infer digitum tuum huc et vide manus meas et adfer manum tuam et mitte in latus meum et noli esse incredulus sed fidelis
JOHN|20|28|respondit Thomas et dixit ei Dominus meus et Deus meus
JOHN|20|29|dicit ei Iesus quia vidisti me credidisti beati qui non viderunt et crediderunt
JOHN|20|30|multa quidem et alia signa fecit Iesus in conspectu discipulorum suorum quae non sunt scripta in libro hoc
JOHN|20|31|haec autem scripta sunt ut credatis quia Iesus est Christus Filius Dei et ut credentes vitam habeatis in nomine eius
JOHN|21|1|postea manifestavit se iterum Iesus ad mare Tiberiadis manifestavit autem sic
JOHN|21|2|erant simul Simon Petrus et Thomas qui dicitur Didymus et Nathanahel qui erat a Cana Galilaeae et filii Zebedaei et alii ex discipulis eius duo
JOHN|21|3|dicit eis Simon Petrus vado piscari dicunt ei venimus et nos tecum et exierunt et ascenderunt in navem et illa nocte nihil prendiderunt
JOHN|21|4|mane autem iam facto stetit Iesus in litore non tamen cognoverunt discipuli quia Iesus est
JOHN|21|5|dicit ergo eis Iesus pueri numquid pulmentarium habetis responderunt ei non
JOHN|21|6|dixit eis mittite in dexteram navigii rete et invenietis miserunt ergo et iam non valebant illud trahere a multitudine piscium
JOHN|21|7|dicit ergo discipulus ille quem diligebat Iesus Petro Dominus est Simon Petrus cum audisset quia Dominus est tunicam succinxit se erat enim nudus et misit se in mare
JOHN|21|8|alii autem discipuli navigio venerunt non enim longe erant a terra sed quasi a cubitis ducentis trahentes rete piscium
JOHN|21|9|ut ergo descenderunt in terram viderunt prunas positas et piscem superpositum et panem
JOHN|21|10|dicit eis Iesus adferte de piscibus quos prendidistis nunc
JOHN|21|11|ascendit Simon Petrus et traxit rete in terram plenum magnis piscibus centum quinquaginta tribus et cum tanti essent non est scissum rete
JOHN|21|12|dicit eis Iesus venite prandete et nemo audebat discentium interrogare eum tu quis es scientes quia Dominus esset
JOHN|21|13|et venit Iesus et accepit panem et dat eis et piscem similiter
JOHN|21|14|hoc iam tertio manifestatus est Iesus discipulis cum surrexisset a mortuis
JOHN|21|15|cum ergo prandissent dicit Simoni Petro Iesus Simon Iohannis diligis me plus his dicit ei etiam Domine tu scis quia amo te dicit ei pasce agnos meos
JOHN|21|16|dicit ei iterum Simon Iohannis diligis me ait illi etiam Domine tu scis quia amo te dicit ei pasce agnos meos
JOHN|21|17|dicit ei tertio Simon Iohannis amas me contristatus est Petrus quia dixit ei tertio amas me et dicit ei Domine tu omnia scis tu scis quia amo te dicit ei pasce oves meas
JOHN|21|18|amen amen dico tibi cum esses iunior cingebas te et ambulabas ubi volebas cum autem senueris extendes manus tuas et alius te cinget et ducet quo non vis
JOHN|21|19|hoc autem dixit significans qua morte clarificaturus esset Deum et hoc cum dixisset dicit ei sequere me
JOHN|21|20|conversus Petrus vidit illum discipulum quem diligebat Iesus sequentem qui et recubuit in cena super pectus eius et dixit Domine quis est qui tradit te
JOHN|21|21|hunc ergo cum vidisset Petrus dicit Iesu Domine hic autem quid
JOHN|21|22|dicit ei Iesus si sic eum volo manere donec veniam quid ad te tu me sequere
JOHN|21|23|exivit ergo sermo iste in fratres quia discipulus ille non moritur et non dixit ei Iesus non moritur sed si sic eum volo manere donec venio quid ad te
JOHN|21|24|hic est discipulus qui testimonium perhibet de his et scripsit haec et scimus quia verum est testimonium eius
JOHN|21|25|sunt autem et alia multa quae fecit Iesus quae si scribantur per singula nec ipsum arbitror mundum capere eos qui scribendi sunt libros amen
ACTS|1|1|primum quidem sermonem feci de omnibus o Theophile quae coepit Iesus facere et docere
ACTS|1|2|usque in diem qua praecipiens apostolis per Spiritum Sanctum quos elegit adsumptus est
ACTS|1|3|quibus et praebuit se ipsum vivum post passionem suam in multis argumentis per dies quadraginta apparens eis et loquens de regno Dei
ACTS|1|4|et convescens praecepit eis ab Hierosolymis ne discederent sed expectarent promissionem Patris quam audistis per os meum
ACTS|1|5|quia Iohannes quidem baptizavit aqua vos autem baptizabimini Spiritu Sancto non post multos hos dies
ACTS|1|6|igitur qui convenerant interrogabant eum dicentes Domine si in tempore hoc restitues regnum Israhel
ACTS|1|7|dixit autem eis non est vestrum nosse tempora vel momenta quae Pater posuit in sua potestate
ACTS|1|8|sed accipietis virtutem supervenientis Spiritus Sancti in vos et eritis mihi testes in Hierusalem et in omni Iudaea et Samaria et usque ad ultimum terrae
ACTS|1|9|et cum haec dixisset videntibus illis elevatus est et nubes suscepit eum ab oculis eorum
ACTS|1|10|cumque intuerentur in caelum eunte illo ecce duo viri adstiterunt iuxta illos in vestibus albis
ACTS|1|11|qui et dixerunt viri galilaei quid statis aspicientes in caelum hic Iesus qui adsumptus est a vobis in caelum sic veniet quemadmodum vidistis eum euntem in caelum
ACTS|1|12|tunc reversi sunt Hierosolymam a monte qui vocatur Oliveti qui est iuxta Hierusalem sabbati habens iter
ACTS|1|13|et cum introissent in cenaculum ascenderunt ubi manebant Petrus et Iohannes Iacobus et Andreas Philippus et Thomas Bartholomeus et Mattheus Iacobus Alphei et Simon Zelotes et Iudas Iacobi
ACTS|1|14|hii omnes erant perseverantes unianimiter in oratione cum mulieribus et Maria matre Iesu et fratribus eius
ACTS|1|15|et in diebus illis exsurgens Petrus in medio fratrum dixit erat autem turba nominum simul fere centum viginti
ACTS|1|16|viri fratres oportet impleri scripturam quam praedixit Spiritus Sanctus per os David de Iuda qui fuit dux eorum qui conprehenderunt Iesum
ACTS|1|17|quia connumeratus erat in nobis et sortitus est sortem ministerii huius
ACTS|1|18|et hic quidem possedit agrum de mercede iniquitatis et suspensus crepuit medius et diffusa sunt omnia viscera eius
ACTS|1|19|et notum factum est omnibus habitantibus Hierusalem ita ut appellaretur ager ille lingua eorum Acheldemach hoc est ager Sanguinis
ACTS|1|20|scriptum est enim in libro Psalmorum fiat commoratio eius deserta et non sit qui inhabitet in ea et episcopatum eius accipiat alius
ACTS|1|21|oportet ergo ex his viris qui nobiscum congregati sunt in omni tempore quo intravit et exivit inter nos Dominus Iesus
ACTS|1|22|incipiens a baptismate Iohannis usque in diem qua adsumptus est a nobis testem resurrectionis eius nobiscum fieri unum ex istis
ACTS|1|23|et statuerunt duos Ioseph qui vocabatur Barsabban qui cognominatus est Iustus et Matthiam
ACTS|1|24|et orantes dixerunt tu Domine qui corda nosti omnium ostende quem elegeris ex his duobus unum
ACTS|1|25|accipere locum ministerii huius et apostolatus de quo praevaricatus est Iudas ut abiret in locum suum
ACTS|1|26|et dederunt sortes eis et cecidit sors super Matthiam et adnumeratus est cum undecim apostolis
ACTS|2|1|et cum conplerentur dies pentecostes erant omnes pariter in eodem loco
ACTS|2|2|et factus est repente de caelo sonus tamquam advenientis spiritus vehementis et replevit totam domum ubi erant sedentes
ACTS|2|3|et apparuerunt illis dispertitae linguae tamquam ignis seditque supra singulos eorum
ACTS|2|4|et repleti sunt omnes Spiritu Sancto et coeperunt loqui aliis linguis prout Spiritus Sanctus dabat eloqui illis
ACTS|2|5|erant autem in Hierusalem habitantes Iudaei viri religiosi ex omni natione quae sub caelo sunt
ACTS|2|6|facta autem hac voce convenit multitudo et mente confusa est quoniam audiebat unusquisque lingua sua illos loquentes
ACTS|2|7|stupebant autem omnes et mirabantur dicentes nonne omnes ecce isti qui loquuntur Galilaei sunt
ACTS|2|8|et quomodo nos audivimus unusquisque lingua nostra in qua nati sumus
ACTS|2|9|Parthi et Medi et Elamitae et qui habitant Mesopotamiam et Iudaeam et Cappadociam Pontum et Asiam
ACTS|2|10|Frygiam et Pamphiliam Aegyptum et partes Lybiae quae est circa Cyrenen et advenae romani
ACTS|2|11|Iudaei quoque et proselyti Cretes et Arabes audivimus loquentes eos nostris linguis magnalia Dei
ACTS|2|12|stupebant autem omnes et mirabantur ad invicem dicentes quidnam hoc vult esse
ACTS|2|13|alii autem inridentes dicebant quia musto pleni sunt isti
ACTS|2|14|stans autem Petrus cum undecim levavit vocem suam et locutus est eis viri iudaei et qui habitatis Hierusalem universi hoc vobis notum sit et auribus percipite verba mea
ACTS|2|15|non enim sicut vos aestimatis hii ebrii sunt cum sit hora diei tertia
ACTS|2|16|sed hoc est quod dictum est per prophetam Iohel
ACTS|2|17|et erit in novissimis diebus dicit Dominus effundam de Spiritu meo super omnem carnem et prophetabunt filii vestri et filiae vestrae et iuvenes vestri visiones videbunt et seniores vestri somnia somniabunt
ACTS|2|18|et quidem super servos meos et super ancillas meas in diebus illis effundam de Spiritu meo et prophetabunt
ACTS|2|19|et dabo prodigia in caelo sursum et signa in terra deorsum sanguinem et ignem et vaporem fumi
ACTS|2|20|sol convertetur in tenebras et luna in sanguinem antequam veniat dies Domini magnus et manifestus
ACTS|2|21|et erit omnis quicumque invocaverit nomen Domini salvus erit
ACTS|2|22|viri israhelitae audite verba haec Iesum Nazarenum virum adprobatum a Deo in vobis virtutibus et prodigiis et signis quae fecit per illum Deus in medio vestri sicut vos scitis
ACTS|2|23|hunc definito consilio et praescientia Dei traditum per manus iniquorum adfigentes interemistis
ACTS|2|24|quem Deus suscitavit solutis doloribus inferni iuxta quod inpossibile erat teneri illum ab eo
ACTS|2|25|David enim dicit in eum providebam Dominum coram me semper quoniam a dextris meis est ne commovear
ACTS|2|26|propter hoc laetatum est cor meum et exultavit lingua mea insuper et caro mea requiescet in spe
ACTS|2|27|quoniam non derelinques animam meam in inferno neque dabis Sanctum tuum videre corruptionem
ACTS|2|28|notas fecisti mihi vias vitae replebis me iucunditate cum facie tua
ACTS|2|29|viri fratres liceat audenter dicere ad vos de patriarcha David quoniam et defunctus est et sepultus est et sepulchrum eius est apud nos usque in hodiernum diem
ACTS|2|30|propheta igitur cum esset et sciret quia iureiurando iurasset illi Deus de fructu lumbi eius sedere super sedem eius
ACTS|2|31|providens locutus est de resurrectione Christi quia neque derelictus est in inferno neque caro eius vidit corruptionem
ACTS|2|32|hunc Iesum resuscitavit Deus cui omnes nos testes sumus
ACTS|2|33|dextera igitur Dei exaltatus et promissione Spiritus Sancti accepta a Patre effudit hunc quem vos videtis et audistis
ACTS|2|34|non enim David ascendit in caelos dicit autem ipse dixit Dominus Domino meo sede a dextris meis
ACTS|2|35|donec ponam inimicos tuos scabillum pedum tuorum
ACTS|2|36|certissime ergo sciat omnis domus Israhel quia et Dominum eum et Christum Deus fecit hunc Iesum quem vos crucifixistis
ACTS|2|37|his auditis conpuncti sunt corde et dixerunt ad Petrum et ad reliquos apostolos quid faciemus viri fratres
ACTS|2|38|Petrus vero ad illos paenitentiam inquit agite et baptizetur unusquisque vestrum in nomine Iesu Christi in remissionem peccatorum vestrorum et accipietis donum Sancti Spiritus
ACTS|2|39|vobis enim est repromissio et filiis vestris et omnibus qui longe sunt quoscumque advocaverit Dominus Deus noster
ACTS|2|40|aliis etiam verbis pluribus testificatus est et exhortabatur eos dicens salvamini a generatione ista prava
ACTS|2|41|qui ergo receperunt sermonem eius baptizati sunt et adpositae sunt in illa die animae circiter tria milia
ACTS|2|42|erant autem perseverantes in doctrina apostolorum et communicatione fractionis panis et orationibus
ACTS|2|43|fiebat autem omni animae timor multa quoque prodigia et signa per apostolos fiebant in Hierusalem et metus erat magnus in universis
ACTS|2|44|omnes etiam qui credebant erant pariter et habebant omnia communia
ACTS|2|45|possessiones et substantias vendebant et dividebant illa omnibus prout cuique opus erat
ACTS|2|46|cotidie quoque perdurantes unianimiter in templo et frangentes circa domos panem sumebant cibum cum exultatione et simplicitate cordis
ACTS|2|47|conlaudantes Deum et habentes gratiam ad omnem plebem Dominus autem augebat qui salvi fierent cotidie in id ipsum
ACTS|3|1|Petrus autem et Iohannes ascendebant in templum ad horam orationis nonam
ACTS|3|2|et quidam vir qui erat claudus ex utero matris suae baiulabatur quem ponebant cotidie ad portam templi quae dicitur Speciosa ut peteret elemosynam ab introeuntibus in templum
ACTS|3|3|is cum vidisset Petrum et Iohannem incipientes introire in templum rogabat ut elemosynam acciperet
ACTS|3|4|intuens autem in eum Petrus cum Iohanne dixit respice in nos
ACTS|3|5|at ille intendebat in eos sperans se aliquid accepturum ab eis
ACTS|3|6|Petrus autem dixit argentum et aurum non est mihi quod autem habeo hoc tibi do in nomine Iesu Christi Nazareni surge et ambula
ACTS|3|7|et adprehensa ei manu dextera adlevavit eum et protinus consolidatae sunt bases eius et plantae
ACTS|3|8|et exiliens stetit et ambulabat et intravit cum illis in templum ambulans et exiliens et laudans Dominum
ACTS|3|9|et vidit omnis populus eum ambulantem et laudantem Deum
ACTS|3|10|cognoscebant autem illum quoniam ipse erat qui ad elemosynam sedebat ad Speciosam portam templi et impleti sunt stupore et extasi in eo quod contigerat illi
ACTS|3|11|cum teneret autem Petrum et Iohannem concurrit omnis populus ad eos ad porticum qui appellatur Salomonis stupentes
ACTS|3|12|videns autem Petrus respondit ad populum viri israhelitae quid miramini in hoc aut nos quid intuemini quasi nostra virtute aut pietate fecerimus hunc ambulare
ACTS|3|13|Deus Abraham et Deus Isaac et Deus Iacob Deus patrum nostrorum glorificavit Filium suum Iesum quem vos quidem tradidistis et negastis ante faciem Pilati iudicante illo dimitti
ACTS|3|14|vos autem sanctum et iustum negastis et petistis virum homicidam donari vobis
ACTS|3|15|auctorem vero vitae interfecistis quem Deus suscitavit a mortuis cuius nos testes sumus
ACTS|3|16|et in fide nominis eius hunc quem videtis et nostis confirmavit nomen eius et fides quae per eum est dedit integram sanitatem istam in conspectu omnium vestrum
ACTS|3|17|et nunc fratres scio quia per ignorantiam fecistis sicut et principes vestri
ACTS|3|18|Deus autem quae praenuntiavit per os omnium prophetarum pati Christum suum implevit sic
ACTS|3|19|paenitemini igitur et convertimini ut deleantur vestra peccata
ACTS|3|20|ut cum venerint tempora refrigerii a conspectu Domini et miserit eum qui praedicatus est vobis Iesum Christum
ACTS|3|21|quem oportet caelum quidem suscipere usque in tempora restitutionis omnium quae locutus est Deus per os sanctorum suorum a saeculo prophetarum
ACTS|3|22|Moses quidem dixit quia prophetam vobis suscitabit Dominus Deus vester de fratribus vestris tamquam me ipsum audietis iuxta omnia quaecumque locutus fuerit vobis
ACTS|3|23|erit autem omnis anima quae non audierit prophetam illum exterminabitur de plebe
ACTS|3|24|et omnes prophetae a Samuhel et deinceps qui locuti sunt et adnuntiaverunt dies istos
ACTS|3|25|vos estis filii prophetarum et testamenti quod disposuit Deus ad patres vestros dicens ad Abraham et in semine tuo benedicentur omnes familiae terrae
ACTS|3|26|vobis primum Deus suscitans Filium suum misit eum benedicentem vobis ut convertat se unusquisque a nequitia sua
ACTS|4|1|loquentibus autem illis ad populum supervenerunt sacerdotes et magistratus templi et Sadducaei
ACTS|4|2|dolentes quod docerent populum et adnuntiarent in Iesu resurrectionem ex mortuis
ACTS|4|3|et iniecerunt in eis manus et posuerunt eos in custodiam in crastinum erat enim iam vespera
ACTS|4|4|multi autem eorum qui audierant verbum crediderunt et factus est numerus virorum quinque milia
ACTS|4|5|factum est autem in crastinum ut congregarentur principes eorum et seniores et scribae in Hierusalem
ACTS|4|6|et Annas princeps sacerdotum et Caiphas et Iohannes et Alexander et quotquot erant de genere sacerdotali
ACTS|4|7|et statuentes eos in medio interrogabant in qua virtute aut in quo nomine fecistis hoc vos
ACTS|4|8|tunc Petrus repletus Spiritu Sancto dixit ad eos principes populi et seniores
ACTS|4|9|si nos hodie diiudicamur in benefacto hominis infirmi in quo iste salvus factus est
ACTS|4|10|notum sit omnibus vobis et omni plebi Israhel quia in nomine Iesu Christi Nazareni quem vos crucifixistis quem Deus suscitavit a mortuis in hoc iste adstat coram vobis sanus
ACTS|4|11|hic est lapis qui reprobatus est a vobis aedificantibus qui factus est in caput anguli
ACTS|4|12|et non est in alio aliquo salus nec enim nomen aliud est sub caelo datum hominibus in quo oportet nos salvos fieri
ACTS|4|13|videntes autem Petri constantiam et Iohannis conperto quod homines essent sine litteris et idiotae admirabantur et cognoscebant eos quoniam cum Iesu fuerant
ACTS|4|14|hominem quoque videntes stantem cum eis qui curatus fuerat nihil poterant contradicere
ACTS|4|15|iusserunt autem eos foras extra concilium secedere et conferebant ad invicem
ACTS|4|16|dicentes quid faciemus hominibus istis quoniam quidem notum signum factum est per eos omnibus habitantibus in Hierusalem manifestum et non possumus negare
ACTS|4|17|sed ne amplius divulgetur in populum comminemur eis ne ultra loquantur in nomine hoc ulli hominum
ACTS|4|18|et vocantes eos denuntiaverunt ne omnino loquerentur neque docerent in nomine Iesu
ACTS|4|19|Petrus vero et Iohannes respondentes dixerunt ad eos si iustum est in conspectu Dei vos potius audire quam Deum iudicate
ACTS|4|20|non enim possumus quae vidimus et audivimus non loqui
ACTS|4|21|at illi comminantes dimiserunt eos non invenientes quomodo punirent eos propter populum quia omnes clarificabant Deum in eo quod acciderat
ACTS|4|22|annorum enim erat amplius quadraginta homo in quo factum erat signum istud sanitatis
ACTS|4|23|dimissi autem venerunt ad suos et adnuntiaverunt eis quanta ad eos principes sacerdotum et seniores dixissent
ACTS|4|24|qui cum audissent unianimiter levaverunt vocem ad Deum et dixerunt Domine tu qui fecisti caelum et terram et mare et omnia quae in eis sunt
ACTS|4|25|qui Spiritu Sancto per os patris nostri David pueri tui dixisti quare fremuerunt gentes et populi meditati sunt inania
ACTS|4|26|adstiterunt reges terrae et principes convenerunt in unum adversus Dominum et adversus Christum eius
ACTS|4|27|convenerunt enim vere in civitate ista adversus sanctum puerum tuum Iesum quem unxisti Herodes et Pontius Pilatus cum gentibus et populis Israhel
ACTS|4|28|facere quae manus tua et consilium decreverunt fieri
ACTS|4|29|et nunc Domine respice in minas eorum et da servis tuis cum omni fiducia loqui verbum tuum
ACTS|4|30|in eo cum manum tuam extendas sanitates et signa et prodigia fieri per nomen sancti Filii tui Iesu
ACTS|4|31|et cum orassent motus est locus in quo erant congregati et repleti sunt omnes Spiritu Sancto et loquebantur verbum Dei cum fiducia
ACTS|4|32|multitudinis autem credentium erat cor et anima una nec quisquam eorum quae possidebant aliquid suum esse dicebat sed erant illis omnia communia
ACTS|4|33|et virtute magna reddebant apostoli testimonium resurrectionis Iesu Christi Domini et gratia magna erat in omnibus illis
ACTS|4|34|neque enim quisquam egens erat inter illos quotquot enim possessores agrorum aut domorum erant vendentes adferebant pretia eorum quae vendebant
ACTS|4|35|et ponebant ante pedes apostolorum dividebantur autem singulis prout cuique opus erat
ACTS|4|36|Ioseph autem qui cognominatus est Barnabas ab apostolis quod est interpretatum Filius consolationis Levites Cyprius genere
ACTS|4|37|cum haberet agrum vendidit illum et adtulit pretium et posuit ante pedes apostolorum
ACTS|5|1|vir autem quidam nomine Ananias cum Saffira uxore sua vendidit agrum
ACTS|5|2|et fraudavit de pretio agri conscia uxore sua et adferens partem quandam ad pedes apostolorum posuit
ACTS|5|3|dixit autem Petrus Anania cur temptavit Satanas cor tuum mentiri te Spiritui Sancto et fraudare de pretio agri
ACTS|5|4|nonne manens tibi manebat et venundatum in tua erat potestate quare posuisti in corde tuo hanc rem non es mentitus hominibus sed Deo
ACTS|5|5|audiens autem Ananias haec verba cecidit et exspiravit et factus est timor magnus in omnes qui audierant
ACTS|5|6|surgentes autem iuvenes amoverunt eum et efferentes sepelierunt
ACTS|5|7|factum est autem quasi horarum trium spatium et uxor ipsius nesciens quod factum fuerat introiit
ACTS|5|8|respondit autem ei Petrus dic mihi si tanti agrum vendidistis at illa dixit etiam tanti
ACTS|5|9|Petrus autem ad eam quid utique convenit vobis temptare Spiritum Domini ecce pedes eorum qui sepelierunt virum tuum ad ostium et efferent te
ACTS|5|10|confestim cecidit ante pedes eius et exspiravit intrantes autem iuvenes invenerunt illam mortuam et extulerunt et sepelierunt ad virum suum
ACTS|5|11|et factus est timor magnus in universa ecclesia et in omnes qui audierunt haec
ACTS|5|12|per manus autem apostolorum fiebant signa et prodigia multa in plebe et erant unianimiter omnes in porticu Salomonis
ACTS|5|13|ceterorum autem nemo audebat coniungere se illis sed magnificabat eos populus
ACTS|5|14|magis autem augebatur credentium in Domino multitudo virorum ac mulierum
ACTS|5|15|ita ut in plateas eicerent infirmos et ponerent in lectulis et grabattis ut veniente Petro saltim umbra illius obumbraret quemquam eorum
ACTS|5|16|concurrebat autem et multitudo vicinarum civitatum Hierusalem adferentes aegros et vexatos ab spiritibus inmundis qui curabantur omnes
ACTS|5|17|exsurgens autem princeps sacerdotum et omnes qui cum illo erant quae est heresis Sadducaeorum repleti sunt zelo
ACTS|5|18|et iniecerunt manus in apostolos et posuerunt illos in custodia publica
ACTS|5|19|angelus autem Domini per noctem aperiens ianuas carceris et educens eos dixit
ACTS|5|20|ite et stantes loquimini in templo plebi omnia verba vitae huius
ACTS|5|21|qui cum audissent intraverunt diluculo in templum et docebant adveniens autem princeps sacerdotum et qui cum eo erant convocaverunt concilium et omnes seniores filiorum Israhel et miserunt in carcerem ut adducerentur
ACTS|5|22|cum venissent autem ministri et aperto carcere non invenissent illos reversi nuntiaverunt
ACTS|5|23|dicentes carcerem quidem invenimus clausum cum omni diligentia et custodes stantes ad ianuas aperientes autem neminem intus invenimus
ACTS|5|24|ut audierunt autem hos sermones magistratus templi et principes sacerdotum ambigebant de illis quidnam fieret
ACTS|5|25|adveniens autem quidam nuntiavit eis quia ecce viri quos posuistis in carcere sunt in templo stantes et docentes populum
ACTS|5|26|tunc abiit magistratus cum ministris et adduxit illos sine vi timebant enim populum ne lapidarentur
ACTS|5|27|et cum adduxissent illos statuerunt in concilio et interrogavit eos princeps sacerdotum
ACTS|5|28|dicens praecipiendo praecepimus vobis ne doceretis in nomine isto et ecce replestis Hierusalem doctrina vestra et vultis inducere super nos sanguinem hominis istius
ACTS|5|29|respondens autem Petrus et apostoli dixerunt oboedire oportet Deo magis quam hominibus
ACTS|5|30|Deus patrum nostrorum suscitavit Iesum quem vos interemistis suspendentes in ligno
ACTS|5|31|hunc Deus principem et salvatorem exaltavit dextera sua ad dandam paenitentiam Israhel et remissionem peccatorum
ACTS|5|32|et nos sumus testes horum verborum et Spiritus Sanctus quem dedit Deus omnibus oboedientibus sibi
ACTS|5|33|haec cum audissent dissecabantur et cogitabant interficere illos
ACTS|5|34|surgens autem quidam in concilio Pharisaeus nomine Gamalihel legis doctor honorabilis universae plebi iussit foras ad breve homines fieri
ACTS|5|35|dixitque ad illos viri israhelitae adtendite vobis super hominibus istis quid acturi sitis
ACTS|5|36|ante hos enim dies extitit Theodas dicens esse se aliquem cui consensit virorum numerus circiter quadringentorum qui occisus est et omnes quicumque credebant ei dissipati sunt et redactus est ad nihilum
ACTS|5|37|post hunc extitit Iudas Galilaeus in diebus professionis et avertit populum post se et ipse periit et omnes quotquot consenserunt ei dispersi sunt
ACTS|5|38|et nunc itaque dico vobis discedite ab hominibus istis et sinite illos quoniam si est ex hominibus consilium hoc aut opus dissolvetur
ACTS|5|39|si vero ex Deo est non poteritis dissolvere eos ne forte et Deo repugnare inveniamini consenserunt autem illi
ACTS|5|40|et convocantes apostolos caesis denuntiaverunt ne loquerentur in nomine Iesu et dimiserunt eos
ACTS|5|41|et illi quidem ibant gaudentes a conspectu concilii quoniam digni habiti sunt pro nomine Iesu contumeliam pati
ACTS|5|42|omni autem die in templo et circa domos non cessabant docentes et evangelizantes Christum Iesum
ACTS|6|1|in diebus autem illis crescente numero discipulorum factus est murmur Graecorum adversus Hebraeos eo quod dispicerentur in ministerio cotidiano viduae eorum
ACTS|6|2|convocantes autem duodecim multitudinem discipulorum dixerunt non est aequum nos derelinquere verbum Dei et ministrare mensis
ACTS|6|3|considerate ergo fratres viros ex vobis boni testimonii septem plenos Spiritu et sapientia quos constituamus super hoc opus
ACTS|6|4|nos vero orationi et ministerio verbi instantes erimus
ACTS|6|5|et placuit sermo coram omni multitudine et elegerunt Stephanum virum plenum fide et Spiritu Sancto et Philippum et Prochorum et Nicanorem et Timonem et Parmenam et Nicolaum advenam Antiochenum
ACTS|6|6|hos statuerunt ante conspectum apostolorum et orantes inposuerunt eis manus
ACTS|6|7|et verbum Dei crescebat et multiplicabatur numerus discipulorum in Hierusalem valde multa etiam turba sacerdotum oboediebat fidei
ACTS|6|8|Stephanus autem plenus gratia et fortitudine faciebat prodigia et signa magna in populo
ACTS|6|9|surrexerunt autem quidam de synagoga quae appellatur Libertinorum et Cyrenensium et Alexandrinorum et eorum qui erant a Cilicia et Asia disputantes cum Stephano
ACTS|6|10|et non poterant resistere sapientiae et Spiritui quo loquebatur
ACTS|6|11|tunc submiserunt viros qui dicerent se audisse eum dicentem verba blasphemiae in Mosen et Deum
ACTS|6|12|commoverunt itaque plebem et seniores et scribas et concurrentes rapuerunt eum et adduxerunt in concilium
ACTS|6|13|et statuerunt testes falsos dicentes homo iste non cessat loqui verba adversus locum sanctum et legem
ACTS|6|14|audivimus enim eum dicentem quoniam Iesus Nazarenus hic destruet locum istum et mutabit traditiones quas tradidit nobis Moses
ACTS|6|15|et intuentes eum omnes qui sedebant in concilio viderunt faciem eius tamquam faciem angeli
ACTS|7|1|dixit autem princeps sacerdotum si haec ita se habent
ACTS|7|2|qui ait viri fratres et patres audite Deus gloriae apparuit patri nostro Abraham cum esset in Mesopotamiam priusquam moraretur in Charram
ACTS|7|3|et dixit ad illum exi de terra tua et de cognatione tua et veni in terram quam tibi monstravero
ACTS|7|4|tunc exiit de terra Chaldeorum et habitavit in Charram et inde postquam mortuus est pater eius transtulit illum in terram istam in qua nunc vos habitatis
ACTS|7|5|et non dedit illi hereditatem in ea nec passum pedis et repromisit dare illi eam in possessionem et semini eius post ipsum cum non haberet filium
ACTS|7|6|locutus est autem Deus quia erit semen eius accola in terra aliena et servituti eos subicient et male tractabunt eos annis quadringentis
ACTS|7|7|et gentem cui servierint iudicabo ego dixit Deus et post haec exibunt et deservient mihi in loco isto
ACTS|7|8|et dedit illi testamentum circumcisionis et sic genuit Isaac et circumcidit eum die octava et Isaac Iacob et Iacob duodecim patriarchas
ACTS|7|9|et patriarchae aemulantes Ioseph vendiderunt in Aegyptum et erat Deus cum eo
ACTS|7|10|et eripuit eum ex omnibus tribulationibus eius et dedit ei gratiam et sapientiam in conspectu Pharaonis regis Aegypti et constituit eum praepositum super Aegyptum et super omnem domum suam
ACTS|7|11|venit autem fames in universam Aegyptum et Chanaan et tribulatio magna et non inveniebant cibos patres nostri
ACTS|7|12|cum audisset autem Iacob esse frumentum in Aegypto misit patres nostros primum
ACTS|7|13|et in secundo cognitus est Ioseph a fratribus suis et manifestatum est Pharaoni genus eius
ACTS|7|14|mittens autem Ioseph accersivit Iacob patrem suum et omnem cognationem in animabus septuaginta quinque
ACTS|7|15|et descendit Iacob in Aegyptum et defunctus est ipse et patres nostri
ACTS|7|16|et translati sunt in Sychem et positi sunt in sepulchro quod emit Abraham pretio argenti a filiis Emmor filii Sychem
ACTS|7|17|cum adpropinquaret autem tempus repromissionis quam confessus erat Deus Abrahae crevit populus et multiplicatus est in Aegypto
ACTS|7|18|quoadusque surrexit rex alius in Aegypto qui non sciebat Ioseph
ACTS|7|19|hic circumveniens genus nostrum adflixit patres ut exponerent infantes suos ne vivificarentur
ACTS|7|20|eodem tempore natus est Moses et fuit gratus Deo qui nutritus est tribus mensibus in domo patris sui
ACTS|7|21|exposito autem illo sustulit eum filia Pharaonis et enutrivit eum sibi in filium
ACTS|7|22|et eruditus est Moses omni sapientia Aegyptiorum et erat potens in verbis et in operibus suis
ACTS|7|23|cum autem impleretur ei quadraginta annorum tempus ascendit in cor eius ut visitaret fratres suos filios Israhel
ACTS|7|24|et cum vidisset quendam iniuriam patientem vindicavit illum et fecit ultionem ei qui iniuriam sustinebat percusso Aegyptio
ACTS|7|25|existimabat autem intellegere fratres quoniam Deus per manum ipsius daret salutem illis at illi non intellexerunt
ACTS|7|26|sequenti vero die apparuit illis litigantibus et reconciliabat eos in pacem dicens viri fratres estis ut quid nocetis alterutrum
ACTS|7|27|qui autem iniuriam faciebat proximo reppulit eum dicens quis te constituit principem et iudicem super nos
ACTS|7|28|numquid interficere me tu vis quemadmodum interfecisti heri Aegyptium
ACTS|7|29|fugit autem Moses in verbo isto et factus est advena in terra Madiam ubi generavit filios duos
ACTS|7|30|et expletis annis quadraginta apparuit illi in deserto montis Sina angelus in igne flammae rubi
ACTS|7|31|Moses autem videns admiratus est visum et accedente illo ut consideraret facta est vox Domini
ACTS|7|32|ego Deus patrum tuorum Deus Abraham et Deus Isaac et Deus Iacob tremefactus autem Moses non audebat considerare
ACTS|7|33|dixit autem illi Dominus solve calciamentum pedum tuorum locus enim in quo stas terra sancta est
ACTS|7|34|videns vidi adflictionem populi mei qui est in Aegypto et gemitum eorum audivi et descendi liberare eos et nunc veni et mittam te in Aegyptum
ACTS|7|35|hunc Mosen quem negaverunt dicentes quis te constituit principem et iudicem hunc Deus principem et redemptorem misit cum manu angeli qui apparuit illi in rubo
ACTS|7|36|hic eduxit illos faciens prodigia et signa in terra Aegypti et in Rubro mari et in deserto annis quadraginta
ACTS|7|37|hic est Moses qui dixit filiis Israhel prophetam vobis suscitabit Deus de fratribus vestris tamquam me
ACTS|7|38|hic est qui fuit in ecclesia in solitudine cum angelo qui loquebatur ei in monte Sina et cum patribus nostris qui accepit verba vitae dare nobis
ACTS|7|39|cui noluerunt oboedire patres nostri sed reppulerunt et aversi sunt cordibus suis in Aegyptum
ACTS|7|40|dicentes ad Aaron fac nobis deos qui praecedant nos Moses enim hic qui eduxit nos de terra Aegypti nescimus quid factum sit ei
ACTS|7|41|et vitulum fecerunt in illis diebus et obtulerunt hostiam simulacro et laetabantur in operibus manuum suarum
ACTS|7|42|convertit autem Deus et tradidit eos servire militiae caeli sicut scriptum est in libro Prophetarum numquid victimas aut hostias obtulistis mihi annis quadraginta in deserto domus Israhel
ACTS|7|43|et suscepistis tabernaculum Moloch et sidus dei vestri Rempham figuras quas fecistis adorare eas et transferam vos trans Babylonem
ACTS|7|44|tabernaculum testimonii fuit patribus nostris in deserto sicut disposuit loquens ad Mosen ut faceret illud secundum formam quam viderat
ACTS|7|45|quod et induxerunt suscipientes patres nostri cum Iesu in possessionem gentium quas expulit Deus a facie patrum nostrorum usque in diebus David
ACTS|7|46|qui invenit gratiam ante Deum et petiit ut inveniret tabernaculum Deo Iacob
ACTS|7|47|Salomon autem aedificavit illi domum
ACTS|7|48|sed non Excelsus in manufactis habitat sicut propheta dicit
ACTS|7|49|caelum mihi sedis est terra autem scabillum pedum meorum quam domum aedificabitis mihi dicit Dominus aut quis locus requietionis meae est
ACTS|7|50|nonne manus mea fecit haec omnia
ACTS|7|51|dura cervice et incircumcisi cordibus et auribus vos semper Spiritui Sancto resistitis sicut patres vestri et vos
ACTS|7|52|quem prophetarum non sunt persecuti patres vestri et occiderunt eos qui praenuntiabant de adventu Iusti cuius vos nunc proditores et homicidae fuistis
ACTS|7|53|qui accepistis legem in dispositionem angelorum et non custodistis
ACTS|7|54|audientes autem haec dissecabantur cordibus suis et stridebant dentibus in eum
ACTS|7|55|cum autem esset plenus Spiritu Sancto intendens in caelum vidit gloriam Dei et Iesum stantem a dextris Dei et ait ecce video caelos apertos et Filium hominis a dextris stantem Dei
ACTS|7|56|exclamantes autem voce magna continuerunt aures suas et impetum fecerunt unianimiter in eum
ACTS|7|57|et eicientes eum extra civitatem lapidabant et testes deposuerunt vestimenta sua secus pedes adulescentis qui vocabatur Saulus
ACTS|7|58|et lapidabant Stephanum invocantem et dicentem Domine Iesu suscipe spiritum meum
ACTS|7|59|positis autem genibus clamavit voce magna Domine ne statuas illis hoc peccatum et cum hoc dixisset obdormivit Saulus autem erat consentiens neci eius
ACTS|8|1|facta est autem in illa die persecutio magna in ecclesia quae erat Hierosolymis et omnes dispersi sunt per regiones Iudaeae et Samariae praeter apostolos
ACTS|8|2|curaverunt autem Stephanum viri timorati et fecerunt planctum magnum super illum
ACTS|8|3|Saulus vero devastabat ecclesiam per domos intrans et trahens viros ac mulieres tradebat in custodiam
ACTS|8|4|igitur qui dispersi erant pertransiebant evangelizantes verbum
ACTS|8|5|Philippus autem descendens in civitatem Samariae praedicabat illis Christum
ACTS|8|6|intendebant autem turbae his quae a Philippo dicebantur unianimiter audientes et videntes signa quae faciebat
ACTS|8|7|multi enim eorum qui habebant spiritus inmundos clamantes voce magna exiebant multi autem paralytici et claudi curati sunt
ACTS|8|8|factum est ergo magnum gaudium in illa civitate
ACTS|8|9|vir autem quidam nomine Simon qui ante fuerat in civitate magus seducens gentem Samariae dicens esse se aliquem magnum
ACTS|8|10|cui auscultabant omnes a minimo usque ad maximum dicentes hic est virtus Dei quae vocatur Magna
ACTS|8|11|adtendebant autem eum propter quod multo tempore magicis suis dementasset eos
ACTS|8|12|cum vero credidissent Philippo evangelizanti de regno Dei et nomine Iesu Christi baptizabantur viri ac mulieres
ACTS|8|13|tunc Simon et ipse credidit et cum baptizatus esset adherebat Philippo videns etiam signa et virtutes maximas fieri stupens admirabatur
ACTS|8|14|cum autem audissent apostoli qui erant Hierosolymis quia recepit Samaria verbum Dei miserunt ad illos Petrum et Iohannem
ACTS|8|15|qui cum venissent oraverunt pro ipsis ut acciperent Spiritum Sanctum
ACTS|8|16|nondum enim in quemquam illorum venerat sed baptizati tantum erant in nomine Domini Iesu
ACTS|8|17|tunc inponebant manus super illos et accipiebant Spiritum Sanctum
ACTS|8|18|cum vidisset autem Simon quia per inpositionem manus apostolorum daretur Spiritus Sanctus obtulit eis pecuniam
ACTS|8|19|dicens date et mihi hanc potestatem ut cuicumque inposuero manus accipiat Spiritum Sanctum Petrus autem dixit ad eum
ACTS|8|20|pecunia tua tecum sit in perditionem quoniam donum Dei existimasti pecunia possideri
ACTS|8|21|non est tibi pars neque sors in sermone isto cor enim tuum non est rectum coram Deo
ACTS|8|22|paenitentiam itaque age ab hac nequitia tua et roga Deum si forte remittatur tibi haec cogitatio cordis tui
ACTS|8|23|in felle enim amaritudinis et obligatione iniquitatis video te esse
ACTS|8|24|respondens autem Simon dixit precamini vos pro me ad Dominum ut nihil veniat super me horum quae dixistis
ACTS|8|25|et illi quidem testificati et locuti verbum Domini rediebant Hierosolymam et multis regionibus Samaritanorum evangelizabant
ACTS|8|26|angelus autem Domini locutus est ad Philippum dicens surge et vade contra meridianum ad viam quae descendit ab Hierusalem in Gazam haec est deserta
ACTS|8|27|et surgens abiit et ecce vir aethiops eunuchus potens Candacis reginae Aethiopum qui erat super omnes gazas eius venerat adorare in Hierusalem
ACTS|8|28|et revertebatur sedens super currum suum legensque prophetam Esaiam
ACTS|8|29|dixit autem Spiritus Philippo accede et adiunge te ad currum istum
ACTS|8|30|adcurrens autem Philippus audivit illum legentem Esaiam prophetam et dixit putasne intellegis quae legis
ACTS|8|31|qui ait et quomodo possum si non aliquis ostenderit mihi rogavitque Philippum ut ascenderet et sederet secum
ACTS|8|32|locus autem scripturae quam legebat erat hic tamquam ovis ad occisionem ductus est et sicut agnus coram tondente se sine voce sic non aperuit os suum
ACTS|8|33|in humilitate iudicium eius sublatum est generationem illius quis enarrabit quoniam tollitur de terra vita eius
ACTS|8|34|respondens autem eunuchus Philippo dixit obsecro te de quo propheta dicit hoc de se an de alio aliquo
ACTS|8|35|aperiens autem Philippus os suum et incipiens ab scriptura ista evangelizavit illi Iesum
ACTS|8|36|et dum irent per viam venerunt ad quandam aquam et ait eunuchus ecce aqua quid prohibet me baptizari
ACTS|8|37|
ACTS|8|38|et iussit stare currum et descenderunt uterque in aquam Philippus et eunuchus et baptizavit eum
ACTS|8|39|cum autem ascendissent de aqua Spiritus Domini rapuit Philippum et amplius non vidit eum eunuchus ibat enim per viam suam gaudens
ACTS|8|40|Philippus autem inventus est in Azoto et pertransiens evangelizabat civitatibus cunctis donec veniret Caesaream
ACTS|9|1|Saulus autem adhuc inspirans minarum et caedis in discipulos Domini accessit ad principem sacerdotum
ACTS|9|2|et petiit ab eo epistulas in Damascum ad synagogas ut si quos invenisset huius viae viros ac mulieres vinctos perduceret in Hierusalem
ACTS|9|3|et cum iter faceret contigit ut adpropinquaret Damasco et subito circumfulsit eum lux de caelo
ACTS|9|4|et cadens in terram audivit vocem dicentem sibi Saule Saule quid me persequeris
ACTS|9|5|qui dixit quis es Domine et ille ego sum Iesus quem tu persequeris
ACTS|9|6|
ACTS|9|7|sed surge et ingredere civitatem et dicetur tibi quid te oporteat facere viri autem illi qui comitabantur cum eo stabant stupefacti audientes quidem vocem neminem autem videntes
ACTS|9|8|surrexit autem Saulus de terra apertisque oculis nihil videbat ad manus autem illum trahentes introduxerunt Damascum
ACTS|9|9|et erat tribus diebus non videns et non manducavit neque bibit
ACTS|9|10|erat autem quidam discipulus Damasci nomine Ananias et dixit ad illum in visu Dominus Anania at ille ait ecce ego Domine
ACTS|9|11|et Dominus ad illum surgens vade in vicum qui vocatur Rectus et quaere in domo Iudae Saulum nomine Tarsensem ecce enim orat
ACTS|9|12|et vidit virum Ananiam nomine introeuntem et inponentem sibi manus ut visum recipiat
ACTS|9|13|respondit autem Ananias Domine audivi a multis de viro hoc quanta mala sanctis tuis fecerit in Hierusalem
ACTS|9|14|et hic habet potestatem a principibus sacerdotum alligandi omnes qui invocant nomen tuum
ACTS|9|15|dixit autem ad eum Dominus vade quoniam vas electionis est mihi iste ut portet nomen meum coram gentibus et regibus et filiis Israhel
ACTS|9|16|ego enim ostendam illi quanta oporteat eum pro nomine meo pati
ACTS|9|17|et abiit Ananias et introivit in domum et inponens ei manus dixit Saule frater Dominus misit me Iesus qui apparuit tibi in via qua veniebas ut videas et implearis Spiritu Sancto
ACTS|9|18|et confestim ceciderunt ab oculis eius tamquam squamae et visum recepit et surgens baptizatus est
ACTS|9|19|et cum accepisset cibum confortatus est fuit autem cum discipulis qui erant Damasci per dies aliquot
ACTS|9|20|et continuo in synagogis praedicabat Iesum quoniam hic est Filius Dei
ACTS|9|21|stupebant autem omnes qui audiebant et dicebant nonne hic est qui expugnabat in Hierusalem eos qui invocabant nomen istud et huc ad hoc venit ut vinctos illos duceret ad principes sacerdotum
ACTS|9|22|Saulus autem magis convalescebat et confundebat Iudaeos qui habitabant Damasci adfirmans quoniam hic est Christus
ACTS|9|23|cum implerentur autem dies multi consilium fecerunt Iudaei ut eum interficerent
ACTS|9|24|notae autem factae sunt Saulo insidiae eorum custodiebant autem et portas die ac nocte ut eum interficerent
ACTS|9|25|accipientes autem discipuli eius nocte per murum dimiserunt eum submittentes in sporta
ACTS|9|26|cum autem venisset in Hierusalem temptabat iungere se discipulis et omnes timebant eum non credentes quia esset discipulus
ACTS|9|27|Barnabas autem adprehensum illum duxit ad apostolos et narravit illis quomodo in via vidisset Dominum et quia locutus est ei et quomodo in Damasco fiducialiter egerit in nomine Iesu
ACTS|9|28|et erat cum illis intrans et exiens in Hierusalem et fiducialiter agens in nomine Domini
ACTS|9|29|loquebatur quoque et disputabat cum Graecis illi autem quaerebant occidere eum
ACTS|9|30|quod cum cognovissent fratres deduxerunt eum Caesaream et dimiserunt Tarsum
ACTS|9|31|ecclesia quidem per totam Iudaeam et Galilaeam et Samariam habebat pacem et aedificabatur ambulans in timore Domini et consolatione Sancti Spiritus replebatur
ACTS|9|32|factum est autem Petrum dum pertransiret universos devenire et ad sanctos qui habitabant Lyddae
ACTS|9|33|invenit autem ibi hominem quendam nomine Aeneam ab annis octo iacentem in grabatto qui erat paralyticus
ACTS|9|34|et ait illi Petrus Aeneas sanat te Iesus Christus surge et sterne tibi et continuo surrexit
ACTS|9|35|et viderunt illum omnes qui habitabant Lyddae et Saronae qui conversi sunt ad Dominum
ACTS|9|36|in Ioppe autem fuit quaedam discipula nomine Tabitas quae interpretata dicitur Dorcas haec erat plena operibus bonis et elemosynis quas faciebat
ACTS|9|37|factum est autem in diebus illis ut infirmata moreretur quam cum lavissent posuerunt eam in cenaculo
ACTS|9|38|cum autem prope esset Lydda ab Ioppe discipuli audientes quia Petrus esset in ea miserunt duos viros ad eum rogantes ne pigriteris venire usque ad nos
ACTS|9|39|exsurgens autem Petrus venit cum illis et cum advenisset duxerunt illum in cenaculum et circumsteterunt illum omnes viduae flentes et ostendentes tunicas et vestes quas faciebat illis Dorcas
ACTS|9|40|eiectis autem omnibus foras Petrus ponens genua oravit et conversus ad corpus dixit Tabita surge at illa aperuit oculos suos et viso Petro resedit
ACTS|9|41|dans autem illi manum erexit eam et cum vocasset sanctos et viduas adsignavit eam vivam
ACTS|9|42|notum autem factum est per universam Ioppen et crediderunt multi in Domino
ACTS|9|43|factum est autem ut dies multos moraretur in Ioppe apud quendam Simonem coriarium
ACTS|10|1|vir autem quidam erat in Caesarea nomine Cornelius centurio cohortis quae dicitur Italica
ACTS|10|2|religiosus et timens Deum cum omni domo sua faciens elemosynas multas plebi et deprecans Deum semper
ACTS|10|3|vidit in visu manifeste quasi hora nona diei angelum Dei introeuntem ad se et dicentem sibi Corneli
ACTS|10|4|at ille intuens eum timore correptus dixit quid est domine dixit autem illi orationes tuae et elemosynae tuae ascenderunt in memoriam in conspectu Dei
ACTS|10|5|et nunc mitte viros in Ioppen et accersi Simonem quendam qui cognominatur Petrus
ACTS|10|6|hic hospitatur apud Simonem quendam coriarium cuius est domus iuxta mare
ACTS|10|7|et cum discessisset angelus qui loquebatur illi vocavit duos domesticos suos et militem metuentem Dominum ex his qui illi parebant
ACTS|10|8|quibus cum narrasset omnia misit illos in Ioppen
ACTS|10|9|postera autem die iter illis facientibus et adpropinquantibus civitati ascendit Petrus in superiora ut oraret circa horam sextam
ACTS|10|10|et cum esuriret voluit gustare parantibus autem eis cecidit super eum mentis excessus
ACTS|10|11|et videt caelum apertum et descendens vas quoddam velut linteum magnum quattuor initiis submitti de caelo in terram
ACTS|10|12|in quo erant omnia quadrupedia et serpentia terrae et volatilia caeli
ACTS|10|13|et facta est vox ad eum surge Petre et occide et manduca
ACTS|10|14|ait autem Petrus absit Domine quia numquam manducavi omne commune et inmundum
ACTS|10|15|et vox iterum secundo ad eum quae Deus purificavit ne tu commune dixeris
ACTS|10|16|hoc autem factum est per ter et statim receptum est vas in caelum
ACTS|10|17|et dum intra se haesitaret Petrus quidnam esset visio quam vidisset ecce viri qui missi erant a Cornelio inquirentes domum Simonis adstiterunt ad ianuam
ACTS|10|18|et cum vocassent interrogabant si Simon qui cognominatur Petrus illic haberet hospitium
ACTS|10|19|Petro autem cogitante de visione dixit Spiritus ei ecce viri tres quaerunt te
ACTS|10|20|surge itaque et descende et vade cum eis nihil dubitans quia ego misi illos
ACTS|10|21|descendens autem Petrus ad viros dixit ecce ego sum quem quaeritis quae causa est propter quam venistis
ACTS|10|22|qui dixerunt Cornelius centurio vir iustus et timens Deum et testimonium habens ab universa gente Iudaeorum responsum accepit ab angelo sancto accersire te in domum suam et audire verba abs te
ACTS|10|23|introducens igitur eos recepit hospitio sequenti autem die surgens profectus est cum eis et quidam ex fratribus ab Ioppe comitati sunt eum
ACTS|10|24|altera autem die introivit Caesaream Cornelius vero expectabat illos convocatis cognatis suis et necessariis amicis
ACTS|10|25|et factum est cum introisset Petrus obvius ei Cornelius et procidens ad pedes adoravit
ACTS|10|26|Petrus vero levavit eum dicens surge et ego ipse homo sum
ACTS|10|27|et loquens cum illo intravit et invenit multos qui convenerant
ACTS|10|28|dixitque ad illos vos scitis quomodo abominatum sit viro iudaeo coniungi aut accedere ad alienigenam et mihi ostendit Deus neminem communem aut inmundum dicere hominem
ACTS|10|29|propter quod sine dubitatione veni accersitus interrogo ergo quam ob causam accersistis me
ACTS|10|30|et Cornelius ait a nudius quartana die usque in hanc horam orans eram hora nona in domo mea et ecce vir stetit ante me in veste candida et ait
ACTS|10|31|Corneli exaudita est oratio tua et elemosynae tuae commemoratae sunt in conspectu Dei
ACTS|10|32|mitte ergo in Ioppen et accersi Simonem qui cognominatur Petrus hic hospitatur in domo Simonis coriarii iuxta mare
ACTS|10|33|confestim igitur misi ad te et tu bene fecisti veniendo nunc ergo omnes nos in conspectu tuo adsumus audire omnia quaecumque tibi praecepta sunt a Domino
ACTS|10|34|aperiens autem Petrus os dixit in veritate conperi quoniam non est personarum acceptor Deus
ACTS|10|35|sed in omni gente qui timet eum et operatur iustitiam acceptus est illi
ACTS|10|36|verbum misit filiis Israhel adnuntians pacem per Iesum Christum hic est omnium Dominus
ACTS|10|37|vos scitis quod factum est verbum per universam Iudaeam incipiens enim a Galilaea post baptismum quod praedicavit Iohannes
ACTS|10|38|Iesum a Nazareth quomodo unxit eum Deus Spiritu Sancto et virtute qui pertransivit benefaciendo et sanando omnes oppressos a diabolo quoniam Deus erat cum illo
ACTS|10|39|et nos testes sumus omnium quae fecit in regione Iudaeorum et Hierusalem quem et occiderunt suspendentes in ligno
ACTS|10|40|hunc Deus suscitavit tertia die et dedit eum manifestum fieri
ACTS|10|41|non omni populo sed testibus praeordinatis a Deo nobis qui manducavimus et bibimus cum illo postquam resurrexit a mortuis
ACTS|10|42|et praecepit nobis praedicare populo et testificari quia ipse est qui constitutus est a Deo iudex vivorum et mortuorum
ACTS|10|43|huic omnes prophetae testimonium perhibent remissionem peccatorum accipere per nomen eius omnes qui credunt in eum
ACTS|10|44|adhuc loquente Petro verba haec cecidit Spiritus Sanctus super omnes qui audiebant verbum
ACTS|10|45|et obstipuerunt ex circumcisione fideles qui venerant cum Petro quia et in nationes gratia Spiritus Sancti effusa est
ACTS|10|46|audiebant enim illos loquentes linguis et magnificantes Deum
ACTS|10|47|tunc respondit Petrus numquid aquam quis prohibere potest ut non baptizentur hii qui Spiritum Sanctum acceperunt sicut et nos
ACTS|10|48|et iussit eos in nomine Iesu Christi baptizari tunc rogaverunt eum ut maneret aliquot diebus
ACTS|11|1|audierunt autem apostoli et fratres qui erant in Iudaea quoniam et gentes receperunt verbum Dei
ACTS|11|2|cum ascendisset autem Petrus in Hierosolymam disceptabant adversus illum qui erant ex circumcisione
ACTS|11|3|dicentes quare introisti ad viros praeputium habentes et manducasti cum illis
ACTS|11|4|incipiens autem Petrus exponebat illis ordinem dicens
ACTS|11|5|ego eram in civitate Ioppe orans et vidi in excessu mentis visionem descendens vas quoddam velut linteum magnum quattuor initiis submitti de caelo et venit usque ad me
ACTS|11|6|in quod intuens considerabam et vidi quadrupedia terrae et bestias et reptilia et volatilia caeli
ACTS|11|7|audivi autem et vocem dicentem mihi surgens Petre occide et manduca
ACTS|11|8|dixi autem nequaquam Domine quia commune aut inmundum numquam introivit in os meum
ACTS|11|9|respondit autem vox secundo de caelo quae Deus mundavit tu ne commune dixeris
ACTS|11|10|hoc autem factum est per ter et recepta sunt rursum omnia in caelum
ACTS|11|11|et ecce confestim tres viri adstiterunt in domo in qua eram missi a Caesarea ad me
ACTS|11|12|dixit autem Spiritus mihi ut irem cum illis nihil haesitans venerunt autem mecum et sex fratres isti et ingressi sumus in domum viri
ACTS|11|13|narravit autem nobis quomodo vidisset angelum in domo sua stantem et dicentem sibi mitte in Ioppen et accersi Simonem qui cognominatur Petrus
ACTS|11|14|qui loquetur tibi verba in quibus salvus eris tu et universa domus tua
ACTS|11|15|cum autem coepissem loqui decidit Spiritus Sanctus super eos sicut et in nos in initio
ACTS|11|16|recordatus sum autem verbi Domini sicut dicebat Iohannes quidem baptizavit aqua vos autem baptizabimini Spiritu Sancto
ACTS|11|17|si ergo eandem gratiam dedit illis Deus sicut et nobis qui credidimus in Dominum Iesum Christum ego quis eram qui possem prohibere Deum
ACTS|11|18|his auditis tacuerunt et glorificaverunt Deum dicentes ergo et gentibus Deus paenitentiam ad vitam dedit
ACTS|11|19|et illi quidem qui dispersi fuerant a tribulatione quae facta fuerat sub Stephano perambulaverunt usque Foenicen et Cyprum et Antiochiam nemini loquentes verbum nisi solis Iudaeis
ACTS|11|20|erant autem quidam ex eis viri cyprii et cyrenei qui cum introissent Antiochiam loquebantur et ad Graecos adnuntiantes Dominum Iesum
ACTS|11|21|et erat manus Domini cum eis multusque numerus credentium conversus est ad Dominum
ACTS|11|22|pervenit autem sermo ad aures ecclesiae quae erat Hierosolymis super istis et miserunt Barnaban usque Antiochiam
ACTS|11|23|qui cum pervenisset et vidisset gratiam Dei gavisus est et hortabatur omnes proposito cordis permanere in Domino
ACTS|11|24|quia erat vir bonus et plenus Spiritu Sancto et fide et adposita est turba multa Domino
ACTS|11|25|profectus est autem Tarsum ut quaereret Saulum quem cum invenisset perduxit Antiochiam
ACTS|11|26|et annum totum conversati sunt in ecclesia et docuerunt turbam multam ita ut cognominarentur primum Antiochiae discipuli Christiani
ACTS|11|27|in his autem diebus supervenerunt ab Hierosolymis prophetae Antiochiam
ACTS|11|28|et surgens unus ex eis nomine Agabus significabat per Spiritum famem magnam futuram in universo orbe terrarum quae facta est sub Claudio
ACTS|11|29|discipuli autem prout quis habebat proposuerunt singuli eorum in ministerium mittere habitantibus in Iudaea fratribus
ACTS|11|30|quod et fecerunt mittentes ad seniores per manus Barnabae et Sauli
ACTS|12|1|eodem autem tempore misit Herodes rex manus ut adfligeret quosdam de ecclesia
ACTS|12|2|occidit autem Iacobum fratrem Iohannis gladio
ACTS|12|3|videns autem quia placeret Iudaeis adposuit adprehendere et Petrum erant autem dies azymorum
ACTS|12|4|quem cum adprehendisset misit in carcerem tradens quattuor quaternionibus militum custodire eum volens post pascha producere eum populo
ACTS|12|5|et Petrus quidem servabatur in carcere oratio autem fiebat sine intermissione ab ecclesia ad Deum pro eo
ACTS|12|6|cum autem producturus eum esset Herodes in ipsa nocte erat Petrus dormiens inter duos milites vinctus catenis duabus et custodes ante ostium custodiebant carcerem
ACTS|12|7|et ecce angelus Domini adstitit et lumen refulsit in habitaculo percussoque latere Petri suscitavit eum dicens surge velociter et ceciderunt catenae de manibus eius
ACTS|12|8|dixit autem angelus ad eum praecingere et calcia te gallicas tuas et fecit sic et dixit illi circumda tibi vestimentum tuum et sequere me
ACTS|12|9|et exiens sequebatur et nesciebat quia verum est quod fiebat per angelum aestimabat autem se visum videre
ACTS|12|10|transeuntes autem primam et secundam custodiam venerunt ad portam ferream quae ducit ad civitatem quae ultro aperta est eis et exeuntes processerunt vicum unum et continuo discessit angelus ab eo
ACTS|12|11|et Petrus ad se reversus dixit nunc scio vere quia misit Dominus angelum suum et eripuit me de manu Herodis et de omni expectatione plebis Iudaeorum
ACTS|12|12|consideransque venit ad domum Mariae matris Iohannis qui cognominatus est Marcus ubi erant multi congregati et orantes
ACTS|12|13|pulsante autem eo ostium ianuae processit puella ad audiendum nomine Rhode
ACTS|12|14|et ut cognovit vocem Petri prae gaudio non aperuit ianuam sed intro currens nuntiavit stare Petrum ante ianuam
ACTS|12|15|at illi dixerunt ad eam insanis illa autem adfirmabat sic se habere illi autem dicebant angelus eius est
ACTS|12|16|Petrus autem perseverabat pulsans cum autem aperuissent viderunt eum et obstipuerunt
ACTS|12|17|annuens autem eis manu ut tacerent enarravit quomodo Dominus eduxisset eum de carcere dixitque nuntiate Iacobo et fratribus haec et egressus abiit in alium locum
ACTS|12|18|facta autem die erat non parva turbatio inter milites quidnam de Petro factum esset
ACTS|12|19|Herodes autem cum requisisset eum et non invenisset inquisitione facta de custodibus iussit eos duci descendensque a Iudaea in Caesaream ibi commoratus est
ACTS|12|20|erat autem iratus Tyriis et Sidoniis at illi unianimes venerunt ad eum et persuaso Blasto qui erat super cubiculum regis postulabant pacem eo quod alerentur regiones eorum ab illo
ACTS|12|21|statuto autem die Herodes vestitus veste regia sedit pro tribunali et contionabatur ad eos
ACTS|12|22|populus autem adclamabat dei voces et non hominis
ACTS|12|23|confestim autem percussit eum angelus Domini eo quod non dedisset honorem Deo et consumptus a vermibus exspiravit
ACTS|12|24|verbum autem Domini crescebat et multiplicabatur
ACTS|12|25|Barnabas autem et Saulus reversi sunt ab Hierosolymis expleto ministerio adsumpto Iohanne qui cognominatus est Marcus
ACTS|13|1|erant autem in ecclesia quae erat Antiochiae prophetae et doctores in quibus Barnabas et Symeon qui vocabatur Niger et Lucius Cyrenensis et Manaen qui erat Herodis tetrarchae conlactaneus et Saulus
ACTS|13|2|ministrantibus autem illis Domino et ieiunantibus dixit Spiritus Sanctus separate mihi Barnaban et Saulum in opus quod adsumpsi eos
ACTS|13|3|tunc ieiunantes et orantes inponentesque eis manus dimiserunt illos
ACTS|13|4|et ipsi quidem missi ab Spiritu Sancto abierunt Seleuciam et inde navigaverunt Cyprum
ACTS|13|5|et cum venissent Salamina praedicabant verbum Dei in synagogis Iudaeorum habebant autem et Iohannem in ministerio
ACTS|13|6|et cum perambulassent universam insulam usque Paphum invenerunt quendam virum magum pseudoprophetam Iudaeum cui nomen erat Bariesu
ACTS|13|7|qui erat cum proconsule Sergio Paulo viro prudente hic accitis Barnaba et Saulo desiderabat audire verbum Dei
ACTS|13|8|resistebat autem illis Elymas magus sic enim interpretatur nomen eius quaerens avertere proconsulem a fide
ACTS|13|9|Saulus autem qui et Paulus repletus Spiritu Sancto intuens in eum
ACTS|13|10|dixit o plene omni dolo et omni fallacia fili diaboli inimice omnis iustitiae non desinis subvertere vias Domini rectas
ACTS|13|11|et nunc ecce manus Domini super te et eris caecus non videns solem usque ad tempus et confestim cecidit in eum caligo et tenebrae et circumiens quaerebat qui ei manum daret
ACTS|13|12|tunc proconsul cum vidisset factum credidit admirans super doctrinam Domini
ACTS|13|13|et cum a Papho navigassent Paulus et qui cum eo venerunt Pergen Pamphiliae Iohannes autem discedens ab eis reversus est Hierosolymam
ACTS|13|14|illi vero pertranseuntes Pergen venerunt Antiochiam Pisidiae et ingressi synagogam die sabbatorum sederunt
ACTS|13|15|post lectionem autem legis et prophetarum miserunt principes synagogae ad eos dicentes viri fratres si quis est in vobis sermo exhortationis ad plebem dicite
ACTS|13|16|surgens autem Paulus et manu silentium indicens ait viri israhelitae et qui timetis Deum audite
ACTS|13|17|Deus plebis Israhel elegit patres nostros et plebem exaltavit cum essent incolae in terra Aegypti et in brachio excelso eduxit eos ex ea
ACTS|13|18|et per quadraginta annorum tempus mores eorum sustinuit in deserto
ACTS|13|19|et destruens gentes septem in terra Chanaan sorte distribuit eis terram eorum
ACTS|13|20|quasi post quadringentos et quinquaginta annos et post haec dedit iudices usque ad Samuhel prophetam
ACTS|13|21|et exinde postulaverunt regem et dedit illis Deus Saul filium Cis virum de tribu Beniamin annis quadraginta
ACTS|13|22|et amoto illo suscitavit illis David regem cui et testimonium perhibens dixit inveni David filium Iesse virum secundum cor meum qui faciet omnes voluntates meas
ACTS|13|23|huius Deus ex semine secundum promissionem eduxit Israhel salvatorem Iesum
ACTS|13|24|praedicante Iohanne ante faciem adventus eius baptismum paenitentiae omni populo Israhel
ACTS|13|25|cum impleret autem Iohannes cursum suum dicebat quem me arbitramini esse non sum ego sed ecce venit post me cuius non sum dignus calciamenta pedum solvere
ACTS|13|26|viri fratres filii generis Abraham et qui in vobis timent Deum vobis verbum salutis huius missum est
ACTS|13|27|qui enim habitabant Hierusalem et principes eius hunc ignorantes et voces prophetarum quae per omne sabbatum leguntur iudicantes impleverunt
ACTS|13|28|et nullam causam mortis invenientes in eum petierunt a Pilato ut interficerent eum
ACTS|13|29|cumque consummassent omnia quae de eo scripta erant deponentes eum de ligno posuerunt in monumento
ACTS|13|30|Deus vero suscitavit eum a mortuis qui visus est per dies multos his
ACTS|13|31|qui simul ascenderant cum eo de Galilaea in Hierusalem qui usque nunc sunt testes eius ad plebem
ACTS|13|32|et nos vobis adnuntiamus ea quae ad patres nostros repromissio facta est
ACTS|13|33|quoniam hanc Deus adimplevit filiis nostris resuscitans Iesum sicut et in psalmo secundo scriptum est Filius meus es tu ego hodie genui te
ACTS|13|34|quod autem suscitaverit eum a mortuis amplius iam non reversurum in corruptionem ita dixit quia dabo vobis sancta David fidelia
ACTS|13|35|ideoque et alias dicit non dabis Sanctum tuum videre corruptionem
ACTS|13|36|David enim sua generatione cum administrasset voluntati Dei dormivit et adpositus est ad patres suos et vidit corruptionem
ACTS|13|37|quem vero Deus suscitavit non vidit corruptionem
ACTS|13|38|notum igitur sit vobis viri fratres quia per hunc vobis remissio peccatorum adnuntiatur ab omnibus quibus non potuistis in lege Mosi iustificari
ACTS|13|39|in hoc omnis qui credit iustificatur
ACTS|13|40|videte ergo ne superveniat quod dictum est in prophetis
ACTS|13|41|videte contemptores et admiramini et disperdimini quia opus operor ego in diebus vestris opus quod non credetis si quis enarraverit vobis
ACTS|13|42|exeuntibus autem illis rogabant ut sequenti sabbato loquerentur sibi verba haec
ACTS|13|43|cumque dimissa esset synagoga secuti sunt multi Iudaeorum et colentium advenarum Paulum et Barnaban qui loquentes suadebant eis ut permanerent in gratia Dei
ACTS|13|44|sequenti vero sabbato paene universa civitas convenit audire verbum Domini
ACTS|13|45|videntes autem turbas Iudaei repleti sunt zelo et contradicebant his quae a Paulo dicebantur blasphemantes
ACTS|13|46|tunc constanter Paulus et Barnabas dixerunt vobis oportebat primum loqui verbum Dei sed quoniam repellitis illud et indignos vos iudicastis aeternae vitae ecce convertimur ad gentes
ACTS|13|47|sic enim praecepit nobis Dominus posui te in lumen gentibus ut sis in salutem usque ad extremum terrae
ACTS|13|48|audientes autem gentes gavisae sunt et glorificabant verbum Domini et crediderunt quotquot erant praeordinati ad vitam aeternam
ACTS|13|49|disseminabatur autem verbum Domini per universam regionem
ACTS|13|50|Iudaei autem concitaverunt religiosas mulieres et honestas et primos civitatis et excitaverunt persecutionem in Paulum et Barnaban et eiecerunt eos de finibus suis
ACTS|13|51|at illi excusso pulvere pedum in eos venerunt Iconium
ACTS|13|52|discipuli quoque replebantur gaudio et Spiritu Sancto
ACTS|14|1|factum est autem Iconii ut simul introirent synagogam Iudaeorum et loquerentur ita ut crederet Iudaeorum et Graecorum copiosa multitudo
ACTS|14|2|qui vero increduli fuerunt Iudaei suscitaverunt et ad iracundiam concitaverunt animas gentium adversus fratres
ACTS|14|3|multo igitur tempore demorati sunt fiducialiter agentes in Domino testimonium perhibente verbo gratiae suae dante signa et prodigia fieri per manus eorum
ACTS|14|4|divisa est autem multitudo civitatis et quidam quidem erant cum Iudaeis quidam vero cum apostolis
ACTS|14|5|cum autem factus esset impetus gentilium et Iudaeorum cum principibus suis ut contumeliis adficerent et lapidarent eos
ACTS|14|6|intellegentes confugerunt ad civitates Lycaoniae Lystram et Derben et universam in circuitu regionem et ibi evangelizantes erant
ACTS|14|7|et quidam vir in Lystris infirmus pedibus sedebat claudus ex utero matris suae qui numquam ambulaverat
ACTS|14|8|hic audivit Paulum loquentem qui intuitus eum et videns quia haberet fidem ut salvus fieret
ACTS|14|9|dixit magna voce surge super pedes tuos rectus et exilivit et ambulabat
ACTS|14|10|turbae autem cum vidissent quod fecerat Paulus levaverunt vocem suam lycaonice dicentes dii similes facti hominibus descenderunt ad nos
ACTS|14|11|et vocabant Barnaban Iovem Paulum vero Mercurium quoniam ipse erat dux verbi
ACTS|14|12|sacerdos quoque Iovis qui erat ante civitatem tauros et coronas ante ianuas adferens cum populis volebat sacrificare
ACTS|14|13|quod ubi audierunt apostoli Barnabas et Paulus conscissis tunicis suis exilierunt in turbas clamantes
ACTS|14|14|et dicentes viri quid haec facitis et nos mortales sumus similes vobis homines adnuntiantes vobis ab his vanis converti ad Deum vivum qui fecit caelum et terram et mare et omnia quae in eis sunt
ACTS|14|15|qui in praeteritis generationibus dimisit omnes gentes ingredi in vias suas
ACTS|14|16|et quidem non sine testimonio semet ipsum reliquit benefaciens de caelo dans pluvias et tempora fructifera implens cibo et laetitia corda vestra
ACTS|14|17|et haec dicentes vix sedaverunt turbas ne sibi immolarent
ACTS|14|18|supervenerunt autem quidam ab Antiochia et Iconio Iudaei et persuasis turbis lapidantesque Paulum traxerunt extra civitatem aestimantes eum mortuum esse
ACTS|14|19|circumdantibus autem eum discipulis surgens intravit civitatem et postera die profectus est cum Barnaba in Derben
ACTS|14|20|cumque evangelizassent civitati illi et docuissent multos reversi sunt Lystram et Iconium et Antiochiam
ACTS|14|21|confirmantes animas discipulorum exhortantes ut permanerent in fide et quoniam per multas tribulationes oportet nos intrare in regnum Dei
ACTS|14|22|et cum constituissent illis per singulas ecclesias presbyteros et orassent cum ieiunationibus commendaverunt eos Domino in quem crediderunt
ACTS|14|23|transeuntesque Pisidiam venerunt Pamphiliam
ACTS|14|24|et loquentes in Pergen verbum Domini descenderunt in Attaliam
ACTS|14|25|et inde navigaverunt Antiochiam unde erant traditi gratiae Dei in opus quod conpleverunt
ACTS|14|26|cum autem venissent et congregassent ecclesiam rettulerunt quanta fecisset Deus cum illis quia aperuisset gentibus ostium fidei
ACTS|14|27|morati sunt autem tempus non modicum cum discipulis
ACTS|15|1|et quidam descendentes de Iudaea docebant fratres quia nisi circumcidamini secundum morem Mosi non potestis salvi fieri
ACTS|15|2|facta ergo seditione non minima Paulo et Barnabae adversum illos statuerunt ut ascenderent Paulus et Barnabas et quidam alii ex illis ad apostolos et presbyteros in Hierusalem super hac quaestione
ACTS|15|3|illi igitur deducti ab ecclesia pertransiebant Foenicen et Samariam narrantes conversionem gentium et faciebant gaudium magnum omnibus fratribus
ACTS|15|4|cum autem venissent Hierosolymam suscepti sunt ab ecclesia et ab apostolis et senioribus adnuntiantes quanta Deus fecisset cum illis
ACTS|15|5|surrexerunt autem quidam de heresi Pharisaeorum qui crediderant dicentes quia oportet circumcidi eos praecipere quoque servare legem Mosi
ACTS|15|6|conveneruntque apostoli et seniores videre de verbo hoc
ACTS|15|7|cum autem magna conquisitio fieret surgens Petrus dixit ad eos viri fratres vos scitis quoniam ab antiquis diebus in nobis elegit Deus per os meum audire gentes verbum evangelii et credere
ACTS|15|8|et qui novit corda Deus testimonium perhibuit dans illis Spiritum Sanctum sicut et nobis
ACTS|15|9|et nihil discrevit inter nos et illos fide purificans corda eorum
ACTS|15|10|nunc ergo quid temptatis Deum inponere iugum super cervicem discipulorum quod neque patres nostri neque nos portare potuimus
ACTS|15|11|sed per gratiam Domini Iesu credimus salvari quemadmodum et illi
ACTS|15|12|tacuit autem omnis multitudo et audiebant Barnaban et Paulum narrantes quanta fecisset Deus signa et prodigia in gentibus per eos
ACTS|15|13|et postquam tacuerunt respondit Iacobus dicens viri fratres audite me
ACTS|15|14|Simeon narravit quemadmodum primum Deus visitavit sumere ex gentibus populum nomini suo
ACTS|15|15|et huic concordant verba prophetarum sicut scriptum est
ACTS|15|16|post haec revertar et aedificabo tabernaculum David quod decidit et diruta eius reaedificabo et erigam illud
ACTS|15|17|ut requirant ceteri hominum Dominum et omnes gentes super quas invocatum est nomen meum dicit Dominus faciens haec
ACTS|15|18|notum a saeculo est Domino opus suum
ACTS|15|19|propter quod ego iudico non inquietari eos qui ex gentibus convertuntur ad Deum
ACTS|15|20|sed scribere ad eos ut abstineant se a contaminationibus simulacrorum et fornicatione et suffocatis et sanguine
ACTS|15|21|Moses enim a temporibus antiquis habet in singulis civitatibus qui eum praedicent in synagogis ubi per omne sabbatum legitur
ACTS|15|22|tunc placuit apostolis et senioribus cum omni ecclesia eligere viros ex eis et mittere Antiochiam cum Paulo et Barnaba Iudam qui cognominatur Barsabban et Silam viros primos in fratribus
ACTS|15|23|scribentes per manus eorum apostoli et seniores fratres his qui sunt Antiochiae et Syriae et Ciliciae fratribus ex gentibus salutem
ACTS|15|24|quoniam audivimus quia quidam ex nobis exeuntes turbaverunt vos verbis evertentes animas vestras quibus non mandavimus
ACTS|15|25|placuit nobis collectis in unum eligere viros et mittere ad vos cum carissimis nostris Barnaba et Paulo
ACTS|15|26|hominibus qui tradiderunt animas suas pro nomine Domini nostri Iesu Christi
ACTS|15|27|misimus ergo Iudam et Silam qui et ipsi vobis verbis referent eadem
ACTS|15|28|visum est enim Spiritui Sancto et nobis nihil ultra inponere vobis oneris quam haec necessario
ACTS|15|29|ut abstineatis vos ab immolatis simulacrorum et sanguine suffocato et fornicatione a quibus custodientes vos bene agetis valete
ACTS|15|30|illi igitur dimissi descenderunt Antiochiam et congregata multitudine tradiderunt epistulam
ACTS|15|31|quam cum legissent gavisi sunt super consolatione
ACTS|15|32|Iudas autem et Silas et ipsi cum essent prophetae verbo plurimo consolati sunt fratres et confirmaverunt
ACTS|15|33|facto autem ibi tempore dimissi sunt cum pace a fratribus ad eos qui miserant illos
ACTS|15|34|
ACTS|15|35|Paulus autem et Barnabas demorabantur Antiochiae docentes et evangelizantes cum aliis pluribus verbum Domini
ACTS|15|36|post aliquot autem dies dixit ad Barnaban Paulus revertentes visitemus fratres per universas civitates in quibus praedicavimus verbum Domini quomodo se habeant
ACTS|15|37|Barnabas autem volebat secum adsumere et Iohannem qui cognominatur Marcus
ACTS|15|38|Paulus autem rogabat eum qui discessisset ab eis a Pamphilia et non isset cum eis in opus non debere recipi eum
ACTS|15|39|facta est autem dissensio ita ut discederent ab invicem et Barnabas adsumpto Marco navigaret Cyprum
ACTS|15|40|Paulus vero electo Sila profectus est traditus gratiae Domini a fratribus
ACTS|15|41|perambulabat autem Syriam et Ciliciam confirmans ecclesias
ACTS|16|1|pervenit autem in Derben et Lystram et ecce discipulus quidam erat ibi nomine Timotheus filius mulieris iudaeae fidelis patre gentili
ACTS|16|2|huic testimonium reddebant qui in Lystris erant et Iconii fratres
ACTS|16|3|hunc voluit Paulus secum proficisci et adsumens circumcidit eum propter Iudaeos qui erant in illis locis sciebant enim omnes quod pater eius gentilis esset
ACTS|16|4|cum autem pertransirent civitates tradebant eis custodire dogmata quae erant decreta ab apostolis et senioribus qui essent Hierosolymis
ACTS|16|5|et ecclesiae quidem confirmabantur fide et abundabant numero cotidie
ACTS|16|6|transeuntes autem Frygiam et Galatiae regionem vetati sunt a Sancto Spiritu loqui verbum in Asia
ACTS|16|7|cum venissent autem in Mysiam temptabant ire Bithyniam et non permisit eos Spiritus Iesu
ACTS|16|8|cum autem pertransissent Mysiam descenderunt Troadem
ACTS|16|9|et visio per noctem Paulo ostensa est vir macedo quidam erat stans et deprecans eum et dicens transiens in Macedoniam adiuva nos
ACTS|16|10|ut autem visum vidit statim quaesivimus proficisci in Macedoniam certi facti quia vocasset nos Deus evangelizare eis
ACTS|16|11|navigantes autem a Troade recto cursu venimus Samothraciam et sequenti die Neapolim
ACTS|16|12|et inde Philippis quae est prima partis Macedoniae civitas colonia eramus autem in hac urbe diebus aliquot conferentes
ACTS|16|13|die autem sabbatorum egressi sumus foras portam iuxta flumen ubi videbatur oratio esse et sedentes loquebamur mulieribus quae convenerant
ACTS|16|14|et quaedam mulier nomine Lydia purpuraria civitatis Thyatirenorum colens Deum audivit cuius Dominus aperuit cor intendere his quae dicebantur a Paulo
ACTS|16|15|cum autem baptizata esset et domus eius deprecata est dicens si iudicastis me fidelem Domino esse introite in domum meam et manete et coegit nos
ACTS|16|16|factum est autem euntibus nobis ad orationem puellam quandam habentem spiritum pythonem obviare nobis quae quaestum magnum praestabat dominis suis divinando
ACTS|16|17|haec subsecuta Paulum et nos clamabat dicens isti homines servi Dei excelsi sunt qui adnuntiant vobis viam salutis
ACTS|16|18|hoc autem faciebat multis diebus dolens autem Paulus et conversus spiritui dixit praecipio tibi in nomine Iesu Christi exire ab ea et exiit eadem hora
ACTS|16|19|videntes autem domini eius quia exivit spes quaestus eorum adprehendentes Paulum et Silam perduxerunt in forum ad principes
ACTS|16|20|et offerentes eos magistratibus dixerunt hii homines conturbant civitatem nostram cum sint Iudaei
ACTS|16|21|et adnuntiant morem quem non licet nobis suscipere neque facere cum simus Romani
ACTS|16|22|et concurrit plebs adversus eos et magistratus scissis tunicis eorum iusserunt virgis caedi
ACTS|16|23|et cum multas plagas eis inposuissent miserunt eos in carcerem praecipientes custodi ut diligenter custodiret eos
ACTS|16|24|qui cum tale praeceptum accepisset misit eos in interiorem carcerem et pedes eorum strinxit in ligno
ACTS|16|25|media autem nocte Paulus et Silas adorantes laudabant Deum et audiebant eos qui in custodia erant
ACTS|16|26|subito vero terraemotus factus est magnus ita ut moverentur fundamenta carceris et aperta sunt statim ostia omnia et universorum vincula soluta sunt
ACTS|16|27|expergefactus autem custos carceris et videns apertas ianuas carceris evaginato gladio volebat se interficere aestimans fugisse vinctos
ACTS|16|28|clamavit autem Paulus magna voce dicens nihil feceris tibi mali universi enim hic sumus
ACTS|16|29|petitoque lumine introgressus est et tremefactus procidit Paulo et Silae
ACTS|16|30|et producens eos foras ait domini quid me oportet facere ut salvus fiam
ACTS|16|31|at illi dixerunt crede in Domino Iesu et salvus eris tu et domus tua
ACTS|16|32|et locuti sunt ei verbum Domini cum omnibus qui erant in domo eius
ACTS|16|33|et tollens eos in illa hora noctis lavit plagas eorum et baptizatus est ipse et omnes eius continuo
ACTS|16|34|cumque perduxisset eos in domum suam adposuit eis mensam et laetatus est cum omni domo sua credens Deo
ACTS|16|35|et cum dies factus esset miserunt magistratus lictores dicentes dimitte homines illos
ACTS|16|36|nuntiavit autem custos carceris verba haec Paulo quia miserunt magistratus ut dimittamini nunc igitur exeuntes ite in pace
ACTS|16|37|Paulus autem dixit eis caesos nos publice indemnatos homines romanos miserunt in carcerem et nunc occulte nos eiciunt non ita sed veniant
ACTS|16|38|et ipsi nos eiciant nuntiaverunt autem magistratibus lictores verba haec timueruntque audito quod Romani essent
ACTS|16|39|et venientes deprecati sunt eos et educentes rogabant ut egrederentur urbem
ACTS|16|40|exeuntes autem de carcere introierunt ad Lydiam et visis fratribus consolati sunt eos et profecti sunt
ACTS|17|1|cum autem perambulassent Amphipolim et Apolloniam venerunt Thessalonicam ubi erat synagoga Iudaeorum
ACTS|17|2|secundum consuetudinem autem Paulus introivit ad eos et per sabbata tria disserebat eis de scripturis
ACTS|17|3|adaperiens et insinuans quia Christum oportuit pati et resurgere a mortuis et quia hic est Christus Iesus quem ego adnuntio vobis
ACTS|17|4|et quidam ex eis crediderunt et adiuncti sunt Paulo et Silae et de colentibus gentilibusque multitudo magna et mulieres nobiles non paucae
ACTS|17|5|zelantes autem Iudaei adsumentesque de vulgo viros quosdam malos et turba facta concitaverunt civitatem et adsistentes domui Iasonis quaerebant eos producere in populum
ACTS|17|6|et cum non invenissent eos trahebant Iasonem et quosdam fratres ad principes civitatis clamantes quoniam hii qui orbem concitant et huc venerunt
ACTS|17|7|quos suscepit Iason et hii omnes contra decreta Caesaris faciunt regem alium dicentes esse Iesum
ACTS|17|8|concitaverunt autem plebem et principes civitatis audientes haec
ACTS|17|9|et accepto satis ab Iasone et a ceteris dimiserunt eos
ACTS|17|10|fratres vero confestim per noctem dimiserunt Paulum et Silam in Beroeam qui cum advenissent in synagogam Iudaeorum introierunt
ACTS|17|11|hii autem erant nobiliores eorum qui sunt Thessalonicae qui susceperunt verbum cum omni aviditate cotidie scrutantes scripturas si haec ita se haberent
ACTS|17|12|et multi quidem crediderunt ex eis et gentilium mulierum honestarum et viri non pauci
ACTS|17|13|cum autem cognovissent in Thessalonica Iudaei quia et Beroeae praedicatum est a Paulo verbum Dei venerunt et illuc commoventes et turbantes multitudinem
ACTS|17|14|statimque tunc Paulum dimiserunt fratres ut iret usque ad mare Silas autem et Timotheus remanserunt ibi
ACTS|17|15|qui autem deducebant Paulum perduxerunt usque Athenas et accepto mandato ab eo ad Silam et Timotheum ut quam celeriter venirent ad illum profecti sunt
ACTS|17|16|Paulus autem cum Athenis eos expectaret incitabatur spiritus eius in ipso videns idolatriae deditam civitatem
ACTS|17|17|disputabat igitur in synagoga cum Iudaeis et colentibus et in foro per omnes dies ad eos qui aderant
ACTS|17|18|quidam autem epicurei et stoici philosophi disserebant cum eo et quidam dicebant quid vult seminiverbius hic dicere alii vero novorum daemoniorum videtur adnuntiator esse quia Iesum et resurrectionem adnuntiabat eis
ACTS|17|19|et adprehensum eum ad Ariopagum duxerunt dicentes possumus scire quae est haec nova quae a te dicitur doctrina
ACTS|17|20|nova enim quaedam infers auribus nostris volumus ergo scire quidnam velint haec esse
ACTS|17|21|Athenienses autem omnes et advenae hospites ad nihil aliud vacabant nisi aut dicere aut audire aliquid novi
ACTS|17|22|stans autem Paulus in medio Ariopagi ait viri athenienses per omnia quasi superstitiosiores vos video
ACTS|17|23|praeteriens enim et videns simulacra vestra inveni et aram in qua scriptum erat ignoto deo quod ergo ignorantes colitis hoc ego adnuntio vobis
ACTS|17|24|Deus qui fecit mundum et omnia quae in eo sunt hic caeli et terrae cum sit Dominus non in manufactis templis inhabitat
ACTS|17|25|nec manibus humanis colitur indigens aliquo cum ipse det omnibus vitam et inspirationem et omnia
ACTS|17|26|fecitque ex uno omne genus hominum inhabitare super universam faciem terrae definiens statuta tempora et terminos habitationis eorum
ACTS|17|27|quaerere Deum si forte adtractent eum aut inveniant quamvis non longe sit ab unoquoque nostrum
ACTS|17|28|in ipso enim vivimus et movemur et sumus sicut et quidam vestrum poetarum dixerunt ipsius enim et genus sumus
ACTS|17|29|genus ergo cum simus Dei non debemus aestimare auro aut argento aut lapidi sculpturae artis et cogitationis hominis divinum esse simile
ACTS|17|30|et tempora quidem huius ignorantiae despiciens Deus nunc adnuntiat hominibus ut omnes ubique paenitentiam agant
ACTS|17|31|eo quod statuit diem in qua iudicaturus est orbem in aequitate in viro in quo statuit fidem praebens omnibus suscitans eum a mortuis
ACTS|17|32|cum audissent autem resurrectionem mortuorum quidam quidem inridebant quidam vero dixerunt audiemus te de hoc iterum
ACTS|17|33|sic Paulus exivit de medio eorum
ACTS|17|34|quidam vero viri adherentes ei crediderunt in quibus et Dionisius Ariopagita et mulier nomine Damaris et alii cum eis
ACTS|18|1|post haec egressus ab Athenis venit Corinthum
ACTS|18|2|et inveniens quendam Iudaeum nomine Aquilam Ponticum genere qui nuper venerat ab Italia et Priscillam uxorem eius eo quod praecepisset Claudius discedere omnes Iudaeos a Roma accessit ad eos
ACTS|18|3|et quia eiusdem erat artis manebat apud eos et operabatur erat autem scenofactoriae artis
ACTS|18|4|
ACTS|18|5|cum venissent autem de Macedonia Silas et Timotheus instabat verbo Paulus testificans Iudaeis esse Christum Iesum
ACTS|18|6|contradicentibus autem eis et blasphemantibus excutiens vestimenta dixit ad eos sanguis vester super caput vestrum mundus ego ex hoc ad gentes vadam
ACTS|18|7|et migrans inde intravit in domum cuiusdam nomine Titi Iusti colentis Deum cuius domus erat coniuncta synagogae
ACTS|18|8|Crispus autem archisynagogus credidit Domino cum omni domo sua et multi Corinthiorum audientes credebant et baptizabantur
ACTS|18|9|dixit autem Dominus nocte per visionem Paulo noli timere sed loquere et ne taceas
ACTS|18|10|propter quod ego sum tecum et nemo adponetur tibi ut noceat te quoniam populus est mihi multus in hac civitate
ACTS|18|11|sedit autem annum et sex menses docens apud eos verbum Dei
ACTS|18|12|Gallione autem proconsule Achaiae insurrexerunt uno animo Iudaei in Paulum et adduxerunt eum ad tribunal
ACTS|18|13|dicentes quia contra legem hic persuadet hominibus colere Deum
ACTS|18|14|incipiente autem Paulo aperire os dixit Gallio ad Iudaeos si quidem esset iniquum aliquid aut facinus pessimum o viri iudaei recte vos sustinerem
ACTS|18|15|si vero quaestiones sunt de verbo et nominibus et legis vestrae vos ipsi videritis iudex ego horum nolo esse
ACTS|18|16|et minavit eos a tribunali
ACTS|18|17|adprehendentes autem omnes Sosthenen principem synagogae percutiebant ante tribunal et nihil eorum Gallioni curae erat
ACTS|18|18|Paulus vero cum adhuc sustinuisset dies multos fratribus valefaciens navigavit Syriam et cum eo Priscilla et Aquila qui sibi totonderat in Cencris caput habebat enim votum
ACTS|18|19|devenitque Ephesum et illos ibi reliquit ipse vero ingressus synagogam disputavit cum Iudaeis
ACTS|18|20|rogantibus autem eis ut ampliori tempore maneret non consensit
ACTS|18|21|sed valefaciens et dicens iterum revertar ad vos Deo volente profectus est ab Epheso
ACTS|18|22|et descendens Caesaream ascendit et salutavit ecclesiam et descendit Antiochiam
ACTS|18|23|et facto ibi aliquanto tempore profectus est perambulans ex ordine galaticam regionem et Frygiam confirmans omnes discipulos
ACTS|18|24|Iudaeus autem quidam Apollo nomine Alexandrinus natione vir eloquens devenit Ephesum potens in scripturis
ACTS|18|25|hic erat edoctus viam Domini et fervens spiritu loquebatur et docebat diligenter ea quae sunt Iesu sciens tantum baptisma Iohannis
ACTS|18|26|hic ergo coepit fiducialiter agere in synagoga quem cum audissent Priscilla et Aquila adsumpserunt eum et diligentius exposuerunt ei viam Dei
ACTS|18|27|cum autem vellet ire Achaiam exhortati fratres scripserunt discipulis ut susciperent eum qui cum venisset contulit multum his qui crediderant
ACTS|18|28|vehementer enim Iudaeos revincebat publice ostendens per scripturas esse Christum Iesum
ACTS|19|1|factum est autem cum Apollo esset Corinthi ut Paulus peragratis superioribus partibus veniret Ephesum et inveniret quosdam discipulos
ACTS|19|2|dixitque ad eos si Spiritum Sanctum accepistis credentes at illi ad eum sed neque si Spiritus Sanctus est audivimus
ACTS|19|3|ille vero ait in quo ergo baptizati estis qui dixerunt in Iohannis baptismate
ACTS|19|4|dixit autem Paulus Iohannes baptizavit baptisma paenitentiae populum dicens in eum qui venturus esset post ipsum ut crederent hoc est in Iesum
ACTS|19|5|his auditis baptizati sunt in nomine Domini Iesu
ACTS|19|6|et cum inposuisset illis manum Paulus venit Spiritus Sanctus super eos et loquebantur linguis et prophetabant
ACTS|19|7|erant autem omnes viri fere duodecim
ACTS|19|8|introgressus autem synagogam cum fiducia loquebatur per tres menses disputans et suadens de regno Dei
ACTS|19|9|cum autem quidam indurarentur et non crederent maledicentes viam coram multitudine discedens ab eis segregavit discipulos cotidie disputans in scola Tyranni
ACTS|19|10|hoc autem factum est per biennium ita ut omnes qui habitabant in Asia audirent verbum Domini Iudaei atque gentiles
ACTS|19|11|virtutesque non quaslibet Deus faciebat per manus Pauli
ACTS|19|12|ita ut etiam super languidos deferrentur a corpore eius sudaria vel semicintia et recedebant ab eis languores et spiritus nequam egrediebantur
ACTS|19|13|temptaverunt autem quidam et de circumeuntibus iudaeis exorcistis invocare super eos qui habebant spiritus malos nomen Domini Iesu dicentes adiuro vos per Iesum quem Paulus praedicat
ACTS|19|14|erant autem quidam Scevae Iudaei principis sacerdotum septem filii qui hoc faciebant
ACTS|19|15|respondens autem spiritus nequam dixit eis Iesum novi et Paulum scio vos autem qui estis
ACTS|19|16|et insiliens homo in eos in quo erat daemonium pessimum et dominatus amborum invaluit contra eos ita ut nudi et vulnerati effugerent de domo illa
ACTS|19|17|hoc autem notum factum est omnibus Iudaeis atque gentilibus qui habitabant Ephesi et cecidit timor super omnes illos et magnificabatur nomen Domini Iesu
ACTS|19|18|multique credentium veniebant confitentes et adnuntiantes actus suos
ACTS|19|19|multi autem ex his qui fuerant curiosa sectati contulerunt libros et conbuserunt coram omnibus et conputatis pretiis illorum invenerunt pecuniam denariorum quinquaginta milium
ACTS|19|20|ita fortiter verbum Dei crescebat et confirmabatur
ACTS|19|21|his autem expletis posuit Paulus in Spiritu transita Macedonia et Achaia ire Hierosolymam dicens quoniam postquam fuero ibi oportet me et Romam videre
ACTS|19|22|mittens autem in Macedoniam duos ex ministrantibus sibi Timotheum et Erastum ipse remansit ad tempus in Asia
ACTS|19|23|facta est autem in illo tempore turbatio non minima de via
ACTS|19|24|Demetrius enim quidam nomine argentarius faciens aedes argenteas Dianae praestabat artificibus non modicum quaestum
ACTS|19|25|quos convocans et eos qui eiusmodi erant opifices dixit viri scitis quia de hoc artificio adquisitio est nobis
ACTS|19|26|et videtis et auditis quia non solum Ephesi sed paene totius Asiae Paulus hic suadens avertit multam turbam dicens quoniam non sunt dii qui manibus fiunt
ACTS|19|27|non solum autem haec periclitabitur nobis pars in redargutionem venire sed et magnae deae Dianae templum in nihilum reputabitur sed et destrui incipiet maiestas eius quam tota Asia et orbis colit
ACTS|19|28|his auditis repleti sunt ira et exclamaverunt dicentes magna Diana Ephesiorum
ACTS|19|29|et impleta est civitas confusione et impetum fecerunt uno animo in theatrum rapto Gaio et Aristarcho Macedonibus comitibus Pauli
ACTS|19|30|Paulo autem volente intrare in populum non permiserunt discipuli
ACTS|19|31|quidam autem et de Asiae principibus qui erant amici eius miserunt ad eum rogantes ne se daret in theatrum
ACTS|19|32|alii autem aliud clamabant erat enim ecclesia confusa et plures nesciebant qua ex causa convenissent
ACTS|19|33|de turba autem detraxerunt Alexandrum propellentibus eum Iudaeis Alexander ergo manu silentio postulato volebat rationem reddere populo
ACTS|19|34|quem ut cognoverunt Iudaeum esse vox facta est una omnium quasi per horas duas clamantium magna Diana Ephesiorum
ACTS|19|35|et cum sedasset scriba turbas dixit viri ephesii quis enim est hominum qui nesciat Ephesiorum civitatem cultricem esse magnae Dianae Iovisque prolis
ACTS|19|36|cum ergo his contradici non possit oportet vos sedatos esse et nihil temere agere
ACTS|19|37|adduxistis enim homines istos neque sacrilegos neque blasphemantes deam vestram
ACTS|19|38|quod si Demetrius et qui cum eo sunt artifices habent adversus aliquem causam conventus forenses aguntur et pro consulibus sunt accusent invicem
ACTS|19|39|si quid autem alterius rei quaeritis in legitima ecclesia poterit absolvi
ACTS|19|40|nam et periclitamur argui seditionis hodiernae cum nullus obnoxius sit de quo non possimus reddere rationem concursus istius et cum haec dixisset dimisit ecclesiam
ACTS|20|1|postquam autem cessavit tumultus vocatis Paulus discipulis et exhortatus eos valedixit et profectus est ut iret in Macedoniam
ACTS|20|2|cum autem perambulasset partes illas et exhortatus eos fuisset multo sermone venit ad Graeciam
ACTS|20|3|ubi cum fecisset menses tres factae sunt illi insidiae a Iudaeis navigaturo in Syriam habuitque consilium ut reverteretur per Macedoniam
ACTS|20|4|comitatus est autem eum Sopater Pyrri Beroensis Thessalonicensium vero Aristarchus et Secundus et Gaius Derbeus et Timotheus Asiani vero Tychicus et Trophimus
ACTS|20|5|hii cum praecessissent sustinebant nos Troade
ACTS|20|6|nos vero navigavimus post dies azymorum a Philippis et venimus ad eos Troadem in diebus quinque ubi demorati sumus diebus septem
ACTS|20|7|in una autem sabbati cum convenissemus ad frangendum panem Paulus disputabat eis profecturus in crastinum protraxitque sermonem usque in mediam noctem
ACTS|20|8|erant autem lampades copiosae in cenaculo ubi eramus congregati
ACTS|20|9|sedens autem quidam adulescens nomine Eutychus super fenestram cum mergeretur somno gravi disputante diu Paulo eductus somno cecidit de tertio cenaculo deorsum et sublatus est mortuus
ACTS|20|10|ad quem cum descendisset Paulus incubuit super eum et conplexus dixit nolite turbari anima enim ipsius in eo est
ACTS|20|11|ascendens autem frangensque panem et gustans satisque adlocutus usque in lucem sic profectus est
ACTS|20|12|adduxerunt autem puerum viventem et consolati sunt non minime
ACTS|20|13|nos autem ascendentes navem enavigavimus in Asson inde suscepturi Paulum sic enim disposuerat ipse per terram iter facturus
ACTS|20|14|cum autem convenisset nos in Asson adsumpto eo venimus Mytilenen
ACTS|20|15|et inde navigantes sequenti die venimus contra Chium et alia adplicuimus Samum et sequenti venimus Miletum
ACTS|20|16|proposuerat enim Paulus transnavigare Ephesum ne qua mora illi fieret in Asia festinabat enim si possibile sibi esset ut diem pentecosten faceret Hierosolymis
ACTS|20|17|a Mileto autem mittens Ephesum vocavit maiores natu ecclesiae
ACTS|20|18|qui cum venissent ad eum et simul essent dixit eis vos scitis a prima die qua ingressus sum in Asiam qualiter vobiscum per omne tempus fuerim
ACTS|20|19|serviens Domino cum omni humilitate et lacrimis et temptationibus quae mihi acciderunt ex insidiis Iudaeorum
ACTS|20|20|quomodo nihil subtraxerim utilium quo minus adnuntiarem vobis et docerem vos publice et per domos
ACTS|20|21|testificans Iudaeis atque gentilibus in Deum paenitentiam et fidem in Dominum nostrum Iesum Christum
ACTS|20|22|et nunc ecce alligatus ego Spiritu vado in Hierusalem quae in ea eventura sint mihi ignorans
ACTS|20|23|nisi quod Spiritus Sanctus per omnes civitates protestatur mihi dicens quoniam vincula et tribulationes me manent
ACTS|20|24|sed nihil horum vereor nec facio animam pretiosiorem quam me dummodo consummem cursum meum et ministerium quod accepi a Domino Iesu testificari evangelium gratiae Dei
ACTS|20|25|et nunc ecce ego scio quia amplius non videbitis faciem meam vos omnes per quos transivi praedicans regnum Dei
ACTS|20|26|quapropter contestor vos hodierna die quia mundus sum a sanguine omnium
ACTS|20|27|non enim subterfugi quo minus adnuntiarem omne consilium Dei vobis
ACTS|20|28|adtendite vobis et universo gregi in quo vos Spiritus Sanctus posuit episcopos regere ecclesiam Dei quam adquisivit sanguine suo
ACTS|20|29|ego scio quoniam intrabunt post discessionem meam lupi graves in vos non parcentes gregi
ACTS|20|30|et ex vobis ipsis exsurgent viri loquentes perversa ut abducant discipulos post se
ACTS|20|31|propter quod vigilate memoria retinentes quoniam per triennium nocte et die non cessavi cum lacrimis monens unumquemque vestrum
ACTS|20|32|et nunc commendo vos Deo et verbo gratiae ipsius qui potens est aedificare et dare hereditatem in sanctificatis omnibus
ACTS|20|33|argentum aut aurum aut vestem nullius concupivi
ACTS|20|34|ipsi scitis quoniam ad ea quae mihi opus erant et his qui mecum sunt ministraverunt manus istae
ACTS|20|35|omnia ostendi vobis quoniam sic laborantes oportet suscipere infirmos ac meminisse verbi Domini Iesu quoniam ipse dixit beatius est magis dare quam accipere
ACTS|20|36|et cum haec dixisset positis genibus suis cum omnibus illis oravit
ACTS|20|37|magnus autem fletus factus est omnium et procumbentes super collum Pauli osculabantur eum
ACTS|20|38|dolentes maxime in verbo quo dixerat quoniam amplius faciem eius non essent visuri et deducebant eum ad navem
ACTS|21|1|cum autem factum esset ut navigaremus abstracti ab eis recto cursu venimus Cho et sequenti die Rhodum et inde Patara
ACTS|21|2|et cum invenissemus navem transfretantem in Foenicen ascendentes navigavimus
ACTS|21|3|cum paruissemus autem Cypro et relinquentes eam ad sinistram navigabamus in Syriam et venimus Tyrum ibi enim navis erat expositura onus
ACTS|21|4|inventis autem discipulis mansimus ibi diebus septem qui Paulo dicebant per Spiritum ne ascenderet Hierosolymam
ACTS|21|5|et explicitis diebus profecti ibamus deducentibus nos omnibus cum uxoribus et filiis usque foras civitatem et positis genibus in litore oravimus
ACTS|21|6|et cum valefecissemus invicem ascendimus in navem illi autem redierunt in sua
ACTS|21|7|nos vero navigatione explicita a Tyro descendimus Ptolomaida et salutatis fratribus mansimus die una apud illos
ACTS|21|8|alia autem die profecti venimus Caesaream et intrantes in domum Philippi evangelistae qui erat de septem mansimus apud eum
ACTS|21|9|huic autem erant filiae quattuor virgines prophetantes
ACTS|21|10|et cum moraremur per dies aliquot supervenit quidam a Iudaea propheta nomine Agabus
ACTS|21|11|is cum venisset ad nos tulit zonam Pauli et alligans sibi pedes et manus dixit haec dicit Spiritus Sanctus virum cuius est zona haec sic alligabunt in Hierusalem Iudaei et tradent in manus gentium
ACTS|21|12|quod cum audissemus rogabamus nos et qui loci illius erant ne ascenderet Hierosolymam
ACTS|21|13|tunc respondit Paulus et dixit quid facitis flentes et adfligentes cor meum ego enim non solum alligari sed et mori in Hierusalem paratus sum propter nomen Domini Iesu
ACTS|21|14|et cum ei suadere non possemus quievimus dicentes Domini voluntas fiat
ACTS|21|15|post dies autem istos praeparati ascendebamus Hierusalem
ACTS|21|16|venerunt autem et ex discipulis a Caesarea nobiscum adducentes apud quem hospitaremur Mnasonem quendam Cyprium antiquum discipulum
ACTS|21|17|et cum venissemus Hierosolymam libenter exceperunt nos fratres
ACTS|21|18|sequenti autem die introibat Paulus nobiscum ad Iacobum omnesque collecti sunt seniores
ACTS|21|19|quos cum salutasset narrabat per singula quae fecisset Deus in gentibus per ministerium ipsius
ACTS|21|20|at illi cum audissent magnificabant Deum dixeruntque ei vides frater quot milia sint in Iudaeis qui crediderunt et omnes aemulatores sunt legis
ACTS|21|21|audierunt autem de te quia discessionem doceas a Mose eorum qui per gentes sunt Iudaeorum dicens non debere circumcidere eos filios suos neque secundum consuetudinem ingredi
ACTS|21|22|quid ergo est utique oportet convenire multitudinem audient enim te supervenisse
ACTS|21|23|hoc ergo fac quod tibi dicimus sunt nobis viri quattuor votum habentes super se
ACTS|21|24|his adsumptis sanctifica te cum illis et inpende in illis ut radant capita et scient omnes quia quae de te audierunt falsa sunt sed ambulas et ipse custodiens legem
ACTS|21|25|de his autem qui crediderunt ex gentibus nos scripsimus iudicantes ut abstineant se ab idolis immolato et sanguine et suffocato et fornicatione
ACTS|21|26|tunc Paulus adsumptis viris postera die purificatus cum illis intravit in templum adnuntians expletionem dierum purificationis donec offerretur pro unoquoque eorum oblatio
ACTS|21|27|dum autem septem dies consummarentur hii qui de Asia erant Iudaei cum vidissent eum in templo concitaverunt omnem populum et iniecerunt ei manus clamantes
ACTS|21|28|viri israhelitae adiuvate hic est homo qui adversus populum et legem et locum hunc omnes ubique docens insuper et gentiles induxit in templum et violavit sanctum locum istum
ACTS|21|29|viderant enim Trophimum Ephesium in civitate cum ipso quem aestimaverunt quoniam in templum induxisset Paulus
ACTS|21|30|commotaque est civitas tota et facta est concursio populi et adprehendentes Paulum trahebant eum extra templum et statim clausae sunt ianuae
ACTS|21|31|quaerentibus autem eum occidere nuntiatum est tribuno cohortis quia tota confunditur Hierusalem
ACTS|21|32|qui statim adsumptis militibus et centurionibus decucurrit ad illos qui cum vidissent tribunum et milites cessaverunt percutere Paulum
ACTS|21|33|tunc accedens tribunus adprehendit eum et iussit alligari catenis duabus et interrogabat quis esset et quid fecisset
ACTS|21|34|alii autem aliud clamabant in turba et cum non posset certum cognoscere prae tumultu iussit duci eum in castra
ACTS|21|35|et cum venisset ad gradus contigit ut portaretur a militibus propter vim populi
ACTS|21|36|sequebatur enim multitudo populi clamans tolle eum
ACTS|21|37|et cum coepisset induci in castra Paulus dicit tribuno si licet mihi loqui aliquid ad te qui dixit graece nosti
ACTS|21|38|nonne tu es Aegyptius qui ante hos dies tumultum concitasti et eduxisti in desertum quattuor milia virorum sicariorum
ACTS|21|39|et dixit ad eum Paulus ego homo sum quidem iudaeus a Tarso Ciliciae non ignotae civitatis municeps rogo autem te permitte mihi loqui ad populum
ACTS|21|40|et cum ille permisisset Paulus stans in gradibus annuit manu ad plebem et magno silentio facto adlocutus est hebraea lingua dicens
ACTS|22|1|viri fratres et patres audite quam ad vos nunc reddo rationem
ACTS|22|2|cum audissent autem quia hebraea lingua loquitur ad illos magis praestiterunt silentium
ACTS|22|3|et dixit ego sum vir iudaeus natus Tarso Ciliciae nutritus autem in ista civitate secus pedes Gamalihel eruditus iuxta veritatem paternae legis aemulator legis sicut et vos omnes estis hodie
ACTS|22|4|qui hanc viam persecutus sum usque ad mortem alligans et tradens in custodias viros ac mulieres
ACTS|22|5|sicut princeps sacerdotum testimonium mihi reddit et omnes maiores natu a quibus et epistulas accipiens ad fratres Damascum pergebam ut adducerem inde vinctos in Hierusalem uti punirentur
ACTS|22|6|factum est autem eunte me et adpropinquante Damasco media die subito de caelo circumfulsit me lux copiosa
ACTS|22|7|et decidens in terram audivi vocem dicentem mihi Saule Saule quid me persequeris
ACTS|22|8|ego autem respondi quis es Domine dixitque ad me ego sum Iesus Nazarenus quem tu persequeris
ACTS|22|9|et qui mecum erant lumen quidem viderunt vocem autem non audierunt eius qui loquebatur mecum
ACTS|22|10|et dixi quid faciam Domine Dominus autem dixit ad me surgens vade Damascum et ibi tibi dicetur de omnibus quae te oporteat facere
ACTS|22|11|et cum non viderem prae claritate luminis illius ad manum deductus a comitibus veni Damascum
ACTS|22|12|Ananias autem quidam vir secundum legem testimonium habens ab omnibus habitantibus Iudaeis
ACTS|22|13|veniens ad me et adstans dixit mihi Saule frater respice et ego eadem hora respexi in eum
ACTS|22|14|at ille dixit Deus patrum nostrorum praeordinavit te ut cognosceres voluntatem eius et videres Iustum et audires vocem ex ore eius
ACTS|22|15|quia eris testis illius ad omnes homines eorum quae vidisti et audisti
ACTS|22|16|et nunc quid moraris exsurge baptizare et ablue peccata tua invocato nomine ipsius
ACTS|22|17|factum est autem revertenti mihi in Hierusalem et oranti in templo fieri me in stupore mentis
ACTS|22|18|et videre illum dicentem mihi festina et exi velociter ex Hierusalem quoniam non recipient testimonium tuum de me
ACTS|22|19|et ego dixi Domine ipsi sciunt quia ego eram concludens in carcerem et caedens per synagogas eos qui credebant in te
ACTS|22|20|et cum funderetur sanguis Stephani testis tui ego adstabam et consentiebam et custodiebam vestimenta interficientium illum
ACTS|22|21|et dixit ad me vade quoniam ego in nationes longe mittam te
ACTS|22|22|audiebant autem eum usque ad hoc verbum et levaverunt vocem suam dicentes tolle de terra eiusmodi non enim fas est eum vivere
ACTS|22|23|vociferantibus autem eis et proicientibus vestimenta sua et pulverem iactantibus in aerem
ACTS|22|24|iussit tribunus induci eum in castra et flagellis caedi et torqueri eum ut sciret propter quam causam sic adclamarent ei
ACTS|22|25|et cum adstrinxissent eum loris dixit adstanti sibi centurioni Paulus si hominem romanum et indemnatum licet vobis flagellare
ACTS|22|26|quo audito centurio accessit ad tribunum et nuntiavit dicens quid acturus es hic enim homo civis romanus est
ACTS|22|27|accedens autem tribunus dixit illi dic mihi tu Romanus es at ille dixit etiam
ACTS|22|28|et respondit tribunus ego multa summa civitatem hanc consecutus sum et Paulus ait ego autem et natus sum
ACTS|22|29|protinus ergo discesserunt ab illo qui eum torturi erant tribunus quoque timuit postquam rescivit quia civis romanus esset et quia alligasset eum
ACTS|22|30|postera autem die volens scire diligentius qua ex causa accusaretur a Iudaeis solvit eum et iussit sacerdotes convenire et omne concilium et producens Paulum statuit inter illos
ACTS|23|1|intendens autem concilium Paulus ait viri fratres ego omni conscientia bona conversatus sum ante Deum usque in hodiernum diem
ACTS|23|2|princeps autem sacerdotum Ananias praecepit adstantibus sibi percutere os eius
ACTS|23|3|tunc Paulus ad eum dixit percutiet te Deus paries dealbate et tu sedens iudicas me secundum legem et contra legem iubes me percuti
ACTS|23|4|et qui adstabant dixerunt summum sacerdotem Dei maledicis
ACTS|23|5|dixit autem Paulus nesciebam fratres quia princeps est sacerdotum scriptum est enim principem populi tui non maledices
ACTS|23|6|sciens autem Paulus quia una pars esset Sadducaeorum et altera Pharisaeorum exclamavit in concilio viri fratres ego Pharisaeus sum filius Pharisaeorum de spe et resurrectione mortuorum ego iudicor
ACTS|23|7|et cum haec dixisset facta est dissensio inter Pharisaeos et Sadducaeos et soluta est multitudo
ACTS|23|8|Sadducaei enim dicunt non esse resurrectionem neque angelum neque spiritum Pharisaei autem utrumque confitentur
ACTS|23|9|factus est autem clamor magnus et surgentes quidam Pharisaeorum pugnabant dicentes nihil mali invenimus in homine isto quod si spiritus locutus est ei aut angelus
ACTS|23|10|et cum magna dissensio facta esset timens tribunus ne discerperetur Paulus ab ipsis iussit milites descendere et rapere eum de medio eorum ac deducere eum in castra
ACTS|23|11|sequenti autem nocte adsistens ei Dominus ait constans esto sicut enim testificatus es de me Hierusalem sic te oportet et Romae testificari
ACTS|23|12|facta autem die collegerunt se quidam ex Iudaeis et devoverunt se dicentes neque manducaturos neque bibituros donec occiderent Paulum
ACTS|23|13|erant autem plus quam quadraginta qui hanc coniurationem fecerant
ACTS|23|14|qui accesserunt ad principes sacerdotum et seniores et dixerunt devotione devovimus nos nihil gustaturos donec occidamus Paulum
ACTS|23|15|nunc ergo vos notum facite tribuno cum concilio ut producat illum ad vos tamquam aliquid certius cognituri de eo nos vero priusquam adpropiet parati sumus interficere illum
ACTS|23|16|quod cum audisset filius sororis Pauli insidias venit et intravit in castra nuntiavitque Paulo
ACTS|23|17|vocans autem Paulus ad se unum ex centurionibus ait adulescentem hunc perduc ad tribunum habet enim aliquid indicare illi
ACTS|23|18|et ille quidem adsumens eum duxit ad tribunum et ait vinctus Paulus vocans rogavit me hunc adulescentem perducere ad te habentem aliquid loqui tibi
ACTS|23|19|adprehendens autem tribunus manum illius secessit cum eo seorsum et interrogavit illum quid est quod habes indicare mihi
ACTS|23|20|ille autem dixit Iudaeis convenit rogare te ut crastina die Paulum producas in concilium quasi aliquid certius inquisituri sint de illo
ACTS|23|21|tu vero ne credideris illis insidiantur enim ei ex eis viri amplius quadraginta qui se devoverunt non manducare neque bibere donec interficiant eum et nunc parati sunt expectantes promissum tuum
ACTS|23|22|tribunus igitur dimisit adulescentem praecipiens ne cui loqueretur quoniam haec nota sibi fecisset
ACTS|23|23|et vocatis duobus centurionibus dixit illis parate milites ducentos ut eant usque Caesaream et equites septuaginta et lancearios ducentos a tertia hora noctis
ACTS|23|24|et iumenta praeparate ut inponentes Paulum salvum perducerent ad Felicem praesidem
ACTS|23|25|
ACTS|23|26|scribens epistulam continentem haec Claudius Lysias optimo praesidi Felici salutem
ACTS|23|27|virum hunc conprehensum a Iudaeis et incipientem interfici ab eis superveniens cum exercitu eripui cognito quia Romanus est
ACTS|23|28|volensque scire causam quam obiciebant illi deduxi eum in concilium eorum
ACTS|23|29|quem inveni accusari de quaestionibus legis ipsorum nihil vero dignum morte aut vinculis habentem crimen
ACTS|23|30|et cum mihi perlatum esset de insidiis quas paraverunt ei misi ad te denuntians et accusatoribus ut dicant apud te
ACTS|23|31|milites ergo secundum praeceptum sibi adsumentes Paulum duxerunt per noctem in Antipatridem
ACTS|23|32|et postera die dimissis equitibus ut irent cum eo reversi sunt ad castra
ACTS|23|33|qui cum venissent Caesaream et tradidissent epistulam praesidi statuerunt ante illum et Paulum
ACTS|23|34|cum legisset autem et interrogasset de qua provincia esset et cognoscens quia de Cilicia
ACTS|23|35|audiam te inquit cum et accusatores tui venerint iussitque in praetorio Herodis custodiri eum
ACTS|24|1|post quinque autem dies descendit princeps sacerdotum Ananias cum senioribus quibusdam et Tertullo quodam oratore qui adierunt praesidem adversus Paulum
ACTS|24|2|et citato Paulo coepit accusare Tertullus dicens cum in multa pace agamus per te et multa corrigantur per tuam providentiam
ACTS|24|3|semper et ubique suscipimus optime Felix cum omni gratiarum actione
ACTS|24|4|ne diutius autem te protraham oro breviter audias nos pro tua clementia
ACTS|24|5|invenimus hunc hominem pestiferum et concitantem seditiones omnibus Iudaeis in universo orbe et auctorem seditionis sectae Nazarenorum
ACTS|24|6|qui etiam templum violare conatus est quem et adprehendimus
ACTS|24|7|
ACTS|24|8|a quo poteris ipse iudicans de omnibus istis cognoscere de quibus nos accusamus eum
ACTS|24|9|adiecerunt autem et Iudaei dicentes haec ita se habere
ACTS|24|10|respondit autem Paulus annuente sibi praeside dicere ex multis annis esse te iudicem genti huic sciens bono animo pro me satisfaciam
ACTS|24|11|potes enim cognoscere quia non plus sunt dies mihi quam duodecim ex quo ascendi adorare in Hierusalem
ACTS|24|12|et neque in templo invenerunt me cum aliquo disputantem aut concursum facientem turbae neque in synagogis neque in civitate
ACTS|24|13|neque probare possunt tibi de quibus nunc accusant me
ACTS|24|14|confiteor autem hoc tibi quod secundum sectam quam dicunt heresim sic deservio patrio Deo meo credens omnibus quae in lege et prophetis scripta sunt
ACTS|24|15|spem habens in Deum quam et hii ipsi expectant resurrectionem futuram iustorum et iniquorum
ACTS|24|16|in hoc et ipse studeo sine offendiculo conscientiam habere ad Deum et ad homines semper
ACTS|24|17|post annos autem plures elemosynas facturus in gentem meam veni et oblationes et vota
ACTS|24|18|in quibus invenerunt me purificatum in templo non cum turba neque cum tumultu
ACTS|24|19|quidam autem ex Asia Iudaei quos oportebat apud te praesto esse et accusare si quid haberent adversum me
ACTS|24|20|aut hii ipsi dicant si quid invenerunt in me iniquitatis cum stem in concilio
ACTS|24|21|nisi de una hac solummodo voce qua clamavi inter eos stans quoniam de resurrectione mortuorum ego iudicor hodie a vobis
ACTS|24|22|distulit autem illos Felix certissime sciens de via dicens cum tribunus Lysias descenderit audiam vos
ACTS|24|23|iussitque centurioni custodiri eum et habere requiem nec quemquam prohibere de suis ministrare ei
ACTS|24|24|post aliquot autem dies veniens Felix cum Drusilla uxore sua quae erat Iudaea vocavit Paulum et audivit ab eo fidem quae est in Iesum Christum
ACTS|24|25|disputante autem illo de iustitia et castitate et de iudicio futuro timefactus Felix respondit quod nunc adtinet vade tempore autem oportuno accersiam te
ACTS|24|26|simul et sperans quia pecunia daretur a Paulo propter quod et frequenter accersiens eum loquebatur cum eo
ACTS|24|27|biennio autem expleto accepit successorem Felix Porcium Festum volens autem gratiam praestare Iudaeis Felix reliquit Paulum vinctum
ACTS|25|1|Festus ergo cum venisset in provinciam post triduum ascendit Hierosolymam a Caesarea
ACTS|25|2|adieruntque eum principes sacerdotum et primi Iudaeorum adversus Paulum et rogabant eum
ACTS|25|3|postulantes gratiam adversum eum ut iuberet perduci eum Hierusalem insidias tendentes ut eum interficerent in via
ACTS|25|4|Festus autem respondit servari Paulum in Caesarea se autem maturius profecturum
ACTS|25|5|qui ergo in vobis ait potentes sunt descendentes simul si quod est in viro crimen accusent eum
ACTS|25|6|demoratus autem inter eos dies non amplius quam octo aut decem descendit Caesaream et altera die sedit pro tribunali et iussit Paulum adduci
ACTS|25|7|qui cum perductus esset circumsteterunt eum qui ab Hierosolyma descenderant Iudaei multas et graves causas obicientes quas non poterant probare
ACTS|25|8|Paulo autem rationem reddente quoniam neque in legem Iudaeorum neque in templum neque in Caesarem quicquam peccavi
ACTS|25|9|Festus autem volens Iudaeis gratiam praestare respondens Paulo dixit vis Hierosolymam ascendere et ibi de his iudicari apud me
ACTS|25|10|dixit autem Paulus ad tribunal Caesaris sto ubi me oportet iudicari Iudaeis non nocui sicut tu melius nosti
ACTS|25|11|si enim nocui aut dignum morte aliquid feci non recuso mori si vero nihil est eorum quae hii accusant me nemo potest me illis donare Caesarem appello
ACTS|25|12|tunc Festus cum consilio locutus respondit Caesarem appellasti ad Caesarem ibis
ACTS|25|13|et cum dies aliquot transacti essent Agrippa rex et Bernice descenderunt Caesaream ad salutandum Festum
ACTS|25|14|et cum dies plures ibi demorarentur Festus regi indicavit de Paulo dicens vir quidam est derelictus a Felice vinctus
ACTS|25|15|de quo cum essem Hierosolymis adierunt me principes sacerdotum et seniores Iudaeorum postulantes adversus illum damnationem
ACTS|25|16|ad quos respondi quia non est consuetudo Romanis donare aliquem hominem priusquam is qui accusatur praesentes habeat accusatores locumque defendendi accipiat ad abluenda crimina
ACTS|25|17|cum ergo huc convenissent sine ulla dilatione sequenti die sedens pro tribunali iussi adduci virum
ACTS|25|18|de quo cum stetissent accusatores nullam causam deferebant de quibus ego suspicabar malum
ACTS|25|19|quaestiones vero quasdam de sua superstitione habebant adversus eum et de quodam Iesu defuncto quem adfirmabat Paulus vivere
ACTS|25|20|haesitans autem ego de huiusmodi quaestione dicebam si vellet ire Hierosolymam et ibi iudicari de istis
ACTS|25|21|Paulo autem appellante ut servaretur ad Augusti cognitionem iussi servari eum donec mittam eum ad Caesarem
ACTS|25|22|Agrippa autem ad Festum volebam et ipse hominem audire cras inquit audies eum
ACTS|25|23|altera autem die cum venisset Agrippa et Bernice cum multa ambitione et introissent in auditorium cum tribunis et viris principalibus civitatis et iubente Festo adductus est Paulus
ACTS|25|24|et dixit Festus Agrippa rex et omnes qui simul adestis nobiscum viri videtis hunc de quo omnis multitudo Iudaeorum interpellavit me Hierosolymis petens et hic clamantes non oportere eum vivere amplius
ACTS|25|25|ego vero conperi nihil dignum eum morte admisisse ipso autem hoc appellante Augustum iudicavi mittere
ACTS|25|26|de quo quid certum scribam domino non habeo propter quod produxi eum ad vos et maxime ad te rex Agrippa ut interrogatione facta habeam quid scribam
ACTS|25|27|sine ratione enim mihi videtur mittere vinctum et causas eius non significare
ACTS|26|1|Agrippa vero ad Paulum ait permittitur tibi loqui pro temet ipso tunc Paulus extenta manu coepit rationem reddere
ACTS|26|2|de omnibus quibus accusor a Iudaeis rex Agrippa aestimo me beatum apud te cum sim defensurus me hodie
ACTS|26|3|maxime te sciente omnia quae apud Iudaeos sunt consuetudines et quaestiones propter quod obsecro patienter me audias
ACTS|26|4|et quidem vitam meam a iuventute quae ab initio fuit in gente mea in Hierosolymis noverunt omnes Iudaei
ACTS|26|5|praescientes me ab initio si velint testimonium perhibere quoniam secundum certissimam sectam nostrae religionis vixi Pharisaeus
ACTS|26|6|et nunc in spe quae ad patres nostros repromissionis facta est a Deo sto iudicio subiectus
ACTS|26|7|in quam duodecim tribus nostrae nocte ac die deservientes sperant devenire de qua spe accusor a Iudaeis rex
ACTS|26|8|quid incredibile iudicatur apud vos si Deus mortuos suscitat
ACTS|26|9|et ego quidem existimaveram me adversus nomen Iesu Nazareni debere multa contraria agere
ACTS|26|10|quod et feci Hierosolymis et multos sanctorum ego in carceribus inclusi a principibus sacerdotum potestate accepta et cum occiderentur detuli sententiam
ACTS|26|11|et per omnes synagogas frequenter puniens eos conpellebam blasphemare et amplius insaniens in eos persequebar usque in exteras civitates
ACTS|26|12|in quibus dum irem Damascum cum potestate et permissu principum sacerdotum
ACTS|26|13|die media in via vidi rex de caelo supra splendorem solis circumfulsisse me lumen et eos qui mecum simul erant
ACTS|26|14|omnesque nos cum decidissemus in terram audivi vocem loquentem mihi hebraica lingua Saule Saule quid me persequeris durum est tibi contra stimulum calcitrare
ACTS|26|15|ego autem dixi quis es Domine Dominus autem dixit ego sum Iesus quem tu persequeris
ACTS|26|16|sed exsurge et sta super pedes tuos ad hoc enim apparui tibi ut constituam te ministrum et testem eorum quae vidisti et eorum quibus apparebo tibi
ACTS|26|17|eripiens te de populo et gentibus in quas nunc ego mitto te
ACTS|26|18|aperire oculos eorum ut convertantur a tenebris ad lucem et de potestate Satanae ad Deum ut accipiant remissionem peccatorum et sortem inter sanctos per fidem quae est in me
ACTS|26|19|unde rex Agrippa non fui incredulus caelestis visionis
ACTS|26|20|sed his qui sunt Damasci primum et Hierosolymis et in omnem regionem Iudaeae et gentibus adnuntiabam ut paenitentiam agerent et converterentur ad Deum digna paenitentiae opera facientes
ACTS|26|21|hac ex causa me Iudaei cum essem in templo conprehensum temptabant interficere
ACTS|26|22|auxilio autem adiutus Dei usque in hodiernum diem sto testificans minori atque maiori nihil extra dicens quam ea quae prophetae sunt locuti futura esse et Moses
ACTS|26|23|si passibilis Christus si primus ex resurrectione mortuorum lumen adnuntiaturus est populo et gentibus
ACTS|26|24|haec loquente eo et rationem reddente Festus magna voce dixit insanis Paule multae te litterae ad insaniam convertunt
ACTS|26|25|at Paulus non insanio inquit optime Feste sed veritatis et sobrietatis verba eloquor
ACTS|26|26|scit enim de his rex ad quem et constanter loquor latere enim eum nihil horum arbitror neque enim in angulo quicquam horum gestum est
ACTS|26|27|credis rex Agrippa prophetis scio quia credis
ACTS|26|28|Agrippa autem ad Paulum in modico suades me Christianum fieri
ACTS|26|29|et Paulus opto apud Deum et in modico et in magno non tantum te sed et omnes hos qui audiunt hodie fieri tales qualis et ego sum exceptis vinculis his
ACTS|26|30|et exsurrexit rex et praeses et Bernice et qui adsidebant eis
ACTS|26|31|et cum secessissent loquebantur ad invicem dicentes quia nihil morte aut vinculorum dignum quid facit homo iste
ACTS|26|32|Agrippa autem Festo dixit dimitti poterat homo hic si non appellasset Caesarem
ACTS|27|1|ut autem iudicatum est eum navigare in Italiam et tradi Paulum cum reliquis custodiis centurioni nomine Iulio cohortis Augustae
ACTS|27|2|ascendentes autem navem hadrumetinam incipientem navigare circa Asiae loca sustulimus perseverante nobiscum Aristarcho Macedone Thessalonicense
ACTS|27|3|sequenti autem die devenimus Sidonem humane autem tractans Iulius Paulum permisit ad amicos ire et curam sui agere
ACTS|27|4|et inde cum sustulissemus subnavigavimus Cypro propterea quod essent venti contrarii
ACTS|27|5|et pelagus Ciliciae et Pamphiliae navigantes venimus Lystram quae est Lyciae
ACTS|27|6|et ibi inveniens centurio navem alexandrinam navigantem in Italiam transposuit nos in eam
ACTS|27|7|et cum multis diebus tarde navigaremus et vix devenissemus contra Cnidum prohibente nos vento adnavigavimus Cretae secundum Salmonem
ACTS|27|8|et vix iuxta navigantes venimus in locum quendam qui vocatur Boni portus cui iuxta erat civitas Thalassa
ACTS|27|9|multo autem tempore peracto et cum iam non esset tuta navigatio eo quod et ieiunium iam praeterisset consolabatur Paulus
ACTS|27|10|dicens eis viri video quoniam cum iniuria et multo damno non solum oneris et navis sed etiam animarum nostrarum incipit esse navigatio
ACTS|27|11|centurio autem gubernatori et nauclerio magis credebat quam his quae a Paulo dicebantur
ACTS|27|12|et cum aptus portus non esset ad hiemandum plurimi statuerunt consilium navigare inde si quo modo possent devenientes Phoenice hiemare portum Cretae respicientem ad africum et ad chorum
ACTS|27|13|adspirante autem austro aestimantes propositum se tenere cum sustulissent de Asson legebant Cretam
ACTS|27|14|non post multum autem misit se contra ipsam ventus typhonicus qui vocatur euroaquilo
ACTS|27|15|cumque arrepta esset navis et non posset conari in ventum data nave flatibus ferebamur
ACTS|27|16|insulam autem quandam decurrentes quae vocatur Caudam potuimus vix obtinere scapham
ACTS|27|17|qua sublata adiutoriis utebantur accingentes navem timentes ne in Syrtim inciderent submisso vase sic ferebantur
ACTS|27|18|valide autem nobis tempestate iactatis sequenti die iactum fecerunt
ACTS|27|19|et tertia die suis manibus armamenta navis proiecerunt
ACTS|27|20|neque sole autem neque sideribus apparentibus per plures dies et tempestate non exigua inminente iam ablata erat spes omnis salutis nostrae
ACTS|27|21|et cum multa ieiunatio fuisset tunc stans Paulus in medio eorum dixit oportebat quidem o viri audito me non tollere a Creta lucrique facere iniuriam hanc et iacturam
ACTS|27|22|et nunc suadeo vobis bono animo esse amissio enim nullius animae erit ex vobis praeterquam navis
ACTS|27|23|adstitit enim mihi hac nocte angelus Dei cuius sum ego et cui deservio
ACTS|27|24|dicens ne timeas Paule Caesari te oportet adsistere et ecce donavit tibi Deus omnes qui navigant tecum
ACTS|27|25|propter quod bono animo estote viri credo enim Deo quia sic erit quemadmodum dictum est mihi
ACTS|27|26|in insulam autem quandam oportet nos devenire
ACTS|27|27|sed posteaquam quartadecima nox supervenit navigantibus nobis in Hadria circa mediam noctem suspicabantur nautae apparere sibi aliquam regionem
ACTS|27|28|qui submittentes invenerunt passus viginti et pusillum inde separati invenerunt passus quindecim
ACTS|27|29|timentes autem ne in aspera loca incideremus de puppi mittentes anchoras quattuor optabant diem fieri
ACTS|27|30|nautis vero quaerentibus fugere de navi cum misissent scapham in mare sub obtentu quasi a prora inciperent anchoras extendere
ACTS|27|31|dixit Paulus centurioni et militibus nisi hii in navi manserint vos salvi fieri non potestis
ACTS|27|32|tunc absciderunt milites funes scaphae et passi sunt eam excidere
ACTS|27|33|et cum lux inciperet fieri rogabat Paulus omnes sumere cibum dicens quartadecima hodie die expectantes ieiuni permanetis nihil accipientes
ACTS|27|34|propter quod rogo vos accipere cibum pro salute vestra quia nullius vestrum capillus de capite peribit
ACTS|27|35|et cum haec dixisset sumens panem gratias egit Deo in conspectu omnium et cum fregisset coepit manducare
ACTS|27|36|animaequiores autem facti omnes et ipsi adsumpserunt cibum
ACTS|27|37|eramus vero universae animae in navi ducentae septuaginta sex
ACTS|27|38|et satiati cibo adleviabant navem iactantes triticum in mare
ACTS|27|39|cum autem dies factus esset terram non agnoscebant sinum vero quendam considerabant habentem litus in quem cogitabant si possent eicere navem
ACTS|27|40|et cum anchoras abstulissent committebant se mari simul laxantes iuncturas gubernaculorum et levato artemone secundum flatum aurae tendebant ad litus
ACTS|27|41|et cum incidissemus in locum bithalassum inpegerunt navem et prora quidem fixa manebat inmobilis puppis vero solvebatur a vi maris
ACTS|27|42|militum autem consilium fuit ut custodias occiderent ne quis cum enatasset effugeret
ACTS|27|43|centurio autem volens servare Paulum prohibuit fieri iussitque eos qui possent natare mittere se primos et evadere et ad terram exire
ACTS|27|44|et ceteros alios in tabulis ferebant quosdam super ea quae de navi essent et sic factum est ut omnes animae evaderent ad terram
ACTS|28|1|et cum evasissemus tunc cognovimus quia Militene insula vocatur barbari vero praestabant non modicam humanitatem nobis
ACTS|28|2|accensa enim pyra reficiebant nos omnes propter imbrem qui inminebat et frigus
ACTS|28|3|cum congregasset autem Paulus sarmentorum aliquantam multitudinem et inposuisset super ignem vipera a calore cum processisset invasit manum eius
ACTS|28|4|ut vero viderunt barbari pendentem bestiam de manu eius ad invicem dicebant utique homicida est homo hic qui cum evaserit de mari Ultio non sinit vivere
ACTS|28|5|et ille quidem excutiens bestiam in ignem nihil mali passus est
ACTS|28|6|at illi existimabant eum in tumorem convertendum et subito casurum et mori diu autem illis sperantibus et videntibus nihil mali in eo fieri convertentes se dicebant eum esse deum
ACTS|28|7|in locis autem illis erant praedia principis insulae nomine Publii qui nos suscipiens triduo benigne exhibuit
ACTS|28|8|contigit autem patrem Publii febribus et dysenteria vexatum iacere ad quem Paulus intravit et cum orasset et inposuisset ei manus salvavit eum
ACTS|28|9|quo facto et omnes qui in insula habebant infirmitates accedebant et curabantur
ACTS|28|10|qui etiam multis honoribus nos honoraverunt et navigantibus inposuerunt quae necessaria erant
ACTS|28|11|post menses autem tres navigavimus in nave alexandrina quae in insula hiemaverat cui erat insigne Castorum
ACTS|28|12|et cum venissemus Syracusam mansimus ibi triduo
ACTS|28|13|inde circumlegentes devenimus Regium et post unum diem flante austro secunda die venimus Puteolos
ACTS|28|14|ubi inventis fratribus rogati sumus manere apud eos dies septem et sic venimus Romam
ACTS|28|15|et inde cum audissent fratres occurrerunt nobis usque ad Appii Forum et Tribus Tabernis quos cum vidisset Paulus gratias agens Deo accepit fiduciam
ACTS|28|16|cum venissemus autem Romam permissum est Paulo manere sibimet cum custodiente se milite
ACTS|28|17|post tertium autem diem convocavit primos Iudaeorum cumque convenissent dicebat eis ego viri fratres nihil adversus plebem faciens aut morem paternum vinctus ab Hierosolymis traditus sum in manus Romanorum
ACTS|28|18|qui cum interrogationem de me habuissent voluerunt me dimittere eo quod nulla causa esset mortis in me
ACTS|28|19|contradicentibus autem Iudaeis coactus sum appellare Caesarem non quasi gentem meam habens aliquid accusare
ACTS|28|20|propter hanc igitur causam rogavi vos videre et adloqui propter spem enim Israhel catena hac circumdatus sum
ACTS|28|21|at illi dixerunt ad eum nos neque litteras accepimus de te a Iudaea neque adveniens aliquis fratrum nuntiavit aut locutus est quid de te malum
ACTS|28|22|rogamus autem a te audire quae sentis nam de secta hac notum est nobis quia ubique ei contradicitur
ACTS|28|23|cum constituissent autem illi diem venerunt ad eum in hospitium plures quibus exponebat testificans regnum Dei suadensque eos de Iesu ex lege Mosi et prophetis a mane usque ad vesperam
ACTS|28|24|et quidam credebant his quae dicebantur quidam vero non credebant
ACTS|28|25|cumque invicem non essent consentientes discedebant dicente Paulo unum verbum quia bene Spiritus Sanctus locutus est per Esaiam prophetam ad patres nostros
ACTS|28|26|dicens vade ad populum istum et dic aure audietis et non intellegetis et videntes videbitis et non perspicietis
ACTS|28|27|incrassatum est enim cor populi huius et auribus graviter audierunt et oculos suos conpresserunt ne forte videant oculis et auribus audiant et corde intellegant et convertantur et sanem illos
ACTS|28|28|notum ergo sit vobis quoniam gentibus missum est hoc salutare Dei ipsi et audient
ACTS|28|29|
ACTS|28|30|mansit autem biennio toto in suo conducto et suscipiebat omnes qui ingrediebantur ad eum
ACTS|28|31|praedicans regnum Dei et docens quae sunt de Domino Iesu Christo cum omni fiducia sine prohibitione
ROM|1|1|Paulus servus Christi Iesu vocatus apostolus segregatus in evangelium Dei
ROM|1|2|quod ante promiserat per prophetas suos in scripturis sanctis
ROM|1|3|de Filio suo qui factus est ex semine David secundum carnem
ROM|1|4|qui praedestinatus est Filius Dei in virtute secundum Spiritum sanctificationis ex resurrectione mortuorum Iesu Christi Domini nostri
ROM|1|5|per quem accepimus gratiam et apostolatum ad oboediendum fidei in omnibus gentibus pro nomine eius
ROM|1|6|in quibus estis et vos vocati Iesu Christi
ROM|1|7|omnibus qui sunt Romae dilectis Dei vocatis sanctis gratia vobis et pax a Deo Patre nostro et Domino Iesu Christo
ROM|1|8|primum quidem gratias ago Deo meo per Iesum Christum pro omnibus vobis quia fides vestra adnuntiatur in universo mundo
ROM|1|9|testis enim mihi est Deus cui servio in spiritu meo in evangelio Filii eius quod sine intermissione memoriam vestri facio
ROM|1|10|semper in orationibus meis obsecrans si quo modo tandem aliquando prosperum iter habeam in voluntate Dei veniendi ad vos
ROM|1|11|desidero enim videre vos ut aliquid inpertiar gratiae vobis spiritalis ad confirmandos vos
ROM|1|12|id est simul consolari in vobis per eam quae invicem est fidem vestram atque meam
ROM|1|13|nolo autem vos ignorare fratres quia saepe proposui venire ad vos et prohibitus sum usque adhuc ut aliquem fructum habeam et in vobis sicut et in ceteris gentibus
ROM|1|14|Graecis ac barbaris sapientibus et insipientibus debitor sum
ROM|1|15|ita quod in me promptum est et vobis qui Romae estis evangelizare
ROM|1|16|non enim erubesco evangelium virtus enim Dei est in salutem omni credenti Iudaeo primum et Graeco
ROM|1|17|iustitia enim Dei in eo revelatur ex fide in fidem sicut scriptum est iustus autem ex fide vivit
ROM|1|18|revelatur enim ira Dei de caelo super omnem impietatem et iniustitiam hominum eorum qui veritatem in iniustitiam detinent
ROM|1|19|quia quod notum est Dei manifestum est in illis Deus enim illis manifestavit
ROM|1|20|invisibilia enim ipsius a creatura mundi per ea quae facta sunt intellecta conspiciuntur sempiterna quoque eius virtus et divinitas ut sint inexcusabiles
ROM|1|21|quia cum cognovissent Deum non sicut Deum glorificaverunt aut gratias egerunt sed evanuerunt in cogitationibus suis et obscuratum est insipiens cor eorum
ROM|1|22|dicentes enim se esse sapientes stulti facti sunt
ROM|1|23|et mutaverunt gloriam incorruptibilis Dei in similitudinem imaginis corruptibilis hominis et volucrum et quadrupedum et serpentium
ROM|1|24|propter quod tradidit illos Deus in desideria cordis eorum in inmunditiam ut contumeliis adficiant corpora sua in semet ipsis
ROM|1|25|qui commutaverunt veritatem Dei in mendacio et coluerunt et servierunt creaturae potius quam creatori qui est benedictus in saecula amen
ROM|1|26|propterea tradidit illos Deus in passiones ignominiae nam feminae eorum inmutaverunt naturalem usum in eum usum qui est contra naturam
ROM|1|27|similiter autem et masculi relicto naturali usu feminae exarserunt in desideriis suis in invicem masculi in masculos turpitudinem operantes et mercedem quam oportuit erroris sui in semet ipsis recipientes
ROM|1|28|et sicut non probaverunt Deum habere in notitia tradidit eos Deus in reprobum sensum ut faciant quae non conveniunt
ROM|1|29|repletos omni iniquitate malitia fornicatione avaritia nequitia plenos invidia homicidio contentione dolo malignitate susurrones
ROM|1|30|detractores Deo odibiles contumeliosos superbos elatos inventores malorum parentibus non oboedientes
ROM|1|31|insipientes inconpositos sine affectione absque foedere sine misericordia
ROM|1|32|qui cum iustitiam Dei cognovissent non intellexerunt quoniam qui talia agunt digni sunt morte non solum ea faciunt sed et consentiunt facientibus
ROM|2|1|propter quod inexcusabilis es o homo omnis qui iudicas in quo enim iudicas alterum te ipsum condemnas eadem enim agis qui iudicas
ROM|2|2|scimus enim quoniam iudicium Dei est secundum veritatem in eos qui talia agunt
ROM|2|3|existimas autem hoc o homo qui iudicas eos qui talia agunt et facis ea quia tu effugies iudicium Dei
ROM|2|4|an divitias bonitatis eius et patientiae et longanimitatis contemnis ignorans quoniam benignitas Dei ad paenitentiam te adducit
ROM|2|5|secundum duritiam autem tuam et inpaenitens cor thesaurizas tibi iram in die irae et revelationis iusti iudicii Dei
ROM|2|6|qui reddet unicuique secundum opera eius
ROM|2|7|his quidem qui secundum patientiam boni operis gloriam et honorem et incorruptionem quaerentibus vitam aeternam
ROM|2|8|his autem qui ex contentione et qui non adquiescunt veritati credunt autem iniquitati ira et indignatio
ROM|2|9|tribulatio et angustia in omnem animam hominis operantis malum Iudaei primum et Graeci
ROM|2|10|gloria autem et honor et pax omni operanti bonum Iudaeo primum et Graeco
ROM|2|11|non est enim personarum acceptio apud Deum
ROM|2|12|quicumque enim sine lege peccaverunt sine lege et peribunt et quicumque in lege peccaverunt per legem iudicabuntur
ROM|2|13|non enim auditores legis iusti sunt apud Deum sed factores legis iustificabuntur
ROM|2|14|cum enim gentes quae legem non habent naturaliter quae legis sunt faciunt eiusmodi legem non habentes ipsi sibi sunt lex
ROM|2|15|qui ostendunt opus legis scriptum in cordibus suis testimonium reddente illis conscientia ipsorum et inter se invicem cogitationum accusantium aut etiam defendentium
ROM|2|16|in die cum iudicabit Deus occulta hominum secundum evangelium meum per Iesum Christum
ROM|2|17|si autem tu Iudaeus cognominaris et requiescis in lege et gloriaris in Deo
ROM|2|18|et nosti voluntatem et probas utiliora instructus per legem
ROM|2|19|confidis te ipsum ducem esse caecorum lumen eorum qui in tenebris sunt
ROM|2|20|eruditorem insipientium magistrum infantium habentem formam scientiae et veritatis in lege
ROM|2|21|qui ergo alium doces te ipsum non doces qui praedicas non furandum furaris
ROM|2|22|qui dicis non moechandum moecharis qui abominaris idola sacrilegium facis
ROM|2|23|qui in lege gloriaris per praevaricationem legis Deum inhonoras
ROM|2|24|nomen enim Dei per vos blasphematur inter gentes sicut scriptum est
ROM|2|25|circumcisio quidem prodest si legem observes si autem praevaricator legis sis circumcisio tua praeputium facta est
ROM|2|26|si igitur praeputium iustitias legis custodiat nonne praeputium illius in circumcisionem reputabitur
ROM|2|27|et iudicabit quod ex natura est praeputium legem consummans te qui per litteram et circumcisionem praevaricator legis es
ROM|2|28|non enim qui in manifesto Iudaeus est neque quae in manifesto in carne circumcisio
ROM|2|29|sed qui in abscondito Iudaeus et circumcisio cordis in spiritu non littera cuius laus non ex hominibus sed ex Deo est
ROM|3|1|quid ergo amplius est Iudaeo aut quae utilitas circumcisionis
ROM|3|2|multum per omnem modum primum quidem quia credita sunt illis eloquia Dei
ROM|3|3|quid enim si quidam illorum non crediderunt numquid incredulitas illorum fidem Dei evacuabit absit
ROM|3|4|est autem Deus verax omnis autem homo mendax sicut scriptum est ut iustificeris in sermonibus tuis et vincas cum iudicaris
ROM|3|5|si autem iniquitas nostra iustitiam Dei commendat quid dicemus numquid iniquus Deus qui infert iram secundum hominem dico
ROM|3|6|absit alioquin quomodo iudicabit Deus mundum
ROM|3|7|si enim veritas Dei in meo mendacio abundavit in gloriam ipsius quid adhuc et ego tamquam peccator iudicor
ROM|3|8|et non sicut blasphemamur et sicut aiunt nos quidam dicere faciamus mala ut veniant bona quorum damnatio iusta est
ROM|3|9|quid igitur praecellimus eos nequaquam causati enim sumus Iudaeos et Graecos omnes sub peccato esse
ROM|3|10|sicut scriptum est quia non est iustus quisquam
ROM|3|11|non est intellegens non est requirens Deum
ROM|3|12|omnes declinaverunt simul inutiles facti sunt non est qui faciat bonum non est usque ad unum
ROM|3|13|sepulchrum patens est guttur eorum linguis suis dolose agebant venenum aspidum sub labiis eorum
ROM|3|14|quorum os maledictione et amaritudine plenum est
ROM|3|15|veloces pedes eorum ad effundendum sanguinem
ROM|3|16|contritio et infelicitas in viis eorum
ROM|3|17|et viam pacis non cognoverunt
ROM|3|18|non est timor Dei ante oculos eorum
ROM|3|19|scimus autem quoniam quaecumque lex loquitur his qui in lege sunt loquitur ut omne os obstruatur et subditus fiat omnis mundus Deo
ROM|3|20|quia ex operibus legis non iustificabitur omnis caro coram illo per legem enim cognitio peccati
ROM|3|21|nunc autem sine lege iustitia Dei manifestata est testificata a lege et prophetis
ROM|3|22|iustitia autem Dei per fidem Iesu Christi super omnes qui credunt non enim est distinctio
ROM|3|23|omnes enim peccaverunt et egent gloriam Dei
ROM|3|24|iustificati gratis per gratiam ipsius per redemptionem quae est in Christo Iesu
ROM|3|25|quem proposuit Deus propitiationem per fidem in sanguine ipsius ad ostensionem iustitiae suae propter remissionem praecedentium delictorum
ROM|3|26|in sustentatione Dei ad ostensionem iustitiae eius in hoc tempore ut sit ipse iustus et iustificans eum qui ex fide est Iesu
ROM|3|27|ubi est ergo gloriatio exclusa est per quam legem factorum non sed per legem fidei
ROM|3|28|arbitramur enim iustificari hominem per fidem sine operibus legis
ROM|3|29|an Iudaeorum Deus tantum nonne et gentium immo et gentium
ROM|3|30|quoniam quidem unus Deus qui iustificabit circumcisionem ex fide et praeputium per fidem
ROM|3|31|legem ergo destruimus per fidem absit sed legem statuimus
ROM|4|1|quid ergo dicemus invenisse Abraham patrem nostrum secundum carnem
ROM|4|2|si enim Abraham ex operibus iustificatus est habet gloriam sed non apud Deum
ROM|4|3|quid enim scriptura dicit credidit Abraham Deo et reputatum est illi ad iustitiam
ROM|4|4|ei autem qui operatur merces non inputatur secundum gratiam sed secundum debitum
ROM|4|5|ei vero qui non operatur credenti autem in eum qui iustificat impium reputatur fides eius ad iustitiam
ROM|4|6|sicut et David dicit beatitudinem hominis cui Deus accepto fert iustitiam sine operibus
ROM|4|7|beati quorum remissae sunt iniquitates et quorum tecta sunt peccata
ROM|4|8|beatus vir cui non inputabit Dominus peccatum
ROM|4|9|beatitudo ergo haec in circumcisione an etiam in praeputio dicimus enim quia reputata est Abrahae fides ad iustitiam
ROM|4|10|quomodo ergo reputata est in circumcisione an in praeputio non in circumcisione sed in praeputio
ROM|4|11|et signum accepit circumcisionis signaculum iustitiae fidei quae est in praeputio ut sit pater omnium credentium per praeputium ut reputetur et illis ad iustitiam
ROM|4|12|et sit pater circumcisionis non his tantum qui sunt ex circumcisione sed et his qui sectantur vestigia quae est in praeputio fidei patris nostri Abrahae
ROM|4|13|non enim per legem promissio Abrahae aut semini eius ut heres esset mundi sed per iustitiam fidei
ROM|4|14|si enim qui ex lege heredes sunt exinanita est fides abolita est promissio
ROM|4|15|lex enim iram operatur ubi enim non est lex nec praevaricatio
ROM|4|16|ideo ex fide ut secundum gratiam ut firma sit promissio omni semini non ei qui ex lege est solum sed et ei qui ex fide est Abrahae qui est pater omnium nostrum
ROM|4|17|sicut scriptum est quia patrem multarum gentium posui te ante Deum cui credidit qui vivificat mortuos et vocat quae non sunt tamquam ea quae sunt
ROM|4|18|qui contra spem in spem credidit ut fieret pater multarum gentium secundum quod dictum est sic erit semen tuum
ROM|4|19|et non infirmatus fide consideravit corpus suum emortuum cum fere centum annorum esset et emortuam vulvam Sarrae
ROM|4|20|in repromissione etiam Dei non haesitavit diffidentia sed confortatus est fide dans gloriam Deo
ROM|4|21|plenissime sciens quia quaecumque promisit potens est et facere
ROM|4|22|ideo et reputatum est illi ad iustitiam
ROM|4|23|non est autem scriptum tantum propter ipsum quia reputatum est illi
ROM|4|24|sed et propter nos quibus reputabitur credentibus in eum qui suscitavit Iesum Dominum nostrum a mortuis
ROM|4|25|qui traditus est propter delicta nostra et resurrexit propter iustificationem nostram
ROM|5|1|iustificati igitur ex fide pacem habeamus ad Deum per Dominum nostrum Iesum Christum
ROM|5|2|per quem et accessum habemus fide in gratiam istam in qua stamus et gloriamur in spe gloriae filiorum Dei
ROM|5|3|non solum autem sed et gloriamur in tribulationibus scientes quod tribulatio patientiam operatur
ROM|5|4|patientia autem probationem probatio vero spem
ROM|5|5|spes autem non confundit quia caritas Dei diffusa est in cordibus nostris per Spiritum Sanctum qui datus est nobis
ROM|5|6|ut quid enim Christus cum adhuc infirmi essemus secundum tempus pro impiis mortuus est
ROM|5|7|vix enim pro iusto quis moritur nam pro bono forsitan quis et audeat mori
ROM|5|8|commendat autem suam caritatem Deus in nos quoniam cum adhuc peccatores essemus
ROM|5|9|Christus pro nobis mortuus est multo igitur magis iustificati nunc in sanguine ipsius salvi erimus ab ira per ipsum
ROM|5|10|si enim cum inimici essemus reconciliati sumus Deo per mortem Filii eius multo magis reconciliati salvi erimus in vita ipsius
ROM|5|11|non solum autem sed et gloriamur in Deo per Dominum nostrum Iesum Christum per quem nunc reconciliationem accepimus
ROM|5|12|propterea sicut per unum hominem in hunc mundum peccatum intravit et per peccatum mors et ita in omnes homines mors pertransiit in quo omnes peccaverunt
ROM|5|13|usque ad legem enim peccatum erat in mundo peccatum autem non inputatur cum lex non est
ROM|5|14|sed regnavit mors ab Adam usque ad Mosen etiam in eos qui non peccaverunt in similitudinem praevaricationis Adae qui est forma futuri
ROM|5|15|sed non sicut delictum ita et donum si enim unius delicto multi mortui sunt multo magis gratia Dei et donum in gratiam unius hominis Iesu Christi in plures abundavit
ROM|5|16|et non sicut per unum peccantem ita et donum nam iudicium ex uno in condemnationem gratia autem ex multis delictis in iustificationem
ROM|5|17|si enim in unius delicto mors regnavit per unum multo magis abundantiam gratiae et donationis et iustitiae accipientes in vita regnabunt per unum Iesum Christum
ROM|5|18|igitur sicut per unius delictum in omnes homines in condemnationem sic et per unius iustitiam in omnes homines in iustificationem vitae
ROM|5|19|sicut enim per inoboedientiam unius hominis peccatores constituti sunt multi ita et per unius oboeditionem iusti constituentur multi
ROM|5|20|lex autem subintravit ut abundaret delictum ubi autem abundavit delictum superabundavit gratia
ROM|5|21|ut sicut regnavit peccatum in morte ita et gratia regnet per iustitiam in vitam aeternam per Iesum Christum Dominum nostrum
ROM|6|1|quid ergo dicemus permanebimus in peccato ut gratia abundet
ROM|6|2|absit qui enim mortui sumus peccato quomodo adhuc vivemus in illo
ROM|6|3|an ignoratis quia quicumque baptizati sumus in Christo Iesu in morte ipsius baptizati sumus
ROM|6|4|consepulti enim sumus cum illo per baptismum in mortem ut quomodo surrexit Christus a mortuis per gloriam Patris ita et nos in novitate vitae ambulemus
ROM|6|5|si enim conplantati facti sumus similitudini mortis eius simul et resurrectionis erimus
ROM|6|6|hoc scientes quia vetus homo noster simul crucifixus est ut destruatur corpus peccati ut ultra non serviamus peccato
ROM|6|7|qui enim mortuus est iustificatus est a peccato
ROM|6|8|si autem mortui sumus cum Christo credimus quia simul etiam vivemus cum Christo
ROM|6|9|scientes quod Christus surgens ex mortuis iam non moritur mors illi ultra non dominabitur
ROM|6|10|quod enim mortuus est peccato mortuus est semel quod autem vivit vivit Deo
ROM|6|11|ita et vos existimate vos mortuos quidem esse peccato viventes autem Deo in Christo Iesu
ROM|6|12|non ergo regnet peccatum in vestro mortali corpore ut oboediatis concupiscentiis eius
ROM|6|13|sed neque exhibeatis membra vestra arma iniquitatis peccato sed exhibete vos Deo tamquam ex mortuis viventes et membra vestra arma iustitiae Deo
ROM|6|14|peccatum enim vobis non dominabitur non enim sub lege estis sed sub gratia
ROM|6|15|quid ergo peccavimus quoniam non sumus sub lege sed sub gratia absit
ROM|6|16|nescitis quoniam cui exhibetis vos servos ad oboediendum servi estis eius cui oboeditis sive peccati sive oboeditionis ad iustitiam
ROM|6|17|gratias autem Deo quod fuistis servi peccati oboedistis autem ex corde in eam formam doctrinae in qua traditi estis
ROM|6|18|liberati autem a peccato servi facti estis iustitiae
ROM|6|19|humanum dico propter infirmitatem carnis vestrae sicut enim exhibuistis membra vestra servire inmunditiae et iniquitati ad iniquitatem ita nunc exhibete membra vestra servire iustitiae in sanctificationem
ROM|6|20|cum enim servi essetis peccati liberi fuistis iustitiae
ROM|6|21|quem ergo fructum habuistis tunc in quibus nunc erubescitis nam finis illorum mors est
ROM|6|22|nunc vero liberati a peccato servi autem facti Deo habetis fructum vestrum in sanctificationem finem vero vitam aeternam
ROM|6|23|stipendia enim peccati mors gratia autem Dei vita aeterna in Christo Iesu Domino nostro
ROM|7|1|an ignoratis fratres scientibus enim legem loquor quia lex in homine dominatur quanto tempore vivit
ROM|7|2|nam quae sub viro est mulier vivente viro alligata est legi si autem mortuus fuerit vir soluta est a lege viri
ROM|7|3|igitur vivente viro vocabitur adultera si fuerit cum alio viro si autem mortuus fuerit vir eius liberata est a lege ut non sit adultera si fuerit cum alio viro
ROM|7|4|itaque fratres mei et vos mortificati estis legi per corpus Christi ut sitis alterius qui ex mortuis resurrexit ut fructificaremus Deo
ROM|7|5|cum enim essemus in carne passiones peccatorum quae per legem erant operabantur in membris nostris ut fructificarent morti
ROM|7|6|nunc autem soluti sumus a lege morientes in quo detinebamur ita ut serviamus in novitate spiritus et non in vetustate litterae
ROM|7|7|quid ergo dicemus lex peccatum est absit sed peccatum non cognovi nisi per legem nam concupiscentiam nesciebam nisi lex diceret non concupisces
ROM|7|8|occasione autem accepta peccatum per mandatum operatum est in me omnem concupiscentiam sine lege enim peccatum mortuum erat
ROM|7|9|ego autem vivebam sine lege aliquando sed cum venisset mandatum peccatum revixit
ROM|7|10|ego autem mortuus sum et inventum est mihi mandatum quod erat ad vitam hoc esse ad mortem
ROM|7|11|nam peccatum occasione accepta per mandatum seduxit me et per illud occidit
ROM|7|12|itaque lex quidem sancta et mandatum sanctum et iustum et bonum
ROM|7|13|quod ergo bonum est mihi factum est mors absit sed peccatum ut appareat peccatum per bonum mihi operatum est mortem ut fiat supra modum peccans peccatum per mandatum
ROM|7|14|scimus enim quod lex spiritalis est ego autem carnalis sum venundatus sub peccato
ROM|7|15|quod enim operor non intellego non enim quod volo hoc ago sed quod odi illud facio
ROM|7|16|si autem quod nolo illud facio consentio legi quoniam bona
ROM|7|17|nunc autem iam non ego operor illud sed quod habitat in me peccatum
ROM|7|18|scio enim quia non habitat in me hoc est in carne mea bonum nam velle adiacet mihi perficere autem bonum non invenio
ROM|7|19|non enim quod volo bonum hoc facio sed quod nolo malum hoc ago
ROM|7|20|si autem quod nolo illud facio non ego operor illud sed quod habitat in me peccatum
ROM|7|21|invenio igitur legem volenti mihi facere bonum quoniam mihi malum adiacet
ROM|7|22|condelector enim legi Dei secundum interiorem hominem
ROM|7|23|video autem aliam legem in membris meis repugnantem legi mentis meae et captivantem me in lege peccati quae est in membris meis
ROM|7|24|infelix ego homo quis me liberabit de corpore mortis huius
ROM|7|25|gratia Dei per Iesum Christum Dominum nostrum igitur ego ipse mente servio legi Dei carne autem legi peccati
ROM|8|1|nihil ergo nunc damnationis est his qui sunt in Christo Iesu qui non secundum carnem ambulant
ROM|8|2|lex enim Spiritus vitae in Christo Iesu liberavit me a lege peccati et mortis
ROM|8|3|nam quod inpossibile erat legis in quo infirmabatur per carnem Deus Filium suum mittens in similitudinem carnis peccati et de peccato damnavit peccatum in carne
ROM|8|4|ut iustificatio legis impleretur in nobis qui non secundum carnem ambulamus sed secundum Spiritum
ROM|8|5|qui enim secundum carnem sunt quae carnis sunt sapiunt qui vero secundum Spiritum quae sunt Spiritus sentiunt
ROM|8|6|nam prudentia carnis mors prudentia autem Spiritus vita et pax
ROM|8|7|quoniam sapientia carnis inimicitia est in Deum legi enim Dei non subicitur nec enim potest
ROM|8|8|qui autem in carne sunt Deo placere non possunt
ROM|8|9|vos autem in carne non estis sed in Spiritu si tamen Spiritus Dei habitat in vobis si quis autem Spiritum Christi non habet hic non est eius
ROM|8|10|si autem Christus in vobis est corpus quidem mortuum est propter peccatum spiritus vero vita propter iustificationem
ROM|8|11|quod si Spiritus eius qui suscitavit Iesum a mortuis habitat in vobis qui suscitavit Iesum Christum a mortuis vivificabit et mortalia corpora vestra propter inhabitantem Spiritum eius in vobis
ROM|8|12|ergo fratres debitores sumus non carni ut secundum carnem vivamus
ROM|8|13|si enim secundum carnem vixeritis moriemini si autem Spiritu facta carnis mortificatis vivetis
ROM|8|14|quicumque enim Spiritu Dei aguntur hii filii sunt Dei
ROM|8|15|non enim accepistis spiritum servitutis iterum in timore sed accepistis Spiritum adoptionis filiorum in quo clamamus Abba Pater
ROM|8|16|ipse Spiritus testimonium reddit spiritui nostro quod sumus filii Dei
ROM|8|17|si autem filii et heredes heredes quidem Dei coheredes autem Christi si tamen conpatimur ut et conglorificemur
ROM|8|18|existimo enim quod non sunt condignae passiones huius temporis ad futuram gloriam quae revelabitur in nobis
ROM|8|19|nam expectatio creaturae revelationem filiorum Dei expectat
ROM|8|20|vanitati enim creatura subiecta est non volens sed propter eum qui subiecit in spem
ROM|8|21|quia et ipsa creatura liberabitur a servitute corruptionis in libertatem gloriae filiorum Dei
ROM|8|22|scimus enim quod omnis creatura ingemescit et parturit usque adhuc
ROM|8|23|non solum autem illa sed et nos ipsi primitias Spiritus habentes et ipsi intra nos gemimus adoptionem filiorum expectantes redemptionem corporis nostri
ROM|8|24|spe enim salvi facti sumus spes autem quae videtur non est spes nam quod videt quis quid sperat
ROM|8|25|si autem quod non videmus speramus per patientiam expectamus
ROM|8|26|similiter autem et Spiritus adiuvat infirmitatem nostram nam quid oremus sicut oportet nescimus sed ipse Spiritus postulat pro nobis gemitibus inenarrabilibus
ROM|8|27|qui autem scrutatur corda scit quid desideret Spiritus quia secundum Deum postulat pro sanctis
ROM|8|28|scimus autem quoniam diligentibus Deum omnia cooperantur in bonum his qui secundum propositum vocati sunt sancti
ROM|8|29|nam quos praescivit et praedestinavit conformes fieri imaginis Filii eius ut sit ipse primogenitus in multis fratribus
ROM|8|30|quos autem praedestinavit hos et vocavit et quos vocavit hos et iustificavit quos autem iustificavit illos et glorificavit
ROM|8|31|quid ergo dicemus ad haec si Deus pro nobis quis contra nos
ROM|8|32|qui etiam Filio suo non pepercit sed pro nobis omnibus tradidit illum quomodo non etiam cum illo omnia nobis donabit
ROM|8|33|quis accusabit adversus electos Dei Deus qui iustificat
ROM|8|34|quis est qui condemnet Christus Iesus qui mortuus est immo qui resurrexit qui et est ad dexteram Dei qui etiam interpellat pro nobis
ROM|8|35|quis nos separabit a caritate Christi tribulatio an angustia an persecutio an fames an nuditas an periculum an gladius
ROM|8|36|sicut scriptum est quia propter te mortificamur tota die aestimati sumus ut oves occisionis
ROM|8|37|sed in his omnibus superamus propter eum qui dilexit nos
ROM|8|38|certus sum enim quia neque mors neque vita neque angeli neque principatus neque instantia neque futura neque fortitudines
ROM|8|39|neque altitudo neque profundum neque creatura alia poterit nos separare a caritate Dei quae est in Christo Iesu Domino nostro
ROM|9|1|veritatem dico in Christo non mentior testimonium mihi perhibente conscientia mea in Spiritu Sancto
ROM|9|2|quoniam tristitia est mihi magna et continuus dolor cordi meo
ROM|9|3|optabam enim ipse ego anathema esse a Christo pro fratribus meis qui sunt cognati mei secundum carnem
ROM|9|4|qui sunt Israhelitae quorum adoptio est filiorum et gloria et testamenta et legislatio et obsequium et promissa
ROM|9|5|quorum patres et ex quibus Christus secundum carnem qui est super omnia Deus benedictus in saecula amen
ROM|9|6|non autem quod exciderit verbum Dei non enim omnes qui ex Israhel hii sunt Israhel
ROM|9|7|neque quia semen sunt Abrahae omnes filii sed in Isaac vocabitur tibi semen
ROM|9|8|id est non qui filii carnis hii filii Dei sed qui filii sunt promissionis aestimantur in semine
ROM|9|9|promissionis enim verbum hoc est secundum hoc tempus veniam et erit Sarrae filius
ROM|9|10|non solum autem sed et Rebecca ex uno concubitum habens Isaac patre nostro
ROM|9|11|cum enim nondum nati fuissent aut aliquid egissent bonum aut malum ut secundum electionem propositum Dei maneret
ROM|9|12|non ex operibus sed ex vocante dictum est ei quia maior serviet minori
ROM|9|13|sicut scriptum est Iacob dilexi Esau autem odio habui
ROM|9|14|quid ergo dicemus numquid iniquitas apud Deum absit
ROM|9|15|Mosi enim dicit miserebor cuius misereor et misericordiam praestabo cuius miserebor
ROM|9|16|igitur non volentis neque currentis sed miserentis Dei
ROM|9|17|dicit enim scriptura Pharaoni quia in hoc ipsum excitavi te ut ostendam in te virtutem meam et ut adnuntietur nomen meum in universa terra
ROM|9|18|ergo cuius vult miseretur et quem vult indurat
ROM|9|19|dicis itaque mihi quid adhuc queritur voluntati enim eius quis resistit
ROM|9|20|o homo tu quis es qui respondeas Deo numquid dicit figmentum ei qui se finxit quid me fecisti sic
ROM|9|21|an non habet potestatem figulus luti ex eadem massa facere aliud quidem vas in honorem aliud vero in contumeliam
ROM|9|22|quod si volens Deus ostendere iram et notam facere potentiam suam sustinuit in multa patientia vasa irae aptata in interitum
ROM|9|23|ut ostenderet divitias gloriae suae in vasa misericordiae quae praeparavit in gloriam
ROM|9|24|quos et vocavit nos non solum ex Iudaeis sed etiam ex gentibus
ROM|9|25|sicut in Osee dicit vocabo non plebem meam plebem meam et non misericordiam consecutam misericordiam consecutam
ROM|9|26|et erit in loco ubi dictum est eis non plebs mea vos ibi vocabuntur filii Dei vivi
ROM|9|27|Esaias autem clamat pro Israhel si fuerit numerus filiorum Israhel tamquam harena maris reliquiae salvae fient
ROM|9|28|verbum enim consummans et brevians in aequitate quia verbum breviatum faciet Dominus super terram
ROM|9|29|et sicut praedixit Esaias nisi Dominus Sabaoth reliquisset nobis semen sicut Sodoma facti essemus et sicut Gomorra similes fuissemus
ROM|9|30|quid ergo dicemus quod gentes quae non sectabantur iustitiam adprehenderunt iustitiam iustitiam autem quae ex fide est
ROM|9|31|Israhel vero sectans legem iustitiae in legem iustitiae non pervenit
ROM|9|32|quare quia non ex fide sed quasi ex operibus offenderunt in lapidem offensionis
ROM|9|33|sicut scriptum est ecce pono in Sion lapidem offensionis et petram scandali et omnis qui credit in eum non confundetur
ROM|10|1|fratres voluntas quidem cordis mei et obsecratio ad Deum fit pro illis in salutem
ROM|10|2|testimonium enim perhibeo illis quod aemulationem Dei habent sed non secundum scientiam
ROM|10|3|ignorantes enim Dei iustitiam et suam quaerentes statuere iustitiae Dei non sunt subiecti
ROM|10|4|finis enim legis Christus ad iustitiam omni credenti
ROM|10|5|Moses enim scripsit quoniam iustitiam quae ex lege est qui fecerit homo vivet in ea
ROM|10|6|quae autem ex fide est iustitia sic dicit ne dixeris in corde tuo quis ascendit in caelum id est Christum deducere
ROM|10|7|aut quis descendit in abyssum hoc est Christum ex mortuis revocare
ROM|10|8|sed quid dicit prope est verbum in ore tuo et in corde tuo hoc est verbum fidei quod praedicamus
ROM|10|9|quia si confitearis in ore tuo Dominum Iesum et in corde tuo credideris quod Deus illum excitavit ex mortuis salvus eris
ROM|10|10|corde enim creditur ad iustitiam ore autem confessio fit in salutem
ROM|10|11|dicit enim scriptura omnis qui credit in illum non confundetur
ROM|10|12|non enim est distinctio Iudaei et Graeci nam idem Dominus omnium dives in omnes qui invocant illum
ROM|10|13|omnis enim quicumque invocaverit nomen Domini salvus erit
ROM|10|14|quomodo ergo invocabunt in quem non crediderunt aut quomodo credent ei quem non audierunt quomodo autem audient sine praedicante
ROM|10|15|quomodo vero praedicabunt nisi mittantur sicut scriptum est quam speciosi pedes evangelizantium pacem evangelizantium bona
ROM|10|16|sed non omnes oboedierunt evangelio Esaias enim dicit Domine quis credidit auditui nostro
ROM|10|17|ergo fides ex auditu auditus autem per verbum Christi
ROM|10|18|sed dico numquid non audierunt et quidem in omnem terram exiit sonus eorum et in fines orbis terrae verba eorum
ROM|10|19|sed dico numquid Israhel non cognovit primus Moses dicit ego ad aemulationem vos adducam in non gentem in gentem insipientem in iram vos mittam
ROM|10|20|Esaias autem audet et dicit inventus sum non quaerentibus me palam apparui his qui me non interrogabant
ROM|10|21|ad Israhel autem dicit tota die expandi manus meas ad populum non credentem et contradicentem
ROM|11|1|dico ergo numquid reppulit Deus populum suum absit nam et ego Israhelita sum ex semine Abraham tribu Beniamin
ROM|11|2|non reppulit Deus plebem suam quam praesciit an nescitis in Helia quid dicit scriptura quemadmodum interpellat Deum adversus Israhel
ROM|11|3|Domine prophetas tuos occiderunt altaria tua suffoderunt et ego relictus sum solus et quaerunt animam meam
ROM|11|4|sed quid dicit illi responsum divinum reliqui mihi septem milia virorum qui non curvaverunt genu Baal
ROM|11|5|sic ergo et in hoc tempore reliquiae secundum electionem gratiae factae sunt
ROM|11|6|si autem gratia non ex operibus alioquin gratia iam non est gratia
ROM|11|7|quid ergo quod quaerebat Israhel hoc non est consecutus electio autem consecuta est ceteri vero excaecati sunt
ROM|11|8|sicut scriptum est dedit illis Deus spiritum conpunctionis oculos ut non videant et aures ut non audiant usque in hodiernum diem
ROM|11|9|et David dicit fiat mensa eorum in laqueum et in captionem et in scandalum et in retributionem illis
ROM|11|10|obscurentur oculi eorum ne videant et dorsum illorum semper incurva
ROM|11|11|dico ergo numquid sic offenderunt ut caderent absit sed illorum delicto salus gentibus ut illos aemulentur
ROM|11|12|quod si delictum illorum divitiae sunt mundi et deminutio eorum divitiae gentium quanto magis plenitudo eorum
ROM|11|13|vobis enim dico gentibus quamdiu quidem ego sum gentium apostolus ministerium meum honorificabo
ROM|11|14|si quo modo ad aemulandum provocem carnem meam et salvos faciam aliquos ex illis
ROM|11|15|si enim amissio eorum reconciliatio est mundi quae adsumptio nisi vita ex mortuis
ROM|11|16|quod si delibatio sancta est et massa et si radix sancta et rami
ROM|11|17|quod si aliqui ex ramis fracti sunt tu autem cum oleaster esses insertus es in illis et socius radicis et pinguidinis olivae factus es
ROM|11|18|noli gloriari adversus ramos quod si gloriaris non tu radicem portas sed radix te
ROM|11|19|dices ergo fracti sunt rami ut ego inserar
ROM|11|20|bene propter incredulitatem fracti sunt tu autem fide stas noli altum sapere sed time
ROM|11|21|si enim Deus naturalibus ramis non pepercit ne forte nec tibi parcat
ROM|11|22|vide ergo bonitatem et severitatem Dei in eos quidem qui ceciderunt severitatem in te autem bonitatem Dei si permanseris in bonitate alioquin et tu excideris
ROM|11|23|sed et illi si non permanserint in incredulitate inserentur potens est enim Deus iterum inserere illos
ROM|11|24|nam si tu ex naturali excisus es oleastro et contra naturam insertus es in bonam olivam quanto magis hii secundum naturam inserentur suae olivae
ROM|11|25|nolo enim vos ignorare fratres mysterium hoc ut non sitis vobis ipsis sapientes quia caecitas ex parte contigit in Israhel donec plenitudo gentium intraret
ROM|11|26|et sic omnis Israhel salvus fieret sicut scriptum est veniet ex Sion qui eripiat avertet impietates ab Iacob
ROM|11|27|et hoc illis a me testamentum cum abstulero peccata eorum
ROM|11|28|secundum evangelium quidem inimici propter vos secundum electionem autem carissimi propter patres
ROM|11|29|sine paenitentia enim sunt dona et vocatio Dei
ROM|11|30|sicut enim aliquando et vos non credidistis Deo nunc autem misericordiam consecuti estis propter illorum incredulitatem
ROM|11|31|ita et isti nunc non crediderunt in vestram misericordiam ut et ipsi misericordiam consequantur
ROM|11|32|conclusit enim Deus omnia in incredulitatem ut omnium misereatur
ROM|11|33|o altitudo divitiarum sapientiae et scientiae Dei quam inconprehensibilia sunt iudicia eius et investigabiles viae eius
ROM|11|34|quis enim cognovit sensum Domini aut quis consiliarius eius fuit
ROM|11|35|aut quis prior dedit illi et retribuetur ei
ROM|11|36|quoniam ex ipso et per ipsum et in ipso omnia ipsi gloria in saecula amen
ROM|12|1|obsecro itaque vos fratres per misericordiam Dei ut exhibeatis corpora vestra hostiam viventem sanctam Deo placentem rationabile obsequium vestrum
ROM|12|2|et nolite conformari huic saeculo sed reformamini in novitate sensus vestri ut probetis quae sit voluntas Dei bona et placens et perfecta
ROM|12|3|dico enim per gratiam quae data est mihi omnibus qui sunt inter vos non plus sapere quam oportet sapere sed sapere ad sobrietatem unicuique sicut Deus divisit mensuram fidei
ROM|12|4|sicut enim in uno corpore multa membra habemus omnia autem membra non eundem actum habent
ROM|12|5|ita multi unum corpus sumus in Christo singuli autem alter alterius membra
ROM|12|6|habentes autem donationes secundum gratiam quae data est nobis differentes sive prophetiam secundum rationem fidei
ROM|12|7|sive ministerium in ministrando sive qui docet in doctrina
ROM|12|8|qui exhortatur in exhortando qui tribuit in simplicitate qui praeest in sollicitudine qui miseretur in hilaritate
ROM|12|9|dilectio sine simulatione odientes malum adherentes bono
ROM|12|10|caritatem fraternitatis invicem diligentes honore invicem praevenientes
ROM|12|11|sollicitudine non pigri spiritu ferventes Domino servientes
ROM|12|12|spe gaudentes in tribulatione patientes orationi instantes
ROM|12|13|necessitatibus sanctorum communicantes hospitalitatem sectantes
ROM|12|14|benedicite persequentibus benedicite et nolite maledicere
ROM|12|15|gaudere cum gaudentibus flere cum flentibus
ROM|12|16|id ipsum invicem sentientes non alta sapientes sed humilibus consentientes nolite esse prudentes apud vosmet ipsos
ROM|12|17|nulli malum pro malo reddentes providentes bona non tantum coram Deo sed etiam coram omnibus hominibus
ROM|12|18|si fieri potest quod ex vobis est cum omnibus hominibus pacem habentes
ROM|12|19|non vosmet ipsos defendentes carissimi sed date locum irae scriptum est enim mihi vindictam ego retribuam dicit Dominus
ROM|12|20|sed si esurierit inimicus tuus ciba illum si sitit potum da illi hoc enim faciens carbones ignis congeres super caput eius
ROM|12|21|noli vinci a malo sed vince in bono malum
ROM|13|1|omnis anima potestatibus sublimioribus subdita sit non est enim potestas nisi a Deo quae autem sunt a Deo ordinatae sunt
ROM|13|2|itaque qui resistit potestati Dei ordinationi resistit qui autem resistunt ipsi sibi damnationem adquirunt
ROM|13|3|nam principes non sunt timori boni operis sed mali vis autem non timere potestatem bonum fac et habebis laudem ex illa
ROM|13|4|Dei enim minister est tibi in bonum si autem male feceris time non enim sine causa gladium portat Dei enim minister est vindex in iram ei qui malum agit
ROM|13|5|ideo necessitate subditi estote non solum propter iram sed et propter conscientiam
ROM|13|6|ideo enim et tributa praestatis ministri enim Dei sunt in hoc ipsum servientes
ROM|13|7|reddite omnibus debita cui tributum tributum cui vectigal vectigal cui timorem timorem cui honorem honorem
ROM|13|8|nemini quicquam debeatis nisi ut invicem diligatis qui enim diligit proximum legem implevit
ROM|13|9|nam non adulterabis non occides non furaberis non concupisces et si quod est aliud mandatum in hoc verbo instauratur diliges proximum tuum tamquam te ipsum
ROM|13|10|dilectio proximo malum non operatur plenitudo ergo legis est dilectio
ROM|13|11|et hoc scientes tempus quia hora est iam nos de somno surgere nunc enim propior est nostra salus quam cum credidimus
ROM|13|12|nox praecessit dies autem adpropiavit abiciamus ergo opera tenebrarum et induamur arma lucis
ROM|13|13|sicut in die honeste ambulemus non in comesationibus et ebrietatibus non in cubilibus et inpudicitiis non in contentione et aemulatione
ROM|13|14|sed induite Dominum Iesum Christum et carnis curam ne feceritis in desideriis
ROM|14|1|infirmum autem in fide adsumite non in disceptationibus cogitationum
ROM|14|2|alius enim credit manducare omnia qui autem infirmus est holus manducat
ROM|14|3|is qui manducat non manducantem non spernat et qui non manducat manducantem non iudicet Deus enim illum adsumpsit
ROM|14|4|tu quis es qui iudices alienum servum suo domino stat aut cadit stabit autem potens est enim Deus statuere illum
ROM|14|5|nam alius iudicat diem plus inter diem alius iudicat omnem diem unusquisque in suo sensu abundet
ROM|14|6|qui sapit diem Domino sapit et qui manducat Domino manducat gratias enim agit Deo et qui non manducat Domino non manducat et gratias agit Deo
ROM|14|7|nemo enim nostrum sibi vivit et nemo sibi moritur
ROM|14|8|sive enim vivimus Domino vivimus sive morimur Domino morimur sive ergo vivimus sive morimur Domini sumus
ROM|14|9|in hoc enim Christus et mortuus est et revixit ut et mortuorum et vivorum dominetur
ROM|14|10|tu autem quid iudicas fratrem tuum aut tu quare spernis fratrem tuum omnes enim stabimus ante tribunal Dei
ROM|14|11|scriptum est enim vivo ego dicit Dominus quoniam mihi flectet omne genu et omnis lingua confitebitur Deo
ROM|14|12|itaque unusquisque nostrum pro se rationem reddet Deo
ROM|14|13|non ergo amplius invicem iudicemus sed hoc iudicate magis ne ponatis offendiculum fratri vel scandalum
ROM|14|14|scio et confido in Domino Iesu quia nihil commune per ipsum nisi ei qui existimat quid commune esse illi commune est
ROM|14|15|si enim propter cibum frater tuus contristatur iam non secundum caritatem ambulas noli cibo tuo illum perdere pro quo Christus mortuus est
ROM|14|16|non ergo blasphemetur bonum nostrum
ROM|14|17|non est regnum Dei esca et potus sed iustitia et pax et gaudium in Spiritu Sancto
ROM|14|18|qui enim in hoc servit Christo placet Deo et probatus est hominibus
ROM|14|19|itaque quae pacis sunt sectemur et quae aedificationis sunt in invicem
ROM|14|20|noli propter escam destruere opus Dei omnia quidem munda sunt sed malum est homini qui per offendiculum manducat
ROM|14|21|bonum est non manducare carnem et non bibere vinum neque in quo frater tuus offendit aut scandalizatur aut infirmatur
ROM|14|22|tu fidem habes penes temet ipsum habe coram Deo beatus qui non iudicat semet ipsum in eo quo probat
ROM|14|23|qui autem discernit si manducaverit damnatus est quia non ex fide omne autem quod non ex fide peccatum est
ROM|15|1|debemus autem nos firmiores inbecillitates infirmorum sustinere et non nobis placere
ROM|15|2|unusquisque vestrum proximo suo placeat in bonum ad aedificationem
ROM|15|3|etenim Christus non sibi placuit sed sicut scriptum est inproperia inproperantium tibi ceciderunt super me
ROM|15|4|quaecumque enim scripta sunt ad nostram doctrinam scripta sunt ut per patientiam et consolationem scripturarum spem habeamus
ROM|15|5|Deus autem patientiae et solacii det vobis id ipsum sapere in alterutrum secundum Iesum Christum
ROM|15|6|ut unianimes uno ore honorificetis Deum et Patrem Domini nostri Iesu Christi
ROM|15|7|propter quod suscipite invicem sicut et Christus suscepit vos in honorem Dei
ROM|15|8|dico enim Christum Iesum ministrum fuisse circumcisionis propter veritatem Dei ad confirmandas promissiones patrum
ROM|15|9|gentes autem super misericordiam honorare Deum sicut scriptum est propter hoc confitebor tibi in gentibus et nomini tuo cantabo
ROM|15|10|et iterum dicit laetamini gentes cum plebe eius
ROM|15|11|et iterum laudate omnes gentes Dominum et magnificate eum omnes populi
ROM|15|12|et rursus Esaias ait erit radix Iesse et qui exsurget regere gentes in eo gentes sperabunt
ROM|15|13|Deus autem spei repleat vos omni gaudio et pace in credendo ut abundetis in spe in virtute Spiritus Sancti
ROM|15|14|certus sum autem fratres mei et ego ipse de vobis quoniam et ipsi pleni estis dilectione repleti omni scientia ita ut possitis alterutrum monere
ROM|15|15|audacius autem scripsi vobis fratres ex parte tamquam in memoriam vos reducens propter gratiam quae data est mihi a Deo
ROM|15|16|ut sim minister Christi Iesu in gentibus sanctificans evangelium Dei ut fiat oblatio gentium accepta sanctificata in Spiritu Sancto
ROM|15|17|habeo igitur gloriam in Christo Iesu ad Deum
ROM|15|18|non enim audeo aliquid loqui eorum quae per me non effecit Christus in oboedientiam gentium verbo et factis
ROM|15|19|in virtute signorum et prodigiorum in virtute Spiritus Sancti ita ut ab Hierusalem per circuitum usque in Illyricum repleverim evangelium Christi
ROM|15|20|sic autem hoc praedicavi evangelium non ubi nominatus est Christus ne super alienum fundamentum aedificarem
ROM|15|21|sed sicut scriptum est quibus non est adnuntiatum de eo videbunt et qui non audierunt intellegent
ROM|15|22|propter quod et inpediebar plurimum venire ad vos
ROM|15|23|nunc vero ulterius locum non habens in his regionibus cupiditatem autem habens veniendi ad vos ex multis iam annis
ROM|15|24|cum in Hispaniam proficisci coepero spero quod praeteriens videam vos et a vobis deducar illuc si vobis primum ex parte fruitus fuero
ROM|15|25|nunc igitur proficiscar in Hierusalem ministrare sanctis
ROM|15|26|probaverunt enim Macedonia et Achaia conlationem aliquam facere in pauperes sanctorum qui sunt in Hierusalem
ROM|15|27|placuit enim eis et debitores sunt eorum nam si spiritalium eorum participes facti sunt gentiles debent et in carnalibus ministrare eis
ROM|15|28|hoc igitur cum consummavero et adsignavero eis fructum hunc proficiscar per vos in Hispaniam
ROM|15|29|scio autem quoniam veniens ad vos in abundantia benedictionis Christi veniam
ROM|15|30|obsecro igitur vos fratres per Dominum nostrum Iesum Christum et per caritatem Spiritus ut adiuvetis me in orationibus pro me ad Deum
ROM|15|31|ut liberer ab infidelibus qui sunt in Iudaea et obsequii mei oblatio accepta fiat in Hierosolyma sanctis
ROM|15|32|ut veniam ad vos in gaudio per voluntatem Dei et refrigerer vobiscum
ROM|15|33|Deus autem pacis sit cum omnibus vobis amen
ROM|16|1|commendo autem vobis Phoebem sororem nostram quae est in ministerio ecclesiae quae est Cenchris
ROM|16|2|ut eam suscipiatis in Domino digne sanctis et adsistatis ei in quocumque negotio vestri indiguerit etenim ipsa quoque adstitit multis et mihi ipsi
ROM|16|3|salutate Priscam et Aquilam adiutores meos in Christo Iesu
ROM|16|4|qui pro anima mea suas cervices subposuerunt quibus non solus ego gratias ago sed et cunctae ecclesiae gentium
ROM|16|5|et domesticam eorum ecclesiam salutate Ephaenetum dilectum mihi qui est primitivus Asiae in Christo
ROM|16|6|salutate Mariam quae multum laboravit in vobis
ROM|16|7|salutate Andronicum et Iuniam cognatos et concaptivos meos qui sunt nobiles in apostolis qui et ante me fuerunt in Christo
ROM|16|8|salutate Ampliatum dilectissimum mihi in Domino
ROM|16|9|salutate Urbanum adiutorem nostrum in Christo et Stachyn dilectum meum
ROM|16|10|salutate Apellen probum in Christo
ROM|16|11|salutate eos qui sunt ex Aristoboli salutate Herodionem cognatum meum salutate eos qui sunt ex Narcissi qui sunt in Domino
ROM|16|12|salutate Tryfenam et Tryfosam quae laborant in Domino salutate Persidam carissimam quae multum laboravit in Domino
ROM|16|13|salutate Rufum electum in Domino et matrem eius et meam
ROM|16|14|salutate Asyncritum Flegonta Hermen Patrobam Hermam et qui cum eis sunt fratres
ROM|16|15|salutate Filologum et Iuliam Nereum et sororem eius et Olympiadem et omnes qui cum eis sunt sanctos
ROM|16|16|salutate invicem in osculo sancto salutant vos omnes ecclesiae Christi
ROM|16|17|rogo autem vos fratres ut observetis eos qui dissensiones et offendicula praeter doctrinam quam vos didicistis faciunt et declinate ab illis
ROM|16|18|huiusmodi enim Christo Domino nostro non serviunt sed suo ventri et per dulces sermones et benedictiones seducunt corda innocentium
ROM|16|19|vestra enim oboedientia in omnem locum divulgata est gaudeo igitur in vobis sed volo vos sapientes esse in bono et simplices in malo
ROM|16|20|Deus autem pacis conteret Satanan sub pedibus vestris velociter gratia Domini nostri Iesu Christi vobiscum
ROM|16|21|salutat vos Timotheus adiutor meus et Lucius et Iason et Sosipater cognati mei
ROM|16|22|saluto vos ego Tertius qui scripsi epistulam in Domino
ROM|16|23|salutat vos Gaius hospes meus et universae ecclesiae salutat vos Erastus arcarius civitatis et Quartus frater
ROM|16|24|
ROM|16|25|ei autem qui potens est vos confirmare iuxta evangelium meum et praedicationem Iesu Christi secundum revelationem mysterii temporibus aeternis taciti
ROM|16|26|quod nunc patefactum est per scripturas prophetarum secundum praeceptum aeterni Dei ad oboeditionem fidei in cunctis gentibus cognito
ROM|16|27|solo sapienti Deo per Iesum Christum cui honor in saecula saeculorum amen
1COR|1|1|Paulus vocatus apostolus Christi Iesu per voluntatem Dei et Sosthenes frater
1COR|1|2|ecclesiae Dei quae est Corinthi sanctificatis in Christo Iesu vocatis sanctis cum omnibus qui invocant nomen Domini nostri Iesu Christi in omni loco ipsorum et nostro
1COR|1|3|gratia vobis et pax a Deo Patre nostro et Domino Iesu Christo
1COR|1|4|gratias ago Deo meo semper pro vobis in gratia Dei quae data est vobis in Christo Iesu
1COR|1|5|quia in omnibus divites facti estis in illo in omni verbo et in omni scientia
1COR|1|6|sicut testimonium Christi confirmatum est in vobis
1COR|1|7|ita ut nihil vobis desit in ulla gratia expectantibus revelationem Domini nostri Iesu Christi
1COR|1|8|qui et confirmabit vos usque ad finem sine crimine in die adventus Domini nostri Iesu Christi
1COR|1|9|fidelis Deus per quem vocati estis in societatem Filii eius Iesu Christi Domini nostri
1COR|1|10|obsecro autem vos fratres per nomen Domini nostri Iesu Christi ut id ipsum dicatis omnes et non sint in vobis scismata sitis autem perfecti in eodem sensu et in eadem sententia
1COR|1|11|significatum est enim mihi de vobis fratres mei ab his qui sunt Chloes quia contentiones inter vos sunt
1COR|1|12|hoc autem dico quod unusquisque vestrum dicit ego quidem sum Pauli ego autem Apollo ego vero Cephae ego autem Christi
1COR|1|13|divisus est Christus numquid Paulus crucifixus est pro vobis aut in nomine Pauli baptizati estis
1COR|1|14|gratias ago Deo quod neminem vestrum baptizavi nisi Crispum et Gaium
1COR|1|15|ne quis dicat quod in nomine meo baptizati sitis
1COR|1|16|baptizavi autem et Stephanae domum ceterum nescio si quem alium baptizaverim
1COR|1|17|non enim misit me Christus baptizare sed evangelizare non in sapientia verbi ut non evacuetur crux Christi
1COR|1|18|verbum enim crucis pereuntibus quidem stultitia est his autem qui salvi fiunt id est nobis virtus Dei est
1COR|1|19|scriptum est enim perdam sapientiam sapientium et prudentiam prudentium reprobabo
1COR|1|20|ubi sapiens ubi scriba ubi conquisitor huius saeculi nonne stultam fecit Deus sapientiam huius mundi
1COR|1|21|nam quia in Dei sapientia non cognovit mundus per sapientiam Deum placuit Deo per stultitiam praedicationis salvos facere credentes
1COR|1|22|quoniam et Iudaei signa petunt et Graeci sapientiam quaerunt
1COR|1|23|nos autem praedicamus Christum crucifixum Iudaeis quidem scandalum gentibus autem stultitiam
1COR|1|24|ipsis autem vocatis Iudaeis atque Graecis Christum Dei virtutem et Dei sapientiam
1COR|1|25|quia quod stultum est Dei sapientius est hominibus et quod infirmum est Dei fortius est hominibus
1COR|1|26|videte enim vocationem vestram fratres quia non multi sapientes secundum carnem non multi potentes non multi nobiles
1COR|1|27|sed quae stulta sunt mundi elegit Deus ut confundat sapientes et infirma mundi elegit Deus ut confundat fortia
1COR|1|28|et ignobilia mundi et contemptibilia elegit Deus et quae non sunt ut ea quae sunt destrueret
1COR|1|29|ut non glorietur omnis caro in conspectu eius
1COR|1|30|ex ipso autem vos estis in Christo Iesu qui factus est sapientia nobis a Deo et iustitia et sanctificatio et redemptio
1COR|1|31|ut quemadmodum scriptum est qui gloriatur in Domino glorietur
1COR|2|1|et ego cum venissem ad vos fratres veni non per sublimitatem sermonis aut sapientiae adnuntians vobis testimonium Christi
1COR|2|2|non enim iudicavi scire me aliquid inter vos nisi Iesum Christum et hunc crucifixum
1COR|2|3|et ego in infirmitate et timore et tremore multo fui apud vos
1COR|2|4|et sermo meus et praedicatio mea non in persuasibilibus sapientiae verbis sed in ostensione Spiritus et virtutis
1COR|2|5|ut fides vestra non sit in sapientia hominum sed in virtute Dei
1COR|2|6|sapientiam autem loquimur inter perfectos sapientiam vero non huius saeculi neque principum huius saeculi qui destruuntur
1COR|2|7|sed loquimur Dei sapientiam in mysterio quae abscondita est quam praedestinavit Deus ante saecula in gloriam nostram
1COR|2|8|quam nemo principum huius saeculi cognovit si enim cognovissent numquam Dominum gloriae crucifixissent
1COR|2|9|sed sicut scriptum est quod oculus non vidit nec auris audivit nec in cor hominis ascendit quae praeparavit Deus his qui diligunt illum
1COR|2|10|nobis autem revelavit Deus per Spiritum suum Spiritus enim omnia scrutatur etiam profunda Dei
1COR|2|11|quis enim scit hominum quae sint hominis nisi spiritus hominis qui in ipso est ita et quae Dei sunt nemo cognovit nisi Spiritus Dei
1COR|2|12|nos autem non spiritum mundi accepimus sed Spiritum qui ex Deo est ut sciamus quae a Deo donata sunt nobis
1COR|2|13|quae et loquimur non in doctis humanae sapientiae verbis sed in doctrina Spiritus spiritalibus spiritalia conparantes
1COR|2|14|animalis autem homo non percipit ea quae sunt Spiritus Dei stultitia est enim illi et non potest intellegere quia spiritaliter examinatur
1COR|2|15|spiritalis autem iudicat omnia et ipse a nemine iudicatur
1COR|2|16|quis enim cognovit sensum Domini qui instruat eum nos autem sensum Christi habemus
1COR|3|1|et ego fratres non potui vobis loqui quasi spiritalibus sed quasi carnalibus tamquam parvulis in Christo
1COR|3|2|lac vobis potum dedi non escam nondum enim poteratis sed ne nunc quidem potestis adhuc enim estis carnales
1COR|3|3|cum enim sit inter vos zelus et contentio nonne carnales estis et secundum hominem ambulatis
1COR|3|4|cum enim quis dicit ego quidem sum Pauli alius autem ego Apollo nonne homines estis quid igitur est Apollo quid vero Paulus
1COR|3|5|ministri eius cui credidistis et unicuique sicut Dominus dedit
1COR|3|6|ego plantavi Apollo rigavit sed Deus incrementum dedit
1COR|3|7|itaque neque qui plantat est aliquid neque qui rigat sed qui incrementum dat Deus
1COR|3|8|qui plantat autem et qui rigat unum sunt unusquisque autem propriam mercedem accipiet secundum suum laborem
1COR|3|9|Dei enim sumus adiutores Dei agricultura estis Dei aedificatio estis
1COR|3|10|secundum gratiam Dei quae data est mihi ut sapiens architectus fundamentum posui alius autem superaedificat unusquisque autem videat quomodo superaedificet
1COR|3|11|fundamentum enim aliud nemo potest ponere praeter id quod positum est qui est Christus Iesus
1COR|3|12|si quis autem superaedificat supra fundamentum hoc aurum argentum lapides pretiosos ligna faenum stipulam
1COR|3|13|uniuscuiusque opus manifestum erit dies enim declarabit quia in igne revelabitur et uniuscuiusque opus quale sit ignis probabit
1COR|3|14|si cuius opus manserit quod superaedificavit mercedem accipiet
1COR|3|15|si cuius opus arserit detrimentum patietur ipse autem salvus erit sic tamen quasi per ignem
1COR|3|16|nescitis quia templum Dei estis et Spiritus Dei habitat in vobis
1COR|3|17|si quis autem templum Dei violaverit disperdet illum Deus templum enim Dei sanctum est quod estis vos
1COR|3|18|nemo se seducat si quis videtur inter vos sapiens esse in hoc saeculo stultus fiat ut sit sapiens
1COR|3|19|sapientia enim huius mundi stultitia est apud Deum scriptum est enim conprehendam sapientes in astutia eorum
1COR|3|20|et iterum Dominus novit cogitationes sapientium quoniam vanae sunt
1COR|3|21|itaque nemo glorietur in hominibus omnia enim vestra sunt
1COR|3|22|sive Paulus sive Apollo sive Cephas sive mundus sive vita sive mors sive praesentia sive futura omnia enim vestra sunt
1COR|3|23|vos autem Christi Christus autem Dei
1COR|4|1|sic nos existimet homo ut ministros Christi et dispensatores mysteriorum Dei
1COR|4|2|hic iam quaeritur inter dispensatores ut fidelis quis inveniatur
1COR|4|3|mihi autem pro minimo est ut a vobis iudicer aut ab humano die sed neque me ipsum iudico
1COR|4|4|nihil enim mihi conscius sum sed non in hoc iustificatus sum qui autem iudicat me Dominus est
1COR|4|5|itaque nolite ante tempus iudicare quoadusque veniat Dominus qui et inluminabit abscondita tenebrarum et manifestabit consilia cordium et tunc laus erit unicuique a Deo
1COR|4|6|haec autem fratres transfiguravi in me et Apollo propter vos ut in nobis discatis ne supra quam scriptum est unus adversus alterum infletur pro alio
1COR|4|7|quis enim te discernit quid autem habes quod non accepisti si autem accepisti quid gloriaris quasi non acceperis
1COR|4|8|iam saturati estis iam divites facti estis sine nobis regnastis et utinam regnaretis ut et nos vobiscum regnaremus
1COR|4|9|puto enim Deus nos apostolos novissimos ostendit tamquam morti destinatos quia spectaculum facti sumus mundo et angelis et hominibus
1COR|4|10|nos stulti propter Christum vos autem prudentes in Christo nos infirmi vos autem fortes vos nobiles nos autem ignobiles
1COR|4|11|usque in hanc horam et esurimus et sitimus et nudi sumus et colaphis caedimur et instabiles sumus
1COR|4|12|et laboramus operantes manibus nostris maledicimur et benedicimus persecutionem patimur et sustinemus
1COR|4|13|blasphemamur et obsecramus tamquam purgamenta huius mundi facti sumus omnium peripsima usque adhuc
1COR|4|14|non ut confundam vos haec scribo sed ut filios meos carissimos moneo
1COR|4|15|nam si decem milia pedagogorum habeatis in Christo sed non multos patres nam in Christo Iesu per evangelium ego vos genui
1COR|4|16|rogo ergo vos imitatores mei estote
1COR|4|17|ideo misi ad vos Timotheum qui est filius meus carissimus et fidelis in Domino qui vos commonefaciat vias meas quae sunt in Christo sicut ubique in omni ecclesia doceo
1COR|4|18|tamquam non venturus sim ad vos sic inflati sunt quidam
1COR|4|19|veniam autem cito ad vos si Dominus voluerit et cognoscam non sermonem eorum qui inflati sunt sed virtutem
1COR|4|20|non enim in sermone est regnum Dei sed in virtute
1COR|4|21|quid vultis in virga veniam ad vos an in caritate et spiritu mansuetudinis
1COR|5|1|omnino auditur inter vos fornicatio et talis fornicatio qualis nec inter gentes ita ut uxorem patris aliquis habeat
1COR|5|2|et vos inflati estis et non magis luctum habuistis ut tollatur de medio vestrum qui hoc opus fecit
1COR|5|3|ego quidem absens corpore praesens autem spiritu iam iudicavi ut praesens eum qui sic operatus est
1COR|5|4|in nomine Domini nostri Iesu Christi congregatis vobis et meo spiritu cum virtute Domini Iesu
1COR|5|5|tradere huiusmodi Satanae in interitum carnis ut spiritus salvus sit in die Domini Iesu
1COR|5|6|non bona gloriatio vestra nescitis quia modicum fermentum totam massam corrumpit
1COR|5|7|expurgate vetus fermentum ut sitis nova consparsio sicut estis azymi etenim pascha nostrum immolatus est Christus
1COR|5|8|itaque epulemur non in fermento veteri neque in fermento malitiae et nequitiae sed in azymis sinceritatis et veritatis
1COR|5|9|scripsi vobis in epistula ne commisceamini fornicariis
1COR|5|10|non utique fornicariis huius mundi aut avaris aut rapacibus aut idolis servientibus alioquin debueratis de hoc mundo exisse
1COR|5|11|nunc autem scripsi vobis non commisceri si is qui frater nominatur est fornicator aut avarus aut idolis serviens aut maledicus aut ebriosus aut rapax cum eiusmodi nec cibum sumere
1COR|5|12|quid enim mihi de his qui foris sunt iudicare nonne de his qui intus sunt vos iudicatis
1COR|5|13|nam eos qui foris sunt Deus iudicabit auferte malum ex vobis ipsis
1COR|6|1|audet aliquis vestrum habens negotium adversus alterum iudicari apud iniquos et non apud sanctos
1COR|6|2|an nescitis quoniam sancti de mundo iudicabunt et si in vobis iudicabitur mundus indigni estis qui de minimis iudicetis
1COR|6|3|nescitis quoniam angelos iudicabimus quanto magis saecularia
1COR|6|4|saecularia igitur iudicia si habueritis contemptibiles qui sunt in ecclesia illos constituite ad iudicandum
1COR|6|5|ad verecundiam vestram dico sic non est inter vos sapiens quisquam qui possit iudicare inter fratrem suum
1COR|6|6|sed frater cum fratre iudicio contendit et hoc apud infideles
1COR|6|7|iam quidem omnino delictum est in vobis quod iudicia habetis inter vos quare non magis iniuriam accipitis quare non magis fraudem patimini
1COR|6|8|sed vos iniuriam facitis et fraudatis et hoc fratribus
1COR|6|9|an nescitis quia iniqui regnum Dei non possidebunt nolite errare neque fornicarii neque idolis servientes neque adulteri
1COR|6|10|neque molles neque masculorum concubitores neque fures neque avari neque ebriosi neque maledici neque rapaces regnum Dei possidebunt
1COR|6|11|et haec quidam fuistis sed abluti estis sed sanctificati estis sed iustificati estis in nomine Domini nostri Iesu Christi et in Spiritu Dei nostri
1COR|6|12|omnia mihi licent sed non omnia expediunt omnia mihi licent sed ego sub nullius redigar potestate
1COR|6|13|esca ventri et venter escis Deus autem et hunc et haec destruet corpus autem non fornicationi sed Domino et Dominus corpori
1COR|6|14|Deus vero et Dominum suscitavit et nos suscitabit per virtutem suam
1COR|6|15|nescitis quoniam corpora vestra membra Christi sunt tollens ergo membra Christi faciam membra meretricis absit
1COR|6|16|an nescitis quoniam qui adheret meretrici unum corpus efficitur erunt enim inquit duo in carne una
1COR|6|17|qui autem adheret Domino unus spiritus est
1COR|6|18|fugite fornicationem omne peccatum quodcumque fecerit homo extra corpus est qui autem fornicatur in corpus suum peccat
1COR|6|19|an nescitis quoniam membra vestra templum est Spiritus Sancti qui in vobis est quem habetis a Deo et non estis vestri
1COR|6|20|empti enim estis pretio magno glorificate et portate Deum in corpore vestro
1COR|7|1|de quibus autem scripsistis bonum est homini mulierem non tangere
1COR|7|2|propter fornicationes autem unusquisque suam uxorem habeat et unaquaeque suum virum habeat
1COR|7|3|uxori vir debitum reddat similiter autem et uxor viro
1COR|7|4|mulier sui corporis potestatem non habet sed vir similiter autem et vir sui corporis potestatem non habet sed mulier
1COR|7|5|nolite fraudare invicem nisi forte ex consensu ad tempus ut vacetis orationi et iterum revertimini in id ipsum ne temptet vos Satanas propter incontinentiam vestram
1COR|7|6|hoc autem dico secundum indulgentiam non secundum imperium
1COR|7|7|volo autem omnes homines esse sicut me ipsum sed unusquisque proprium habet donum ex Deo alius quidem sic alius vero sic
1COR|7|8|dico autem non nuptis et viduis bonum est illis si sic maneant sicut et ego
1COR|7|9|quod si non se continent nubant melius est enim nubere quam uri
1COR|7|10|his autem qui matrimonio iuncti sunt praecipio non ego sed Dominus uxorem a viro non discedere
1COR|7|11|quod si discesserit manere innuptam aut viro suo reconciliari et vir uxorem ne dimittat
1COR|7|12|nam ceteris ego dico non Dominus si quis frater uxorem habet infidelem et haec consentit habitare cum illo non dimittat illam
1COR|7|13|et si qua mulier habet virum infidelem et hic consentit habitare cum illa non dimittat virum
1COR|7|14|sanctificatus est enim vir infidelis in muliere fideli et sanctificata est mulier infidelis per virum fidelem alioquin filii vestri inmundi essent nunc autem sancti sunt
1COR|7|15|quod si infidelis discedit discedat non est enim servituti subiectus frater aut soror in eiusmodi in pace autem vocavit nos Deus
1COR|7|16|unde enim scis mulier si virum salvum facies aut unde scis vir si mulierem salvam facies
1COR|7|17|nisi unicuique sicut divisit Dominus unumquemque sicut vocavit Deus ita ambulet et sic in omnibus ecclesiis doceo
1COR|7|18|circumcisus aliquis vocatus est non adducat praeputium in praeputio aliquis vocatus est non circumcidatur
1COR|7|19|circumcisio nihil est et praeputium nihil est sed observatio mandatorum Dei
1COR|7|20|unusquisque in qua vocatione vocatus est in ea permaneat
1COR|7|21|servus vocatus es non sit tibi curae sed et si potes liber fieri magis utere
1COR|7|22|qui enim in Domino vocatus est servus libertus est Domini similiter qui liber vocatus est servus est Christi
1COR|7|23|pretio empti estis nolite fieri servi hominum
1COR|7|24|unusquisque in quo vocatus est fratres in hoc maneat apud Deum
1COR|7|25|de virginibus autem praeceptum Domini non habeo consilium autem do tamquam misericordiam consecutus a Domino ut sim fidelis
1COR|7|26|existimo ergo hoc bonum esse propter instantem necessitatem quoniam bonum est homini sic esse
1COR|7|27|alligatus es uxori noli quaerere solutionem solutus es ab uxore noli quaerere uxorem
1COR|7|28|si autem acceperis uxorem non peccasti et si nupserit virgo non peccavit tribulationem tamen carnis habebunt huiusmodi ego autem vobis parco
1COR|7|29|hoc itaque dico fratres tempus breve est reliquum est ut qui habent uxores tamquam non habentes sint
1COR|7|30|et qui flent tamquam non flentes et qui gaudent tamquam non gaudentes et qui emunt tamquam non possidentes
1COR|7|31|et qui utuntur hoc mundo tamquam non utantur praeterit enim figura huius mundi
1COR|7|32|volo autem vos sine sollicitudine esse qui sine uxore est sollicitus est quae Domini sunt quomodo placeat Deo
1COR|7|33|qui autem cum uxore est sollicitus est quae sunt mundi quomodo placeat uxori et divisus est
1COR|7|34|et mulier innupta et virgo cogitat quae Domini sunt ut sit sancta et corpore et spiritu quae autem nupta est cogitat quae sunt mundi quomodo placeat viro
1COR|7|35|porro hoc ad utilitatem vestram dico non ut laqueum vobis iniciam sed ad id quod honestum est et quod facultatem praebeat sine inpedimento Dominum observandi
1COR|7|36|si quis autem turpem se videri existimat super virgine sua quod sit superadulta et ita oportet fieri quod vult faciat non peccat nubat
1COR|7|37|nam qui statuit in corde suo firmus non habens necessitatem potestatem autem habet suae voluntatis et hoc iudicavit in corde suo servare virginem suam bene facit
1COR|7|38|igitur et qui matrimonio iungit virginem suam bene facit et qui non iungit melius facit
1COR|7|39|mulier alligata est quanto tempore vir eius vivit quod si dormierit vir eius liberata est cui vult nubat tantum in Domino
1COR|7|40|beatior autem erit si sic permanserit secundum meum consilium puto autem quod et ego Spiritum Dei habeo
1COR|8|1|de his autem quae idolis sacrificantur scimus quia omnes scientiam habemus scientia inflat caritas vero aedificat
1COR|8|2|si quis se existimat scire aliquid nondum cognovit quemadmodum oporteat eum scire
1COR|8|3|si quis autem diligit Deum hic cognitus est ab eo
1COR|8|4|de escis autem quae idolis immolantur scimus quia nihil est idolum in mundo et quod nullus Deus nisi unus
1COR|8|5|nam et si sunt qui dicantur dii sive in caelo sive in terra siquidem sunt dii multi et domini multi
1COR|8|6|nobis tamen unus Deus Pater ex quo omnia et nos in illum et unus Dominus Iesus Christus per quem omnia et nos per ipsum
1COR|8|7|sed non in omnibus est scientia quidam autem conscientia usque nunc idoli quasi idolothytum manducant et conscientia ipsorum cum sit infirma polluitur
1COR|8|8|esca autem nos non commendat Deo neque si non manducaverimus deficiemus neque si manducaverimus abundabimus
1COR|8|9|videte autem ne forte haec licentia vestra offendiculum fiat infirmibus
1COR|8|10|si enim quis viderit eum qui habet scientiam in idolio recumbentem nonne conscientia eius cum sit infirma aedificabitur ad manducandum idolothyta
1COR|8|11|et peribit infirmus in tua scientia frater propter quem Christus mortuus est
1COR|8|12|sic autem peccantes in fratres et percutientes conscientiam eorum infirmam in Christo peccatis
1COR|8|13|quapropter si esca scandalizat fratrem meum non manducabo carnem in aeternum ne fratrem meum scandalizem
1COR|9|1|non sum liber non sum apostolus nonne Iesum Dominum nostrum vidi non opus meum vos estis in Domino
1COR|9|2|si aliis non sum apostolus sed tamen vobis sum nam signaculum apostolatus mei vos estis in Domino
1COR|9|3|mea defensio apud eos qui me interrogant haec est
1COR|9|4|numquid non habemus potestatem manducandi et bibendi
1COR|9|5|numquid non habemus potestatem sororem mulierem circumducendi sicut et ceteri apostoli et fratres Domini et Cephas
1COR|9|6|aut solus ego et Barnabas non habemus potestatem hoc operandi
1COR|9|7|quis militat suis stipendiis umquam quis plantat vineam et fructum eius non edit quis pascit gregem et de lacte gregis non manducat
1COR|9|8|numquid secundum hominem haec dico an et lex haec non dicit
1COR|9|9|scriptum est enim in lege Mosi non alligabis os bovi trituranti numquid de bubus cura est Deo
1COR|9|10|an propter nos utique dicit nam propter nos scripta sunt quoniam debet in spe qui arat arare et qui triturat in spe fructus percipiendi
1COR|9|11|si nos vobis spiritalia seminavimus magnum est si nos carnalia vestra metamus
1COR|9|12|si alii potestatis vestrae participes sunt non potius nos sed non usi sumus hac potestate sed omnia sustinemus ne quod offendiculum demus evangelio Christi
1COR|9|13|nescitis quoniam qui in sacrario operantur quae de sacrario sunt edunt qui altario deserviunt cum altario participantur
1COR|9|14|ita et Dominus ordinavit his qui evangelium adnuntiant de evangelio vivere
1COR|9|15|ego autem nullo horum usus sum non scripsi autem haec ut ita fiant in me bonum est enim mihi magis mori quam ut gloriam meam quis evacuet
1COR|9|16|nam si evangelizavero non est mihi gloria necessitas enim mihi incumbit vae enim mihi est si non evangelizavero
1COR|9|17|si enim volens hoc ago mercedem habeo si autem invitus dispensatio mihi credita est
1COR|9|18|quae est ergo merces mea ut evangelium praedicans sine sumptu ponam evangelium ut non abutar potestate mea in evangelio
1COR|9|19|nam cum liber essem ex omnibus omnium me servum feci ut plures lucri facerem
1COR|9|20|et factus sum Iudaeis tamquam Iudaeus ut Iudaeos lucrarer
1COR|9|21|his qui sub lege sunt quasi sub lege essem cum ipse non essem sub lege ut eos qui sub lege erant lucri facerem his qui sine lege erant tamquam sine lege essem cum sine lege Dei non essem sed in lege essem Christi ut lucri facerem eos qui sine lege erant
1COR|9|22|factus sum infirmis infirmus ut infirmos lucri facerem omnibus omnia factus sum ut omnes facerem salvos
1COR|9|23|omnia autem facio propter evangelium ut particeps eius efficiar
1COR|9|24|nescitis quod hii qui in stadio currunt omnes quidem currunt sed unus accipit bravium sic currite ut conprehendatis
1COR|9|25|omnis autem qui in agone contendit ab omnibus se abstinet et illi quidem ut corruptibilem coronam accipiant nos autem incorruptam
1COR|9|26|ego igitur sic curro non quasi in incertum sic pugno non quasi aerem verberans
1COR|9|27|sed castigo corpus meum et in servitutem redigo ne forte cum aliis praedicaverim ipse reprobus efficiar
1COR|10|1|nolo enim vos ignorare fratres quoniam patres nostri omnes sub nube fuerunt et omnes mare transierunt
1COR|10|2|et omnes in Mose baptizati sunt in nube et in mari
1COR|10|3|et omnes eandem escam spiritalem manducaverunt
1COR|10|4|et omnes eundem potum spiritalem biberunt bibebant autem de spiritali consequenti eos petra petra autem erat Christus
1COR|10|5|sed non in pluribus eorum beneplacitum est Deo nam prostrati sunt in deserto
1COR|10|6|haec autem in figura facta sunt nostri ut non simus concupiscentes malorum sicut et illi concupierunt
1COR|10|7|neque idolorum cultores efficiamini sicut quidam ex ipsis quemadmodum scriptum est sedit populus manducare et bibere et surrexerunt ludere
1COR|10|8|neque fornicemur sicut quidam ex ipsis fornicati sunt et ceciderunt una die viginti tria milia
1COR|10|9|neque temptemus Christum sicut quidam eorum temptaverunt et a serpentibus perierunt
1COR|10|10|neque murmuraveritis sicut quidam eorum murmuraverunt et perierunt ab exterminatore
1COR|10|11|haec autem omnia in figura contingebant illis scripta sunt autem ad correptionem nostram in quos fines saeculorum devenerunt
1COR|10|12|itaque qui se existimat stare videat ne cadat
1COR|10|13|temptatio vos non adprehendat nisi humana fidelis autem Deus qui non patietur vos temptari super id quod potestis sed faciet cum temptatione etiam proventum ut possitis sustinere
1COR|10|14|propter quod carissimi mihi fugite ab idolorum cultura
1COR|10|15|ut prudentibus loquor vos iudicate quod dico
1COR|10|16|calicem benedictionis cui benedicimus nonne communicatio sanguinis Christi est et panis quem frangimus nonne participatio corporis Domini est
1COR|10|17|quoniam unus panis unum corpus multi sumus omnes quidem de uno pane participamur
1COR|10|18|videte Israhel secundum carnem nonne qui edunt hostias participes sunt altaris
1COR|10|19|quid ergo dico quod idolis immolatum sit aliquid aut quod idolum sit aliquid
1COR|10|20|sed quae immolant gentes daemoniis immolant et non Deo nolo autem vos socios fieri daemoniorum non potestis calicem Domini bibere et calicem daemoniorum
1COR|10|21|non potestis mensae Domini participes esse et mensae daemoniorum
1COR|10|22|an aemulamur Dominum numquid fortiores illo sumus omnia licent sed non omnia expediunt
1COR|10|23|omnia licent sed non omnia aedificant
1COR|10|24|nemo quod suum est quaerat sed quod alterius
1COR|10|25|omne quod in macello venit manducate nihil interrogantes propter conscientiam
1COR|10|26|Domini est terra et plenitudo eius
1COR|10|27|si quis vocat vos infidelium et vultis ire omne quod vobis adponitur manducate nihil interrogantes propter conscientiam
1COR|10|28|si quis autem dixerit hoc immolaticium est idolis nolite manducare propter illum qui indicavit et propter conscientiam
1COR|10|29|conscientiam autem dico non tuam sed alterius ut quid enim libertas mea iudicatur ab alia conscientia
1COR|10|30|si ego cum gratia participo quid blasphemor pro eo quod gratias ago
1COR|10|31|sive ergo manducatis sive bibitis vel aliud quid facitis omnia in gloriam Dei facite
1COR|10|32|sine offensione estote Iudaeis et gentilibus et ecclesiae Dei
1COR|10|33|sicut et ego per omnia omnibus placeo non quaerens quod mihi utile est sed quod multis ut salvi fiant
1COR|11|1|imitatores mei estote sicut et ego Christi
1COR|11|2|laudo autem vos fratres quod omnia mei memores estis et sicut tradidi vobis praecepta mea tenetis
1COR|11|3|volo autem vos scire quod omnis viri caput Christus est caput autem mulieris vir caput vero Christi Deus
1COR|11|4|omnis vir orans aut prophetans velato capite deturpat caput suum
1COR|11|5|omnis autem mulier orans aut prophetans non velato capite deturpat caput suum unum est enim atque si decalvetur
1COR|11|6|nam si non velatur mulier et tondeatur si vero turpe est mulieri tonderi aut decalvari velet caput suum
1COR|11|7|vir quidem non debet velare caput quoniam imago et gloria est Dei mulier autem gloria viri est
1COR|11|8|non enim vir ex muliere est sed mulier ex viro
1COR|11|9|etenim non est creatus vir propter mulierem sed mulier propter virum
1COR|11|10|ideo debet mulier potestatem habere supra caput propter angelos
1COR|11|11|verumtamen neque vir sine muliere neque mulier sine viro in Domino
1COR|11|12|nam sicut mulier de viro ita et vir per mulierem omnia autem ex Deo
1COR|11|13|vos ipsi iudicate decet mulierem non velatam orare Deum
1COR|11|14|nec ipsa natura docet vos quod vir quidem si comam nutriat ignominia est illi
1COR|11|15|mulier vero si comam nutriat gloria est illi quoniam capilli pro velamine ei dati sunt
1COR|11|16|si quis autem videtur contentiosus esse nos talem consuetudinem non habemus neque ecclesiae Dei
1COR|11|17|hoc autem praecipio non laudans quod non in melius sed in deterius convenitis
1COR|11|18|primum quidem convenientibus vobis in ecclesia audio scissuras esse et ex parte credo
1COR|11|19|nam oportet et hereses esse ut et qui probati sunt manifesti fiant in vobis
1COR|11|20|convenientibus ergo vobis in unum iam non est dominicam cenam manducare
1COR|11|21|unusquisque enim suam cenam praesumit ad manducandum et alius quidem esurit alius autem ebrius est
1COR|11|22|numquid domos non habetis ad manducandum et bibendum aut ecclesiam Dei contemnitis et confunditis eos qui non habent quid dicam vobis laudo vos in hoc non laudo
1COR|11|23|ego enim accepi a Domino quod et tradidi vobis quoniam Dominus Iesus in qua nocte tradebatur accepit panem
1COR|11|24|et gratias agens fregit et dixit hoc est corpus meum pro vobis hoc facite in meam commemorationem
1COR|11|25|similiter et calicem postquam cenavit dicens hic calix novum testamentum est in meo sanguine hoc facite quotienscumque bibetis in meam commemorationem
1COR|11|26|quotienscumque enim manducabitis panem hunc et calicem bibetis mortem Domini adnuntiatis donec veniat
1COR|11|27|itaque quicumque manducaverit panem vel biberit calicem Domini indigne reus erit corporis et sanguinis Domini
1COR|11|28|probet autem se ipsum homo et sic de pane illo edat et de calice bibat
1COR|11|29|qui enim manducat et bibit indigne iudicium sibi manducat et bibit non diiudicans corpus
1COR|11|30|ideo inter vos multi infirmes et inbecilles et dormiunt multi
1COR|11|31|quod si nosmet ipsos diiudicaremus non utique iudicaremur
1COR|11|32|dum iudicamur autem a Domino corripimur ut non cum hoc mundo damnemur
1COR|11|33|itaque fratres mei cum convenitis ad manducandum invicem expectate
1COR|11|34|si quis esurit domi manducet ut non in iudicium conveniatis cetera autem cum venero disponam
1COR|12|1|de spiritalibus autem nolo vos ignorare fratres
1COR|12|2|scitis quoniam cum gentes essetis ad simulacra muta prout ducebamini euntes
1COR|12|3|ideo notum vobis facio quod nemo in Spiritu Dei loquens dicit anathema Iesu et nemo potest dicere Dominus Iesus nisi in Spiritu Sancto
1COR|12|4|divisiones vero gratiarum sunt idem autem Spiritus
1COR|12|5|et divisiones ministrationum sunt idem autem Dominus
1COR|12|6|et divisiones operationum sunt idem vero Deus qui operatur omnia in omnibus
1COR|12|7|unicuique autem datur manifestatio Spiritus ad utilitatem
1COR|12|8|alii quidem per Spiritum datur sermo sapientiae alii autem sermo scientiae secundum eundem Spiritum
1COR|12|9|alteri fides in eodem Spiritu alii gratia sanitatum in uno Spiritu
1COR|12|10|alii operatio virtutum alii prophetatio alii discretio spirituum alii genera linguarum alii interpretatio sermonum
1COR|12|11|haec autem omnia operatur unus atque idem Spiritus dividens singulis prout vult
1COR|12|12|sicut enim corpus unum est et membra habet multa omnia autem membra corporis cum sint multa unum corpus sunt ita et Christus
1COR|12|13|etenim in uno Spiritu omnes nos in unum corpus baptizati sumus sive Iudaei sive gentiles sive servi sive liberi et omnes unum Spiritum potati sumus
1COR|12|14|nam et corpus non est unum membrum sed multa
1COR|12|15|si dixerit pes quoniam non sum manus non sum de corpore non ideo non est de corpore
1COR|12|16|et si dixerit auris quia non sum oculus non sum de corpore non ideo non est de corpore
1COR|12|17|si totum corpus oculus ubi auditus si totum auditus ubi odoratus
1COR|12|18|nunc autem posuit Deus membra unumquodque eorum in corpore sicut voluit
1COR|12|19|quod si essent omnia unum membrum ubi corpus
1COR|12|20|nunc autem multa quidem membra unum autem corpus
1COR|12|21|non potest dicere oculus manui opera tua non indigeo aut iterum caput pedibus non estis mihi necessarii
1COR|12|22|sed multo magis quae videntur membra corporis infirmiora esse necessariora sunt
1COR|12|23|et quae putamus ignobiliora membra esse corporis his honorem abundantiorem circumdamus et quae inhonesta sunt nostra abundantiorem honestatem habent
1COR|12|24|honesta autem nostra nullius egent sed Deus temperavit corpus ei cui deerat abundantiorem tribuendo honorem
1COR|12|25|ut non sit scisma in corpore sed id ipsum pro invicem sollicita sint membra
1COR|12|26|et si quid patitur unum membrum conpatiuntur omnia membra sive gloriatur unum membrum congaudent omnia membra
1COR|12|27|vos autem estis corpus Christi et membra de membro
1COR|12|28|et quosdam quidem posuit Deus in ecclesia primum apostolos secundo prophetas tertio doctores deinde virtutes exin gratias curationum opitulationes gubernationes genera linguarum
1COR|12|29|numquid omnes apostoli numquid omnes prophetae numquid omnes doctores
1COR|12|30|numquid omnes virtutes numquid omnes gratiam habent curationum numquid omnes linguis loquuntur numquid omnes interpretantur
1COR|12|31|aemulamini autem charismata maiora et adhuc excellentiorem viam vobis demonstro
1COR|13|1|si linguis hominum loquar et angelorum caritatem autem non habeam factus sum velut aes sonans aut cymbalum tinniens
1COR|13|2|et si habuero prophetiam et noverim mysteria omnia et omnem scientiam et habuero omnem fidem ita ut montes transferam caritatem autem non habuero nihil sum
1COR|13|3|et si distribuero in cibos pauperum omnes facultates meas et si tradidero corpus meum ut ardeam caritatem autem non habuero nihil mihi prodest
1COR|13|4|caritas patiens est benigna est caritas non aemulatur non agit perperam non inflatur
1COR|13|5|non est ambitiosa non quaerit quae sua sunt non inritatur non cogitat malum
1COR|13|6|non gaudet super iniquitatem congaudet autem veritati
1COR|13|7|omnia suffert omnia credit omnia sperat omnia sustinet
1COR|13|8|caritas numquam excidit sive prophetiae evacuabuntur sive linguae cessabunt sive scientia destruetur
1COR|13|9|ex parte enim cognoscimus et ex parte prophetamus
1COR|13|10|cum autem venerit quod perfectum est evacuabitur quod ex parte est
1COR|13|11|cum essem parvulus loquebar ut parvulus sapiebam ut parvulus cogitabam ut parvulus quando factus sum vir evacuavi quae erant parvuli
1COR|13|12|videmus nunc per speculum in enigmate tunc autem facie ad faciem nunc cognosco ex parte tunc autem cognoscam sicut et cognitus sum
1COR|13|13|nunc autem manet fides spes caritas tria haec maior autem his est caritas
1COR|14|1|sectamini caritatem aemulamini spiritalia magis autem ut prophetetis
1COR|14|2|qui enim loquitur lingua non hominibus loquitur sed Deo nemo enim audit Spiritu autem loquitur mysteria
1COR|14|3|nam qui prophetat hominibus loquitur aedificationem et exhortationem et consolationes
1COR|14|4|qui loquitur lingua semet ipsum aedificat qui autem prophetat ecclesiam aedificat
1COR|14|5|volo autem omnes vos loqui linguis magis autem prophetare nam maior est qui prophetat quam qui loquitur linguis nisi si forte ut interpretetur ut ecclesia aedificationem accipiat
1COR|14|6|nunc autem fratres si venero ad vos linguis loquens quid vobis prodero nisi si vobis loquar aut in revelatione aut scientia aut prophetia aut in doctrina
1COR|14|7|tamen quae sine anima sunt vocem dantia sive tibia sive cithara nisi distinctionem sonituum dederint quomodo scietur quod canitur aut quod citharizatur
1COR|14|8|etenim si incertam vocem det tuba quis parabit se ad bellum
1COR|14|9|ita et vos per linguam nisi manifestum sermonem dederitis quomodo scietur id quod dicitur eritis enim in aera loquentes
1COR|14|10|tam multa ut puta genera linguarum sunt in mundo et nihil sine voce est
1COR|14|11|si ergo nesciero virtutem vocis ero ei cui loquor barbarus et qui loquitur mihi barbarus
1COR|14|12|sic et vos quoniam aemulatores estis spirituum ad aedificationem ecclesiae quaerite ut abundetis
1COR|14|13|et ideo qui loquitur lingua oret ut interpretetur
1COR|14|14|nam si orem lingua spiritus meus orat mens autem mea sine fructu est
1COR|14|15|quid ergo est orabo spiritu orabo et mente psallam spiritu psallam et mente
1COR|14|16|ceterum si benedixeris spiritu qui supplet locum idiotae quomodo dicet amen super tuam benedictionem quoniam quid dicas nescit
1COR|14|17|nam tu quidem bene gratias agis sed alter non aedificatur
1COR|14|18|gratias ago Deo quod omnium vestrum lingua loquor
1COR|14|19|sed in ecclesia volo quinque verba sensu meo loqui ut et alios instruam quam decem milia verborum in lingua
1COR|14|20|fratres nolite pueri effici sensibus sed malitia parvuli estote sensibus autem perfecti estote
1COR|14|21|in lege scriptum est quoniam in aliis linguis et labiis aliis loquar populo huic et nec sic exaudient me dicit Dominus
1COR|14|22|itaque linguae in signum sunt non fidelibus sed infidelibus prophetia autem non infidelibus sed fidelibus
1COR|14|23|si ergo conveniat universa ecclesia in unum et omnes linguis loquantur intrent autem idiotae aut infideles nonne dicent quod insanitis
1COR|14|24|si autem omnes prophetent intret autem quis infidelis vel idiota convincitur ab omnibus diiudicatur ab omnibus
1COR|14|25|occulta cordis eius manifesta fiunt et ita cadens in faciem adorabit Deum pronuntians quod vere Deus in vobis est
1COR|14|26|quid ergo est fratres cum convenitis unusquisque vestrum psalmum habet doctrinam habet apocalypsin habet linguam habet interpretationem habet omnia ad aedificationem fiant
1COR|14|27|sive lingua quis loquitur secundum duos aut ut multum tres et per partes et unus interpretetur
1COR|14|28|si autem non fuerit interpres taceat in ecclesia sibi autem loquatur et Deo
1COR|14|29|prophetae duo aut tres dicant et ceteri diiudicent
1COR|14|30|quod si alii revelatum fuerit sedenti prior taceat
1COR|14|31|potestis enim omnes per singulos prophetare ut omnes discant et omnes exhortentur
1COR|14|32|et spiritus prophetarum prophetis subiecti sunt
1COR|14|33|non enim est dissensionis Deus sed pacis sicut in omnibus ecclesiis sanctorum
1COR|14|34|mulieres in ecclesiis taceant non enim permittitur eis loqui sed subditas esse sicut et lex dicit
1COR|14|35|si quid autem volunt discere domi viros suos interrogent turpe est enim mulieri loqui in ecclesia
1COR|14|36|an a vobis verbum Dei processit aut in vos solos pervenit
1COR|14|37|si quis videtur propheta esse aut spiritalis cognoscat quae scribo vobis quia Domini sunt mandata
1COR|14|38|si quis autem ignorat ignorabitur
1COR|14|39|itaque fratres aemulamini prophetare et loqui linguis nolite prohibere
1COR|14|40|omnia autem honeste et secundum ordinem fiant
1COR|15|1|notum autem vobis facio fratres evangelium quod praedicavi vobis quod et accepistis in quo et statis
1COR|15|2|per quod et salvamini qua ratione praedicaverim vobis si tenetis nisi si frustra credidistis
1COR|15|3|tradidi enim vobis in primis quod et accepi quoniam Christus mortuus est pro peccatis nostris secundum scripturas
1COR|15|4|et quia sepultus est et quia resurrexit tertia die secundum scripturas
1COR|15|5|et quia visus est Cephae et post haec undecim
1COR|15|6|deinde visus est plus quam quingentis fratribus simul ex quibus multi manent usque adhuc quidam autem dormierunt
1COR|15|7|deinde visus est Iacobo deinde apostolis omnibus
1COR|15|8|novissime autem omnium tamquam abortivo visus est et mihi
1COR|15|9|ego enim sum minimus apostolorum qui non sum dignus vocari apostolus quoniam persecutus sum ecclesiam Dei
1COR|15|10|gratia autem Dei sum id quod sum et gratia eius in me vacua non fuit sed abundantius illis omnibus laboravi non ego autem sed gratia Dei mecum
1COR|15|11|sive enim ego sive illi sic praedicamus et sic credidistis
1COR|15|12|si autem Christus praedicatur quod resurrexit a mortuis quomodo quidam dicunt in vobis quoniam resurrectio mortuorum non est
1COR|15|13|si autem resurrectio mortuorum non est neque Christus resurrexit
1COR|15|14|si autem Christus non resurrexit inanis est ergo praedicatio nostra inanis est et fides vestra
1COR|15|15|invenimur autem et falsi testes Dei quoniam testimonium diximus adversus Deum quod suscitaverit Christum quem non suscitavit si mortui non resurgunt
1COR|15|16|nam si mortui non resurgunt neque Christus resurrexit
1COR|15|17|quod si Christus non resurrexit vana est fides vestra adhuc enim estis in peccatis vestris
1COR|15|18|ergo et qui dormierunt in Christo perierunt
1COR|15|19|si in hac vita tantum in Christo sperantes sumus miserabiliores sumus omnibus hominibus
1COR|15|20|nunc autem Christus resurrexit a mortuis primitiae dormientium
1COR|15|21|quoniam enim per hominem mors et per hominem resurrectio mortuorum
1COR|15|22|et sicut in Adam omnes moriuntur ita et in Christo omnes vivificabuntur
1COR|15|23|unusquisque autem in suo ordine primitiae Christus deinde hii qui sunt Christi in adventu eius
1COR|15|24|deinde finis cum tradiderit regnum Deo et Patri cum evacuaverit omnem principatum et potestatem et virtutem
1COR|15|25|oportet autem illum regnare donec ponat omnes inimicos sub pedibus eius
1COR|15|26|novissima autem inimica destruetur mors omnia enim subiecit sub pedibus eius cum autem dicat
1COR|15|27|omnia subiecta sunt sine dubio praeter eum qui subiecit ei omnia
1COR|15|28|cum autem subiecta fuerint illi omnia tunc ipse Filius subiectus erit illi qui sibi subiecit omnia ut sit Deus omnia in omnibus
1COR|15|29|alioquin quid facient qui baptizantur pro mortuis si omnino mortui non resurgunt ut quid et baptizantur pro illis
1COR|15|30|ut quid et nos periclitamur omni hora
1COR|15|31|cotidie morior per vestram gloriam fratres quam habeo in Christo Iesu Domino nostro
1COR|15|32|si secundum hominem ad bestias pugnavi Ephesi quid mihi prodest si mortui non resurgunt manducemus et bibamus cras enim moriemur
1COR|15|33|nolite seduci corrumpunt mores bonos conloquia mala
1COR|15|34|evigilate iuste et nolite peccare ignorantiam enim Dei quidam habent ad reverentiam vobis loquor
1COR|15|35|sed dicet aliquis quomodo resurgunt mortui quali autem corpore veniunt
1COR|15|36|insipiens tu quod seminas non vivificatur nisi prius moriatur
1COR|15|37|et quod seminas non corpus quod futurum est seminas sed nudum granum ut puta tritici aut alicuius ceterorum
1COR|15|38|Deus autem dat illi corpus sicut voluit et unicuique seminum proprium corpus
1COR|15|39|non omnis caro eadem caro sed alia hominum alia pecorum alia caro volucrum alia autem piscium
1COR|15|40|et corpora caelestia et corpora terrestria sed alia quidem caelestium gloria alia autem terrestrium
1COR|15|41|alia claritas solis alia claritas lunae et alia claritas stellarum stella enim ab stella differt in claritate
1COR|15|42|sic et resurrectio mortuorum seminatur in corruptione surgit in incorruptione
1COR|15|43|seminatur in ignobilitate surgit in gloria seminatur in infirmitate surgit in virtute
1COR|15|44|seminatur corpus animale surgit corpus spiritale si est corpus animale est et spiritale sic et scriptum est
1COR|15|45|factus est primus homo Adam in animam viventem novissimus Adam in spiritum vivificantem
1COR|15|46|sed non prius quod spiritale est sed quod animale est deinde quod spiritale
1COR|15|47|primus homo de terra terrenus secundus homo de caelo caelestis
1COR|15|48|qualis terrenus tales et terreni et qualis caelestis tales et caelestes
1COR|15|49|igitur sicut portavimus imaginem terreni portemus et imaginem caelestis
1COR|15|50|hoc autem dico fratres quoniam caro et sanguis regnum Dei possidere non possunt neque corruptio incorruptelam possidebit
1COR|15|51|ecce mysterium vobis dico omnes quidem resurgemus sed non omnes inmutabimur
1COR|15|52|in momento in ictu oculi in novissima tuba canet enim et mortui resurgent incorrupti et nos inmutabimur
1COR|15|53|oportet enim corruptibile hoc induere incorruptelam et mortale hoc induere inmortalitatem
1COR|15|54|cum autem mortale hoc induerit inmortalitatem tunc fiet sermo qui scriptus est absorta est mors in victoria
1COR|15|55|ubi est mors victoria tua ubi est mors stimulus tuus
1COR|15|56|stimulus autem mortis peccatum est virtus vero peccati lex
1COR|15|57|Deo autem gratias qui dedit nobis victoriam per Dominum nostrum Iesum Christum
1COR|15|58|itaque fratres mei dilecti stabiles estote et inmobiles abundantes in opere Domini semper scientes quod labor vester non est inanis in Domino
1COR|16|1|de collectis autem quae fiunt in sanctos sicut ordinavi ecclesiis Galatiae ita et vos facite
1COR|16|2|per unam sabbati unusquisque vestrum apud se ponat recondens quod ei beneplacuerit ut non cum venero tunc collectae fiant
1COR|16|3|cum autem praesens fuero quos probaveritis per epistulas hos mittam perferre gratiam vestram in Hierusalem
1COR|16|4|quod si dignum fuerit ut et ego eam mecum ibunt
1COR|16|5|veniam autem ad vos cum Macedoniam pertransiero nam Macedoniam pertransibo
1COR|16|6|apud vos autem forsitan manebo vel etiam hiemabo ut vos me deducatis quocumque iero
1COR|16|7|nolo enim vos modo in transitu videre spero enim me aliquantum temporis manere apud vos si Dominus permiserit
1COR|16|8|permanebo autem Ephesi usque ad pentecosten
1COR|16|9|ostium enim mihi apertum est magnum et evidens et adversarii multi
1COR|16|10|si autem venerit Timotheus videte ut sine timore sit apud vos opus enim Domini operatur sicut et ego
1COR|16|11|ne quis ergo illum spernat deducite autem illum in pace ut veniat ad me expecto enim illum cum fratribus
1COR|16|12|de Apollo autem fratre multum rogavi eum ut veniret ad vos cum fratribus et utique non fuit voluntas ut nunc veniret veniet autem cum ei vacuum fuerit
1COR|16|13|vigilate state in fide viriliter agite et confortamini
1COR|16|14|omnia vestra in caritate fiant
1COR|16|15|obsecro autem vos fratres nostis domum Stephanae et Fortunati quoniam sunt primitiae Achaiae et in ministerium sanctorum ordinaverunt se ipsos
1COR|16|16|ut et vos subditi sitis eiusmodi et omni cooperanti et laboranti
1COR|16|17|gaudeo autem in praesentia Stephanae et Fortunati et Achaici quoniam id quod vobis deerat ipsi suppleverunt
1COR|16|18|refecerunt enim et meum spiritum et vestrum cognoscite ergo qui eiusmodi sunt
1COR|16|19|salutant vos ecclesiae Asiae salutant vos in Domino multum Aquila et Prisca cum domestica sua ecclesia
1COR|16|20|salutant vos fratres omnes salutate invicem in osculo sancto
1COR|16|21|salutatio mea manu Pauli
1COR|16|22|si quis non amat Dominum Iesum Christum sit anathema maranatha
1COR|16|23|gratia Domini Iesu vobiscum
1COR|16|24|caritas mea cum omnibus vobis in Christo Iesu amen
2COR|1|1|Paulus apostolus Iesu Christi per voluntatem Dei et Timotheus frater ecclesiae Dei quae est Corinthi cum sanctis omnibus qui sunt in universa Achaia
2COR|1|2|gratia vobis et pax a Deo Patre nostro et Domino Iesu Christo
2COR|1|3|benedictus Deus et Pater Domini nostri Iesu Christi Pater misericordiarum et Deus totius consolationis
2COR|1|4|qui consolatur nos in omni tribulatione nostra ut possimus et ipsi consolari eos qui in omni pressura sunt per exhortationem qua exhortamur et ipsi a Deo
2COR|1|5|quoniam sicut abundant passiones Christi in nobis ita et per Christum abundat consolatio nostra
2COR|1|6|sive autem tribulamur pro vestra exhortatione et salute sive exhortamur pro vestra exhortatione quae operatur in tolerantia earundem passionum quas et nos patimur
2COR|1|7|et spes nostra firma pro vobis scientes quoniam sicut socii passionum estis sic eritis et consolationis
2COR|1|8|non enim volumus ignorare vos fratres de tribulatione nostra quae facta est in Asia quoniam supra modum gravati sumus supra virtutem ita ut taederet nos etiam vivere
2COR|1|9|sed ipsi in nobis ipsis responsum mortis habuimus ut non simus fidentes in nobis sed in Deo qui suscitat mortuos
2COR|1|10|qui de tantis periculis eripuit nos et eruet in quem speramus quoniam et adhuc eripiet
2COR|1|11|adiuvantibus et vobis in oratione pro nobis ut ex multis personis eius quae in nobis est donationis per multos gratiae agantur pro nobis
2COR|1|12|nam gloria nostra haec est testimonium conscientiae nostrae quod in simplicitate et sinceritate Dei et non in sapientia carnali sed in gratia Dei conversati sumus in mundo abundantius autem ad vos
2COR|1|13|non enim alia scribimus vobis quam quae legistis et cognoscitis spero autem quod usque in finem cognoscetis
2COR|1|14|sicut et cognovistis nos ex parte quia gloria vestra sumus sicut et vos nostra in die Domini nostri Iesu Christi
2COR|1|15|et hac confidentia volui prius venire ad vos ut secundam gratiam haberetis
2COR|1|16|et per vos transire in Macedoniam et iterum a Macedonia venire ad vos et a vobis deduci in Iudaeam
2COR|1|17|cum hoc ergo voluissem numquid levitate usus sum aut quae cogito secundum carnem cogito ut sit apud me est et non
2COR|1|18|fidelis autem Deus quia sermo noster qui fit apud vos non est in illo est et non
2COR|1|19|Dei enim Filius Iesus Christus qui in vobis per nos praedicatus est per me et Silvanum et Timotheum non fuit est et non sed est in illo fuit
2COR|1|20|quotquot enim promissiones Dei sunt in illo est ideo et per ipsum amen Deo ad gloriam nostram
2COR|1|21|qui autem confirmat nos vobiscum in Christum et qui unxit nos Deus
2COR|1|22|et qui signavit nos et dedit pignus Spiritus in cordibus nostris
2COR|1|23|ego autem testem Deum invoco in animam meam quod parcens vobis non veni ultra Corinthum
2COR|1|24|non quia dominamur fidei vestrae sed adiutores sumus gaudii vestri nam fide stetistis
2COR|2|1|statui autem hoc ipse apud me ne iterum in tristitia venirem ad vos
2COR|2|2|si enim ego contristo vos et quis est qui me laetificet nisi qui contristatur ex me
2COR|2|3|et hoc ipsum scripsi ut non cum venero tristitiam super tristitiam habeam de quibus oportuerat me gaudere confidens in omnibus vobis quia meum gaudium omnium vestrum est
2COR|2|4|nam ex multa tribulatione et angustia cordis scripsi vobis per multas lacrimas non ut contristemini sed ut sciatis quam caritatem habeo abundantius in vobis
2COR|2|5|si quis autem contristavit non me contristavit sed ex parte ut non onerem omnes vos
2COR|2|6|sufficit illi qui eiusmodi est obiurgatio haec quae fit a pluribus
2COR|2|7|ita ut e contra magis donetis et consolemini ne forte abundantiori tristitia absorbeatur qui eiusmodi est
2COR|2|8|propter quod obsecro vos ut confirmetis in illum caritatem
2COR|2|9|ideo enim et scripsi ut cognoscam experimentum vestrum an in omnibus oboedientes sitis
2COR|2|10|cui autem aliquid donatis et ego nam et ego quod donavi si quid donavi propter vos in persona Christi
2COR|2|11|ut non circumveniamur a Satana non enim ignoramus cogitationes eius
2COR|2|12|cum venissem autem Troadem propter evangelium Christi et ostium mihi apertum esset in Domino
2COR|2|13|non habui requiem spiritui meo eo quod non invenerim Titum fratrem meum sed valefaciens eis profectus sum in Macedoniam
2COR|2|14|Deo autem gratias qui semper triumphat nos in Christo Iesu et odorem notitiae suae manifestat per nos in omni loco
2COR|2|15|quia Christi bonus odor sumus Deo in his qui salvi fiunt et in his qui pereunt
2COR|2|16|aliis quidem odor mortis in mortem aliis autem odor vitae in vitam et ad haec quis tam idoneus
2COR|2|17|non enim sumus sicut plurimi adulterantes verbum Dei sed ex sinceritate sed sicut ex Deo coram Deo in Christo loquimur
2COR|3|1|incipimus iterum nosmet ipsos commendare aut numquid egemus sicut quidam commendaticiis epistulis ad vos aut ex vobis
2COR|3|2|epistula nostra vos estis scripta in cordibus nostris quae scitur et legitur ab omnibus hominibus
2COR|3|3|manifestati quoniam epistula estis Christi ministrata a nobis et scripta non atramento sed Spiritu Dei vivi non in tabulis lapideis sed in tabulis cordis carnalibus
2COR|3|4|fiduciam autem talem habemus per Christum ad Deum
2COR|3|5|non quod sufficientes simus cogitare aliquid a nobis quasi ex nobis sed sufficientia nostra ex Deo est
2COR|3|6|qui et idoneos nos fecit ministros novi testamenti non litterae sed Spiritus littera enim occidit Spiritus autem vivificat
2COR|3|7|quod si ministratio mortis litteris deformata in lapidibus fuit in gloria ita ut non possent intendere filii Israhel in faciem Mosi propter gloriam vultus eius quae evacuatur
2COR|3|8|quomodo non magis ministratio Spiritus erit in gloria
2COR|3|9|nam si ministratio damnationis gloria est multo magis abundat ministerium iustitiae in gloria
2COR|3|10|nam nec glorificatum est quod claruit in hac parte propter excellentem gloriam
2COR|3|11|si enim quod evacuatur per gloriam est multo magis quod manet in gloria est
2COR|3|12|habentes igitur talem spem multa fiducia utimur
2COR|3|13|et non sicut Moses ponebat velamen super faciem suam ut non intenderent filii Israhel in faciem eius quod evacuatur
2COR|3|14|sed obtusi sunt sensus eorum usque in hodiernum enim diem id ipsum velamen in lectione veteris testamenti manet non revelatum quoniam in Christo evacuatur
2COR|3|15|sed usque in hodiernum diem cum legitur Moses velamen est positum super cor eorum
2COR|3|16|cum autem conversus fuerit ad Deum aufertur velamen
2COR|3|17|Dominus autem Spiritus est ubi autem Spiritus Domini ibi libertas
2COR|3|18|nos vero omnes revelata facie gloriam Domini speculantes in eandem imaginem transformamur a claritate in claritatem tamquam a Domini Spiritu
2COR|4|1|ideo habentes hanc ministrationem iuxta quod misericordiam consecuti sumus non deficimus
2COR|4|2|sed abdicamus occulta dedecoris non ambulantes in astutia neque adulterantes verbum Dei sed in manifestatione veritatis commendantes nosmet ipsos ad omnem conscientiam hominum coram Deo
2COR|4|3|quod si etiam opertum est evangelium nostrum in his qui pereunt est opertum
2COR|4|4|in quibus deus huius saeculi excaecavit mentes infidelium ut non fulgeat inluminatio evangelii gloriae Christi qui est imago Dei
2COR|4|5|non enim nosmet ipsos praedicamus sed Iesum Christum Dominum nos autem servos vestros per Iesum
2COR|4|6|quoniam Deus qui dixit de tenebris lucem splendescere qui inluxit in cordibus nostris ad inluminationem scientiae claritatis Dei in facie Christi Iesu
2COR|4|7|habemus autem thesaurum istum in vasis fictilibus ut sublimitas sit virtutis Dei et non ex nobis
2COR|4|8|in omnibus tribulationem patimur sed non angustiamur aporiamur sed non destituimur
2COR|4|9|persecutionem patimur sed non derelinquimur deicimur sed non perimus
2COR|4|10|semper mortificationem Iesu in corpore nostro circumferentes ut et vita Iesu in corporibus nostris manifestetur
2COR|4|11|semper enim nos qui vivimus in mortem tradimur propter Iesum ut et vita Iesu manifestetur in carne nostra mortali
2COR|4|12|ergo mors in nobis operatur vita autem in vobis
2COR|4|13|habentes autem eundem spiritum fidei sicut scriptum est credidi propter quod locutus sum et nos credimus propter quod et loquimur
2COR|4|14|scientes quoniam qui suscitavit Iesum et nos cum Iesu suscitabit et constituet vobiscum
2COR|4|15|omnia enim propter vos ut gratia abundans per multos gratiarum actione abundet in gloriam Dei
2COR|4|16|propter quod non deficimus sed licet is qui foris est noster homo corrumpitur tamen is qui intus est renovatur de die in diem
2COR|4|17|id enim quod in praesenti est momentaneum et leve tribulationis nostrae supra modum in sublimitatem aeternum gloriae pondus operatur nobis
2COR|4|18|non contemplantibus nobis quae videntur sed quae non videntur quae enim videntur temporalia sunt quae autem non videntur aeterna sunt
2COR|5|1|scimus enim quoniam si terrestris domus nostra huius habitationis dissolvatur quod aedificationem ex Deo habeamus domum non manufactam aeternam in caelis
2COR|5|2|nam et in hoc ingemescimus habitationem nostram quae de caelo est superindui cupientes
2COR|5|3|si tamen vestiti non nudi inveniamur
2COR|5|4|nam et qui sumus in tabernaculo ingemescimus gravati eo quod nolumus expoliari sed supervestiri ut absorbeatur quod mortale est a vita
2COR|5|5|qui autem efficit nos in hoc ipsum Deus qui dedit nobis pignus Spiritus
2COR|5|6|audentes igitur semper et scientes quoniam dum sumus in corpore peregrinamur a Domino
2COR|5|7|per fidem enim ambulamus et non per speciem
2COR|5|8|audemus autem et bonam voluntatem habemus magis peregrinari a corpore et praesentes esse ad Deum
2COR|5|9|et ideo contendimus sive absentes sive praesentes placere illi
2COR|5|10|omnes enim nos manifestari oportet ante tribunal Christi ut referat unusquisque propria corporis prout gessit sive bonum sive malum
2COR|5|11|scientes ergo timorem Domini hominibus suademus Deo autem manifesti sumus spero autem et in conscientiis vestris manifestos nos esse
2COR|5|12|non iterum nos commendamus vobis sed occasionem damus vobis gloriandi pro nobis ut habeatis ad eos qui in facie gloriantur et non in corde
2COR|5|13|sive enim mente excedimus Deo sive sobrii sumus vobis
2COR|5|14|caritas enim Christi urget nos aestimantes hoc quoniam si unus pro omnibus mortuus est ergo omnes mortui sunt
2COR|5|15|et pro omnibus mortuus est ut et qui vivunt iam non sibi vivant sed ei qui pro ipsis mortuus est et resurrexit
2COR|5|16|itaque nos ex hoc neminem novimus secundum carnem et si cognovimus secundum carnem Christum sed nunc iam non novimus
2COR|5|17|si qua ergo in Christo nova creatura vetera transierunt ecce facta sunt nova
2COR|5|18|omnia autem ex Deo qui reconciliavit nos sibi per Christum et dedit nobis ministerium reconciliationis
2COR|5|19|quoniam quidem Deus erat in Christo mundum reconcilians sibi non reputans illis delicta ipsorum et posuit in nobis verbum reconciliationis
2COR|5|20|pro Christo ergo legationem fungimur tamquam Deo exhortante per nos obsecramus pro Christo reconciliamini Deo
2COR|5|21|eum qui non noverat peccatum pro nobis peccatum fecit ut nos efficeremur iustitia Dei in ipso
2COR|6|1|adiuvantes autem et exhortamur ne in vacuum gratiam Dei recipiatis
2COR|6|2|ait enim tempore accepto exaudivi te et in die salutis adiuvavi te ecce nunc tempus acceptabile ecce nunc dies salutis
2COR|6|3|nemini dantes ullam offensionem ut non vituperetur ministerium
2COR|6|4|sed in omnibus exhibeamus nosmet ipsos sicut Dei ministros in multa patientia in tribulationibus in necessitatibus in angustiis
2COR|6|5|in plagis in carceribus in seditionibus in laboribus in vigiliis in ieiuniis
2COR|6|6|in castitate in scientia in longanimitate in suavitate in Spiritu Sancto in caritate non ficta
2COR|6|7|in verbo veritatis in virtute Dei per arma iustitiae a dextris et sinistris
2COR|6|8|per gloriam et ignobilitatem per infamiam et bonam famam ut seductores et veraces sicut qui ignoti et cogniti
2COR|6|9|quasi morientes et ecce vivimus ut castigati et non mortificati
2COR|6|10|quasi tristes semper autem gaudentes sicut egentes multos autem locupletantes tamquam nihil habentes et omnia possidentes
2COR|6|11|os nostrum patet ad vos o Corinthii cor nostrum dilatatum est
2COR|6|12|non angustiamini in nobis angustiamini autem in visceribus vestris
2COR|6|13|eandem autem habentes remunerationem tamquam filiis dico dilatamini et vos
2COR|6|14|nolite iugum ducere cum infidelibus quae enim participatio iustitiae cum iniquitate aut quae societas luci ad tenebras
2COR|6|15|quae autem conventio Christi ad Belial aut quae pars fideli cum infidele
2COR|6|16|qui autem consensus templo Dei cum idolis vos enim estis templum Dei vivi sicut dicit Deus quoniam inhabitabo in illis et inambulabo et ero illorum Deus et ipsi erunt mihi populus
2COR|6|17|propter quod exite de medio eorum et separamini dicit Dominus et inmundum ne tetigeritis
2COR|6|18|et ego recipiam vos et ero vobis in patrem et vos eritis mihi in filios et filias dicit Dominus omnipotens
2COR|7|1|has igitur habentes promissiones carissimi mundemus nos ab omni inquinamento carnis et spiritus perficientes sanctificationem in timore Dei
2COR|7|2|capite nos neminem laesimus neminem corrupimus neminem circumvenimus
2COR|7|3|non ad condemnationem dico praedixi enim quod in cordibus nostris estis ad conmoriendum et ad convivendum
2COR|7|4|multa mihi fiducia est apud vos multa mihi gloriatio pro vobis repletus sum consolatione superabundo gaudio in omni tribulatione nostra
2COR|7|5|nam et cum venissemus Macedoniam nullam requiem habuit caro nostra sed omnem tribulationem passi foris pugnae intus timores
2COR|7|6|sed qui consolatur humiles consolatus est nos Deus in adventu Titi
2COR|7|7|non solum autem in adventu eius sed etiam in solacio quo consolatus est in vobis referens nobis vestrum desiderium vestrum fletum vestram aemulationem pro me ita ut magis gauderem
2COR|7|8|quoniam et si contristavi vos in epistula non me paenitet et si paeniteret videns quod epistula illa et si ad horam vos contristavit
2COR|7|9|nunc gaudeo non quia contristati estis sed quia contristati estis ad paenitentiam contristati enim estis secundum Deum ut in nullo detrimentum patiamini ex nobis
2COR|7|10|quae enim secundum Deum tristitia est paenitentiam in salutem stabilem operatur saeculi autem tristitia mortem operatur
2COR|7|11|ecce enim hoc ipsum secundum Deum contristari vos quantam in vobis operatur sollicitudinem sed defensionem sed indignationem sed timorem sed desiderium sed aemulationem sed vindictam in omnibus exhibuistis vos incontaminatos esse negotio
2COR|7|12|igitur et si scripsi vobis non propter eum qui fecit iniuriam nec propter eum qui passus est sed ad manifestandam sollicitudinem nostram quam pro vobis habemus ad vos coram Deo
2COR|7|13|ideo consolati sumus in consolatione autem nostra abundantius magis gavisi sumus super gaudium Titi quia refectus est spiritus eius ab omnibus vobis
2COR|7|14|et si quid apud illum de vobis gloriatus sum non sum confusus sed sicut omnia vobis in veritate locuti sumus ita et gloriatio nostra quae fuit ad Titum veritas facta est
2COR|7|15|et viscera eius abundantius in vos sunt reminiscentis omnium vestrum oboedientiam quomodo cum timore et tremore excepistis eum
2COR|7|16|gaudeo quod in omnibus confido in vobis
2COR|8|1|notam autem facimus vobis fratres gratiam Dei quae data est in ecclesiis Macedoniae
2COR|8|2|quod in multo experimento tribulationis abundantia gaudii ipsorum et altissima paupertas eorum abundavit in divitias simplicitatis eorum
2COR|8|3|quia secundum virtutem testimonium illis reddo et supra virtutem voluntarii fuerunt
2COR|8|4|cum multa exhortatione obsecrantes nos gratiam et communicationem ministerii quod fit in sanctos
2COR|8|5|et non sicut speravimus sed semet ipsos dederunt primum Domino deinde nobis per voluntatem Dei
2COR|8|6|ita ut rogaremus Titum ut quemadmodum coepit ita et perficiat in vos etiam gratiam istam
2COR|8|7|sed sicut in omnibus abundatis fide et sermone et scientia et omni sollicitudine et caritate vestra in nos ut et in hac gratia abundetis
2COR|8|8|non quasi imperans dico sed per aliorum sollicitudinem etiam vestrae caritatis ingenitum bonum conprobans
2COR|8|9|scitis enim gratiam Domini nostri Iesu Christi quoniam propter vos egenus factus est cum esset dives ut illius inopia vos divites essetis
2COR|8|10|et consilium in hoc do hoc enim vobis utile est qui non solum facere sed et velle coepistis ab anno priore
2COR|8|11|nunc vero et facto perficite ut quemadmodum promptus est animus voluntatis ita sit et perficiendi ex eo quod habetis
2COR|8|12|si enim voluntas prompta est secundum id quod habet accepta est non secundum quod non habet
2COR|8|13|non enim ut aliis sit remissio vobis autem tribulatio sed ex aequalitate
2COR|8|14|in praesenti tempore vestra abundantia illorum inopiam suppleat ut et illorum abundantia vestrae inopiae sit supplementum ut fiat aequalitas sicut scriptum est
2COR|8|15|qui multum non abundavit et qui modicum non minoravit
2COR|8|16|gratias autem Deo qui dedit eandem sollicitudinem pro vobis in corde Titi
2COR|8|17|quoniam exhortationem quidem suscepit sed cum sollicitior esset sua voluntate profectus est ad vos
2COR|8|18|misimus etiam cum illo fratrem cuius laus est in evangelio per omnes ecclesias
2COR|8|19|non solum autem sed et ordinatus ab ecclesiis comes peregrinationis nostrae in hac gratia quae ministratur a nobis ad Domini gloriam et destinatam voluntatem nostram
2COR|8|20|devitantes hoc ne quis nos vituperet in hac plenitudine quae ministratur a nobis
2COR|8|21|providemus enim bona non solum coram Deo sed etiam coram hominibus
2COR|8|22|misimus autem cum illis et fratrem nostrum quem probavimus in multis saepe sollicitum esse nunc autem multo sollicitiorem confidentia multa in vos
2COR|8|23|sive pro Tito qui est socius meus et in vos adiutor sive fratres nostri apostoli ecclesiarum gloriae Christi
2COR|8|24|ostensionem ergo quae est caritatis vestrae et nostrae gloriae pro vobis in illos ostendite in faciem ecclesiarum
2COR|9|1|nam de ministerio quod fit in sanctos ex abundanti est mihi scribere vobis
2COR|9|2|scio enim promptum animum vestrum pro quo de vobis glorior apud Macedonas quoniam Achaia parata est ab anno praeterito et vestra aemulatio provocavit plurimos
2COR|9|3|misi autem fratres ut ne quod gloriamur de vobis evacuetur in hac parte ut quemadmodum dixi parati sitis
2COR|9|4|ne cum venerint mecum Macedones et invenerint vos inparatos erubescamus nos ut non dicamus vos in hac substantia
2COR|9|5|necessarium ergo existimavi rogare fratres ut praeveniant ad vos et praeparent repromissam benedictionem hanc paratam esse sic quasi benedictionem non quasi avaritiam
2COR|9|6|hoc autem qui parce seminat parce et metet et qui seminat in benedictionibus de benedictionibus et metet
2COR|9|7|unusquisque prout destinavit corde suo non ex tristitia aut ex necessitate hilarem enim datorem diligit Deus
2COR|9|8|potens est autem Deus omnem gratiam abundare facere in vobis ut in omnibus semper omnem sufficientiam habentes abundetis in omne opus bonum
2COR|9|9|sicut scriptum est dispersit dedit pauperibus iustitia eius manet in aeternum
2COR|9|10|qui autem administrat semen seminanti et panem ad manducandum praestabit et multiplicabit semen vestrum et augebit incrementa frugum iustitiae vestrae
2COR|9|11|ut in omnibus locupletati abundetis in omnem simplicitatem quae operatur per nos gratiarum actionem Deo
2COR|9|12|quoniam ministerium huius officii non solum supplet ea quae desunt sanctis sed etiam abundat per multas gratiarum actiones in Domino
2COR|9|13|per probationem ministerii huius glorificantes Deum in oboedientia confessionis vestrae in evangelium Christi et simplicitate communicationis in illos et in omnes
2COR|9|14|et ipsorum obsecratione pro vobis desiderantium vos propter eminentem gratiam Dei in vobis
2COR|9|15|gratias Deo super inenarrabili dono eius
2COR|10|1|ipse autem ego Paulus obsecro vos per mansuetudinem et modestiam Christi qui in facie quidem humilis inter vos absens autem confido in vobis
2COR|10|2|rogo autem ne praesens audeam per eam confidentiam qua existimo audere in quosdam qui arbitrantur nos tamquam secundum carnem ambulemus
2COR|10|3|in carne enim ambulantes non secundum carnem militamus
2COR|10|4|nam arma militiae nostrae non carnalia sed potentia Deo ad destructionem munitionum consilia destruentes
2COR|10|5|et omnem altitudinem extollentem se adversus scientiam Dei et in captivitatem redigentes omnem intellectum in obsequium Christi
2COR|10|6|et in promptu habentes ulcisci omnem inoboedientiam cum impleta fuerit vestra oboedientia
2COR|10|7|quae secundum faciem sunt videte si quis confidit sibi Christi se esse hoc cogitet iterum apud se quia sicut ipse Christi est ita et nos
2COR|10|8|nam et si amplius aliquid gloriatus fuero de potestate nostra quam dedit Dominus in aedificationem et non in destructionem vestram non erubescam
2COR|10|9|ut autem non existimer tamquam terrere vos per epistulas
2COR|10|10|quoniam quidem epistulae inquiunt graves sunt et fortes praesentia autem corporis infirma et sermo contemptibilis
2COR|10|11|hoc cogitet qui eiusmodi est quia quales sumus verbo per epistulas absentes tales et praesentes in facto
2COR|10|12|non enim audemus inserere aut conparare nos quibusdam qui se ipsos commendant sed ipsi in nobis nosmet ipsos metientes et conparantes nosmet ipsos nobis
2COR|10|13|nos autem non in inmensum gloriabimur sed secundum mensuram regulae quam mensus est nobis Deus mensuram pertingendi usque ad vos
2COR|10|14|non enim quasi non pertingentes ad vos superextendimus nos usque ad vos enim pervenimus in evangelio Christi
2COR|10|15|non in inmensum gloriantes in alienis laboribus spem autem habentes crescentis fidei vestrae in vobis magnificari secundum regulam nostram in abundantiam
2COR|10|16|etiam in illa quae ultra vos sunt evangelizare non in aliena regula in his quae praeparata sunt gloriari
2COR|10|17|qui autem gloriatur in Domino glorietur
2COR|10|18|non enim qui se ipsum commendat ille probatus est sed quem Dominus commendat
2COR|11|1|utinam sustineretis modicum quid insipientiae meae sed et subportate me
2COR|11|2|aemulor enim vos Dei aemulatione despondi enim vos uni viro virginem castam exhibere Christo
2COR|11|3|timeo autem ne sicut serpens Evam seduxit astutia sua ita corrumpantur sensus vestri et excidant a simplicitate quae est in Christo
2COR|11|4|nam si is qui venit alium Christum praedicat quem non praedicavimus aut alium spiritum accipitis quem non accepistis aut aliud evangelium quod non recepistis recte pateremini
2COR|11|5|existimo enim nihil me minus fecisse magnis apostolis
2COR|11|6|et si inperitus sermone sed non scientia in omnibus autem manifestatus sum vobis
2COR|11|7|aut numquid peccatum feci me ipsum humilians ut vos exaltemini quoniam gratis evangelium Dei evangelizavi vobis
2COR|11|8|alias ecclesias expoliavi accipiens stipendium ad ministerium vestrum
2COR|11|9|et cum essem apud vos et egerem nulli onerosus fui nam quod mihi deerat suppleverunt fratres qui venerunt a Macedonia et in omnibus sine onere me vobis servavi et servabo
2COR|11|10|est veritas Christi in me quoniam haec gloria non infringetur in me in regionibus Achaiae
2COR|11|11|quare quia non diligo vos Deus scit
2COR|11|12|quod autem facio et faciam ut amputem occasionem eorum qui volunt occasionem ut in quo gloriantur inveniantur sicut et nos
2COR|11|13|nam eiusmodi pseudoapostoli operarii subdoli transfigurantes se in apostolos Christi
2COR|11|14|et non mirum ipse enim Satanas transfigurat se in angelum lucis
2COR|11|15|non est ergo magnum si ministri eius transfigurentur velut ministri iustitiae quorum finis erit secundum opera ipsorum
2COR|11|16|iterum dico ne quis me putet insipientem alioquin velut insipientem accipite me ut et ego modicum quid glorier
2COR|11|17|quod loquor non loquor secundum Dominum sed quasi in insipientia in hac substantia gloriae
2COR|11|18|quoniam multi gloriantur secundum carnem et ego gloriabor
2COR|11|19|libenter enim suffertis insipientes cum sitis ipsi sapientes
2COR|11|20|sustinetis enim si quis vos in servitutem redigit si quis devorat si quis accipit si quis extollitur si quis in faciem vos caedit
2COR|11|21|secundum ignobilitatem dico quasi nos infirmi fuerimus in quo quis audet in insipientia dico audeo et ego
2COR|11|22|Hebraei sunt et ego Israhelitae sunt et ego semen Abrahae sunt et ego
2COR|11|23|ministri Christi sunt minus sapiens dico plus ego in laboribus plurimis in carceribus abundantius in plagis supra modum in mortibus frequenter
2COR|11|24|a Iudaeis quinquies quadragenas una minus accepi
2COR|11|25|ter virgis caesus sum semel lapidatus sum ter naufragium feci nocte et die in profundo maris fui
2COR|11|26|in itineribus saepe periculis fluminum periculis latronum periculis ex genere periculis ex gentibus periculis in civitate periculis in solitudine periculis in mari periculis in falsis fratribus
2COR|11|27|in labore et aerumna in vigiliis multis in fame et siti in ieiuniis multis in frigore et nuditate
2COR|11|28|praeter illa quae extrinsecus sunt instantia mea cotidiana sollicitudo omnium ecclesiarum
2COR|11|29|quis infirmatur et non infirmor quis scandalizatur et ego non uror
2COR|11|30|si gloriari oportet quae infirmitatis meae sunt gloriabor
2COR|11|31|Deus et Pater Domini Iesu scit qui est benedictus in saecula quod non mentior
2COR|11|32|Damasci praepositus gentis Aretae regis custodiebat civitatem Damascenorum ut me conprehenderet
2COR|11|33|et per fenestram in sporta dimissus sum per murum et effugi manus eius
2COR|12|1|si gloriari oportet non expedit quidem veniam autem ad visiones et revelationes Domini
2COR|12|2|scio hominem in Christo ante annos quattuordecim sive in corpore nescio sive extra corpus nescio Deus scit raptum eiusmodi usque ad tertium caelum
2COR|12|3|et scio huiusmodi hominem sive in corpore sive extra corpus nescio Deus scit
2COR|12|4|quoniam raptus est in paradisum et audivit arcana verba quae non licet homini loqui
2COR|12|5|pro eiusmodi gloriabor pro me autem nihil gloriabor nisi in infirmitatibus meis
2COR|12|6|nam et si voluero gloriari non ero insipiens veritatem enim dicam parco autem ne quis in me existimet supra id quod videt me aut audit ex me
2COR|12|7|et ne magnitudo revelationum extollat me datus est mihi stimulus carnis meae angelus Satanae ut me colaphizet
2COR|12|8|propter quod ter Dominum rogavi ut discederet a me
2COR|12|9|et dixit mihi sufficit tibi gratia mea nam virtus in infirmitate perficitur libenter igitur gloriabor in infirmitatibus meis ut inhabitet in me virtus Christi
2COR|12|10|propter quod placeo mihi in infirmitatibus in contumeliis in necessitatibus in persecutionibus in angustiis pro Christo cum enim infirmor tunc potens sum
2COR|12|11|factus sum insipiens vos me coegistis ego enim debui a vobis commendari nihil enim minus fui ab his qui sunt supra modum apostoli tametsi nihil sum
2COR|12|12|signa tamen apostoli facta sunt super vos in omni patientia signis et prodigiis et virtutibus
2COR|12|13|quid est enim quod minus habuistis prae ceteris ecclesiis nisi quod ego ipse non gravavi vos donate mihi hanc iniuriam
2COR|12|14|ecce tertio hoc paratus sum venire ad vos et non ero gravis vobis non enim quaero quae vestra sunt sed vos nec enim debent filii parentibus thesaurizare sed parentes filiis
2COR|12|15|ego autem libentissime inpendam et superinpendar ipse pro animabus vestris licet plus vos diligens minus diligar
2COR|12|16|sed esto ego vos non gravavi sed cum essem astutus dolo vos cepi
2COR|12|17|numquid per aliquem eorum quos misi ad vos circumveni vos
2COR|12|18|rogavi Titum et misi cum illo fratrem numquid Titus vos circumvenit nonne eodem spiritu ambulavimus nonne hisdem vestigiis
2COR|12|19|olim putatis quod excusemus nos apud vos coram Deo in Christo loquimur omnia autem carissimi propter vestram aedificationem
2COR|12|20|timeo enim ne forte cum venero non quales volo inveniam vos et ego inveniar a vobis qualem non vultis ne forte contentiones aemulationes animositates dissensiones detractiones susurrationes inflationes seditiones sint inter vos
2COR|12|21|ne iterum cum venero humiliet me Deus apud vos et lugeam multos ex his qui ante peccaverunt et non egerunt paenitentiam super inmunditia et fornicatione et inpudicitia quam gesserunt
2COR|13|1|ecce tertio hoc venio ad vos in ore duorum vel trium testium stabit omne verbum
2COR|13|2|praedixi et praedico ut praesens bis et nunc absens his qui ante peccaverunt et ceteris omnibus quoniam si venero iterum non parcam
2COR|13|3|an experimentum quaeritis eius qui in me loquitur Christi qui in vos non infirmatur sed potens est in vobis
2COR|13|4|nam et si crucifixus est ex infirmitate sed vivit ex virtute Dei nam et nos infirmi sumus in illo sed vivemus cum eo ex virtute Dei in vobis
2COR|13|5|vosmet ipsos temptate si estis in fide ipsi vos probate an non cognoscitis vos ipsos quia Christus Iesus in vobis est nisi forte reprobi estis
2COR|13|6|spero autem quod cognoscetis quia nos non sumus reprobi
2COR|13|7|oramus autem Deum ut nihil mali faciatis non ut nos probati pareamus sed ut vos quod bonum est faciatis nos autem ut reprobi simus
2COR|13|8|non enim possumus aliquid adversus veritatem sed pro veritate
2COR|13|9|gaudemus enim quando nos infirmi sumus vos autem potentes estis hoc et oramus vestram consummationem
2COR|13|10|ideo haec absens scribo ut non praesens durius agam secundum potestatem quam Dominus dedit mihi in aedificationem et non in destructionem
2COR|13|11|de cetero fratres gaudete perfecti estote exhortamini idem sapite pacem habete et Deus dilectionis et pacis erit vobiscum
2COR|13|12|salutate invicem in osculo sancto salutant vos sancti omnes
2COR|13|13|gratia Domini nostri Iesu Christi et caritas Dei et communicatio Sancti Spiritus cum omnibus vobis amen
GAL|1|1|Paulus apostolus non ab hominibus neque per hominem sed per Iesum Christum et Deum Patrem qui suscitavit eum a mortuis
GAL|1|2|et qui mecum sunt omnes fratres ecclesiis Galatiae
GAL|1|3|gratia vobis et pax a Deo Patre et Domino nostro Iesu Christo
GAL|1|4|qui dedit semet ipsum pro peccatis nostris ut eriperet nos de praesenti saeculo nequam secundum voluntatem Dei et Patris nostri
GAL|1|5|cui est gloria in saecula saeculorum amen
GAL|1|6|miror quod sic tam cito transferimini ab eo qui vos vocavit in gratiam Christi in aliud evangelium
GAL|1|7|quod non est aliud nisi sunt aliqui qui vos conturbant et volunt convertere evangelium Christi
GAL|1|8|sed licet nos aut angelus de caelo evangelizet vobis praeterquam quod evangelizavimus vobis anathema sit
GAL|1|9|sicut praediximus et nunc iterum dico si quis vobis evangelizaverit praeter id quod accepistis anathema sit
GAL|1|10|modo enim hominibus suadeo aut Deo aut quaero hominibus placere si adhuc hominibus placerem Christi servus non essem
GAL|1|11|notum enim vobis facio fratres evangelium quod evangelizatum est a me quia non est secundum hominem
GAL|1|12|neque enim ego ab homine accepi illud neque didici sed per revelationem Iesu Christi
GAL|1|13|audistis enim conversationem meam aliquando in iudaismo quoniam supra modum persequebar ecclesiam Dei et expugnabam illam
GAL|1|14|et proficiebam in iudaismo supra multos coetaneos in genere meo abundantius aemulator existens paternarum mearum traditionum
GAL|1|15|cum autem placuit ei qui me segregavit de utero matris meae et vocavit per gratiam suam
GAL|1|16|ut revelaret Filium suum in me ut evangelizarem illum in gentibus continuo non adquievi carni et sanguini
GAL|1|17|neque veni Hierosolyma ad antecessores meos apostolos sed abii in Arabiam et iterum reversus sum Damascum
GAL|1|18|deinde post annos tres veni Hierosolyma videre Petrum et mansi apud eum diebus quindecim
GAL|1|19|alium autem apostolorum vidi neminem nisi Iacobum fratrem Domini
GAL|1|20|quae autem scribo vobis ecce coram Deo quia non mentior
GAL|1|21|deinde veni in partes Syriae et Ciliciae
GAL|1|22|eram autem ignotus facie ecclesiis Iudaeae quae erant in Christo
GAL|1|23|tantum autem auditum habebant quoniam qui persequebatur nos aliquando nunc evangelizat fidem quam aliquando expugnabat
GAL|1|24|et in me clarificabant Deum
GAL|2|1|deinde post annos quattuordecim iterum ascendi Hierosolyma cum Barnaba adsumpto et Tito
GAL|2|2|ascendi autem secundum revelationem et contuli cum illis evangelium quod praedico in gentibus seorsum autem his qui videbantur ne forte in vacuum currerem aut cucurrissem
GAL|2|3|sed neque Titus qui mecum erat cum esset gentilis conpulsus est circumcidi
GAL|2|4|sed propter subintroductos falsos fratres qui subintroierunt explorare libertatem nostram quam habemus in Christo Iesu ut nos in servitutem redigerent
GAL|2|5|quibus neque ad horam cessimus subiectioni ut veritas evangelii permaneat apud vos
GAL|2|6|ab his autem qui videbantur esse aliquid quales aliquando fuerint nihil mea interest Deus personam hominis non accipit mihi enim qui videbantur nihil contulerunt
GAL|2|7|sed e contra cum vidissent quod creditum est mihi evangelium praeputii sicut Petro circumcisionis
GAL|2|8|qui enim operatus est Petro in apostolatum circumcisionis operatus est et mihi inter gentes
GAL|2|9|et cum cognovissent gratiam quae data est mihi Iacobus et Cephas et Iohannes qui videbantur columnae esse dextras dederunt mihi et Barnabae societatis ut nos in gentes ipsi autem in circumcisionem
GAL|2|10|tantum ut pauperum memores essemus quod etiam sollicitus fui hoc ipsum facere
GAL|2|11|cum autem venisset Cephas Antiochiam in faciem ei restiti quia reprehensibilis erat
GAL|2|12|prius enim quam venirent quidam ab Iacobo cum gentibus edebat cum autem venissent subtrahebat et segregabat se timens eos qui ex circumcisione erant
GAL|2|13|et simulationi eius consenserunt ceteri Iudaei ita ut et Barnabas duceretur ab eis in illa simulatione
GAL|2|14|sed cum vidissem quod non recte ambularent ad veritatem evangelii dixi Cephae coram omnibus si tu cum Iudaeus sis gentiliter et non iudaice vivis quomodo gentes cogis iudaizare
GAL|2|15|nos natura Iudaei et non ex gentibus peccatores
GAL|2|16|scientes autem quod non iustificatur homo ex operibus legis nisi per fidem Iesu Christi et nos in Christo Iesu credidimus ut iustificemur ex fide Christi et non ex operibus legis propter quod ex operibus legis non iustificabitur omnis caro
GAL|2|17|quod si quaerentes iustificari in Christo inventi sumus et ipsi peccatores numquid Christus peccati minister est absit
GAL|2|18|si enim quae destruxi haec iterum aedifico praevaricatorem me constituo
GAL|2|19|ego enim per legem legi mortuus sum ut Deo vivam Christo confixus sum cruci
GAL|2|20|vivo autem iam non ego vivit vero in me Christus quod autem nunc vivo in carne in fide vivo Filii Dei qui dilexit me et tradidit se ipsum pro me
GAL|2|21|non abicio gratiam Dei si enim per legem iustitia ergo Christus gratis mortuus est
GAL|3|1|o insensati Galatae quis vos fascinavit ante quorum oculos Iesus Christus proscriptus est crucifixus
GAL|3|2|hoc solum volo a vobis discere ex operibus legis Spiritum accepistis an ex auditu fidei
GAL|3|3|sic stulti estis cum Spiritu coeperitis nunc carne consummamini
GAL|3|4|tanta passi estis sine causa si tamen sine causa
GAL|3|5|qui ergo tribuit vobis Spiritum et operatur virtutes in vobis ex operibus legis an ex auditu fidei
GAL|3|6|sicut Abraham credidit Deo et reputatum est ei ad iustitiam
GAL|3|7|cognoscitis ergo quia qui ex fide sunt hii sunt filii Abrahae
GAL|3|8|providens autem scriptura quia ex fide iustificat gentes Deus praenuntiavit Abrahae quia benedicentur in te omnes gentes
GAL|3|9|igitur qui ex fide sunt benedicentur cum fideli Abraham
GAL|3|10|quicumque enim ex operibus legis sunt sub maledicto sunt scriptum est enim maledictus omnis qui non permanserit in omnibus quae scripta sunt in libro legis ut faciat ea
GAL|3|11|quoniam autem in lege nemo iustificatur apud Deum manifestum est quia iustus ex fide vivit
GAL|3|12|lex autem non est ex fide sed qui fecerit ea vivet in illis
GAL|3|13|Christus nos redemit de maledicto legis factus pro nobis maledictum quia scriptum est maledictus omnis qui pendet in ligno
GAL|3|14|ut in gentibus benedictio Abrahae fieret in Christo Iesu ut pollicitationem Spiritus accipiamus per fidem
GAL|3|15|fratres secundum hominem dico tamen hominis confirmatum testamentum nemo spernit aut superordinat
GAL|3|16|Abrahae dictae sunt promissiones et semini eius non dicit et seminibus quasi in multis sed quasi in uno et semini tuo qui est Christus
GAL|3|17|hoc autem dico testamentum confirmatum a Deo quae post quadringentos et triginta annos facta est lex non irritam facit ad evacuandam promissionem
GAL|3|18|nam si ex lege hereditas iam non ex repromissione Abrahae autem per promissionem donavit Deus
GAL|3|19|quid igitur lex propter transgressiones posita est donec veniret semen cui promiserat ordinata per angelos in manu mediatoris
GAL|3|20|mediator autem unius non est Deus autem unus est
GAL|3|21|lex ergo adversus promissa Dei absit si enim data esset lex quae posset vivificare vere ex lege esset iustitia
GAL|3|22|sed conclusit scriptura omnia sub peccato ut promissio ex fide Iesu Christi daretur credentibus
GAL|3|23|prius autem quam veniret fides sub lege custodiebamur conclusi in eam fidem quae revelanda erat
GAL|3|24|itaque lex pedagogus noster fuit in Christo ut ex fide iustificemur
GAL|3|25|at ubi venit fides iam non sumus sub pedagogo
GAL|3|26|omnes enim filii Dei estis per fidem in Christo Iesu
GAL|3|27|quicumque enim in Christo baptizati estis Christum induistis
GAL|3|28|non est Iudaeus neque Graecus non est servus neque liber non est masculus neque femina omnes enim vos unum estis in Christo Iesu
GAL|3|29|si autem vos Christi ergo Abrahae semen estis secundum promissionem heredes
GAL|4|1|dico autem quanto tempore heres parvulus est nihil differt servo cum sit dominus omnium
GAL|4|2|sed sub tutoribus est et actoribus usque ad praefinitum tempus a patre
GAL|4|3|ita et nos cum essemus parvuli sub elementis mundi eramus servientes
GAL|4|4|at ubi venit plenitudo temporis misit Deus Filium suum factum ex muliere factum sub lege
GAL|4|5|ut eos qui sub lege erant redimeret ut adoptionem filiorum reciperemus
GAL|4|6|quoniam autem estis filii misit Deus Spiritum Filii sui in corda nostra clamantem Abba Pater
GAL|4|7|itaque iam non es servus sed filius quod si filius et heres per Deum
GAL|4|8|sed tunc quidem ignorantes Deum his qui natura non sunt dii serviebatis
GAL|4|9|nunc autem cum cognoveritis Deum immo cogniti sitis a Deo quomodo convertimini iterum ad infirma et egena elementa quibus denuo servire vultis
GAL|4|10|dies observatis et menses et tempora et annos
GAL|4|11|timeo vos ne forte sine causa laboraverim in vobis
GAL|4|12|estote sicut et ego quia et ego sicut vos fratres obsecro vos nihil me laesistis
GAL|4|13|scitis autem quia per infirmitatem carnis evangelizavi vobis iam pridem
GAL|4|14|et temptationem vestram in carne mea non sprevistis neque respuistis sed sicut angelum Dei excepistis me sicut Christum Iesum
GAL|4|15|ubi est ergo beatitudo vestra testimonium enim perhibeo vobis quia si fieri posset oculos vestros eruissetis et dedissetis mihi
GAL|4|16|ergo inimicus vobis factus sum verum dicens vobis
GAL|4|17|aemulantur vos non bene sed excludere vos volunt ut illos aemulemini
GAL|4|18|bonum autem aemulamini in bono semper et non tantum cum praesens sum apud vos
GAL|4|19|filioli mei quos iterum parturio donec formetur Christus in vobis
GAL|4|20|vellem autem esse apud vos modo et mutare vocem meam quoniam confundor in vobis
GAL|4|21|dicite mihi qui sub lege vultis esse legem non legistis
GAL|4|22|scriptum est enim quoniam Abraham duos filios habuit unum de ancilla et unum de libera
GAL|4|23|sed qui de ancilla secundum carnem natus est qui autem de libera per repromissionem
GAL|4|24|quae sunt per allegoriam dicta haec enim sunt duo testamenta unum quidem a monte Sina in servitutem generans quae est Agar
GAL|4|25|Sina enim mons est in Arabia qui coniunctus est ei quae nunc est Hierusalem et servit cum filiis eius
GAL|4|26|illa autem quae sursum est Hierusalem libera est quae est mater nostra
GAL|4|27|scriptum est enim laetare sterilis quae non paris erumpe et exclama quae non parturis quia multi filii desertae magis quam eius quae habet virum
GAL|4|28|nos autem fratres secundum Isaac promissionis filii sumus
GAL|4|29|sed quomodo tunc qui secundum carnem natus fuerat persequebatur eum qui secundum spiritum ita et nunc
GAL|4|30|sed quid dicit scriptura eice ancillam et filium eius non enim heres erit filius ancillae cum filio liberae
GAL|4|31|itaque fratres non sumus ancillae filii sed liberae qua libertate nos Christus liberavit
GAL|5|1|state et nolite iterum iugo servitutis contineri
GAL|5|2|ecce ego Paulus dico vobis quoniam si circumcidamini Christus vobis nihil proderit
GAL|5|3|testificor autem rursum omni homini circumcidenti se quoniam debitor est universae legis faciendae
GAL|5|4|evacuati estis a Christo qui in lege iustificamini a gratia excidistis
GAL|5|5|nos enim spiritu ex fide spem iustitiae expectamus
GAL|5|6|nam in Christo Iesu neque circumcisio aliquid valet neque praeputium sed fides quae per caritatem operatur
GAL|5|7|currebatis bene quis vos inpedivit veritati non oboedire
GAL|5|8|persuasio non est ex eo qui vocat vos
GAL|5|9|modicum fermentum totam massam corrumpit
GAL|5|10|ego confido in vobis in Domino quod nihil aliud sapietis qui autem conturbat vos portabit iudicium quicumque est ille
GAL|5|11|ego autem fratres si circumcisionem adhuc praedico quid adhuc persecutionem patior ergo evacuatum est scandalum crucis
GAL|5|12|utinam et abscidantur qui vos conturbant
GAL|5|13|vos enim in libertatem vocati estis fratres tantum ne libertatem in occasionem detis carnis sed per caritatem servite invicem
GAL|5|14|omnis enim lex in uno sermone impletur diliges proximum tuum sicut te ipsum
GAL|5|15|quod si invicem mordetis et comeditis videte ne ab invicem consumamini
GAL|5|16|dico autem spiritu ambulate et desiderium carnis non perficietis
GAL|5|17|caro enim concupiscit adversus spiritum spiritus autem adversus carnem haec enim invicem adversantur ut non quaecumque vultis illa faciatis
GAL|5|18|quod si spiritu ducimini non estis sub lege
GAL|5|19|manifesta autem sunt opera carnis quae sunt fornicatio inmunditia luxuria
GAL|5|20|idolorum servitus veneficia inimicitiae contentiones aemulationes irae rixae dissensiones sectae
GAL|5|21|invidiae homicidia ebrietates comesationes et his similia quae praedico vobis sicut praedixi quoniam qui talia agunt regnum Dei non consequentur
GAL|5|22|fructus autem Spiritus est caritas gaudium pax longanimitas bonitas benignitas
GAL|5|23|fides modestia continentia adversus huiusmodi non est lex
GAL|5|24|qui autem sunt Christi carnem crucifixerunt cum vitiis et concupiscentiis
GAL|5|25|si vivimus spiritu spiritu et ambulemus
GAL|5|26|non efficiamur inanis gloriae cupidi invicem provocantes invicem invidentes
GAL|6|1|fratres et si praeoccupatus fuerit homo in aliquo delicto vos qui spiritales estis huiusmodi instruite in spiritu lenitatis considerans te ipsum ne et tu tempteris
GAL|6|2|alter alterius onera portate et sic adimplebitis legem Christi
GAL|6|3|nam si quis existimat se aliquid esse cum sit nihil ipse se seducit
GAL|6|4|opus autem suum probet unusquisque et sic in semet ipso tantum gloriam habebit et non in altero
GAL|6|5|unusquisque enim onus suum portabit
GAL|6|6|communicet autem is qui catecizatur verbum ei qui se catecizat in omnibus bonis
GAL|6|7|nolite errare Deus non inridetur
GAL|6|8|quae enim seminaverit homo haec et metet quoniam qui seminat in carne sua de carne et metet corruptionem qui autem seminat in spiritu de spiritu metet vitam aeternam
GAL|6|9|bonum autem facientes non deficiamus tempore enim suo metemus non deficientes
GAL|6|10|ergo dum tempus habemus operemur bonum ad omnes maxime autem ad domesticos fidei
GAL|6|11|videte qualibus litteris scripsi vobis mea manu
GAL|6|12|quicumque volunt placere in carne hii cogunt vos circumcidi tantum ut crucis Christi persecutionem non patiantur
GAL|6|13|neque enim qui circumciduntur legem custodiunt sed volunt vos circumcidi ut in carne vestra glorientur
GAL|6|14|mihi autem absit gloriari nisi in cruce Domini nostri Iesu Christi per quem mihi mundus crucifixus est et ego mundo
GAL|6|15|in Christo enim Iesu neque circumcisio aliquid valet neque praeputium sed nova creatura
GAL|6|16|et quicumque hanc regulam secuti fuerint pax super illos et misericordia et super Israhel Dei
GAL|6|17|de cetero nemo mihi molestus sit ego enim stigmata Iesu in corpore meo porto
GAL|6|18|gratia Domini nostri Iesu Christi cum spiritu vestro fratres amen
EPH|1|1|Paulus apostolus Christi Iesu per voluntatem Dei sanctis omnibus qui sunt Ephesi et fidelibus in Christo Iesu
EPH|1|2|gratia vobis et pax a Deo Patre nostro et Domino Iesu Christo
EPH|1|3|benedictus Deus et Pater Domini nostri Iesu Christi qui benedixit nos in omni benedictione spiritali in caelestibus in Christo
EPH|1|4|sicut elegit nos in ipso ante mundi constitutionem ut essemus sancti et inmaculati in conspectu eius in caritate
EPH|1|5|qui praedestinavit nos in adoptionem filiorum per Iesum Christum in ipsum secundum propositum voluntatis suae
EPH|1|6|in laudem gloriae gratiae suae in qua gratificavit nos in dilecto
EPH|1|7|in quo habemus redemptionem per sanguinem eius remissionem peccatorum secundum divitias gratiae eius
EPH|1|8|quae superabundavit in nobis in omni sapientia et prudentia
EPH|1|9|ut notum faceret nobis sacramentum voluntatis suae secundum bonum placitum eius quod proposuit in eo
EPH|1|10|in dispensationem plenitudinis temporum instaurare omnia in Christo quae in caelis et quae in terra sunt in ipso
EPH|1|11|in quo etiam sorte vocati sumus praedestinati secundum propositum eius qui omnia operatur secundum consilium voluntatis suae
EPH|1|12|ut simus in laudem gloriae eius qui ante speravimus in Christo
EPH|1|13|in quo et vos cum audissetis verbum veritatis evangelium salutis vestrae in quo et credentes signati estis Spiritu promissionis Sancto
EPH|1|14|qui est pignus hereditatis nostrae in redemptionem adquisitionis in laudem gloriae ipsius
EPH|1|15|propterea et ego audiens fidem vestram quae est in Domino Iesu et dilectionem in omnes sanctos
EPH|1|16|non cesso gratias agens pro vobis memoriam vestri faciens in orationibus meis
EPH|1|17|ut Deus Domini nostri Iesu Christi Pater gloriae det vobis spiritum sapientiae et revelationis in agnitione eius
EPH|1|18|inluminatos oculos cordis vestri ut sciatis quae sit spes vocationis eius quae divitiae gloriae hereditatis eius in sanctis
EPH|1|19|et quae sit supereminens magnitudo virtutis eius in nos qui credidimus secundum operationem potentiae virtutis eius
EPH|1|20|quam operatus est in Christo suscitans illum a mortuis et constituens ad dexteram suam in caelestibus
EPH|1|21|supra omnem principatum et potestatem et virtutem et dominationem et omne nomen quod nominatur non solum in hoc saeculo sed et in futuro
EPH|1|22|et omnia subiecit sub pedibus eius et ipsum dedit caput supra omnia ecclesiae
EPH|1|23|quae est corpus ipsius plenitudo eius qui omnia in omnibus adimpletur
EPH|2|1|et vos cum essetis mortui delictis et peccatis vestris
EPH|2|2|in quibus aliquando ambulastis secundum saeculum mundi huius secundum principem potestatis aeris huius spiritus qui nunc operatur in filios diffidentiae
EPH|2|3|in quibus et nos omnes aliquando conversati sumus in desideriis carnis nostrae facientes voluntates carnis et cogitationum et eramus natura filii irae sicut et ceteri
EPH|2|4|Deus autem qui dives est in misericordia propter nimiam caritatem suam qua dilexit nos
EPH|2|5|et cum essemus mortui peccatis convivificavit nos Christo gratia estis salvati
EPH|2|6|et conresuscitavit et consedere fecit in caelestibus in Christo Iesu
EPH|2|7|ut ostenderet in saeculis supervenientibus abundantes divitias gratiae suae in bonitate super nos in Christo Iesu
EPH|2|8|gratia enim estis salvati per fidem et hoc non ex vobis Dei enim donum est
EPH|2|9|non ex operibus ut ne quis glorietur
EPH|2|10|ipsius enim sumus factura creati in Christo Iesu in operibus bonis quae praeparavit Deus ut in illis ambulemus
EPH|2|11|propter quod memores estote quod aliquando vos gentes in carne qui dicimini praeputium ab ea quae dicitur circumcisio in carne manufacta
EPH|2|12|quia eratis illo in tempore sine Christo alienati a conversatione Israhel et hospites testamentorum promissionis spem non habentes et sine Deo in mundo
EPH|2|13|nunc autem in Christo Iesu vos qui aliquando eratis longe facti estis prope in sanguine Christi
EPH|2|14|ipse est enim pax nostra qui fecit utraque unum et medium parietem maceriae solvens inimicitiam in carne sua
EPH|2|15|legem mandatorum decretis evacuans ut duos condat in semet ipsum in unum novum hominem faciens pacem
EPH|2|16|et reconciliet ambos in uno corpore Deo per crucem interficiens inimicitiam in semet ipso
EPH|2|17|et veniens evangelizavit pacem vobis qui longe fuistis et pacem his qui prope
EPH|2|18|quoniam per ipsum habemus accessum ambo in uno Spiritu ad Patrem
EPH|2|19|ergo iam non estis hospites et advenae sed estis cives sanctorum et domestici Dei
EPH|2|20|superaedificati super fundamentum apostolorum et prophetarum ipso summo angulari lapide Christo Iesu
EPH|2|21|in quo omnis aedificatio constructa crescit in templum sanctum in Domino
EPH|2|22|in quo et vos coaedificamini in habitaculum Dei in Spiritu
EPH|3|1|huius rei gratia ego Paulus vinctus Christi Iesu pro vobis gentibus
EPH|3|2|si tamen audistis dispensationem gratiae Dei quae data est mihi in vobis
EPH|3|3|quoniam secundum revelationem notum mihi factum est sacramentum sicut supra scripsi in brevi
EPH|3|4|prout potestis legentes intellegere prudentiam meam in mysterio Christi
EPH|3|5|quod aliis generationibus non est agnitum filiis hominum sicuti nunc revelatum est sanctis apostolis eius et prophetis in Spiritu
EPH|3|6|esse gentes coheredes et concorporales et conparticipes promissionis in Christo Iesu per evangelium
EPH|3|7|cuius factus sum minister secundum donum gratiae Dei quae data est mihi secundum operationem virtutis eius
EPH|3|8|mihi omnium sanctorum minimo data est gratia haec in gentibus evangelizare ininvestigabiles divitias Christi
EPH|3|9|et inluminare omnes quae sit dispensatio sacramenti absconditi a saeculis in Deo qui omnia creavit
EPH|3|10|ut innotescat principibus et potestatibus in caelestibus per ecclesiam multiformis sapientia Dei
EPH|3|11|secundum praefinitionem saeculorum quam fecit in Christo Iesu Domino nostro
EPH|3|12|in quo habemus fiduciam et accessum in confidentia per fidem eius
EPH|3|13|propter quod peto ne deficiatis in tribulationibus meis pro vobis quae est gloria vestra
EPH|3|14|huius rei gratia flecto genua mea ad Patrem Domini nostri Iesu Christi
EPH|3|15|ex quo omnis paternitas in caelis et in terra nominatur
EPH|3|16|ut det vobis secundum divitias gloriae suae virtute corroborari per Spiritum eius in interiore homine
EPH|3|17|habitare Christum per fidem in cordibus vestris in caritate radicati et fundati
EPH|3|18|ut possitis conprehendere cum omnibus sanctis quae sit latitudo et longitudo et sublimitas et profundum
EPH|3|19|scire etiam supereminentem scientiae caritatem Christi ut impleamini in omnem plenitudinem Dei
EPH|3|20|ei autem qui potens est omnia facere superabundanter quam petimus aut intellegimus secundum virtutem quae operatur in nobis
EPH|3|21|ipsi gloria in ecclesia et in Christo Iesu in omnes generationes saeculi saeculorum amen
EPH|4|1|obsecro itaque vos ego vinctus in Domino ut digne ambuletis vocatione qua vocati estis
EPH|4|2|cum omni humilitate et mansuetudine cum patientia subportantes invicem in caritate
EPH|4|3|solliciti servare unitatem spiritus in vinculo pacis
EPH|4|4|unum corpus et unus spiritus sicut vocati estis in una spe vocationis vestrae
EPH|4|5|unus Dominus una fides unum baptisma
EPH|4|6|unus Deus et Pater omnium qui super omnes et per omnia et in omnibus nobis
EPH|4|7|unicuique autem nostrum data est gratia secundum mensuram donationis Christi
EPH|4|8|propter quod dicit ascendens in altum captivam duxit captivitatem dedit dona hominibus
EPH|4|9|quod autem ascendit quid est nisi quia et descendit primum in inferiores partes terrae
EPH|4|10|qui descendit ipse est et qui ascendit super omnes caelos ut impleret omnia
EPH|4|11|et ipse dedit quosdam quidem apostolos quosdam autem prophetas alios vero evangelistas alios autem pastores et doctores
EPH|4|12|ad consummationem sanctorum in opus ministerii in aedificationem corporis Christi
EPH|4|13|donec occurramus omnes in unitatem fidei et agnitionis Filii Dei in virum perfectum in mensuram aetatis plenitudinis Christi
EPH|4|14|ut iam non simus parvuli fluctuantes et circumferamur omni vento doctrinae in nequitia hominum in astutia ad circumventionem erroris
EPH|4|15|veritatem autem facientes in caritate crescamus in illo per omnia qui est caput Christus
EPH|4|16|ex quo totum corpus conpactum et conexum per omnem iuncturam subministrationis secundum operationem in mensuram uniuscuiusque membri augmentum corporis facit in aedificationem sui in caritate
EPH|4|17|hoc igitur dico et testificor in Domino ut iam non ambuletis sicut gentes ambulant in vanitate sensus sui
EPH|4|18|tenebris obscuratum habentes intellectum alienati a vita Dei per ignorantiam quae est in illis propter caecitatem cordis ipsorum
EPH|4|19|qui desperantes semet ipsos tradiderunt inpudicitiae in operationem inmunditiae omnis in avaritia
EPH|4|20|vos autem non ita didicistis Christum
EPH|4|21|si tamen illum audistis et in ipso edocti estis sicut est veritas in Iesu
EPH|4|22|deponere vos secundum pristinam conversationem veterem hominem qui corrumpitur secundum desideria erroris
EPH|4|23|renovamini autem spiritu mentis vestrae
EPH|4|24|et induite novum hominem qui secundum Deum creatus est in iustitia et sanctitate veritatis
EPH|4|25|propter quod deponentes mendacium loquimini veritatem unusquisque cum proximo suo quoniam sumus invicem membra
EPH|4|26|irascimini et nolite peccare sol non occidat super iracundiam vestram
EPH|4|27|nolite locum dare diabolo
EPH|4|28|qui furabatur iam non furetur magis autem laboret operando manibus quod bonum est ut habeat unde tribuat necessitatem patienti
EPH|4|29|omnis sermo malus ex ore vestro non procedat sed si quis bonus ad aedificationem oportunitatis ut det gratiam audientibus
EPH|4|30|et nolite contristare Spiritum Sanctum Dei in quo signati estis in die redemptionis
EPH|4|31|omnis amaritudo et ira et indignatio et clamor et blasphemia tollatur a vobis cum omni malitia
EPH|4|32|estote autem invicem benigni misericordes donantes invicem sicut et Deus in Christo donavit nobis
EPH|5|1|estote ergo imitatores Dei sicut filii carissimi
EPH|5|2|et ambulate in dilectione sicut et Christus dilexit nos et tradidit se ipsum pro nobis oblationem et hostiam Deo in odorem suavitatis
EPH|5|3|fornicatio autem et omnis inmunditia aut avaritia nec nominetur in vobis sicut decet sanctos
EPH|5|4|aut turpitudo aut stultiloquium aut scurrilitas quae ad rem non pertinent sed magis gratiarum actio
EPH|5|5|hoc enim scitote intellegentes quod omnis fornicator aut inmundus aut avarus quod est idolorum servitus non habet hereditatem in regno Christi et Dei
EPH|5|6|nemo vos seducat inanibus verbis propter haec enim venit ira Dei in filios diffidentiae
EPH|5|7|nolite ergo effici participes eorum
EPH|5|8|eratis enim aliquando tenebrae nunc autem lux in Domino ut filii lucis ambulate
EPH|5|9|fructus enim lucis est in omni bonitate et iustitia et veritate
EPH|5|10|probantes quid sit beneplacitum Deo
EPH|5|11|et nolite communicare operibus infructuosis tenebrarum magis autem et redarguite
EPH|5|12|quae enim in occulto fiunt ab ipsis turpe est et dicere
EPH|5|13|omnia autem quae arguuntur a lumine manifestantur omne enim quod manifestatur lumen est
EPH|5|14|propter quod dicit surge qui dormis et exsurge a mortuis et inluminabit tibi Christus
EPH|5|15|videte itaque fratres quomodo caute ambuletis non quasi insipientes sed ut sapientes
EPH|5|16|redimentes tempus quoniam dies mali sunt
EPH|5|17|propterea nolite fieri inprudentes sed intellegentes quae sit voluntas Domini
EPH|5|18|et nolite inebriari vino in quo est luxuria sed implemini Spiritu
EPH|5|19|loquentes vobismet ipsis in psalmis et hymnis et canticis spiritalibus cantantes et psallentes in cordibus vestris Domino
EPH|5|20|gratias agentes semper pro omnibus in nomine Domini nostri Iesu Christi Deo et Patri
EPH|5|21|subiecti invicem in timore Christi
EPH|5|22|mulieres viris suis subditae sint sicut Domino
EPH|5|23|quoniam vir caput est mulieris sicut Christus caput est ecclesiae ipse salvator corporis
EPH|5|24|sed ut ecclesia subiecta est Christo ita et mulieres viris suis in omnibus
EPH|5|25|viri diligite uxores sicut et Christus dilexit ecclesiam et se ipsum tradidit pro ea
EPH|5|26|ut illam sanctificaret mundans lavacro aquae in verbo
EPH|5|27|ut exhiberet ipse sibi gloriosam ecclesiam non habentem maculam aut rugam aut aliquid eiusmodi sed ut sit sancta et inmaculata
EPH|5|28|ita et viri debent diligere uxores suas ut corpora sua qui suam uxorem diligit se ipsum diligit
EPH|5|29|nemo enim umquam carnem suam odio habuit sed nutrit et fovet eam sicut et Christus ecclesiam
EPH|5|30|quia membra sumus corporis eius de carne eius et de ossibus eius
EPH|5|31|propter hoc relinquet homo patrem et matrem suam et adherebit uxori suae et erunt duo in carne una
EPH|5|32|sacramentum hoc magnum est ego autem dico in Christo et in ecclesia
EPH|5|33|verumtamen et vos singuli unusquisque suam uxorem sicut se ipsum diligat uxor autem ut timeat virum
EPH|6|1|filii oboedite parentibus vestris in Domino hoc enim est iustum
EPH|6|2|honora patrem tuum et matrem quod est mandatum primum in promissione
EPH|6|3|ut bene sit tibi et sis longevus super terram
EPH|6|4|et patres nolite ad iracundiam provocare filios vestros sed educate illos in disciplina et correptione Domini
EPH|6|5|servi oboedite dominis carnalibus cum timore et tremore in simplicitate cordis vestri sicut Christo
EPH|6|6|non ad oculum servientes quasi hominibus placentes sed ut servi Christi facientes voluntatem Dei ex animo
EPH|6|7|cum bona voluntate servientes sicut Domino et non hominibus
EPH|6|8|scientes quoniam unusquisque quodcumque fecerit bonum hoc percipiet a Domino sive servus sive liber
EPH|6|9|et domini eadem facite illis remittentes minas scientes quia et illorum et vester Dominus est in caelis et personarum acceptio non est apud eum
EPH|6|10|de cetero fratres confortamini in Domino et in potentia virtutis eius
EPH|6|11|induite vos arma Dei ut possitis stare adversus insidias diaboli
EPH|6|12|quia non est nobis conluctatio adversus carnem et sanguinem sed adversus principes et potestates adversus mundi rectores tenebrarum harum contra spiritalia nequitiae in caelestibus
EPH|6|13|propterea accipite armaturam Dei ut possitis resistere in die malo et omnibus perfectis stare
EPH|6|14|state ergo succincti lumbos vestros in veritate et induti loricam iustitiae
EPH|6|15|et calciati pedes in praeparatione evangelii pacis
EPH|6|16|in omnibus sumentes scutum fidei in quo possitis omnia tela nequissimi ignea extinguere
EPH|6|17|et galeam salutis adsumite et gladium Spiritus quod est verbum Dei
EPH|6|18|per omnem orationem et obsecrationem orantes omni tempore in Spiritu et in ipso vigilantes in omni instantia et obsecratione pro omnibus sanctis
EPH|6|19|et pro me ut detur mihi sermo in apertione oris mei cum fiducia notum facere mysterium evangelii
EPH|6|20|pro quo legatione fungor in catena ita ut in ipso audeam prout oportet me loqui
EPH|6|21|ut autem et vos sciatis quae circa me sunt quid agam omnia nota vobis faciet Tychicus carissimus frater et fidelis minister in Domino
EPH|6|22|quem misi ad vos in hoc ipsum ut cognoscatis quae circa nos sunt et consoletur corda vestra
EPH|6|23|pax fratribus et caritas cum fide a Deo Patre et Domino Iesu Christo
EPH|6|24|gratia cum omnibus qui diligunt Dominum nostrum Iesum Christum in incorruptione
PHIL|1|1|Paulus et Timotheus servi Iesu Christi omnibus sanctis in Christo Iesu qui sunt Philippis cum episcopis et diaconis
PHIL|1|2|gratia vobis et pax a Deo Patre nostro et Domino Iesu Christo
PHIL|1|3|gratias ago Deo meo in omni memoria vestri
PHIL|1|4|semper in cunctis orationibus meis pro omnibus vobis cum gaudio deprecationem faciens
PHIL|1|5|super communicatione vestra in evangelio a prima die usque nunc
PHIL|1|6|confidens hoc ipsum quia qui coepit in vobis opus bonum perficiet usque in diem Christi Iesu
PHIL|1|7|sicut est mihi iustum hoc sentire pro omnibus vobis eo quod habeam in corde vos et in vinculis meis et in defensione et confirmatione evangelii socios gaudii mei omnes vos esse
PHIL|1|8|testis enim mihi est Deus quomodo cupiam omnes vos in visceribus Christi Iesu
PHIL|1|9|et hoc oro ut caritas vestra magis ac magis abundet in scientia et omni sensu
PHIL|1|10|ut probetis potiora ut sitis sinceres et sine offensa in diem Christi
PHIL|1|11|repleti fructu iustitiae per Christum Iesum in gloriam et laudem Dei
PHIL|1|12|scire autem vos volo fratres quia quae circa me sunt magis ad profectum venerunt evangelii
PHIL|1|13|ita ut vincula mea manifesta fierent in Christo in omni praetorio et in ceteris omnibus
PHIL|1|14|et plures e fratribus in Domino confidentes vinculis meis abundantius audere sine timore verbum Dei loqui
PHIL|1|15|quidam quidem et propter invidiam et contentionem quidam autem et propter bonam voluntatem Christum praedicant
PHIL|1|16|quidam ex caritate scientes quoniam in defensionem evangelii positus sum
PHIL|1|17|quidam autem ex contentione Christum adnuntiant non sincere existimantes pressuram se suscitare vinculis meis
PHIL|1|18|quid enim dum omni modo sive per occasionem sive per veritatem Christus adnuntiatur et in hoc gaudeo sed et gaudebo
PHIL|1|19|scio enim quia hoc mihi proveniet in salutem per vestram orationem et subministrationem Spiritus Iesu Christi
PHIL|1|20|secundum expectationem et spem meam quia in nullo confundar sed in omni fiducia sicut semper et nunc magnificabitur Christus in corpore meo sive per vitam sive per mortem
PHIL|1|21|mihi enim vivere Christus est et mori lucrum
PHIL|1|22|quod si vivere in carne hic mihi fructus operis est et quid eligam ignoro
PHIL|1|23|coartor autem e duobus desiderium habens dissolvi et cum Christo esse multo magis melius
PHIL|1|24|permanere autem in carne magis necessarium est propter vos
PHIL|1|25|et hoc confidens scio quia manebo et permanebo omnibus vobis ad profectum vestrum et gaudium fidei
PHIL|1|26|ut gratulatio vestra abundet in Christo Iesu in me per meum adventum iterum ad vos
PHIL|1|27|tantum digne evangelio Christi conversamini ut sive cum venero et videro vos sive absens audiam de vobis quia stetistis uno spiritu unianimes conlaborantes fide evangelii
PHIL|1|28|et in nullo terreamini ab adversariis quae est illis causa perditionis vobis autem salutis et hoc a Deo
PHIL|1|29|quia vobis donatum est pro Christo non solum ut in eum credatis sed ut etiam pro illo patiamini
PHIL|1|30|eundem certamen habentes qualem et vidistis in me et nunc audistis de me
PHIL|2|1|si qua ergo consolatio in Christo si quod solacium caritatis si qua societas spiritus si quid viscera et miserationes
PHIL|2|2|implete gaudium meum ut idem sapiatis eandem caritatem habentes unianimes id ipsum sentientes
PHIL|2|3|nihil per contentionem neque per inanem gloriam sed in humilitate superiores sibi invicem arbitrantes
PHIL|2|4|non quae sua sunt singuli considerantes sed et ea quae aliorum
PHIL|2|5|hoc enim sentite in vobis quod et in Christo Iesu
PHIL|2|6|qui cum in forma Dei esset non rapinam arbitratus est esse se aequalem Deo
PHIL|2|7|sed semet ipsum exinanivit formam servi accipiens in similitudinem hominum factus et habitu inventus ut homo
PHIL|2|8|humiliavit semet ipsum factus oboediens usque ad mortem mortem autem crucis
PHIL|2|9|propter quod et Deus illum exaltavit et donavit illi nomen super omne nomen
PHIL|2|10|ut in nomine Iesu omne genu flectat caelestium et terrestrium et infernorum
PHIL|2|11|et omnis lingua confiteatur quia Dominus Iesus Christus in gloria est Dei Patris
PHIL|2|12|itaque carissimi mei sicut semper oboedistis non ut in praesentia mei tantum sed multo magis nunc in absentia mea cum metu et tremore vestram salutem operamini
PHIL|2|13|Deus est enim qui operatur in vobis et velle et perficere pro bona voluntate
PHIL|2|14|omnia autem facite sine murmurationibus et haesitationibus
PHIL|2|15|ut sitis sine querella et simplices filii Dei sine reprehensione in medio nationis pravae et perversae inter quos lucetis sicut luminaria in mundo
PHIL|2|16|verbum vitae continentes ad gloriam meam in die Christi quia non in vacuum cucurri neque in vacuum laboravi
PHIL|2|17|sed et si immolor supra sacrificium et obsequium fidei vestrae gaudeo et congratulor omnibus vobis
PHIL|2|18|id ipsum autem et vos gaudete et congratulamini mihi
PHIL|2|19|spero autem in Domino Iesu Timotheum cito me mittere ad vos ut et ego bono animo sim cognitis quae circa vos sunt
PHIL|2|20|neminem enim habeo tam unianimem qui sincera affectione pro vobis sollicitus sit
PHIL|2|21|omnes enim sua quaerunt non quae sunt Christi Iesu
PHIL|2|22|experimentum autem eius cognoscite quoniam sicut patri filius mecum servivit in evangelium
PHIL|2|23|hunc igitur spero me mittere mox ut videro quae circa me sunt
PHIL|2|24|confido autem in Domino quoniam et ipse veniam ad vos cito
PHIL|2|25|necessarium autem existimavi Epafroditum fratrem et cooperatorem et commilitonem meum vestrum autem apostolum et ministrum necessitatis meae mittere ad vos
PHIL|2|26|quoniam quidem omnes vos desiderabat et maestus erat propterea quod audieratis illum infirmatum
PHIL|2|27|nam et infirmatus est usque ad mortem sed Deus misertus est eius non solum autem eius verum etiam et mei ne tristitiam super tristitiam haberem
PHIL|2|28|festinantius ergo misi illum ut viso eo iterum gaudeatis et ego sine tristitia sim
PHIL|2|29|excipite itaque illum cum omni gaudio in Domino et eiusmodi cum honore habetote
PHIL|2|30|quoniam propter opus Christi usque ad mortem accessit tradens animam suam ut impleret id quod ex vobis deerat erga meum obsequium
PHIL|3|1|de cetero fratres mei gaudete in Domino eadem vobis scribere mihi quidem non pigrum vobis autem necessarium
PHIL|3|2|videte canes videte malos operarios videte concisionem
PHIL|3|3|nos enim sumus circumcisio qui spiritu Deo servimus et gloriamur in Christo Iesu et non in carne fiduciam habentes
PHIL|3|4|quamquam ego habeam confidentiam et in carne si quis alius videtur confidere in carne ego magis
PHIL|3|5|circumcisus octava die ex genere Israhel de tribu Beniamin Hebraeus ex Hebraeis secundum legem Pharisaeus
PHIL|3|6|secundum aemulationem persequens ecclesiam Dei secundum iustitiam quae in lege est conversatus sine querella
PHIL|3|7|sed quae mihi fuerunt lucra haec arbitratus sum propter Christum detrimenta
PHIL|3|8|verumtamen existimo omnia detrimentum esse propter eminentem scientiam Iesu Christi Domini mei propter quem omnia detrimentum feci et arbitror ut stercora ut Christum lucri faciam
PHIL|3|9|et inveniar in illo non habens meam iustitiam quae ex lege est sed illam quae ex fide est Christi quae ex Deo est iustitia in fide
PHIL|3|10|ad agnoscendum illum et virtutem resurrectionis eius et societatem passionum illius configuratus morti eius
PHIL|3|11|si quo modo occurram ad resurrectionem quae est ex mortuis
PHIL|3|12|non quod iam acceperim aut iam perfectus sim sequor autem si conprehendam in quo et conprehensus sum a Christo Iesu
PHIL|3|13|fratres ego me non arbitror conprehendisse unum autem quae quidem retro sunt obliviscens ad ea vero quae sunt in priora extendens me
PHIL|3|14|ad destinatum persequor ad bravium supernae vocationis Dei in Christo Iesu
PHIL|3|15|quicumque ergo perfecti hoc sentiamus et si quid aliter sapitis et hoc vobis Deus revelabit
PHIL|3|16|verumtamen ad quod pervenimus ut idem sapiamus et in eadem permaneamus regula
PHIL|3|17|imitatores mei estote fratres et observate eos qui ita ambulant sicut habetis formam nos
PHIL|3|18|multi enim ambulant quos saepe dicebam vobis nunc autem et flens dico inimicos crucis Christi
PHIL|3|19|quorum finis interitus quorum deus venter et gloria in confusione ipsorum qui terrena sapiunt
PHIL|3|20|nostra autem conversatio in caelis est unde etiam salvatorem expectamus Dominum Iesum Christum
PHIL|3|21|qui reformabit corpus humilitatis nostrae configuratum corpori claritatis suae secundum operationem qua possit etiam subicere sibi omnia
PHIL|4|1|itaque fratres mei carissimi et desiderantissimi gaudium meum et corona mea sic state in Domino carissimi
PHIL|4|2|Euhodiam rogo et Syntychen deprecor id ipsum sapere in Domino
PHIL|4|3|etiam rogo et te germane conpar adiuva illas quae mecum laboraverunt in evangelio cum Clemente et ceteris adiutoribus meis quorum nomina sunt in libro vitae
PHIL|4|4|gaudete in Domino semper iterum dico gaudete
PHIL|4|5|modestia vestra nota sit omnibus hominibus Dominus prope
PHIL|4|6|nihil solliciti sitis sed in omni oratione et obsecratione cum gratiarum actione petitiones vestrae innotescant apud Deum
PHIL|4|7|et pax Dei quae exsuperat omnem sensum custodiat corda vestra et intellegentias vestras in Christo Iesu
PHIL|4|8|de cetero fratres quaecumque sunt vera quaecumque pudica quaecumque iusta quaecumque sancta quaecumque amabilia quaecumque bonae famae si qua virtus si qua laus haec cogitate
PHIL|4|9|quae et didicistis et accepistis et audistis et vidistis in me haec agite et Deus pacis erit vobiscum
PHIL|4|10|gavisus sum autem in Domino vehementer quoniam tandem aliquando refloruistis pro me sentire sicut et sentiebatis occupati autem eratis
PHIL|4|11|non quasi propter penuriam dico ego enim didici in quibus sum sufficiens esse
PHIL|4|12|scio et humiliari scio et abundare ubique et in omnibus institutus sum et satiari et esurire et abundare et penuriam pati
PHIL|4|13|omnia possum in eo qui me confortat
PHIL|4|14|verumtamen bene fecistis communicantes tribulationi meae
PHIL|4|15|scitis autem et vos Philippenses quod in principio evangelii quando profectus sum a Macedonia nulla mihi ecclesia communicavit in ratione dati et accepti nisi vos soli
PHIL|4|16|quia et Thessalonicam et semel et bis in usum mihi misistis
PHIL|4|17|non quia quaero datum sed requiro fructum abundantem in rationem vestram
PHIL|4|18|habeo autem omnia et abundo repletus sum acceptis ab Epafrodito quae misistis odorem suavitatis hostiam acceptam placentem Deo
PHIL|4|19|Deus autem meus impleat omne desiderium vestrum secundum divitias suas in gloria in Christo Iesu
PHIL|4|20|Deo autem et Patri nostro gloria in saecula saeculorum amen
PHIL|4|21|salutate omnem sanctum in Christo Iesu salutant vos qui mecum sunt fratres
PHIL|4|22|salutant vos omnes sancti maxime autem qui de Caesaris domo sunt
PHIL|4|23|gratia Domini Iesu Christi cum spiritu vestro amen
COL|1|1|Paulus apostolus Christi Iesu per voluntatem Dei et Timotheus frater
COL|1|2|his qui sunt Colossis sanctis et fidelibus fratribus in Christo Iesu gratia vobis et pax a Deo Patre nostro
COL|1|3|gratias agimus Deo et Patri Domini nostri Iesu Christi semper pro vobis orantes
COL|1|4|audientes fidem vestram in Christo Iesu et dilectionem quam habetis in sanctos omnes
COL|1|5|propter spem quae reposita est vobis in caelis quam audistis in verbo veritatis evangelii
COL|1|6|quod pervenit ad vos sicut et in universo mundo est et fructificat et crescit sicut in vobis ex ea die qua audistis et cognovistis gratiam Dei in veritate
COL|1|7|sicut didicistis ab Epaphra carissimo conservo nostro qui est fidelis pro vobis minister Christi Iesu
COL|1|8|qui etiam manifestavit nobis dilectionem vestram in Spiritu
COL|1|9|ideo et nos ex qua die audivimus non cessamus pro vobis orantes et postulantes ut impleamini agnitione voluntatis eius in omni sapientia et intellectu spiritali
COL|1|10|ut ambuletis digne Deo per omnia placentes in omni opere bono fructificantes et crescentes in scientia Dei
COL|1|11|in omni virtute confortati secundum potentiam claritatis eius in omni patientia et longanimitate cum gaudio
COL|1|12|gratias agentes Patri qui dignos nos fecit in partem sortis sanctorum in lumine
COL|1|13|qui eripuit nos de potestate tenebrarum et transtulit in regnum Filii dilectionis suae
COL|1|14|in quo habemus redemptionem remissionem peccatorum
COL|1|15|qui est imago Dei invisibilis primogenitus omnis creaturae
COL|1|16|quia in ipso condita sunt universa in caelis et in terra visibilia et invisibilia sive throni sive dominationes sive principatus sive potestates omnia per ipsum et in ipso creata sunt
COL|1|17|et ipse est ante omnes et omnia in ipso constant
COL|1|18|et ipse est caput corporis ecclesiae qui est principium primogenitus ex mortuis ut sit in omnibus ipse primatum tenens
COL|1|19|quia in ipso conplacuit omnem plenitudinem habitare
COL|1|20|et per eum reconciliare omnia in ipsum pacificans per sanguinem crucis eius sive quae in terris sive quae in caelis sunt
COL|1|21|et vos cum essetis aliquando alienati et inimici sensu in operibus malis
COL|1|22|nunc autem reconciliavit in corpore carnis eius per mortem exhibere vos sanctos et inmaculatos et inreprehensibiles coram ipso
COL|1|23|si tamen permanetis in fide fundati et stabiles et inmobiles ab spe evangelii quod audistis quod praedicatum est in universa creatura quae sub caelo est cuius factus sum ego Paulus minister
COL|1|24|qui nunc gaudeo in passionibus pro vobis et adimpleo ea quae desunt passionum Christi in carne mea pro corpore eius quod est ecclesia
COL|1|25|cuius factus sum ego minister secundum dispensationem Dei quae data est mihi in vos ut impleam verbum Dei
COL|1|26|mysterium quod absconditum fuit a saeculis et generationibus nunc autem manifestatum est sanctis eius
COL|1|27|quibus voluit Deus notas facere divitias gloriae sacramenti huius in gentibus quod est Christus in vobis spes gloriae
COL|1|28|quem nos adnuntiamus corripientes omnem hominem et docentes omnem hominem in omni sapientia ut exhibeamus omnem hominem perfectum in Christo Iesu
COL|1|29|in quo et laboro certando secundum operationem eius quam operatur in me in virtute
COL|2|1|volo enim vos scire qualem sollicitudinem habeam pro vobis et pro his qui sunt Laodiciae et quicumque non viderunt faciem meam in carne
COL|2|2|ut consolentur corda ipsorum instructi in caritate et in omnes divitias plenitudinis intellectus in agnitionem mysterii Dei Patris Christi Iesu
COL|2|3|in quo sunt omnes thesauri sapientiae et scientiae absconditi
COL|2|4|hoc autem dico ut nemo vos decipiat in subtilitate sermonum
COL|2|5|nam et si corpore absens sum sed spiritu vobiscum sum gaudens et videns ordinem vestrum et firmamentum eius quae in Christo est fidei vestrae
COL|2|6|sicut ergo accepistis Christum Iesum Dominum in ipso ambulate
COL|2|7|radicati et superaedificati in ipso et confirmati fide sicut et didicistis abundantes in gratiarum actione
COL|2|8|videte ne quis vos decipiat per philosophiam et inanem fallaciam secundum traditionem hominum secundum elementa mundi et non secundum Christum
COL|2|9|quia in ipso inhabitat omnis plenitudo divinitatis corporaliter
COL|2|10|et estis in illo repleti qui est caput omnis principatus et potestatis
COL|2|11|in quo et circumcisi estis circumcisione non manufacta in expoliatione corporis carnis in circumcisione Christi
COL|2|12|consepulti ei in baptismo in quo et resurrexistis per fidem operationis Dei qui suscitavit illum a mortuis
COL|2|13|et vos cum mortui essetis in delictis et praeputio carnis vestrae convivificavit cum illo donans vobis omnia delicta
COL|2|14|delens quod adversum nos erat chirografum decretis quod erat contrarium nobis et ipsum tulit de medio adfigens illud cruci
COL|2|15|expolians principatus et potestates traduxit palam triumphans illos in semet ipso
COL|2|16|nemo ergo vos iudicet in cibo aut in potu aut in parte diei festi aut neomeniae aut sabbatorum
COL|2|17|quae sunt umbra futurorum corpus autem Christi
COL|2|18|nemo vos seducat volens in humilitate et religione angelorum quae non vidit ambulans frustra inflatus sensu carnis suae
COL|2|19|et non tenens caput ex quo totum corpus per nexus et coniunctiones subministratum et constructum crescit in augmentum Dei
COL|2|20|si mortui estis cum Christo ab elementis mundi quid adhuc tamquam viventes in mundo decernitis
COL|2|21|ne tetigeris neque gustaveris neque contrectaveris
COL|2|22|quae sunt omnia in interitu ipso usu secundum praecepta et doctrinas hominum
COL|2|23|quae sunt rationem quidem habentia sapientiae in superstitione et humilitate et ad non parcendum corpori non in honore aliquo ad saturitatem carnis
COL|3|1|igitur si conresurrexistis Christo quae sursum sunt quaerite ubi Christus est in dextera Dei sedens
COL|3|2|quae sursum sunt sapite non quae supra terram
COL|3|3|mortui enim estis et vita vestra abscondita est cum Christo in Deo
COL|3|4|cum Christus apparuerit vita vestra tunc et vos apparebitis cum ipso in gloria
COL|3|5|mortificate ergo membra vestra quae sunt super terram fornicationem inmunditiam libidinem concupiscentiam malam et avaritiam quae est simulacrorum servitus
COL|3|6|propter quae venit ira Dei super filios incredulitatis
COL|3|7|in quibus et vos ambulastis aliquando cum viveretis in illis
COL|3|8|nunc autem deponite et vos omnia iram indignationem malitiam blasphemiam turpem sermonem de ore vestro
COL|3|9|nolite mentiri invicem expoliantes vos veterem hominem cum actibus eius
COL|3|10|et induentes novum eum qui renovatur in agnitionem secundum imaginem eius qui creavit eum
COL|3|11|ubi non est gentilis et Iudaeus circumcisio et praeputium barbarus et Scytha servus et liber sed omnia et in omnibus Christus
COL|3|12|induite vos ergo sicut electi Dei sancti et dilecti viscera misericordiae benignitatem humilitatem modestiam patientiam
COL|3|13|subportantes invicem et donantes vobis ipsis si quis adversus aliquem habet querellam sicut et Dominus donavit vobis ita et vos
COL|3|14|super omnia autem haec caritatem quod est vinculum perfectionis
COL|3|15|et pax Christi exultet in cordibus vestris in qua et vocati estis in uno corpore et grati estote
COL|3|16|verbum Christi habitet in vobis abundanter in omni sapientia docentes et commonentes vosmet ipsos psalmis hymnis canticis spiritalibus in gratia cantantes in cordibus vestris Deo
COL|3|17|omne quodcumque facitis in verbo aut in opere omnia in nomine Domini Iesu gratias agentes Deo et Patri per ipsum
COL|3|18|mulieres subditae estote viris sicut oportet in Domino
COL|3|19|viri diligite uxores et nolite amari esse ad illas
COL|3|20|filii oboedite parentibus per omnia hoc enim placitum est in Domino
COL|3|21|patres nolite ad indignationem provocare filios vestros ut non pusillo animo fiant
COL|3|22|servi oboedite per omnia dominis carnalibus non ad oculum servientes quasi hominibus placentes sed in simplicitate cordis timentes Dominum
COL|3|23|quodcumque facitis ex animo operamini sicut Domino et non hominibus
COL|3|24|scientes quod a Domino accipietis retributionem hereditatis Domino Christo servite
COL|3|25|qui enim iniuriam facit recipiet id quod inique gessit et non est personarum acceptio
COL|4|1|domini quod iustum est et aequum servis praestate scientes quoniam et vos Dominum habetis in caelo
COL|4|2|orationi instate vigilantes in ea in gratiarum actione
COL|4|3|orantes simul et pro nobis ut Deus aperiat nobis ostium sermonis ad loquendum mysterium Christi propter quod etiam vinctus sum
COL|4|4|ut manifestem illud ita ut oportet me loqui
COL|4|5|in sapientia ambulate ad eos qui foris sunt tempus redimentes
COL|4|6|sermo vester semper in gratia sale sit conditus ut sciatis quomodo oporteat vos unicuique respondere
COL|4|7|quae circa me sunt omnia vobis nota faciet Tychicus carissimus frater et fidelis minister et conservus in Domino
COL|4|8|quem misi ad vos ad hoc ipsum ut cognoscat quae circa vos sunt et consoletur corda vestra
COL|4|9|cum Onesimo carissimo et fideli fratre qui est ex vobis omnia quae hic aguntur nota facient vobis
COL|4|10|salutat vos Aristarchus concaptivus meus et Marcus consobrinus Barnabae de quo accepistis mandata si venerit ad vos excipite illum
COL|4|11|et Iesus qui dicitur Iustus qui sunt ex circumcisione hii soli sunt adiutores in regno Dei qui mihi fuerunt solacio
COL|4|12|salutat vos Epaphras qui ex vobis est servus Christi Iesu semper sollicitus pro vobis in orationibus ut stetis perfecti et pleni in omni voluntate Dei
COL|4|13|testimonium enim illi perhibeo quod habet multum laborem pro vobis et pro his qui sunt Laodiciae et qui Hierapoli
COL|4|14|salutat vos Lucas medicus carissimus et Demas
COL|4|15|salutate fratres qui sunt Laodiciae et Nympham et quae in domo eius est ecclesiam
COL|4|16|et cum lecta fuerit apud vos epistula facite ut et in Laodicensium ecclesia legatur et eam quae Laodicensium est vos legatis
COL|4|17|et dicite Archippo vide ministerium quod accepisti in Domino ut illud impleas
COL|4|18|salutatio mea manu Pauli memores estote vinculorum meorum gratia vobiscum amen
1THESS|1|1|Paulus et Silvanus et Timotheus ecclesiae Thessalonicensium in Deo Patre et Domino Iesu Christo gratia vobis et pax
1THESS|1|2|gratias agimus Deo semper pro omnibus vobis memoriam facientes in orationibus nostris sine intermissione
1THESS|1|3|memores operis fidei vestrae et laboris et caritatis et sustinentiae spei Domini nostri Iesu Christi ante Deum et Patrem nostrum
1THESS|1|4|scientes fratres dilecti a Deo electionem vestram
1THESS|1|5|quia evangelium nostrum non fuit ad vos in sermone tantum sed et in virtute et in Spiritu Sancto et in plenitudine multa sicut scitis quales fuerimus vobis propter vos
1THESS|1|6|et vos imitatores nostri facti estis et Domini excipientes verbum in tribulatione multa cum gaudio Spiritus Sancti
1THESS|1|7|ita ut facti sitis forma omnibus credentibus in Macedonia et in Achaia
1THESS|1|8|a vobis enim diffamatus est sermo Domini non solum in Macedonia et in Achaia sed in omni loco fides vestra quae est ad Deum profecta est ita ut non sit nobis necesse quicquam loqui
1THESS|1|9|ipsi enim de nobis adnuntiant qualem introitum habuerimus ad vos et quomodo conversi estis ad Deum a simulacris servire Deo vivo et vero
1THESS|1|10|et expectare Filium eius de caelis quem suscitavit ex mortuis Iesum qui eripuit nos ab ira ventura
1THESS|2|1|nam ipsi scitis fratres introitum nostrum ad vos quia non inanis fuit
1THESS|2|2|sed ante passi et contumeliis affecti sicut scitis in Philippis fiduciam habuimus in Deo nostro loqui ad vos evangelium Dei in multa sollicitudine
1THESS|2|3|exhortatio enim nostra non de errore neque de inmunditia neque in dolo
1THESS|2|4|sed sicut probati sumus a Deo ut crederetur nobis evangelium ita loquimur non quasi hominibus placentes sed Deo qui probat corda nostra
1THESS|2|5|neque enim aliquando fuimus in sermone adulationis sicut scitis neque in occasione avaritiae Deus testis est
1THESS|2|6|nec quaerentes ab hominibus gloriam neque a vobis neque ab aliis
1THESS|2|7|cum possimus oneri esse ut Christi apostoli sed facti sumus lenes in medio vestrum tamquam si nutrix foveat filios suos
1THESS|2|8|ita desiderantes vos cupide volebamus tradere vobis non solum evangelium Dei sed etiam animas nostras quoniam carissimi nobis facti estis
1THESS|2|9|memores enim estis fratres laborem nostrum et fatigationem nocte et die operantes ne quem vestrum gravaremus praedicavimus in vobis evangelium Dei
1THESS|2|10|vos testes estis et Deus quam sancte et iuste et sine querella vobis qui credidistis fuimus
1THESS|2|11|sicut scitis qualiter unumquemque vestrum tamquam pater filios suos
1THESS|2|12|deprecantes vos et consolantes testificati sumus ut ambularetis digne Deo qui vocavit vos in suum regnum et gloriam
1THESS|2|13|ideo et nos gratias agimus Deo sine intermissione quoniam cum accepissetis a nobis verbum auditus Dei accepistis non ut verbum hominum sed sicut est vere verbum Dei qui operatur in vobis qui credidistis
1THESS|2|14|vos enim imitatores facti estis fratres ecclesiarum Dei quae sunt in Iudaea in Christo Iesu quia eadem passi estis et vos a contribulibus vestris sicut et ipsi a Iudaeis
1THESS|2|15|qui et Dominum occiderunt Iesum et prophetas et nos persecuti sunt et Deo non placent et omnibus hominibus adversantur
1THESS|2|16|prohibentes nos gentibus loqui ut salvae fiant ut impleant peccata sua semper praevenit autem ira Dei super illos usque in finem
1THESS|2|17|nos autem fratres desolati a vobis ad tempus horae aspectu non corde abundantius festinavimus faciem vestram videre cum multo desiderio
1THESS|2|18|quoniam voluimus venire ad vos ego quidem Paulus et semel et iterum et inpedivit nos Satanas
1THESS|2|19|quae est enim nostra spes aut gaudium aut corona gloriae nonne vos ante Dominum nostrum Iesum estis in adventu eius
1THESS|2|20|vos enim estis gloria nostra et gaudium
1THESS|3|1|propter quod non sustinentes amplius placuit nobis remanere Athenis solis
1THESS|3|2|et misimus Timotheum fratrem nostrum et ministrum Dei in evangelio Christi ad confirmandos vos et exhortandos pro fide vestra
1THESS|3|3|ut nemo moveatur in tribulationibus istis ipsi enim scitis quod in hoc positi sumus
1THESS|3|4|nam et cum apud vos essemus praedicebamus vobis passuros nos tribulationes sicut et factum est et scitis
1THESS|3|5|propterea et ego amplius non sustinens misi ad cognoscendam fidem vestram ne forte temptaverit vos is qui temptat et inanis fiat labor noster
1THESS|3|6|nunc autem veniente Timotheo ad nos a vobis et adnuntiante nobis fidem et caritatem vestram et quia memoriam nostri habetis bonam semper desiderantes nos videre sicut nos quoque vos
1THESS|3|7|ideo consolati sumus fratres in vobis in omni necessitate et tribulatione nostra per vestram fidem
1THESS|3|8|quoniam nunc vivimus si vos statis in Domino
1THESS|3|9|quam enim gratiarum actionem possumus Deo retribuere pro vobis in omni gaudio quo gaudemus propter vos ante Deum nostrum
1THESS|3|10|nocte et die abundantius orantes ut videamus faciem vestram et conpleamus ea quae desunt fidei vestrae
1THESS|3|11|ipse autem Deus et Pater noster et Dominus Iesus dirigat viam nostram ad vos
1THESS|3|12|vos autem Dominus multiplicet et abundare faciat caritatem in invicem et in omnes quemadmodum et nos in vobis
1THESS|3|13|ad confirmanda corda vestra sine querella in sanctitate ante Deum et Patrem nostrum in adventu Domini nostri Iesu cum omnibus sanctis eius amen
1THESS|4|1|de cetero ergo fratres rogamus vos et obsecramus in Domino Iesu ut quemadmodum accepistis a nobis quomodo vos oporteat ambulare et placere Deo sicut et ambulatis ut abundetis magis
1THESS|4|2|scitis enim quae praecepta dederimus vobis per Dominum Iesum
1THESS|4|3|haec est enim voluntas Dei sanctificatio vestra
1THESS|4|4|ut abstineatis vos a fornicatione ut sciat unusquisque vestrum suum vas possidere in sanctificatione et honore
1THESS|4|5|non in passione desiderii sicut et gentes quae ignorant Deum
1THESS|4|6|ut ne quis supergrediatur neque circumveniat in negotio fratrem suum quoniam vindex est Dominus de his omnibus sicut et praediximus vobis et testificati sumus
1THESS|4|7|non enim vocavit nos Deus in inmunditia sed in sanctificatione
1THESS|4|8|itaque qui spernit non hominem spernit sed Deum qui etiam dedit Spiritum suum Sanctum in vobis
1THESS|4|9|de caritate autem fraternitatis non necesse habemus scribere vobis ipsi enim vos a Deo didicistis ut diligatis invicem
1THESS|4|10|etenim facitis illud in omnes fratres in universa Macedonia rogamus autem vos fratres ut abundetis magis
1THESS|4|11|et operam detis ut quieti sitis et ut vestrum negotium agatis et operemini manibus vestris sicut praecepimus vobis
1THESS|4|12|et ut honeste ambuletis ad eos qui foris sunt et nullius aliquid desideretis
1THESS|4|13|nolumus autem vos ignorare fratres de dormientibus ut non contristemini sicut et ceteri qui spem non habent
1THESS|4|14|si enim credimus quod Iesus mortuus est et resurrexit ita et Deus eos qui dormierunt per Iesum adducet cum eo
1THESS|4|15|hoc enim vobis dicimus in verbo Domini quia nos qui vivimus qui residui sumus in adventum Domini non praeveniemus eos qui dormierunt
1THESS|4|16|quoniam ipse Dominus in iussu et in voce archangeli et in tuba Dei descendet de caelo et mortui qui in Christo sunt resurgent primi
1THESS|4|17|deinde nos qui vivimus qui relinquimur simul rapiemur cum illis in nubibus obviam Domino in aera et sic semper cum Domino erimus
1THESS|4|18|itaque consolamini invicem in verbis istis
1THESS|5|1|de temporibus autem et momentis fratres non indigetis ut scribamus vobis
1THESS|5|2|ipsi enim diligenter scitis quia dies Domini sicut fur in nocte ita veniet
1THESS|5|3|cum enim dixerint pax et securitas tunc repentinus eis superveniet interitus sicut dolor in utero habenti et non effugient
1THESS|5|4|vos autem fratres non estis in tenebris ut vos dies ille tamquam fur conprehendat
1THESS|5|5|omnes enim vos filii lucis estis et filii diei non sumus noctis neque tenebrarum
1THESS|5|6|igitur non dormiamus sicut ceteri sed vigilemus et sobrii simus
1THESS|5|7|qui enim dormiunt nocte dormiunt et qui ebrii sunt nocte ebrii sunt
1THESS|5|8|nos autem qui diei sumus sobrii simus induti loricam fidei et caritatis et galeam spem salutis
1THESS|5|9|quoniam non posuit nos Deus in iram sed in adquisitionem salutis per Dominum nostrum Iesum Christum
1THESS|5|10|qui mortuus est pro nobis ut sive vigilemus sive dormiamus simul cum illo vivamus
1THESS|5|11|propter quod consolamini invicem et aedificate alterutrum sicut et facitis
1THESS|5|12|rogamus autem vos fratres ut noveritis eos qui laborant inter vos et praesunt vobis in Domino et monent vos
1THESS|5|13|ut habeatis illos abundantius in caritate propter opus illorum pacem habete cum eis
1THESS|5|14|rogamus autem vos fratres corripite inquietos consolamini pusillianimes suscipite infirmos patientes estote ad omnes
1THESS|5|15|videte ne quis malum pro malo alicui reddat sed semper quod bonum est sectamini et in invicem et in omnes
1THESS|5|16|semper gaudete
1THESS|5|17|sine intermissione orate
1THESS|5|18|in omnibus gratias agite haec enim voluntas Dei est in Christo Iesu in omnibus vobis
1THESS|5|19|Spiritum nolite extinguere
1THESS|5|20|prophetias nolite spernere
1THESS|5|21|omnia autem probate quod bonum est tenete
1THESS|5|22|ab omni specie mala abstinete vos
1THESS|5|23|ipse autem Deus pacis sanctificet vos per omnia et integer spiritus vester et anima et corpus sine querella in adventu Domini nostri Iesu Christi servetur
1THESS|5|24|fidelis est qui vocavit vos qui etiam faciet
1THESS|5|25|fratres orate pro nobis
1THESS|5|26|salutate fratres omnes in osculo sancto
1THESS|5|27|adiuro vos per Dominum ut legatur epistula omnibus sanctis fratribus
1THESS|5|28|gratia Domini nostri Iesu Christi vobiscum amen
2THESS|1|1|Paulus et Silvanus et Timotheus ecclesiae Thessalonicensium in Deo Patre nostro et Domino Iesu Christo
2THESS|1|2|gratia vobis et pax a Deo Patre nostro et Domino Iesu Christo
2THESS|1|3|gratias agere debemus Deo semper pro vobis fratres ita ut dignum est quoniam supercrescit fides vestra et abundat caritas uniuscuiusque omnium vestrum in invicem
2THESS|1|4|ita ut et nos ipsi in vobis gloriemur in ecclesiis Dei pro patientia vestra et fide in omnibus persecutionibus vestris et tribulationibus quas sustinetis
2THESS|1|5|in exemplum iusti iudicii Dei ut digni habeamini regno Dei pro quo et patimini
2THESS|1|6|si tamen iustum est apud Deum retribuere tribulationem his qui vos tribulant
2THESS|1|7|et vobis qui tribulamini requiem nobiscum in revelatione Domini Iesu de caelo cum angelis virtutis eius
2THESS|1|8|in flamma ignis dantis vindictam his qui non noverunt Deum et qui non oboediunt evangelio Domini nostri Iesu
2THESS|1|9|qui poenas dabunt in interitu aeternas a facie Domini et a gloria virtutis eius
2THESS|1|10|cum venerit glorificari in sanctis suis et admirabilis fieri in omnibus qui crediderunt quia creditum est testimonium nostrum super vos in die illo
2THESS|1|11|in quo etiam oramus semper pro vobis ut dignetur vos vocatione sua Deus et impleat omnem voluntatem bonitatis et opus fidei in virtute
2THESS|1|12|ut clarificetur nomen Domini nostri Iesu Christi in vobis et vos in illo secundum gratiam Dei nostri et Domini Iesu Christi
2THESS|2|1|rogamus autem vos fratres per adventum Domini nostri Iesu Christi et nostrae congregationis in ipsum
2THESS|2|2|ut non cito moveamini a sensu neque terreamini neque per spiritum neque per sermonem neque per epistulam tamquam per nos quasi instet dies Domini
2THESS|2|3|ne quis vos seducat ullo modo quoniam nisi venerit discessio primum et revelatus fuerit homo peccati filius perditionis
2THESS|2|4|qui adversatur et extollitur supra omne quod dicitur Deus aut quod colitur ita ut in templo Dei sedeat ostendens se quia sit Deus
2THESS|2|5|non retinetis quod cum adhuc essem apud vos haec dicebam vobis
2THESS|2|6|et nunc quid detineat scitis ut reveletur in suo tempore
2THESS|2|7|nam mysterium iam operatur iniquitatis tantum ut qui tenet nunc donec de medio fiat
2THESS|2|8|et tunc revelabitur ille iniquus quem Dominus Iesus interficiet spiritu oris sui et destruet inlustratione adventus sui
2THESS|2|9|eum cuius est adventus secundum operationem Satanae in omni virtute et signis et prodigiis mendacibus
2THESS|2|10|et in omni seductione iniquitatis his qui pereunt eo quod caritatem veritatis non receperunt ut salvi fierent
2THESS|2|11|ideo mittit illis Deus operationem erroris ut credant mendacio
2THESS|2|12|ut iudicentur omnes qui non crediderunt veritati sed consenserunt iniquitati
2THESS|2|13|nos autem debemus gratias agere Deo semper pro vobis fratres dilecti a Deo quod elegerit nos Deus primitias in salutem in sanctificatione Spiritus et fide veritatis
2THESS|2|14|ad quod et vocavit vos per evangelium nostrum in adquisitionem gloriae Domini nostri Iesu Christi
2THESS|2|15|itaque fratres state et tenete traditiones quas didicistis sive per sermonem sive per epistulam nostram
2THESS|2|16|ipse autem Dominus noster Iesus Christus et Deus et Pater noster qui dilexit nos et dedit consolationem aeternam et spem bonam in gratia
2THESS|2|17|exhortetur corda vestra et confirmet in omni opere et sermone bono
2THESS|3|1|de cetero fratres orate pro nobis ut sermo Domini currat et clarificetur sicut et apud vos
2THESS|3|2|et ut liberemur ab inportunis et malis hominibus non enim omnium est fides
2THESS|3|3|fidelis autem Dominus est qui confirmabit vos et custodiet a malo
2THESS|3|4|confidimus autem de vobis in Domino quoniam quae praecipimus et facitis et facietis
2THESS|3|5|Dominus autem dirigat corda vestra in caritate Dei et patientia Christi
2THESS|3|6|denuntiamus autem vobis fratres in nomine Domini nostri Iesu Christi ut subtrahatis vos ab omni fratre ambulante inordinate et non secundum traditionem quam acceperunt a nobis
2THESS|3|7|ipsi enim scitis quemadmodum oporteat imitari nos quoniam non inquieti fuimus inter vos
2THESS|3|8|neque gratis panem manducavimus ab aliquo sed in labore et fatigatione nocte et die operantes ne quem vestrum gravaremus
2THESS|3|9|non quasi non habuerimus potestatem sed ut nosmet ipsos formam daremus vobis ad imitandum nos
2THESS|3|10|nam et cum essemus apud vos hoc denuntiabamus vobis quoniam si quis non vult operari nec manducet
2THESS|3|11|audimus enim inter vos quosdam ambulare inquiete nihil operantes sed curiose agentes
2THESS|3|12|his autem qui eiusmodi sunt denuntiamus et obsecramus in Domino Iesu Christo ut cum silentio operantes suum panem manducent
2THESS|3|13|vos autem fratres nolite deficere benefacientes
2THESS|3|14|quod si quis non oboedit verbo nostro per epistulam hunc notate et non commisceamini cum illo ut confundatur
2THESS|3|15|et nolite quasi inimicum existimare sed corripite ut fratrem
2THESS|3|16|ipse autem Dominus pacis det vobis pacem sempiternam in omni loco Dominus cum omnibus vobis
2THESS|3|17|salutatio mea manu Pauli quod est signum in omni epistula ita scribo
2THESS|3|18|gratia Domini nostri Iesu Christi cum omnibus vobis amen
1TIM|1|1|Paulus apostolus Christi Iesu secundum imperium Dei salvatoris nostri et Christi Iesu spei nostrae
1TIM|1|2|Timotheo dilecto filio in fide gratia misericordia pax a Deo Patre et Christo Iesu Domino nostro
1TIM|1|3|sicut rogavi te ut remaneres Ephesi cum irem in Macedoniam ut denuntiares quibusdam ne aliter docerent
1TIM|1|4|neque intenderent fabulis et genealogiis interminatis quae quaestiones praestant magis quam aedificationem Dei quae est in fide
1TIM|1|5|finis autem praecepti est caritas de corde puro et conscientia bona et fide non ficta
1TIM|1|6|a quibus quidam aberrantes conversi sunt in vaniloquium
1TIM|1|7|volentes esse legis doctores non intellegentes neque quae loquuntur neque de quibus adfirmant
1TIM|1|8|scimus autem quia bona est lex si quis ea legitime utatur
1TIM|1|9|sciens hoc quia iusto lex non est posita sed iniustis et non subditis impiis et peccatoribus sceleratis et contaminatis patricidis et matricidis homicidis
1TIM|1|10|fornicariis masculorum concubitoribus plagiariis mendacibus periuris et si quid aliud sanae doctrinae adversatur
1TIM|1|11|quae est secundum evangelium gloriae beati Dei quod creditum est mihi
1TIM|1|12|gratias ago ei qui me confortavit Christo Iesu Domino nostro quia fidelem me existimavit ponens in ministerio
1TIM|1|13|qui prius fui blasphemus et persecutor et contumeliosus sed misericordiam consecutus sum quia ignorans feci in incredulitate
1TIM|1|14|superabundavit autem gratia Domini nostri cum fide et dilectione quae est in Christo Iesu
1TIM|1|15|fidelis sermo et omni acceptione dignus quia Christus Iesus venit in mundum peccatores salvos facere quorum primus ego sum
1TIM|1|16|sed ideo misericordiam consecutus sum ut in me primo ostenderet Christus Iesus omnem patientiam ad deformationem eorum qui credituri sunt illi in vitam aeternam
1TIM|1|17|regi autem saeculorum inmortali invisibili soli Deo honor et gloria in saecula saeculorum amen
1TIM|1|18|hoc praeceptum commendo tibi fili Timothee secundum praecedentes in te prophetias ut milites in illis bonam militiam
1TIM|1|19|habens fidem et bonam conscientiam quam quidam repellentes circa fidem naufragaverunt
1TIM|1|20|ex quibus est Hymeneus et Alexander quos tradidi Satanae ut discant non blasphemare
1TIM|2|1|obsecro igitur primo omnium fieri obsecrationes orationes postulationes gratiarum actiones pro omnibus hominibus
1TIM|2|2|pro regibus et omnibus qui in sublimitate sunt ut quietam et tranquillam vitam agamus in omni pietate et castitate
1TIM|2|3|hoc enim bonum est et acceptum coram salutari nostro Deo
1TIM|2|4|qui omnes homines vult salvos fieri et ad agnitionem veritatis venire
1TIM|2|5|unus enim Deus unus et mediator Dei et hominum homo Christus Iesus
1TIM|2|6|qui dedit redemptionem semet ipsum pro omnibus testimonium temporibus suis
1TIM|2|7|in quo positus sum ego praedicator et apostolus veritatem dico non mentior doctor gentium in fide et veritate
1TIM|2|8|volo ergo viros orare in omni loco levantes puras manus sine ira et disceptatione
1TIM|2|9|similiter et mulieres in habitu ornato cum verecundia et sobrietate ornantes se non in tortis crinibus aut auro aut margaritis vel veste pretiosa
1TIM|2|10|sed quod decet mulieres promittentes pietatem per opera bona
1TIM|2|11|mulier in silentio discat cum omni subiectione
1TIM|2|12|docere autem mulieri non permitto neque dominari in virum sed esse in silentio
1TIM|2|13|Adam enim primus formatus est deinde Eva
1TIM|2|14|et Adam non est seductus mulier autem seducta in praevaricatione fuit
1TIM|2|15|salvabitur autem per filiorum generationem si permanserint in fide et dilectione et sanctificatione cum sobrietate
1TIM|3|1|fidelis sermo si quis episcopatum desiderat bonum opus desiderat
1TIM|3|2|oportet ergo episcopum inreprehensibilem esse unius uxoris virum sobrium prudentem ornatum hospitalem doctorem
1TIM|3|3|non vinolentum non percussorem sed modestum non litigiosum non cupidum
1TIM|3|4|suae domui bene praepositum filios habentem subditos cum omni castitate
1TIM|3|5|si quis autem domui suae praeesse nescit quomodo ecclesiae Dei diligentiam habebit
1TIM|3|6|non neophytum ne in superbia elatus in iudicium incidat diaboli
1TIM|3|7|oportet autem illum et testimonium habere bonum ab his qui foris sunt ut non in obprobrium incidat et laqueum diaboli
1TIM|3|8|diaconos similiter pudicos non bilingues non multo vino deditos non turpe lucrum sectantes
1TIM|3|9|habentes mysterium fidei in conscientia pura
1TIM|3|10|et hii autem probentur primum et sic ministrent nullum crimen habentes
1TIM|3|11|mulieres similiter pudicas non detrahentes sobrias fideles in omnibus
1TIM|3|12|diacones sint unius uxoris viri qui filiis suis bene praesunt et suis domibus
1TIM|3|13|qui enim bene ministraverint gradum sibi bonum adquirent et multam fiduciam in fide quae est in Christo Iesu
1TIM|3|14|haec tibi scribo sperans venire ad te cito
1TIM|3|15|si autem tardavero ut scias quomodo oporteat te in domo Dei conversari quae est ecclesia Dei vivi columna et firmamentum veritatis
1TIM|3|16|et manifeste magnum est pietatis sacramentum quod manifestatum est in carne iustificatum est in spiritu apparuit angelis praedicatum est gentibus creditum est in mundo adsumptum est in gloria
1TIM|4|1|Spiritus autem manifeste dicit quia in novissimis temporibus discedent quidam a fide adtendentes spiritibus erroris et doctrinis daemoniorum
1TIM|4|2|in hypocrisi loquentium mendacium et cauteriatam habentium suam conscientiam
1TIM|4|3|prohibentium nubere abstinere a cibis quos Deus creavit ad percipiendum cum gratiarum actione fidelibus et his qui cognoverunt veritatem
1TIM|4|4|quia omnis creatura Dei bona et nihil reiciendum quod cum gratiarum actione percipitur
1TIM|4|5|sanctificatur enim per verbum Dei et orationem
1TIM|4|6|haec proponens fratribus bonus eris minister Christi Iesu enutritus verbis fidei et bonae doctrinae quam adsecutus es
1TIM|4|7|ineptas autem et aniles fabulas devita exerce te ipsum ad pietatem
1TIM|4|8|nam corporalis exercitatio ad modicum utilis est pietas autem ad omnia utilis est promissionem habens vitae quae nunc est et futurae
1TIM|4|9|fidelis sermo et omni acceptione dignus
1TIM|4|10|in hoc enim laboramus et maledicimur quia speravimus in Deum vivum qui est salvator omnium hominum maxime fidelium
1TIM|4|11|praecipe haec et doce
1TIM|4|12|nemo adulescentiam tuam contemnat sed exemplum esto fidelium in verbo in conversatione in caritate in fide in castitate
1TIM|4|13|dum venio adtende lectioni exhortationi doctrinae
1TIM|4|14|noli neglegere gratiam quae in te est quae data est tibi per prophetiam cum inpositione manuum presbyterii
1TIM|4|15|haec meditare in his esto ut profectus tuus manifestus sit omnibus
1TIM|4|16|adtende tibi et doctrinae insta in illis hoc enim faciens et te ipsum salvum facies et qui te audiunt
1TIM|5|1|seniorem ne increpaveris sed obsecra ut patrem iuvenes ut fratres
1TIM|5|2|anus ut matres iuvenculas ut sorores in omni castitate
1TIM|5|3|viduas honora quae vere viduae sunt
1TIM|5|4|si qua autem vidua filios aut nepotes habet discant primum domum suam regere et mutuam vicem reddere parentibus hoc enim acceptum est coram Deo
1TIM|5|5|quae autem vere vidua est et desolata speravit in Deum et instat obsecrationibus et orationibus nocte ac die
1TIM|5|6|nam quae in deliciis est vivens mortua est
1TIM|5|7|et hoc praecipe ut inreprehensibiles sint
1TIM|5|8|si quis autem suorum et maxime domesticorum curam non habet fidem negavit et est infideli deterior
1TIM|5|9|vidua eligatur non minus sexaginta annorum quae fuerit unius viri uxor
1TIM|5|10|in operibus bonis testimonium habens si filios educavit si hospitio recepit si sanctorum pedes lavit si tribulationem patientibus subministravit si omne opus bonum subsecuta est
1TIM|5|11|adulescentiores autem viduas devita cum enim luxuriatae fuerint in Christo nubere volunt
1TIM|5|12|habentes damnationem quia primam fidem irritam fecerunt
1TIM|5|13|simul autem et otiosae discunt circumire domos non solum otiosae sed et verbosae et curiosae loquentes quae non oportet
1TIM|5|14|volo ergo iuveniores nubere filios procreare matres familias esse nullam occasionem dare adversario maledicti gratia
1TIM|5|15|iam enim quaedam conversae sunt retro Satanan
1TIM|5|16|si qua fidelis habet viduas subministret illis et non gravetur ecclesia ut his quae vere viduae sunt sufficiat
1TIM|5|17|qui bene praesunt presbyteri duplici honore digni habeantur maxime qui laborant in verbo et doctrina
1TIM|5|18|dicit enim scriptura non infrenabis os bovi trituranti et dignus operarius mercede sua
1TIM|5|19|adversus presbyterum accusationem noli recipere nisi sub duobus et tribus testibus
1TIM|5|20|peccantes coram omnibus argue ut et ceteri timorem habeant
1TIM|5|21|testor coram Deo et Christo Iesu et electis angelis ut haec custodias sine praeiudicio nihil faciens in aliam partem declinando
1TIM|5|22|manus cito nemini inposueris neque communicaveris peccatis alienis te ipsum castum custodi
1TIM|5|23|noli adhuc aquam bibere sed vino modico utere propter stomachum tuum et frequentes tuas infirmitates
1TIM|5|24|quorundam hominum peccata manifesta sunt praecedentia ad iudicium quosdam autem et subsequuntur
1TIM|5|25|similiter et facta bona manifesta sunt et quae aliter se habent abscondi non possunt
1TIM|6|1|quicumque sunt sub iugo servi dominos suos omni honore dignos arbitrentur ne nomen Domini et doctrina blasphemetur
1TIM|6|2|qui autem fideles habent dominos non contemnant quia fratres sunt sed magis serviant quia fideles sunt et dilecti qui beneficii participes sunt haec doce et exhortare
1TIM|6|3|si quis aliter docet et non adquiescit sanis sermonibus Domini nostri Iesu Christi et ei quae secundum pietatem est doctrinae
1TIM|6|4|superbus nihil sciens sed languens circa quaestiones et pugnas verborum ex quibus oriuntur invidiae contentiones blasphemiae suspiciones malae
1TIM|6|5|conflictationes hominum mente corruptorum et qui veritate privati sunt existimantium quaestum esse pietatem
1TIM|6|6|est autem quaestus magnus pietas cum sufficientia
1TIM|6|7|nihil enim intulimus in mundum haut dubium quia nec auferre quid possumus
1TIM|6|8|habentes autem alimenta et quibus tegamur his contenti sumus
1TIM|6|9|nam qui volunt divites fieri incidunt in temptationem et laqueum et desideria multa inutilia et nociva quae mergunt homines in interitum et perditionem
1TIM|6|10|radix enim omnium malorum est cupiditas quam quidam appetentes erraverunt a fide et inseruerunt se doloribus multis
1TIM|6|11|tu autem o homo Dei haec fuge sectare vero iustitiam pietatem fidem caritatem patientiam mansuetudinem
1TIM|6|12|certa bonum certamen fidei adprehende vitam aeternam in qua vocatus es et confessus bonam confessionem coram multis testibus
1TIM|6|13|praecipio tibi coram Deo qui vivificat omnia et Christo Iesu qui testimonium reddidit sub Pontio Pilato bonam confessionem
1TIM|6|14|ut serves mandatum sine macula inreprehensibile usque in adventum Domini nostri Iesu Christi
1TIM|6|15|quem suis temporibus ostendet beatus et solus potens rex regum et Dominus dominantium
1TIM|6|16|qui solus habet inmortalitatem lucem habitans inaccessibilem quem vidit nullus hominum sed nec videre potest cui honor et imperium sempiternum amen
1TIM|6|17|divitibus huius saeculi praecipe non sublime sapere neque sperare in incerto divitiarum sed in Deo qui praestat nobis omnia abunde ad fruendum
1TIM|6|18|bene agere divites fieri in operibus bonis facile tribuere communicare
1TIM|6|19|thesaurizare sibi fundamentum bonum in futurum ut adprehendant veram vitam
1TIM|6|20|o Timothee depositum custodi devitans profanas vocum novitates et oppositiones falsi nominis scientiae
1TIM|6|21|quam quidam promittentes circa fidem exciderunt gratia tecum
2TIM|1|1|Paulus apostolus Christi Iesu per voluntatem Dei secundum promissionem vitae quae est in Christo Iesu
2TIM|1|2|Timotheo carissimo filio gratia misericordia pax a Deo Patre et Christo Iesu Domino nostro
2TIM|1|3|gratias ago Deo cui servio a progenitoribus in conscientia pura quam sine intermissione habeam tui memoriam in orationibus meis nocte ac die
2TIM|1|4|desiderans te videre memor lacrimarum tuarum ut gaudio implear
2TIM|1|5|recordationem accipiens eius fidei quae est in te non ficta quae et habitavit primum in avia tua Loide et matre tua Eunice certus sum autem quod et in te
2TIM|1|6|propter quam causam admoneo te ut resuscites gratiam Dei quae est in te per inpositionem manuum mearum
2TIM|1|7|non enim dedit nobis Deus spiritum timoris sed virtutis et dilectionis et sobrietatis
2TIM|1|8|noli itaque erubescere testimonium Domini nostri neque me vinctum eius sed conlabora evangelio secundum virtutem Dei
2TIM|1|9|qui nos liberavit et vocavit vocatione sancta non secundum opera nostra sed secundum propositum suum et gratiam quae data est nobis in Christo Iesu ante tempora saecularia
2TIM|1|10|manifestata est autem nunc per inluminationem salvatoris nostri Iesu Christi qui destruxit quidem mortem inluminavit autem vitam et incorruptionem per evangelium
2TIM|1|11|in quo positus sum ego praedicator et apostolus et magister gentium
2TIM|1|12|ob quam causam etiam haec patior sed non confundor scio enim cui credidi et certus sum quia potens est depositum meum servare in illum diem
2TIM|1|13|formam habe sanorum verborum quae a me audisti in fide et dilectione in Christo Iesu
2TIM|1|14|bonum depositum custodi per Spiritum Sanctum qui habitat in nobis
2TIM|1|15|scis hoc quod aversi sunt a me omnes qui in Asia sunt ex quibus est Phygelus et Hermogenes
2TIM|1|16|det misericordiam Dominus Onesifori domui quia saepe me refrigeravit et catenam meam non erubuit
2TIM|1|17|sed cum Romam venisset sollicite me quaesivit et invenit
2TIM|1|18|det illi Dominus invenire misericordiam a Domino in illa die et quanta Ephesi ministravit melius tu nosti
2TIM|2|1|tu ergo fili mi confortare in gratia quae est in Christo Iesu
2TIM|2|2|et quae audisti a me per multos testes haec commenda fidelibus hominibus qui idonei erunt et alios docere
2TIM|2|3|labora sicut bonus miles Christi Iesu
2TIM|2|4|nemo militans inplicat se negotiis saecularibus ut ei placeat cui se probavit
2TIM|2|5|nam et qui certat in agone non coronatur nisi legitime certaverit
2TIM|2|6|laborantem agricolam oportet primum de fructibus accipere
2TIM|2|7|intellege quae dico dabit enim tibi Dominus in omnibus intellectum
2TIM|2|8|memor esto Iesum Christum resurrexisse a mortuis ex semine David secundum evangelium meum
2TIM|2|9|in quo laboro usque ad vincula quasi male operans sed verbum Dei non est alligatum
2TIM|2|10|ideo omnia sustineo propter electos ut et ipsi salutem consequantur quae est in Christo Iesu cum gloria caelesti
2TIM|2|11|fidelis sermo nam si conmortui sumus et convivemus
2TIM|2|12|si sustinemus et conregnabimus si negabimus et ille negabit nos
2TIM|2|13|si non credimus ille fidelis manet negare se ipsum non potest
2TIM|2|14|haec commone testificans coram Domino noli verbis contendere in nihil utile ad subversionem audientium
2TIM|2|15|sollicite cura te ipsum probabilem exhibere Deo operarium inconfusibilem recte tractantem verbum veritatis
2TIM|2|16|profana autem inaniloquia devita multum enim proficient ad impietatem
2TIM|2|17|et sermo eorum ut cancer serpit ex quibus est Hymeneus et Philetus
2TIM|2|18|qui a veritate exciderunt dicentes resurrectionem iam factam et subvertunt quorundam fidem
2TIM|2|19|sed firmum fundamentum Dei stetit habens signaculum hoc cognovit Dominus qui sunt eius et discedat ab iniquitate omnis qui nominat nomen Domini
2TIM|2|20|in magna autem domo non solum sunt vasa aurea et argentea sed et lignea et fictilia et quaedam quidem in honorem quaedam autem in contumeliam
2TIM|2|21|si quis ergo emundaverit se ab istis erit vas in honorem sanctificatum et utile Domino ad omne opus bonum paratum
2TIM|2|22|iuvenilia autem desideria fuge sectare vero iustitiam fidem caritatem pacem cum his qui invocant Dominum de corde puro
2TIM|2|23|stultas autem et sine disciplina quaestiones devita sciens quia generant lites
2TIM|2|24|servum autem Domini non oportet litigare sed mansuetum esse ad omnes docibilem patientem
2TIM|2|25|cum modestia corripientem eos qui resistunt nequando det illis Deus paenitentiam ad cognoscendam veritatem
2TIM|2|26|et resipiscant a diaboli laqueis a quo capti tenentur ad ipsius voluntatem
2TIM|3|1|hoc autem scito quod in novissimis diebus instabunt tempora periculosa
2TIM|3|2|et erunt homines se ipsos amantes cupidi elati superbi blasphemi parentibus inoboedientes ingrati scelesti
2TIM|3|3|sine affectione sine pace criminatores incontinentes inmites sine benignitate
2TIM|3|4|proditores protervi tumidi voluptatium amatores magis quam Dei
2TIM|3|5|habentes speciem quidem pietatis virtutem autem eius abnegantes et hos devita
2TIM|3|6|ex his enim sunt qui penetrant domos et captivas ducunt mulierculas oneratas peccatis quae ducuntur variis desideriis
2TIM|3|7|semper discentes et numquam ad scientiam veritatis pervenientes
2TIM|3|8|quemadmodum autem Iannes et Mambres restiterunt Mosi ita et hii resistunt veritati homines corrupti mente reprobi circa fidem
2TIM|3|9|sed ultra non proficient insipientia enim eorum manifesta erit omnibus sicut et illorum fuit
2TIM|3|10|tu autem adsecutus es meam doctrinam institutionem propositum fidem longanimitatem dilectionem patientiam
2TIM|3|11|persecutiones passiones qualia mihi facta sunt Antiochiae Iconii Lystris quales persecutiones sustinui et ex omnibus me eripuit Dominus
2TIM|3|12|et omnes qui volunt pie vivere in Christo Iesu persecutionem patientur
2TIM|3|13|mali autem homines et seductores proficient in peius errantes et in errorem mittentes
2TIM|3|14|tu vero permane in his quae didicisti et credita sunt tibi sciens a quo didiceris
2TIM|3|15|et quia ab infantia sacras litteras nosti quae te possint instruere ad salutem per fidem quae est in Christo Iesu
2TIM|3|16|omnis scriptura divinitus inspirata et utilis ad docendum ad arguendum ad corrigendum ad erudiendum in iustitia
2TIM|3|17|ut perfectus sit homo Dei ad omne opus bonum instructus
2TIM|4|1|testificor coram Deo et Christo Iesu qui iudicaturus est vivos ac mortuos et adventum ipsius et regnum eius
2TIM|4|2|praedica verbum insta oportune inportune argue obsecra increpa in omni patientia et doctrina
2TIM|4|3|erit enim tempus cum sanam doctrinam non sustinebunt sed ad sua desideria coacervabunt sibi magistros prurientes auribus
2TIM|4|4|et a veritate quidem auditum avertent ad fabulas autem convertentur
2TIM|4|5|tu vero vigila in omnibus labora opus fac evangelistae ministerium tuum imple
2TIM|4|6|ego enim iam delibor et tempus meae resolutionis instat
2TIM|4|7|bonum certamen certavi cursum consummavi fidem servavi
2TIM|4|8|in reliquo reposita est mihi iustitiae corona quam reddet mihi Dominus in illa die iustus iudex non solum autem mihi sed et his qui diligunt adventum eius
2TIM|4|9|festina venire ad me cito
2TIM|4|10|Demas enim me dereliquit diligens hoc saeculum et abiit Thessalonicam Crescens in Galliam Titus in Dalmatiam
2TIM|4|11|Lucas est mecum solus Marcum adsume et adduc tecum est enim mihi utilis in ministerium
2TIM|4|12|Tychicum autem misi Ephesum
2TIM|4|13|paenulam quam reliqui Troade apud Carpum veniens adfers et libros maxime autem membranas
2TIM|4|14|Alexander aerarius multa mala mihi ostendit reddat ei Dominus secundum opera eius
2TIM|4|15|quem et tu devita valde enim restitit verbis nostris
2TIM|4|16|in prima mea defensione nemo mihi adfuit sed omnes me dereliquerunt non illis reputetur
2TIM|4|17|Dominus autem mihi adstitit et confortavit me ut per me praedicatio impleatur et audiant omnes gentes et liberatus sum de ore leonis
2TIM|4|18|liberabit me Dominus ab omni opere malo et salvum faciet in regnum suum caeleste cui gloria in saecula saeculorum amen
2TIM|4|19|saluta Priscam et Aquilam et Onesifori domum
2TIM|4|20|Erastus remansit Corinthi Trophimum autem reliqui infirmum Mileti
2TIM|4|21|festina ante hiemem venire salutat te Eubulus et Pudens et Linus et Claudia et fratres omnes
2TIM|4|22|Dominus Iesus cum spiritu tuo gratia nobiscum amen
TITUS|1|1|Paulus servus Dei apostolus autem Iesu Christi secundum fidem electorum Dei et agnitionem veritatis quae secundum pietatem est
TITUS|1|2|in spem vitae aeternae quam promisit qui non mentitur Deus ante tempora saecularia
TITUS|1|3|manifestavit autem temporibus suis verbum suum in praedicatione quae credita est mihi secundum praeceptum salvatoris nostri Dei
TITUS|1|4|Tito dilecto filio secundum communem fidem gratia et pax a Deo Patre et Christo Iesu salvatore nostro
TITUS|1|5|huius rei gratia reliqui te Cretae ut ea quae desunt corrigas et constituas per civitates presbyteros sicut ego tibi disposui
TITUS|1|6|si quis sine crimine est unius uxoris vir filios habens fideles non in accusatione luxuriae aut non subditos
TITUS|1|7|oportet enim episcopum sine crimine esse sicut Dei dispensatorem non superbum non iracundum non vinolentum non percussorem non turpilucri cupidum
TITUS|1|8|sed hospitalem benignum sobrium iustum sanctum continentem
TITUS|1|9|amplectentem eum qui secundum doctrinam est fidelem sermonem ut potens sit et exhortari in doctrina sana et eos qui contradicunt arguere
TITUS|1|10|sunt enim multi et inoboedientes vaniloqui et seductores maxime qui de circumcisione sunt
TITUS|1|11|quos oportet redargui qui universas domos subvertunt docentes quae non oportet turpis lucri gratia
TITUS|1|12|dixit quidam ex illis proprius ipsorum propheta Cretenses semper mendaces malae bestiae ventres pigri
TITUS|1|13|testimonium hoc verum est quam ob causam increpa illos dure ut sani sint in fide
TITUS|1|14|non intendentes iudaicis fabulis et mandatis hominum aversantium se a veritate
TITUS|1|15|omnia munda mundis coinquinatis autem et infidelibus nihil mundum sed inquinatae sunt eorum et mens et conscientia
TITUS|1|16|confitentur se nosse Deum factis autem negant cum sunt abominati et incredibiles et ad omne opus bonum reprobi
TITUS|2|1|tu autem loquere quae decet sanam doctrinam
TITUS|2|2|senes ut sobrii sint pudici prudentes sani fide dilectione patientia
TITUS|2|3|anus similiter in habitu sancto non criminatrices non vino multo servientes bene docentes
TITUS|2|4|ut prudentiam doceant adulescentulas ut viros suos ament filios diligant
TITUS|2|5|prudentes castas domus curam habentes benignas subditas suis viris ut non blasphemetur verbum Dei
TITUS|2|6|iuvenes similiter hortare ut sobrii sint
TITUS|2|7|in omnibus te ipsum praebe exemplum bonorum operum in doctrina integritatem gravitatem
TITUS|2|8|verbum sanum inreprehensibilem ut is qui ex adverso est vereatur nihil habens malum dicere de nobis
TITUS|2|9|servos dominis suis subditos esse in omnibus placentes non contradicentes
TITUS|2|10|non fraudantes, sed in omnibus fidem bonam ostendentes ut doctrinam salutaris nostri Dei ornent in omnibus
TITUS|2|11|apparuit enim gratia Dei salutaris omnibus hominibus
TITUS|2|12|erudiens nos ut abnegantes impietatem et saecularia desideria sobrie et iuste et pie vivamus in hoc saeculo
TITUS|2|13|expectantes beatam spem et adventum gloriae magni Dei et salvatoris nostri Iesu Christi
TITUS|2|14|qui dedit semet ipsum pro nobis ut nos redimeret ab omni iniquitate et mundaret sibi populum acceptabilem sectatorem bonorum operum
TITUS|2|15|haec loquere et exhortare et argue cum omni imperio nemo te contemnat
TITUS|3|1|admone illos principibus et potestatibus subditos esse dicto oboedire ad omne opus bonum paratos esse
TITUS|3|2|neminem blasphemare non litigiosos esse modestos omnem ostendentes mansuetudinem ad omnes homines
TITUS|3|3|eramus enim et nos aliquando insipientes increduli errantes servientes desideriis et voluptatibus variis in malitia et invidia agentes odibiles odientes invicem
TITUS|3|4|cum autem benignitas et humanitas apparuit salvatoris nostri Dei
TITUS|3|5|non ex operibus iustitiae quae fecimus nos sed secundum suam misericordiam salvos nos fecit per lavacrum regenerationis et renovationis Spiritus Sancti
TITUS|3|6|quem effudit in nos abunde per Iesum Christum salvatorem nostrum
TITUS|3|7|ut iustificati gratia ipsius heredes simus secundum spem vitae aeternae
TITUS|3|8|fidelis sermo est et de his volo te confirmare ut curent bonis operibus praeesse qui credunt Deo haec sunt bona et utilia hominibus
TITUS|3|9|stultas autem quaestiones et genealogias et contentiones et pugnas legis devita sunt enim inutiles et vanae
TITUS|3|10|hereticum hominem post unam et secundam correptionem devita
TITUS|3|11|sciens quia subversus est qui eiusmodi est et delinquit proprio iudicio condemnatus
TITUS|3|12|cum misero ad te Arteman aut Tychicum festina ad me venire Nicopolim ibi enim statui hiemare
TITUS|3|13|Zenan legis peritum et Apollo sollicite praemitte ut nihil illis desit
TITUS|3|14|discant autem et nostri bonis operibus praeesse ad usus necessarios ut non sint infructuosi
TITUS|3|15|salutant te qui mecum sunt omnes saluta qui nos amant in fide gratia Dei cum omnibus vobis amen
PHLM|1|1|Paulus vinctus Iesu Christi et Timotheus frater Philemoni dilecto et adiutori nostro
PHLM|1|2|et Appiae sorori et Archippo commilitoni nostro et ecclesiae quae in domo tua est
PHLM|1|3|gratia vobis et pax a Deo Patre nostro et Domino Iesu Christo
PHLM|1|4|gratias ago Deo meo semper memoriam tui faciens in orationibus meis
PHLM|1|5|audiens caritatem tuam et fidem quam habes in Domino Iesu et in omnes sanctos
PHLM|1|6|ut communicatio fidei tuae evidens fiat in agnitione omnis boni in nobis in Christo Iesu
PHLM|1|7|gaudium enim magnum habui et consolationem in caritate tua quia viscera sanctorum requieverunt per te frater
PHLM|1|8|propter quod multam fiduciam habentes in Christo Iesu imperandi tibi quod ad rem pertinet
PHLM|1|9|propter caritatem magis obsecro cum sis talis ut Paulus senex nunc autem et vinctus Iesu Christi
PHLM|1|10|obsecro te de meo filio quem genui in vinculis Onesimo
PHLM|1|11|qui tibi aliquando inutilis fuit nunc autem et tibi et mihi utilis
PHLM|1|12|quem remisi tu autem illum id est mea viscera suscipe
PHLM|1|13|quem ego volueram mecum detinere ut pro te mihi ministraret in vinculis evangelii
PHLM|1|14|sine consilio autem tuo nihil volui facere uti ne velut ex necessitate bonum tuum esset sed voluntarium
PHLM|1|15|forsitan enim ideo discessit ad horam a te ut aeternum illum recipere
PHLM|1|16|iam non ut servum sed plus servo carissimum fratrem maxime mihi quanto autem magis tibi et in carne et in Domino
PHLM|1|17|si ergo habes me socium suscipe illum sicut me
PHLM|1|18|si autem aliquid nocuit tibi aut debet hoc mihi inputa
PHLM|1|19|ego Paulus scripsi mea manu ego reddam ut non dicam tibi quod et te ipsum mihi debes
PHLM|1|20|ita frater ego te fruar in Domino refice viscera mea in Domino
PHLM|1|21|confidens oboedientia tua scripsi tibi sciens quoniam et super id quod dico facies
PHLM|1|22|simul autem et para mihi hospitium nam spero per orationes vestras donari me vobis
PHLM|1|23|salutat te Epaphras concaptivus meus in Christo Iesu
PHLM|1|24|Marcus Aristarchus Demas Lucas adiutores mei
PHLM|1|25|gratia Domini nostri Iesu Christi cum spiritu vestro amen
HEB|1|1|multifariam et multis modis olim Deus loquens patribus in prophetis
HEB|1|2|novissime diebus istis locutus est nobis in Filio quem constituit heredem universorum per quem fecit et saecula
HEB|1|3|qui cum sit splendor gloriae et figura substantiae eius portansque omnia verbo virtutis suae purgationem peccatorum faciens sedit ad dexteram Maiestatis in excelsis
HEB|1|4|tanto melior angelis effectus quanto differentius prae illis nomen hereditavit
HEB|1|5|cui enim dixit aliquando angelorum Filius meus es tu ego hodie genui te et rursum ego ero illi in Patrem et ipse erit mihi in Filium
HEB|1|6|et cum iterum introducit primogenitum in orbem terrae dicit et adorent eum omnes angeli Dei
HEB|1|7|et ad angelos quidem dicit qui facit angelos suos spiritus et ministros suos flammam ignis
HEB|1|8|ad Filium autem thronus tuus Deus in saeculum saeculi et virga aequitatis virga regni tui
HEB|1|9|dilexisti iustitiam et odisti iniquitatem propterea unxit te Deus Deus tuus oleo exultationis prae participibus tuis
HEB|1|10|et tu in principio Domine terram fundasti et opera manuum tuarum sunt caeli
HEB|1|11|ipsi peribunt tu autem permanebis et omnes ut vestimentum veterescent
HEB|1|12|et velut amictum involves eos et mutabuntur tu autem idem es et anni tui non deficient
HEB|1|13|ad quem autem angelorum dixit aliquando sede a dextris meis quoadusque ponam inimicos tuos scabillum pedum tuorum
HEB|1|14|nonne omnes sunt administratorii spiritus in ministerium missi propter eos qui hereditatem capient salutis
HEB|2|1|propterea abundantius oportet observare nos ea quae audivimus ne forte pereffluamus
HEB|2|2|si enim qui per angelos dictus est sermo factus est firmus et omnis praevaricatio et inoboedientia accepit iustam mercedis retributionem
HEB|2|3|quomodo nos effugiemus si tantam neglexerimus salutem quae cum initium accepisset enarrari per Dominum ab eis qui audierunt in nos confirmata est
HEB|2|4|contestante Deo signis et portentis et variis virtutibus et Spiritus Sancti distributionibus secundum suam voluntatem
HEB|2|5|non enim angelis subiecit orbem terrae futurum de quo loquimur
HEB|2|6|testatus est autem in quodam loco quis dicens quid est homo quod memor es eius aut filius hominis quoniam visitas eum
HEB|2|7|minuisti eum paulo minus ab angelis gloria et honore coronasti eum et constituisti eum super opera manuum tuarum
HEB|2|8|omnia subiecisti sub pedibus eius in eo enim quod ei omnia subiecit nihil dimisit non subiectum ei nunc autem necdum videmus omnia subiecta ei
HEB|2|9|eum autem qui modico quam angeli minoratus est videmus Iesum propter passionem mortis gloria et honore coronatum ut gratia Dei pro omnibus gustaret mortem
HEB|2|10|decebat enim eum propter quem omnia et per quem omnia qui multos filios in gloriam adduxerat auctorem salutis eorum per passiones consummare
HEB|2|11|qui enim sanctificat et qui sanctificantur ex uno omnes propter quam causam non confunditur fratres eos vocare dicens
HEB|2|12|nuntiabo nomen tuum fratribus meis in medio ecclesiae laudabo te
HEB|2|13|et iterum ego ero fidens in eum et iterum ecce ego et pueri mei quos mihi dedit Deus
HEB|2|14|quia ergo pueri communicaverunt sanguini et carni et ipse similiter participavit hisdem ut per mortem destrueret eum qui habebat mortis imperium id est diabolum
HEB|2|15|et liberaret eos qui timore mortis per totam vitam obnoxii erant servituti
HEB|2|16|nusquam enim angelos adprehendit sed semen Abrahae adprehendit
HEB|2|17|unde debuit per omnia fratribus similare ut misericors fieret et fidelis pontifex ad Deum ut repropitiaret delicta populi
HEB|2|18|in eo enim in quo passus est ipse temptatus potens est eis qui temptantur auxiliari
HEB|3|1|unde fratres sancti vocationis caelestis participes considerate apostolum et pontificem confessionis nostrae Iesum
HEB|3|2|qui fidelis est ei qui fecit illum sicut et Moses in omni domo illius
HEB|3|3|amplioris enim gloriae iste prae Mose dignus habitus est quanto ampliorem honorem habet domus qui fabricavit illam
HEB|3|4|omnis namque domus fabricatur ab aliquo qui autem omnia creavit Deus
HEB|3|5|et Moses quidem fidelis erat in tota domo eius tamquam famulus in testimonium eorum quae dicenda erant
HEB|3|6|Christus vero tamquam filius in domo sua quae domus sumus nos si fiduciam et gloriam spei usque ad finem firmam retineamus
HEB|3|7|quapropter sicut dicit Spiritus Sanctus hodie si vocem eius audieritis
HEB|3|8|nolite obdurare corda vestra sicut in exacerbatione secundum diem temptationis in deserto
HEB|3|9|ubi temptaverunt me patres vestri probaverunt et viderunt opera mea
HEB|3|10|quadraginta annos propter quod infensus fui generationi huic et dixi semper errant corde ipsi autem non cognoverunt vias meas
HEB|3|11|sicut iuravi in ira mea si introibunt in requiem meam
HEB|3|12|videte fratres ne forte sit in aliquo vestrum cor malum incredulitatis discedendi a Deo vivo
HEB|3|13|sed adhortamini vosmet ipsos per singulos dies donec hodie cognominatur ut non obduretur quis ex vobis fallacia peccati
HEB|3|14|participes enim Christi effecti sumus si tamen initium substantiae usque ad finem firmum retineamus
HEB|3|15|dum dicitur hodie si vocem eius audieritis nolite obdurare corda vestra quemadmodum in illa exacerbatione
HEB|3|16|quidam enim audientes exacerbaverunt sed non universi qui profecti sunt ab Aegypto per Mosen
HEB|3|17|quibus autem infensus est quadraginta annos nonne illis qui peccaverunt quorum cadavera prostrata sunt in deserto
HEB|3|18|quibus autem iuravit non introire in requiem ipsius nisi illis qui increduli fuerunt
HEB|3|19|et videmus quia non potuerunt introire propter incredulitatem
HEB|4|1|timeamus ergo ne forte relicta pollicitatione introeundi in requiem eius existimetur aliqui ex vobis deesse
HEB|4|2|etenim et nobis nuntiatum est quemadmodum et illis sed non profuit illis sermo auditus non admixtis fidei ex his quae audierunt
HEB|4|3|ingrediemur enim in requiem qui credidimus quemadmodum dixit sicut iuravi in ira mea si introibunt in requiem meam et quidem operibus ab institutione mundi factis
HEB|4|4|dixit enim quodam loco de die septima sic et requievit Deus die septima ab omnibus operibus suis
HEB|4|5|et in isto rursum si introibunt in requiem meam
HEB|4|6|quoniam ergo superest quosdam introire in illam et hii quibus prioribus adnuntiatum est non introierunt propter incredulitatem
HEB|4|7|iterum terminat diem quendam hodie in David dicendo post tantum temporis sicut supra dictum est hodie si vocem eius audieritis nolite obdurare corda vestra
HEB|4|8|nam si eis Iesus requiem praestitisset numquam de alio loqueretur posthac die
HEB|4|9|itaque relinquitur sabbatismus populo Dei
HEB|4|10|qui enim ingressus est in requiem eius etiam ipse requievit ab operibus suis sicut a suis Deus
HEB|4|11|festinemus ergo ingredi in illam requiem ut ne in id ipsum quis incidat incredulitatis exemplum
HEB|4|12|vivus est enim Dei sermo et efficax et penetrabilior omni gladio ancipiti et pertingens usque ad divisionem animae ac spiritus conpagum quoque et medullarum et discretor cogitationum et intentionum cordis
HEB|4|13|et non est ulla creatura invisibilis in conspectu eius omnia autem nuda et aperta sunt oculis eius ad quem nobis sermo
HEB|4|14|habentes ergo pontificem magnum qui penetraverit caelos Iesum Filium Dei teneamus confessionem
HEB|4|15|non enim habemus pontificem qui non possit conpati infirmitatibus nostris temptatum autem per omnia pro similitudine absque peccato
HEB|4|16|adeamus ergo cum fiducia ad thronum gratiae ut misericordiam consequamur et gratiam inveniamus in auxilio oportuno
HEB|5|1|omnis namque pontifex ex hominibus adsumptus pro hominibus constituitur in his quae sunt ad Deum ut offerat dona et sacrificia pro peccatis
HEB|5|2|qui condolere possit his qui ignorant et errant quoniam et ipse circumdatus est infirmitate
HEB|5|3|et propter eam debet quemadmodum et pro populo ita etiam pro semet ipso offerre pro peccatis
HEB|5|4|nec quisquam sumit sibi honorem sed qui vocatur a Deo tamquam Aaron
HEB|5|5|sic et Christus non semet ipsum clarificavit ut pontifex fieret sed qui locutus est ad eum Filius meus es tu ego hodie genui te
HEB|5|6|quemadmodum et in alio dicit tu es sacerdos in aeternum secundum ordinem Melchisedech
HEB|5|7|qui in diebus carnis suae preces supplicationesque ad eum qui possit salvum illum a morte facere cum clamore valido et lacrimis offerens et exauditus pro sua reverentia
HEB|5|8|et quidem cum esset Filius didicit ex his quae passus est oboedientiam
HEB|5|9|et consummatus factus est omnibus obtemperantibus sibi causa salutis aeternae
HEB|5|10|appellatus a Deo pontifex iuxta ordinem Melchisedech
HEB|5|11|de quo grandis nobis sermo et ininterpretabilis ad dicendum quoniam inbecilles facti estis ad audiendum
HEB|5|12|etenim cum deberetis magistri esse propter tempus rursum indigetis ut vos doceamini quae sint elementa exordii sermonum Dei et facti estis quibus lacte opus sit non solido cibo
HEB|5|13|omnis enim qui lactis est particeps expers est sermonis iustitiae parvulus enim est
HEB|5|14|perfectorum autem est solidus cibus eorum qui pro consuetudine exercitatos habent sensus ad discretionem boni ac mali
HEB|6|1|quapropter intermittentes inchoationis Christi sermonem ad perfectionem feramur non rursum iacientes fundamentum paenitentiae ab operibus mortuis et fidei ad Deum
HEB|6|2|baptismatum doctrinae inpositionis quoque manuum ac resurrectionis mortuorum et iudicii aeterni
HEB|6|3|et hoc faciemus siquidem permiserit Deus
HEB|6|4|inpossibile est enim eos qui semel sunt inluminati gustaverunt etiam donum caeleste et participes sunt facti Spiritus Sancti
HEB|6|5|gustaverunt nihilominus bonum Dei verbum virtutesque saeculi venturi
HEB|6|6|et prolapsi sunt renovari rursus ad paenitentiam rursum crucifigentes sibimet ipsis Filium Dei et ostentui habentes
HEB|6|7|terra enim saepe venientem super se bibens imbrem et generans herbam oportunam illis a quibus colitur accipit benedictionem a Deo
HEB|6|8|proferens autem spinas ac tribulos reproba est et maledicto proxima cuius consummatio in conbustionem
HEB|6|9|confidimus autem de vobis dilectissimi meliora et viciniora saluti tametsi ita loquimur
HEB|6|10|non enim iniustus Deus ut obliviscatur operis vestri et dilectionis quam ostendistis in nomine ipsius qui ministrastis sanctis et ministratis
HEB|6|11|cupimus autem unumquemque vestrum eandem ostentare sollicitudinem ad expletionem spei usque in finem
HEB|6|12|ut non segnes efficiamini verum imitatores eorum qui fide et patientia hereditabunt promissiones
HEB|6|13|Abrahae namque promittens Deus quoniam neminem habuit per quem iuraret maiorem iuravit per semet ipsum
HEB|6|14|dicens nisi benedicens benedicam te et multiplicans multiplicabo te
HEB|6|15|et sic longanimiter ferens adeptus est repromissionem
HEB|6|16|homines enim per maiorem sui iurant et omnis controversiae eorum finis ad confirmationem est iuramentum
HEB|6|17|in quo abundantius volens Deus ostendere pollicitationis heredibus inmobilitatem consilii sui interposuit iusiurandum
HEB|6|18|ut per duas res inmobiles quibus inpossibile est mentiri Deum fortissimum solacium habeamus qui confugimus ad tenendam propositam spem
HEB|6|19|quam sicut anchoram habemus animae tutam ac firmam et incedentem usque in interiora velaminis
HEB|6|20|ubi praecursor pro nobis introiit Iesus secundum ordinem Melchisedech pontifex factus in aeternum
HEB|7|1|hic enim Melchisedech rex Salem sacerdos Dei summi qui obviavit Abrahae regresso a caede regum et benedixit ei
HEB|7|2|cui decimas omnium divisit Abraham primum quidem qui interpretatur rex iustitiae deinde autem et rex Salem quod est rex pacis
HEB|7|3|sine patre sine matre sine genealogia neque initium dierum neque finem vitae habens adsimilatus autem Filio Dei manet sacerdos in perpetuum
HEB|7|4|intuemini autem quantus sit hic cui et decimam dedit de praecipuis Abraham patriarcha
HEB|7|5|et quidem de filiis Levi sacerdotium accipientes mandatum habent decimas sumere a populo secundum legem id est a fratribus suis quamquam et ipsi exierunt de lumbis Abrahae
HEB|7|6|cuius autem generatio non adnumeratur in eis decimas sumpsit Abraham et hunc qui habebat repromissiones benedixit
HEB|7|7|sine ulla autem contradictione quod minus est a meliore benedicitur
HEB|7|8|et hic quidem decimas morientes homines accipiunt ibi autem contestatus quia vivit
HEB|7|9|et ut ita dictum sit per Abraham et Levi qui decimas accipit decimatus est
HEB|7|10|adhuc enim in lumbis patris erat quando obviavit ei Melchisedech
HEB|7|11|si ergo consummatio per sacerdotium leviticum erat populus enim sub ipso legem accepit quid adhuc necessarium secundum ordinem Melchisedech alium surgere sacerdotem et non secundum ordinem Aaron dici
HEB|7|12|translato enim sacerdotio necesse est ut et legis translatio fiat
HEB|7|13|in quo enim haec dicuntur de alia tribu est de qua nullus altario praesto fuit
HEB|7|14|manifestum enim quod ex Iuda ortus sit Dominus noster in qua tribu nihil de sacerdotibus Moses locutus est
HEB|7|15|et amplius adhuc manifestum est si secundum similitudinem Melchisedech exsurgit alius sacerdos
HEB|7|16|qui non secundum legem mandati carnalis factus est sed secundum virtutem vitae insolubilis
HEB|7|17|contestatur enim quoniam tu es sacerdos in aeternum secundum ordinem Melchisedech
HEB|7|18|reprobatio quidem fit praecedentis mandati propter infirmitatem eius et inutilitatem
HEB|7|19|nihil enim ad perfectum adduxit lex introductio vero melioris spei per quam proximamus ad Deum
HEB|7|20|et quantum est non sine iureiurando alii quidem sine iureiurando sacerdotes facti sunt
HEB|7|21|hic autem cum iureiurando per eum qui dixit ad illum iuravit Dominus et non paenitebit tu es sacerdos in aeternum
HEB|7|22|in tantum melioris testamenti sponsor factus est Iesus
HEB|7|23|et alii quidem plures facti sunt sacerdotes idcirco quod morte prohiberentur permanere
HEB|7|24|hic autem eo quod maneat in aeternum sempiternum habet sacerdotium
HEB|7|25|unde et salvare in perpetuo potest accedentes per semet ipsum ad Deum semper vivens ad interpellandum pro eis
HEB|7|26|talis enim decebat ut nobis esset pontifex sanctus innocens inpollutus segregatus a peccatoribus et excelsior caelis factus
HEB|7|27|qui non habet cotidie necessitatem quemadmodum sacerdotes prius pro suis delictis hostias offerre deinde pro populi hoc enim fecit semel se offerendo
HEB|7|28|lex enim homines constituit sacerdotes infirmitatem habentes sermo autem iurisiurandi qui post legem est Filium in aeternum perfectum
HEB|8|1|capitulum autem super ea quae dicuntur talem habemus pontificem qui consedit in dextera sedis Magnitudinis in caelis
HEB|8|2|sanctorum minister et tabernaculi veri quod fixit Dominus et non homo
HEB|8|3|omnis enim pontifex ad offerenda munera et hostias constituitur unde necesse est et hunc habere aliquid quod offerat
HEB|8|4|si ergo esset super terram nec esset sacerdos cum essent qui offerrent secundum legem munera
HEB|8|5|qui exemplari et umbrae deserviunt caelestium sicut responsum est Mosi cum consummaret tabernaculum vide inquit omnia facito secundum exemplar quod tibi ostensum est in monte
HEB|8|6|nunc autem melius sortitus est ministerium quanto et melioris testamenti mediator est quod in melioribus repromissionibus sanctum est
HEB|8|7|nam si illud prius culpa vacasset non utique secundi locus inquireretur
HEB|8|8|vituperans enim eos dicit ecce dies veniunt dicit Dominus et consummabo super domum Israhel et super domum Iuda testamentum novum
HEB|8|9|non secundum testamentum quod feci patribus eorum in die qua adprehendi manum illorum ut educerem illos de terra Aegypti quoniam ipsi non permanserunt in testamento meo et ego neglexi eos dicit Dominus
HEB|8|10|quia hoc testamentum quod disponam domui Israhel post dies illos dicit Dominus dando leges meas in mentem eorum et in corde eorum superscribam eas et ero eis in Deum et ipsi erunt mihi in populum
HEB|8|11|et non docebit unusquisque proximum suum et unusquisque fratrem suum dicens cognosce Dominum quoniam omnes scient me a minore usque ad maiorem eorum
HEB|8|12|quia propitius ero iniquitatibus eorum et peccatorum illorum iam non memorabor
HEB|8|13|dicendo autem novum veteravit prius quod autem antiquatur et senescit prope interitum est
HEB|9|1|habuit quidem et prius iustificationes culturae et sanctum saeculare
HEB|9|2|tabernaculum enim factum est primum in quo inerant candelabra et mensa et propositio panum quae dicitur sancta
HEB|9|3|post velamentum autem secundum tabernaculum quod dicitur sancta sanctorum
HEB|9|4|aureum habens turibulum et arcam testamenti circumtectam ex omni parte auro in qua urna aurea habens manna et virga Aaron quae fronduerat et tabulae testamenti
HEB|9|5|superque eam cherubin gloriae obumbrantia propitiatorium de quibus non est modo dicendum per singula
HEB|9|6|his vero ita conpositis in priori quidem tabernaculo semper introibant sacerdotes sacrificiorum officia consummantes
HEB|9|7|in secundo autem semel in anno solus pontifex non sine sanguine quem offert pro sua et populi ignorantia
HEB|9|8|hoc significante Spiritu Sancto nondum propalatam esse sanctorum viam adhuc priore tabernaculo habente statum
HEB|9|9|quae parabola est temporis instantis iuxta quam munera et hostiae offeruntur quae non possunt iuxta conscientiam perfectum facere servientem
HEB|9|10|solummodo in cibis et in potibus et variis baptismis et iustitiis carnis usque ad tempus correctionis inpositis
HEB|9|11|Christus autem adsistens pontifex futurorum bonorum per amplius et perfectius tabernaculum non manufactum id est non huius creationis
HEB|9|12|neque per sanguinem hircorum et vitulorum sed per proprium sanguinem introivit semel in sancta aeterna redemptione inventa
HEB|9|13|si enim sanguis hircorum et taurorum et cinis vitulae aspersus inquinatos sanctificat ad emundationem carnis
HEB|9|14|quanto magis sanguis Christi qui per Spiritum Sanctum semet ipsum obtulit inmaculatum Deo emundabit conscientiam vestram ab operibus mortuis ad serviendum Deo viventi
HEB|9|15|et ideo novi testamenti mediator est ut morte intercedente in redemptionem earum praevaricationum quae erant sub priore testamento repromissionem accipiant qui vocati sunt aeternae hereditatis
HEB|9|16|ubi enim testamentum mors necesse est intercedat testatoris
HEB|9|17|testamentum enim in mortuis confirmatum est alioquin nondum valet dum vivit qui testatus est
HEB|9|18|unde ne primum quidem sine sanguine dedicatum est
HEB|9|19|lecto enim omni mandato legis a Mose universo populo accipiens sanguinem vitulorum et hircorum cum aqua et lana coccinea et hysopo ipsum quoque librum et omnem populum aspersit
HEB|9|20|dicens hic sanguis testamenti quod mandavit ad vos Deus
HEB|9|21|etiam tabernaculum et omnia vasa ministerii sanguine similiter aspersit
HEB|9|22|et omnia paene in sanguine mundantur secundum legem et sine sanguinis fusione non fit remissio
HEB|9|23|necesse est ergo exemplaria quidem caelestium his mundari ipsa autem caelestia melioribus hostiis quam istis
HEB|9|24|non enim in manufactis sanctis Iesus introiit exemplaria verorum sed in ipsum caelum ut appareat nunc vultui Dei pro nobis
HEB|9|25|neque ut saepe offerat semet ipsum quemadmodum pontifex intrat in sancta per singulos annos in sanguine alieno
HEB|9|26|alioquin oportebat eum frequenter pati ab origine mundi nunc autem semel in consummatione saeculorum ad destitutionem peccati per hostiam suam apparuit
HEB|9|27|et quemadmodum statutum est hominibus semel mori post hoc autem iudicium
HEB|9|28|sic et Christus semel oblatus ad multorum exhaurienda peccata secundo sine peccato apparebit expectantibus se in salutem
HEB|10|1|umbram enim habens lex bonorum futurorum non ipsam imaginem rerum per singulos annos hisdem ipsis hostiis quas offerunt indesinenter numquam potest accedentes perfectos facere
HEB|10|2|alioquin non cessassent offerri ideo quod nullam haberent ultra conscientiam peccati cultores semel mundati
HEB|10|3|sed in ipsis commemoratio peccatorum per singulos annos fit
HEB|10|4|inpossibile enim est sanguine taurorum et hircorum auferri peccata
HEB|10|5|ideo ingrediens mundum dicit hostiam et oblationem noluisti corpus autem aptasti mihi
HEB|10|6|holocaustomata et pro peccato non tibi placuit
HEB|10|7|tunc dixi ecce venio in capitulo libri scriptum est de me ut faciam Deus voluntatem tuam
HEB|10|8|superius dicens quia hostias et oblationes et holocaustomata et pro peccato noluisti nec placita sunt tibi quae secundum legem offeruntur
HEB|10|9|tunc dixit ecce venio ut faciam Deus voluntatem tuam aufert primum ut sequens statuat
HEB|10|10|in qua voluntate sanctificati sumus per oblationem corporis Christi Iesu in semel
HEB|10|11|et omnis quidem sacerdos praesto est cotidie ministrans et easdem saepe offerens hostias quae numquam possunt auferre peccata
HEB|10|12|hic autem unam pro peccatis offerens hostiam in sempiternum sedit in dextera Dei
HEB|10|13|de cetero expectans donec ponantur inimici eius scabillum pedum eius
HEB|10|14|una enim oblatione consummavit in sempiternum sanctificatos
HEB|10|15|contestatur autem nos et Spiritus Sanctus postquam enim dixit
HEB|10|16|hoc autem testamentum quod testabor ad illos post dies illos dicit Dominus dando leges meas in cordibus eorum et in mente eorum superscribam eas
HEB|10|17|et peccatorum et iniquitatium eorum iam non recordabor amplius
HEB|10|18|ubi autem horum remissio iam non oblatio pro peccato
HEB|10|19|habentes itaque fratres fiduciam in introitu sanctorum in sanguine Christi
HEB|10|20|quam initiavit nobis viam novam et viventem per velamen id est carnem suam
HEB|10|21|et sacerdotem magnum super domum Dei
HEB|10|22|accedamus cum vero corde in plenitudine fidei aspersi corda a conscientia mala et abluti corpus aqua munda
HEB|10|23|teneamus spei nostrae confessionem indeclinabilem fidelis enim est qui repromisit
HEB|10|24|et consideremus invicem in provocationem caritatis et bonorum operum
HEB|10|25|non deserentes collectionem nostram sicut est consuetudinis quibusdam sed consolantes et tanto magis quanto videritis adpropinquantem diem
HEB|10|26|voluntarie enim peccantibus nobis post acceptam notitiam veritatis iam non relinquitur pro peccatis hostia
HEB|10|27|terribilis autem quaedam expectatio iudicii et ignis aemulatio quae consumptura est adversarios
HEB|10|28|irritam quis faciens legem Mosi sine ulla miseratione duobus vel tribus testibus moritur
HEB|10|29|quanto magis putatis deteriora mereri supplicia qui Filium Dei conculcaverit et sanguinem testamenti pollutum duxerit in quo sanctificatus est et Spiritui gratiae contumeliam fecerit
HEB|10|30|scimus enim qui dixit mihi vindictam ego reddam et iterum quia iudicabit Dominus populum suum
HEB|10|31|horrendum est incidere in manus Dei viventis
HEB|10|32|rememoramini autem pristinos dies in quibus inluminati magnum certamen sustinuistis passionum
HEB|10|33|et in altero quidem obprobriis et tribulationibus spectaculum facti in altero autem socii taliter conversantium effecti
HEB|10|34|nam et vinctis conpassi estis et rapinam bonorum vestrorum cum gaudio suscepistis cognoscentes vos habere meliorem et manentem substantiam
HEB|10|35|nolite itaque amittere confidentiam vestram quae magnam habet remunerationem
HEB|10|36|patientia enim vobis necessaria est ut voluntatem Dei facientes reportetis promissionem
HEB|10|37|adhuc enim modicum quantulum qui venturus est veniet et non tardabit
HEB|10|38|iustus autem meus ex fide vivit quod si subtraxerit se non placebit animae meae
HEB|10|39|nos autem non sumus subtractionis in perditionem sed fidei in adquisitionem animae
HEB|11|1|est autem fides sperandorum substantia rerum argumentum non parentum
HEB|11|2|in hac enim testimonium consecuti sunt senes
HEB|11|3|fide intellegimus aptata esse saecula verbo Dei ut ex invisibilibus visibilia fierent
HEB|11|4|fide plurimam hostiam Abel quam Cain obtulit Deo per quam testimonium consecutus est esse iustus testimonium perhibente muneribus eius Deo et per illam defunctus adhuc loquitur
HEB|11|5|fide Enoch translatus est ne videret mortem et non inveniebatur quia transtulit illum Deus ante translationem enim testimonium habebat placuisse Deo
HEB|11|6|sine fide autem inpossibile placere credere enim oportet accedentem ad Deum quia est et inquirentibus se remunerator fit
HEB|11|7|fide Noe responso accepto de his quae adhuc non videbantur metuens aptavit arcam in salutem domus suae per quam damnavit mundum et iustitiae quae per fidem est heres est institutus
HEB|11|8|fide qui vocatur Abraham oboedivit in locum exire quem accepturus erat in hereditatem et exiit nesciens quo iret
HEB|11|9|fide moratus est in terra repromissionis tamquam in aliena in casulis habitando cum Isaac et Iacob coheredibus repromissionis eiusdem
HEB|11|10|expectabat enim fundamenta habentem civitatem cuius artifex et conditor Deus
HEB|11|11|fide et ipsa Sarra sterilis virtutem in conceptionem seminis accepit etiam praeter tempus aetatis quoniam fidelem credidit esse qui promiserat
HEB|11|12|propter quod et ab uno orti sunt et haec emortuo tamquam sidera caeli in multitudinem et sicut harena quae est ad oram maris innumerabilis
HEB|11|13|iuxta fidem defuncti sunt omnes isti non acceptis repromissionibus sed a longe eas aspicientes et salutantes et confitentes quia peregrini et hospites sunt supra terram
HEB|11|14|qui enim haec dicunt significant se patriam inquirere
HEB|11|15|et si quidem illius meminissent de qua exierunt habebant utique tempus revertendi
HEB|11|16|nunc autem meliorem appetunt id est caelestem ideo non confunditur Deus vocari Deus eorum paravit enim illis civitatem
HEB|11|17|fide obtulit Abraham Isaac cum temptaretur et unigenitum offerebat qui susceperat repromissiones
HEB|11|18|ad quem dictum est quia in Isaac vocabitur tibi semen
HEB|11|19|arbitrans quia et a mortuis suscitare potens est Deus unde eum et in parabola accepit
HEB|11|20|fide et de futuris benedixit Isaac Iacob et Esau
HEB|11|21|fide Iacob moriens singulis filiorum Ioseph benedixit et adoravit fastigium virgae eius
HEB|11|22|fide Ioseph moriens de profectione filiorum Israhel memoratus est et de ossibus suis mandavit
HEB|11|23|fide Moses natus occultatus est mensibus tribus a parentibus suis eo quod vidissent elegantem infantem et non timuerunt regis edictum
HEB|11|24|fide Moses grandis factus negavit se esse filium filiae Pharaonis
HEB|11|25|magis eligens adfligi cum populo Dei quam temporalis peccati habere iucunditatem
HEB|11|26|maiores divitias aestimans thesauro Aegyptiorum inproperium Christi aspiciebat enim in remunerationem
HEB|11|27|fide reliquit Aegyptum non veritus animositatem regis invisibilem enim tamquam videns sustinuit
HEB|11|28|fide celebravit pascha et sanguinis effusionem ne qui vastabat primitiva tangeret eos
HEB|11|29|fide transierunt mare Rubrum tamquam per aridam terram quod experti Aegyptii devorati sunt
HEB|11|30|fide muri Hiericho ruerunt circuiti dierum septem
HEB|11|31|fide Raab meretrix non periit cum incredulis excipiens exploratores cum pace
HEB|11|32|et quid adhuc dicam deficiet enim me tempus enarrantem de Gedeon Barac Samson Iepthae David et Samuhel et prophetis
HEB|11|33|qui per fidem devicerunt regna operati sunt iustitiam adepti sunt repromissiones obturaverunt ora leonum
HEB|11|34|extinxerunt impetum ignis effugerunt aciem gladii convaluerunt de infirmitate fortes facti sunt in bello castra verterunt exterorum
HEB|11|35|acceperunt mulieres de resurrectione mortuos suos alii autem distenti sunt non suscipientes redemptionem ut meliorem invenirent resurrectionem
HEB|11|36|alii vero ludibria et verbera experti insuper et vincula et carceres
HEB|11|37|lapidati sunt secti sunt temptati sunt in occisione gladii mortui sunt circumierunt in melotis in pellibus caprinis egentes angustiati adflicti
HEB|11|38|quibus dignus non erat mundus in solitudinibus errantes et montibus et speluncis et in cavernis terrae
HEB|11|39|et hii omnes testimonio fidei probati non acceperunt repromissionem
HEB|11|40|Deo pro nobis melius aliquid providente ut ne sine nobis consummarentur
HEB|12|1|ideoque et nos tantam habentes inpositam nubem testium deponentes omne pondus et circumstans nos peccatum per patientiam curramus propositum nobis certamen
HEB|12|2|aspicientes in auctorem fidei et consummatorem Iesum qui pro proposito sibi gaudio sustinuit crucem confusione contempta atque in dextera sedis Dei sedit
HEB|12|3|recogitate enim eum qui talem sustinuit a peccatoribus adversum semet ipsos contradictionem ut ne fatigemini animis vestris deficientes
HEB|12|4|nondum usque ad sanguinem restitistis adversus peccatum repugnantes
HEB|12|5|et obliti estis consolationis quae vobis tamquam filiis loquitur dicens fili mi noli neglegere disciplinam Domini neque fatigeris dum ab eo argueris
HEB|12|6|quem enim diligit Dominus castigat flagellat autem omnem filium quem recipit
HEB|12|7|in disciplina perseverate tamquam filiis vobis offert Deus quis enim filius quem non corripit pater
HEB|12|8|quod si extra disciplinam estis cuius participes facti sunt omnes ergo adulteri et non filii estis
HEB|12|9|deinde patres quidem carnis nostrae habuimus eruditores et reverebamur non multo magis obtemperabimus Patri spirituum et vivemus
HEB|12|10|et illi quidem in tempore paucorum dierum secundum voluntatem suam erudiebant nos hic autem ad id quod utile est in recipiendo sanctificationem eius
HEB|12|11|omnis autem disciplina in praesenti quidem videtur non esse gaudii sed maeroris postea autem fructum pacatissimum exercitatis per eam reddit iustitiae
HEB|12|12|propter quod remissas manus et soluta genua erigite
HEB|12|13|et gressus rectos facite pedibus vestris ut non claudicans erret magis autem sanetur
HEB|12|14|pacem sequimini cum omnibus et sanctimoniam sine qua nemo videbit Dominum
HEB|12|15|contemplantes ne quis desit gratiae Dei ne qua radix amaritudinis sursum germinans inpediat et per illam inquinentur multi
HEB|12|16|ne quis fornicator aut profanus ut Esau qui propter unam escam vendidit primitiva sua
HEB|12|17|scitote enim quoniam et postea cupiens hereditare benedictionem reprobatus est non enim invenit paenitentiae locum quamquam cum lacrimis inquisisset eam
HEB|12|18|non enim accessistis ad tractabilem et accensibilem ignem et turbinem et caliginem et procellam
HEB|12|19|et tubae sonum et vocem verborum quam qui audierunt excusaverunt se ne eis fieret verbum
HEB|12|20|non enim portabant quod dicebatur et si bestia tetigerit montem lapidabitur
HEB|12|21|et ita terribile erat quod videbatur Moses dixit exterritus sum et tremebundus
HEB|12|22|sed accessistis ad Sion montem et civitatem Dei viventis Hierusalem caelestem et multorum milium angelorum frequentiae
HEB|12|23|et ecclesiam primitivorum qui conscripti sunt in caelis et iudicem omnium Deum et spiritus iustorum perfectorum
HEB|12|24|et testamenti novi mediatorem Iesum et sanguinis sparsionem melius loquentem quam Abel
HEB|12|25|videte ne recusetis loquentem si enim illi non effugerunt recusantes eum qui super terram loquebatur multo magis nos qui de caelis loquentem nobis avertimur
HEB|12|26|cuius vox movit terram tunc modo autem repromittit dicens adhuc semel ego movebo non solum terram sed et caelum
HEB|12|27|quod autem adhuc semel dicit declarat mobilium translationem tamquam factorum ut maneant ea quae sunt inmobilia
HEB|12|28|itaque regnum inmobile suscipientes habemus gratiam per quam serviamus placentes Deo cum metu et reverentia
HEB|12|29|etenim Deus noster ignis consumens est
HEB|13|1|caritas fraternitatis maneat
HEB|13|2|hospitalitatem nolite oblivisci per hanc enim latuerunt quidam angelis hospitio receptis
HEB|13|3|mementote vinctorum tamquam simul vincti et laborantium tamquam et ipsi in corpore morantes
HEB|13|4|honorabile conubium in omnibus et torus inmaculatus fornicatores enim et adulteros iudicabit Deus
HEB|13|5|sint mores sine avaritia contenti praesentibus ipse enim dixit non te deseram neque derelinquam
HEB|13|6|ita ut confidenter dicamus Dominus mihi adiutor non timebo quid faciat mihi homo
HEB|13|7|mementote praepositorum vestrorum qui vobis locuti sunt verbum Dei quorum intuentes exitum conversationis imitamini fidem
HEB|13|8|Iesus Christus heri et hodie ipse et in saecula
HEB|13|9|doctrinis variis et peregrinis nolite abduci optimum enim est gratia stabiliri cor non escis quae non profuerunt ambulantibus in eis
HEB|13|10|habemus altare de quo edere non habent potestatem qui tabernaculo deserviunt
HEB|13|11|quorum enim animalium infertur sanguis pro peccato in sancta per pontificem horum corpora cremantur extra castra
HEB|13|12|propter quod et Iesus ut sanctificaret per suum sanguinem populum extra portam passus est
HEB|13|13|exeamus igitur ad eum extra castra inproperium eius portantes
HEB|13|14|non enim habemus hic manentem civitatem sed futuram inquirimus
HEB|13|15|per ipsum ergo offeramus hostiam laudis semper Deo id est fructum labiorum confitentium nomini eius
HEB|13|16|beneficientiae autem et communionis nolite oblivisci talibus enim hostiis promeretur Deus
HEB|13|17|oboedite praepositis vestris et subiacete eis ipsi enim pervigilant quasi rationem pro animabus vestris reddituri ut cum gaudio hoc faciant et non gementes hoc enim non expedit vobis
HEB|13|18|orate pro nobis confidimus enim quia bonam conscientiam habemus in omnibus bene volentes conversari
HEB|13|19|amplius autem deprecor vos hoc facere ut quo celerius restituar vobis
HEB|13|20|Deus autem pacis qui eduxit de mortuis pastorem magnum ovium in sanguine testamenti aeterni Dominum nostrum Iesum
HEB|13|21|aptet vos in omni bono ut faciatis voluntatem eius faciens in vobis quod placeat coram se per Iesum Christum cui gloria in saecula saeculorum amen
HEB|13|22|rogo autem vos fratres sufferatis verbum solacii etenim perpaucis scripsi vobis
HEB|13|23|cognoscite fratrem nostrum Timotheum dimissum cum quo si celerius venerit videbo vos
HEB|13|24|salutate omnes praepositos vestros et omnes sanctos salutant vos de Italia
HEB|13|25|gratia cum omnibus vobis amen
JAS|1|1|Iacobus Dei et Domini nostri Iesu Christi servus duodecim tribubus quae sunt in dispersione salutem
JAS|1|2|omne gaudium existimate fratres mei cum in temptationibus variis incideritis
JAS|1|3|scientes quod probatio fidei vestrae patientiam operatur
JAS|1|4|patientia autem opus perfectum habeat ut sitis perfecti et integri in nullo deficientes
JAS|1|5|si quis autem vestrum indiget sapientiam postulet a Deo qui dat omnibus affluenter et non inproperat et dabitur ei
JAS|1|6|postulet autem in fide nihil haesitans qui enim haesitat similis est fluctui maris qui a vento movetur et circumfertur
JAS|1|7|non ergo aestimet homo ille quod accipiat aliquid a Domino
JAS|1|8|vir duplex animo inconstans in omnibus viis suis
JAS|1|9|glorietur autem frater humilis in exaltatione sua
JAS|1|10|dives autem in humilitate sua quoniam sicut flos faeni transibit
JAS|1|11|exortus est enim sol cum ardore et arefecit faenum et flos eius decidit et decor vultus eius deperiit ita et dives in itineribus suis marcescet
JAS|1|12|beatus vir qui suffert temptationem quia cum probatus fuerit accipiet coronam vitae quam repromisit Deus diligentibus se
JAS|1|13|nemo cum temptatur dicat quoniam a Deo temptor Deus enim intemptator malorum est ipse autem neminem temptat
JAS|1|14|unusquisque vero temptatur a concupiscentia sua abstractus et inlectus
JAS|1|15|dein concupiscentia cum conceperit parit peccatum peccatum vero cum consummatum fuerit generat mortem
JAS|1|16|nolite itaque errare fratres mei dilectissimi
JAS|1|17|omne datum optimum et omne donum perfectum desursum est descendens a Patre luminum apud quem non est transmutatio nec vicissitudinis obumbratio
JAS|1|18|voluntarie genuit nos verbo veritatis ut simus initium aliquod creaturae eius
JAS|1|19|scitis fratres mei dilecti sit autem omnis homo velox ad audiendum tardus autem ad loquendum et tardus ad iram
JAS|1|20|ira enim viri iustitiam Dei non operatur
JAS|1|21|propter quod abicientes omnem inmunditiam et abundantiam malitiae in mansuetudine suscipite insitum verbum quod potest salvare animas vestras
JAS|1|22|estote autem factores verbi et non auditores tantum fallentes vosmet ipsos
JAS|1|23|quia si quis auditor est verbi et non factor hic conparabitur viro consideranti vultum nativitatis suae in speculo
JAS|1|24|consideravit enim se et abiit et statim oblitus est qualis fuerit
JAS|1|25|qui autem perspexerit in lege perfecta libertatis et permanserit non auditor obliviosus factus sed factor operis hic beatus in facto suo erit
JAS|1|26|si quis autem putat se religiosum esse non refrenans linguam suam sed seducens cor suum huius vana est religio
JAS|1|27|religio munda et inmaculata apud Deum et Patrem haec est visitare pupillos et viduas in tribulatione eorum inmaculatum se custodire ab hoc saeculo
JAS|2|1|fratres mei nolite in personarum acceptione habere fidem Domini nostri Iesu Christi gloriae
JAS|2|2|etenim si introierit in conventu vestro vir aureum anulum habens in veste candida introierit autem et pauper in sordido habitu
JAS|2|3|et intendatis in eum qui indutus est veste praeclara et dixeritis tu sede hic bene pauperi autem dicatis tu sta illic aut sede sub scabillo pedum meorum
JAS|2|4|nonne iudicatis apud vosmet ipsos et facti estis iudices cogitationum iniquarum
JAS|2|5|audite fratres mei dilectissimi nonne Deus elegit pauperes in hoc mundo divites in fide et heredes regni quod repromisit Deus diligentibus se
JAS|2|6|vos autem exhonorastis pauperem nonne divites per potentiam opprimunt vos et ipsi trahunt vos ad iudicia
JAS|2|7|nonne ipsi blasphemant bonum nomen quod invocatum est super vos
JAS|2|8|si tamen legem perficitis regalem secundum scripturas diliges proximum tuum sicut te ipsum bene facitis
JAS|2|9|si autem personas accipitis peccatum operamini redarguti a lege quasi transgressores
JAS|2|10|quicumque autem totam legem servaverit offendat autem in uno factus est omnium reus
JAS|2|11|qui enim dixit non moechaberis dixit et non occides quod si non moechaberis occides autem factus es transgressor legis
JAS|2|12|sic loquimini et sic facite sicut per legem libertatis incipientes iudicari
JAS|2|13|iudicium enim sine misericordia illi qui non fecit misericordiam superexultat autem misericordia iudicio
JAS|2|14|quid proderit fratres mei si fidem quis dicat se habere opera autem non habeat numquid poterit fides salvare eum
JAS|2|15|si autem frater aut soror nudi sunt et indigent victu cotidiano
JAS|2|16|dicat autem aliquis de vobis illis ite in pace calefacimini et saturamini non dederitis autem eis quae necessaria sunt corporis quid proderit
JAS|2|17|sic et fides si non habeat opera mortua est in semet ipsam
JAS|2|18|sed dicet quis tu fidem habes et ego opera habeo ostende mihi fidem tuam sine operibus et ego ostendam tibi ex operibus fidem meam
JAS|2|19|tu credis quoniam unus est Deus bene facis et daemones credunt et contremescunt
JAS|2|20|vis autem scire o homo inanis quoniam fides sine operibus otiosa est
JAS|2|21|Abraham pater noster nonne ex operibus iustificatus est offerens Isaac filium suum super altare
JAS|2|22|vides quoniam fides cooperabatur operibus illius et ex operibus fides consummata est
JAS|2|23|et suppleta est scriptura dicens credidit Abraham Deo et reputatum est illi ad iustitiam et amicus Dei appellatus est
JAS|2|24|videtis quoniam ex operibus iustificatur homo et non ex fide tantum
JAS|2|25|similiter autem et Raab meretrix nonne ex operibus iustificata est suscipiens nuntios et alia via eiciens
JAS|2|26|sicut enim corpus sine spiritu emortuum est ita et fides sine operibus mortua est
JAS|3|1|nolite plures magistri fieri fratres mei scientes quoniam maius iudicium sumitis
JAS|3|2|in multis enim offendimus omnes si quis in verbo non offendit hic perfectus est vir potens etiam freno circumducere totum corpus
JAS|3|3|si autem equorum frenos in ora mittimus ad consentiendum nobis et omne corpus illorum circumferimus
JAS|3|4|ecce et naves cum magnae sint et a ventis validis minentur circumferuntur a modico gubernaculo ubi impetus dirigentis voluerit
JAS|3|5|ita et lingua modicum quidem membrum est et magna exultat ecce quantus ignis quam magnam silvam incendit
JAS|3|6|et lingua ignis est universitas iniquitatis lingua constituitur in membris nostris quae maculat totum corpus et inflammat rotam nativitatis nostrae inflammata a gehenna
JAS|3|7|omnis enim natura bestiarum et volucrum et serpentium etiam ceterorum domantur et domita sunt a natura humana
JAS|3|8|linguam autem nullus hominum domare potest inquietum malum plena veneno mortifero
JAS|3|9|in ipsa benedicimus Dominum et Patrem et in ipsa maledicimus homines qui ad similitudinem Dei facti sunt
JAS|3|10|ex ipso ore procedit benedictio et maledictio non oportet fratres mei haec ita fieri
JAS|3|11|numquid fons de eodem foramine emanat dulcem et amaram aquam
JAS|3|12|numquid potest fratres mei ficus olivas facere aut vitis ficus sic neque salsa dulcem potest facere aquam
JAS|3|13|quis sapiens et disciplinatus inter vos ostendat ex bona conversatione operationem suam in mansuetudine sapientiae
JAS|3|14|quod si zelum amarum habetis et contentiones in cordibus vestris nolite gloriari et mendaces esse adversus veritatem
JAS|3|15|non est ista sapientia desursum descendens sed terrena animalis diabolica
JAS|3|16|ubi enim zelus et contentio ibi inconstantia et omne opus pravum
JAS|3|17|quae autem desursum est sapientia primum quidem pudica est deinde pacifica modesta suadibilis plena misericordia et fructibus bonis non iudicans sine simulatione
JAS|3|18|fructus autem iustitiae in pace seminatur facientibus pacem
JAS|4|1|unde bella et lites in vobis nonne hinc ex concupiscentiis vestris quae militant in membris vestris
JAS|4|2|concupiscitis et non habetis occiditis et zelatis et non potestis adipisci litigatis et belligeratis non habetis propter quod non postulatis
JAS|4|3|petitis et non accipitis eo quod male petatis ut in concupiscentiis vestris insumatis
JAS|4|4|adulteri nescitis quia amicitia huius mundi inimica est Dei quicumque ergo voluerit amicus esse saeculi huius inimicus Dei constituitur
JAS|4|5|aut putatis quia inaniter scriptura dicat ad invidiam concupiscit Spiritus qui inhabitat in nobis
JAS|4|6|maiorem autem dat gratiam propter quod dicit Deus superbis resistit humilibus autem dat gratiam
JAS|4|7|subditi igitur estote Deo resistite autem diabolo et fugiet a vobis
JAS|4|8|adpropiate Domino et adpropinquabit vobis emundate manus peccatores et purificate corda duplices animo
JAS|4|9|miseri estote et lugete et plorate risus vester in luctum convertatur et gaudium in maerorem
JAS|4|10|humiliamini in conspectu Domini et exaltabit vos
JAS|4|11|nolite detrahere de alterutrum fratres qui detrahit fratri aut qui iudicat fratrem suum detrahit legi et iudicat legem si autem iudicas legem non es factor legis sed iudex
JAS|4|12|unus est legislator et iudex qui potest perdere et liberare tu autem quis es qui iudicas proximum
JAS|4|13|ecce nunc qui dicitis hodie aut crastino ibimus in illam civitatem et faciemus quidem ibi annum et mercabimur et lucrum faciemus
JAS|4|14|qui ignoratis quid erit in crastinum quae enim est vita vestra vapor est ad modicum parens deinceps exterminatur
JAS|4|15|pro eo ut dicatis si Dominus voluerit et vixerimus faciemus hoc aut illud
JAS|4|16|nunc autem exultatis in superbiis vestris omnis exultatio talis maligna est
JAS|4|17|scienti igitur bonum facere et non facienti peccatum est illi
JAS|5|1|age nunc divites plorate ululantes in miseriis quae advenient vobis
JAS|5|2|divitiae vestrae putrefactae sunt et vestimenta vestra a tineis comesta sunt
JAS|5|3|aurum et argentum vestrum eruginavit et erugo eorum in testimonium vobis erit et manducabit carnes vestras sicut ignis thesaurizastis in novissimis diebus
JAS|5|4|ecce merces operariorum qui messuerunt regiones vestras qui fraudatus est a vobis clamat et clamor ipsorum in aures Domini Sabaoth introiit
JAS|5|5|epulati estis super terram et in luxuriis enutristis corda vestra in die occisionis
JAS|5|6|addixistis occidistis iustum non resistit vobis
JAS|5|7|patientes igitur estote fratres usque ad adventum Domini ecce agricola expectat pretiosum fructum terrae patienter ferens donec accipiat temporivum et serotinum
JAS|5|8|patientes estote et vos confirmate corda vestra quoniam adventus Domini adpropinquavit
JAS|5|9|nolite ingemescere fratres in alterutrum ut non iudicemini ecce iudex ante ianuam adsistit
JAS|5|10|exemplum accipite fratres laboris et patientiae prophetas qui locuti sunt in nomine Domini
JAS|5|11|ecce beatificamus qui sustinuerunt sufferentiam Iob audistis et finem Domini vidistis quoniam misericors est Dominus et miserator
JAS|5|12|ante omnia autem fratres mei nolite iurare neque per caelum neque per terram neque aliud quodcumque iuramentum sit autem vestrum est est non non uti non sub iudicio decidatis
JAS|5|13|tristatur aliquis vestrum oret aequo animo est psallat
JAS|5|14|infirmatur quis in vobis inducat presbyteros ecclesiae et orent super eum unguentes eum oleo in nomine Domini
JAS|5|15|et oratio fidei salvabit infirmum et adlevabit eum Dominus et si in peccatis sit dimittentur ei
JAS|5|16|confitemini ergo alterutrum peccata vestra et orate pro invicem ut salvemini multum enim valet deprecatio iusti adsidua
JAS|5|17|Helias homo erat similis nobis passibilis et oratione oravit ut non plueret super terram et non pluit annos tres et menses sex
JAS|5|18|et rursum oravit et caelum dedit pluviam et terra dedit fructum suum
JAS|5|19|fratres mei si quis ex vobis erraverit a veritate et converterit quis eum
JAS|5|20|scire debet quoniam qui converti fecerit peccatorem ab errore viae suae salvabit animam eius a morte et operit multitudinem peccatorum
1PET|1|1|Petrus apostolus Iesu Christi electis advenis dispersionis Ponti Galatiae Cappadociae Asiae et Bithyniae
1PET|1|2|secundum praescientiam Dei Patris in sanctificatione Spiritus in oboedientiam et aspersionem sanguinis Iesu Christi gratia vobis et pax multiplicetur
1PET|1|3|benedictus Deus et Pater Domini nostri Iesu Christi qui secundum magnam misericordiam suam regeneravit nos in spem vivam per resurrectionem Iesu Christi ex mortuis
1PET|1|4|in hereditatem incorruptibilem et incontaminatam et inmarcescibilem conservatam in caelis in vobis
1PET|1|5|qui in virtute Dei custodimini per fidem in salutem paratam revelari in tempore novissimo
1PET|1|6|in quo exultatis modicum nunc si oportet contristati in variis temptationibus
1PET|1|7|ut probatum vestrae fidei multo pretiosius sit auro quod perit per ignem probato inveniatur in laudem et gloriam et honorem in revelatione Iesu Christi
1PET|1|8|quem cum non videritis diligitis in quem nunc quoque non videntes credentes autem exultatis laetitia inenarrabili et glorificata
1PET|1|9|reportantes finem fidei vestrae salutem animarum
1PET|1|10|de qua salute exquisierunt atque scrutati sunt prophetae qui de futura in vobis gratia prophetaverunt
1PET|1|11|scrutantes in quod vel quale tempus significaret in eis Spiritus Christi praenuntians eas quae in Christo sunt passiones et posteriores glorias
1PET|1|12|quibus revelatum est quia non sibi ipsis vobis autem ministrabant ea quae nunc nuntiata sunt vobis per eos qui evangelizaverunt vos Spiritu Sancto misso de caelo in quae desiderant angeli prospicere
1PET|1|13|propter quod succincti lumbos mentis vestrae sobrii perfecte sperate in eam quae offertur vobis gratiam in revelatione Iesu Christi
1PET|1|14|quasi filii oboedientiae non configurati prioribus ignorantiae vestrae desideriis
1PET|1|15|sed secundum eum qui vocavit vos sanctum et ipsi sancti in omni conversatione sitis
1PET|1|16|quoniam scriptum est sancti eritis quia ego sanctus sum
1PET|1|17|et si Patrem invocatis eum qui sine acceptione personarum iudicat secundum uniuscuiusque opus in timore incolatus vestri tempore conversamini
1PET|1|18|scientes quod non corruptibilibus argento vel auro redempti estis de vana vestra conversatione paternae traditionis
1PET|1|19|sed pretioso sanguine quasi agni incontaminati et inmaculati Christi
1PET|1|20|praecogniti quidem ante constitutionem mundi manifestati autem novissimis temporibus propter vos
1PET|1|21|qui per ipsum fideles estis in Deo qui suscitavit eum a mortuis et dedit ei gloriam ut fides vestra et spes esset in Deo
1PET|1|22|animas vestras castificantes in oboedientia caritatis in fraternitatis amore simplici ex corde invicem diligite adtentius
1PET|1|23|renati non ex semine corruptibili sed incorruptibili per verbum Dei vivi et permanentis
1PET|1|24|quia omnis caro ut faenum et omnis gloria eius tamquam flos faeni exaruit faenum et flos decidit
1PET|1|25|verbum autem Domini manet in aeternum hoc est autem verbum quod evangelizatum est in vos
1PET|2|1|deponentes igitur omnem malitiam et omnem dolum et simulationes et invidias et omnes detractiones
1PET|2|2|sicut modo geniti infantes rationale sine dolo lac concupiscite ut in eo crescatis in salutem
1PET|2|3|si gustastis quoniam dulcis Dominus
1PET|2|4|ad quem accedentes lapidem vivum ab hominibus quidem reprobatum a Deo autem electum honorificatum
1PET|2|5|et ipsi tamquam lapides vivi superaedificamini domus spiritalis sacerdotium sanctum offerre spiritales hostias acceptabiles Deo per Iesum Christum
1PET|2|6|propter quod continet in scriptura ecce pono in Sion lapidem summum angularem electum pretiosum et qui crediderit in eo non confundetur
1PET|2|7|vobis igitur honor credentibus non credentibus autem lapis quem reprobaverunt aedificantes hic factus est in caput anguli
1PET|2|8|et lapis offensionis et petra scandali qui offendunt verbo nec credunt in quod et positi sunt
1PET|2|9|vos autem genus electum regale sacerdotium gens sancta populus adquisitionis ut virtutes adnuntietis eius qui de tenebris vos vocavit in admirabile lumen suum
1PET|2|10|qui aliquando non populus nunc autem populus Dei qui non consecuti misericordiam nunc autem misericordiam consecuti
1PET|2|11|carissimi obsecro tamquam advenas et peregrinos abstinere vos a carnalibus desideriis quae militant adversus animam
1PET|2|12|conversationem vestram inter gentes habentes bonam ut in eo quod detractant de vobis tamquam de malefactoribus ex bonis operibus considerantes glorificent Deum in die visitationis
1PET|2|13|subiecti estote omni humanae creaturae propter Dominum sive regi quasi praecellenti
1PET|2|14|sive ducibus tamquam ab eo missis ad vindictam malefactorum laudem vero bonorum
1PET|2|15|quia sic est voluntas Dei ut benefacientes obmutescere faciatis inprudentium hominum ignorantiam
1PET|2|16|quasi liberi et non quasi velamen habentes malitiae libertatem sed sicut servi Dei
1PET|2|17|omnes honorate fraternitatem diligite Deum timete regem honorificate
1PET|2|18|servi subditi in omni timore dominis non tantum bonis et modestis sed etiam discolis
1PET|2|19|haec est enim gratia si propter conscientiam Dei sustinet quis tristitias patiens iniuste
1PET|2|20|quae enim gloria est si peccantes et colaphizati suffertis sed si benefacientes et patientes sustinetis haec est gratia apud Deum
1PET|2|21|in hoc enim vocati estis quia et Christus passus est pro vobis vobis relinquens exemplum ut sequamini vestigia eius
1PET|2|22|qui peccatum non fecit nec inventus est dolus in ore ipsius
1PET|2|23|qui cum malediceretur non maledicebat cum pateretur non comminabatur tradebat autem iudicanti se iniuste
1PET|2|24|qui peccata nostra ipse pertulit in corpore suo super lignum ut peccatis mortui iustitiae viveremus cuius livore sanati estis
1PET|2|25|eratis enim sicut oves errantes sed conversi estis nunc ad pastorem et episcopum animarum vestrarum
1PET|3|1|similiter mulieres subditae suis viris ut et si qui non credunt verbo per mulierum conversationem sine verbo lucri fiant
1PET|3|2|considerantes in timore castam conversationem vestram
1PET|3|3|quarum sit non extrinsecus capillaturae aut circumdatio auri aut indumenti vestimentorum cultus
1PET|3|4|sed qui absconditus cordis est homo in incorruptibilitate quieti et modesti spiritus quod est in conspectu Dei locuples
1PET|3|5|sic enim aliquando et sanctae mulieres sperantes in Deo ornabant se subiectae propriis viris
1PET|3|6|sicut Sarra oboediebat Abrahae dominum eum vocans cuius estis filiae benefacientes et non timentes ullam perturbationem
1PET|3|7|viri similiter cohabitantes secundum scientiam quasi infirmiori vaso muliebri inpertientes honorem tamquam et coheredibus gratiae vitae uti ne inpediantur orationes vestrae
1PET|3|8|in fine autem omnes unianimes conpatientes fraternitatis amatores misericordes humiles
1PET|3|9|non reddentes malum pro malo vel maledictum pro maledicto sed e contrario benedicentes quia in hoc vocati estis ut benedictionem hereditate possideatis
1PET|3|10|qui enim vult vitam diligere et videre dies bonos coerceat linguam suam a malo et labia eius ne loquantur dolum
1PET|3|11|declinet autem a malo et faciat bonum inquirat pacem et persequatur eam
1PET|3|12|quia oculi Domini super iustos et aures eius in preces eorum vultus autem Domini super facientes mala
1PET|3|13|et quis est qui vobis noceat si boni aemulatores fueritis
1PET|3|14|sed et si quid patimini propter iustitiam beati timorem autem eorum ne timueritis et non conturbemini
1PET|3|15|Dominum autem Christum sanctificate in cordibus vestris parati semper ad satisfactionem omni poscenti vos rationem de ea quae in vobis est spe
1PET|3|16|sed cum modestia et timore conscientiam habentes bonam ut in eo quod detrahunt vobis confundantur qui calumniantur vestram bonam in Christo conversationem
1PET|3|17|melius est enim benefacientes si velit voluntas Dei pati quam malefacientes
1PET|3|18|quia et Christus semel pro peccatis mortuus est iustus pro iniustis ut nos offerret Deo mortificatus carne vivificatus autem spiritu
1PET|3|19|in quo et his qui in carcere erant spiritibus veniens praedicavit
1PET|3|20|qui increduli fuerant aliquando quando expectabat Dei patientia in diebus Noe cum fabricaretur arca in qua pauci id est octo animae salvae factae sunt per aquam
1PET|3|21|quod et vos nunc similis formae salvos facit baptisma non carnis depositio sordium sed conscientiae bonae interrogatio in Deum per resurrectionem Iesu Christi
1PET|3|22|qui est in dextera Dei profectus in caelum subiectis sibi angelis et potestatibus et virtutibus
1PET|4|1|Christo igitur passo in carne et vos eadem cogitatione armamini quia qui passus est carne desiit a peccatis
1PET|4|2|ut iam non hominum desideriis sed voluntate Dei quod reliquum est in carne vivat temporis
1PET|4|3|sufficit enim praeteritum tempus ad voluntatem gentium consummandam qui ambulaverunt in luxuriis desideriis vinolentiis comesationibus potationibus et inlicitis idolorum cultibus
1PET|4|4|in quo peregrinantur non concurrentibus vobis in eandem luxuriae confusionem blasphemantes
1PET|4|5|qui reddent rationem ei qui paratus est iudicare vivos et mortuos
1PET|4|6|propter hoc enim et mortuis evangelizatum est ut iudicentur quidem secundum homines in carne vivant autem secundum Deum spiritu
1PET|4|7|omnium autem finis adpropinquavit estote itaque prudentes et vigilate in orationibus
1PET|4|8|ante omnia mutuam in vosmet ipsos caritatem continuam habentes quia caritas operit multitudinem peccatorum
1PET|4|9|hospitales invicem sine murmuratione
1PET|4|10|unusquisque sicut accepit gratiam in alterutrum illam administrantes sicut boni dispensatores multiformis gratiae Dei
1PET|4|11|si quis loquitur quasi sermones Dei si quis ministrat tamquam ex virtute quam administrat Deus ut in omnibus honorificetur Deus per Iesum Christum cui est gloria et imperium in saecula saeculorum amen
1PET|4|12|carissimi nolite peregrinari in fervore qui ad temptationem vobis fit quasi novi aliquid vobis contingat
1PET|4|13|sed communicantes Christi passionibus gaudete ut et in revelatione gloriae eius gaudeatis exultantes
1PET|4|14|si exprobramini in nomine Christi beati quoniam gloriae Dei Spiritus in vobis requiescit
1PET|4|15|nemo enim vestrum patiatur quasi homicida aut fur aut maledicus aut alienorum appetitor
1PET|4|16|si autem ut Christianus non erubescat glorificet autem Deum in isto nomine
1PET|4|17|quoniam tempus ut incipiat iudicium de domo Dei si autem primum a nobis qui finis eorum qui non credunt Dei evangelio
1PET|4|18|et si iustus vix salvatur impius et peccator ubi parebit
1PET|4|19|itaque et hii qui patiuntur secundum voluntatem Dei fideli creatori commendant animas suas in benefactis
1PET|5|1|seniores ergo qui in vobis sunt obsecro consenior et testis Christi passionum qui et eius quae in futuro revelanda est gloriae communicator
1PET|5|2|pascite qui est in vobis gregem Dei providentes non coacto sed spontanee secundum Deum neque turpis lucri gratia sed voluntarie
1PET|5|3|neque ut dominantes in cleris sed formae facti gregi et ex animo
1PET|5|4|et cum apparuerit princeps pastorum percipietis inmarcescibilem gloriae coronam
1PET|5|5|similiter adulescentes subditi estote senioribus omnes autem invicem humilitatem insinuate quia Deus superbis resistit humilibus autem dat gratiam
1PET|5|6|humiliamini igitur sub potenti manu Dei ut vos exaltet in tempore visitationis
1PET|5|7|omnem sollicitudinem vestram proicientes in eum quoniam ipsi cura est de vobis
1PET|5|8|sobrii estote vigilate quia adversarius vester diabolus tamquam leo rugiens circuit quaerens quem devoret
1PET|5|9|cui resistite fortes fide scientes eadem passionum ei quae in mundo est vestrae fraternitati fieri
1PET|5|10|Deus autem omnis gratiae qui vocavit nos in aeternam suam gloriam in Christo Iesu modicum passos ipse perficiet confirmabit solidabit
1PET|5|11|ipsi imperium in saecula saeculorum amen
1PET|5|12|per Silvanum vobis fidelem fratrem ut arbitror breviter scripsi obsecrans et contestans hanc esse veram gratiam Dei in qua state
1PET|5|13|salutat vos quae est in Babylone cumelecta et Marcus filius meus
1PET|5|14|salutate invicem in osculo sancto gratia vobis omnibus qui estis in Christo
2PET|1|1|Simon Petrus servus et apostolus Iesu Christi his qui coaequalem nobis sortiti sunt fidem in iustitia Dei nostri et salvatoris Iesu Christi
2PET|1|2|gratia vobis et pax adimpleatur in cognitione Domini nostri
2PET|1|3|quomodo omnia nobis divinae virtutis suae quae ad vitam et pietatem donata est per cognitionem eius qui vocavit nos propria gloria et virtute
2PET|1|4|per quae maxima et pretiosa nobis promissa donavit ut per haec efficiamini divinae consortes naturae fugientes eius quae in mundo est concupiscentiae corruptionem
2PET|1|5|vos autem curam omnem subinferentes ministrate in fide vestra virtutem in virtute autem scientiam
2PET|1|6|in scientia autem abstinentiam in abstinentia autem patientiam in patientia autem pietatem
2PET|1|7|in pietate autem amorem fraternitatis in amore autem fraternitatis caritatem
2PET|1|8|haec enim vobis cum adsint et superent non vacuos nec sine fructu vos constituent in Domini nostri Iesu Christi cognitione
2PET|1|9|cui enim non praesto sunt haec caecus est et manu temptans oblivionem accipiens purgationis veterum suorum delictorum
2PET|1|10|quapropter fratres magis satagite ut per bona opera certam vestram vocationem et electionem faciatis haec enim facientes non peccabitis aliquando
2PET|1|11|sic enim abundanter ministrabitur vobis introitus in aeternum regnum Domini nostri et salvatoris Iesu Christi
2PET|1|12|propter quod incipiam vos semper commonere de his et quidem scientes et confirmatos in praesenti veritate
2PET|1|13|iustum autem arbitror quamdiu sum in hoc tabernaculo suscitare vos in commonitione
2PET|1|14|certus quod velox est depositio tabernaculi mei secundum quod et Dominus noster Iesus Christus significavit mihi
2PET|1|15|dabo autem operam et frequenter habere vos post obitum meum ut horum memoriam faciatis
2PET|1|16|non enim doctas fabulas secuti notam fecimus vobis Domini nostri Iesu Christi virtutem et praesentiam sed speculatores facti illius magnitudinis
2PET|1|17|accipiens enim a Deo Patre honorem et gloriam voce delapsa ad eum huiuscemodi a magnifica gloria hic est Filius meus dilectus in quo mihi conplacui
2PET|1|18|et hanc vocem nos audivimus de caelo adlatam cum essemus cum ipso in monte sancto
2PET|1|19|et habemus firmiorem propheticum sermonem cui bene facitis adtendentes quasi lucernae lucenti in caliginoso loco donec dies inlucescat et lucifer oriatur in cordibus vestris
2PET|1|20|hoc primum intellegentes quod omnis prophetia scripturae propria interpretatione non fit
2PET|1|21|non enim voluntate humana adlata est aliquando prophetia sed Spiritu Sancto inspirati locuti sunt sancti Dei homines
2PET|2|1|fuerunt vero et pseudoprophetae in populo sicut et in vobis erunt magistri mendaces qui introducent sectas perditionis et eum qui emit eos Dominum negant superducentes sibi celerem perditionem
2PET|2|2|et multi sequentur eorum luxurias per quos via veritatis blasphemabitur
2PET|2|3|et in avaritia fictis verbis de vobis negotiabuntur quibus iudicium iam olim non cessat et perditio eorum non dormitat
2PET|2|4|si enim Deus angelis peccantibus non pepercit sed rudentibus inferni detractos in tartarum tradidit in iudicium cruciatos reservari
2PET|2|5|et originali mundo non pepercit sed octavum Noe iustitiae praeconem custodivit diluvium mundo impiorum inducens
2PET|2|6|et civitates Sodomorum et Gomorraeorum in cinerem redigens eversione damnavit exemplum eorum qui impie acturi sunt ponens
2PET|2|7|et iustum Loth oppressum a nefandorum iniuria conversatione eruit
2PET|2|8|aspectu enim et auditu iustus erat habitans apud eos qui diem de die animam iustam iniquis operibus cruciabant
2PET|2|9|novit Dominus pios de temptatione eripere iniquos vero in diem iudicii cruciandos reservare
2PET|2|10|magis autem eos qui post carnem in concupiscentia inmunditiae ambulant dominationemque contemnunt audaces sibi placentes sectas non metuunt blasphemantes
2PET|2|11|ubi angeli fortitudine et virtute cum sint maiores non portant adversum se execrabile iudicium
2PET|2|12|hii vero velut inrationabilia pecora naturaliter in captionem et in perniciem in his quae ignorant blasphemantes in corruptione sua et peribunt
2PET|2|13|percipientes mercedem iniustitiae voluptatem existimantes diei delicias coinquinationes et maculae deliciis affluentes in conviviis suis luxuriantes vobiscum
2PET|2|14|oculos habentes plenos adulterio et incessabiles delicti pellicentes animas instabiles cor exercitatum avaritiae habentes maledictionis filii
2PET|2|15|derelinquentes rectam viam erraverunt secuti viam Balaam ex Bosor qui mercedem iniquitatis amavit
2PET|2|16|correptionem vero habuit suae vesaniae subiugale mutum in hominis voce loquens prohibuit prophetae insipientiam
2PET|2|17|hii sunt fontes sine aqua et nebulae turbinibus exagitatae quibus caligo tenebrarum reservatur
2PET|2|18|superba enim vanitatis loquentes pellicent in desideriis carnis luxuriae eos qui paululum effugiunt qui in errore conversantur
2PET|2|19|libertatem illis promittentes cum ipsi servi sint corruptionis a quo enim quis superatus est huius et servus est
2PET|2|20|si enim refugientes coinquinationes mundi in cognitione Domini nostri et salvatoris Iesu Christi his rursus inpliciti superantur facta sunt eis posteriora deteriora prioribus
2PET|2|21|melius enim erat illis non cognoscere viam iustitiae quam post agnitionem retrorsum converti ab eo quod illis traditum est sancto mandato
2PET|2|22|contigit enim eis illud veri proverbii canis reversus ad suum vomitum et sus lota in volutabro luti
2PET|3|1|hanc ecce vobis carissimi secundam scribo epistulam in quibus excito vestram in commonitione sinceram mentem
2PET|3|2|ut memores sitis eorum quae praedixi verborum a sanctis prophetis et apostolorum vestrorum praeceptorum Domini et salvatoris
2PET|3|3|hoc primum scientes quod venient in novissimis diebus in deceptione inlusores iuxta proprias concupiscentias ambulantes
2PET|3|4|dicentes ubi est promissio aut adventus eius ex quo enim patres dormierunt omnia sic perseverant ab initio creaturae
2PET|3|5|latet enim eos hoc volentes quod caeli erant prius et terra de aqua et per aquam consistens Dei verbo
2PET|3|6|per quae ille tunc mundus aqua inundatus periit
2PET|3|7|caeli autem qui nunc sunt et terra eodem verbo repositi sunt igni servati in diem iudicii et perditionis impiorum hominum
2PET|3|8|unum vero hoc non lateat vos carissimi quia unus dies apud Dominum sicut mille anni et mille anni sicut dies unus
2PET|3|9|non tardat Dominus promissi sed patienter agit propter vos nolens aliquos perire sed omnes ad paenitentiam reverti
2PET|3|10|adveniet autem dies Domini ut fur in qua caeli magno impetu transient elementa vero calore solventur
2PET|3|11|cum haec igitur omnia dissolvenda sint quales oportet esse vos in sanctis conversationibus et pietatibus
2PET|3|12|expectantes et properantes in adventum Dei diei per quam caeli ardentes solventur et elementa ignis ardore tabescent
2PET|3|13|novos vero caelos et novam terram et promissa ipsius expectamus in quibus iustitia habitat
2PET|3|14|propter quod carissimi haec expectantes satis agite inmaculati et inviolati ei inveniri in pace
2PET|3|15|et Domini nostri longanimitatem salutem arbitramini sicut et carissimus frater noster Paulus secundum datam sibi sapientiam scripsit vobis
2PET|3|16|sicut et in omnibus epistulis loquens in eis de his in quibus sunt quaedam difficilia intellectu quae indocti et instabiles depravant sicut et ceteras scripturas ad suam ipsorum perditionem
2PET|3|17|vos igitur fratres praescientes custodite ne insipientium errore transducti excidatis a propria firmitate
2PET|3|18|crescite vero in gratia et in cognitione Domini nostri et salvatoris Iesu Christi ipsi gloria et nunc et in die aeternitatis amen
1JOHN|1|1|quod fuit ab initio quod audivimus quod vidimus oculis nostris quod perspeximus et manus nostrae temptaverunt de verbo vitae
1JOHN|1|2|et vita manifestata est et vidimus et testamur et adnuntiamus vobis vitam aeternam quae erat apud Patrem et apparuit nobis
1JOHN|1|3|quod vidimus et audivimus adnuntiamus et vobis ut et vos societatem habeatis nobiscum et societas nostra sit cum Patre et cum Filio eius Iesu Christo
1JOHN|1|4|et haec scribimus vobis ut gaudium nostrum sit plenum
1JOHN|1|5|et haec est adnuntiatio quam audivimus ab eo et adnuntiamus vobis quoniam Deus lux est et tenebrae in eo non sunt ullae
1JOHN|1|6|si dixerimus quoniam societatem habemus cum eo et in tenebris ambulamus mentimur et non facimus veritatem
1JOHN|1|7|si autem in luce ambulemus sicut et ipse est in luce societatem habemus ad invicem et sanguis Iesu Filii eius mundat nos ab omni peccato
1JOHN|1|8|si dixerimus quoniam peccatum non habemus ipsi nos seducimus et veritas in nobis non est
1JOHN|1|9|si confiteamur peccata nostra fidelis est et iustus ut remittat nobis peccata et emundet nos ab omni iniquitate
1JOHN|1|10|si dixerimus quoniam non peccavimus mendacem facimus eum et verbum eius non est in nobis
1JOHN|2|1|filioli mei haec scribo vobis ut non peccetis sed et si quis peccaverit advocatum habemus apud Patrem Iesum Christum iustum
1JOHN|2|2|et ipse est propitiatio pro peccatis nostris non pro nostris autem tantum sed etiam pro totius mundi
1JOHN|2|3|et in hoc scimus quoniam cognovimus eum si mandata eius observemus
1JOHN|2|4|qui dicit se nosse eum et mandata eius non custodit mendax est in hoc veritas non est
1JOHN|2|5|qui autem servat verbum eius vere in hoc caritas Dei perfecta est in hoc scimus quoniam in ipso sumus
1JOHN|2|6|qui dicit se in ipso manere debet sicut ille ambulavit et ipse ambulare
1JOHN|2|7|carissimi non mandatum novum scribo vobis sed mandatum vetus quod habuistis ab initio mandatum vetus est verbum quod audistis
1JOHN|2|8|iterum mandatum novum scribo vobis quod est verum et in ipso et in vobis quoniam tenebrae transeunt et lumen verum iam lucet
1JOHN|2|9|qui dicit se in luce esse et fratrem suum odit in tenebris est usque adhuc
1JOHN|2|10|qui diligit fratrem suum in lumine manet et scandalum in eo non est
1JOHN|2|11|qui autem odit fratrem suum in tenebris est et in tenebris ambulat et nescit quo eat quoniam tenebrae obcaecaverunt oculos eius
1JOHN|2|12|scribo vobis filioli quoniam remittuntur vobis peccata propter nomen eius
1JOHN|2|13|scribo vobis patres quoniam cognovistis eum qui ab initio est scribo vobis adulescentes quoniam vicistis malignum
1JOHN|2|14|scripsi vobis infantes quoniam cognovistis Patrem scripsi vobis patres quia cognovistis eum qui ab initio scripsi vobis adulescentes quia fortes estis et verbum Dei in vobis manet et vicistis malignum
1JOHN|2|15|nolite diligere mundum neque ea quae in mundo sunt si quis diligit mundum non est caritas Patris in eo
1JOHN|2|16|quoniam omne quod est in mundo concupiscentia carnis et concupiscentia oculorum est et superbia vitae quae non est ex Patre sed ex mundo est
1JOHN|2|17|et mundus transit et concupiscentia eius qui autem facit voluntatem Dei manet in aeternum
1JOHN|2|18|filioli novissima hora est et sicut audistis quia antichristus venit nunc antichristi multi facti sunt unde scimus quoniam novissima hora est
1JOHN|2|19|ex nobis prodierunt sed non erant ex nobis nam si fuissent ex nobis permansissent utique nobiscum sed ut manifesti sint quoniam non sunt omnes ex nobis
1JOHN|2|20|sed vos unctionem habetis a Sancto et nostis omnia
1JOHN|2|21|non scripsi vobis quasi ignorantibus veritatem sed quasi scientibus eam et quoniam omne mendacium ex veritate non est
1JOHN|2|22|quis est mendax nisi is qui negat quoniam Iesus non est Christus hic est antichristus qui negat Patrem et Filium
1JOHN|2|23|omnis qui negat Filium nec Patrem habet qui confitetur Filium et Patrem habet
1JOHN|2|24|vos quod audistis ab initio in vobis permaneat si in vobis permanserit quod ab initio audistis et vos in Filio et Patre manebitis
1JOHN|2|25|et haec est repromissio quam ipse pollicitus est nobis vitam aeternam
1JOHN|2|26|haec scripsi vobis de eis qui seducunt vos
1JOHN|2|27|et vos unctionem quam accepistis ab eo manet in vobis et non necesse habetis ut aliquis doceat vos sed sicut unctio eius docet vos de omnibus et verum est et non est mendacium et sicut docuit vos manete in eo
1JOHN|2|28|et nunc filioli manete in eo ut cum apparuerit habeamus fiduciam et non confundamur ab eo in adventu eius
1JOHN|2|29|si scitis quoniam iustus est scitote quoniam et omnis qui facit iustitiam ex ipso natus est
1JOHN|3|1|videte qualem caritatem dedit nobis Pater ut filii Dei nominemur et sumus propter hoc mundus non novit nos quia non novit eum
1JOHN|3|2|carissimi nunc filii Dei sumus et nondum apparuit quid erimus scimus quoniam cum apparuerit similes ei erimus quoniam videbimus eum sicuti est
1JOHN|3|3|et omnis qui habet spem hanc in eo sanctificat se sicut et ille sanctus est
1JOHN|3|4|omnis qui facit peccatum et iniquitatem facit et peccatum est iniquitas
1JOHN|3|5|et scitis quoniam ille apparuit ut peccata tolleret et peccatum in eo non est
1JOHN|3|6|omnis qui in eo manet non peccat omnis qui peccat non vidit eum nec cognovit eum
1JOHN|3|7|filioli nemo vos seducat qui facit iustitiam iustus est sicut et ille iustus est
1JOHN|3|8|qui facit peccatum ex diabolo est quoniam ab initio diabolus peccat in hoc apparuit Filius Dei ut dissolvat opera diaboli
1JOHN|3|9|omnis qui natus est ex Deo peccatum non facit quoniam semen ipsius in eo manet et non potest peccare quoniam ex Deo natus est
1JOHN|3|10|in hoc manifesti sunt filii Dei et filii diaboli omnis qui non est iustus non est de Deo et qui non diligit fratrem suum
1JOHN|3|11|quoniam haec est adnuntiatio quam audistis ab initio ut diligamus alterutrum
1JOHN|3|12|non sicut Cain ex maligno erat et occidit fratrem suum et propter quid occidit eum quoniam opera eius maligna erant fratris autem eius iusta
1JOHN|3|13|nolite mirari fratres si odit vos mundus
1JOHN|3|14|nos scimus quoniam translati sumus de morte in vitam quoniam diligimus fratres qui non diligit manet in morte
1JOHN|3|15|omnis qui odit fratrem suum homicida est et scitis quoniam omnis homicida non habet vitam aeternam in se manentem
1JOHN|3|16|in hoc cognovimus caritatem quoniam ille pro nobis animam suam posuit et nos debemus pro fratribus animas ponere
1JOHN|3|17|qui habuerit substantiam mundi et viderit fratrem suum necesse habere et clauserit viscera sua ab eo quomodo caritas Dei manet in eo
1JOHN|3|18|filioli non diligamus verbo nec lingua sed opere et veritate
1JOHN|3|19|in hoc cognoscimus quoniam ex veritate sumus et in conspectu eius suadeamus corda nostra
1JOHN|3|20|quoniam si reprehenderit nos cor maior est Deus corde nostro et novit omnia
1JOHN|3|21|carissimi si cor non reprehenderit nos fiduciam habemus ad Deum
1JOHN|3|22|et quodcumque petierimus accipiemus ab eo quoniam mandata eius custodimus et ea quae sunt placita coram eo facimus
1JOHN|3|23|et hoc est mandatum eius ut credamus in nomine Filii eius Iesu Christi et diligamus alterutrum sicut dedit mandatum nobis
1JOHN|3|24|et qui servat mandata eius in illo manet et ipse in eo et in hoc scimus quoniam manet in nobis de Spiritu quem nobis dedit
1JOHN|4|1|carissimi nolite omni spiritui credere sed probate spiritus si ex Deo sint quoniam multi pseudoprophetae exierunt in mundum
1JOHN|4|2|in hoc cognoscitur Spiritus Dei omnis spiritus qui confitetur Iesum Christum in carne venisse ex Deo est
1JOHN|4|3|et omnis spiritus qui solvit Iesum ex Deo non est et hoc est antichristi quod audistis quoniam venit et nunc iam in mundo est
1JOHN|4|4|vos ex Deo estis filioli et vicistis eos quoniam maior est qui in vobis est quam qui in mundo
1JOHN|4|5|ipsi de mundo sunt ideo de mundo loquuntur et mundus eos audit
1JOHN|4|6|nos ex Deo sumus qui novit Deum audit nos qui non est ex Deo non audit nos in hoc cognoscimus Spiritum veritatis et spiritum erroris
1JOHN|4|7|carissimi diligamus invicem quoniam caritas ex Deo est et omnis qui diligit ex Deo natus est et cognoscit Deum
1JOHN|4|8|qui non diligit non novit Deum quoniam Deus caritas est
1JOHN|4|9|in hoc apparuit caritas Dei in nobis quoniam Filium suum unigenitum misit Deus in mundum ut vivamus per eum
1JOHN|4|10|in hoc est caritas non quasi nos dilexerimus Deum sed quoniam ipse dilexit nos et misit Filium suum propitiationem pro peccatis nostris
1JOHN|4|11|carissimi si sic Deus dilexit nos et nos debemus alterutrum diligere
1JOHN|4|12|Deum nemo vidit umquam si diligamus invicem Deus in nobis manet et caritas eius in nobis perfecta est
1JOHN|4|13|in hoc intellegimus quoniam in eo manemus et ipse in nobis quoniam de Spiritu suo dedit nobis
1JOHN|4|14|et nos vidimus et testificamur quoniam Pater misit Filium salvatorem mundi
1JOHN|4|15|quisque confessus fuerit quoniam Iesus est Filius Dei Deus in eo manet et ipse in Deo
1JOHN|4|16|et nos cognovimus et credidimus caritati quam habet Deus in nobis Deus caritas est et qui manet in caritate in Deo manet et Deus in eo
1JOHN|4|17|in hoc perfecta est caritas nobiscum ut fiduciam habeamus in die iudicii quia sicut ille est et nos sumus in hoc mundo
1JOHN|4|18|timor non est in caritate sed perfecta caritas foras mittit timorem quoniam timor poenam habet qui autem timet non est perfectus in caritate
1JOHN|4|19|nos ergo diligamus quoniam Deus prior dilexit nos
1JOHN|4|20|si quis dixerit quoniam diligo Deum et fratrem suum oderit mendax est qui enim non diligit fratrem suum quem vidit Deum quem non vidit quomodo potest diligere
1JOHN|4|21|et hoc mandatum habemus ab eo ut qui diligit Deum diligat et fratrem suum
1JOHN|5|1|omnis qui credit quoniam Iesus est Christus ex Deo natus est et omnis qui diligit eum qui genuit diligit eum qui natus est ex eo
1JOHN|5|2|in hoc cognoscimus quoniam diligimus natos Dei cum Deum diligamus et mandata eius faciamus
1JOHN|5|3|haec est enim caritas Dei ut mandata eius custodiamus et mandata eius gravia non sunt
1JOHN|5|4|quoniam omne quod natum est ex Deo vincit mundum et haec est victoria quae vincit mundum fides nostra
1JOHN|5|5|quis est qui vincit mundum nisi qui credit quoniam Iesus est Filius Dei
1JOHN|5|6|hic est qui venit per aquam et sanguinem Iesus Christus non in aqua solum sed in aqua et sanguine et Spiritus est qui testificatur quoniam Christus est veritas
1JOHN|5|7|quia tres sunt qui testimonium dant
1JOHN|5|8|Spiritus et aqua et sanguis et tres unum sunt
1JOHN|5|9|si testimonium hominum accipimus testimonium Dei maius est quoniam hoc est testimonium Dei quod maius est quia testificatus est de Filio suo
1JOHN|5|10|qui credit in Filio Dei habet testimonium Dei in se qui non credit Filio mendacem facit eum quoniam non credidit in testimonio quod testificatus est Deus de Filio suo
1JOHN|5|11|et hoc est testimonium quoniam vitam aeternam dedit nobis Deus et haec vita in Filio eius est
1JOHN|5|12|qui habet Filium habet vitam qui non habet Filium Dei vitam non habet
1JOHN|5|13|haec scripsi vobis ut sciatis quoniam vitam habetis aeternam qui creditis in nomine Filii Dei
1JOHN|5|14|et haec est fiducia quam habemus ad eum quia quodcumque petierimus secundum voluntatem eius audit nos
1JOHN|5|15|et scimus quoniam audit nos quicquid petierimus scimus quoniam habemus petitiones quas postulavimus ab eo
1JOHN|5|16|qui scit fratrem suum peccare peccatum non ad mortem petet et dabit ei vitam peccantibus non ad mortem est peccatum ad mortem non pro illo dico ut roget
1JOHN|5|17|omnis iniquitas peccatum est et est peccatum non ad mortem
1JOHN|5|18|scimus quoniam omnis qui natus est ex Deo non peccat sed generatio Dei conservat eum et malignus non tangit eum
1JOHN|5|19|scimus quoniam ex Deo sumus et mundus totus in maligno positus est
1JOHN|5|20|et scimus quoniam Filius Dei venit et dedit nobis sensum ut cognoscamus verum Deum et simus in vero Filio eius hic est verus Deus et vita aeterna
1JOHN|5|21|filioli custodite vos a simulacris
2JOHN|1|1|senior electae dominae et natis eius quos ego diligo in veritate et non ego solus sed et omnes qui cognoverunt veritatem
2JOHN|1|2|propter veritatem quae permanet in nobis et nobiscum erit in aeternum
2JOHN|1|3|sit nobiscum gratia misericordia pax a Deo Patre et a Christo Iesu Filio Patris in veritate et caritate
2JOHN|1|4|gavisus sum valde quoniam inveni de filiis tuis ambulantes in veritate sicut mandatum accepimus a Patre
2JOHN|1|5|et nunc rogo te domina non tamquam mandatum novum scribens tibi sed quod habuimus ab initio ut diligamus alterutrum
2JOHN|1|6|et haec est caritas ut ambulemus secundum mandata eius hoc mandatum est ut quemadmodum audistis ab initio in eo ambuletis
2JOHN|1|7|quoniam multi seductores exierunt in mundum qui non confitentur Iesum Christum venientem in carne hic est seductor et antichristus
2JOHN|1|8|videte vosmet ipsos ne perdatis quae operati estis sed ut mercedem plenam accipiatis
2JOHN|1|9|omnis qui praecedit et non manet in doctrina Christi Deum non habet qui permanet in doctrina hic et Filium et Patrem habet
2JOHN|1|10|si quis venit ad vos et hanc doctrinam non adfert nolite recipere eum in domum nec have ei dixeritis
2JOHN|1|11|qui enim dicit illi have communicat operibus illius malignis
2JOHN|1|12|plura habens vobis scribere nolui per cartam et atramentum spero enim me futurum apud vos et os ad os loqui ut gaudium vestrum plenum sit
2JOHN|1|13|salutant te filii sororis tuae electae
3JOHN|1|1|senior Gaio carissimo quem ego diligo in veritate
3JOHN|1|2|carissime de omnibus orationem facio prospere te ingredi et valere sicut prospere agit anima tua
3JOHN|1|3|gavisus sum valde venientibus fratribus et testimonium perhibentibus veritati tuae sicut tu in veritate ambulas
3JOHN|1|4|maiorem horum non habeo gratiam quam ut audiam filios meos in veritate ambulantes
3JOHN|1|5|carissime fideliter facis quicquid operaris in fratres et hoc in peregrinos
3JOHN|1|6|qui testimonium reddiderunt caritati tuae in conspectu ecclesiae quos bene facies deducens digne Deo
3JOHN|1|7|pro nomine enim profecti sunt nihil accipientes a gentibus
3JOHN|1|8|nos ergo debemus suscipere huiusmodi ut cooperatores simus veritatis
3JOHN|1|9|scripsissem forsitan ecclesiae sed is qui amat primatum gerere in eis Diotrepes non recipit nos
3JOHN|1|10|propter hoc si venero commoneam eius opera quae facit verbis malignis garriens in nos et quasi non ei ista sufficiant nec ipse suscipit fratres et eos qui cupiunt prohibet et de ecclesia eicit
3JOHN|1|11|carissime noli imitari malum sed quod bonum est qui benefacit ex Deo est qui malefacit non vidit Deum
3JOHN|1|12|Demetrio testimonium redditur ab omnibus et ab ipsa veritate et nos autem testimonium perhibemus et nosti quoniam testimonium nostrum verum est
3JOHN|1|13|multa habui scribere tibi sed nolui per atramentum et calamum scribere tibi
3JOHN|1|14|spero autem protinus te videre et os ad os loquemur
3JOHN|1|15|pax tibi salutant te amici saluta amicos per nomen
JUDE|1|1|Iudas Iesu Christi servus frater autem Iacobi his qui in Deo Patre dilectis et Iesu Christo conservatis vocatis
JUDE|1|2|misericordia vobis et pax et caritas adimpleatur
JUDE|1|3|carissimi omnem sollicitudinem faciens scribendi vobis de communi vestra salute necesse habui scribere vobis deprecans supercertari semel traditae sanctis fidei
JUDE|1|4|subintroierunt enim quidam homines qui olim praescripti sunt in hoc iudicium impii Dei nostri gratiam transferentes in luxuriam et solum Dominatorem et Dominum nostrum Iesum Christum negantes
JUDE|1|5|commonere autem vos volo scientes semel omnia quoniam Iesus populum de terra Aegypti salvans secundo eos qui non crediderunt perdidit
JUDE|1|6|angelos vero qui non servaverunt suum principatum sed dereliquerunt suum domicilium in iudicium magni diei vinculis aeternis sub caligine reservavit
JUDE|1|7|sicut Sodoma et Gomorra et finitimae civitates simili modo exfornicatae et abeuntes post carnem alteram factae sunt exemplum ignis aeterni poenam sustinentes
JUDE|1|8|similiter et hii carnem quidem maculant dominationem autem spernunt maiestates autem blasphemant
JUDE|1|9|cum Michahel archangelus cum diabolo disputans altercaretur de Mosi corpore non est ausus iudicium inferre blasphemiae sed dixit imperet tibi Dominus
JUDE|1|10|hii autem quaecumque quidem ignorant blasphemant quaecumque autem naturaliter tamquam muta animalia norunt in his corrumpuntur
JUDE|1|11|vae illis quia via Cain abierunt et errore Balaam mercede effusi sunt et contradictione Core perierunt
JUDE|1|12|hii sunt in epulis suis maculae convivantes sine timore semet ipsos pascentes nubes sine aqua quae a ventis circumferuntur arbores autumnales infructuosae bis mortuae eradicatae
JUDE|1|13|fluctus feri maris despumantes suas confusiones sidera errantia quibus procella tenebrarum in aeternum servata est
JUDE|1|14|prophetavit autem et his septimus ab Adam Enoc dicens ecce venit Dominus in sanctis milibus suis
JUDE|1|15|facere iudicium contra omnes et arguere omnes impios de omnibus operibus impietatis eorum quibus impie egerunt et de omnibus duris quae locuti sunt contra eum peccatores impii
JUDE|1|16|hii sunt murmuratores querellosi secundum desideria sua ambulantes et os illorum loquitur superba mirantes personas quaestus causa
JUDE|1|17|vos autem carissimi memores estote verborum quae praedicta sunt ab apostolis Domini nostri Iesu Christi
JUDE|1|18|quia dicebant vobis quoniam in novissimo tempore venient inlusores secundum sua desideria ambulantes impietatum
JUDE|1|19|hii sunt qui segregant animales Spiritum non habentes
JUDE|1|20|vos autem carissimi superaedificantes vosmet ipsos sanctissimae vestrae fidei in Spiritu Sancto orantes
JUDE|1|21|ipsos vos in dilectione Dei servate
JUDE|1|22|et hos quidem arguite iudicatos
JUDE|1|23|illos vero salvate de igne rapientes aliis autem miseremini in timore odientes et eam quae carnalis est maculatam tunicam
JUDE|1|24|ei autem qui potest vos conservare sine peccato et constituere ante conspectum gloriae suae inmaculatos in exultatione
JUDE|1|25|soli Deo salvatori nostro per Iesum Christum Dominum nostrum gloria magnificentia imperium et potestas ante omne saeculum et nunc et in omnia saecula amen
REV|1|1|apocalypsis Iesu Christi quam dedit illi Deus palam facere servis suis quae oportet fieri cito et significavit mittens per angelum suum servo suo Iohanni
REV|1|2|qui testimonium perhibuit verbo Dei et testimonium Iesu Christi quaecumque vidit
REV|1|3|beatus qui legit et qui audiunt verba prophetiae et servant ea quae in ea scripta sunt tempus enim prope est
REV|1|4|Iohannes septem ecclesiis quae sunt in Asia gratia vobis et pax ab eo qui est et qui erat et qui venturus est et a septem spiritibus qui in conspectu throni eius sunt
REV|1|5|et ab Iesu Christo qui est testis fidelis primogenitus mortuorum et princeps regum terrae qui dilexit nos et lavit nos a peccatis nostris in sanguine suo
REV|1|6|et fecit nostrum regnum sacerdotes Deo et Patri suo ipsi gloria et imperium in saecula saeculorum amen
REV|1|7|ecce venit cum nubibus et videbit eum omnis oculus et qui eum pupugerunt et plangent se super eum omnes tribus terrae etiam amen
REV|1|8|ego sum Alpha et Omega principium et finis dicit Dominus Deus qui est et qui erat et qui venturus est Omnipotens
REV|1|9|ego Iohannes frater vester et particeps in tribulatione et regno et patientia in Iesu fui in insula quae appellatur Patmos propter verbum Dei et testimonium Iesu
REV|1|10|fui in spiritu in dominica die et audivi post me vocem magnam tamquam tubae
REV|1|11|dicentis quod vides scribe in libro et mitte septem ecclesiis Ephesum et Zmyrnam et Pergamum et Thyatiram et Sardis et Philadelphiam et Laodiciam
REV|1|12|et conversus sum ut viderem vocem quae loquebatur mecum et conversus vidi septem candelabra aurea
REV|1|13|et in medio septem candelabrorum similem Filio hominis vestitum podere et praecinctum ad mamillas zonam auream
REV|1|14|caput autem eius et capilli erant candidi tamquam lana alba tamquam nix et oculi eius velut flamma ignis
REV|1|15|et pedes eius similes orichalco sicut in camino ardenti et vox illius tamquam vox aquarum multarum
REV|1|16|et habebat in dextera sua stellas septem et de ore eius gladius utraque parte acutus exiebat et facies eius sicut sol lucet in virtute sua
REV|1|17|et cum vidissem eum cecidi ad pedes eius tamquam mortuus et posuit dexteram suam super me dicens noli timere ego sum primus et novissimus
REV|1|18|et vivus et fui mortuus et ecce sum vivens in saecula saeculorum et habeo claves mortis et inferni
REV|1|19|scribe ergo quae vidisti et quae sunt et quae oportet fieri post haec
REV|1|20|sacramentum septem stellarum quas vidisti in dextera mea et septem candelabra aurea septem stellae angeli sunt septem ecclesiarum et candelabra septem septem ecclesiae sunt
REV|2|1|angelo Ephesi ecclesiae scribe haec dicit qui tenet septem stellas in dextera sua qui ambulat in medio septem candelabrorum aureorum
REV|2|2|scio opera tua et laborem et patientiam tuam et quia non potes sustinere malos et temptasti eos qui se dicunt apostolos et non sunt et invenisti eos mendaces
REV|2|3|et patientiam habes et sustinuisti propter nomen meum et non defecisti
REV|2|4|sed habeo adversus te quod caritatem tuam primam reliquisti
REV|2|5|memor esto itaque unde excideris et age paenitentiam et prima opera fac sin autem venio tibi et movebo candelabrum tuum de loco suo nisi paenitentiam egeris
REV|2|6|sed hoc habes quia odisti facta Nicolaitarum quae et ego odi
REV|2|7|qui habet aurem audiat quid Spiritus dicat ecclesiis vincenti dabo ei edere de ligno vitae quod est in paradiso Dei mei
REV|2|8|et angelo Zmyrnae ecclesiae scribe haec dicit primus et novissimus qui fuit mortuus et vivit
REV|2|9|scio tribulationem tuam et paupertatem tuam sed dives es et blasphemaris ab his qui se dicunt Iudaeos esse et non sunt sed sunt synagoga Satanae
REV|2|10|nihil horum timeas quae passurus es ecce missurus est diabolus ex vobis in carcerem ut temptemini et habebitis tribulationem diebus decem esto fidelis usque ad mortem et dabo tibi coronam vitae
REV|2|11|qui habet aurem audiat quid Spiritus dicat ecclesiis qui vicerit non laedetur a morte secunda
REV|2|12|et angelo Pergami ecclesiae scribe haec dicit qui habet rompheam utraque parte acutam
REV|2|13|scio ubi habitas ubi sedes est Satanae et tenes nomen meum et non negasti fidem meam et in diebus Antipas testis meus fidelis qui occisus est apud vos ubi Satanas habitat
REV|2|14|sed habeo adversus te pauca quia habes illic tenentes doctrinam Balaam qui docebat Balac mittere scandalum coram filiis Israhel edere et fornicari
REV|2|15|ita habes et tu tenentes doctrinam Nicolaitarum
REV|2|16|similiter paenitentiam age si quo minus venio tibi cito et pugnabo cum illis in gladio oris mei
REV|2|17|qui habet aurem audiat quid Spiritus dicat ecclesiis vincenti dabo ei manna absconditum et dabo illi calculum candidum et in calculo nomen novum scriptum quod nemo scit nisi qui accipit
REV|2|18|et angelo Thyatirae ecclesiae scribe haec dicit Filius Dei qui habet oculos ut flammam ignis et pedes eius similes orichalco
REV|2|19|novi opera tua et caritatem et fidem et ministerium et patientiam tuam et opera tua novissima plura prioribus
REV|2|20|sed habeo adversus te quia permittis mulierem Hiezabel quae se dicit propheten docere et seducere servos meos fornicari et manducare de idolothytis
REV|2|21|et dedi illi tempus ut paenitentiam ageret et non vult paeniteri a fornicatione sua
REV|2|22|ecce mitto eam in lectum et qui moechantur cum ea in tribulationem maximam nisi paenitentiam egerint ab operibus eius
REV|2|23|et filios eius interficiam in morte et scient omnes ecclesiae quia ego sum scrutans renes et corda et dabo unicuique vestrum secundum opera vestra
REV|2|24|vobis autem dico ceteris qui Thyatirae estis quicumque non habent doctrinam hanc qui non cognoverunt altitudines Satanae quemadmodum dicunt non mittam super vos aliud pondus
REV|2|25|tamen id quod habetis tenete donec veniam
REV|2|26|et qui vicerit et qui custodierit usque in finem opera mea dabo illi potestatem super gentes
REV|2|27|et reget illas in virga ferrea tamquam vas figuli confringentur
REV|2|28|sicut et ego accepi a Patre meo et dabo illi stellam matutinam
REV|2|29|qui habet aurem audiat quid Spiritus dicat ecclesiis
REV|3|1|et angelo ecclesiae Sardis scribe haec dicit qui habet septem spiritus Dei et septem stellas scio opera tua quia nomen habes quod vivas et mortuus es
REV|3|2|esto vigilans et confirma cetera quae moritura erant non enim invenio opera tua plena coram Deo meo
REV|3|3|in mente ergo habe qualiter acceperis et audieris et serva et paenitentiam age si ergo non vigilaveris veniam tamquam fur et nescies qua hora veniam ad te
REV|3|4|sed habes pauca nomina in Sardis qui non inquinaverunt vestimenta sua et ambulabunt mecum in albis quia digni sunt
REV|3|5|qui vicerit sic vestietur vestimentis albis et non delebo nomen eius de libro vitae et confitebor nomen eius coram Patre meo et coram angelis eius
REV|3|6|qui habet aurem audiat quid Spiritus dicat ecclesiis
REV|3|7|et angelo Philadelphiae ecclesiae scribe haec dicit sanctus et verus qui habet clavem David qui aperit et nemo cludit et cludit et nemo aperit
REV|3|8|scio opera tua ecce dedi coram te ostium apertum quod nemo potest cludere quia modicam habes virtutem et servasti verbum meum et non negasti nomen meum
REV|3|9|ecce dabo de synagoga Satanae qui dicunt se Iudaeos esse et non sunt sed mentiuntur ecce faciam illos ut veniant et adorent ante pedes tuos et scient quia ego dilexi te
REV|3|10|quoniam servasti verbum patientiae meae et ego te servabo ab hora temptationis quae ventura est in orbem universum temptare habitantes in terra
REV|3|11|venio cito tene quod habes ut nemo accipiat coronam tuam
REV|3|12|qui vicerit faciam illum columnam in templo Dei mei et foras non egredietur amplius et scribam super eum nomen Dei mei et nomen civitatis Dei mei novae Hierusalem quae descendit de caelo a Deo meo et nomen meum novum
REV|3|13|qui habet aurem audiat quid Spiritus dicat ecclesiis
REV|3|14|et angelo Laodiciae ecclesiae scribe haec dicit Amen testis fidelis et verus qui est principium creaturae Dei
REV|3|15|scio opera tua quia neque frigidus es neque calidus utinam frigidus esses aut calidus
REV|3|16|sed quia tepidus es et nec frigidus nec calidus incipiam te evomere ex ore meo
REV|3|17|quia dicis quod dives sum et locupletatus et nullius egeo et nescis quia tu es miser et miserabilis et pauper et caecus et nudus
REV|3|18|suadeo tibi emere a me aurum ignitum probatum ut locuples fias et vestimentis albis induaris et non appareat confusio nuditatis tuae et collyrio inungue oculos tuos ut videas
REV|3|19|ego quos amo arguo et castigo aemulare ergo et paenitentiam age
REV|3|20|ecce sto ad ostium et pulso si quis audierit vocem meam et aperuerit ianuam introibo ad illum et cenabo cum illo et ipse mecum
REV|3|21|qui vicerit dabo ei sedere mecum in throno meo sicut et ego vici et sedi cum Patre meo in throno eius
REV|3|22|qui habet aurem audiat quid Spiritus dicat ecclesiis
REV|4|1|post haec vidi et ecce ostium apertum in caelo et vox prima quam audivi tamquam tubae loquentis mecum dicens ascende huc et ostendam tibi quae oportet fieri post haec
REV|4|2|statim fui in spiritu et ecce sedis posita erat in caelo et supra sedem sedens
REV|4|3|et qui sedebat similis erat aspectui lapidis iaspidis et sardini et iris erat in circuitu sedis similis visioni zmaragdinae
REV|4|4|et in circuitu sedis sedilia viginti quattuor et super thronos viginti quattuor seniores sedentes circumamictos vestimentis albis et in capitibus eorum coronas aureas
REV|4|5|et de throno procedunt fulgura et voces et tonitrua et septem lampades ardentes ante thronum quae sunt septem spiritus Dei
REV|4|6|et in conspectu sedis tamquam mare vitreum simile cristallo et in medio sedis et in circuitu sedis quattuor animalia plena oculis ante et retro
REV|4|7|et animal primum simile leoni et secundum animal simile vitulo et tertium animal habens faciem quasi hominis et quartum animal simile aquilae volanti
REV|4|8|et quattuor animalia singula eorum habebant alas senas et in circuitu et intus plena sunt oculis et requiem non habent die et nocte dicentia sanctus sanctus sanctus Dominus Deus omnipotens qui erat et qui est et qui venturus est
REV|4|9|et cum darent illa animalia gloriam et honorem et benedictionem sedenti super thronum viventi in saecula saeculorum
REV|4|10|procident viginti quattuor seniores ante sedentem in throno et adorabunt viventem in saecula saeculorum et mittent coronas suas ante thronum dicentes
REV|4|11|dignus es Domine et Deus noster accipere gloriam et honorem et virtutem quia tu creasti omnia et propter voluntatem tuam erant et creata sunt
REV|5|1|et vidi in dextera sedentis super thronum librum scriptum intus et foris signatum sigillis septem
REV|5|2|et vidi angelum fortem praedicantem voce magna quis est dignus aperire librum et solvere signacula eius
REV|5|3|et nemo poterat in caelo neque in terra neque subtus terram aperire librum neque respicere illum
REV|5|4|et ego flebam multum quoniam nemo dignus inventus est aperire librum nec videre eum
REV|5|5|et unus de senioribus dicit mihi ne fleveris ecce vicit leo de tribu Iuda radix David aperire librum et septem signacula eius
REV|5|6|et vidi et ecce in medio throni et quattuor animalium et in medio seniorum agnum stantem tamquam occisum habentem cornua septem et oculos septem qui sunt spiritus Dei missi in omnem terram
REV|5|7|et venit et accepit de dextera sedentis de throno
REV|5|8|et cum aperuisset librum quattuor animalia et viginti quattuor seniores ceciderunt coram agno habentes singuli citharas et fialas aureas plenas odoramentorum quae sunt orationes sanctorum
REV|5|9|et cantant novum canticum dicentes dignus es accipere librum et aperire signacula eius quoniam occisus es et redemisti nos Deo in sanguine tuo ex omni tribu et lingua et populo et natione
REV|5|10|et fecisti eos Deo nostro regnum et sacerdotes et regnabunt super terram
REV|5|11|et vidi et audivi vocem angelorum multorum in circuitu throni et animalium et seniorum et erat numerus eorum milia milium
REV|5|12|dicentium voce magna dignus est agnus qui occisus est accipere virtutem et divinitatem et sapientiam et fortitudinem et honorem et gloriam et benedictionem
REV|5|13|et omnem creaturam quae in caelo est et super terram et sub terram et quae sunt in mari et quae in ea omnes audivi dicentes sedenti in throno et agno benedictio et honor et gloria et potestas in saecula saeculorum
REV|5|14|et quattuor animalia dicebant amen et seniores ceciderunt et adoraverunt
REV|6|1|et vidi quod aperuisset agnus unum de septem signaculis et audivi unum de quattuor animalibus dicentem tamquam vocem tonitrui veni
REV|6|2|et vidi et ecce equus albus et qui sedebat super illum habebat arcum et data est ei corona et exivit vincens ut vinceret
REV|6|3|et cum aperuisset sigillum secundum audivi secundum animal dicens veni
REV|6|4|et exivit alius equus rufus et qui sedebat super illum datum est ei ut sumeret pacem de terra et ut invicem se interficiant et datus est illi gladius magnus
REV|6|5|et cum aperuisset sigillum tertium audivi tertium animal dicens veni et vidi et ecce equus niger et qui sedebat super eum habebat stateram in manu sua
REV|6|6|et audivi tamquam vocem in medio quattuor animalium dicentem bilibris tritici denario et tres bilibres hordei denario et vinum et oleum ne laeseris
REV|6|7|et cum aperuisset sigillum quartum audivi vocem quarti animalis dicentis veni et vidi
REV|6|8|et ecce equus pallidus et qui sedebat desuper nomen illi Mors et inferus sequebatur eum et data est illi potestas super quattuor partes terrae interficere gladio fame et morte et bestiis terrae
REV|6|9|et cum aperuisset quintum sigillum vidi subtus altare animas interfectorum propter verbum Dei et propter testimonium quod habebant
REV|6|10|et clamabant voce magna dicentes usquequo Domine sanctus et verus non iudicas et vindicas sanguinem nostrum de his qui habitant in terra
REV|6|11|et datae sunt illis singulae stolae albae et dictum est illis ut requiescerent tempus adhuc modicum donec impleantur conservi eorum et fratres eorum qui interficiendi sunt sicut et illi
REV|6|12|et vidi cum aperuisset sigillum sextum et terraemotus factus est magnus et sol factus est niger tamquam saccus cilicinus et luna tota facta est sicut sanguis
REV|6|13|et stellae caeli ceciderunt super terram sicut ficus mittit grossos suos cum vento magno movetur
REV|6|14|et caelum recessit sicut liber involutus et omnis mons et insulae de locis suis motae sunt
REV|6|15|et reges terrae et principes et tribuni et divites et fortes et omnis servus et liber absconderunt se in speluncis et petris montium
REV|6|16|et dicunt montibus et petris cadite super nos et abscondite nos a facie sedentis super thronum et ab ira agni
REV|6|17|quoniam venit dies magnus irae ipsorum et quis poterit stare
REV|7|1|post haec vidi quattuor angelos stantes super quattuor angulos terrae tenentes quattuor ventos terrae ne flaret ventus super terram neque super mare neque in ullam arborem
REV|7|2|et vidi alterum angelum ascendentem ab ortu solis habentem signum Dei vivi et clamavit voce magna quattuor angelis quibus datum est nocere terrae et mari
REV|7|3|dicens nolite nocere terrae neque mari neque arboribus quoadusque signemus servos Dei nostri in frontibus eorum
REV|7|4|et audivi numerum signatorum centum quadraginta quattuor milia signati ex omni tribu filiorum Israhel
REV|7|5|ex tribu Iuda duodecim milia signati ex tribu Ruben duodecim milia ex tribu Gad duodecim milia
REV|7|6|ex tribu Aser duodecim milia ex tribu Nepthalim duodecim milia ex tribu Manasse duodecim milia
REV|7|7|ex tribu Symeon duodecim milia ex tribu Levi duodecim milia ex tribu Issachar duodecim milia
REV|7|8|ex tribu Zabulon duodecim milia ex tribu Ioseph duodecim milia ex tribu Beniamin duodecim milia signati
REV|7|9|post haec vidi turbam magnam quam dinumerare nemo poterat ex omnibus gentibus et tribubus et populis et linguis stantes ante thronum et in conspectu agni amicti stolas albas et palmae in manibus eorum
REV|7|10|et clamabant voce magna dicentes salus Deo nostro qui sedet super thronum et agno
REV|7|11|et omnes angeli stabant in circuitu throni et seniorum et quattuor animalium et ceciderunt in conspectu throni in facies suas et adoraverunt Deum
REV|7|12|dicentes amen benedictio et claritas et sapientia et gratiarum actio et honor et virtus et fortitudo Deo nostro in saecula saeculorum amen
REV|7|13|et respondit unus de senioribus dicens mihi hii qui amicti sunt stolis albis qui sunt et unde venerunt
REV|7|14|et dixi illi domine mi tu scis et dixit mihi hii sunt qui veniunt de tribulatione magna et laverunt stolas suas et dealbaverunt eas in sanguine agni
REV|7|15|ideo sunt ante thronum Dei et serviunt ei die ac nocte in templo eius et qui sedet in throno habitabit super illos
REV|7|16|non esurient neque sitient amplius neque cadet super illos sol neque ullus aestus
REV|7|17|quoniam agnus qui in medio throni est reget illos et deducet eos ad vitae fontes aquarum et absterget Deus omnem lacrimam ex oculis eorum
REV|8|1|et cum aperuisset sigillum septimum factum est silentium in caelo quasi media hora
REV|8|2|et vidi septem angelos stantes in conspectu Dei et datae sunt illis septem tubae
REV|8|3|et alius angelus venit et stetit ante altare habens turibulum aureum et data sunt illi incensa multa ut daret orationibus sanctorum omnium super altare aureum quod est ante thronum
REV|8|4|et ascendit fumus incensorum de orationibus sanctorum de manu angeli coram Deo
REV|8|5|et accepit angelus turibulum et implevit illud de igne altaris et misit in terram et facta sunt tonitrua et voces et fulgora et terraemotus
REV|8|6|et septem angeli qui habebant septem tubas paraverunt se ut tuba canerent
REV|8|7|et primus tuba cecinit et facta est grando et ignis mixta in sanguine et missum est in terram et tertia pars terrae conbusta est et tertia pars arborum conbusta est et omne faenum viride conbustum est
REV|8|8|et secundus angelus tuba cecinit et tamquam mons magnus igne ardens missus est in mare et facta est tertia pars maris sanguis
REV|8|9|et mortua est tertia pars creaturae quae habent animas et tertia pars navium interiit
REV|8|10|et tertius angelus tuba cecinit et cecidit de caelo stella magna ardens tamquam facula et cecidit in tertiam partem fluminum et in fontes aquarum
REV|8|11|et nomen stellae dicitur Absinthius et facta est tertia pars aquarum in absinthium et multi hominum mortui sunt de aquis quia amarae factae sunt
REV|8|12|et quartus angelus tuba cecinit et percussa est tertia pars solis et tertia pars lunae et tertia pars stellarum ut obscuraretur tertia pars eorum et diei non luceret pars tertia et nox similiter
REV|8|13|et vidi et audivi vocem unius aquilae volantis per medium caelum dicentis voce magna vae vae vae habitantibus in terra de ceteris vocibus tubae trium angelorum qui erant tuba canituri
REV|9|1|et quintus angelus tuba cecinit et vidi stellam de caelo cecidisse in terram et data est illi clavis putei abyssi
REV|9|2|et aperuit puteum abyssi et ascendit fumus putei sicut fumus fornacis magnae et obscuratus est sol et aer de fumo putei
REV|9|3|et de fumo exierunt lucustae in terram et data est illis potestas sicut habent potestatem scorpiones terrae
REV|9|4|et praeceptum est illis ne laederent faenum terrae neque omne viride neque omnem arborem nisi tantum homines qui non habent signum Dei in frontibus
REV|9|5|et datum est illis ne occiderent eos sed ut cruciarentur mensibus quinque et cruciatus eorum ut cruciatus scorpii cum percutit hominem
REV|9|6|et in diebus illis quaerent homines mortem et non invenient eam et desiderabunt mori et fugiet mors ab ipsis
REV|9|7|et similitudines lucustarum similes equis paratis in proelium et super capita earum tamquam coronae similes auro et facies earum sicut facies hominum
REV|9|8|et habebant capillos sicut capillos mulierum et dentes earum sicut leonum erant
REV|9|9|et habebant loricas sicut loricas ferreas et vox alarum earum sicut vox curruum equorum multorum currentium in bellum
REV|9|10|et habebant caudas similes scorpionum et aculei in caudis earum potestas earum nocere hominibus mensibus quinque
REV|9|11|et habebant super se regem angelum abyssi cui nomen hebraice Abaddon graece autem Apollyon et latine habet nomen Exterminans
REV|9|12|vae unum abiit ecce veniunt adhuc duo vae post haec
REV|9|13|et sextus angelus tuba cecinit et audivi vocem unum ex cornibus altaris aurei quod est ante oculos Dei
REV|9|14|dicentem sexto angelo qui habebat tubam solve quattuor angelos qui alligati sunt in flumine magno Eufrate
REV|9|15|et soluti sunt quattuor angeli qui parati erant in horam et diem et mensem et annum ut occiderent tertiam partem hominum
REV|9|16|et numerus equestris exercitus vicies milies dena milia audivi numerum eorum
REV|9|17|et ita vidi equos in visione et qui sedebant super eos habentes loricas igneas et hyacinthinas et sulphureas et capita equorum erant tamquam capita leonum et de ore ipsorum procedit ignis et fumus et sulphur
REV|9|18|ab his tribus plagis occisa est tertia pars hominum de igne et fumo et sulphure qui procedebat ex ore ipsorum
REV|9|19|potestas enim equorum in ore eorum est et in caudis eorum nam caudae illorum similes serpentibus habentes capita et in his nocent
REV|9|20|et ceteri homines qui non sunt occisi in his plagis neque paenitentiam egerunt de operibus manuum suarum ut non adorarent daemonia et simulacra aurea et argentea et aerea et lapidea et lignea quae neque videre possunt neque audire neque ambulare
REV|9|21|et non egerunt paenitentiam ab homicidiis suis neque a veneficiis suis neque a fornicatione sua neque a furtis suis
REV|10|1|et vidi alium angelum fortem descendentem de caelo amictum nube et iris in capite eius et facies eius erat ut sol et pedes eius tamquam columna ignis
REV|10|2|et habebat in manu sua libellum apertum et posuit pedem suum dextrum supra mare sinistrum autem super terram
REV|10|3|et clamavit voce magna quemadmodum cum leo rugit et cum clamasset locuta sunt septem tonitrua voces suas
REV|10|4|et cum locuta fuissent septem tonitrua scripturus eram et audivi vocem de caelo dicentem signa quae locuta sunt septem tonitrua et noli ea scribere
REV|10|5|et angelum quem vidi stantem supra mare et supra terram levavit manum suam ad caelum
REV|10|6|et iuravit per viventem in saecula saeculorum qui creavit caelum et ea quae in illo sunt et terram et ea quae in ea sunt et mare et quae in eo sunt quia tempus amplius non erit
REV|10|7|sed in diebus vocis septimi angeli cum coeperit tuba canere et consummabitur mysterium Dei sicut evangelizavit per servos suos prophetas
REV|10|8|et vox quam audivi de caelo iterum loquentem mecum et dicentem vade accipe librum apertum de manu angeli stantis supra mare et supra terram
REV|10|9|et abii ad angelum dicens ei ut daret mihi librum et dicit mihi accipe et devora illum et faciet amaricare ventrem tuum sed in ore tuo erit dulce tamquam mel
REV|10|10|et accepi librum de manu angeli et devoravi eum et erat in ore meo tamquam mel dulce et cum devorassem eum amaricatus est venter meus
REV|10|11|et dicunt mihi oportet te iterum prophetare populis et gentibus et linguis et regibus multis
REV|11|1|et datus est mihi calamus similis virgae dicens surge et metire templum Dei et altare et adorantes in eo
REV|11|2|atrium autem quod est foris templum eice foras et ne metieris eum quoniam datum est gentibus et civitatem sanctam calcabunt mensibus quadraginta duobus
REV|11|3|et dabo duobus testibus meis et prophetabunt diebus mille ducentis sexaginta amicti saccos
REV|11|4|hii sunt duo olivae et duo candelabra in conspectu Domini terrae stantes
REV|11|5|et si quis eos voluerit nocere ignis exiet de ore illorum et devorabit inimicos eorum et si quis voluerit eos laedere sic oportet eum occidi
REV|11|6|hii habent potestatem cludendi caelum ne pluat diebus prophetiae ipsorum et potestatem habent super aquas convertendi eas in sanguinem et percutere terram omni plaga quotienscumque voluerint
REV|11|7|et cum finierint testimonium suum bestia quae ascendit de abysso faciet adversus illos bellum et vincet eos et occidet illos
REV|11|8|et corpora eorum in plateis civitatis magnae quae vocatur spiritaliter Sodoma et Aegyptus ubi et Dominus eorum crucifixus est
REV|11|9|et videbunt de populis et tribubus et linguis et gentibus corpora eorum per tres dies et dimidium et corpora eorum non sinunt poni in monumentis
REV|11|10|et inhabitantes terram gaudebunt super illis et iucundabuntur et munera mittent invicem quoniam hii duo prophetae cruciaverunt eos qui inhabitant super terram
REV|11|11|et post dies tres et dimidium spiritus vitae a Deo intravit in eos et steterunt super pedes suos et timor magnus cecidit super eos qui viderunt eos
REV|11|12|et audierunt vocem magnam de caelo dicentem illis ascendite huc et ascenderunt in caelum in nube et viderunt illos inimici eorum
REV|11|13|et in illa hora factus est terraemotus magnus et decima pars civitatis cecidit et occisi sunt in terraemotu nomina hominum septem milia et reliqui in timore sunt missi et dederunt gloriam Deo caeli
REV|11|14|vae secundum abiit ecce vae tertium veniet cito
REV|11|15|et septimus angelus tuba cecinit et factae sunt voces magnae in caelo dicentes factum est regnum huius mundi Domini nostri et Christi eius et regnabit in saecula saeculorum
REV|11|16|et viginti quattuor seniores qui in conspectu Dei sedent in sedibus suis ceciderunt in facies suas et adoraverunt Deum
REV|11|17|dicentes gratias agimus tibi Domine Deus omnipotens qui es et qui eras quia accepisti virtutem tuam magnam et regnasti
REV|11|18|et iratae sunt gentes et advenit ira tua et tempus mortuorum iudicari et reddere mercedem servis tuis prophetis et sanctis et timentibus nomen tuum pusillis et magnis et exterminandi eos qui corruperunt terram
REV|11|19|et apertum est templum Dei in caelo et visa est arca testamenti eius in templo eius et facta sunt fulgora et voces et terraemotus et grando magna
REV|12|1|et signum magnum paruit in caelo mulier amicta sole et luna sub pedibus eius et in capite eius corona stellarum duodecim
REV|12|2|et in utero habens et clamat parturiens et cruciatur ut pariat
REV|12|3|et visum est aliud signum in caelo et ecce draco magnus rufus habens capita septem et cornua decem et in capitibus suis septem diademata
REV|12|4|et cauda eius trahebat tertiam partem stellarum caeli et misit eas in terram et draco stetit ante mulierem quae erat paritura ut cum peperisset filium eius devoraret
REV|12|5|et peperit filium masculum qui recturus erit omnes gentes in virga ferrea et raptus est filius eius ad Deum et ad thronum eius
REV|12|6|et mulier fugit in solitudinem ubi habet locum paratum a Deo ut ibi pascant illam diebus mille ducentis sexaginta
REV|12|7|et factum est proelium in caelo Michahel et angeli eius proeliabantur cum dracone et draco pugnabat et angeli eius
REV|12|8|et non valuerunt neque locus inventus est eorum amplius in caelo
REV|12|9|et proiectus est draco ille magnus serpens antiquus qui vocatur Diabolus et Satanas qui seducit universum orbem proiectus est in terram et angeli eius cum illo missi sunt
REV|12|10|et audivi vocem magnam in caelo dicentem nunc facta est salus et virtus et regnum Dei nostri et potestas Christi eius quia proiectus est accusator fratrum nostrorum qui accusabat illos ante conspectum Dei nostri die ac nocte
REV|12|11|et ipsi vicerunt illum propter sanguinem agni et propter verbum testimonii sui et non dilexerunt animam suam usque ad mortem
REV|12|12|propterea laetamini caeli et qui habitatis in eis vae terrae et mari quia descendit diabolus ad vos habens iram magnam sciens quod modicum tempus habet
REV|12|13|et postquam vidit draco quod proiectus est in terram persecutus est mulierem quae peperit masculum
REV|12|14|et datae sunt mulieri duae alae aquilae magnae ut volaret in desertum in locum suum ubi alitur per tempus et tempora et dimidium temporis a facie serpentis
REV|12|15|et misit serpens ex ore suo post mulierem aquam tamquam flumen ut eam faceret trahi a flumine
REV|12|16|et adiuvit terra mulierem et aperuit terra os suum et absorbuit flumen quod misit draco de ore suo
REV|12|17|et iratus est draco in mulierem et abiit facere proelium cum reliquis de semine eius qui custodiunt mandata Dei et habent testimonium Iesu
REV|12|18|et stetit super harenam maris
REV|13|1|et vidi de mare bestiam ascendentem habentem capita septem et cornua decem et super cornua eius decem diademata et super capita eius nomina blasphemiae
REV|13|2|et bestiam quam vidi similis erat pardo et pedes eius sicut ursi et os eius sicut os leonis et dedit illi draco virtutem suam et potestatem magnam
REV|13|3|et unum de capitibus suis quasi occisum in mortem et plaga mortis eius curata est et admirata est universa terra post bestiam
REV|13|4|et adoraverunt draconem quia dedit potestatem bestiae et adoraverunt bestiam dicentes quis similis bestiae et quis poterit pugnare cum ea
REV|13|5|et datum est ei os loquens magna et blasphemiae et data est illi potestas facere menses quadraginta duo
REV|13|6|et aperuit os suum in blasphemias ad Deum blasphemare nomen eius et tabernaculum eius et eos qui in caelo habitant
REV|13|7|et datum est illi bellum facere cum sanctis et vincere illos et data est ei potestas in omnem tribum et populum et linguam et gentem
REV|13|8|et adorabunt eum omnes qui inhabitant terram quorum non sunt scripta nomina in libro vitae agni qui occisus est ab origine mundi
REV|13|9|si quis habet aurem audiat
REV|13|10|qui in captivitatem in captivitatem vadit qui in gladio occiderit oportet eum gladio occidi hic est patientia et fides sanctorum
REV|13|11|et vidi aliam bestiam ascendentem de terra et habebat cornua duo similia agni et loquebatur sicut draco
REV|13|12|et potestatem prioris bestiae omnem faciebat in conspectu eius et facit terram et inhabitantes in eam adorare bestiam primam cuius curata est plaga mortis
REV|13|13|et fecit signa magna ut etiam ignem faceret de caelo descendere in terram in conspectu hominum
REV|13|14|et seducit habitantes terram propter signa quae data sunt illi facere in conspectu bestiae dicens habitantibus in terra ut faciant imaginem bestiae quae habet plagam gladii et vixit
REV|13|15|et datum est illi ut daret spiritum imagini bestiae ut et loquatur imago bestiae et faciat quicumque non adoraverint imaginem bestiae occidantur
REV|13|16|et faciet omnes pusillos et magnos et divites et pauperes et liberos et servos habere caracter in dextera manu aut in frontibus suis
REV|13|17|et ne quis possit emere aut vendere nisi qui habet caracter nomen bestiae aut numerum nominis eius
REV|13|18|hic sapientia est qui habet intellectum conputet numerum bestiae numerus enim hominis est et numerus eius est sescenti sexaginta sex
REV|14|1|et vidi et ecce agnus stabat supra montem Sion et cum illo centum quadraginta quattuor milia habentes nomen eius et nomen Patris eius scriptum in frontibus suis
REV|14|2|et audivi vocem de caelo tamquam vocem aquarum multarum et tamquam vocem tonitrui magni et vocem quam audivi sicut citharoedorum citharizantium in citharis suis
REV|14|3|et cantabant quasi canticum novum ante sedem et ante quattuor animalia et seniores et nemo poterat discere canticum nisi illa centum quadraginta quattuor milia qui empti sunt de terra
REV|14|4|hii sunt qui cum mulieribus non sunt coinquinati virgines enim sunt hii qui sequuntur agnum quocumque abierit hii empti sunt ex hominibus primitiae Deo et agno
REV|14|5|et in ore ipsorum non est inventum mendacium sine macula sunt
REV|14|6|et vidi alterum angelum volantem per medium caelum habentem evangelium aeternum ut evangelizaret sedentibus super terram et super omnem gentem et tribum et linguam et populum
REV|14|7|dicens magna voce timete Deum et date illi honorem quia venit hora iudicii eius et adorate eum qui fecit caelum et terram et mare et fontes aquarum
REV|14|8|et alius angelus secutus est dicens cecidit cecidit Babylon illa magna quae a vino irae fornicationis suae potionavit omnes gentes
REV|14|9|et alius angelus tertius secutus est illos dicens voce magna si quis adoraverit bestiam et imaginem eius et acceperit caracterem in fronte sua aut in manu sua
REV|14|10|et hic bibet de vino irae Dei qui mixtus est mero in calice irae ipsius et cruciabitur igne et sulphure in conspectu angelorum sanctorum et ante conspectum agni
REV|14|11|et fumus tormentorum eorum in saecula saeculorum ascendit nec habent requiem die ac nocte qui adoraverunt bestiam et imaginem eius et si quis acceperit caracterem nominis eius
REV|14|12|hic patientia sanctorum est qui custodiunt mandata Dei et fidem Iesu
REV|14|13|et audivi vocem de caelo dicentem scribe beati mortui qui in Domino moriuntur amodo iam dicit Spiritus ut requiescant a laboribus suis opera enim illorum sequuntur illos
REV|14|14|et vidi et ecce nubem candidam et supra nubem sedentem similem Filio hominis habentem in capite suo coronam auream et in manu sua falcem acutam
REV|14|15|et alter angelus exivit de templo clamans voce magna ad sedentem super nubem mitte falcem tuam et mete quia venit hora ut metatur quoniam aruit messis terrae
REV|14|16|et misit qui sedebat supra nubem falcem suam in terram et messa est terra
REV|14|17|et alius angelus exivit de templo quod est in caelo habens et ipse falcem acutam
REV|14|18|et alius angelus de altari qui habet potestatem supra ignem et clamavit voce magna qui habebat falcem acutam dicens mitte falcem tuam acutam et vindemia botros vineae terrae quoniam maturae sunt uvae eius
REV|14|19|et misit angelus falcem suam in terram et vindemiavit vineam terrae et misit in lacum irae Dei magnum
REV|14|20|et calcatus est lacus extra civitatem et exivit sanguis de lacu usque ad frenos equorum per stadia mille sescenta
REV|15|1|et vidi aliud signum in caelo magnum et mirabile angelos septem habentes plagas septem novissimas quoniam in illis consummata est ira Dei
REV|15|2|et vidi tamquam mare vitreum mixtum igne et eos qui vicerunt bestiam et imaginem illius et numerum nominis eius stantes supra mare vitreum habentes citharas Dei
REV|15|3|et cantant canticum Mosi servi Dei et canticum agni dicentes magna et mirabilia opera tua Domine Deus omnipotens iustae et verae viae tuae rex saeculorum
REV|15|4|quis non timebit Domine et magnificabit nomen tuum quia solus pius quoniam omnes gentes venient et adorabunt in conspectu tuo quoniam iudicia tua manifestata sunt
REV|15|5|et post haec vidi et ecce apertum est templum tabernaculi testimonii in caelo
REV|15|6|et exierunt septem angeli habentes septem plagas de templo vestiti lapide mundo candido et praecincti circa pectora zonis aureis
REV|15|7|et unus ex quattuor animalibus dedit septem angelis septem fialas aureas plenas iracundiae Dei viventis in saecula saeculorum
REV|15|8|et impletum est templum fumo a maiestate Dei et de virtute eius et nemo poterat introire in templum donec consummarentur septem plagae septem angelorum
REV|16|1|et audivi vocem magnam de templo dicentem septem angelis ite et effundite septem fialas irae Dei in terram
REV|16|2|et abiit primus et effudit fialam suam in terram et factum est vulnus saevum ac pessimum in homines qui habent caracterem bestiae et eos qui adoraverunt imaginem eius
REV|16|3|et secundus effudit fialam suam in mare et factus est sanguis tamquam mortui et omnis anima vivens mortua est in mari
REV|16|4|et tertius effudit fialam suam super flumina et super fontes aquarum et factus est sanguis
REV|16|5|et audivi angelum aquarum dicentem iustus es qui es et qui eras sanctus quia haec iudicasti
REV|16|6|quia sanguinem sanctorum et prophetarum fuderunt et sanguinem eis dedisti bibere digni sunt
REV|16|7|et audivi altare dicens etiam Domine Deus omnipotens vera et iusta iudicia tua
REV|16|8|et quartus effudit fialam suam in solem et datum est illi aestu adficere homines et igni
REV|16|9|et aestuaverunt homines aestu magno et blasphemaverunt nomen Dei habentis potestatem super has plagas neque egerunt paenitentiam ut darent illi gloriam
REV|16|10|et quintus effudit fialam suam super sedem bestiae et factum est regnum eius tenebrosum et conmanducaverunt linguas suas prae dolore
REV|16|11|et blasphemaverunt Deum caeli prae doloribus et vulneribus suis et non egerunt paenitentiam ex operibus suis
REV|16|12|et sextus effudit fialam suam in flumen illud magnum Eufraten et siccavit aquam eius ut praepararetur via regibus ab ortu solis
REV|16|13|et vidi de ore draconis et de ore bestiae et de ore pseudoprophetae spiritus tres inmundos in modum ranarum
REV|16|14|sunt enim spiritus daemoniorum facientes signa et procedunt ad reges totius terrae congregare illos in proelium ad diem magnum Dei omnipotentis
REV|16|15|ecce venio sicut fur beatus qui vigilat et custodit vestimenta sua ne nudus ambulet et videant turpitudinem eius
REV|16|16|et congregavit illos in locum qui vocatur hebraice Hermagedon
REV|16|17|et septimus effudit fialam suam in aerem et exivit vox magna de templo a throno dicens factum est
REV|16|18|et facta sunt fulgora et voces et tonitrua et terraemotus factus est magnus qualis numquam fuit ex quo homines fuerunt super terram talis terraemotus sic magnus
REV|16|19|et facta est civitas magna in tres partes et civitates gentium ceciderunt et Babylon magna venit in memoriam ante Deum dare ei calicem vini indignationis irae eius
REV|16|20|et omnis insula fugit et montes non sunt inventi
REV|16|21|et grando magna sicut talentum descendit de caelo in homines et blasphemaverunt homines Deum propter plagam grandinis quoniam magna facta est vehementer
REV|17|1|et venit unus de septem angelis qui habebant septem fialas et locutus est mecum dicens veni ostendam tibi damnationem meretricis magnae quae sedet super aquas multas
REV|17|2|cum qua fornicati sunt reges terrae et inebriati sunt qui inhabitant terram de vino prostitutionis eius
REV|17|3|et abstulit me in desertum in spiritu et vidi mulierem sedentem super bestiam coccineam plenam nominibus blasphemiae habentem capita septem et cornua decem
REV|17|4|et mulier erat circumdata purpura et coccino et inaurata auro et lapide pretioso et margaritis habens poculum aureum in manu sua plenum abominationum et inmunditia fornicationis eius
REV|17|5|et in fronte eius nomen scriptum mysterium Babylon magna mater fornicationum et abominationum terrae
REV|17|6|et vidi mulierem ebriam de sanguine sanctorum et de sanguine martyrum Iesu et miratus sum cum vidissem illam admiratione magna
REV|17|7|et dixit mihi angelus quare miraris ego tibi dicam sacramentum mulieris et bestiae quae portat eam quae habet capita septem et decem cornua
REV|17|8|bestiam quam vidisti fuit et non est et ascensura est de abysso et in interitum ibit et mirabuntur inhabitantes terram quorum non sunt scripta nomina in libro vitae a constitutione mundi videntes bestiam quia erat et non est
REV|17|9|et hic est sensus qui habet sapientiam septem capita septem montes sunt super quos mulier sedet et reges septem sunt
REV|17|10|quinque ceciderunt unus est alius nondum venit et cum venerit oportet illum breve tempus manere
REV|17|11|et bestia quae erat et non est et ipsa octava est et de septem est et in interitum vadit
REV|17|12|et decem cornua quae vidisti decem reges sunt qui regnum nondum acceperunt sed potestatem tamquam reges una hora accipiunt post bestiam
REV|17|13|hii unum consilium habent et virtutem et potestatem suam bestiae tradunt
REV|17|14|hii cum agno pugnabunt et agnus vincet illos quoniam Dominus dominorum est et rex regum et qui cum illo sunt vocati et electi et fideles
REV|17|15|et dixit mihi aquas quas vidisti ubi meretrix sedet populi sunt et gentes et linguae
REV|17|16|et decem cornua quae vidisti et bestiam hii odient fornicariam et desolatam facient illam et nudam et carnes eius manducabunt et ipsam igni concremabunt
REV|17|17|Deus enim dedit in corda eorum ut faciant quod illi placitum est ut dent regnum suum bestiae donec consummentur verba Dei
REV|17|18|et mulier quam vidisti est civitas magna quae habet regnum super reges terrae
REV|18|1|et post haec vidi alium angelum descendentem de caelo habentem potestatem magnam et terra inluminata est a gloria eius
REV|18|2|et exclamavit in forti voce dicens cecidit cecidit Babylon magna et facta est habitatio daemoniorum et custodia omnis spiritus inmundi et custodia omnis volucris inmundae
REV|18|3|quia de ira fornicationis eius biberunt omnes gentes et reges terrae cum illa fornicati sunt et mercatores terrae de virtute deliciarum eius divites facti sunt
REV|18|4|et audivi aliam vocem de caelo dicentem exite de illa populus meus ut ne participes sitis delictorum eius et de plagis eius non accipiatis
REV|18|5|quoniam pervenerunt peccata eius usque ad caelum et recordatus est Deus iniquitatum eius
REV|18|6|reddite illi sicut ipsa reddidit et duplicate duplicia secundum opera eius in poculo quo miscuit miscite illi duplum
REV|18|7|quantum glorificavit se et in deliciis fuit tantum date illi tormentum et luctum quia in corde suo dicit sedeo regina et vidua non sum et luctum non videbo
REV|18|8|ideo in una die venient plagae eius mors et luctus et fames et igni conburetur quia fortis est Deus qui iudicavit illam
REV|18|9|et flebunt et plangent se super illam reges terrae qui cum illa fornicati sunt et in deliciis vixerunt cum viderint fumum incendii eius
REV|18|10|longe stantes propter timorem tormentorum eius dicentes vae vae civitas illa magna Babylon civitas illa fortis quoniam una hora venit iudicium tuum
REV|18|11|et negotiatores terrae flebunt et lugebunt super illam quoniam merces eorum nemo emet amplius
REV|18|12|mercem auri et argenti et lapidis pretiosi et margaritis et byssi et purpurae et serici et cocci et omne lignum thyinum et omnia vasa eboris et omnia vasa de lapide pretioso et aeramento et ferro et marmore
REV|18|13|et cinnamomum et amomum et odoramentorum et unguenti et turis et vini et olei et similae et tritici et iumentorum et ovium et equorum et raedarum et mancipiorum et animarum hominum
REV|18|14|et poma tua desiderii animae discessit a te et omnia pinguia et clara perierunt a te et amplius illa iam non invenient
REV|18|15|mercatores horum qui divites facti sunt ab ea longe stabunt propter timorem tormentorum eius flentes ac lugentes
REV|18|16|et dicentes vae vae civitas illa magna quae amicta erat byssino et purpura et cocco et deaurata est auro et lapide pretioso et margaritis
REV|18|17|quoniam una hora destitutae sunt tantae divitiae et omnis gubernator et omnis qui in locum navigat et nautae et qui maria operantur longe steterunt
REV|18|18|et clamaverunt videntes locum incendii eius dicentes quae similis civitati huic magnae
REV|18|19|et miserunt pulverem super capita sua et clamaverunt flentes et lugentes dicentes vae vae civitas magna in qua divites facti sunt omnes qui habent naves in mari de pretiis eius quoniam una hora desolata est
REV|18|20|exulta super eam caelum et sancti et apostoli et prophetae quoniam iudicavit Deus iudicium vestrum de illa
REV|18|21|et sustulit unus angelus fortis lapidem quasi molarem magnum et misit in mare dicens hoc impetu mittetur Babylon magna illa civitas et ultra iam non invenietur
REV|18|22|et vox citharoedorum et musicorum et tibia canentium et tuba non audietur in te amplius et omnis artifex omnis artis non invenietur in te amplius et vox molae non audietur in te amplius
REV|18|23|et lux lucernae non lucebit tibi amplius et vox sponsi et sponsae non audietur adhuc in te quia mercatores tui erant principes terrae quia in veneficiis tuis erraverunt omnes gentes
REV|18|24|et in ea sanguis prophetarum et sanctorum inventus est et omnium qui interfecti sunt in terra
REV|19|1|post haec audivi quasi vocem magnam turbarum multarum in caelo dicentium alleluia salus et gloria et virtus Deo nostro est
REV|19|2|quia vera et iusta iudicia sunt eius quia iudicavit de meretrice magna quae corrupit terram in prostitutione sua et vindicavit sanguinem servorum suorum de manibus eius
REV|19|3|et iterum dixerunt alleluia et fumus eius ascendit in saecula saeculorum
REV|19|4|et ceciderunt seniores viginti quattuor et quattuor animalia et adoraverunt Deum sedentem super thronum dicentes amen alleluia
REV|19|5|et vox de throno exivit dicens laudem dicite Deo nostro omnes servi eius et qui timetis eum pusilli et magni
REV|19|6|et audivi quasi vocem turbae magnae et sicut vocem aquarum multarum et sicut vocem tonitruum magnorum dicentium alleluia quoniam regnavit Dominus Deus noster omnipotens
REV|19|7|gaudeamus et exultemus et demus gloriam ei quia venerunt nuptiae agni et uxor eius praeparavit se
REV|19|8|et datum est illi ut cooperiat se byssinum splendens candidum byssinum enim iustificationes sunt sanctorum
REV|19|9|et dicit mihi scribe beati qui ad cenam nuptiarum agni vocati sunt et dicit mihi haec verba vera Dei sunt
REV|19|10|et cecidi ante pedes eius ut adorarem eum et dicit mihi vide ne feceris conservus tuus sum et fratrum tuorum habentium testimonium Iesu Deum adora testimonium enim Iesu est spiritus prophetiae
REV|19|11|et vidi caelum apertum et ecce equus albus et qui sedebat super eum vocabatur Fidelis et Verax vocatur et iustitia iudicat et pugnat
REV|19|12|oculi autem eius sicut flamma ignis et in capite eius diademata multa habens nomen scriptum quod nemo novit nisi ipse
REV|19|13|et vestitus erat vestem aspersam sanguine et vocatur nomen eius Verbum Dei
REV|19|14|et exercitus qui sunt in caelo sequebantur eum in equis albis vestiti byssinum album mundum
REV|19|15|et de ore ipsius procedit gladius acutus ut in ipso percutiat gentes et ipse reget eos in virga ferrea et ipse calcat torcular vini furoris irae Dei omnipotentis
REV|19|16|et habet in vestimento et in femore suo scriptum rex regum et Dominus dominantium
REV|19|17|et vidi unum angelum stantem in sole et clamavit voce magna dicens omnibus avibus quae volabant per medium caeli venite congregamini ad cenam magnam Dei
REV|19|18|ut manducetis carnes regum et carnes tribunorum et carnes fortium et carnes equorum et sedentium in ipsis et carnes omnium liberorum ac servorum et pusillorum ac magnorum
REV|19|19|et vidi bestiam et reges terrae et exercitus eorum congregatos ad faciendum proelium cum illo qui sedebat in equo et cum exercitu eius
REV|19|20|et adprehensa est bestia et cum illo pseudopropheta qui fecit signa coram ipso quibus seduxit eos qui acceperunt caracterem bestiae qui et adorant imaginem eius vivi missi sunt hii duo in stagnum ignis ardentis sulphure
REV|19|21|et ceteri occisi sunt in gladio sedentis super equum qui procedit de ore ipsius et omnes aves saturatae sunt carnibus eorum
REV|20|1|et vidi angelum descendentem de caelo habentem clavem abyssi et catenam magnam in manu sua
REV|20|2|et adprehendit draconem serpentem antiquum qui est diabolus et Satanas et ligavit eum per annos mille
REV|20|3|et misit eum in abyssum et clusit et signavit super illum ut non seducat amplius gentes donec consummentur mille anni post haec oportet illum solvi modico tempore
REV|20|4|et vidi sedes et sederunt super eas et iudicium datum est illis et animas decollatorum propter testimonium Iesu et propter verbum Dei et qui non adoraverunt bestiam neque imaginem eius nec acceperunt caracterem in frontibus aut in manibus suis et vixerunt et regnaverunt cum Christo mille annis
REV|20|5|ceteri mortuorum non vixerunt donec consummentur mille anni haec est resurrectio prima
REV|20|6|beatus et sanctus qui habet partem in resurrectione prima in his secunda mors non habet potestatem sed erunt sacerdotes Dei et Christi et regnabunt cum illo mille annis
REV|20|7|et cum consummati fuerint mille anni solvetur Satanas de carcere suo et exibit et seducet gentes quae sunt super quattuor angulos terrae Gog et Magog et congregabit eos in proelium quorum numerus est sicut harena maris
REV|20|8|et ascenderunt super latitudinem terrae et circumierunt castra sanctorum et civitatem dilectam
REV|20|9|et descendit ignis a Deo de caelo et devoravit eos et diabolus qui seducebat eos missus est in stagnum ignis et sulphuris ubi et bestia
REV|20|10|et pseudoprophetes et cruciabuntur die ac nocte in saecula saeculorum
REV|20|11|et vidi thronum magnum candidum et sedentem super eum a cuius aspectu fugit terra et caelum et locus non est inventus ab eis
REV|20|12|et vidi mortuos magnos et pusillos stantes in conspectu throni et libri aperti sunt et alius liber apertus est qui est vitae et iudicati sunt mortui ex his quae scripta erant in libris secundum opera ipsorum
REV|20|13|et dedit mare mortuos qui in eo erant et mors et inferus dederunt mortuos qui in ipsis erant et iudicatum est de singulis secundum opera ipsorum
REV|20|14|et inferus et mors missi sunt in stagnum ignis haec mors secunda est stagnum ignis
REV|20|15|et qui non est inventus in libro vitae scriptus missus est in stagnum ignis
REV|21|1|et vidi caelum novum et terram novam primum enim caelum et prima terra abiit et mare iam non est
REV|21|2|et civitatem sanctam Hierusalem novam vidi descendentem de caelo a Deo paratam sicut sponsam ornatam viro suo
REV|21|3|et audivi vocem magnam de throno dicentem ecce tabernaculum Dei cum hominibus et habitabit cum eis et ipsi populus eius erunt et ipse Deus cum eis erit eorum Deus
REV|21|4|et absterget Deus omnem lacrimam ab oculis eorum et mors ultra non erit neque luctus neque clamor neque dolor erit ultra quae prima abierunt
REV|21|5|et dixit qui sedebat in throno ecce nova facio omnia et dicit scribe quia haec verba fidelissima sunt et vera
REV|21|6|et dixit mihi factum est ego sum Alpha et Omega initium et finis ego sitienti dabo de fonte aquae vivae gratis
REV|21|7|qui vicerit possidebit haec et ero illi Deus et ille erit mihi filius
REV|21|8|timidis autem et incredulis et execratis et homicidis et fornicatoribus et veneficis et idolatris et omnibus mendacibus pars illorum erit in stagno ardenti igne et sulphure quod est mors secunda
REV|21|9|et venit unus de septem angelis habentibus fialas plenas septem plagis novissimis et locutus est mecum dicens veni ostendam tibi sponsam uxorem agni
REV|21|10|et sustulit me in spiritu in montem magnum et altum et ostendit mihi civitatem sanctam Hierusalem descendentem de caelo a Deo
REV|21|11|habentem claritatem Dei lumen eius simile lapidi pretioso tamquam lapidi iaspidis sicut cristallum
REV|21|12|et habebat murum magnum et altum habens portas duodecim et in portis angelos duodecim et nomina inscripta quae sunt nomina duodecim tribuum filiorum Israhel
REV|21|13|ab oriente portae tres et ab aquilone portae tres et ab austro portae tres et ab occasu portae tres
REV|21|14|et murus civitatis habens fundamenta duodecim et in ipsis duodecim nomina duodecim apostolorum agni
REV|21|15|et qui loquebatur mecum habebat mensuram harundinem auream ut metiretur civitatem et portas eius et murum
REV|21|16|et civitas in quadro posita est et longitudo eius tanta est quanta et latitudo et mensus est civitatem de harundine per stadia duodecim milia longitudo et latitudo et altitudo eius aequalia sunt
REV|21|17|et mensus est murus eius centum quadraginta quattuor cubitorum mensura hominis quae est angeli
REV|21|18|et erat structura muri eius ex lapide iaspide ipsa vero civitas auro mundo simile vitro mundo
REV|21|19|fundamenta muri civitatis omni lapide pretioso ornata fundamentum primum iaspis secundus sapphyrus tertius carcedonius quartus zmaragdus
REV|21|20|quintus sardonix sextus sardinus septimus chrysolitus octavus berillus nonus topazius decimus chrysoprassus undecimus hyacinthus duodecimus amethistus
REV|21|21|et duodecim portae duodecim margaritae sunt per singulas et singulae portae erant ex singulis margaritis et platea civitatis aurum mundum tamquam vitrum perlucidum
REV|21|22|et templum non vidi in ea Dominus enim Deus omnipotens templum illius est et agnus
REV|21|23|et civitas non eget sole neque luna ut luceant in ea nam claritas Dei inluminavit eam et lucerna eius est agnus
REV|21|24|et ambulabunt gentes per lumen eius et reges terrae adferent gloriam suam et honorem in illam
REV|21|25|et portae eius non cludentur per diem nox enim non erit illic
REV|21|26|et adferent gloriam et honorem gentium in illam
REV|21|27|nec intrabit in ea aliquid coinquinatum et faciens abominationem et mendacium nisi qui scripti sunt in libro vitae agni
REV|22|1|et ostendit mihi fluvium aquae vitae splendidum tamquam cristallum procedentem de sede Dei et agni
REV|22|2|in medio plateae eius et ex utraque parte fluminis lignum vitae adferens fructus duodecim per menses singula reddentia fructum suum et folia ligni ad sanitatem gentium
REV|22|3|et omne maledictum non erit amplius et sedes Dei et agni in illa erunt et servi eius servient illi
REV|22|4|et videbunt faciem eius et nomen eius in frontibus eorum
REV|22|5|et nox ultra non erit et non egebunt lumine lucernae neque lumine solis quoniam Dominus Deus inluminat illos et regnabunt in saecula saeculorum
REV|22|6|et dixit mihi haec verba fidelissima et vera sunt et Dominus Deus spirituum prophetarum misit angelum suum ostendere servis suis quae oportet fieri cito
REV|22|7|et ecce venio velociter beatus qui custodit verba prophetiae libri huius
REV|22|8|et ego Iohannes qui audivi et vidi haec et postquam audissem et vidissem cecidi ut adorarem ante pedes angeli qui mihi haec ostendebat
REV|22|9|et dicit mihi vide ne feceris conservus tuus sum et fratrum tuorum prophetarum et eorum qui servant verba libri huius Deum adora
REV|22|10|et dicit mihi ne signaveris verba prophetiae libri huius tempus enim prope est
REV|22|11|qui nocet noceat adhuc et qui in sordibus est sordescat adhuc et iustus iustitiam faciat adhuc et sanctus sanctificetur adhuc
REV|22|12|ecce venio cito et merces mea mecum est reddere unicuique secundum opera sua
REV|22|13|ego Alpha et Omega primus et novissimus principium et finis
REV|22|14|beati qui lavant stolas suas ut sit potestas eorum in ligno vitae et portis intrent in civitatem
REV|22|15|foris canes et venefici et inpudici et homicidae et idolis servientes et omnis qui amat et facit mendacium
REV|22|16|ego Iesus misi angelum meum testificari vobis haec in ecclesiis ego sum radix et genus David stella splendida et matutina
REV|22|17|et Spiritus et sponsa dicunt veni et qui audit dicat veni et qui sitit veniat qui vult accipiat aquam vitae gratis
REV|22|18|contestor ego omni audienti verba prophetiae libri huius si quis adposuerit ad haec adponet Deus super illum plagas scriptas in libro isto
REV|22|19|et si quis deminuerit de verbis libri prophetiae huius auferet Deus partem eius de ligno vitae et de civitate sancta et de his quae scripta sunt in libro isto
REV|22|20|dicit qui testimonium perhibet istorum etiam venio cito amen veni Domine Iesu
REV|22|21|gratia Domini nostri Iesu Christi cum omnibus
