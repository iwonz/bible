LEV|1|1|Vocavit autem Moysen et locu tus est ei Dominus de tabernacu lo conventus dicens:
LEV|1|2|" Loquere filiis Israel et dices ad eos: Homo, qui obtulerit ex vobis hostiam Domino de animalibus domesticis, de bobus et pecoribus offerens victimas,
LEV|1|3|si holocaustum fuerit eius oblatio de armento, masculum immaculatum offeret ad ostium tabernaculi conventus ad placandum sibi Dominum;
LEV|1|4|ponetque manum super caput hostiae, et acceptabilis erit atque in expiationem eius proficiens.
LEV|1|5|Immolabitque vitulum coram Domino, et offerent filii Aaron sacerdotes sanguinem eius aspergentes per altaris circuitum, quod est ante ostium tabernaculi conventus.
LEV|1|6|Detracta pelle, hostiam offerens in frusta concidet;
LEV|1|7|et filii Aaron sacerdotis ponent in altari ignem, strueque lignorum super ignem composita,
LEV|1|8|membra, quae caesa sunt, desuper ordinabunt, caput videlicet et adipem.
LEV|1|9|Intestina autem et crura offerens lavabit aqua adolebitque ea sacerdos super altare in holocaustum, incensum suavissimi odoris Domino.
LEV|1|10|Quod si de pecoribus eius oblatio est, de ovibus sive de capris holocaustum, masculum absque macula offeret;
LEV|1|11|immolabitque ad latus altaris, quod respicit ad aquilonem, coram Domino. Sanguinem vero illius aspergent contra altare filii Aaron sacerdotes per circuitum;
LEV|1|12|dividetque offerens membra, caput et adipem, et sacerdos imponet ea super ligna, quibus subest ignis in altari.
LEV|1|13|Intestina vero et crura lavabit offerens aqua, et oblata omnia adolebit sacerdos super altare: holocaustum est et incensum odoris suavissimi Domino.
LEV|1|14|Sin autem de avibus holocausti oblatio fuerit Domino, offeret de turturibus aut pullis columbae oblationem suam.
LEV|1|15|Et sacerdos afferet eam ad altare; retortum ad collum caput adolebit in altari, sanguisque eius exprimetur contra parietem altaris.
LEV|1|16|Vesiculam vero gutturis et plumas proiciet offerens prope altare ad orientalem plagam in loco, in quo cineres effundi solent;
LEV|1|17|confringetque eam inter alas, quas non secabit, et adolebit eam sacerdos super altare, lignis super ignem positis: holocaustum est et incensum suavissimi odoris Domino.
LEV|2|1|Anima cum obtulerit oblationem sacrificii farinae Domino, simila erit eius oblatio, fundetque super eam oleum et ponet tus
LEV|2|2|ac deferet ad filios Aaron sacerdotes, tolletque ex eo pugillum plenum similae et olei ac totum tus, et sacerdos adolebit memoriale super altare, incensum odoris suavissimi Domino.
LEV|2|3|Quod autem reliquum fuerit de sacrificio, erit Aaron et filiorum eius: sanctum sanctorum de incensis Domini.
LEV|2|4|Cum autem obtuleris sacrificium similae coctum in clibano: de simila erunt panes, scilicet absque fermento conspersi oleo et lagana azyma oleo lita;
LEV|2|5|si oblatio tua fuerit de sartagine, simila erit, conspersa oleo et absque fermento;
LEV|2|6|divides eam minutatim et fundes super eam oleum: oblatio similae est.
LEV|2|7|Sin autem de frixorio fuerit sacrificium, aeque simila oleo conspergetur.
LEV|2|8|Et deferes oblationem ex his Domino factam tradens manibus sacerdotis,
LEV|2|9|qui afferet eam ad altare, tollet memoriale de sacrificio et adolebit super altare: incensum odoris suavissimi Domino.
LEV|2|10|Quidquid autem reliquum est, erit Aaron et filiorum eius: sanctum sanctorum de incensis Domini.
LEV|2|11|Omnis oblatio similae, quam offeretis Domino, absque fermento fiet, quia nihil fermenti ac mellis adolebitis incensum Domino.
LEV|2|12|Primitias tantum eorum offeretis tamquam munera Domino; super altare vero non ponentur in odorem suavitatis.
LEV|2|13|Quidquid obtuleris sacrificii, similae sale condies nec auferes sal foederis Dei tui de sacrificio tuo: in omni oblatione tua offeres sal.
LEV|2|14|Sin autem obtuleris munus primarum frugum tuarum Domino, spicas tostas igni et grana fracta farris recentis offeres in sacrificium primarum frugum tuarum
LEV|2|15|fundens supra oleum et tus imponens: similae oblatio est.
LEV|2|16|De qua adolebit sacerdos tamquam memoriale partem farris fracti et olei ac totum tus.
LEV|3|1|Quod si hostia pacificorum fue rit eius oblatio et de bobus vo luerit offerre marem sive feminam, immaculata offeret coram Domino.
LEV|3|2|Ponetque manum super caput victimae suae, quam immolabit ad ostium tabernaculi conventus, fundentque filii Aaron sacerdotes sanguinem per circuitum altaris
LEV|3|3|et offerent de hostia pacificorum tamquam incensum Domino adipem, qui operit vitalia, et quidquid pinguedinis eis adhaeret,
LEV|3|4|duos renes cum adipe, quo teguntur iuxta ilia, et reticulum iecoris, quem iuxta renes, auferet.
LEV|3|5|Adolebuntque ea filii Aaron in altari super holocausto, quod est super lignis et igne: incensum suavissimi odoris Domino.
LEV|3|6|Si vero de pecoribus fuerit Domino eius oblatio, pacificorum scilicet hostia, sive masculum sive feminam obtulerit, immaculata erunt.
LEV|3|7|Si agnum obtulerit coram Domino,
LEV|3|8|ponet manum super caput victimae suae, quam immolabit coram tabernaculo conventus; fundentque filii Aaron sanguinem eius per altaris circuitum;
LEV|3|9|et offeret de pacificorum hostia incensum Domino adipem et caudam totam, quam iuxta tergum, auferet, et pinguedinem, quae operit ventrem, atque universum adipem, qui vitalibus adhaeret,
LEV|3|10|et utrumque renunculum cum adipe, qui est iuxta ilia, reticulumque iecoris, quem iuxta renunculos, auferet.
LEV|3|11|Et adolebit ea sacerdos super altare: panis et incensum Domino.
LEV|3|12|Si capra fuerit eius oblatio, offeret eam coram Domino,
LEV|3|13|ponet manum suam super caput eius immolabitque eam coram tabernaculo conventus. Et fundent filii Aaron sanguinem eius per altaris circuitum,
LEV|3|14|tolletque ex ea oblationem suam, incensum Domino, adipem scilicet, qui operit ventrem, et universum, qui vitalibus adhaeret,
LEV|3|15|duos renunculos cum adipe, qui est super eos iuxta ilia, et reticulum iecoris, quem iuxta renunculos, auferet;
LEV|3|16|adolebitque ea sacerdos super altare: panis et incensum suavissimi odoris omnis adeps Domino.
LEV|3|17|Iure perpetuo in generationibus et cunctis habitaculis vestris, nec adipem nec sanguinem omnino comedetis ".
LEV|4|1|Locutusque est Dominus ad Moysen dicens:
LEV|4|2|" Loquere filiis Israel: Anima cum peccaverit per ignorantiam et de universis mandatis Domini, quae praecepit ut non fierent, quippiam fecerit,
LEV|4|3|si sacerdos, qui est unctus, peccaverit, delinquere faciens populum, offeret pro peccato suo vitulum immaculatum Domino sacrificium pro peccato;
LEV|4|4|et adducet illum ad ostium tabernaculi conventus coram Domino ponetque manum super caput eius et immolabit eum coram Domino.
LEV|4|5|Hauriet quoque sacerdos unctus de sanguine vituli inferens illum in tabernaculum conventus;
LEV|4|6|cumque intinxerit digitum in sanguinem, asperget eo septies coram Domino contra velum sanctuarii;
LEV|4|7|ponetque de eodem sanguine super cornua altaris thymiamatis gratissimi coram Domino, quod est in tabernaculo conventus; omnem autem reliquum sanguinem fundet in basim altaris holocausti in introitu tabernaculi.
LEV|4|8|Et omnem adipem vituli pro peccato auferet tam eum, qui operit vitalia, quam omnem, qui vitalibus adhaeret,
LEV|4|9|duos renunculos et adipem, qui est super eos iuxta ilia, et reticulum iecoris, quem iuxta renunculos, auferet,
LEV|4|10|sicut aufertur de vitulo hostiae pacificorum; et adolebit ea sacerdos super altare holocausti.
LEV|4|11|Pellem vero et omnes carnes cum capite et pedibus et intestinis et fimo,
LEV|4|12|totum vitulum efferet extra castra in locum mundum, ubi cineres effundi solent; incendetque eum super lignorum struem igne: in loco effusorum cinerum cremabitur.
LEV|4|13|Quod si omnis coetus Israel ignoraverit, et res abscondita fuerit ab oculis congregationis, feceritque quod contra mandatum Domini est et deliquerit,
LEV|4|14|et postea intellexerit peccatum suum, offeret congregatio vitulum pro peccato adducetque eum ad ostium tabernaculi conventus.
LEV|4|15|Et ponent seniores coetus populi manus super caput eius coram Domino, immolatoque vitulo in conspectu Domini,
LEV|4|16|inferet sacerdos, qui unctus est, de sanguine eius in tabernaculum conventus,
LEV|4|17|tincto digito aspergens septies contra velum;
LEV|4|18|ponetque de eodem sanguine in cornibus altaris, quod est coram Domino in tabernaculo conventus. Reliquum autem sanguinem fundet iuxta basim altaris holocaustorum, quod est in ostio tabernaculi conventus;
LEV|4|19|omnemque eius adipem tollet et adolebit super altare.
LEV|4|20|Sic faciens et de hoc vitulo quomodo fecit de vitulo pro peccato; sic faciet ei. Expiante eos sacerdote, propitius erit Dominus.
LEV|4|21|Ipsum autem vitulum efferet extra castra atque comburet sicut et priorem vitulum: sacrificium pro peccato est congregationis.
LEV|4|22|Si peccaverit princeps et fecerit unum ex omnibus per ignorantiam, quod Domini Dei sui lege prohibetur, deliqueritque,
LEV|4|23|aut indicatum ei fuerit peccatum suum, offeret hostiam Domino hircum de capris immaculatum
LEV|4|24|ponetque manum suam super caput eius et immolabit eum in loco, ubi solet mactari holocaustum coram Domino: sacrificium pro peccato est.
LEV|4|25|Et tinguat sacerdos digitum in sanguine hostiae pro peccato ponetque super cornua altaris holocausti et reliquum fundet ad basim eius.
LEV|4|26|Adipem vero adolebit supra, sicut in victimis pacificorum fieri solet; expiabitque eum a peccato eius, ac dimittetur ei.
LEV|4|27|Quod si peccaverit anima per ignorantiam de populo terrae, ut faciat quidquam ex his, quae Domini lege prohibentur, atque delinquat,
LEV|4|28|aut indicatum ei fuerit peccatum suum, offeret capram immaculatam;
LEV|4|29|ponetque manum super caput hostiae pro peccato et immolabit eam in loco holocausti.
LEV|4|30|Tolletque sacerdos de sanguine in digito suo et ponet super cornua altaris holocausti et reliquum fundet ad basim eius.
LEV|4|31|Omnem autem auferens adipem, sicut auferri solet de victimis pacificorum, adolebit super altare in odorem suavitatis Domino, expiabitque eum, et propitius erit Dominus.
LEV|4|32|Sin autem de ovibus obtulerit victimam pro peccato, adducet agnam immaculatam;
LEV|4|33|ponet manum super caput eius et immolabit eam in loco, ubi solent holocaustorum caedi hostiae.
LEV|4|34|Sumetque sacerdos de sanguine eius digito suo et ponens super cornua altaris holocausti reliquum fundet ad basim eius.
LEV|4|35|Omnem quoque auferens adipem, sicut auferri solet adeps agni, qui immolatur pro pacificis, cremabit in altari super incensis Domini; expiabitque eum et peccatum eius, et dimittetur illi.
LEV|5|1|Si peccaverit anima et audiverit vocem iurantis testisque fuerit, quod aut ipse vidit aut comperit, si non indicaverit, iniquitatem portabit;
LEV|5|2|vel si anima tetigerit aliquid immundum, sive cadaver bestiae sit aut iumenti vel reptilis, et absconditum fuerit ab eo, ipse immundus et reus erit;
LEV|5|3|aut si tetigerit quidquam de immunditia hominis iuxta omnem impuritatem, qua pollui solet, absconditumque fuerit ab eo, sed ipse cognoverit postea, subiacebit delicto;
LEV|5|4|aut si anima temere iuraverit et protulerit labiis suis, ut vel male quid faceret vel bene iuxta omnia, quae homines temere iurant, absconditumque fuerit ab eo, sed ipse postea intellexerit, delicto subiacebit;
LEV|5|5|si ergo reus factus fuerit uno ex istis, confiteatur peccatum suum
LEV|5|6|et offerat Domino sacrificium delicti pro peccato suo agnam de gregibus sive capram ut sacrificium pro peccato; expiabitque eum sacerdos a peccato eius.
LEV|5|7|Sin autem non potuerit offerre pecus, offerat ut sacrificium pro delicto duos turtures vel duos pullos columbarum Domino: unum in sacrificium pro peccato et alterum in holocaustum;
LEV|5|8|dabitque eos sacerdoti, qui primum offerens ut sacrificium pro peccato retorquebit caput eius ad pennulas, ita ut collo haereat et non penitus abrumpatur;
LEV|5|9|et asperget de sanguine eius parietem altaris; quidquid autem reliquum fuerit, faciet destillare ad fundamentum eius: sacrificium pro peccato est.
LEV|5|10|Alterum vero adolebit holocaustum, ut fieri solet; expiabitque eum sacerdos a peccato eius, et dimittetur ei.
LEV|5|11|Quod si non quiverit manus eius offerre duos turtures aut duos pullos columbarum, offeret pro peccato suo similae partem ephi decimam in sacrificium pro peccato; non mittet in eam oleum, nec turis aliquid imponet, quia sacrificium pro peccato est.
LEV|5|12|Tradetque eam sacerdoti, qui, plenum ex toto pugillum in memoriale hauriens, cremabit in altari super incensis Domini: sacrificium pro peccato est.
LEV|5|13|Et expiabit eum sacerdos et peccatum eius in uno ex his casibus, et propitius erit Dominus. Reliquam vero partem sacerdos habebit sicut in oblatione similae ".
LEV|5|14|Locutus est Dominus ad Moysen dicens:
LEV|5|15|" Anima, si praevaricans per errorem in his, quae Domino sunt sanctificata, peccaverit, offeret sacrificium pro delicto arietem immaculatum de gregibus iuxta aestimationem argenti siclorum pondere sanctuarii in paenitentiam;
LEV|5|16|ipsumque, quod intulit damni, restituet et quintam partem ponet supra tradens sacerdoti, qui expiabit eum offerens arietem, et dimittetur ei.
LEV|5|17|Anima, si peccaverit per ignorantiam feceritque unum ex his, quae Domini lege prohibentur, et peccati rea portaverit iniquitatem suam,
LEV|5|18|offeret arietem immaculatum de gregibus iuxta aestimationem sacerdoti, qui expiabit eum ab eo, quod nesciens fecerit, et dimittetur ei:
LEV|5|19|sacrificium pro delicto est, delinquens deliquit in Dominum ".
LEV|5|20|Locutus est Dominus ad Moysen dicens:
LEV|5|21|" Anima, quae peccaverit et, contempto Domino, negaverit proximo suo depositum, quod fidei eius creditum fuerat, vel vi aliquid extorserit aut calumniam fecerit,
LEV|5|22|sive rem perditam invenerit et infitians insuper peierarit in uno ex omnibus, in quibus peccare solent homines,
LEV|5|23|si quis sic peccaverit et deliquerit, reddet omnia, quae per rapinam vel calumniam abstulerit vel deposita retinuerit vel perdita invenerit
LEV|5|24|vel de quibus peierarit, et restituet integra et quintam insuper addet partem domino, cui damnum intulerat, in die sacrificii pro delicto.
LEV|5|25|Sacrificium pro delicto offeret Domino: arietem immaculatum de grege iuxta aestimationem;
LEV|5|26|qui expiabit eum coram Domino, et dimittetur illi pro singulis, quae faciendo peccaverit ".
LEV|6|1|Locutus est Dominus ad Moysen dicens:
LEV|6|2|" Praecipe Aaron et filiis eius: Haec est lex holocausti: cremabitur in foco altaris tota nocte usque mane; ignis altaris in eo ardebit.
LEV|6|3|Vestietur sacerdos tunica et feminalibus lineis super verecunda sua; tolletque cineres, quos vorans ignis exussit, et ponet iuxta altare.
LEV|6|4|Porro spoliabitur prioribus vestimentis; indutusque aliis efferet cineres extra castra in locum mundum.
LEV|6|5|Ignis autem in altari semper ardebit, non exstinguetur, quem nutriet sacerdos subiciens ligna mane per singulos dies et, imposito holocausto, desuper adolebit adipes pacificorum.
LEV|6|6|Ignis est iste perpetuus, qui numquam deficiet in altari.
LEV|6|7|Haec est lex sacrificii similae, quod offerent filii Aaron coram Domino et coram altare:
LEV|6|8|tollet sacerdos ex eo pugillum similae, quae conspersa est oleo, et totum tus, quod super similam positum est; adolebitque illud in altari in odorem suavissimum, memoriale Domino.
LEV|6|9|Reliquam autem partem similae comedet Aaron cum filiis suis, et panis absque fermento comedetur in loco sancto; in atrio tabernaculi conventus comedent illam.
LEV|6|10|Ideo autem non coquetur fermentata, quia ut partem eorum dedi illam ex incensis meis: sanctum sanctorum est, sicut sacrificium pro peccato atque pro delicto;
LEV|6|11|mares tantum stirpis Aaron comedent illud. Legitimum sempiternum est in generationibus vestris de incensis Domini; omnis, qui tetigerit illa, sanctificabitur ".
LEV|6|12|Et locutus est Dominus ad Moysen dicens:
LEV|6|13|" Haec est oblatio Aaron et filiorum eius, quam offerre debent Domino in die unctionis ipsius: decimam partem ephi offerent similae in sacrificio sempiterno medium eius mane et medium vespere;
LEV|6|14|quae in sartagine oleo conspersa frigetur. Afferes eam calidam et offeres divisam minutatim, sacrificium in odorem suavissimum Domino.
LEV|6|15|Sacerdos unctus, qui patri iure successerit, faciet illud. Legitimum sempiternum: Domino tota cremabitur;
LEV|6|16|omne enim sacrificium similae sacerdotum igne consumetur, nec quisquam comedet ex eo ".
LEV|6|17|Locutus est Dominus ad Moysen dicens:
LEV|6|18|" Loquere Aaron et filiis eius: Ista est lex sacrificii pro peccato: in loco, ubi mactatur holocaustum, mactabitur coram Domino: sanctum sanctorum est.
LEV|6|19|Sacerdos, qui offert, comedet illud in loco sancto, in atrio tabernaculi conventus.
LEV|6|20|Quidquid tetigerit carnes eius, sanctificabitur: si de sanguine illius vestis fuerit aspersa, lavabitur in loco sancto;
LEV|6|21|vas autem fictile, in quo coctum est, confringetur; quod si vas aeneum fuerit, defricabitur et lavabitur aqua.
LEV|6|22|Omnis masculus de genere sacerdotali vescetur carnibus eius, quia sanctum sanctorum est.
LEV|6|23|Omne autem sacrificium pro peccato, de cuius sanguine infertur in tabernaculum conventus ad expiandum in sanctuario, non comedetur, sed comburetur igni.
LEV|7|1|Haec quoque est lex sacrificii pro delicto: sanctum sanctorum est,
LEV|7|2|idcirco, ubi immolatur holocaustum, mactabitur et victima pro delicto; sanguis eius per gyrum fundetur altaris.
LEV|7|3|Omnemque adipem offeret ex ea, caudam scilicet et adipem, qui operit vitalia,
LEV|7|4|duos renunculos et pinguedinem, quae super eos iuxta ilia est, reticulumque iecoris, quem iuxta renunculos, auferet;
LEV|7|5|et adolebit ea sacerdos super altare ut incensum Domino: sacrificium pro delicto est.
LEV|7|6|Omnis masculus de sacerdotali genere in loco sancto vescetur his carnibus, quia sanctum sanctorum est.
LEV|7|7|Sicut sacrificium pro peccato, ita et sacrificium pro delicto, utriusque hostiae lex una est; ad sacerdotem, qui eam obtulerit, pertinebit.
LEV|7|8|Sacerdos, qui offert holocaustum cuiusdam viri, habebit pellem victimae,
LEV|7|9|et omne sacrificium similae, quod coquitur in clibano, et, quidquid in frixorio vel in sartagine praeparatur, eius erit sacerdotis, a quo offertur;
LEV|7|10|et omne sacrificium similae sive oleo conspersum sive aridum fuerit, cunctis filiis Aaron aequa mensura per singulos dividetur.
LEV|7|11|Haec est lex hostiae pacificorum quae offertur Domino;
LEV|7|12|si pro gratiarum actione fuerit oblatio, offerent panes absque fermento conspersos oleo et lagana azyma uncta oleo coctamque similam ut collyridas olei admixtione conspersas,
LEV|7|13|panes quoque fermentatos cum hostia pacificorum pro gratiarum actione,
LEV|7|14|ex quibus unus offeretur munus Domino et erit sacerdotis, qui fundet hostiae sanguinem.
LEV|7|15|Cuius carnes eadem comedentur die, nec remanebit ex eis quidquam usque mane.
LEV|7|16|Si voto vel sponte quisquam obtulerit hostiam, eadem similiter edetur die; sed et si quid in crastinum remanserit, vesci licitum est;
LEV|7|17|quidquid autem tertius invenerit dies, ignis absumet.
LEV|7|18|Si quis de carnibus victimae pacificorum die tertio comederit, irrita fiet oblatio nec proderit offerenti; quin potius, quaecumque anima tali se edulio contaminarit, praevaricationis rea erit.
LEV|7|19|Caro, quae aliquid tetigerit immundum, non comedetur, sed comburetur igni; ceterum carne, qui fuerit mundus, vescetur.
LEV|7|20|Anima polluta, quae ederit de carnibus hostiae pacificorum, quae oblata est Domino, peribit de populis suis;
LEV|7|21|et, quae tetigerit immunditiam hominis vel iumenti, sive omnis rei abominabilis, quae polluere potest, et comederit de huiuscemodi carnibus, interibit de populis suis ".
LEV|7|22|Locutusque est Dominus ad Moysen dicens:
LEV|7|23|" Loquere filiis Israel: Adipem bovis et ovis et caprae non comedetis.
LEV|7|24|Adipem cadaveris morticini et eius animalis, quod a bestia laceratum est, habebitis in usus varios, sed non comedetis.
LEV|7|25|Si quis adipem, qui offertur in incensum Domini, comederit, peribit de populo suo.
LEV|7|26|Sanguinem quoque omnis animalis non sumetis in cibo, tam de avibus quam de pecoribus;
LEV|7|27|omnis anima, quae ederit sanguinem, peribit de populis suis ".
LEV|7|28|Locutus est Dominus ad Moysen dicens:
LEV|7|29|" Loquere filiis Israel: Qui offert victimam pacificorum Domino, afferat oblationem suam Domino de victima pacificorum.
LEV|7|30|Tenebit manibus incensa Domini, adipem scilicet et pectusculum afferet; pectusculum, ut elevetur coram Domino.
LEV|7|31|Et sacerdos adolebit adipem super altare; pectusculum autem erit Aaron et filiorum eius.
LEV|7|32|Armus quoque dexter de pacificorum hostiis cedet in munus sacerdotis.
LEV|7|33|Qui de filiis Aaron obtulerit sanguinem et adipem victimae pacificorum, ipse habebit armum dextrum in portione sua;
LEV|7|34|pectusculum enim elationis et armum donationis tuli a filiis Israel de hostiis eorum pacificis et dedi Aaron sacerdoti ac filiis eius, lege perpetua, ab omni populo Israel ".
LEV|7|35|Haec est portio Aaron et filiorum eius de incensis Domini die, qua applicavit eos, ut sacerdotio fungerentur;
LEV|7|36|et quae praecepit dari eis Dominus a filiis Israel die, qua unxit eos, religione perpetua in generationibus eorum.
LEV|7|37|Ista est lex holocausti et oblationis similae et sacrificii pro peccato atque delicto et pro consecratione et pacificorum victimis,
LEV|7|38|quam constituit Dominus Moysi in monte Sinai, quando mandavit filiis Israel, ut offerrent oblationes suas Domino in deserto Sinai.
LEV|8|1|Locutusque est Dominus ad Moysen dicens:
LEV|8|2|" Tolle Aaron cum filiis suis, vestes eorum et unctionis oleum, vitulum pro peccato, duos arietes, canistrum cum azymis;
LEV|8|3|et congregabis omnem coetum ad ostium tabernaculi conventus ".
LEV|8|4|Fecit Moyses, ut Dominus imperarat; congregatoque omni coetu ante fores tabernaculi conventus,
LEV|8|5|ait: " Iste est sermo, quem iussit Dominus fieri ".
LEV|8|6|Statimque applicavit Aaron et filios eius. Cumque lavisset eos aqua,
LEV|8|7|vestivit pontificem subucula linea accingens eum balteo et induens tunica hyacinthina et desuper ephod imposuit,
LEV|8|8|quod astrinxit cingulo ephod firmiter; et imposuit ei pectorale, in quo dedit Urim et Tummim.
LEV|8|9|Cidari quoque texit caput et super eam contra frontem posuit laminam auream, diadema sanctum, sicut praeceperat Dominus Moysi.
LEV|8|10|Tulit et unctionis oleum, quo levit habitaculum cum omni supellectili sua et sanctificavit ea.
LEV|8|11|Cumque de eo aspersisset altare septem vicibus, unxit illud et omnia vasa eius labrumque cum basi sua sanctificavit oleo.
LEV|8|12|Quod fundens super caput Aaron, unxit eum et consecravit;
LEV|8|13|filios quoque eius applicatos vestivit subuculis lineis et cinxit balteo imposuitque mitras, ut iusserat Dominus Moysi.
LEV|8|14|Adduxit et vitulum pro peccato; cumque super caput eius posuissent Aaron et filii eius manus suas,
LEV|8|15|immolavit eum; et hauriens Moyses sanguinem tincto digito tetigit cornua altaris per gyrum et mundavit illud; fuditque reliquum sanguinem ad fundamenta eius et sanctificavit illud expiando.
LEV|8|16|Adipem autem, qui erat super vitalia, et reticulum iecoris duosque renunculos cum arvinulis suis adolevit super altare;
LEV|8|17|vitulum cum pelle, carnibus et fimo cremans extra castra, sicut praeceperat Dominus Moysi.
LEV|8|18|Attulit et arietem in holocaustum, super cuius caput cum imposuissent Aaron et filii eius manus suas,
LEV|8|19|immolavit eum et fudit sanguinem eius per altaris circuitum.
LEV|8|20|Ipsumque arietem in frusta concidens, caput eius et artus et adipem adolevit igni;
LEV|8|21|lotis prius intestinis et pedibus, totumque simul arietem adolevit super altare, eo quod esset holocaustum suavissimi odoris, incensum Domino, sicut praeceperat Dominus Moysi.
LEV|8|22|Attulit et arietem secundum in consecrationem sacerdotum; posueruntque super caput illius Aaron et filii eius manus suas.
LEV|8|23|Quem cum immolasset Moyses, sumens de sanguine tetigit extremum auriculae dextrae Aaron et pollicem manus eius dextrae, similiter et pedis.
LEV|8|24|Applicavit et filios Aaron; cumque de sanguine arietis immolati tetigisset extremum auriculae singulorum dextrae et pollices manus ac pedis dextri, reliquum fudit super altare per circuitum.
LEV|8|25|Tulitque adipem et caudam omnemque pinguedinem, quae operit intestina reticulumque iecoris, et duos renes cum adipibus suis et armo dextro.
LEV|8|26|Tollens autem de canistro azymorum, quod erat coram Domino, panem absque fermento et collyridam conspersam oleo laganumque posuit super adipes et armum dextrum,
LEV|8|27|tradens simul omnia super manus Aaron et filiorum eius. Qui, postquam levaverunt ea coram Domino,
LEV|8|28|rursum suscepta de manibus eorum adolevit in altari super holocausto, eo quod illa essent consecrationis oblatio, in odorem suavitatis: incensum erat Domino.
LEV|8|29|Tulit et pectusculum elevans illud coram Domino de ariete consecrationis in partem suam, sicut praeceperat Dominus Moysi.
LEV|8|30|Assumensque de unguento et sanguine, qui erat in altari, aspersit super Aaron et vestimenta eius et super filios illius ac vestes eorum.
LEV|8|31|Cumque sanctificasset eos in vestitu suo, praecepit eis dicens: " Coquite carnes ante fores tabernaculi et ibi comedite eas; panes quoque consecrationis edite, qui positi sunt in canistro, sicut mihi praeceptum est: "Aaron et filii eius comedent eos;
LEV|8|32|quidquid autem reliquum fuerit de carne et panibus, ignis absumet".
LEV|8|33|De ostio quoque tabernaculi conventus non exibitis septem diebus usque ad diem, quo complebitur tempus consecrationis vestrae; septem enim diebus finitur consecratio.
LEV|8|34|Sicut et impraesentiarum factum est, praecepit Dominus, ut fieret in expiationem eorum.
LEV|8|35|Die ac nocte manebitis in ostio tabernaculi conventus observantes observationem Domini, ne moriamini: sic enim mihi praeceptum est ".
LEV|8|36|Feceruntque Aaron et filii eius cuncta, quae locutus est Dominus per manum Moysi.
LEV|9|1|Facto autem octavo die, vocavit Moyses Aaron et filios eius ac maiores natu Israel dixitque ad Aaron:
LEV|9|2|" Tolle de armento vitulum pro peccato et arietem in holocaustum, utrumque immaculatum, et affer illos coram Domino.
LEV|9|3|Et ad filios Israel loqueris: "Tollite hircum pro peccato et vitulum atque agnum anniculos et sine macula in holocaustum,
LEV|9|4|bovem et arietem pro pacificis, et immolate eos coram Domino, et sacrificium similae oleo conspersae: hodie enim Dominus apparebit vobis" ".
LEV|9|5|Tulerunt ergo cuncta, quae iusserat Moyses, ad ostium tabernaculi conventus; ubi, cum omnis coetus accessisset et staret coram Domino,
LEV|9|6|ait Moyses: " Iste est sermo, quem praecepit Dominus: facite, et apparebit vobis gloria eius ".
LEV|9|7|Dixit et ad Aaron: " Accede ad altare et immola pro peccato tuo; offer holocaustum et expia te et populum. Et fac hostiam populi et expia eum, sicut praecepit Dominus ".
LEV|9|8|Statimque Aaron accedens ad altare immolavit vitulum pro peccato suo,
LEV|9|9|cuius sanguinem obtulerunt ei filii sui; in quo tinguens digitum tetigit cornua altaris et fudit residuum ad basim eius.
LEV|9|10|Adipemque et renunculos ac reticulum iecoris, quae sunt de sacrificio pro peccato, adolevit super altare, sicut praeceperat Dominus Moysi.
LEV|9|11|Carnes vero et pellem eius extra castra combussit igni.
LEV|9|12|Immolavit et holocausti victimam; obtuleruntque ei filii sui sanguinem eius, quem fudit per altaris circuitum.
LEV|9|13|Ipsam etiam hostiam in frusta concisam cum capite ei obtulerunt, quae omnia super altare cremavit igni;
LEV|9|14|lavit quoque aqua intestina cruraque et adolevit super holocausto in altari.
LEV|9|15|Et applicavit oblationem populi sumensque hircum pro peccato populi mactavit et obtulit in expiationem sicut priorem;
LEV|9|16|fecit quoque holocaustum secundum ritum
LEV|9|17|et addens sacrificium similae implevit manum ex illa et adolevit super altare praeter holocaustum matutinum.
LEV|9|18|Immolavit et bovem atque arietem, hostias pacificas populi; obtuleruntque ei filii sui sanguinem, quem fudit super altare in circuitu.
LEV|9|19|Adipes autem bovis et caudam arietis renunculosque cum adipibus suis et reticulum iecoris
LEV|9|20|posuerunt super pectora; cumque cremati essent adipes in altari,
LEV|9|21|pectora eorum et armos dextros Aaron elevavit coram Domino, sicut praeceperat Moyses.
LEV|9|22|Et elevans Aaron manus ad populum benedixit eis. Sicque, completis hostiis pro peccato et holocaustis et pacificis, descendit.
LEV|9|23|Ingressi autem Moyses et Aaron tabernaculum conventus et deinceps egressi benedixerunt populo. Apparuitque gloria Domini omni populo;
LEV|9|24|et ecce egressus ignis a Domino devoravit holocaustum et adipes, qui erant super altare. Quod cum vidissent turbae, exultaverunt ruentes in facies suas.
LEV|10|1|Arreptisque Nadab et Abiu filii Aaron turibulis, posue runt ignem et incensum desuper offerentes coram Domino ignem alienum, qui eis praeceptus non erat.
LEV|10|2|Egressusque ignis a Domino devoravit eos, et mortui sunt coram Domino.
LEV|10|3|Dixitque Moyses ad Aaron: " Hoc est, quod locutus est Dominus: "Sanctificabor in his, qui appropinquant mihi, et in conspectu omnis populi glorificabor" ". Quod audiens tacuit Aaron.
LEV|10|4|Vocatis autem Moyses Misael et Elisaphan filiis Oziel patrui Aaron, ait ad eos: " Ite et tollite fratres vestros de conspectu sanctuarii et asportate extra castra ".
LEV|10|5|Confestimque pergentes tulerunt eos, sicut iacebant vestitos subuculis suis, foras, ut sibi fuerat imperatum.
LEV|10|6|Locutus est Moyses ad Aaron et ad Eleazar atque Ithamar filios eius: " Comas vestras nolite excutere et vestimenta nolite scindere, ne moriamini, et super omnem coetum oriatur indignatio. Fratres vestri, omnis domus Israel, plangant incendium, quod Dominus suscitavit.
LEV|10|7|Vos autem non egredimini fores tabernaculi conventus, alioquin peribitis; oleum quippe unctionis Domini est super vos ". Qui fecerunt omnia iuxta praeceptum Moysi.
LEV|10|8|Dixit quoque Dominus ad Aaron:
LEV|10|9|" Vinum et omne, quod inebriare potest, non bibetis tu et filii tui, quando intratis tabernaculum conventus, ne moriamini ­ praeceptum est sempiternum in generationes vestras ­
LEV|10|10|et ut habeatis scientiam discernendi inter sanctum et profanum, inter pollutum et mundum,
LEV|10|11|doceatisque filios Israel omnia legitima mea, quae locutus est Dominus ad eos per manum Moysi ".
LEV|10|12|Locutusque est Moyses ad Aaron et ad Eleazar atque Ithamar filios eius, qui residui erant: " Tollite oblationem similae, quae remansit de incensis Domini, et comedite illam absque fermento iuxta altare, quia sanctum sanctorum est.
LEV|10|13|Comedetis autem in loco sancto, quia data est tibi et filiis tuis de incensis Domini, sicut praeceptum est mihi.
LEV|10|14|Pectusculum quoque elationis et armum donationis edetis in loco mundissimo, tu et filii tui ac filiae tuae tecum; tibi enim ac liberis tuis reposita sunt de hostiis pacificis filiorum Israel.
LEV|10|15|Armum et pectus cum incensis adipum afferent ad elationem coram Domino, et pertineant ad te et ad filios tuos lege perpetua, sicut praecepit Dominus ".
LEV|10|16|De hirco autem pro peccato cum quaereret Moyses, exustum repperit; iratusque contra Eleazar et Ithamar filios Aaron, qui remanserant, ait:
LEV|10|17|" Cur non comedistis sacrificium pro peccato in loco sancto? Quod sanctum sanctorum est, et datum vobis, ut portetis iniquitatem coetus in expiationem eorum in conspectu Domini;
LEV|10|18|praesertim cum de sanguine illius non sit illatum intra sancta, comedere eam debuistis in sanctuario, sicut praeceptum est mihi ".
LEV|10|19|Respondit Aaron: " Oblata est hodie victima pro peccato et holocaustum eorum coram Domino; mihi autem accidit, quod vides. Quomodo potui comedere eam et placere Domino? ".
LEV|10|20|Quod cum audisset Moyses, recepit satisfactionem.
LEV|11|1|Locutus est Dominus ad Moysen et Aaron dicens:
LEV|11|2|" Dicite filiis Israel: Haec sunt animalia, quae comedere debetis de cunctis animantibus terrae.
LEV|11|3|Omne, quod habet plene divisam ungulam et ruminat in pecoribus, comedetis.
LEV|11|4|Haec autem non comedetis ex ruminantibus vel dividentibus ungulam: camelum, quia ruminat quidem, sed non dividit ungulam, inter immunda reputabis;
LEV|11|5|hyracem, qui ruminat ungulamque non dividit, immundus est;
LEV|11|6|leporem quoque, nam et ipse ruminat, sed ungulam non dividit;
LEV|11|7|et suem, qui, cum ungulam plene dividat, non ruminat.
LEV|11|8|Horum carnibus non vescemini nec cadavera contingetis, quia immunda sunt vobis.
LEV|11|9|Haec sunt, quae gignuntur in aquis et vesci licitum est: omne, quod habet pinnulas et squamas, tam in mari quam in fluminibus et torrentibus, comedetis.
LEV|11|10|Quidquid autem pinnulas et squamas non habet, reptilium vel quorumlibet aliorum animalium, quae in aquis moventur, abominabile vobis
LEV|11|11|et execrandum erit; carnes eorum non comedetis et morticina vitabitis.
LEV|11|12|Cuncta, quae non habent pinnulas et squamas in aquis, polluta erunt vobis.
LEV|11|13|Haec sunt, quae de avibus comedere non debetis, et vitanda sunt vobis: aquilam et grypem et haliaeetum,
LEV|11|14|milvum ac vulturem iuxta genus suum
LEV|11|15|et omne corvini generis,
LEV|11|16|struthionem et noctuam et larum et accipitrem iuxta genus suum,
LEV|11|17|bubonem et mergulum et ibin,
LEV|11|18|cycnum et nyctocoracem et porphyrionem,
LEV|11|19|erodionem et charadrion iuxta genus suum, upupam quoque et vespertilionem.
LEV|11|20|Omne de volucribus, quod reptat super quattuor pedes, abominabile erit vobis.
LEV|11|21|Quidquid autem ambulat quidem super quattuor pedes, sed habet longiora retro crura, per quae salit super terram,
LEV|11|22|comedere debetis; ut est bruchus in genere suo et attacus atque ophiomachus ac locusta, singula iuxta genus suum.
LEV|11|23|Quidquid autem ex volucribus reptantibus quattuor tantum habet pedes, execrabile erit vobis.
LEV|11|24|Et quicumque morticina eorum tetigerit, polluetur et erit immundus usque ad vesperum.
LEV|11|25|Et si necesse fuerit, ut portet quippiam horum mortuum, lavabit vestimenta sua et immundus erit usque ad solis occasum.
LEV|11|26|Omne animal, quod habet quidem ungulam, sed non dividit eam nec ruminat, immundum erit vobis; et, qui tetigerit illud, contaminabitur.
LEV|11|27|Quod ambulat super plantas pedum ex cunctis animantibus, quae incedunt quadrupedia, immundum erit; qui tetigerit morticina eorum, polluetur usque ad vesperum.
LEV|11|28|Et, qui portaverit huiuscemodi cadavera, lavabit vestimenta sua et immundus erit usque ad vesperum; quia omnia haec immunda sunt vobis.
LEV|11|29|Haec quoque inter polluta reputabuntur de his, quae reptant in terra: mustela et mus et lacerta iuxta genus suum,
LEV|11|30|mygale et testudo et stellio et talpa et chamaeleon:
LEV|11|31|omnia haec immunda sunt.Qui tetigerit morticina eorum, immundus erit usque ad vesperum;
LEV|11|32|et super quod ceciderit quidquam de morticinis eorum, polluetur tam vas ligneum et vestimentum quam pelles et cilicia, et in quocumque fit opus; tinguentur aqua et polluta erunt usque ad vesperum et postea munda.
LEV|11|33|Vas autem fictile, in quo horum quidquam intro ceciderit, polluetur et frangendum est.
LEV|11|34|Omnis cibus, quem comedetis, si fusa fuerit exinde super eum aqua, immundus erit; et omne liquens, quod bibitur de tali vase, immundum erit.
LEV|11|35|Et quidquid de morticinis istiusmodi ceciderit super illud, immundum erit; sive clibani sive chytropodes destruentur: immundi sunt et immundi erunt vobis.
LEV|11|36|Fontes tamen et cisternae et omnis aquarum congregatio munda erit. Qui vero morticinum eorum tetigerit, polluetur.
LEV|11|37|Si ceciderint super sementem, non polluent eam;
LEV|11|38|sin autem quispiam aqua sementem perfuderit, et postea morticinis tacta fuerit, immunda erit vobis.
LEV|11|39|Si mortuum fuerit animal, quod licet vobis comedere, qui cadaver eius tetigerit, immundus erit usque ad vesperum;
LEV|11|40|et, qui comederit ex eo quippiam sive portaverit cadaver eius, lavabit vestimenta sua et immundus erit usque ad vesperum.
LEV|11|41|Omne, quod reptat super terram, abominabile erit nec assumetur in cibum.
LEV|11|42|Quidquid super pectus et quidquid quadrupes graditur, vel multos habet pedes sive per humum trahitur, non comedetis, quia abominabile est.
LEV|11|43|Nolite contaminare animas vestras nec tangatis quidquam eorum, ne immundi sitis.
LEV|11|44|Ego enim sum Dominus Deus vester; sanctificamini et sancti estote, quoniam et ego sanctus sum. Ne polluatis animas vestras in omni reptili, quod movetur super terram.
LEV|11|45|Ego enim sum Dominus, qui eduxi vos de terra Aegypti, ut essem vobis in Deum: sancti eritis, quia et ego sanctus sum.
LEV|11|46|Ista est lex animantium et volucrum et omnis animae viventis, quae movetur in aqua et reptat in terra,
LEV|11|47|ut differentias noveritis mundi et immundi, et sciatis quid comedere et quid respuere debeatis ".
LEV|12|1|Locutus est Dominus ad Moysen dicens:
LEV|12|2|" Loquere fi liis Israel et dices ad eos: Mulier, si, suscepto semine, pepererit masculum, immunda erit septem diebus iuxta dies separationis menstruae,
LEV|12|3|et die octavo circumcidetur infantulus;
LEV|12|4|ipsa vero triginta tribus diebus manebit in sanguine purificationis suae; omne sanctum non tanget nec ingredietur sanctuarium, donec impleantur dies purificationis eius.
LEV|12|5|Sin autem feminam pepererit, immunda erit duabus hebdomadibus iuxta ritum fluxus menstrui, et sexaginta ac sex diebus manebit in sanguine purificationis suae.
LEV|12|6|Cumque expleti fuerint dies purificationis suae pro filio sive pro filia, deferet agnum anniculum in holocaustum et pullum columbae sive turturem pro peccato ad ostium tabernaculi conventus et tradet sacerdoti.
LEV|12|7|Qui offeret illa coram Domino et expiabit eam; et sic mundabitur a profluvio sanguinis sui: ista est lex parientis masculum aut feminam.
LEV|12|8|Quod si non invenerit manus eius, nec potuerit offerre agnum, sumet duos turtures vel duos pullos columbae, unum in holocaustum et alterum pro peccato; expiabitque eam sacerdos, et sic mundabitur ".
LEV|13|1|Locutus est Dominus ad Moysen et Aaron dicens:
LEV|13|2|" Homo, in cuius carne et cute ortus fuerit tumor sive pustula aut quasi lucens quippiam, id est plaga leprae, adducetur ad Aaron sacerdotem vel ad unum quemlibet filiorum eius sacerdotum.
LEV|13|3|Qui cum viderit plagam in cute et pilos in album mutatos colorem ipsamque speciem plagae humiliorem cute et carne reliqua: plaga leprae est; quod cum viderit sacerdos, eum immundum esse decernet.
LEV|13|4|Sin autem lucens candor fuerit in cute nec humilior carne reliqua, et pili coloris pristini, recludet eum sacerdos septem diebus.
LEV|13|5|Et considerabit eum die septimo: et, siquidem plaga ultra non creverit nec transierit in cute priores terminos, rursum recludet eum septem diebus aliis.
LEV|13|6|Et die septimo contemplabitur eum iterum: si obscurior fuerit plaga et non creverit in cute, eum mundum esse decernet, quia scabies est. Lavabitque homo vestimenta sua et mundus erit.
LEV|13|7|Quod si, postquam a sacerdote visus est et redditus munditiae, iterum scabies creverit, adducetur ad eum;
LEV|13|8|et, si viderit ita esse, immunditiae condemnabitur: est lepra.
LEV|13|9|Plaga leprae si fuerit in homine, adducetur ad sacerdotem,
LEV|13|10|et videbit eum. Cumque tumor albus in cute fuerit et capillorum mutaverit aspectum in album, caro quoque viva creverit in tumore,
LEV|13|11|lepra vetustissima iudicabitur atque inolita cuti. Contaminabit itaque eum sacerdos et non recludet, quia perspicue immunditia est.
LEV|13|12|Sin autem effloruerit discurrens lepra in cute et operuerit omnem cutem a capite usque ad pedes, quidquid sub aspectu oculorum cadit,
LEV|13|13|considerabit eum sacerdos et teneri lepra mundissima iudicabit, eo quod omnis in candorem versa sit, et idcirco homo mundus erit.
LEV|13|14|Quando vero caro vivens in eo apparuerit, immundus erit.
LEV|13|15|Quod cum sacerdos viderit, inter immundos reputabit; caro enim viva immunda est: lepra est.
LEV|13|16|Quod si rursum versa fuerit in alborem, veniet ad sacerdotem,
LEV|13|17|qui cum hoc consideraverit, eum mundum esse decernet.
LEV|13|18|Caro et cutis, in qua ulcus natum est et sanatum,
LEV|13|19|et in loco ulceris tumor apparuerit albus sive macula subrufa, ostendet se homo sacerdoti.
LEV|13|20|Qui cum viderit locum maculae humiliorem carne reliqua et pilos versos in candorem, contaminabit eum: plaga enim leprae orta est in ulcere.
LEV|13|21|Quod si pilus coloris est pristini et cicatrix subobscura et vicina carne non est humilior, recludet eum septem diebus.
LEV|13|22|Et, siquidem creverit, adiudicabit eum leprae;
LEV|13|23|sin autem steterit in loco suo macula nec creverit, ulceris est cicatrix, et sacerdos eum mundum esse decernet.
LEV|13|24|Vel si alicuius cutem ignis exusserit, et locus exustionis subrufam sive albam habuerit maculam,
LEV|13|25|considerabit eam sacerdos; et ecce pilus versus est in alborem, et locus eius reliqua cute humilior, contaminabit eum, quia plaga leprae in cicatrice orta est.
LEV|13|26|Quod si pilorum color non fuerit immutatus, nec humilior macula carne reliqua, et ipsa leprae species fuerit subobscura, recludet eum septem diebus.
LEV|13|27|Et die septimo contemplabitur eum; si creverit in cute macula, contaminabit eum: plaga est leprae;
LEV|13|28|sin autem in loco suo macula steterit non satis clara, tumor combustionis est, et idcirco mundabit eum, quia cicatrix est combusturae.
LEV|13|29|Vir sive mulier, in cuius capite vel barba germinarit plaga, videbit eam sacerdos.
LEV|13|30|Et, siquidem humilior fuerit locus carne reliqua, et capillus flavus solitoque subtilior, contaminabit eos, quia scabies est, lepra capitis vel barbae.
LEV|13|31|Sin autem viderit plagam scabiei aequalem vicinae carni nec capillum nigrum in ea, recludet eos septem diebus.
LEV|13|32|Et die septimo intuebitur plagam: si non creverit scabies, nec capillus flavus fuerit in ea, et locus plagae carni reliquae aequalis,
LEV|13|33|radetur homo absque loco maculae, et includet eum sacerdos septem diebus aliis.
LEV|13|34|Si die septimo visa fuerit stetisse plaga in loco suo nec humilior carne reliqua, mundabit eum sacerdos; lotisque vestibus mundus erit.
LEV|13|35|Sin autem post emundationem rursus creverit scabies in cute,
LEV|13|36|non quaeret amplius utrum capillus in flavum colorem sit commutatus, quia aperte immundus est.
LEV|13|37|Porro si steterit macula, et capilli nigri fuerint, noverit hominem esse sanatum et confidenter eum pronuntiet mundum.
LEV|13|38|Vir et mulier, in cuius cute maculae, maculae albae apparuerint,
LEV|13|39|intuebitur eos sacerdos. Si deprehenderit subobscurum alborem lucere in cute, sciat impetiginem ortam esse in cute; mundus est.
LEV|13|40|Vir, de cuius capite capilli fluunt, calvus ac mundus est;
LEV|13|41|et, si a fronte ceciderint pili, recalvaster et mundus est.
LEV|13|42|Sin autem in calvitio sive in recalvatione plaga alba vel subrufa fuerit exorta, lepra est capitis.
LEV|13|43|Sacerdos eum videbit, et ecce tumor plagae subrufus secundum aspectum leprae cutis carnis.
LEV|13|44|Vir maculatus est lepra, et sacerdos omnino decernet eum esse immundum; plaga est in capite eius.
LEV|13|45|Leprosus hac plaga percussus habebit vestimenta dissuta, comam capitis excussam, barbam contectam; clamabit: "Immundus! Immundus!".
LEV|13|46|Omni tempore, quo leprosus est immundus, immundus est et solus habitabit extra castra.
LEV|13|47|Si in veste lanea sive linea lepra fuerit,
LEV|13|48|in stamine sive subtemine lineo vel laneo aut in pelle vel quolibet ex pelle confecto,
LEV|13|49|si macula pallida aut rufa fuerit, lepra reputabitur ostendeturque sacerdoti.
LEV|13|50|Qui considerabit macula infectum et recludet septem diebus;
LEV|13|51|et die septimo rursus aspiciens, si crevisse deprehenderit, lepra maligna est; pollutum iudicabit vestimentum et omne, in quo fuerit inventa,
LEV|13|52|et idcirco comburetur flammis.
LEV|13|53|Quod si eam viderit non crevisse,
LEV|13|54|praecipiet, et lavabunt id, in quo plaga est; recludetque illud septem diebus aliis.
LEV|13|55|Et cum viderit post lavationem faciem quidem pristinam non mutatam, nec tamen crevisse plagam, immunda est res, et igne combures eam, eo quod infusa sit plaga in superficie rei vel in parte aversa.
LEV|13|56|Sin autem obscurior fuerit locus plagae, postquam res est lota, sacerdos abrumpet eum et a solido dividet.
LEV|13|57|Quod si macula ultra apparuerit in his rebus, quae prius immaculata erant, lepra volatilis et vaga, igne combures illas.
LEV|13|58|Quas vero laveris et a quibus cessaverit plaga, illas lavabis secundo, et mundae erunt.
LEV|13|59|Ista est lex leprae vestimenti lanei et linei, staminis atque subteminis, omnisque supellectilis pelliceae, quomodo mundari debeat vel contaminari ".
LEV|14|1|Locutusque est Dominus ad Moysen dicens:
LEV|14|2|" Hic est ri tus leprosi, quando mundandus est: adducetur ad sacerdotem,
LEV|14|3|qui egressus e castris, cum invenerit lepram esse sanatam,
LEV|14|4|praecipiet, ut sumant pro eo, qui purificatur, duas aves vivas, mundas et lignum cedrinum vermiculumque et hyssopum.
LEV|14|5|Et unam ex avibus immolari iubebit in vase fictili super aquas viventes.
LEV|14|6|Aliam autem vivam cum ligno cedrino et cocco et hyssopo tinguet in sanguine avis super aquas viventes immolatae,
LEV|14|7|quo asperget illum, qui a lepra mundandus est, septies, ut iure purgetur; et dimittet avem vivam, ut in agrum avolet.
LEV|14|8|Cumque laverit homo vestimenta sua, radet omnes pilos corporis, et lavabitur aqua; purificatusque ingredietur castra, ita dumtaxat ut maneat extra tabernaculum suum septem diebus.
LEV|14|9|Et die septimo radet capillos capitis barbamque et supercilia ac totius corporis pilos et lavabit vestimenta carnemque suam aqua, et mundus erit.
LEV|14|10|Die octavo assumet duos agnos immaculatos et ovem anniculam absque macula et tres decimas ephi similae in sacrificium, quae conspersa sit oleo, et log olei.
LEV|14|11|Cumque sacerdos purificans hominem statuerit eum et haec omnia coram Domino in ostio tabernaculi conventus,
LEV|14|12|tollet agnum unum et offeret eum in sacrificium pro delicto, oleique log et, elevatis ante Dominum omnibus,
LEV|14|13|immolabit agnum, ubi immolari solet hostia pro peccato et holocaustum, id est in loco sancto. Sicut enim pro peccato ita et pro delicto ad sacerdotem pertinet sacrificium: sanctum sanctorum est.
LEV|14|14|Assumensque sacerdos de sanguine hostiae pro delicto ponet super extremum auriculae dextrae eius, qui mundatur, et super pollices manus dextrae et pedis;
LEV|14|15|et de olei log mittet in manum suam sinistram
LEV|14|16|tinguetque digitum dextrum in eo et asperget septies coram Domino.
LEV|14|17|Quod autem reliquum est olei in laeva manu, fundet super extremum auriculae dextrae eius, qui mundatur, et super pollices manus ac pedis dextri et super sanguinem sacrificii pro delicto
LEV|14|18|et super caput eius, qui mundatur; expiabitque eum coram Domino
LEV|14|19|et faciet sacrificium pro peccato. Tunc immolabit holocaustum
LEV|14|20|et ponet illud in altari cum sacrificio similae, et homo rite mundabitur.
LEV|14|21|Quod si pauper est, et non potest manus eius invenire, quae dicta sunt, assumet agnum pro delicto ad elationem, ut expiet eum sacerdos, decimamque partem similae conspersae oleo in sacrificium et olei log
LEV|14|22|duosque turtures sive duos pullos columbae, quos manus eius invenire poterit, unum pro peccato et alterum in holocaustum.
LEV|14|23|Offeretque ea die octavo purificationis suae sacerdoti ad ostium tabernaculi conventus coram Domino.
LEV|14|24|Qui suscipiens agnum pro delicto et log olei levabit simul coram Domino;
LEV|14|25|immolatoque agno pro delicto, de sanguine eius ponet super extremum auriculae dextrae illius, qui mundatur, et super pollices manus eius ac pedis dextri;
LEV|14|26|olei vero partem mittet in manum suam sinistram.
LEV|14|27|In quo tinguens digitum dextrae manus asperget septies coram Domino;
LEV|14|28|tangetque extremum auriculae dextrae illius, qui mundatur, et pollices manus ac pedis dextri super locum sanguinis, qui effusus est pro delicto.
LEV|14|29|Reliquam autem partem olei, quae est in sinistra manu, mittet super caput hominis, qui purificatur, in expiationem eius coram Domino;
LEV|14|30|et turtures sive pullos columbae, quos manus illius invenerit, offeret,
LEV|14|31|unum pro delicto et alterum in holocaustum cum sacrificio similae, et sic expiabit eum sacerdos coram Domino.
LEV|14|32|Hoc est sacrificium leprosi, qui habere non potest omnia in emundationem sui ".
LEV|14|33|Locutus est Dominus ad Moysen et Aaron dicens:
LEV|14|34|" Cum ingressi fueritis terram Chanaan, quam ego dabo vobis in possessionem, si fuerit plaga leprae in aedibus terrae possessionis vestrae,
LEV|14|35|ibit, cuius est domus, nuntians sacerdoti et dicet: "Quasi plaga videtur mihi esse in domo mea".
LEV|14|36|At ille praecipiet, ut efferant universa de domo, priusquam ingrediatur eam, et videat plagam, ne immunda fiant omnia, quae in domo sunt. Intrabitque postea, ut consideret domum;
LEV|14|37|et, cum viderit in parietibus illius quasi valliculas pallore sive rubore deformes et humiliores superficie reliqua,
LEV|14|38|egredietur ostium domus et statim claudet eam septem diebus.
LEV|14|39|Reversusque die septimo considerabit eam; si invenerit crevisse plagam,
LEV|14|40|iubebit erui lapides, in quibus plaga est, et proici eos extra civitatem in loco immundo;
LEV|14|41|domum autem ipsam radi intrinsecus per circuitum et spargi pulverem rasurae extra urbem in locum immundum
LEV|14|42|lapidesque alios reponi pro his, qui ablati fuerint, et luto alio liniri domum.
LEV|14|43|Sin autem plaga rursum effloruerit in domo, postquam eruti sunt lapides et pulvis erasus et alia terra lita,
LEV|14|44|et ingressus sacerdos viderit crevisse plagam in domo: lepra est maligna et domus immunda.
LEV|14|45|Quam statim destruent et lapides eius ac ligna atque universum pulverem domus proicient extra oppidum in loco immundo.
LEV|14|46|Qui intraverit domum, quando clausa est, immundus erit usque ad vesperum;
LEV|14|47|et, qui dormierit in ea vel comederit quippiam, lavabit vestimenta sua.
LEV|14|48|Quod si introiens sacerdos viderit plagam non crevisse in domo, postquam denuo lita est, mundam eam esse decernet, reddita sanitate.
LEV|14|49|Et in purificationem eius sumet duas aves lignumque cedrinum et vermiculum atque hyssopum
LEV|14|50|et, immolata una avi in vase fictili super aquas vivas,
LEV|14|51|tollet lignum cedrinum et hyssopum et coccum et avem vivam et intinguet omnia in sanguine avis immolatae atque in aquis viventibus et asperget domum septies;
LEV|14|52|purificabitque eam tam in sanguine avis quam in aquis viventibus et in avi viva lignoque cedrino et hyssopo atque vermiculo;
LEV|14|53|cumque dimiserit avem avolare extra urbem in agrum libere, expiabit domum, et erit munda.
LEV|14|54|Ista est lex omnis leprae et scabiei,
LEV|14|55|leprae vestium et domorum,
LEV|14|56|tumoris et pustulae et lucentis maculae,
LEV|14|57|ut possit sciri quo tempore immundum quid vel mundum sit ".
LEV|15|1|Locutus est Dominus ad Moysen et Aaron dicens:
LEV|15|2|" Loquimini filiis Israel et dicite eis: Vir, si patitur fluxum seminis, immundus erit.
LEV|15|3|Et tunc iudicabitur huic vitio subiacere: sive emiserit caro eius fluxum suum vel occluserit se a fluxu.
LEV|15|4|Omne stratum, in quo iacuerit, immundum erit, et ubicumque sederit.
LEV|15|5|Si quis hominum tetigerit lectum eius, lavabit vestimenta sua, et ipse lotus aqua immundus erit usque ad vesperum.
LEV|15|6|Si sederit, ubi ille sederat, et ipse lavabit vestimenta sua et lotus aqua immundus erit usque ad vesperum.
LEV|15|7|Qui tetigerit carnem eius, lavabit vestimenta sua et ipse lotus aqua immundus erit usque ad vesperum.
LEV|15|8|Si salivam huiuscemodi homo iecerit super eum, qui mundus est, hic lavabit vestem suam et lotus aqua immundus erit usque ad vesperum.
LEV|15|9|Sagma, super quo sederit, immundum erit;
LEV|15|10|et quicumque tetigerit omne, quod sub eo fuerit, qui fluxum seminis patitur, pollutus erit usque ad vesperum. Qui portaverit horum aliquid, lavabit vestem suam et ipse lotus aqua immundus erit usque ad vesperum.
LEV|15|11|Omnis, quem tetigerit, qui fluxum patitur, non lotis ante manibus, lavabit vestimenta sua et lotus aqua immundus erit usque ad vesperum.
LEV|15|12|Vas fictile, quod tetigerit, confringetur; vas autem ligneum lavabitur aqua.
LEV|15|13|Si sanatus fuerit, qui huiuscemodi sustinet passionem, numerabit septem dies ad emundationem sui et, lotis vestibus ac toto corpore in aquis viventibus, erit mundus.
LEV|15|14|Die autem octavo sumet duos turtures aut duos pullos columbae et veniet in conspectu Domini ad ostium tabernaculi conventus dabitque eos sacerdoti.
LEV|15|15|Qui faciet unum in sacrificium pro peccato et alterum in holocaustum; expiabitque eum coram Domino et emundabitur a fluxu seminis sui.
LEV|15|16|Vir, de quo egreditur semen, lavabit aqua omne corpus suum et immundus erit usque ad vesperum.
LEV|15|17|Vestem et pellem, super quam fuerit semen effusum, lavabitur aqua et immunda erit usque ad vesperum.
LEV|15|18|Si cum muliere coierit vir, lavabunt se aqua et immundi erunt usque ad vesperum.
LEV|15|19|Mulier, quae redeunte mense patitur fluxum sanguinis, septem diebus separabitur. Omnis, qui tetigerit eam, immundus erit usque ad vesperum;
LEV|15|20|et in quo iacuerit vel sederit diebus separationis suae, polluetur.
LEV|15|21|Qui tetigerit lectum eius, lavabit vestimenta sua et ipse lotus aqua immundus erit usque ad vesperum.
LEV|15|22|Omne vas, super quo illa sederit, quisquis attigerit, lavabit vestimenta sua et ipse lotus aqua pollutus erit usque ad vesperum.
LEV|15|23|Et quicumque tetigerit omne, quod fuerit super lectum vel supellectilem, in qua illa sederit, immundus erit usque ad vesperum.
LEV|15|24|Si coierit cum ea vir tempore sanguinis menstrualis, immundus erit septem diebus, et omne stratum, in quo dormierit, polluetur.
LEV|15|25|Mulier, quae patitur multis diebus fluxum sanguinis non in tempore menstruali vel quae post menstruum sanguinem fluere non cessat, quamdiu huic subiacet passioni, immunda erit quasi sit in tempore menstruo.
LEV|15|26|Omne stratum, in quo dormierit, et vas, in quo sederit, pollutum erit.
LEV|15|27|Quicumque tetigerit ea, polluetur; lavabit vestimenta sua et ipse lotus aqua immundus erit usque ad vesperum.
LEV|15|28|Si steterit sanguis et fluere cessarit, numerabit septem dies et deinde munda erit.
LEV|15|29|Et octavo die assumet pro se duos turtures vel duos pullos columbae afferetque sacerdoti ad ostium tabernaculi conventus.
LEV|15|30|Qui unum faciet in sacrificium pro peccato et alterum in holocaustum; expiabitque eam coram Domino a fluxu immunditiae eius.
LEV|15|31|Docebitis ergo filios Israel, ut caveant immunditiam, ne moriantur in sordibus suis, cum polluerint habitaculum meum, quod est inter eos.
LEV|15|32|Ista est lex eius, qui patitur fluxum seminis et de quo egreditur semen et polluitur,
LEV|15|33|et quae menstruis temporibus separatur vel quae iugi fluit sanguine, et hominis, qui dormierit cum immunda ".
LEV|16|1|Locutusque est Dominus ad Moysen post mortem duum filiorum Aaron, quando appropinquantes in conspectum Domini interfecti sunt,
LEV|16|2|et praecepit ei dicens: " Loquere ad Aaron fratrem tuum, ne omni tempore ingrediatur sanctuarium, quod est intra velum coram propitiatorio, quo tegitur arca, ut non moriatur, quia in nube apparebo super propitiatorium;
LEV|16|3|sed hoc modo ingrediatur: vitulum offeret pro peccato et arietem in holocaustum;
LEV|16|4|subucula linea sancta vestietur, feminalibus lineis verecunda celabit, accingetur zona linea, cidarim lineam imponet capiti. Haec enim vestimenta sunt sancta, quibus cunctis, cum lotus fuerit, induetur.
LEV|16|5|Suscipietque a coetu filiorum Israel duos hircos in sacrificium pro peccato et unum arietem in holocaustum.
LEV|16|6|Cumque obtulerit vitulum in sacrificium suum pro peccato et expiaverit se et domum suam,
LEV|16|7|duos hircos stare faciet coram Domino in ostio tabernaculi conventus,
LEV|16|8|mittens super utrumque sortem, unam Domino et alteram Azazel.
LEV|16|9|Cuius sors exierit Domino, offeret illum pro peccato;
LEV|16|10|cuius autem in Azazel, statuet eum vivum coram Domino in expiationem, ut emittat illum ad Azazel in solitudinem.
LEV|16|11|Afferet ergo Aaron vitulum pro peccato et expians se et domum suam immolabit eum;
LEV|16|12|assumptoque turibulo, quod de prunis altaris coram Domino impleverit, et hauriens manu compositum thymiama in incensum ultra velum intrabit in sancta,
LEV|16|13|ut, positis super ignem aromatibus coram Domino, nebula eorum et vapor operiat propitiatorium, quod est super testimonium, et non moriatur.
LEV|16|14|Tollet quoque de sanguine vituli et asperget digito septies contra frontem propitiatorii.
LEV|16|15|Cumque mactaverit hircum pro peccato populi, inferet sanguinem eius intra velum, sicut praeceptum est de sanguine vituli, ut aspergat e regione propitiatorii
LEV|16|16|et expiet sanctuarium ab immunditiis filiorum Israel et a praevaricationibus eorum cunctisque peccatis. Iuxta hunc ritum faciet tabernaculo conventus, quod fixum est inter eos in medio sordium habitationis eorum.
LEV|16|17|Nullus hominum sit in tabernaculo conventus, quando pontifex ingreditur sanctuarium, ut expiet se et domum suam et universam congregationem Israel, donec egrediatur.
LEV|16|18|Cum autem exierit ad altare, quod coram Domino est, expiabit illud et sumptum sanguinem vituli atque hirci fundet super cornua eius per gyrum;
LEV|16|19|aspergensque de sanguine digito septies mundabit sanctificabitque illud ab immunditiis filiorum Israel.
LEV|16|20|Et postquam compleverit expiationem sanctuarii et tabernaculi conventus et altaris, tunc afferat hircum viventem;
LEV|16|21|et, posita utraque manu super caput eius, confiteatur Aaron super eum omnes iniquitates filiorum Israel et universa delicta atque peccata eorum; quae ponens super caput eius emittet illum per hominem paratum in desertum.
LEV|16|22|Cumque portaverit hircus super se omnes iniquitates eorum in terram solitariam et dimissus fuerit in desertum,
LEV|16|23|ingredietur Aaron in tabernaculum conventus; et, depositis vestibus lineis, quibus prius indutus erat, cum intraret sanctuarium, relictisque ibi,
LEV|16|24|lavabit carnem suam aqua in loco sancto indueturque vestimentis suis. Et postquam egressus obtulerit holocaustum suum ac plebis, expiabit se et populum;
LEV|16|25|et adipem sacrificii pro peccato adolebit super altare.
LEV|16|26|Ille vero, qui dimiserit caprum emissarium ad Azazel, lavabit vestimenta sua et corpus aqua et postea ingredietur in castra.
LEV|16|27|Vitulum autem et hircum, qui pro peccato fuerant immolati, et quorum sanguis illatus est, ut in sanctuario expiatio compleretur, asportabunt foras castra et comburent igni tam pelles quam carnes eorum et fimum;
LEV|16|28|et quicumque combusserit ea, lavabit vestimenta sua et carnem aqua et postea ingredietur in castra.
LEV|16|29|Eritque hoc vobis legitimum sempiternum: mense septimo, decima die mensis affligetis animas vestras nullumque facietis opus sive indigena sive advena, qui peregrinatur inter vos.
LEV|16|30|In hac die expiatio erit vestri atque mundatio; ab omnibus peccatis vestris coram Domino mundabimini.
LEV|16|31|Sabbatum requietionis est vobis, et affligetis animas vestras religione perpetua.
LEV|16|32|Expiabit autem sacerdos, qui unctus fuerit, et cuius initiatae manus, ut sacerdotio fungatur pro patre suo; indueturque vestimentis lineis, vestibus sanctis,
LEV|16|33|et expiabit sanctuarium sanctissimum et tabernaculum conventus atque altare, sacerdotes quoque et universum populum congregationis.
LEV|16|34|Eritque hoc vobis legitimum sempiternum, ut expietis filios Israel a cunctis peccatis eorum semel in anno ".Fecit igitur, sicut praeceperat Dominus Moysi.
LEV|17|1|Et locutus est Dominus ad Moysen dicens:
LEV|17|2|" Loquere Aaron et filiis eius et cunctis filiis Israel et dices ad eos: Iste est sermo, quem mandavit Dominus dicens:
LEV|17|3|Homo quilibet de domo Israel, si occiderit bovem aut ovem sive capram in castris vel extra castra
LEV|17|4|et non attulerit ad ostium tabernaculi conventus in oblationem Domino coram habitaculo Domini, sanguinis reus erit; sanguinem fudit et peribit de medio populi sui.
LEV|17|5|Ideo offerre debent sacerdoti filii Israel hostias suas, quas occidunt in agro, ut afferant Domino ante ostium tabernaculi conventus et immolent eas hostias pacificas Domino.
LEV|17|6|Fundetque sacerdos sanguinem super altare Domini ad ostium tabernaculi conventus et adolebit adipem in odorem suavitatis Domino;
LEV|17|7|et nequaquam ultra immolabunt hostias suas daemonibus, cum quibus fornicati sunt: legitimum sempiternum erit hoc illis et posteris eorum ".
LEV|17|8|Et ad ipsos dices: " Homo de domo Israel et de advenis, qui peregrinantur apud vos, qui obtulerit holocaustum sive sacrificium
LEV|17|9|et ad ostium tabernaculi conventus non adduxerit victimam, ut offeratur Domino, interibit de populo suo.
LEV|17|10|Homo quilibet de domo Israel et de advenis, qui peregrinantur inter eos, si comederit sanguinem, confirmabo faciem meam contra talem animam et disperdam eam de populo suo.
LEV|17|11|Quia anima carnis in sanguine est, et ego dedi illum vobis, ut super altare in eo expietis pro animabus vestris, quia sanguis ipse per animam expiat.
LEV|17|12|Idcirco dixi filiis Israel: Omnis anima ex vobis non comedet sanguinem, nec ex advenis, qui peregrinantur inter vos.
LEV|17|13|Homo quicumque de filiis Israel et de advenis, qui peregrinantur apud vos, si venatione ceperit feram vel avem, quibus vesci licitum est, fundat sanguinem eius et operiat illum terra.
LEV|17|14|Anima enim omnis carnis, sanguis est anima eius, unde dixi filiis Israel: Sanguinem universae carnis non comedetis, quia anima omnis carnis sanguis eius est; et, quicumque comederit illum, interibit.
LEV|17|15|Anima, quae comederit morticinum vel captum a bestia, tam de indigenis quam de advenis, lavabit vestes suas et semetipsum aqua, et contaminatus erit usque ad vesperum; et hoc ordine mundus fiet.
LEV|17|16|Quod si non laverit vestimenta sua nec corpus, portabit iniquitatem suam ".
LEV|18|1|Locutus est Dominus ad Moysen dicens:
LEV|18|2|" Loquere fi liis Israel et dices ad eos: Ego Dominus Deus vester.
LEV|18|3|Iuxta consuetudinem terrae Aegypti, in qua habitastis, non facietis; et iuxta morem regionis Chanaan, ad quam ego introducturus sum vos, non agetis nec in legitimis eorum ambulabitis.
LEV|18|4|Facietis iudicia mea et praecepta mea servabitis et ambulabitis in eis. Ego Dominus Deus vester.
LEV|18|5|Custodite leges meas atque iudicia; quae faciens homo vivet in eis. Ego Dominus.
LEV|18|6|Omnis homo ad consanguineum suum non accedet, ut revelet turpitudinem eius. Ego Dominus.
LEV|18|7|Turpitudinem patris et turpitudinem matris tuae non discooperies: mater tua est, non revelabis turpitudinem eius.
LEV|18|8|Turpitudinem uxoris patris tui non discooperies, turpitudo enim patris tui est.
LEV|18|9|Turpitudinem sororis tuae ex patre sive ex matre, quae domi vel foris genita est, non revelabis.
LEV|18|10|Turpitudinem filiae filii tui vel neptis ex filia non revelabis, quia turpitudo tua est.
LEV|18|11|Turpitudinem filiae uxoris patris tui, quam peperit patri tuo et est soror tua, non revelabis.
LEV|18|12|Turpitudinem sororis patris tui non discooperies, quia caro est patris tui.
LEV|18|13|Turpitudinem sororis matris tuae non revelabis, eo quod caro sit matris tuae.
LEV|18|14|Turpitudinem patrui tui non revelabis nec accedes ad uxorem eius, quae tibi affinitate coniungitur.
LEV|18|15|Turpitudinem nurus tuae non revelabis, quia uxor filii tui est, nec discooperies ignominiam eius.
LEV|18|16|Turpitudinem uxoris fratris tui non revelabis, quia turpitudo fratris tui est.
LEV|18|17|Turpitudinem mulieris et filiae eius non revelabis. Filiam filii eius et filiam filiae illius non sumes, ut reveles ignominiam eius, quia caro illius sunt: nefas est.
LEV|18|18|Sororem uxoris tuae aemulam illius non accipies nec revelabis turpitudinem eius, adhuc illa vivente.
LEV|18|19|Ad mulierem, quae patitur menstrua, non accedes nec revelabis foeditatem eius.
LEV|18|20|Cum uxore proximi tui non coibis nec seminis commixtione maculaberis.
LEV|18|21|De semine tuo non dabis, ut consecretur idolo Moloch, nec pollues nomen Dei tui. Ego Dominus.
LEV|18|22|Cum masculo non commisceberis coitu femineo: abominatio est.
LEV|18|23|Cum omni pecore non coibis nec maculaberis cum eo. Mulier non succumbet iumento nec miscebitur ei, quia scelus est.
LEV|18|24|Ne polluamini in omnibus his, quibus contaminatae sunt universae gentes, quas ego eiciam ante conspectum vestrum
LEV|18|25|et quibus polluta est terra, cuius ego scelera visitavi, et evomuit habitatores suos.
LEV|18|26|Vos autem custodite legitima mea atque iudicia et non faciatis ex omnibus abominationibus istis tam indigena quam colonus, qui peregrinatur apud vos.
LEV|18|27|Omnes enim execrationes istas fecerunt accolae terrae, qui fuerunt ante vos, et polluerunt eam.
LEV|18|28|Cavete ergo, ne et vos similiter evomat, cum pollueritis eam, sicut evomuit gentem, quae fuit ante vos.
LEV|18|29|Omnis enim anima, quae fecerit de abominationibus his quippiam, peribit de medio populi sui.
LEV|18|30|Custodite mandata mea. Nolite facere legitima abominabilia, quae fecerunt hi, qui fuerunt ante vos, et ne polluamini in eis. Ego Dominus Deus vester ".
LEV|19|1|Locutus est Dominus ad Moysen dicens:
LEV|19|2|" Loquere ad omnem coetum filiorum Israel et dices ad eos: Sancti estote, quia sanctus sum ego, Dominus Deus vester.
LEV|19|3|Unusquisque matrem et patrem suum timeat. Sabbata mea custodite. Ego Dominus Deus vester.
LEV|19|4|Nolite converti ad idola nec deos conflatiles faciatis vobis. Ego Dominus Deus vester.
LEV|19|5|Si immolaveritis hostiam pacificorum Domino, immolabitis eam ita ut sit vobis placabilis.
LEV|19|6|Eo die, quo fuerit immolata, comedetur et die altero; quidquid autem residuum fuerit in diem tertium, igne comburetur.
LEV|19|7|Si quid post biduum comestum fuerit, profanum erit neque acceptabile.
LEV|19|8|Qui manducaverit illud, portabit iniquitatem suam, quia sanctum Domini polluit, et peribit anima illa de populo suo.
LEV|19|9|Cum messueris segetes terrae tuae, non tondebis usque ad marginem agri tui nec remanentes spicas colliges.
LEV|19|10|Neque in vinea tua racemos et grana decidentia congregabis, sed pauperibus et peregrinis carpenda dimittes. Ego Dominus Deus vester.
LEV|19|11|Non facietis furtum. Non mentiemini, nec decipiet unusquisque proximum suum.
LEV|19|12|Non periurabis in nomine meo nec pollues nomen Dei tui. Ego Dominus.
LEV|19|13|Non facies calumniam proximo tuo nec spoliabis eum. Non morabitur merces mercennarii apud te usque mane.
LEV|19|14|Non maledices surdo nec coram caeco pones offendiculum; sed timebis Deum tuum. Ego Dominus.
LEV|19|15|Non facietis, quod iniquum est in iudicio. Non consideres personam pauperis nec honores vultum potentis. Iuste iudica proximo tuo.
LEV|19|16|Non eris criminator et susurro in populo tuo. Non stabis contra sanguinem proximi tui. Ego Dominus.
LEV|19|17|Ne oderis fratrem tuum in corde tuo; argue eum, ne habeas super illo peccatum.
LEV|19|18|Non quaeres ultionem nec irasceris civibus tuis. Diliges proximum tuum sicut teipsum. Ego Dominus.
LEV|19|19|Leges meas custodite.Iumenta tua non facies coire cum alterius generis animantibus. Agrum tuum non seres diverso semine. Veste, quae ex duobus texta est, non indueris.
LEV|19|20|Homo, si dormierit cum muliere coitu seminis, quae sit ancilla destinata viro et tamen pretio non redempta nec libertate donata, vapulabunt ambo et non morientur, quia non fuit libera.
LEV|19|21|Et in sacrificium suum pro delicto offeret Domino ad ostium tabernaculi conventus arietem;
LEV|19|22|expiabitque eum sacerdos ariete a peccato eius coram Domino, et dimittetur ei peccatum, quod peccavit.
LEV|19|23|Quando ingressi fueritis terram et plantaveritis omnimoda ligna pomifera, non auferetis praeputia eorum, id est poma, quae germinant; tribus annis erunt vobis immunda ut praeputia, nec edetis ex eis.
LEV|19|24|Quarto anno omnis fructus eorum sanctificabitur laudabilis Domino.
LEV|19|25|Quinto autem anno comedetis fructus eorum, ut augeatur vobis proventus eorum. Ego Dominus Deus vester.
LEV|19|26|Non comedetis cum sanguine.Non augurabimini nec observabitis omina.
LEV|19|27|Neque in rotundum attondebitis marginem comae nec truncabis barbam.
LEV|19|28|Et super mortuo non incidetis carnem vestram neque figuras aliquas in cute incidetis vobis. Ego Dominus.
LEV|19|29|Ne polluas et prostituas filiam tuam, ne contaminetur terra et impleatur piaculo.
LEV|19|30|Sabbata mea custodite et sanctuarium meum metuite. Ego Dominus.
LEV|19|31|Non declinetis ad pythones nec ab hariolis aliquid sciscitemini, ut polluamini per eos. Ego Dominus Deus vester.
LEV|19|32|Coram cano capite consurge et honora personam senis; et time Deum tuum. Ego Dominus.
LEV|19|33|Si habitaverit tecum advena in terra vestra, non opprimetis eum;
LEV|19|34|sed sit inter vos quasi indigena, et diliges eum sicut teipsum: fuistis enim et vos advenae in terra Aegypti. Ego Dominus Deus vester.
LEV|19|35|Nolite facere iniquum aliquid in iudicio, in regula, in pondere, in mensura.
LEV|19|36|Statera iusta, aequa pondera, iustum ephi aequumque hin sint vobis. Ego Dominus Deus vester, qui eduxi vos de terra Aegypti.
LEV|19|37|Custodite omnia praecepta mea et universa iudicia et facite ea. Ego Dominus ".
LEV|20|1|Locutusque est Dominus ad Moysen dicens:
LEV|20|2|" Haec lo queris filiis Israel: Homo de filiis Israel et de advenis, qui habitant in Israel, si dederit de semine suo idolo Moloch, morte moriatur: populus terrae lapidabit eum.
LEV|20|3|Et ego ponam faciem meam contra illum; succidamque eum de medio populi sui, eo quod dederit de semine suo Moloch et contaminaverit sanctuarium meum ac polluerit nomen sanctum meum.
LEV|20|4|Quod si clauserit populus terrae oculos suos, ne videat hominem illum, qui dederit de semine suo Moloch, nec voluerit eum occidere,
LEV|20|5|ponam ego faciem meam super hominem illum et cognationem eius succidamque et ipsum et omnes, qui consenserunt ei, ut fornicarentur cum Moloch, de medio populi sui.
LEV|20|6|Anima, quae declinaverit ad pythones et hariolos et fornicata fuerit cum eis, ponam faciem meam contra eam et interficiam illam de medio populi sui.
LEV|20|7|Sanctificamini et estote sancti, quia ego Dominus Deus vester.
LEV|20|8|Custodite praecepta mea et facite ea. Ego Dominus, qui sanctifico vos.
LEV|20|9|Qui maledixerit patri suo et matri, morte moriatur; qui patri matrique maledixit, sanguis eius sit super eum.
LEV|20|10|Si moechatus quis fuerit cum uxore alterius et adulterium perpetrarit cum coniuge proximi sui, morte moriantur et moechus et adultera.
LEV|20|11|Qui dormierit cum noverca sua et revelaverit ignominiam patris sui, morte moriantur ambo: sanguis eorum sit super eos.
LEV|20|12|Si quis dormierit cum nuru sua, uterque moriatur, quia scelus operati sunt: sanguis eorum sit super eos.
LEV|20|13|Qui dormierit cum masculo coitu femineo, uterque operatus est nefas, morte moriantur: sit sanguis eorum super eos.
LEV|20|14|Qui supra uxorem filiam duxerit matrem eius, scelus operatus est: vivus ardebit cum eis, nec permanebit tantum nefas in medio vestri.
LEV|20|15|Qui cum iumento et pecore coierit, morte moriatur; pecus quoque occidite.
LEV|20|16|Mulier, quae succubuerit cuilibet iumento, simul interficies illam cum eo, morte moriantur: sanguis eorum sit super eos.
LEV|20|17|Qui acceperit sororem suam filiam patris sui vel filiam matris suae et viderit turpitudinem eius, illaque conspexerit fratris ignominiam, nefaria res est; occidentur in conspectu populi sui, eo quod turpitudinem sororis suae revelaverit, portabit iniquitatem suam.
LEV|20|18|Qui coierit cum muliere in fluxu menstruo et revelaverit turpitudinem eius ­ fontem eius nudavit, ipsaque aperuit fontem sanguinis sui ­ interficientur ambo de medio populi sui.
LEV|20|19|Turpitudinem materterae et amitae tuae non discooperies; qui hoc fecerit, ignominiam carnis suae nudavit; portabunt ambo iniquitatem suam.
LEV|20|20|Qui coierit cum uxore patrui vel avunculi sui et revelaverit ignominiam cognationis suae, portabunt ambo peccatum suum: absque liberis morientur.
LEV|20|21|Qui duxerit uxorem fratris sui, immunditia est, turpitudinem fratris sui revelavit: absque liberis erunt.
LEV|20|22|Custodite omnes leges meas atque omnia iudicia et facite ea, ne et vos evomat terra, quam intraturi estis et habitaturi.
LEV|20|23|Nolite ambulare in legitimis nationum, quas ego expulsurus sum ante vos. Omnia enim haec fecerunt, et abominatus sum eas
LEV|20|24|locutusque sum vobis: Vos possidebitis terram eorum, et ego dabo eam vobis in hereditatem, terram fluentem lacte et melle. Ego Dominus Deus vester, qui separavi vos a ceteris populis.
LEV|20|25|Separate ergo et vos iumentum mundum ab immundo et avem immundam a munda, ne polluatis animas vestras in pecore et in avibus et cunctis, quae moventur in terra, et quae vobis separavi tamquam immunda.
LEV|20|26|Eritis mihi sancti, quia sanctus sum ego Dominus et separavi vos a ceteris populis, ut essetis mei.
LEV|20|27|Vir sive mulier, in quibus pythonicus vel divinationis fuerit spiritus, morte moriantur; lapidibus obruent eos: sanguis eorum sit super illos ".
LEV|21|1|Dixit quoque Dominus ad Moysen: " Loquere ad sacer dotes filios Aaron et dices eis: Ne contaminetur sacerdos in mortibus civium suorum,
LEV|21|2|nisi tantum in consanguineis propinquis, id est super matre et patre et filio ac filia, fratre quoque
LEV|21|3|et sorore virgine propinqua, quae non est nupta viro; in ipsa contaminabitur.
LEV|21|4|Non contaminabitur ut maritus in cognatis suis, ne profanetur.
LEV|21|5|Non radent caput nec barbam neque in carne sua facient incisuras.
LEV|21|6|Sancti erunt Deo suo et non polluent nomen eius: incensa enim Domini et panem Dei sui offerunt et ideo sancti erunt.
LEV|21|7|Scortum et oppressam non ducent uxorem nec eam, quae repudiata est a marito, quia consecratus est Deo suo.
LEV|21|8|Et sanctificabis eum, quia panem Dei sui offert. Sit ergo sanctus tibi, quia ego sanctus sum, Dominus, qui sanctifico vos.
LEV|21|9|Sacerdotis filia, si profanaverit se stupro, profanat nomen patris sui; flammis exuretur.
LEV|21|10|Sacerdos maximus inter fratres suos, super cuius caput fusum est unctionis oleum, et cuius manus in sacerdotio consecratae sunt, vestitusque est sanctis vestibus, comam suam non excutiet, vestimenta non scindet
LEV|21|11|et ad omnem mortuum non ingredietur omnino; super patre quoque suo et matre non contaminabitur.
LEV|21|12|Nec egredietur de sanctuario, ne polluat sanctuarium Domini, quia consecratus est oleo unctionis Dei sui. Ego Dominus.
LEV|21|13|Virginem ducet uxorem;
LEV|21|14|viduam et repudiatam et oppressam atque meretricem non accipiet, sed virginem de cognatis suis ducet uxorem.
LEV|21|15|Ne profanet stirpem suam inter cognatos suos, quia ego Dominus, qui sanctifico eum ".
LEV|21|16|Locutusque est Dominus ad Moysen dicens:
LEV|21|17|" Loquere ad Aaron: Homo de semine tuo in generationibus suis, qui habuerit maculam, non accedet, ut offerat panem Dei sui;
LEV|21|18|quia quicumque habuerit maculam, non accedet: si caecus fuerit vel claudus, si mutilo naso vel deformis,
LEV|21|19|si fracto pede vel manu,
LEV|21|20|si gibbus, si pusillus, si albuginem habens in oculo, si iugem scabiem, si impetiginem in corpore vel contritos testiculos.
LEV|21|21|Omnis, qui habuerit maculam de semine Aaron sacerdotis, non accedet offerre incensa Domini nec panem Dei sui.
LEV|21|22|Vescetur tamen pane Dei sui de sanctissimis et de sanctis.
LEV|21|23|Sed ad velum non ingrediatur nec accedat ad altare, quia maculam habet et contaminare non debet sanctuaria mea, quia ego Dominus, qui sanctifico ea ".
LEV|21|24|Locutus est ergo Moyses ad Aaron et filios eius et ad omnem Israel.
LEV|22|1|Locutus quoque est Dominus ad Moysen dicens:
LEV|22|2|" Loquere ad Aaron et ad filios eius, ut caveant ab his, quae consecrata sunt filiorum Israel, et non contaminent nomen sanctum meum, quae ipsi offerunt mihi. Ego Dominus.
LEV|22|3|Dic ad eos pro posteris vestris: Omnis homo, qui accesserit de omni stirpe vestra ad sancta, quae consecraverunt filii Israel Domino, in immunditia sua, peribit coram me. Ego Dominus.
LEV|22|4|Homo de semine Aaron, qui fuerit leprosus aut patiens fluxum, non vescetur de his, quae sanctificata sunt, donec sanetur. Qui tetigerit omne, quod immundum est ex mor tuo, vel vir, ex quo egreditur semen,
LEV|22|5|et qui tangit reptile, quo polluitur, vel hominem, quo polluitur qualibet immunditia illius,
LEV|22|6|immundus erit usque ad vesperum et non vescetur his, quae sanctificata sunt; sed cum laverit carnem suam aqua,
LEV|22|7|et occubuerit sol, tunc mundatus vescetur de sanctificatis, quia cibus illius est.
LEV|22|8|Morticinum et dilaceratum a bestia non comedent, nec polluentur in eis. Ego Dominus.
LEV|22|9|Custodient praeceptum meum, ut non habeant super illo peccatum et propterea moriantur, cum polluerint illud; ego Dominus, qui sanctifico eos.
LEV|22|10|Omnis alienigena non comedet de sanctificatis, inquilinus sacerdotis et mercennarius non vescentur ex eis.
LEV|22|11|Quem autem sacerdos emerit, et qui vernaculus domus eius fuerit, hi comedent ex eis.
LEV|22|12|Si filia sacerdotis cuilibet ex populo nupta fuerit, de muneribus, quae sanctificata sunt, non vescetur;
LEV|22|13|sin autem vidua vel repudiata et absque liberis reversa fuerit ad domum patris sui, sicut puella consueverat, aletur cibo patris sui. Omnis alienigena comedendi ex eo non habet potestatem.
LEV|22|14|Qui comederit de sanctificatis per ignorantiam, addet quintam partem cum eo, quod comedit, et dabit sacerdoti sanctificatum.
LEV|22|15|Nec contaminabunt sanctificata filiorum Israel, quae tamquam munus offerunt Domino,
LEV|22|16|ne inducant super eos iniquitatem delicti, cum illi sanctificata sua comederint. Ego Dominus, qui sanctifico ".
LEV|22|17|Locutus est Dominus ad Moysen dicens:
LEV|22|18|" Loquere ad Aaron et filios eius et ad omnes filios Israel dicesque ad eos: Homo de domo Israel et de advenis, qui habitant apud vos, qui obtulerit oblationem suam vel vota solvens vel sponte offerens, quidquid illud obtulerit in holocaustum Domino,
LEV|22|19|in beneplacitum pro vobis offeratur masculus immaculatus ex bobus et ex ovibus et ex capris;
LEV|22|20|si maculam habuerit, non offeretis, quia non erit vobis acceptabile.
LEV|22|21|Homo, qui obtulerit victimam pacificorum Domino, vel vota solvens vel sponte offerens tam de bobus quam de ovibus immaculatum offeret, ut acceptabile sit; omnis macula non erit in eo.
LEV|22|22|Si caecum fuerit, si fractum, si mutilum, si verrucam habens aut scabiem vel impetiginem, non offeretis ea Domino nec in incensum dabitis ex eis super altare Domino.
LEV|22|23|Bovem et ovem deformem et debilem voluntarie offerre potes; votum autem ex his solvi non potest.
LEV|22|24|Omne animal, quod vel contritis vel tusis vel sectis ablatisque testiculis est, non offeretis Domino, et in terra vestra hoc omnino ne faciatis.
LEV|22|25|De manu alienigenae non offeretis cibum Dei vestri ex omnibus his animalibus, quia corrupta et maculata sunt omnia; non erunt in beneplacitum pro vobis ".
LEV|22|26|Locutusque est Dominus ad Moysen dicens:
LEV|22|27|" Bos, ovis et capra, cum genita fuerint, septem diebus erunt sub ubere matris suae; die autem octavo et deinceps erunt acceptabile munus incensi Domino.
LEV|22|28|Sive illa bos sive ovis non immolabuntur una die cum fetibus suis.
LEV|22|29|Si sacrificaveritis hostiam pro gratiarum actione Domino, sacrificabitis, ut possit esse placabilis.
LEV|22|30|Eodem die comedetis eam; non remanebit quidquam in mane alterius diei. Ego Dominus.
LEV|22|31|Custodite mandata mea et facite ea. Ego Dominus.
LEV|22|32|Ne polluatis nomen meum sanctum, ut sanctificer in medio filiorum Israel. Ego Dominus, qui sanctifico vos
LEV|22|33|et eduxi de terra Aegypti, ut essem vobis in Deum. Ego Dominus ".
LEV|23|1|Locutus est Dominus ad Moysen dicens:
LEV|23|2|" Loquere filiis Israel et dices ad eos: Hae sunt feriae Domini, quas vocabitis conventus sanctos; hae sunt feriae meae.
LEV|23|3|Sex diebus facietis opus; dies septimus sabbatum requiei est, conventus sanctus; omne opus non facietis; sabbatum est Domino in cunctis habitationibus vestris.
LEV|23|4|Hae sunt ergo feriae Domini, conventus sancti, quas celebrare debetis temporibus suis.
LEV|23|5|Mense primo, quarta decima die mensis, ad vesperum Pascha Domini est.
LEV|23|6|Et quinta decima die mensis huius sollemnitas Azymorum Domini est. Septem diebus azyma comedetis.
LEV|23|7|Die primo erit vobis conventus sanctus; omne opus servile non facietis in eo,
LEV|23|8|sed offeretis incensum Domino septem diebus. Die autem septimo erit conventus sanctus, nullumque servile opus facietis in eo ".
LEV|23|9|Locutusque est Dominus ad Moysen dicens:
LEV|23|10|" Loquere filiis Israel et dices ad eos: Cum ingressi fueritis terram, quam ego dabo vobis, et messueritis segetem, feretis manipulum spicarum primitias messis vestrae ad sacerdotem,
LEV|23|11|qui elevabit fasciculum coram Domino, ut acceptabile sit pro vobis; altero die sabbati sanctificabit illum.
LEV|23|12|Atque in eodem die, quo manipulum consecrabitis, facietis agnum immaculatum anniculum in holocaustum Domino,
LEV|23|13|et oblationem cum eo duas decimas similae conspersae oleo in incensum Domino odoremque suavissimum et libamentum eius vini quartam partem hin.
LEV|23|14|Panem et grana tosta farrem recentem non comedetis ex segete usque ad diem, qua offeretis ex ea munus Deo vestro. Praeceptum est sempiternum generationibus vestris in cunctis habitaculis vestris.
LEV|23|15|Numerabitis vobis ab altero die sabbati, in quo obtulistis manipulum elationis, septem hebdomadas plenas
LEV|23|16|usque ad alteram diem expletionis hebdomadae septimae, id est quinquaginta dies; et sic offeretis oblationem novam Domino
LEV|23|17|ex habitaculis vestris panes elationis duos de duabus decimis similae fermentatae, quos coquetis in primitias Domino;
LEV|23|18|offeretisque cum panibus septem agnos immaculatos anniculos et vitulum de armento unum et arietes duos, et erunt holocaustum Domino cum oblatione similae et libamentis suis in odorem suavissimum Domino.
LEV|23|19|Facietis et hircum in sacrificium pro peccato duosque agnos anniculos, hostias pacificorum.
LEV|23|20|Cumque elevaverit eos sacerdos cum panibus primitiarum coram Domino, cum duobus agnis sanctum erunt Domino in usum sacerdotis.
LEV|23|21|Et vocabitis hoc ipso die conventum, conventus sanctus erit vobis; omne opus servile non facietis in eo. Legitimum sempiternum erit in cunctis habitaculis generationibus vestris.
LEV|23|22|Cum autem metatis segetem terrae vestrae, non secabis eam usque ad oram agri nec remanentes spicas colliges, sed pauperibus et peregrinis dimittes eas. Ego Dominus Deus vester ".
LEV|23|23|Locutusque est Dominus ad Moysen dicens:
LEV|23|24|" Loquere filiis Israel: Mense septimo, prima die mensis, erit vobis requies, memoriale, clangentibus tubis, conventus sanctus.
LEV|23|25|Omne opus servile non facietis in eo et offeretis incensum Domino ".
LEV|23|26|Locutusque est Dominus ad Moysen dicens:
LEV|23|27|" Attamen decimo die mensis huius septimi dies Expiationum est, conventus sanctus erit vobis; affligetisque animas vestras in eo et offeretis incensum Domino.
LEV|23|28|Omne opus non facietis in tempore diei huius, quia dies expiationum est in expiationem vestram coram Domino Deo vestro.
LEV|23|29|Omnis anima, quae afflicta non fuerit die hoc, peribit de populis suis;
LEV|23|30|et,quae operis quippiam fecerit die hac, delebo eam de populo suo.
LEV|23|31|Nihil ergo operis facietis in eo: legitimum sempiternum erit vestris generationibus in cunctis habitationibus vestris.
LEV|23|32|Sabbatum requietionis est vobis, et affligetis animas vestras; die nono mensis a vespero usque ad vesperum servabitis sabbatum vestrum ".
LEV|23|33|Et locutus est Dominus ad Moysen dicens:
LEV|23|34|" Loquere filiis Israel: Quinto decimo die mensis huius septimi erit festum Tabernaculorum septem diebus Domino.
LEV|23|35|Die primo conventus sanctus, omne opus servile non facietis in eo;
LEV|23|36|septem diebus offeretis incensum Domino. Die octavo conventus sanctus erit vobis et offeretis incensum Domino; est enim coetus: omne opus servile non facietis.
LEV|23|37|Hae sunt feriae Domini, quas vocabitis conventus sanctos, offeretisque in eis incensum Domino, holocausta et oblationes similae, sacrificia et libamenta iuxta ritum uniuscuiusque diei;
LEV|23|38|praeter sabbata Domini donaque vestra et omnia, quae offeretis ex voto vel quae sponte tribuetis Domino.
LEV|23|39|Sed quinto decimo die mensis septimi, quando congregaveritis omnes fructus terrae, celebrabitis festum Domini septem diebus; die primo et die octavo erit requies.
LEV|23|40|Sumetisque vobis die primo fructus arboris pulcherrimos spatulasque palmarum et ramos ligni densarum frondium et salices de torrente et laetabimini coram Domino Deo vestro.
LEV|23|41|Celebrabitisque sollemnitatem eius septem diebus per annum: legitimum sempiternum erit generationibus vestris. Mense septimo festum celebrabitis
LEV|23|42|et habitabitis in umbraculis septem diebus; omnis, qui de genere est Israel, manebit in tabernaculis,
LEV|23|43|ut discant posteri vestri quod in tabernaculis habitare fecerim filios Israel, cum educerem eos de terra Aegypti. Ego Dominus Deus vester ".
LEV|23|44|Locutusque est Moyses super sollemnitatibus Domini ad filios Israel.
LEV|24|1|Et locutus est Dominus ad Moysen dicens:
LEV|24|2|" Praecipe fi liis Israel, ut afferant tibi oleum de olivis purissimum ac lucidum ad concinnandas lucernas candelabri iugiter.
LEV|24|3|Extra velum testimonii in tabernaculo conventus parabit illud Aaron a vespere usque ad mane coram Domino iugiter, ritu perpetuo in generationibus vestris.
LEV|24|4|Super candelabro mundissimo parabit lucernas semper in conspectu Domini.
LEV|24|5|Accipies quoque similam et coques ex ea duodecim panes, qui singuli habebunt duas decimas,
LEV|24|6|quorum senos altrinsecus super mensam purissimam coram Domino statues.
LEV|24|7|Et pones super ambas strues tus lucidissimum, ut sit panis in memoriale, incensum Domino.
LEV|24|8|Per singula sabbata mutabuntur coram Domino suscepti a filiis Israel; foedus sempiternum.
LEV|24|9|Eruntque Aaron et filiorum eius, ut comedant eos in loco sancto, quia sanctum sanctorum est ei de incensis Domini; iure perpetuo ".
LEV|24|10|Ecce autem egressus filius mulieris Israelitis, quem pepererat de viro Aegyptio inter filios Israel, iurgatus est in castris cum viro Israelita.
LEV|24|11|Cumque blasphemasset nomen et maledixisset ei, adductus est ad Moysen; vocabatur autem mater eius Salomith filia Dabri de tribu Dan.
LEV|24|12|Miseruntque eum in custodiam, donec nossent quid iuberet Dominus.
LEV|24|13|Qui locutus est ad Moysen dicens:
LEV|24|14|" Educ blasphemum extra castra, et ponant omnes, qui audierunt, manus suas super caput eius, et lapidet eum coetus universus.
LEV|24|15|Et ad filios Israel loqueris:Homo, qui maledixerit Deo suo, portabit peccatum suum;
LEV|24|16|et, qui blasphemaverit nomen Domini, morte moriatur: lapidibus opprimet eum omnis coetus, sive ille peregrinus sive civis fuerit. Qui blasphemaverit nomen Domini, morte moriatur.
LEV|24|17|Qui percusserit et occiderit hominem, morte moriatur.
LEV|24|18|Qui percusserit animal, reddet vicarium, id est animam pro anima.
LEV|24|19|Qui irrogaverit maculam cuilibet civium suorum, sicut fecit, sic fiet ei:
LEV|24|20|fracturam pro fractura, oculum pro oculo, dentem pro dente restituet; qualem inflixerit maculam, talem sustinere cogetur.
LEV|24|21|Qui percusserit iumentum, reddet aliud. Qui percusserit hominem, morietur.
LEV|24|22|Aequum iudicium sit inter vos, sive peregrinus sive civis peccaverit; quia ego sum Dominus Deus vester ".
LEV|24|23|Locutusque est Moyses ad filios Israel, et eduxerunt eum, qui blasphemaverat, extra castra, ac lapidibus oppresserunt. Feceruntque filii Israel, sicut praeceperat Dominus Moysi.
LEV|25|1|Locutusque est Dominus ad Moysen in monte Sinai di cens:
LEV|25|2|" Loquere filiis Israel et dices ad eos: Quando ingressi fueritis terram, quam ego dabo vobis, sabbatizet terra sabbatum Domino.
LEV|25|3|Sex annis seres agrum tuum et sex annis putabis vineam tuam colligesque fructus eius;
LEV|25|4|septimo autem anno, sabbatum requietionis erit terrae, sabbatum Domino: agrum tuum non seres et vineam tuam non putabis.
LEV|25|5|Quae sponte gignit humus, non metes et uvas vineae tuae non putatae non colliges quasi vindemiam; annus enim requietionis erit terrae.
LEV|25|6|Et erit sabbatum terrae vobis in cibum: tibi et servo tuo, ancillae et mercennario tuo et advenis, qui peregrinantur apud te,
LEV|25|7|iumentis tuis et animalibus, quae in terra tua sunt, omnia, quae nascuntur, praebebunt cibum.
LEV|25|8|Numerabis quoque tibi septem hebdomadas annorum, id est septem septies, quae simul faciunt annos quadraginta novem;
LEV|25|9|et clanges bucina mense septimo, decima die mensis expiationis die clangetis tuba in universa terra vestra.
LEV|25|10|Sanctificabitisque annum quinquagesimum et vocabitis remissionem in terra cunctis habitatoribus eius: ipse est enim iobeleus. Revertemini unusquisque ad possessionem suam, et unusquisque rediet ad familiam pristinam.
LEV|25|11|Iobeleus erit vobis quinquagesimus annus. Non seretis neque metetis sponte in agro nascentia neque vineas non putatas vindemiabitis
LEV|25|12|ob sanctificationem iobelei; sed de agro statim ablatas comedetis fruges.
LEV|25|13|Hoc anno iobelei rediet unusquisque vestrum ad possessionem suam.
LEV|25|14|Quando vendes quippiam civi tuo vel emes ab eo, ne contristet unusquisque fratrem suum; sed iuxta numerum annorum post iobeleum emes ab eo,
LEV|25|15|et iuxta supputationem annorum frugum vendet tibi.
LEV|25|16|Quanto plures anni remanserint post iobeleum, tanto crescet et pretium; et quanto minus temporis numeraveris, tanto minoris et emptio constabit: tempus enim frugum vendet tibi.
LEV|25|17|Nolite affligere contribules vestros, sed timeas Deum tuum, quia ego Dominus Deus vester.
LEV|25|18|Facite praecepta mea et iudicia, custodite et implete ea, ut habitare possitis in terra absque ullo pavore,
LEV|25|19|et gignat vobis humus fructus suos, quibus vescamini usque ad saturitatem, et habitabitis super terram, nullius impetum formidantes.
LEV|25|20|Quod si dixeritis: "Quid comedemus anno septimo, si non seruerimus neque collegerimus fruges nostras?".
LEV|25|21|Dabo benedictionem meam vobis anno sexto, et faciet fructus trium annorum,
LEV|25|22|seretisque anno octavo et comedetis veteres fruges usque ad nonum annum; donec nova nascantur, edetis vetera.
LEV|25|23|Terra quoque non veniet in perpetuum, quia mea est, et vos advenae et coloni mei estis.
LEV|25|24|Unde cuncta regio possessionis vestrae sub redemptionis condicione a vobis vendetur.
LEV|25|25|Si attenuatus frater tuus vendiderit partem possessionis suae, veniet ut redemptor propinquus eius, et redimet, quod ille vendiderat.
LEV|25|26|Sin autem non habuerit redemptorem et ipse pretium ad redimendum potuerit invenire,
LEV|25|27|computabuntur fructus ex eo tempore, quo vendidit; et, quod reliquum est, reddet emptori sicque recipiet possessionem suam.
LEV|25|28|Quod si non invenerit manus eius, ut reddat pretium, habebit emptor, quod emerat, usque ad annum iobeleum. In ipso enim omnis venditio rediet ad dominum et ad possessorem pristinum.
LEV|25|29|Qui vendiderit domum intra urbis muros, habebit licentiam redimendi, donec unus impleatur annus.
LEV|25|30|Si non redemerit, et anni circulus fuerit evolutus, emptor possidebit eam et posteri eius in perpetuum; et redimi non poterit, etiam in iobeleo.
LEV|25|31|Sin autem in villa fuerit domus, quae muros non habet, agrorum iure vendetur: potest redimi et in iobeleo revertetur ad dominum.
LEV|25|32|Aedes Levitarum, quae in urbibus possessionis eorum sunt, semper possunt ab eis redimi.
LEV|25|33|Si autem quis redemerit a Levitis, domus et urbs in iobeleo revertentur ad dominos; quia domus urbium leviticarum pro possessionibus eorum sunt inter filios Israel.
LEV|25|34|Suburbana autem pascua eorum non venient, quia possessio sempiterna est eis.
LEV|25|35|Si attenuatus fuerit frater tuus, et infirma manus eius apud te, suscipies eum quasi advenam et peregrinum, et vivet tecum.
LEV|25|36|Ne accipias usuras ab eo nec amplius quam dedisti: time Deum tuum, ut vivere possit frater tuus apud te.
LEV|25|37|Pecuniam tuam non dabis ei ad usuram nec plus aequo exiges pro cibo tuo.
LEV|25|38|Ego Dominus Deus vester, qui eduxi vos de terra Aegypti, ut darem vobis terram Chanaan et essem vester Deus.
LEV|25|39|Si paupertate compulsus vendiderit se tibi frater tuus, non eum opprimes servitute servorum,
LEV|25|40|sed quasi mercennarius et colonus erit tecum. Usque ad annum iobeleum operabitur apud te
LEV|25|41|et postea egredietur cum liberis suis et revertetur ad cognationem suam et ad possessionem patrum suorum.
LEV|25|42|Mei enim servi sunt, et ego eduxi eos de terra Aegypti: non venient condicione servorum;
LEV|25|43|ne affligas eum per po tentiam, sed metuito Deum tuum.
LEV|25|44|Servus et ancilla sint tibi de nationibus, quae in circuitu vestro sunt; de illis emetis servum et ancillam.
LEV|25|45|De filiis quoque advenarum, qui peregrinantur apud vos, emetis et de cognatione eorum, quae est apud vos et quam genuerint in terra vestra, hos habebitis in possessionem
LEV|25|46|et hereditario iure transmittetis ad posteros ac possidebitis in aeternum ut servos; fratres autem vestros filios Israel ne opprimatis cum potentia.
LEV|25|47|Si invaluerit apud vos manus advenae atque peregrini, et attenuatus frater tuus vendiderit se ei aut cuiquam de stirpe eius,
LEV|25|48|post venditionem potest redimi. Unus ex fratribus suis redimet eum
LEV|25|49|et patruus et patruelis et consanguineus et affinis. Sin autem et ipse potuerit, redimat se,
LEV|25|50|supputatis dumtaxat cum emptore annis a tempore venditionis suae usque ad annum iobeleum, et pecunia, qua venditus fuerat, iuxta annorum numerum et rationem mercennarii supputata.
LEV|25|51|Si plures fuerint anni, qui remanent usque ad iobeleum, secundum hos reddet et pretium redemptionis de pecunia emptionis;
LEV|25|52|si pauci, ponet rationem cum eo; iuxta annorum numerum reddet emptori, quod reliquum est annorum,
LEV|25|53|quibus ante servivit, mercedibus mercennarii imputatis. Non affliget eum violenter in conspectu tuo.
LEV|25|54|Quod si per haec redimi non potuerit, anno iobeleo egredietur cum liberis suis:
LEV|25|55|mei sunt enim servi filii Israel, quos eduxi de terra Aegypti. Ego Dominus Deus vester ".
LEV|26|1|" Non facietis vobis idolum et sculptile nec lapidem eri getis nec imaginem sculptam in petra ponetis in terra vestra, ut adoretis eam. Ego enim sum Dominus Deus vester.
LEV|26|2|Custodite sabbata mea et pavete sanctuarium meum. Ego Dominus.
LEV|26|3|Si in praeceptis meis ambulaveritis et mandata mea custodieritis et feceritis ea,
LEV|26|4|dabo vobis pluvias temporibus suis, et terra gignet germen suum, et pomis arbores replebuntur.
LEV|26|5|Apprehendet messium tritura vindemiam, et vindemia occupabit sementem; et comedetis panem vestrum in saturitatem et absque pavore habitabitis in terra vestra.
LEV|26|6|Dabo pacem in finibus vestris, dormietis, et non erit qui exterreat. Auferam malas bestias, et gladius non transibit per terminos vestros.
LEV|26|7|Persequemini inimicos vestros, et corruent coram vobis gladio.
LEV|26|8|Persequentur quinque de vestris centum alienos, et centum ex vobis decem milia; cadent inimici vestri in conspectu vestro gladio.
LEV|26|9|Respiciam vos et crescere faciam; multiplicabimini, et firmabo pactum meum vobiscum.
LEV|26|10|Comedetis vetusta congregata priorum messium; et vetera, novis supervenientibus, proicietis.
LEV|26|11|Ponam habitaculum meum in medio vestri, et non abominabitur vos anima mea.
LEV|26|12|Ambulabo inter vos et ero vester Deus, vosque eritis populus meus.
LEV|26|13|Ego Dominus Deus vester, qui eduxi vos de terra Aegyptiorum, ne serviretis eis, et qui confregi vectes iugi vestri, ut incederetis erecti.
LEV|26|14|Quod si non audieritis me nec feceritis omnia mandata haec,
LEV|26|15|si spreveritis leges meas, et iudicia mea contempserit anima vestra, ut non faciatis omnia, quae a me constituta sunt, et ad irritum perducatis pactum meum,
LEV|26|16|ego quoque haec faciam vobis: visitabo vos in terrore repentino, in tabe et ardore, qui conficiant oculos et consumant animam, frustra seretis sementem, quae ab hostibus devorabitur.
LEV|26|17|Ponam faciem meam contra vos, et corruetis coram hostibus vestris et subiciemini his, qui oderunt vos, et fugietis, nemine persequente.
LEV|26|18|Sin autem nec sic oboedieritis mihi, addam correptiones vestras septuplum propter peccata vestra
LEV|26|19|et conteram superbiam duritiae vestrae. Daboque caelum vobis desuper sicut ferrum et terram aeneam.
LEV|26|20|Consumetur incassum robur vestrum: non proferet terra germen, nec arbores poma praebebunt.
LEV|26|21|Si ambulaveritis ex adverso mihi nec volueritis audire me, addam plagas vestras usque in septuplum propter peccata vestra;
LEV|26|22|emittamque in vos bestias agri, quae absque liberis vos faciant et deleant pecora vestra et ad paucitatem vos redigant, desertaeque fiant viae vestrae.
LEV|26|23|Quod si nec sic volueritis recipere disciplinam, sed ambulaveritis ex adverso mihi,
LEV|26|24|ego quoque contra vos adversus incedam et percutiam vos septies propter peccata vestra.
LEV|26|25|inducamque super vos gladium ultorem foederis mei; cumque confugeritis in urbes vestras, mittam pestilentiam in medio vestri, et trademini hostium manibus.
LEV|26|26|Postquam confregero vobis baculum panis, coquent decem mulieres in uno clibano panem vestrum et reddent eum ad pondus, et comedetis et non saturabimini.
LEV|26|27|Sin autem nec per haec audieritis me, sed ambulaveritis contra me,
LEV|26|28|et ego incedam adversus vos in furore contrario; et corripiam vos septem plagis propter peccata vestra,
LEV|26|29|ita ut comedatis carnes filiorum et filiarum vestrarum.
LEV|26|30|Destruam excelsa vestra et thymiamateria confringam et ponam cadavera vestra super cadavera idolorum vestrorum, et abominabitur vos anima mea,
LEV|26|31|in tantum ut urbes vestras redigam in solitudinem et deserta faciam sanctuaria vestra nec recipiam ultra odorem suavissimum.
LEV|26|32|Disperdamque terram vestram; et stupebunt super ea inimici vestri, cum habitatores illius fuerint.
LEV|26|33|Vos autem dispergam in gentes et evaginabo post vos gladium; eritque terra vestra deserta et civitates dirutae.
LEV|26|34|Tunc placebunt terrae sabbata sua cunctis diebus solitudinis suae; quando fueritis in terra hostili, sabbatizabit et sabbata sua supplebit.
LEV|26|35|Cunctis diebus solitudinis sabbatizabit, eo quod non requieverit in sabbatis vestris, quando habitabatis in ea.
LEV|26|36|Et, qui de vobis remanserint, dabo pavorem in cordibus eorum in regionibus hostium; terrebit eos sonitus folii volantis, et ita fugient quasi gladium; cadent, nullo persequente.
LEV|26|37|Et corruent singuli super fratres suos quasi bella fugientes, nemine persequente. Nemo vestrum inimicis audebit resistere.
LEV|26|38|Peribitis inter gentes, et hostilis vos terra consumet.
LEV|26|39|Quod si et de vobis aliqui remanserint, tabescent in iniquitatibus suis in terris inimicorum vestrorum et propter peccata patrum suorum cum ipsis tabescent.
LEV|26|40|Et confitebuntur iniquitates suas et maiorum suorum, quibus praevaricati sunt in me et ambulaverunt ex adverso mihi,
LEV|26|41|ut et ego ambularem contra eos et inducerem illos in terram hostilem; vel tunc humiliabitur incircumcisum cor eorum, et tunc expiabunt pro impietatibus suis.
LEV|26|42|Et recordabor foederis mei, quod pepigi cum Iacob et Isaac et Abraham. Terrae quoque memor ero,
LEV|26|43|quae, cum relicta fuerit ab eis, complacebit sibi in sabbatis suis patiens solitudinem propter illos. Ipsi vero expiabunt pro peccatis suis, eo quod abiecerint iudicia mea et leges meas despexerint.
LEV|26|44|Et tamen, etiam cum essent in terra hostili, non penitus abieci eos neque sic despexi, ut consumerentur, et irritum facerem pactum meum cum eis. Ego enim sum Dominus, Deus eorum.
LEV|26|45|Et recordabor eis foederis cum maioribus, quos eduxi de terra Aegypti in conspectu gentium, ut essem Deus eorum. Ego Dominus ".
LEV|26|46|Haec sunt iudicia atque praecepta et leges, quas dedit Dominus inter se et inter filios Israel in monte Sinai per manum Moysi.
LEV|27|1|Locutusque est Dominus ad Moysen dicens:
LEV|27|2|" Loquere fi liis Israel et dices ad eos: Homo, qui votum fecerit et spoponderit Deo animas, sub aestimatione dabit pretium:
LEV|27|3|si fuerit masculus a vicesimo usque ad sexagesimum annum, dabit quinquaginta siclos argenti ad mensuram sanctuarii;
LEV|27|4|si mulier, triginta.
LEV|27|5|A quinto autem anno usque ad vicesimum masculus dabit viginti siclos, femina decem;
LEV|27|6|ab uno mense usque ad annum quintum pro masculo dabuntur quinque sicli, pro femina tres;
LEV|27|7|sexagenarius et ultra masculus dabit quindecim siclos, femina decem.
LEV|27|8|Si pauper fuerit et aestimationem reddere non valebit, sistet eum coram sacerdote, et quantum ille aestimaverit et viderit posse reddere, tantum dabit.
LEV|27|9|Animal autem, quod immolari potest Domino, si quis voverit, sanctum erit
LEV|27|10|et mutari non poterit, id est nec melius malo nec peius bono. Quod si mutaverit, et ipsum quod mutatum est et illud pro quo mutatum est, consecratum erit Domino.
LEV|27|11|Animal immundum, quod immolari Domino non potest, si quis voverit, adducetur ante sacerdotem,
LEV|27|12|qui diiudicans utrum bonum an malum sit, sicut statuet pretium, sic erit.
LEV|27|13|Quod si redimere illud voluerit is qui offert, addet supra aestimationem quintam partem.
LEV|27|14|Homo si voverit domum suam et sanctificaverit Domino, considerabit eam sacerdos utrum bona an mala sit, et iuxta pretium, quod ab eo fuerit constitutum, stabit.
LEV|27|15|Sin autem ille, qui voverat, voluerit redimere eam, dabit quintam partem aestimationis supra et habebit domum.
LEV|27|16|Quod si agrum possessionis suae voverit et consecraverit Domino, iuxta mensuram sementis aestimabitur pretium: si triginta homer hordei seritur terra, quinquaginta siclis aestimabitur argenti.
LEV|27|17|Si statim ab anno iobelei voverit agrum, quanto valere potest, tanto aestimabitur.
LEV|27|18|Sin autem post aliquantum temporis, supputabit ei sacerdos pecuniam iuxta annorum, qui reliqui sunt, numerum usque ad iobeleum, et detrahetur ex pretio.
LEV|27|19|Quod si voluerit redimere agrum ille, qui voverat, addet quintam partem aestimatae pecuniae et possidebit eum.
LEV|27|20|Sin autem noluerit redimere, sed alteri cuilibet vendiderit, ultra redimi non poterit;
LEV|27|21|sed, cum iobelei venerit dies, sanctum erit Domino sicut ager anathematis; sacerdotis erit possessio eius.
LEV|27|22|Quod si agrum emptum, qui non est de possessione maiorum, sanctificare voluerit Domino,
LEV|27|23|supputabit ei sacerdos iuxta annorum numerum usque ad iobeleum pretium, quod dabit ille, qui voverat, in ipso die ut sanctum Domino.
LEV|27|24|In anno autem iobelei revertetur ager ad priorem dominum, qui vendiderat eum et habuerat in sortem possessionis suae.
LEV|27|25|Omnis aestimatio siclo sanctuarii ponderabitur; siclus viginti gera habet.
LEV|27|26|Primogenita, quae de animalibus ad Dominum pertinent, nemo sanctificare poterit et vovere: sive bos sive ovis fuerit, Domini sunt.
LEV|27|27|Quod si immundum est animal, redimet, qui obtulit, iuxta aestimationem et addet quintam partem pretii; si redimere noluerit, vendetur quanto fuerit.
LEV|27|28|Omne anathema, quod aliquis vir consecrat Domino de omni possessione sua, sive homo fuerit sive animal sive ager, non veniet nec redimi poterit; quidquid semel fuerit consecratum, sanctum sanctorum erit Domino.
LEV|27|29|Et omnis homo, qui ut anathema offertur, non redimetur, sed morte morietur.
LEV|27|30|Omnes decimae terrae sive de frugibus sive de pomis arborum Domini sunt, sanctum Domino.
LEV|27|31|Si quis autem voluerit redimere aliquid de decimis suis, addet quintam partem.
LEV|27|32|Omnes decimae boves et oves et caprae, quae sub pastoris virga transeunt, quidquid decimum venerit, erit sanctum Domino.
LEV|27|33|Non discernetur inter bonum et malum nec altero commutabitur; si quis mutaverit, et quod mutatum est et pro quo mutatum est, sanctum erit et non redimetur ".
LEV|27|34|Haec sunt praecepta, quae mandavit Dominus Moysi ad filios Israel in monte Sinai.
