MIC|1|1|Слово Господнє, що було до морешетського Михея за днів Йотама, Ахаза та Єзекії, Юдиних царів, яке він бачив на Самарію та Єрусалим.
MIC|1|2|Почуйте оце, всі народи, послухай, ти земле та все, що на ній! і хай буде за свідка на вас Господь Бог, Господь з храму святого Свого!
MIC|1|3|Бо Господь ось виходить із місця Свого, і Він сходить і ступає по висотах землі.
MIC|1|4|І топляться гори під Ним, і тануть долини, мов віск від огню, мов ті води, що ллються з узбіччя.
MIC|1|5|Усе це за провинення Якова, за гріхи дому Ізраїля. Хто провинення Якова, чи ж не Самарія? А хто гріх дому Юдиного, чи ж не Єрусалим?
MIC|1|6|І зроблю Самарію руїною в полі, за місце садити виноград, і повикидаю в долину каміння її, і відкрию основи її.
MIC|1|7|І потовчені будуть усі її ідоли, всі ж дарунки її за розпусту попалені будуть в огні, і всіх бовванів її Я віддам на спустошення. Бо зібрала вона від дарунків за блуд, і на подарунки за блуд це повернеться.
MIC|1|8|Над оцим голоситиму я та ридатиму, ходитиму босий й нагий, заводити буду, немов ті шакали, і буду тужити, як струсі!
MIC|1|9|Бо рани її невигойні, бо це аж до Юди прийшло, воно досягло аж до брами народу Мого, аж до Єрусалиму.
MIC|1|10|Цього не оголошуйте в Ґаті, і плакати не плачте, качайтесь по поросі в Бет-Леафрі.
MIC|1|11|Переходь собі ти, о мешканко Шафіру, нага, осоромлена, вже бо не вийде мешканка Цаанану, голосіння Бет-Гаецелу не дасть вам спинитися в ньому.
MIC|1|12|Бо мешканка Мароту чекала добра, та до єрусалимської брами зійшло оце лихо від Господа.
MIC|1|13|Запряжи баскі коні до воза, мешканко Лахішу! Ти початок гріха для сіонської доньки, бо знайшлись серед тебе провини Ізраїлеві,
MIC|1|14|тому то даси розводові листи на Морешет-Ґат. Доми Ахзіва омана для Ізраїлевих царів.
MIC|1|15|Спроваджу тобі ще спадкоємця Я, о мешканко Мареші, Аж по Адуллам прийде слава Ізраїля.
MIC|1|16|Зроби собі лисину та острижися за синів своїх любих, пошир свою лисину, мов ув орла, бо пішли на вигнання від тебе вони!
MIC|2|1|Горе тим, що задумують кривду і на ложах своїх учиняють лихе! За світла поранку виконують це, бо їхня рука має силу.
MIC|2|2|Якщо піль жадають, то грабують вони, а домів то хапають. І вони переслідують мужа та дома його, і чоловіка й спадки його.
MIC|2|3|Тому так промовляє Господь: Ось Я замишляю на цей рід лихе, що ший своїх з нього не визволите, і ходити не будете гордо, бо це час лихий.
MIC|2|4|Того дня проголосять на вас приповістку, і співатимуть пісню жалобну, говорячи: Сталось! До пня опустошені ми, уділ народу мого змінився, як це діткнуло мене! Наше поле поділене буде чужинцями,
MIC|2|5|тому в тебе не буде нікого, хто кидав би шнура мірничого, як жеребка на Господнім зібранні.
MIC|2|6|Не проповідуйте, та вони проповідують! Хай нам не проповідують, не досягне нас ганьба.
MIC|2|7|О ти, що звешся Яковів дім, чи змалів Дух Господній? Чи ці чини Його? Хіба добре не роблять слова Мої тому, хто ходить правдиво?
MIC|2|8|Ще вчора були ви народом Моїм, тепер же стаєте за ворога, з одежі верхньої плаща ви стягаєте з тих, хто проходить безпечно, як здобич війни.
MIC|2|9|Жінок Мого народу з приємного дому її виганяєте кожну, з дітей славу Мою ви берете навіки.
MIC|2|10|Устаньте й ідіть, бо тут не спочинок, це за занечищення ваше, що загладу для вас принесе, вирішальну загладу.
MIC|2|11|Коли б чоловік, який ходить за вітром, і брехню набрехав, говорячи: Буду тобі проповідувати про вино та про напій п'янкий, то був би він любим пророком оцьому народові.
MIC|2|12|Невідмінно зберу тебе всього, о Якове, невідмінно згромаджу останок Ізраїлів, разом поставлю його, як отару в Боцрі, як ту череду на пасовищі, і будуть гомоніти вони від многолюдства!
MIC|2|13|Перед ними виламувач піде, вони продеруться та браму перейдуть і вийдуть із неї. І піде їхній цар перед ними, а Господь на чолі їх!
MIC|3|1|А я відказав: Послухайте ж, голови Якова та начальники дому Ізраїля, чи ж не вам знати право?
MIC|3|2|Добро ви ненавидите та кохаєте зло, шкіру їхню здираєте з них, а їхнє тіло з костей їхніх.
MIC|3|3|Ви останок народу Мого їсте та стягаєте з них їхню шкіру, а їхні кості ламаєте, і січете, немов до горняти, і мов м'ясо в котел.
MIC|3|4|Вони тоді кликати будуть до Господа, та Він відповіді їм не дасть, і заховає обличчя Своє того часу від них, коли будуть робити лихі свої вчинки.
MIC|3|5|Так говорить Господь на пророків, що вводять народ Мій у блуд, що зубами своїми гризуть та покликують: Мир! А на того, хто їм не дає що до рота, на нього святую війну оголошують.
MIC|3|6|Тому буде вам ніч, щоб не стало видіння, і стемніє вам, щоб не чарувати. І над тими пророками сонце закотиться, і над ними потемніє день.
MIC|3|7|І посоромлені будуть такі прозорливці, і будуть застиджені чарівники, і всі вони свої уста закриють, бо не буде їм Божої відповіді.
MIC|3|8|А я повний сили й Господнього Духа, і правди й відваги, щоб представити Якову прогріх його, а Ізраїлеві його гріх.
MIC|3|9|Почуйте ж це, голови дому Якового та начальники дому Ізраїля, які нехтують справедливість, а все просте викривлюють,
MIC|3|10|вони кров'ю будують Сіона, а кривдою Єрусалима.
MIC|3|11|Його голови судять за хабара, і навчають за плату його ті священики, і за срібло ворожать пророки його, хоч на Господа вони опираються, кажучи: Хіба не Господь серед нас? Зло не прийде на нас!
MIC|3|12|О так, через вас Сіон буде на поле заораний, а Єрусалим на руїни обернеться, а гора храмова стане взгір'ями лісу...
MIC|4|1|Та буде наприкінці днів, гора дому Господнього міцно поставлена буде вершиною гір, і піднесена буде вона понад узгір'я, і будуть народи до неї пливсти.
MIC|4|2|І підуть численні народи та й скажуть: Ходімо, і вийдім на гору Господню та до дому Якового, і Він буде навчати доріг Своїх нас, і ми будемо ходити стежками Його. Бо вийде Закон із Сіону, а слово Господнє із Єрусалиму.
MIC|4|3|І Він буде судити численні племена, і розсуджувати буде народи міцні аж у далечині. І вони перекують мечі свої на лемеші, а списи свої на серпи. Не підійме меча народ на народ, і більше не будуть навчатись війни!
MIC|4|4|І буде кожен сидіти під своїм виноградником, і під своєю фіґовницею, і не буде того, хто б страшив, бо уста Господа Саваота оце прорекли.
MIC|4|5|Усі бо народи ходитимуть кожен ім'ям свого бога, а ми будем ходити Ім'ям Господа, нашого Бога, на віки віків!
MIC|4|6|Того дня промовляє Господь позбираю кульгаве й згромаджу розігнане, і те, що на нього навів коли лихо.
MIC|4|7|І зроблю Я кульгаве останком, а віддалене потужним народом, і зацарює над ними Господь на Сіонській горі відтепер й аж навіки!
MIC|4|8|А ти, башто Черідна, підгірку Сіонської доньки, прийде до тебе і дійде старе панування, царювання для донечки Єрусалиму.
MIC|4|9|Тепер нащо здіймаєш ти окрик? Чи в тебе немає царя? Чи ж загинув твій радник, що ти корчишся, мов породілля?
MIC|4|10|Вийся та корчся, о дочко Сіону, немов породілля, бо тепер вийдеш із міста та перебуватимеш у полі, і прийдеш аж до Вавилону. Та будеш ти там урятована, там Господь тебе викупить з рук твоїх ворогів!
MIC|4|11|А зараз зібрались на тебе численні народи, говорячи: Нехай він зневажений буде, і нехай наше око побачить нещастя Сіону!
MIC|4|12|Та не знають вони Господніх думок, і не розуміють поради Його, бо Він їх позбирав, як до клуні снопи.
MIC|4|13|Ставай та молоти, дочко Сіону, бо Я ріг твій залізом учиню, а копита твої вчиню міддю, і ти розпорошиш численні народи та вчиниш закляттям для Господа несправедливий їхній зиск, а їхнє багатство Владиці всієї землі.
MIC|5|1|(4-14) І згромаджуйсь тепер, дочко товпищ! Облогу вчинили на нас, тростиною б'ють по щоці Ізраїлевого суддю...
MIC|5|2|(5-1) А ти, Віфлеєме-Єфрате, хоч малий ти у тисячах Юди, із тебе Мені вийде Той, що буде Владика в Ізраїлі, і віддавна постання Його, від днів віковічних.
MIC|5|3|(5-2) Тому Він їх видасть до часу, аж поки ота не породить, що має родити, а останок братів Його вернеться до Ізраїлевих синів.
MIC|5|4|(5-3) І стане, і буде Він пасти Господньою силою, величністю Ймення Господа Бога Свого. І осядуть вони, бо Він стане великий тепер аж до кінців землі!
MIC|5|5|(5-4) І Він буде миром. Як прийде до нашого краю Ашшур, і буде топтатись по наших палатах, то поставимо на нього сім пастирів та восьмеро людських княжат.
MIC|5|6|(5-5) І вони будуть пасти мечем край Ашшура, край же Німрода у воротях його. Та Він від Ашшура врятує, як той прийде в наш Край, і коли буде топтатись по наших границях.
MIC|5|7|(5-6) І Яковів залишок буде посеред численних народів, як роса та від Господа, як той дощ на траві, і він надії не кластиме на чоловіка, і не буде надії складати на людських синів.
MIC|5|8|(5-7) І Яковів залишок буде між людами, серед численних народів, як лев між лісною худобою, як левчук між отарами овець, що як він переходить, то топче й шматує, і немає нікого, хто б зміг урятувати.
MIC|5|9|(5-8) Хай зведеться рука твоя на твоїх ненависників, і хай всі вороги твої витяті будуть!
MIC|5|10|(5-9) І станеться в день той, говорить Господь, і витну Я коні твої з-серед тебе, і колесниці твої повигублюю.
MIC|5|11|(5-10) І понищу міста твого Краю, і всі твердині твої порозвалюю.
MIC|5|12|(5-11) І повиполюю чари з твоєї руки, і ворожбитів у тебе не буде.
MIC|5|13|(5-12) І понищу боввани твої та жертовні стовпи твої з-посеред тебе, і ти чинові рук своїх більше не будеш вклонятися.
MIC|5|14|(5-13) І повитинаю дерева жертовні твої з-серед тебе, і міста твої вигублю.
MIC|5|15|(5-14) І в гніві та в лютості помсту вчиню над народами, що Мене не послухались!
MIC|6|1|Послухайте, що промовляє Господь: Устань, сперечайсь перед горами, і хай узгір'я почують твій голос!
MIC|6|2|Послухайте, гори, Господнього суду, і візьміть до вух, ви, основи землі, бо в Господа пря із народом Своїм, і з Ізраїлем буде судитися Він!
MIC|6|3|Народе ти Мій, що тобі Я зробив і чим мучив тебе, свідчи на Мене!
MIC|6|4|Бо Я з краю єгипетського тебе вивів, і тебе викупив з дому рабів, і перед тобою послав Я Мойсея, Аарона та Маріям.
MIC|6|5|Мій народе, згадай, що Балак, цар моавський, задумував був, і що йому відповів Валаам, син Беорів, від Шіттіму аж по Ґілґал, щоб пізнати тобі справедливості Господа.
MIC|6|6|З чим піду перед Господа, схилюсь перед Богом Високости? Чи піду перед Нього з цілопаленнями, з річними телятами?
MIC|6|7|Чи Господь уподобає тисячі баранів, десятитисячки потоків оливи? Чи дам за свій гріх свого первенця, плід утроби моєї за гріх моєї душі?
MIC|6|8|Було тобі виявлено, о людино, що добре, і чого пожадає від тебе Господь, нічого, а тільки чинити правосуддя, і милосердя любити, і з твоїм Богом ходити сумирно.
MIC|6|9|Голос Господній кличе до міста, а хто мудрий, боїться той Ймення Твого: Послухайте жезла й Того, Хто призначив його:
MIC|6|10|Чи є ще у домі безбожного коштовності несправедливі, та неповна й неправна ефа?
MIC|6|11|Чи Я всправедливлю вагу неправдиву, і калитку з важками обманними?
MIC|6|12|Що повні насильства його багачі, мешканці ж його говорили неправду, а їхній язик в їхніх устах омана,
MIC|6|13|то теж бити зачну Я тебе, пустошити тебе за гріхи твої.
MIC|6|14|Будеш ти їсти, але не наситишся, і буде голод у нутрі твоїм, і станеш ховати, але не врятуєш, а що ти врятуєш мечеві віддам.
MIC|6|15|Ти сіяти будеш, але не пожнеш, ти будеш оливку топтати, та не будеш маститись оливою, і молодий виноград, та вина ти не питимеш!
MIC|6|16|Бо ще переховуються всі устави Омрі та всі вчинки дому Ахава, і за їхніми радами ходите ви, тому то Я видам тебе на спустошення, і на посміх мешканців його, і ви ганьбу народу Мого понесете!
MIC|7|1|Горе мені, бо я став, мов недобірки літні, як залишки по винобранні; нема грона на їжу, немає доспілої фіґи, якої жадає душа моя!
MIC|7|2|Згинув побожний з землі, і нема поміж людьми правдивого. Вони всі чатують на кров, один одного ловлять у сітку.
MIC|7|3|Наставлені руки на зло, щоб вправно чинити його, начальник жадає дарунків, суддя ж судить за плату, а великий говорить жадання своєї душі, і викривлюють все.
MIC|7|4|Найліпший із них як будяк, найправдивіший гірший від терену. Настає день Твоїх сторожів, Твоїх відвідин, тепер буде збентеження їхнє!
MIC|7|5|І другові не довіряйте, не надійтесь на приятеля, від тієї, що при лоні твоєму лежить, пильнуй двері уст своїх!
MIC|7|6|Бо гордує син батьком своїм, дочка повстає проти неньки своєї, невістка проти свекрухи своєї, вороги чоловіку домашні його!
MIC|7|7|А я виглядаю на Господа, надіюсь на Бога спасіння мого, Бог мій почує мене!
MIC|7|8|Не тішся, моя супротивнице, з мене, хоч я впала, Сіонська дочка, проте встану, хоч сиджу в темноті, та Господь мені світло!
MIC|7|9|Буду зносити я гнів Господній, бо згрішила Йому, аж поки не вирішить справи моєї, та суду не вчинить мені. Він на світло мене попровадить, побачу Його справедливість!
MIC|7|10|І побачить оце все моя супротивниця, і сором покриє її, бо казала мені: Де Він, Господь, Бог твій? Приглядатимуться мої очі до неї, її топчуть тепер, як болото на вулицях.
MIC|7|11|Настане той день, щоб мури твої будувати, тоді віддалиться границя твоя цього дня!
MIC|7|12|Це той день, коли прийдуть до тебе з Асирії та аж до Єгипту, і від Єгипту та аж до Ріки, і від моря до моря, і від гори до гори.
MIC|7|13|І спустошенням стане земля на мешканців її, через плід їхніх учинків.
MIC|7|14|Паси Мій народ своїм берлом, отару спадку Твого; що пробуває в лісі самотно, у середині саду, хай пасуться вони на Башані й Ґілеаді, як за днів стародавніх.
MIC|7|15|Як за днів твого виходу з краю єгипетського, покажу йому чуда.
MIC|7|16|Народи побачать оце, і посоромлені будуть при всій своїй силі, руку покладуть на уста, їхні вуха оглухнуть.
MIC|7|17|Будуть порох лизати вони, як той гад, як плазюче землі, повилазять з дрижанням з укріплень своїх, вони будуть тремтіти перед Господом, Богом нашим, і будуть боятись Тебе!
MIC|7|18|Хто Бог інший, як Ти, що прощає провину і пробачує прогріх останку спадку Свого, Свого гніву не держить назавжди, бо кохається в милості?
MIC|7|19|Знов над нами Він змилується, наші провини потопче, Ти кинеш у морську глибочінь усі наші гріхи.
MIC|7|20|Ти даси правду Яковові, Авраамові милість, яку присягнув Він для наших батьків від днів стародавніх.
