DEUT|1|1|以下是 摩西 在 约旦河 东的旷野， 疏弗 对面的 亚拉巴 ，就是在 巴兰 、 陀弗 、 拉班 、 哈洗录 、 底撒哈 之间，向 以色列 众人所说的话。
DEUT|1|2|从 何烈山 经过 西珥山 到 加低斯．巴尼亚 要十一天的路程。
DEUT|1|3|第四十年十一月初一， 摩西 照耶和华所吩咐他一切有关 以色列 人的话，都告诉他们。
DEUT|1|4|那时，他已经击败了住 希实本 的 亚摩利 王 西宏 和住 亚斯她录 、 以得来 的 巴珊 王 噩 。
DEUT|1|5|摩西 在 约旦河 东的 摩押 地讲解这律法，说：
DEUT|1|6|“耶和华－我们的上帝在 何烈山 吩咐我们说：你们住在这山上已经够久了。
DEUT|1|7|要起行，转到 亚摩利 人的山区和附近的地区，就是 亚拉巴 、山区、 谢非拉 、 尼革夫 、沿海一带， 迦南 人的地和 黎巴嫩 ，直到 大河 ，就是 幼发拉底河 。
DEUT|1|8|看，我将这地摆在你们面前。你们要进去得这地，就是耶和华向你们列祖 亚伯拉罕 、 以撒 、 雅各 起誓要赐给他们和他们后裔为业之地。”
DEUT|1|9|“那时，我对你们说：‘我独自一人无法承担你们的事。
DEUT|1|10|耶和华－你们的上帝使你们增多。看哪，你们今日好像天上的星那样多。
DEUT|1|11|惟愿耶和华－你们列祖的上帝使你们更增加千倍，照他所应许你们的赐福给你们。
DEUT|1|12|但你们的担子，你们的重任，以及你们的争讼，我独自一人怎能承担呢？
DEUT|1|13|你们要按着各支派选出有智慧、明辨是非、为人所知的人来，我就立他们为你们的领袖。’
DEUT|1|14|你们回答我说：‘你说要做的事很好！’
DEUT|1|15|我就将你们各支派的领袖，就是有智慧、为人所知的人，立他们为领袖，作你们各支派的千夫长、百夫长、五十夫长、十夫长等官长，来管理你们。
DEUT|1|16|“当时，我吩咐你们的审判官说：‘你们听讼，无论是弟兄之间的诉讼，或与寄居者之间的诉讼，都要秉公判断。
DEUT|1|17|审判的时候不可看人的情面；无论大小，你们都要听讼。不可因人而惧怕，因为审判是上帝的事。你们当中若有难断的案件，可以呈到我这里，让我来听讼。’
DEUT|1|18|那时，我已经把你们所当做的事都吩咐你们了。”
DEUT|1|19|“我们照着耶和华－我们上帝所吩咐的，从 何烈山 起行，经过你们所看见那一切大而可怕的旷野，往 亚摩利 人的山区去，到了 加低斯．巴尼亚 。
DEUT|1|20|我对你们说：‘你们已经到了耶和华－我们上帝所赐给我们的 亚摩利 人之山区。
DEUT|1|21|看，耶和华－你的上帝已将那地摆在你面前，你要照耶和华－你列祖的上帝所说的，上去得那地为业。不要惧怕，也不要惊惶。’
DEUT|1|22|你们都来到我这里，说：‘让我们先派人去，为我们窥探那地，把我们上去该走的路线和该进的城镇回报我们。’
DEUT|1|23|这话我看为美，就从你们中间选取十二个人，每支派一人。
DEUT|1|24|于是他们起身上山区去，到 以实各谷 ，窥探那地。
DEUT|1|25|他们的手带着那地的一些果子，下到我们这里，回报我们说：‘耶和华－我们的上帝所赐给我们的是美地。’
DEUT|1|26|“你们却不肯上去，竟违背了耶和华─你们上帝的指示，
DEUT|1|27|在帐棚内发怨言说：‘耶和华因为恨我们，所以将我们从 埃及 地领出来，要把我们交在 亚摩利 人的手中，除灭我们。
DEUT|1|28|我们上哪里去呢？我们的弟兄使我们胆战心惊 ，说那里的百姓比我们又大又高 ，那里的城镇又大，城墙又坚固，如天一样高，并且我们在那里看见 亚衲 族人。’
DEUT|1|29|我就对你们说：‘不要惊惶，也不要怕他们。
DEUT|1|30|在你们前面行的耶和华－你们的上帝必为你们争战，正如他在 埃及 ，在你们眼前为你们所做的一样；
DEUT|1|31|并且你们在旷野所行的一切路上，也看见了耶和华─你们的上帝背着你们，如同人背自己的儿子一样，直到你们来到这地方。’
DEUT|1|32|你们在这事上却不信耶和华─你们的上帝。
DEUT|1|33|他一路行在你们前面，为你们寻找安营的地方；他夜间在火中，日间在云中，指示你们当走的路。”
DEUT|1|34|“耶和华听见你们的怨言，就发怒，起誓说：
DEUT|1|35|‘这邪恶世代的人，一个也不得看见我起誓要赐给你们列祖的美地；
DEUT|1|36|惟有 耶孚尼 的儿子 迦勒 必得看见，并且我要将他所踏过的地赐给他和他的子孙，因为他专心跟从我。’
DEUT|1|37|耶和华也因你们的缘故向我发怒，说：‘你也不得进入那地。
DEUT|1|38|那侍候你， 嫩 的儿子 约书亚 必得进入那地。你要勉励他，因为他要使 以色列 承受那地为业。
DEUT|1|39|你们的孩子，你们说要成为掳物的，就是今日尚不知善恶的儿女，必进入那地。我要将那地赐给他们，他们必得为业。
DEUT|1|40|至于你们，要转回，从 红海 的路往旷野去。’
DEUT|1|41|“你们回答我说：‘我们得罪了耶和华！现在我们愿遵照耶和华─我们上帝一切所吩咐的上去争战。’于是你们各人带着兵器，以为很容易就能上到山区去。
DEUT|1|42|耶和华对我说：‘你对他们说：不要上去，也不要争战，因我不在你们中间，恐怕你们在仇敌面前被击败。’
DEUT|1|43|我就告诉了你们，你们却不听从，竟违背耶和华的指示，擅自上到山区去。
DEUT|1|44|住在那山区的 亚摩利 人像蜂群一样出来迎击你们，追赶你们，在 西珥 击败你们，直到 何珥玛 。
DEUT|1|45|你们就回来，在耶和华面前哭泣；耶和华却不听你们的声音，也不向你们侧耳。
DEUT|1|46|你们照着所停留的日子，在 加低斯 停留了许多日子。”
DEUT|2|1|“我们转回，从 红海 的路往旷野去，正如耶和华所吩咐我的。我们在 西珥山 绕行了许多日子。
DEUT|2|2|耶和华对我说：
DEUT|2|3|‘你们绕行这山已经够久了，要转向北方。
DEUT|2|4|你要吩咐百姓说：你们弟兄 以扫 的子孙住在 西珥 ，你们要经过他们的边界。他们必惧怕你们，但你们要分外谨慎。
DEUT|2|5|不可向他们挑战；他们的地，连脚掌可踏之处，我都不给你们，因我已将 西珥山 赐给 以扫 为业。
DEUT|2|6|你们要用钱向他们买粮吃，也要用钱向他们买水喝。
DEUT|2|7|因为耶和华─你的上帝在你手里所做的一切事上已赐福给你。你走这大旷野，他都知道。这四十年，耶和华─你的上帝与你同在，因此你一无所缺。’
DEUT|2|8|“于是，我们经过我们弟兄 以扫 子孙所住的 西珥 ，从 亚拉巴 的路，经过 以拉他 、 以旬．迦别 ，转向 摩押 旷野的路去。
DEUT|2|9|耶和华对我说：‘不可侵犯 摩押 ，也不可向他们挑战。他们的地，我不赐给你为业，因我已将 亚珥 赐给 罗得 的子孙为业。’
DEUT|2|10|先前， 以米 人住在那里，百姓又大又多，像 亚衲 人一样高大。
DEUT|2|11|他们跟 亚衲 人一样，也算是 利乏音 人，但 摩押 人却称他们为 以米 人。
DEUT|2|12|从前， 何利 人也住在 西珥 ，但 以扫 的子孙把他们除灭，占领了他们的地，接续他们在那里居住，如同 以色列 在耶和华赐给他们为业之地所做的一样。
DEUT|2|13|‘现在，起来，过 撒烈溪 ！’于是我们过了 撒烈溪 。
DEUT|2|14|从离开 加低斯．巴尼亚 到渡过 撒烈溪 ，这段时期共三十八年，直到这一代的战士都从营中灭尽，正如耶和华向他们所起的誓。
DEUT|2|15|耶和华的手也攻击他们，将他们从营中除灭，直到灭尽。
DEUT|2|16|“百姓中所有的战士灭尽死亡以后，
DEUT|2|17|耶和华吩咐我说：
DEUT|2|18|‘你今日要经过 摩押 的边界 亚珥 ，
DEUT|2|19|走到 亚扪 人之地。不可侵犯他们，也不可向他们挑战。 亚扪 人的地，我不赐给你们为业，因我已将那地赐给 罗得 的子孙为业。’
DEUT|2|20|那地也算是 利乏音 人之地，因为先前 利乏音 人住在那里， 亚扪 人称他们为 散送冥 人。
DEUT|2|21|那里的百姓又大又多，像 亚衲 人一样高大，但耶和华从 亚扪 人面前除灭他们， 亚扪 人就占领他们的地，接续他们在那里居住。
DEUT|2|22|这正如耶和华从前为住在 西珥 的 以扫 子孙，将 何利 人从他们面前除灭，使他们得了 何利 人的地，接续他们在那里居住，直到今日一样。
DEUT|2|23|亚卫 人先前住在乡村直到 迦萨 ；从 迦斐托 出来的 迦斐托 人将 亚卫 人除灭，接续他们在那里居住。
DEUT|2|24|你们起来往前去，过 亚嫩谷 。看哪，我已将 亚摩利 人 希实本 王 西宏 和他的地交在你手中，你要开始去得他的地为业，向他挑战。
DEUT|2|25|从今日起，我要让天下万民因你惊慌惧怕，听见你的名声，就因你发颤伤恸。”
DEUT|2|26|“我从 基底莫 的旷野派遣使者到 希实本 王 西宏 那里，用和平的话说：
DEUT|2|27|‘求你让我穿越你的地，我走路的时候，只走大路，不偏左右。
DEUT|2|28|你可以卖粮给我吃，卖水给我喝；只要让我步行过去，
DEUT|2|29|就如住在 西珥 的 以扫 子孙和住在 亚珥 的 摩押 人待我一样，等我过了 约旦河 ，进入耶和华－我们上帝所赐给我们的地。’
DEUT|2|30|但 希实本 王 西宏 不肯让我们从他那里经过，因为耶和华－你的上帝使他性情顽梗，内心刚硬，为要把他交在你手中，像今日一样。
DEUT|2|31|耶和华对我说：‘看，我已开始把 西宏 和他的地交给你了，你要开始得他的地为业。’
DEUT|2|32|“ 西宏 和他的众百姓出来迎击我们，在 雅杂 与我们交战。
DEUT|2|33|耶和华－我们的上帝把他交给我们，我们就杀了他和他的众儿子，以及他所有的百姓。
DEUT|2|34|那时，我们夺了他一切的城镇，毁灭各城的男人、女人、孩子，没有留下一个幸存者。
DEUT|2|35|只有牲畜和所夺各城的财物，我们都取为自己的掠物。
DEUT|2|36|从 亚嫩谷 旁的 亚罗珥 和谷中的城，直到 基列 ，没有一座城是高得我们不能攻取的；耶和华－我们的上帝把它们全都交给我们了。
DEUT|2|37|只有 亚扪 人之地， 雅博河 沿岸，以及山区的城镇，你没有挨近，这全是耶和华－我们上帝所吩咐的。”
DEUT|3|1|“我们又转回，朝 巴珊 的路上去。 巴珊 王 噩 和他的众百姓出来迎击我们，在 以得来 与我们交战。
DEUT|3|2|耶和华对我说：‘不要怕他！因我已把他和他的众百姓，以及他的地，都交在你手中；你要待他像从前待住在 希实本 的 亚摩利 王 西宏 一样。’
DEUT|3|3|于是耶和华－我们的上帝也把 巴珊 王 噩 和他的众百姓都交在我们手中；我们杀了他，没有给他留下一个幸存者。
DEUT|3|4|那时，我们夺了他一切的城镇，共六十座，没有一座城不被我们所夺，这是 亚珥歌伯 的全境， 巴珊 王 噩 的国度。
DEUT|3|5|这些坚固的城都有高的城墙，有门有闩，此外，还有许多无城墙的乡村。
DEUT|3|6|我们把这些都毁灭了，像从前待 希实本 王 西宏 一样，毁灭各城的男人、女人、孩子；
DEUT|3|7|只有一切牲畜和城中的财物，我们取为自己的掠物。
DEUT|3|8|那时，我们从两个 亚摩利 王的手里把 约旦河 东边的地夺过来，从 亚嫩谷 直到 黑门山 ，
DEUT|3|9|这 黑门山 ， 西顿 人称为 西连 ， 亚摩利 人称为 示尼珥 。
DEUT|3|10|我们夺了平原的各城、 基列 全地、 巴珊 全地，直到 撒迦 和 以得来 ，都是 巴珊 王 噩 国内的城镇。
DEUT|3|11|利乏音 人所剩下的只有 巴珊 王 噩 。看哪，他的床是铁床，按照人肘的度量，长九肘，宽四肘，现今不是在 亚扪 人的 拉巴 吗？”
DEUT|3|12|“那时，我们得了这地。从 亚嫩谷 旁的 亚罗珥 起，连同 基列 山区的一半和境内的城镇，我都给了 吕便 人和 迦得 人。
DEUT|3|13|基列 其余的地和 巴珊 全地，就是 噩 的国度，我给了 玛拿西 半支派。 亚珥歌伯 全境就是 巴珊 全地，也称为 利乏音 人之地。
DEUT|3|14|玛拿西 的子孙 睚珥 占领了 亚珥歌伯 全境，直到 基述 人和 玛迦 人的边界，就按自己的名字称这些地，就是 巴珊 ，为 哈倭特．睚珥 ，直到今日。
DEUT|3|15|我又将 基列 给了 玛吉 。
DEUT|3|16|我给了 吕便 人和 迦得 人从 基列 到 亚嫩谷 ，以谷的中央为界，直到 亚扪 人边界的 雅博河 ；
DEUT|3|17|还有 亚拉巴 和靠近 约旦河 之地，从 基尼烈 直到 亚拉巴海 ，就是 盐海 ，以及 毗斯迦山 斜坡的山脚东边之地。
DEUT|3|18|“那时，我吩咐你们说：‘耶和华－你们的上帝已将这地赐给你们为业；你们所有的勇士都要带着兵器，在你们的弟兄 以色列 人前面过去。
DEUT|3|19|但你们的妻子、孩子、牲畜，可以住在我所赐给你们的各城里，我知道你们有许多牲畜。
DEUT|3|20|等到耶和华让你们的弟兄像你们一样，得享太平，他们在 约旦河 另一边，也得了耶和华－你们的上帝所赐给他们的地，你们各人才可以回到我所赐给你们为业之地。’
DEUT|3|21|那时，我吩咐 约书亚 说：‘你亲眼看见了耶和华－你们的上帝向这两个王一切所做的事，耶和华也必向你所要去的各国照样做。
DEUT|3|22|不要怕他们，因为那为你们争战的是耶和华－你们的上帝。’”
DEUT|3|23|“那时，我恳求耶和华说：
DEUT|3|24|‘主耶和华啊，你已开始将你的伟大和你大能的手显给你仆人看。在天上，在地下，有什么神明能像你行事，像你有大能的作为呢？
DEUT|3|25|求你让我过去，看 约旦河 另一边的美地，就是那佳美的山区和 黎巴嫩 。’
DEUT|3|26|但耶和华因你们的缘故向我发怒，不应允我。耶和华对我说：‘你够了吧！不要再向我提这事。
DEUT|3|27|你上 毗斯迦山 顶去，向东、西、南、北举目，用你的眼睛观看，因为你必不能过这 约旦河 。
DEUT|3|28|你却要吩咐 约书亚 ，勉励他，使他壮胆，因为他必在这百姓前面过去，使他们承受你所要观看之地。’
DEUT|3|29|于是我们停留在 伯．毗珥 对面的谷中。”
DEUT|4|1|“现在， 以色列 啊，听我所教导你们的律例典章，要遵行，好使你们存活，得以进入耶和华－你们列祖之上帝所赐给你们的地，承受为业。
DEUT|4|2|我吩咐你们的话，你们不可加添，也不可删减，好叫你们遵守耶和华－你们上帝的命令，就是我所吩咐你们的。
DEUT|4|3|你们已亲眼看见耶和华因 巴力．毗珥 所做的。凡随从 巴力．毗珥 的人，耶和华－你的上帝都从你中间除灭了。
DEUT|4|4|只有你们这紧紧跟随耶和华－你们上帝的人，今日全都存活。
DEUT|4|5|看，我照着耶和华－我的上帝所吩咐我的，将律例和典章教导你们，使你们在所要进去得为业的地上遵行。
DEUT|4|6|你们要谨守遵行；这就是你们在万民眼前的智慧和聪明。他们听见这一切律例，必说：‘这大国的人真是有智慧，有聪明！’
DEUT|4|7|哪一大国有神明与他们相近，像耶和华－我们的上帝在我们求告他的时候与我们相近呢？
DEUT|4|8|哪一大国有这样公义的律例典章，像我今日在你们面前所颁布的这一切律法呢？
DEUT|4|9|“但你要谨慎，殷勤保守你的心灵，免得忘记你亲眼所看见的事，又免得在你一生的年日这些事离开你的心，总要把它们传给你的子子孙孙。
DEUT|4|10|你在 何烈山 站在耶和华－你上帝面前的那日，耶和华对我说：‘你为我召集百姓，我要叫他们听见我的话，使他们活在世上的日子，可以学习敬畏我，又可以教导他们的儿女。’
DEUT|4|11|那时，你们近前来，站在山下；山上有火燃烧，直冲天顶，并有黑暗、密云、幽暗。
DEUT|4|12|耶和华从火焰中对你们说话，你们听见说话的声音，只有声音，却没有看见形像。
DEUT|4|13|他将所吩咐你们当守的约指示你们，就是十条诫命 ，并将诫命写在两块石版上。
DEUT|4|14|那时，耶和华吩咐我将律例典章教导你们，使你们在所要过去得为业的地上遵行。”
DEUT|4|15|“所以，你们为自己的缘故要分外谨慎；因为耶和华在 何烈山 ，从火中对你们说话的那日，你们没有看见任何形像。
DEUT|4|16|惟恐你们的行为败坏，为自己雕刻任何形状的偶像，无论是男像或女像，
DEUT|4|17|或地上任何走兽的像，或任何飞在空中有翅膀的鸟的像，
DEUT|4|18|或地上任何爬行动物的像，或地底下任何水中鱼的像。
DEUT|4|19|又恐怕你向天举目，看见耶和华－你的上帝为天下万民所摆列的日月星辰，就是天上的万象，就被诱惑去敬拜它们，事奉它们。
DEUT|4|20|耶和华将你们从 埃及 带领出来，脱离铁炉，是要你们成为他产业的子民，像今日一样。
DEUT|4|21|“耶和华又因你们的缘故向我发怒，起誓不容我过 约旦河 ，不让我进入耶和华－你上帝所赐你为业的那美地。
DEUT|4|22|我只好死在这地，不能过 约旦河 ；但你们必过去得那美地。
DEUT|4|23|你们要谨慎，免得忘记耶和华－你们的上帝与你们所立的约，为自己雕刻任何形状的偶像，就是耶和华－你上帝所禁止的，
DEUT|4|24|因为耶和华－你的上帝是吞灭的火，是忌邪 的上帝。
DEUT|4|25|“你们在那地住久了，生子生孙，若行为败坏，为自己雕刻任何形状的偶像，行耶和华－你上帝眼中看为恶的事，惹他发怒，
DEUT|4|26|我今日呼天唤地向你们作见证，你们在过 约旦河 得为业的地上必迅速灭亡！你们在那地的日子必不长久，必全然灭绝。
DEUT|4|27|耶和华必将你们分散在万民中；在耶和华领你们到的列国中，你们剩下的人丁稀少。
DEUT|4|28|在那里，你们必事奉人手所造的神明，它们是木头，是石头，不能看，不能听，不能吃，不能闻。
DEUT|4|29|你们在那里必寻求耶和华－你的上帝。你若尽心尽性寻求他，就必寻见。
DEUT|4|30|日后你在患难中，当这一切的事临到你，你必归回耶和华－你的上帝，听从他的话。
DEUT|4|31|耶和华－你的上帝是有怜悯的上帝，他不撇下你，不灭绝你，也不忘记他起誓与你列祖所立的约。
DEUT|4|32|“你去问，在你先前的时代，自从上帝造人在地上以来，从天这边到天那边，曾有过或听过这样的大事吗？
DEUT|4|33|有哪些百姓听见上帝在火中说话的声音，像你听见了还能存活呢？
DEUT|4|34|上帝何曾为自己尝试从别的国中领出一国的子民来，用考验、神迹、奇事、战争、大能的手、伸出来的膀臂和大可畏的事，像耶和华－你们的上帝在 埃及 ，在你们眼前为你们所做的一切事呢？
DEUT|4|35|这是要显给你看，使你知道，惟有耶和华他是上帝，除他以外，再没有别的了。
DEUT|4|36|他从天上使你听见他的声音，为要教导你，又在地上使你看见他的烈火，并且听见他从火中所说的话。
DEUT|4|37|因为他爱你的列祖，拣选他们的后裔 ，亲自用大能领你出了 埃及 ，
DEUT|4|38|要将比你强大的列国从你面前赶出，领你进去，把他们的地赐你为业，像今日一样。
DEUT|4|39|所以，今日你要知道，也要记在心里，天上地下惟有耶和华他是上帝，再没有别的了。
DEUT|4|40|我今日吩咐你的律例诫命，你要遵守，使你和你的后裔可以得福，并使你的日子一直在耶和华－你上帝赐你的地上得以长久。”
DEUT|4|41|“那时， 摩西 在 约旦河 东边，向日出的方向，指定三座城，
DEUT|4|42|使那素无仇恨、无意中杀了邻舍的凶手，可以逃到这三座城中的一座，就得存活：
DEUT|4|43|属 吕便 人的是旷野平坦之地的 比悉 ，属 迦得 人的是 基列 的 拉末 ，属 玛拿西 人的是 巴珊 的 哥兰 。”
DEUT|4|44|这是 摩西 在 以色列 人面前颁布的律法。
DEUT|4|45|这些法度、律例、典章是 摩西 在 以色列 人出 埃及 后对他们说的，
DEUT|4|46|在 约旦河 东 伯毗珥 对面的谷中，在住 希实本 的 亚摩利 王 西宏 之地；这 西宏 是 摩西 和 以色列 人出 埃及 后所击杀的。
DEUT|4|47|他们得了他的地，又得了 巴珊 王 噩 的地，就是两个 亚摩利 王，在 约旦河 东，向日出方向的地：
DEUT|4|48|从 亚嫩谷 旁的 亚罗珥 ，直到 西云山 ，就是 黑门山 ，
DEUT|4|49|还有 约旦河 东的整个 亚拉巴 ，向日出方向，直到 亚拉巴海 ，靠近 毗斯迦山 斜坡的山脚。
DEUT|5|1|摩西 召集 以色列 众人，对他们说：“ 以色列 啊，要听我今日在你们耳中所吩咐的律例典章，要学习，谨守遵行。
DEUT|5|2|耶和华－我们的上帝在 何烈山 与我们立约。
DEUT|5|3|这约耶和华不是与我们列祖立的，而是与我们，就是今日在这里还活着的人立的。
DEUT|5|4|耶和华在山上，从火中，面对面与你们说话。
DEUT|5|5|那时我站在耶和华和你们之间，要将耶和华的话传给你们，因为你们惧怕那火，没有上山。他说：
DEUT|5|6|“‘我是耶和华－你的上帝，曾将你从 埃及 地为奴之家领出来。
DEUT|5|7|“‘除了我以外，你不可有别的神。
DEUT|5|8|“‘不可为自己雕刻偶像，也不可做什么形像，仿佛上天、下地和地底下水中的百物。
DEUT|5|9|不可跪拜那些像，也不可事奉它们，因为我耶和华－你的上帝是忌邪 的上帝。恨我的，我必惩罚他们的罪，自父及子，直到三、四代；
DEUT|5|10|爱我、守我诫命的，我必向他们施慈爱，直到千代。
DEUT|5|11|“‘不可妄称耶和华－你上帝的名，因为妄称耶和华名的，耶和华必不以他为无罪。
DEUT|5|12|“‘当守安息日为圣日，正如耶和华－你上帝所吩咐的。
DEUT|5|13|六日要劳碌做你一切的工，
DEUT|5|14|但第七日是向耶和华－你的上帝当守的安息日。这一日，你和你的儿女、仆婢、牛、驴、牲畜，以及你城里寄居的客旅，都不可做任何的工，使你的仆婢可以和你一样休息。
DEUT|5|15|你要记念你在 埃及 地作过奴仆，耶和华－你的上帝用大能的手和伸出来的膀臂领你从那里出来。因此，耶和华－你的上帝吩咐你守安息日。
DEUT|5|16|“‘当孝敬父母，正如耶和华－你上帝所吩咐的，使你得福，并使你的日子在耶和华－你上帝所赐给你的地上得以长久。
DEUT|5|17|“‘不可杀人。
DEUT|5|18|“‘不可奸淫。
DEUT|5|19|“‘不可偷盗。
DEUT|5|20|“‘不可做假见证陷害你的邻舍。
DEUT|5|21|“‘不可贪恋你邻舍的妻子；也不可贪图你邻舍的房屋、田地、仆婢、牛驴，以及他一切所有的。’
DEUT|5|22|“这些话是耶和华在山上，从火焰、密云、幽暗中，大声吩咐你们全会众的，再没有加添别的话了。他把这些话写在两块石版上，交给我。
DEUT|5|23|山被火焰烧着，你们听见从黑暗中发出的声音，那时，你们各支派的领袖和长老都挨近我。
DEUT|5|24|你们说：‘看哪，耶和华－我们的上帝将他的荣耀和他的伟大显给我们看，我们也听见他从火中发出的声音。今日我们看到上帝与人说话，人还活着。
DEUT|5|25|现在这大火将要吞灭我们，我们何必死呢？若再听见耶和华我们上帝的声音，我们就必死。
DEUT|5|26|凡血肉之躯，有谁像我们一样，听见了永生上帝从火中讲话的声音还能活着呢？
DEUT|5|27|求你近前去，听耶和华－我们上帝所要说的一切话，将耶和华－我们上帝对你说的话都传给我们，我们就听从遵行。’
DEUT|5|28|“你们对我说的话，耶和华都听见了。耶和华对我说：‘这百姓对你说的话，我听见了；他们所说的都对。
DEUT|5|29|惟愿他们存这样的心敬畏我，常遵守我一切的诫命，使他们和他们的子孙永远得福。
DEUT|5|30|你去对他们说：你们回帐棚去吧！
DEUT|5|31|至于你，可以站在我这里，我要将一切诫命、律例、典章传给你。你要教导他们，使他们在我赐他们为业的地上遵行。’
DEUT|5|32|所以，你们要照耶和华－你们上帝所吩咐的谨守遵行，不可偏离左右。
DEUT|5|33|你们要走耶和华－你们的上帝所吩咐的一切道路，使你们可以存活得福，并使你们的日子在所要承受的地上得以长久。”
DEUT|6|1|“这是耶和华－你们的上帝所吩咐要教导你们的诫命、律例、典章，叫你们在所要过去得为业的地上遵行，
DEUT|6|2|好叫你和你的子孙在一生的日子都敬畏耶和华－你的上帝，谨守他的一切律例、诫命，就是我所吩咐你的，使你的日子得以长久。
DEUT|6|3|以色列 啊，你要听，要谨守遵行，使你可以在那流奶与蜜之地得福，人数极其增多，正如耶和华－你列祖的上帝所应许你的。
DEUT|6|4|“ 以色列 啊，你要听！耶和华－我们的上帝是独一的主 。
DEUT|6|5|你要尽心、尽性、尽力爱耶和华－你的上帝。
DEUT|6|6|我今日吩咐你的这些话都要记在心上，
DEUT|6|7|也要殷勤教导你的儿女。无论你坐在家里，走在路上，躺下，起来，都要吟诵。
DEUT|6|8|要系在手上作记号，戴在额上 作经匣 ；
DEUT|6|9|又要写在你房屋的门框上和你的城门上。
DEUT|6|10|“耶和华－你的上帝必领你进他向你列祖 亚伯拉罕 、 以撒 、 雅各 起誓要给你的地。那里有又大又美的城镇，不是你建造的；
DEUT|6|11|有装满各样美物的房屋，不是你装满的；有挖成的水井，不是你挖的；有葡萄园、橄榄园，不是你栽植的；你吃了而且饱足。
DEUT|6|12|你要谨慎，免得你忘记领你从 埃及 地为奴之家出来的耶和华。
DEUT|6|13|你要敬畏耶和华－你的上帝，事奉他，奉他的名起誓。
DEUT|6|14|不可随从别神，就是你们四围民族的众神明，
DEUT|6|15|因为在你中间的耶和华－你的上帝是忌邪 的上帝，恐怕耶和华－你上帝的怒气向你发作，把你从地上除灭。
DEUT|6|16|“你们不可试探耶和华－你们的上帝，像你们在 玛撒 那样试探他。
DEUT|6|17|要谨慎遵守耶和华－你们上帝的诫命，和他所吩咐的法度、律例。
DEUT|6|18|耶和华眼中看为正直和美善的事，你都要遵行，使你得福，可以进去得耶和华向你列祖起誓应许的美地，
DEUT|6|19|可以从你面前赶出你所有的仇敌，正如耶和华所说的。
DEUT|6|20|“日后，你的儿子问你说：‘耶和华－我们上帝吩咐你们的法度、律例、典章是什么意思呢？’
DEUT|6|21|你要告诉你的儿子说：‘我们在 埃及 作过法老的奴仆，耶和华用大能的手将我们从 埃及 领出来。
DEUT|6|22|在我们眼前，他施行重大可怕的神迹奇事对付 埃及 、法老和他的全家。
DEUT|6|23|他将我们从那里领出来，为要领我们进入他向我们列祖起誓应许之地，把这地赐给我们。
DEUT|6|24|耶和华又吩咐我们遵行这一切的律例，敬畏耶和华－我们的上帝，使我们一生得福，得以存活，像今日一样。
DEUT|6|25|我们若照耶和华－我们上帝所吩咐的，在他面前谨守遵行这一切诫命，这就是我们的义了。’”
DEUT|7|1|“耶和华－你的上帝领你进入你要得为业之地，从你面前赶出许多国家，就是比你更强大的七个国家： 赫 人、 革迦撒 人、 亚摩利 人、 迦南 人、 比利洗 人、 希未 人、 耶布斯 人。
DEUT|7|2|当耶和华－你的上帝把他们交给你，你击杀他们的时候，你要完全消灭他们，不可与他们立约，也不可怜惜他们。
DEUT|7|3|不可与他们结亲；不可将你的女儿嫁给他的儿子，也不可叫你的儿子娶他的女儿。
DEUT|7|4|因为他必使你的儿女离弃我，去事奉别神，以致耶和华的怒气向你们发作，迅速将你除灭。
DEUT|7|5|你们却要这样处置他们：拆毁他们的祭坛，打碎他们的柱像，砍断他们的 亚舍拉 ，用火焚烧他们雕刻的偶像。
DEUT|7|6|“因为你是属于耶和华－你上帝神圣的子民；耶和华－你的上帝从地面上的万民中拣选你，作自己宝贵的子民。
DEUT|7|7|耶和华专爱你们，拣选你们，并非因你们人数比任何民族多，其实你们的人数在各民族中是最少的。
DEUT|7|8|因为耶和华爱你们，又因要遵守他向你们列祖所起的誓，耶和华就用大能的手领你们出来，救赎你脱离为奴之家，脱离 埃及 王法老的手。
DEUT|7|9|所以，你知道耶和华－你的上帝，他是上帝，是信实的上帝。他向爱他、守他诫命的人守约施慈爱，直到千代；
DEUT|7|10|向恨他的人，他必当面报应，消灭他们。凡恨他的，他必当面报应，绝不迟延。
DEUT|7|11|所以，你要谨守我今日所吩咐你的诫命、律例、典章，遵行它们。”
DEUT|7|12|“你们若听从这些典章，谨守遵行，耶和华－你的上帝必照他向你列祖所起的誓，对你守约，施慈爱。
DEUT|7|13|他必爱你，赐福给你，使你人数增多，也必在他向你列祖起誓要给你的地上赐福给你身所生的，你地所产的，你的五谷、新酒和新的油，以及你的牛犊、羔羊。
DEUT|7|14|你必蒙福胜过万民；你没有不育的男人和不孕的女人，牲畜也没有不生育的。
DEUT|7|15|耶和华必使一切的疾病远离你；你所知道 埃及 各样的恶疾，他不加在你身上，反要加在所有恨你的人身上。
DEUT|7|16|你要吞灭耶和华－你的上帝交给你的各民族，你的眼目不可顾惜他们。你也不可事奉他们的神明，因为这必成为你的圈套。
DEUT|7|17|“你若心里说，这些国的人数比我多，我怎能赶出他们呢？
DEUT|7|18|你不必怕他们，要牢牢记住耶和华－你上帝向法老和 埃及 全地所行的事，
DEUT|7|19|你亲眼见过的大考验、神迹、奇事、大能的手和伸出来的膀臂，都是耶和华－你上帝领你出来所施行的。耶和华－你的上帝也必照样处置你所惧怕的各民族，
DEUT|7|20|并且耶和华－你的上帝必派瘟疫 攻击他们，直到那剩下而躲起来的人都从你面前灭亡。
DEUT|7|21|不要因他们惊恐，因为耶和华－你的上帝在你中间是大而可畏的上帝。
DEUT|7|22|耶和华－你的上帝必将这些国从你面前渐渐赶出；你不可迅速把他们消灭，免得野地的走兽多起来危害你。
DEUT|7|23|耶和华－你的上帝必将他们交给你，大大扰乱他们，直到他们被除灭。
DEUT|7|24|他又要将他们的君王交在你手中，你必从天下除去他们的名；必无一人能在你面前站立得住，直到你把他们除灭了。
DEUT|7|25|你们要用火焚烧他们神明的雕刻偶像；不可贪爱偶像上的金银，也不可私自收起来，免得你因此陷入圈套，因为这是耶和华－你上帝所憎恶的。
DEUT|7|26|你不可把可憎之物带进你的家，否则，你就像它一样成为当毁灭的。你要彻底憎恨它，极其厌恶它，因为这是当毁灭的。”
DEUT|8|1|“我今日所吩咐你的一切诫命，你们要谨守遵行，好使你们存活，人数增多，可以进去得耶和华向你们列祖起誓应许的那地。
DEUT|8|2|你要记得，这四十年耶和华─你的上帝在旷野一路引导你，是要磨炼你，考验你，为要知道你的心如何，是否愿意遵守他的诫命。
DEUT|8|3|他磨炼你，任你饥饿，将你和你列祖所不认识的吗哪赐给你吃，使你知道，人活着，不是单靠食物，乃是靠耶和华口里所出的一切话。
DEUT|8|4|这四十年，你身上的衣服没有穿破，你的脚也没有肿。
DEUT|8|5|你心里要知道，耶和华─你的上帝管教你，像人管教儿女一样。
DEUT|8|6|你要谨守耶和华─你上帝的诫命，遵行他的道，敬畏他。
DEUT|8|7|“耶和华─你的上帝必领你进入美地，那地有河流，有泉源和深渊的水从谷中和山上流出。
DEUT|8|8|那地有小麦、大麦、葡萄树、无花果树、石榴树，那地也有橄榄油和蜂蜜。
DEUT|8|9|那地没有缺乏，你在那里有食物吃，一无所缺；那地的石头是铁，山中可以挖铜。
DEUT|8|10|你吃得饱足，要称颂耶和华─你的上帝，因为他将那美地赐给你。”
DEUT|8|11|“你要谨慎，免得忘记耶和华─你的上帝，不守他的诫命、典章、律例，就是我今日吩咐你的。
DEUT|8|12|免得你吃得饱足，建造上好的房屋，住在其中，
DEUT|8|13|你的牛羊增多，你的金银增多，你拥有的一切全都增多，
DEUT|8|14|于是你的心高傲，忘记耶和华─你的上帝。他曾将你从 埃及 地为奴之家领出来，
DEUT|8|15|曾引领你经过那大而可怕的旷野，有火蛇、蝎子、干旱无水之地。他也曾为你使水从坚硬的磐石中流出来，
DEUT|8|16|又在旷野将你列祖所不认识的吗哪赐给你吃，为要磨炼你，考验你，终久使你享福。
DEUT|8|17|你心里说：‘这财富是我的力量、我手的能力得来的。’
DEUT|8|18|你要记得耶和华─你的上帝，因为得财富的能力是他给你的，为要坚守他向你列祖起誓所立的约，像今日一样。
DEUT|8|19|你若忘记耶和华─你的上帝，随从别神，事奉它们，敬拜它们，我今日警告你们，你们必定灭亡。
DEUT|8|20|耶和华在你们面前怎样使列国灭亡，你们也必照样灭亡，因为你们不听从耶和华─你们上帝的话。”
DEUT|9|1|“ 以色列 啊，你要听！你今日要过 约旦河 ，进去占领比你更强大的列国，那里的城镇又大，城墙又坚固，如天一样高。
DEUT|9|2|那里的百姓是 亚衲 族人，又高又壮，是你所知道的；你也听说过：‘谁能在 亚衲 族人面前站立得住呢？’
DEUT|9|3|你今日应当知道，耶和华─你的上帝在你前面渡过去，如同吞噬的火，要除灭他们，并要在你面前将他们制伏，使你可以赶出他们，速速消灭他们，正如耶和华向你所说的。
DEUT|9|4|“耶和华─你的上帝将他们从你面前赶出以后，你心里不可说：‘耶和华领我得这地是因我的义。’其实，耶和华将这些国家从你面前赶出去是因他们的恶。
DEUT|9|5|你能进去得他们的地，并不是因你的义，也不是因你心里正直，而是因这些国家的恶，耶和华─你的上帝才把他们从你面前赶出去，为了应验耶和华向你列祖 亚伯拉罕 、 以撒 、 雅各 起誓应许的话。
DEUT|9|6|“你当知道，耶和华─你的上帝将这美地赐你为业，并不是因你的义；你本是硬着颈项的百姓。
DEUT|9|7|你要记得，不要忘记，你在旷野怎样惹耶和华－你的上帝发怒。自从你出了 埃及 地的那日，直到你们来到这地方，你们常常悖逆耶和华。
DEUT|9|8|你们在 何烈山 惹耶和华发怒，耶和华对你们动怒，甚至要除灭你们。
DEUT|9|9|我上了山，要领受两块石版，就是耶和华与你们立约的版。那时我在山上住了四十昼夜，没有吃饭，也没有喝水。
DEUT|9|10|耶和华把那两块石版交给我，是上帝用指头写成的；版上是耶和华在大会的那一天，在山上从火中对你们所说的一切话。
DEUT|9|11|过了四十昼夜，耶和华把那两块石版，就是约版，交给我。
DEUT|9|12|耶和华对我说：‘起来，赶快从这里下去！因为你从 埃及 领出来的百姓已经败坏了；他们这么快偏离了我所吩咐的道，为自己铸造偶像。’
DEUT|9|13|“耶和华对我说：‘我看这百姓，看哪，他们是硬着颈项的百姓。
DEUT|9|14|你且由着我，我要除灭他们，从天下涂去他们的名，我要使你成为比他们更大更强的国。’
DEUT|9|15|于是我转身下山，山上有火燃烧，两块约版在我双手中。
DEUT|9|16|我观看，看哪，你们得罪了耶和华－你们的上帝，为自己铸成了一头牛犊，迅速偏离了耶和华所吩咐你们的道，
DEUT|9|17|我拿着那两块石版，从我双手中扔出去，在你们眼前把它们摔碎了。
DEUT|9|18|因为你们所犯的一切罪，做了耶和华眼中看为恶的事，惹他发怒，我就像从前一样俯伏在耶和华面前四十昼夜，没有吃饭，没有喝水。
DEUT|9|19|我很害怕，因为耶和华向你们大发烈怒，要除灭你们。但那一次耶和华又应允了我。
DEUT|9|20|耶和华也向 亚伦 非常生气，甚至要除灭他；那时我也为 亚伦 祈祷。
DEUT|9|21|我把那使你们犯罪所铸的牛犊拿来，用火焚烧，捣碎后再磨成粉末，好像灰尘。我把这灰尘撒在从山上流下来的溪水中。
DEUT|9|22|“你们在 他备拉 、 玛撒 、 基博罗．哈他瓦 又惹耶和华发怒。
DEUT|9|23|耶和华叫你们离开 加低斯．巴尼亚 ，说：‘你们上去得我所赐给你们的地。’那时，你们违背了耶和华－你们上帝的指示，不信服他，不听从他的话。
DEUT|9|24|自从我认识你们的日子以来，你们常常悖逆耶和华。
DEUT|9|25|“我因耶和华说要除灭你们，就在耶和华面前俯伏四十昼夜，像我以前俯伏一样。
DEUT|9|26|我向耶和华祈祷，说：‘主耶和华啊，求你不要灭绝你的百姓，你的产业。他们是你用大能救赎，用你强有力的手从 埃及 领出来的。
DEUT|9|27|求你记念你的仆人 亚伯拉罕 、 以撒 、 雅各 ，不看这百姓的顽梗、邪恶、罪愆，
DEUT|9|28|免得你领我们出来的那地之人说：耶和华因为不能将这百姓领进他所应许之地，又因恨他们，所以领他们出去，要在旷野杀他们。
DEUT|9|29|其实他们是你的百姓，你的产业，是你用大能和伸出的膀臂领出来的。’”
DEUT|10|1|“那时，耶和华对我说：‘你要凿出两块石版，和先前的一样，上山到我这里来。你也要造一个木柜。
DEUT|10|2|我要把你先前摔碎的版上所写的字，写在这版上；你要把这版放在柜里。’
DEUT|10|3|于是我用金合欢木造了一个柜子，又凿出两块石版，和先前的一样。我手里拿着这两块版上山。
DEUT|10|4|耶和华将那大会之日、在山上从火中所吩咐你们的十条诫命，照先前所写的写在这版上。耶和华把它们交给我。
DEUT|10|5|我转身下山，将这版放在我所造的柜里，现今这版还在那里，正如耶和华所吩咐我的。
DEUT|10|6|（ 以色列 人从 比罗比尼．亚干 起行，来到 摩西拉 ， 亚伦 死在那里，就葬在那里。他的儿子 以利亚撒 接续他担任祭司的职分。
DEUT|10|7|他们从那里起行，来到 谷歌大 ，又从 谷歌大 来到 约巴他 ，有溪水之地。
DEUT|10|8|那时，耶和华将 利未 支派分别出来，抬耶和华的约柜，又侍立在耶和华面前事奉他，奉他的名祝福，直到今日。
DEUT|10|9|因此， 利未 没有像他的弟兄有产业，耶和华是他的产业，正如耶和华－你上帝所应许他的。）
DEUT|10|10|“我又像先前一样在山上停留了四十昼夜。这一次耶和华也应允我，不将你灭绝。
DEUT|10|11|耶和华对我说：‘起来，走在百姓前面，领他们进去得我向他们列祖起誓要给他们的地。’”
DEUT|10|12|“ 以色列 啊，现在耶和华－你的上帝向你要的是什么呢？只要你敬畏耶和华－你的上帝，遵行他一切的道，爱他，尽心尽性事奉耶和华－你的上帝，
DEUT|10|13|遵守耶和华的诫命律例，就是我今日所吩咐你的，为要使你得福。
DEUT|10|14|看哪，天和天上的天，地和地上所有的，都属耶和华－你的上帝。
DEUT|10|15|然而，耶和华专爱你的列祖，爱他们，从万民中拣选你们，就是他们的后裔，像今日一样。
DEUT|10|16|所以你们的心要受割礼，不可再硬着颈项。
DEUT|10|17|因为耶和华－你们的上帝是万神之神，万主之主，是伟大、强有力、可畏的上帝，不看人的情面，也不受贿赂。
DEUT|10|18|他为孤儿寡妇伸冤，爱护寄居的，赐给他衣食。
DEUT|10|19|所以你们要爱护寄居的，因为你们在 埃及 地也作过寄居的。
DEUT|10|20|你要敬畏耶和华－你的上帝，事奉他，紧紧跟随他，奉他的名起誓。
DEUT|10|21|他是你当赞美的，是你的上帝，为你做了大而可畏的事，这些是你亲眼见过的。
DEUT|10|22|你的列祖七十人下 埃及 ，现在耶和华－你的上帝却使你如同天上的星那样多。”
DEUT|11|1|“你要爱耶和华－你的上帝，天天遵守他的吩咐、律例、典章、诫命。
DEUT|11|2|今日你们应当知道，而不是你们的儿女，因为他们不知道，也没有见过耶和华─你们上帝的管教、他的伟大、他大能的手和伸出来的膀臂，
DEUT|11|3|以及他在 埃及 向 埃及 王法老和其全地所行的神迹奇事；
DEUT|11|4|他怎样对待 埃及 的军队、马和战车，他们追赶你们的时候，耶和华怎样用 红海 的水淹没他们，消灭了他们，直到今日；
DEUT|11|5|他在旷野怎样待你们，直到你们来到这地方，
DEUT|11|6|以及他怎样待 吕便 子孙， 以利押 的儿子 大坍 、 亚比兰 ，地怎样在 以色列 人中开了裂口，吞了他们和他们的家眷，帐棚，以及跟他们在一起所有活着的。
DEUT|11|7|惟有你们亲眼见过耶和华所做的一切大事。”
DEUT|11|8|“所以，你们要遵守我今日所吩咐的一切诫命，使你们刚强，可以进去得你们所要得的那地，就是你们将过河到那里要得的，
DEUT|11|9|也使你们的日子，在耶和华向你们列祖起誓要给他们和他们后裔的地上得以长久，那是流奶与蜜之地。
DEUT|11|10|你要进去得为业的那地，不像你出来的 埃及 地。在 埃及 ，你撒种后，要用脚浇灌，像浇灌菜园一样。
DEUT|11|11|你们要过去得为业的那地乃是有山有谷、天上的雨水滋润之地，
DEUT|11|12|是耶和华－你上帝所眷顾的地；从岁首到年终，耶和华－你上帝的眼目时常看顾那地。
DEUT|11|13|“你们若留心听从我今日所吩咐你们的诫命，爱耶和华－你们的上帝，尽心尽性事奉他，
DEUT|11|14|我 必按时降下雨水在你们的地上，就是秋雨和春雨，使你们可以收藏五谷、新酒和新的油，
DEUT|11|15|也必使田野为你的牲畜长出草来；这样，你必吃得饱足。
DEUT|11|16|你们要谨慎，免得心受诱惑，转去事奉别神，敬拜它们，
DEUT|11|17|以致耶和华的怒气向你们发作，使天封闭不下雨，使地不出产，使你们在耶和华所赐给你们的美地上速速灭亡。
DEUT|11|18|“你们要将我这些话存在心里，留在意念中，系在手上作记号，戴在额上 作经匣。
DEUT|11|19|你们也要将这些话教导你们的儿女，无论坐在家里，行在路上，躺下，起来，都要讲论，
DEUT|11|20|又要写在房屋的门框上和你的城门上。
DEUT|11|21|这样，你们和你们子孙的日子必在耶和华向你们列祖起誓要给他们的地上得以增多，如天地之长久。
DEUT|11|22|你们若留心谨守遵行我所吩咐这一切的诫命，爱耶和华－你们的上帝，遵行他一切的道，紧紧跟随他，
DEUT|11|23|他必从你们面前赶出这一切国家，你们也要占领比你们更大更强的国家。
DEUT|11|24|凡你们脚掌所踏之地都必归于你们；从旷野到 黎巴嫩 ，从 幼发拉底 大河，直到西边的海，都要成为你们的疆土。
DEUT|11|25|必无一人能在你们面前站立得住；耶和华－你们的上帝必照他所说的，使惧怕惊恐临到你们所踏的全地。
DEUT|11|26|“看，我今日将祝福与诅咒都陈明在你们面前。
DEUT|11|27|你们若听从耶和华─你们上帝的诫命，就是我今日所吩咐你们的，就必蒙福。
DEUT|11|28|你们若不听从耶和华─你们上帝的诫命，偏离我今日所吩咐你们的道，去随从你们所不认识的别神，就必受诅咒。
DEUT|11|29|当耶和华－你的上帝领你进入要得为业的那地，你就要在 基利心山 上宣布祝福，在 以巴路山 上宣布诅咒。
DEUT|11|30|这二座山岂不是在 约旦河 的那边，日落的方向，在住 亚拉巴 的 迦南 人之地， 吉甲 的前面，靠近 摩利 橡树吗？
DEUT|11|31|你们过 约旦河 ，进去得耶和华－你们的上帝所赐你们为业之地；当你们占领它，在那地居住的时候，
DEUT|11|32|你们要谨守遵行我今日在你们面前颁布的一切律例典章。”
DEUT|12|1|“你们活在世上的日子，在耶和华─你列祖的上帝所赐你为业的地上，你们要谨守遵行这些律例典章：
DEUT|12|2|你们占领的国家所事奉他们众神明的地方，无论是在高山，在小山，在一切的青翠树下，你们要彻底毁坏；
DEUT|12|3|要拆毁他们的祭坛，打碎他们的柱像，用火焚烧他们的 亚舍拉 ，砍断他们神明的雕刻偶像，并要从那地方除去他们的名。
DEUT|12|4|你们不可那样敬拜耶和华－你们的上帝。
DEUT|12|5|但耶和华－你们的上帝在你们各支派中选择何处作为立他名的居所，你们就要到那里求问，
DEUT|12|6|将你们的燔祭、祭物、十一奉献、手中的举祭、还愿祭、甘心祭，以及牛群羊群中头生的，都带到那里。
DEUT|12|7|在那里，你们和你们的全家都可以在耶和华─你们上帝的面前吃，并且因你们手所做的一切蒙耶和华－你的上帝赐福而欢乐。
DEUT|12|8|你们不可做像我们今日在这里所做的，各人行自己眼中看为正的一切事；
DEUT|12|9|因为你们现在还没有进入耶和华－你上帝所赐你的安息，所给你的产业。
DEUT|12|10|你们过了 约旦河 ，住在耶和华─你们上帝给你们承受为业的地；他又使你们得享太平，不受四围一切仇敌扰乱，使你们安然居住。
DEUT|12|11|那时你们要将我所吩咐你们的燔祭、祭物、十一奉献、手中的举祭，和向耶和华许愿的一切上好的祭，都带到耶和华─你们上帝所选择立他名的居所。
DEUT|12|12|你们和儿女、仆婢，以及住在你们城里，没有与你们一起分得产业的 利未 人，都要在耶和华－你们的上帝面前欢乐。
DEUT|12|13|你要谨慎，不可在自己所看中的各处献燔祭。
DEUT|12|14|惟独耶和华从你的一个支派中所选择的地方，你要在那里献燔祭，在那里遵行我一切所吩咐你的。
DEUT|12|15|“然而，你在各城里都可以照着耶和华－你上帝所赐给你的福分，随心所欲宰牲吃肉；无论洁净的人不洁净的人都可以吃，就如吃羚羊和鹿的肉一样。
DEUT|12|16|只是血，你不可吃，要把它倒在地上，如同倒水一样。
DEUT|12|17|你的五谷、新酒和新油的十分之一，或是牛群羊群中头生的，或是你的许愿祭、甘心祭和手中的举祭，都不可在你的城里吃，
DEUT|12|18|必须在耶和华－你的上帝面前吃，在耶和华－你上帝所选择的地方，你和儿女、仆婢，以及住在你城里的 利未 人都可以吃，并要因你手所做的一切，在耶和华－你上帝面前欢乐。
DEUT|12|19|你要谨慎，在你所住的地上，你永不可离弃 利未 人。
DEUT|12|20|“耶和华－你的上帝照他的应许扩张你疆土的时候，你心里想要吃肉，说：‘我要吃肉’，就可以随心所欲吃肉。
DEUT|12|21|耶和华－你上帝选择立他名的地方若离你太远，你可以照我所吩咐的，将耶和华赐给你的牛羊取些宰了，随心所欲在你的城里吃。
DEUT|12|22|其实，就如吃羚羊和鹿的肉一样，你要这样吃它，无论洁净的人不洁净的人都可以一起吃。
DEUT|12|23|但是你要坚定，不可吃血，因为血是生命；不可将生命与肉一起吃。
DEUT|12|24|你不可吃血，要把它倒在地上，如同倒水一样。
DEUT|12|25|不可吃血，好让你和你的子孙可以得福，因为你行了耶和华眼中看为正的事。
DEUT|12|26|只是你分别为圣的物和你所还的愿，都要带到耶和华所选择的地方去。
DEUT|12|27|你的燔祭，连肉带血，都要献在耶和华－你上帝的坛上。祭物的血要倒在耶和华－你上帝的坛上；肉你可以吃。
DEUT|12|28|你要谨守听从我所吩咐的一切话，好让你和你的子孙可以永远得福，因为你行耶和华－你上帝眼中看为善、看为正的事。”
DEUT|12|29|“耶和华－你上帝把你要进去赶出的列国从你面前剪除，并且你得了他们的地为业居住，
DEUT|12|30|那时你要谨慎，在他们从你面前被除灭之后，你不可受引诱随从他们，也不可求问他们的神明，说：‘这些国家怎样事奉他们的神明，我也要照样做。’
DEUT|12|31|你不可向耶和华－你的上帝这样做，因为他们向他们的神明做了耶和华所憎恨、所厌恶的一切事，甚至将自己的儿女用火焚烧，献给他们的神明。
DEUT|12|32|凡我所吩咐你们的事，你们都要谨守遵行，不可加添，也不可删减。”
DEUT|13|1|“你中间若有先知或是做梦的人起来，向你显神迹奇事，
DEUT|13|2|他对你说的神迹奇事应验了，说：‘我们去随从别神，事奉它们吧。’那是你不认识的。
DEUT|13|3|你不可听那先知或是那做梦之人的话，因为这是耶和华－你们的上帝考验你们，要知道你们是否尽心尽性爱耶和华－你们的上帝。
DEUT|13|4|你们要顺从耶和华－你们的上帝，敬畏他，谨守他的诫命，听从他的话，事奉他，紧紧跟随他。
DEUT|13|5|那先知或那做梦的人要被处死，因为他出言悖逆那领你们出 埃及 地、救赎你脱离为奴之家的耶和华－你们的上帝，要引诱你离开耶和华－你上帝吩咐你要行的道。这样，你就把恶从你中间除掉。
DEUT|13|6|“你的同胞兄弟，或是你的儿女，或是你怀中的妻，或是如同自己性命的朋友，若暗中引诱你，说：‘我们去事奉别神吧。’那是你和你列祖所不认识的，
DEUT|13|7|你四围列国的神明，无论是离你近或离你远，从地这边到地那边，
DEUT|13|8|你都不可附和他，也不要听从他。你的眼不可顾惜他，不可怜悯他，也不可袒护他。
DEUT|13|9|你务必杀他；你先下手，然后众百姓才下手，把他处死。
DEUT|13|10|要用石头打死他，因为他想引诱你离开那领你出 埃及 地为奴之家的耶和华－你的上帝。
DEUT|13|11|全 以色列 都要听见而害怕，不敢在你中间再行这样的恶事了。
DEUT|13|12|“若你听见人说，在耶和华－你上帝所赐给你居住的城镇中的一座，
DEUT|13|13|有些无赖之徒从你中间出来，引诱本城的居民，说：‘我们去事奉别神吧。’那是你们不认识的，
DEUT|13|14|你就要调查，探听，细心询问。看哪，是真的，确实有这可憎的事在你中间发生，
DEUT|13|15|你务必用刀杀那城里的居民，把城里所有的，连牲畜都用刀灭尽。
DEUT|13|16|你要把从城里所夺取的一切财物堆在广场中，用火将那城和其中夺取的一切财物全烧给耶和华－你的上帝。那城要永远成为废墟，不得重建。
DEUT|13|17|那当毁灭的物一点都不可粘你的手，好让耶和华转回，不向你发烈怒，却恩待你，怜悯你，照他向你列祖所起的誓使你人数增多；
DEUT|13|18|因为你听从耶和华－你上帝的话，遵守我今日所吩咐你的一切诫命，行耶和华－你上帝眼中看为正的事。”
DEUT|14|1|“你们是耶和华─你们上帝的儿女。不可为了死人割划自己，也不可使额上 光秃；
DEUT|14|2|因为你是属于耶和华－你上帝神圣的子民，耶和华从地面上的万民中拣选了你，作自己宝贵的子民。”
DEUT|14|3|“凡可憎的物， 你都不可吃。
DEUT|14|4|可吃的牲畜是：牛、绵羊、山羊、
DEUT|14|5|鹿、羚、麃子、野山羊、瞪羚、羚羊、山绵羊。
DEUT|14|6|凡蹄分两瓣，分趾蹄而又反刍食物的牲畜，你们都可以吃。
DEUT|14|7|但那反刍或分蹄之中不可吃的是：骆驼、兔子、石獾，虽然反刍却不分蹄，对你们是不洁净的；
DEUT|14|8|猪，虽然分蹄却不反刍，对你们也是不洁净的。它们的肉，你们一点都不可吃；它们的尸体，你们也不可摸。
DEUT|14|9|“水中可吃的是这些：凡有鳍有鳞的都可以吃；
DEUT|14|10|凡无鳍无鳞的都不可吃，对你们是不洁净的。
DEUT|14|11|“凡洁净的鸟，你们都可以吃。
DEUT|14|12|不可吃的是：雕、狗头雕、红头雕、
DEUT|14|13|鹯、小鹰、鹞鹰的类群，
DEUT|14|14|各种乌鸦的类群、
DEUT|14|15|鸵鸟、夜鹰、鱼鹰、鹰的类群、
DEUT|14|16|鸮鸟、猫头鹰、角鸱、
DEUT|14|17|鹈鹕、秃雕、鸬鹚、
DEUT|14|18|鹳、鹭鸶的类群、戴鵀与蝙蝠。
DEUT|14|19|凡有翅膀却爬行的群聚动物对你们是不洁净的，都不可吃。
DEUT|14|20|凡洁净的鸟，你们都可以吃。
DEUT|14|21|“凡自然死去的动物，你们都不可吃，可以给城里寄居的人吃，或卖给外人，因为你是属于耶和华－你上帝神圣的子民。 “不可用母山羊的奶来煮它的小山羊。”
DEUT|14|22|“每年，你务必从你播种的一切收成，田地所出产的，取十分之一献上。
DEUT|14|23|要在耶和华－你上帝面前，就是他选择那里作为他名居所的地方，吃你所献十分之一的五谷、新酒和新的油，以及牛群羊群中头生的，好让你天天学习敬畏耶和华－你的上帝。
DEUT|14|24|当耶和华－你的上帝赐福给你的时候，耶和华－你上帝选择立他名的地方若离你太远，路途太长，使你不能把这东西带到那里去，
DEUT|14|25|你可以把它换成银子，把银子包起来，拿在手中，往耶和华－你上帝所选择的地方去。
DEUT|14|26|在那里，你可以随心所欲用银子或买牛羊，或买清酒烈酒，或买任何你心所想的。你和你的全家要在耶和华－你上帝面前吃喝欢乐。
DEUT|14|27|“住在你城里的 利未 人，你不可离弃他，因为他在你那里没有分得产业。
DEUT|14|28|每三年的最后一年，你要把那一年收成的十分之一取出来，积存在你的城中；
DEUT|14|29|那没有与你一起分得产业的 利未 人，和城里的寄居者，以及孤儿寡妇，都可以前来，吃得饱足，好让耶和华－你的上帝在你手里所做的一切事上赐福给你。”
DEUT|15|1|“每七年的最后一年，你要施行豁免。
DEUT|15|2|豁免的方式是这样：凡债主要把手里所借给邻舍的全豁免，不可向邻舍和弟兄追讨，因为耶和华的豁免已经宣告了。
DEUT|15|3|你可以向外邦人追讨；但你弟兄欠你的，无论是什么，你都要放手豁免。
DEUT|15|4|其实，在你中间不会有贫穷人；因为在耶和华－你上帝所赐你为业的地上，耶和华必大大赐福给你。
DEUT|15|5|只要你留心听从耶和华－你上帝的话，谨守遵行我今日所吩咐你这一切的命令，
DEUT|15|6|因为耶和华－你的上帝会照他所应许你的赐福给你，你必借给许多国家，却不需要去借贷；你要管辖许多国家，它们却不能管辖你。
DEUT|15|7|“在耶和华－你上帝所赐给你的地上，任何一座城里，你弟兄中若有一个贫穷人，你不可硬着心，袖手不帮助你贫穷的弟兄。
DEUT|15|8|你总要伸手帮助他，照他所缺乏的借给他，补他的不足。
DEUT|15|9|你要谨慎，不可心起恶念，说：‘第七年的豁免年快到了’，你就冷眼看你贫穷的弟兄，什么都不给他。他若为你的缘故求告耶和华，你就有罪了。
DEUT|15|10|你要慷慨解囊，给他的时候不要心疼，因为耶和华－你的上帝必为这事，在你一切的工作上和你手所做的一切赐福给你。
DEUT|15|11|因为地上的贫穷人永远不会断绝，所以我吩咐你说：‘总要伸手帮助你地上困苦贫穷的弟兄。’”
DEUT|15|12|“你弟兄中，若有一个 希伯来 男人或 希伯来 女人卖给你，已服事你六年，到了第七年就要让他自由离开你。
DEUT|15|13|你让他自由离开的时候，不可让他空手而去，
DEUT|15|14|要从你的羊群、禾场、压酒池中取一些，慷慨地送给他；耶和华－你的上帝怎样赐福给你，你也要照样给他。
DEUT|15|15|要记得你在 埃及 地作过奴仆，耶和华－你的上帝救赎了你。为此，我今日将这事吩咐你。
DEUT|15|16|他若对你说：‘我不愿意离开你’，因为他爱你和你的家，并且他在你那里很好，
DEUT|15|17|你要拿锥子在门上穿透他的耳朵，他就永远成为你的奴仆了。你待婢女也要这样。
DEUT|15|18|你让他从你那里自由离开的时候，不要看作困难，因为他已服事你六年，相当于雇工双倍的工钱。这样，耶和华－你的上帝必在你所做的一切事上赐福给你。”
DEUT|15|19|“你牛群羊群中头生的，凡是公的，都要分别为圣，归给耶和华－你的上帝。头生的牛，不可用它来耕作；头生的羊，不可剪它的毛。
DEUT|15|20|这头生的，你和你全家每年要到耶和华所选择的地方，在耶和华－你上帝面前吃。
DEUT|15|21|这头生的若有残疾，瘸腿的或瞎眼的，若有任何严重缺陷，都不可献给耶和华－你的上帝。
DEUT|15|22|你们可以在城里吃，洁净的人和不洁净的人都可以吃，就如吃羚羊和鹿一样。
DEUT|15|23|只是它的血，你不可吃，要倒在地上，如同倒水一样。”
DEUT|16|1|“你要守亚笔月，向耶和华－你的上帝守逾越节，因为在亚笔月，耶和华－你的上帝在夜间领你出 埃及 。
DEUT|16|2|你当在那里，耶和华选择作为他名居所的地方，从羊群牛群中，将逾越节的祭牲献给耶和华－你的上帝。
DEUT|16|3|这祭牲不可和有酵的东西一起吃。因为你曾匆忙离开 埃及 地，你要吃无酵饼，就是困苦饼七日，好让你一生的年日记得你从 埃及 地出来的那一日。
DEUT|16|4|在你全境内，七日不可见到酵母。第一日晚上所献的肉，一点也不可留到早晨。
DEUT|16|5|你不可在耶和华－你上帝所赐的各城中，任何一座城里，献逾越节的祭，
DEUT|16|6|只可在那里，耶和华－你上帝选择作为他名居所的地方，在晚上日落的时候，就是你出 埃及 的时候，献逾越节的祭。
DEUT|16|7|你要在耶和华－你上帝所选择的地方把肉烤来吃，次日早晨就回到你的帐棚去。
DEUT|16|8|你要吃无酵饼六日，第七日要向耶和华－你的上帝守严肃会，不可做工。”
DEUT|16|9|“你要计算七个七日：从你用镰刀开始收割庄稼时算起，一共七个七日。
DEUT|16|10|你要向耶和华－你的上帝守七七节，按照耶和华－你上帝所赐你的福，献上你手里的甘心祭。
DEUT|16|11|你和你的儿女、仆婢，以及住在你城里的 利未 人、在你中间寄居的和孤儿寡妇，都要在那里，耶和华－你上帝选择作为他名居所的地方，在耶和华－你上帝面前欢乐。
DEUT|16|12|你要记得你在 埃及 作过奴仆，也要谨守遵行这些律例。”
DEUT|16|13|“你收藏了禾场和压酒池的出产以后，就要守住棚节七日。
DEUT|16|14|在节期中，你和你的儿女、仆婢，以及住在你城里的 利未 人、寄居的和孤儿寡妇，都要欢乐。
DEUT|16|15|在耶和华所选择的地方，你要向耶和华－你的上帝守节七日，因为耶和华－你的上帝要在你一切的收成上和你手里所做的一切赐福给你，你就非常欢乐。
DEUT|16|16|“你所有的男丁要在除酵节、七七节、住棚节，一年三次，在耶和华－你上帝所选择的地方朝见他，不可空手朝见耶和华。
DEUT|16|17|各人要按自己手中的能力，照耶和华－你上帝所赐你的福，奉献礼物。”
DEUT|16|18|“你要在耶和华－你上帝所赐的各城中，为各支派设立审判官和官长。他们要按公义的判断审判百姓，
DEUT|16|19|不可屈枉正直，不可看人的情面，也不可接受贿赂，因为贿赂能使智慧人的眼睛变瞎，又能曲解义人的证词。
DEUT|16|20|公正！你要追求公正，好使你存活，承受耶和华－你上帝所赐你的地。”
DEUT|16|21|“你为耶和华－你的上帝筑坛，不可在坛旁栽种任何树木作 亚舍拉 ，
DEUT|16|22|也不可为自己设立柱像，这是耶和华－你的上帝所憎恨的。”
DEUT|17|1|“凡有残疾，有任何恶疾的牛羊，你都不可献给耶和华－你的上帝，因为这是耶和华－你上帝所憎恶的。
DEUT|17|2|“在你中间，在耶和华－你上帝所赐你的各城中，任何一座城里，若有男人或女人做了耶和华－你上帝眼中看为恶的事，违背了他的约，
DEUT|17|3|去事奉别神，敬拜它们，或拜太阳，或拜月亮，或拜天上的万象，是我 不曾吩咐的。
DEUT|17|4|有人告诉你，你也听见了，就要细心探听。看哪，是真的，确实有这可憎的事在 以色列 中发生，
DEUT|17|5|你就要将行这恶事的男人或女人拉到城门外，用石头把这男人或女人处死。
DEUT|17|6|要凭两个证人或三个证人的口，才可以把他处死，不可只凭一个证人的口处死他。
DEUT|17|7|证人要先动手，然后众百姓也动手把他处死。这样，你就把恶从你中间除掉。
DEUT|17|8|“你城中若有难以判断的案件，涉及流血，诉讼，或殴打等争讼的事，你就要起来，上到那里，耶和华－你上帝所选择的地方，
DEUT|17|9|去见 利未 家的祭司和当时的审判官，求问他们，他们必将判决指示你。
DEUT|17|10|他们在耶和华所选择的地方指示你的判决，你要执行，谨守遵行他们一切所教导你的。
DEUT|17|11|要按照所教导你的律法、所告诉你的典章去执行；他们指示你的判决，你不可偏离左右。
DEUT|17|12|若有人擅自行事，不听从那侍立在耶和华－你上帝那里事奉的祭司，或不听从审判官，那人就要处死。这样，你就把恶从 以色列 中除掉。
DEUT|17|13|众百姓听见了都要害怕，不再擅自行事了。”
DEUT|17|14|“你到了耶和华－你上帝所赐你的地，得了那地居住在其中的时候，若说：‘我要立王治理我，像我四围所有的国家一样’，
DEUT|17|15|你一定要立耶和华－你上帝所拣选的人为你的王。要从你弟兄中立一人为你的王，不可立你弟兄之外的外邦人治理你。
DEUT|17|16|只是王不可为自己加添马匹，也不可为加添马匹使百姓回 埃及 去，因耶和华曾对你们说：‘不可再回那条路去。’
DEUT|17|17|王不可为自己多立妃嫔，免得他的心偏离；也不可为自己多积金银。
DEUT|17|18|他登了国度的王位之后，要在 利未 家的祭司面前，将这律法书为自己抄写一份在书卷上。
DEUT|17|19|这书要存在他那里，他一生的年日要诵读，好使他学习敬畏耶和华－他的上帝，谨守遵行这律法书上的一切话和这些律例，
DEUT|17|20|免得他的心向弟兄高傲，偏离了这诫命，或向右或向左。这样，他和他的子孙就可以长久作王治理 以色列 。”
DEUT|18|1|“ 利未 家的祭司和 利未 全支派在 以色列 中没有分得产业；他们可以吃耶和华的火祭，那是他的产业。
DEUT|18|2|他在弟兄中没有产业；耶和华是他的产业，正如耶和华所应许他的。
DEUT|18|3|祭司从百姓当得的权益是这样：凡献牛或羊为祭物的，要把前腿、两腮和胃给祭司。
DEUT|18|4|初收的五谷、新酒和新的油，以及初剪的羊毛，也要给他。
DEUT|18|5|因为耶和华－你的上帝从你众支派中拣选他，使他和他子孙永远奉耶和华的名侍立，事奉。
DEUT|18|6|“ 利未 人若离开他在 以色列 中所居住的任何一座城，一心愿意到耶和华所选择的地方，
DEUT|18|7|就要在那里奉耶和华－他上帝的名事奉，正如他的众弟兄 利未 人在耶和华面前侍立一样。
DEUT|18|8|除了卖祖产所得的以外，他们 要吃同等分量的祭物。”
DEUT|18|9|“你到了耶和华－你上帝所赐你之地，不可学那些国家行可憎恶的事。
DEUT|18|10|你中间不可有人使儿女经火，也不可有占卜的、观星象的、行法术的 、行邪术的、
DEUT|18|11|施符咒的、招魂的、行巫术的和求问死人的。
DEUT|18|12|凡做这些事的都是耶和华所憎恶的；因这可憎恶的事，耶和华－你的上帝把他们从你面前赶出去。
DEUT|18|13|你要向耶和华－你的上帝作完全人。
DEUT|18|14|你所要赶出的那些国家都听从观星象的和占卜的，但是耶和华－你的上帝从来不准你这样做。”
DEUT|18|15|“耶和华－你的上帝要从你弟兄中给你兴起一位先知像我，你们要听他。
DEUT|18|16|这正如你在 何烈山 大会的那日向耶和华－你的上帝所求的一切，说：‘求你不要再叫我听见耶和华－我上帝的声音，也不要再叫我看见这大火，免得我死亡。’
DEUT|18|17|耶和华对我说：‘他们说得对。
DEUT|18|18|我必在他们弟兄中给他们兴起一位先知像你。我要将当说的话放在他口里；他要将我一切所吩咐的都告诉他们。
DEUT|18|19|谁不听从他奉我名所说的话，我必亲自向他追究。
DEUT|18|20|若有先知擅自奉我的名说了我未曾吩咐他说的话，或是奉别神的名说话，那先知就必处死。’
DEUT|18|21|你心里若说：‘我们怎能知道那话是耶和华未曾吩咐的呢？’
DEUT|18|22|先知奉耶和华的名说话，所说的若没有实现，或不应验，这话就是耶和华未曾吩咐的，而是那先知擅自说的，你不必怕他。”
DEUT|19|1|“耶和华－你的上帝将列国剪除，他们的地耶和华－你上帝已赐给你，你又赶出他们，并且住在他们的城镇和房屋，
DEUT|19|2|那时，你要在耶和华－你上帝所赐你为业的地上，为自己指定三座城。
DEUT|19|3|你要预备道路，将耶和华－你上帝使你承受为业的地分为三区，使任何一个杀人的可以逃到那里去。
DEUT|19|4|“杀人的逃到那里得以存活的案例是这样：凡素无仇恨，无意中杀了邻舍的，
DEUT|19|5|就如人与邻舍同入林中伐木，手拿斧子一砍，本想砍下树木，斧头却脱了把，飞落在邻舍身上，以致那人死去，这人就可以逃到那些城中的一座，得以存活，
DEUT|19|6|免得报血仇的心中发火，去追赶那杀了人的，因为路途遥远就能追上他，把他杀死。其实他是不该死的，因为他与被杀者素无仇恨。
DEUT|19|7|所以我吩咐你说，要为自己指定三座城。
DEUT|19|8|耶和华－你的上帝若照他向你列祖所起的誓扩张你的疆土，将所应许赐你列祖的全地给你，
DEUT|19|9|你若谨守遵行我今日所吩咐的这一切诫命，爱耶和华－你的上帝，天天遵行他的道，就要在这三座城之外，再添三座城，
DEUT|19|10|免得无辜人的血流在耶和华－你上帝所赐你为业的地中间，血就归到你身上了。
DEUT|19|11|“若有人恨他的邻舍，埋伏等着，起来击杀他，把他杀死，然后逃到这些城中的一座，
DEUT|19|12|他本城的长老就要派人去，从那里把他带出来，交在报血仇者的手中，把他处死。
DEUT|19|13|你的眼不可顾惜他，要从 以色列 中除掉流无辜血的罪，使你得福。”
DEUT|19|14|“在耶和华－你上帝所赐你承受为业，所分得的地上，不可挪移你邻舍的地界，因为这是前人所定的。”
DEUT|19|15|“人无论犯什么罪，作什么恶，不可单凭一个人的见证，总要凭两个证人的口或三个证人的口才可定案。
DEUT|19|16|若有人怀恶意，起来作证，控告他人犯法，
DEUT|19|17|这两个争讼的人就要站在耶和华面前，和当时的祭司与审判官面前，
DEUT|19|18|审判官要细心调查。看哪，证人作的是伪证，要用伪证陷害弟兄，
DEUT|19|19|你们就要对付他如同他想要对付的弟兄一样。这样，你就把恶从你中间除掉。
DEUT|19|20|其他的人听见就害怕，不敢在你中间再行这样的恶事了。
DEUT|19|21|你的眼不可顾惜，要以命偿命，以眼还眼，以牙还牙，以手还手，以脚还脚。”
DEUT|20|1|“你出去与仇敌作战，若看见马匹、战车，以及比你更多的士兵，不要怕他们，因为领你出 埃及 地的耶和华－你的上帝与你同在。
DEUT|20|2|你们将要上阵的时候，祭司要来，向士兵宣告，
DEUT|20|3|对他们说：‘ 以色列 啊，要听！你们今日将要与仇敌作战，不要心惊胆战，不要惧怕战兢，也不要因他们惊慌，
DEUT|20|4|因为与你们同去的是耶和华－你们的上帝，他要为你们与仇敌作战，拯救你们。’
DEUT|20|5|官长也要向士兵宣告说：‘谁建了新的房屋尚未奉献，他可以回家去，免得他阵亡，别人去奉献。
DEUT|20|6|谁栽植了葡萄园尚未享用所结的果子，他可以回家去，免得他阵亡，别人去享用。
DEUT|20|7|谁与女子订了婚尚未迎娶，他可以回家去，免得他阵亡，别人去娶。’
DEUT|20|8|官长要继续对士兵说：‘谁惧怕，心惊胆战，可以回家去，免得他弟兄的心像他的心一样消沉。’
DEUT|20|9|官长向士兵宣告完毕，军官就率领士兵去了。
DEUT|20|10|“你来到一座城，要攻城之前，先向它宣告和平。
DEUT|20|11|那城若愿意以和平回应，给你开城，城里所有的人就要为你做苦工，服事你。
DEUT|20|12|若那城拒绝和平，却要与你打仗，你就要围困那城。
DEUT|20|13|耶和华－你的上帝把那城交在你手里时，你就要用刀杀尽城里的男丁。
DEUT|20|14|至于妇女、孩童、牲畜和城里所有的，你都可以取为自己的掠物。从仇敌所掠夺的，就是耶和华－你上帝所赐给你的，你都可以享用。
DEUT|20|15|离你很远的各城，就是不属于这些国家的城镇，你都要这样对待他们。
DEUT|20|16|但是这些民族的城镇，就是耶和华－你上帝所赐给你的产业，其中凡有气息的，一个都不可存留。
DEUT|20|17|你要照耶和华－你上帝所吩咐的，将这些 赫 人、 亚摩利 人、 迦南 人、 比利洗 人、 希未 人、 耶布斯 人全都灭绝，
DEUT|20|18|免得他们教导你们去行一切可憎恶的事，就是他们向自己神明所行的，使你们得罪耶和华－你们的上帝。
DEUT|20|19|“你若围困一座城，需要攻打许多日子才能夺取，就不可用斧头砍坏树木。你可以吃树上的果子，却不可把树砍下来。田间的树木岂是人，让你去围攻的吗？
DEUT|20|20|只有那些你知道不能生产食物的树才可以毁坏；你可以把它们砍下来造攻城的工具，攻打那与你打仗的城，直到把城攻下。”
DEUT|21|1|“在耶和华－你上帝所赐你为业的地上，若发现有人被杀，暴尸野地，不知道是谁杀的，
DEUT|21|2|长老和审判官 就要出去，从尸体那里量起，量到四围的城镇，
DEUT|21|3|看哪一座城最靠近这尸体，那城的几位长老就要取一头未曾耕地、未曾负轭的母牛犊；
DEUT|21|4|那城的长老要把这母牛犊牵到流着溪水、未曾耕耘、未曾撒种的山谷去，在谷中打断它的颈项。
DEUT|21|5|利未 人祭司要近前来，因为耶和华－你的上帝拣选他们来事奉他，奉耶和华的名祝福，并且有任何的争讼和殴打，都由他们的口判决。
DEUT|21|6|离尸体最近的那座城的每位长老要在山谷中，在颈项被打断的母牛犊上面洗手，
DEUT|21|7|声明说：‘我们的手未曾流这人的血；我们的眼也未曾看见这事。
DEUT|21|8|耶和华啊，求你赦免你所救赎的百姓 以色列 ，不要让无辜的血归在你的百姓 以色列 中间。’这样，他们流血的罪就必得赦免。
DEUT|21|9|你行了耶和华眼中看为正的事，就可以从你中间除掉无辜的血。”
DEUT|21|10|“你出去与仇敌作战的时候，耶和华－你的上帝将他交在你手中，你就掳了他为俘虏。
DEUT|21|11|若你在被掳的人中看见美丽的女子，喜欢她，要娶她为妻，
DEUT|21|12|就可以带她到你家去。她要剪头发，修指甲，
DEUT|21|13|脱去被掳时所穿的衣服，住在你家里为自己父母哀哭一个月。然后，你就可以与她同房；你作她的丈夫，她作你的妻子。
DEUT|21|14|以后你若不喜欢她，就要让她自由离开，绝不可为钱把她卖了，也不可把她当奴隶看待，因为你已经占有过她。”
DEUT|21|15|“人若有两个妻子，一个是他宠爱的，另一个是失宠的 ，她们都给他生了儿子，但长子是他失宠妻子生的；
DEUT|21|16|到了分产业给儿子的时候，不可将自己宠爱的妻子所生的儿子立为长子，在他失宠妻子所生的长子之上。
DEUT|21|17|他必须认失宠妻子所生的儿子为长子，在所有的产业中给他双分，因为这儿子是他壮年时生的，长子的名分应当是他的。”
DEUT|21|18|“人若有顽梗忤逆的儿子，不听从父母的话，他们虽然惩戒他，他还是不听从他们，
DEUT|21|19|父母就要抓住他，带他出去到当地的城门，本城的长老那里，
DEUT|21|20|对本城的长老说：‘我们这个儿子顽梗忤逆，不听从我们的话，是贪食好酒的人。’
DEUT|21|21|然后，城里的众人就要用石头将他打死。这样，你就把恶从你中间除掉，全 以色列 听见了都要害怕。”
DEUT|21|22|“人若犯了死罪被处死，你把他挂在木头上，
DEUT|21|23|不可让尸体留在木头上过夜，一定要当日把他埋葬，因为被挂的人是上帝所诅咒的。你不可玷污耶和华－你上帝所赐你为业的地。”
DEUT|22|1|“你若看见弟兄的牛或羊迷了路，不可避开它们，总要把它们牵回来交给你的弟兄。
DEUT|22|2|你弟兄若离你远，或是你不认识他，你就要牵到你家，留在你那里，等你的弟兄来寻找就还给他。
DEUT|22|3|你弟兄所失落的，无论是驴，衣服，或任何东西，你若发现，都要这样做，不能避开。
DEUT|22|4|你若看见你弟兄的牛或驴在路上跌倒了，不可避开它们，总要帮助他把牛或驴拉起来。
DEUT|22|5|“妇女不可穿戴男子所穿戴的，男人也不可穿妇女的衣服，因为这样做是耶和华－你上帝所憎恶的。
DEUT|22|6|“你若路上看见鸟窝，无论在树上或地上，里头有小鸟或有蛋，母鸟伏在小鸟或蛋上，你不可连母鸟带小鸟一起拿去。
DEUT|22|7|总要放母鸟走，只可以取小鸟。这样你就可以享福，日子得以长久。
DEUT|22|8|“你若建造新房屋，要在屋顶安栏杆，免得有人从屋顶掉下来，血就归于你家。
DEUT|22|9|“不可在你的葡萄园里栽种别的种子，免得你栽种所结的和葡萄园的果子都成了圣物。
DEUT|22|10|不可并用牛和驴来耕地。
DEUT|22|11|不可穿羊毛和细麻混合做成的衣服。
DEUT|22|12|“你要在所披外衣的四个边上缝繸子。”
DEUT|22|13|“人若娶妻，与她同房后恨恶她，
DEUT|22|14|捏造她行可耻的事，把丑名加在她身上，说：‘我娶了这女人，亲近她，却发现她没有贞洁的凭据’。
DEUT|22|15|女方的父母就要把这女子贞洁的凭据拿出去，到城门的本城长老那里。
DEUT|22|16|女方的父亲要对长老说：‘我把女儿嫁给这人，他却恨恶她，
DEUT|22|17|看哪，他捏造可耻的事，说：我发现你女儿没有贞洁的凭据。但是，这就是我女儿贞洁的凭据。’父母要把那布铺在本城长老的面前。
DEUT|22|18|那城的长老要拿住那人，惩罚他，
DEUT|22|19|罚他一百银子，给女方的父亲，因为他把丑名加在 以色列 一个少女身上。这女子仍是他的妻子，那人终身不可休她。
DEUT|22|20|但若这事是真的，找不到女子贞洁的凭据，
DEUT|22|21|他们就要把这女子带到她父家的门口，城里的人要用石头打死她，因为她在父家犯了淫乱，在 以色列 中做了可耻的事。这样，你就把恶从你中间除掉。
DEUT|22|22|“若发现有人与有夫之妇同寝，就要将奸夫淫妇一起处死。这样，你就把恶从 以色列 中除掉。
DEUT|22|23|“若一女子是处女，已经许配了人，有男子在城里遇见她，与她同寝，
DEUT|22|24|你们就要把这二人带到那城的城门口，用石头打死他们。处死女子是因为她虽然在城里， 却没有喊叫；处死男子是因为他玷污了邻舍的妻子。这样，你就把恶从你中间除掉。
DEUT|22|25|“若有男子在野地遇见已经许配人的女子，抓住她与她同寝，只要处死那与女子同寝的男子。
DEUT|22|26|不可对女子处刑，这女子没有该死的罪。这案件就好比人起来攻击邻舍，把他杀了一样。
DEUT|22|27|因为男子是在野地遇见她，这已经许配了人的女子虽然喊叫，却没有人救她。
DEUT|22|28|“若有男子遇见没有许配人的少女，抓住她与她同寝，被人发现，
DEUT|22|29|这男子就要拿五十银子给女子的父亲，并要娶她为妻，终身不可休她，因为他玷污了这女子。
DEUT|22|30|“人不可娶继母为妻，不可掀开父亲衣服的下边 。”
DEUT|23|1|“凡外肾损伤的，或被阉割的，不可入耶和华的会。
DEUT|23|2|“私生子不可入耶和华的会；甚至到第十代，也不可入耶和华的会。
DEUT|23|3|“ 亚扪 人或 摩押 人不可入耶和华的会；甚至到第十代，也永不可入耶和华的会。
DEUT|23|4|因为你们出 埃及 的时候，他们没有拿食物和水在路上迎接你们，并且雇了 美索不达米亚 的 毗夺 人， 比珥 的儿子 巴兰 来诅咒你。
DEUT|23|5|然而耶和华－你的上帝不愿听 巴兰 ，耶和华－你的上帝为你使诅咒变为祝福，因为耶和华－你的上帝爱你。
DEUT|23|6|你一生一世永不可为他们求平安和福气。
DEUT|23|7|“不可憎恶 以东 人，因为他是你的弟兄。不可憎恶 埃及 人，因为你曾在他的地上作过寄居的。
DEUT|23|8|他们所生的第三代子孙可以入耶和华的会。”
DEUT|23|9|“你出兵攻打敌人，要远离一切恶事。
DEUT|23|10|“你中间若有人因夜间梦遗而不洁净，就要出到营外，不可入营。
DEUT|23|11|到了傍晚，他要用水洗澡，等到日落才可以入营。
DEUT|23|12|“你要在营外划定一个地方，你可以出去在那里方便。
DEUT|23|13|在你器械中当有一把锹；你出营外便溺以后，要用它挖洞，转身掩盖排泄物。
DEUT|23|14|因为耶和华－你的上帝在你营中走动，要拯救你，将仇敌交给你，所以你的营应当圣洁，免得他见你那里有污秽之物就转身离开你。”
DEUT|23|15|“你不可把从主人身边逃到你那里的奴仆，交回给他的主人，
DEUT|23|16|要让他在你那里与你同住，由他在你的城镇中选择一个自己喜欢的地方居住，不可欺负他。
DEUT|23|17|“ 以色列 的女子中不可作神庙娼妓； 以色列 的男子中也不可作神庙娼妓。
DEUT|23|18|妓女和男娼 的赏金，都不可带进耶和华－你上帝的殿中还愿，因为两者都是耶和华－你上帝所憎恶的。
DEUT|23|19|“你借给你弟兄的，无论是钱财是粮食，或任何可生利息的财物，都不可取利。
DEUT|23|20|借给外邦人可以取利，但借给你的弟兄就不可取利；好让耶和华－你的上帝在你去得为业的地上和你手里所做的一切，赐福给你。
DEUT|23|21|“你向耶和华－你的上帝许愿，不可迟延还愿，因为耶和华－你的上帝必定向你追讨，你就有罪了。
DEUT|23|22|你若不许愿，倒没有罪。
DEUT|23|23|你嘴唇所说的，你亲口承诺的，要照你甘心向耶和华－你上帝许的愿谨守遵行。
DEUT|23|24|“你进入邻舍的葡萄园，可以随意吃葡萄，直到饱足，却不可装在器皿中。
DEUT|23|25|你进入邻舍的庄稼中，可以用手摘麦穗，却不可用镰刀割取庄稼。”
DEUT|24|1|“人若娶妻，作了她的丈夫，发现她有不合宜的事不喜欢她，而写休书交在她手中，打发她离开夫家，
DEUT|24|2|妇人若离开夫家以后，去嫁别人，
DEUT|24|3|后夫若恨恶她，写休书交在她手中，打发她离开夫家，又或者娶她为妻的后夫死了，
DEUT|24|4|那休她的前夫就不可在妇人玷污之后再娶她为妻，因为这是耶和华所憎恶的。不可使耶和华－你上帝所赐为业之地蒙受玷污。
DEUT|24|5|“人若娶了新娘，不可从军出征，也不可派他办理任何事情。他可以在家清闲一年，使他所娶的妻快活。
DEUT|24|6|“不可拿人的石磨或上面的磨石作抵押，因为这是拿人的命作抵押。
DEUT|24|7|“若发现有人绑架 以色列 人中的一个弟兄，把他当奴隶对待，或把他卖了，那绑架人的就必处死。这样，你就把恶从你中间除掉。
DEUT|24|8|“关于痲疯 的灾病，你们要谨慎，照 利未 家的祭司一切所指教你们的留心遵行。我怎样吩咐他们，你们要照样遵行。
DEUT|24|9|要记得，在你们出 埃及 后的路途中，耶和华－你的上帝向 米利暗 所做的事。
DEUT|24|10|“你借给邻舍，无论是什么，不可进他家拿抵押品。
DEUT|24|11|要站在外面，等那借贷的人把抵押品拿出来交给你。
DEUT|24|12|他若是困苦的人，你不可用他的抵押品盖着睡觉。
DEUT|24|13|日落的时候，总要把抵押品还给他，让他用那件外衣盖着睡觉，他就为你祝福。这在耶和华－你的上帝面前就是你的义行了。
DEUT|24|14|“困苦贫穷的雇工，无论是你的弟兄，或是住在你境内，在你城里寄居的，你都不可欺负他 。
DEUT|24|15|要当日给他工钱，不可等到日落，因为他困苦，需要靠工钱过活，免得他因你的缘故求告耶和华，罪就归于你了。
DEUT|24|16|“不可因儿子处死父亲，也不可因父亲处死儿子；各人要因自己的罪被处死。
DEUT|24|17|“不可对寄居的和孤儿屈枉正直，也不可拿寡妇的衣服作抵押。
DEUT|24|18|要记得你曾在 埃及 作过奴仆，耶和华－你的上帝从那里救赎了你，所以我吩咐你遵行这事。
DEUT|24|19|“你在田间收割庄稼，若忘了一捆在田间，就不要再回去拿，要留给寄居的、孤儿和寡妇；好让耶和华－你的上帝在你手里所做的一切，赐福给你。
DEUT|24|20|你打了橄榄树，枝上剩下的不可再打，要留给寄居的、孤儿和寡妇。
DEUT|24|21|你摘葡萄园的葡萄，掉落的不可拾取，要留给寄居的、孤儿和寡妇。
DEUT|24|22|你要记得你曾在 埃及 地作过奴仆，所以我吩咐你遵行这事。
DEUT|25|1|“人与人若有争讼，要求审判，当宣判义人为义，恶人有罪的时候，
DEUT|25|2|恶人若该受责打，审判官就要叫他当着面，伏在地上，按他的罪照数责打。
DEUT|25|3|只能打四十下，不可加多；多过这数目就是在你眼中作贱你的弟兄了。
DEUT|25|4|“牛在踹谷的时候，不可笼住它的嘴。”
DEUT|25|5|“兄弟住在一起，若其中一个死了，没有儿子，死者的妻子就不可出去嫁给陌生人。她丈夫的兄弟应当尽兄弟的本分，娶她为妻，与她同房。
DEUT|25|6|妇人生的长子要归在已故兄弟的名下，免得他的名在 以色列 中涂去了。
DEUT|25|7|那人若不情愿娶他兄弟的妻子，他兄弟的妻子就要上到城门长老那里，说：‘我丈夫的兄弟拒绝在 以色列 中为他的兄弟留名，不愿意为我尽兄弟的本分。’
DEUT|25|8|本城的长老就要召那人来，跟他谈话。若他坚持说：‘我不情愿娶她。’
DEUT|25|9|他兄弟的妻子就要在长老眼前来到那人跟前，脱下他脚上的鞋，吐唾沫在他脸上，回应说：‘凡不为兄弟建立家室的都要这样待他。’
DEUT|25|10|在 以色列 中，他要以‘脱鞋之家’闻名。”
DEUT|25|11|“若有人和弟兄争斗，其中一人的妻子近前去，为了救丈夫脱离那打丈夫之人的手，伸手抓住那人的下体，
DEUT|25|12|你就要砍断妇人的手，你的眼不可顾惜。
DEUT|25|13|“你袋中不可有一大一小两样的法码。
DEUT|25|14|你家里不可有一大一小两样的伊法 。
DEUT|25|15|当用准确公正的法码和伊法，好使你的日子在耶和华－你上帝所赐你的地上得以长久。
DEUT|25|16|因为行这一切不义之事的人都是耶和华－你上帝所憎恶的。”
DEUT|25|17|“你要记得你们出 埃及 的时候， 亚玛力 在路上怎样对待你，
DEUT|25|18|在路上迎击你，趁你疲乏困倦时击杀所有在你后面软弱的人；并不敬畏上帝。
DEUT|25|19|所以，当耶和华－你的上帝使你不被四围一切仇敌扰乱，在耶和华－你上帝赐你为业的地上得享平静的时候，你要把 亚玛力 的名从天下涂去；你不可忘记这事。”
DEUT|26|1|“你进去得了耶和华－你上帝所赐你为业的地，并且居住在那里的时候，
DEUT|26|2|就要从耶和华－你上帝所赐你的地上，将收成的各种初熟土产取一些来，盛在筐子里，带到那里，耶和华－你上帝选择作为他名居所的地方，
DEUT|26|3|到当时的祭司那里，对他说：‘我今日向耶和华－你的上帝宣认，我已来到耶和华向我们列祖起誓要赐给我们的地。’
DEUT|26|4|祭司就从你手里把筐子接过来，供在耶和华－你上帝的祭坛前。
DEUT|26|5|你要在耶和华－你上帝面前告白说：‘我的祖先原是一个流亡的 亚兰 人，带着稀少的人丁下到 埃及 寄居。在那里，他却成了又大又强、人数众多的国。
DEUT|26|6|埃及 人恶待我们，迫害我们，将苦工加在我们身上。
DEUT|26|7|于是我们哀求耶和华我们列祖的上帝。耶和华听见我们的声音，看见我们所受的困苦、劳役和欺压，
DEUT|26|8|耶和华就用大能的手和伸出来的膀臂，以及大而可畏的事和神迹奇事，领我们出了 埃及 ，
DEUT|26|9|将我们领进这地方，把这流奶与蜜之地赐给我们。
DEUT|26|10|耶和华啊，看哪，现在我把你所赐我地上初熟的土产供上。’随后你要把筐子供在耶和华－你上帝面前，向耶和华－你的上帝下拜。
DEUT|26|11|你和 利未 人，以及在你中间寄居的，要因耶和华－你上帝所赐你和你家的一切福分欢乐。
DEUT|26|12|“每逢第三年，就是捐十分之一的那年，你从你一切土产中取了十分之一，要分给 利未 人、寄居的、孤儿和寡妇，使他们在你的城镇中可以吃得饱足。
DEUT|26|13|你又要在耶和华－你上帝面前说：‘我已将圣物从家里拿出来，给了 利未 人、寄居的、孤儿和寡妇，是遵照你吩咐我的一切命令。你的命令，我没有违背，也没有忘记。
DEUT|26|14|我守丧的时候，没有吃这圣物，不洁净的时候，也没有拿出来，又没有把它献给死人。我听从了耶和华－我上帝的话，都照你一切所吩咐的做了。
DEUT|26|15|求你从天上，从你的圣所垂看，赐福给你的百姓 以色列 和你向我们列祖起誓所赐给我们的这片土地，就是流奶与蜜之地。’”
DEUT|26|16|“耶和华－你的上帝今日吩咐你遵行这些律例典章，所以你要尽心尽性谨守遵行。
DEUT|26|17|你今日宣认耶和华为你的上帝，承诺遵行他的道，谨守他的律例、诫命、典章，听从他的话。
DEUT|26|18|耶和华今日照他所应许你的，也认你为他宝贵的子民，叫你谨守他的一切诫命，
DEUT|26|19|要使你得称赞、美名、尊荣，超乎他所造的万国之上，并且照他所应许的，使你归耶和华－你的上帝为神圣的子民。”
DEUT|27|1|摩西 和 以色列 的众长老吩咐百姓说：“你们要遵守我今日所吩咐的一切诫命。
DEUT|27|2|你们过了 约旦河 ，到耶和华－你上帝所赐给你的地，当日要竖立几块大石头，涂上石灰。
DEUT|27|3|当你过了河，进入耶和华－你上帝所赐给你流奶与蜜之地，正如耶和华－你列祖的上帝所应许你的，你要把这律法的一切话写在石头上。
DEUT|27|4|你们过了 约旦河 ，就要在 基利心山 上照我今日所吩咐的，把这些石头竖立起来，涂上石灰。
DEUT|27|5|你在那里要为耶和华－你的上帝筑一座石坛，却不可动用铁器在石头上。
DEUT|27|6|要用没有凿过的石头筑耶和华－你上帝的坛，在坛上将燔祭献给耶和华－你的上帝，
DEUT|27|7|又要献平安祭，在那里吃，在耶和华－你的上帝面前欢乐。
DEUT|27|8|你要将这律法的一切话清楚地写在石头上。”
DEUT|27|9|摩西 和 利未 家的祭司吩咐 以色列 众人说：“ 以色列 啊，你要静默倾听！你今日已成为耶和华－你上帝的子民了。
DEUT|27|10|你要听从耶和华－你上帝的话，遵行他的诫命律例，就是我今日所吩咐你的。”
DEUT|27|11|当日， 摩西 吩咐百姓说：
DEUT|27|12|“你们过了 约旦河 ， 西缅 、 利未 、 犹大 、 以萨迦 、 约瑟 和 便雅悯 等支派的人要站在 基利心山 上为百姓祝福。
DEUT|27|13|吕便 、 迦得 、 亚设 、 西布伦 、 但 和 拿弗他利 等支派的人要站在 以巴路山 上宣布诅咒。
DEUT|27|14|利未 人要大声对 以色列 众人说：
DEUT|27|15|“‘凡制造耶和华所憎恶的偶像，无论是雕刻的，是铸造的，就是工匠用手造的，或暗中设置的，这人必受诅咒！’众百姓要回应说：‘阿们！’
DEUT|27|16|“‘轻慢父母的，必受诅咒！’众百姓要说：‘阿们！’
DEUT|27|17|“‘挪移邻舍地界的，必受诅咒！’众百姓要说：‘阿们！’
DEUT|27|18|“‘引领瞎子走错路的，必受诅咒！’众百姓要说：‘阿们！’
DEUT|27|19|“‘对寄居的、孤儿和寡妇屈枉正直的，必受诅咒！’众百姓要说：‘阿们！’
DEUT|27|20|“‘与继母同寝的，必受诅咒！因为他掀开父亲衣服的下边。’众百姓要说：‘阿们！’
DEUT|27|21|“‘与兽交合的，必受诅咒！’众百姓要说：‘阿们！’
DEUT|27|22|“‘与同父异母，或同母异父的姊妹同寝的，必受诅咒！’众百姓要说：‘阿们！’
DEUT|27|23|“‘与岳母同寝的，必受诅咒！’众百姓要说：‘阿们！’
DEUT|27|24|“‘暗中击杀邻舍的，必受诅咒！’众百姓要说：‘阿们！’
DEUT|27|25|“‘受贿赂击杀人而流无辜之血的，必受诅咒！’众百姓要说：‘阿们！’
DEUT|27|26|“‘不坚守遵行这律法之话的，必受诅咒！’众百姓要说：‘阿们！’”
DEUT|28|1|“你若留心听从耶和华－你上帝的话，谨守遵行他的一切诫命，就是我今日所吩咐你的，他必使你超乎地上的万国之上。
DEUT|28|2|你若听从耶和华－你上帝的话，这一切的福气必临到你身上，追随你：
DEUT|28|3|你在城里必蒙福，在田间也必蒙福。
DEUT|28|4|你身所生的，你地所产的，你牲畜所生的，牛犊、羔羊，都必蒙福。
DEUT|28|5|你的筐子和你的揉面盆都必蒙福。
DEUT|28|6|你出也蒙福，入也蒙福。
DEUT|28|7|“耶和华必使那起来攻击你的仇敌在你面前溃败。他们从一条路来攻击你，必在你面前从七条路逃跑。
DEUT|28|8|在你仓房里，以及你手所做的一切，耶和华必发令赐福给你。耶和华－你上帝也必在所赐你的地上赐福给你。
DEUT|28|9|你若谨守耶和华－你上帝的诫命，遵行他的道，他必照他向你所起的誓立你为自己神圣的子民。
DEUT|28|10|地上的万民见你归在耶和华的名下，就必惧怕你。
DEUT|28|11|在耶和华向你列祖起誓应许赐你的土地上，他必使你身所生的，牲畜所生的，地所产的，都丰富有余。
DEUT|28|12|耶和华必为你敞开天上的宝库，按时降雨在你的地上。他必赐福你手里所做的一切。你必借给许多国家，却不必去借贷。
DEUT|28|13|你若听从耶和华－你上帝的诫命，就是我今日所吩咐你的，谨守遵行，耶和华就必使你作首不作尾，居上不居下，
DEUT|28|14|只要你不偏左右，不背离我今日所吩咐你的一切话，也不随从别神，事奉它们。”
DEUT|28|15|“你若不听从耶和华－你上帝的话，不谨守遵行他的一切诫命律例，就是我今日所吩咐你的，这一切的诅咒必临到你身上，追随你：
DEUT|28|16|你在城里必受诅咒，在田间也必受诅咒。
DEUT|28|17|你的筐子和你的揉面盆都必受诅咒。
DEUT|28|18|你身所生的，你地所产的，以及牛犊、羔羊，都必受诅咒。
DEUT|28|19|你出也受诅咒，入也受诅咒。
DEUT|28|20|耶和华因你作恶离弃他，必在你手里所做的一切，使诅咒、困扰、责罚临到你，直到你被除灭，直到你迅速灭亡。
DEUT|28|21|耶和华必使瘟疫紧贴着你，直到他把你从所进去得为业的地上灭绝。
DEUT|28|22|耶和华要用痨病、热病、发炎、高烧、刀剑 、焚风 和霉烂攻击你；这些要追赶你，直到你灭亡。
DEUT|28|23|你头上的天要变成铜，下面的地要化为铁。
DEUT|28|24|耶和华要使那降在你地上的雨变为灰尘，尘土从天落在你身上，直到你被除灭。
DEUT|28|25|“耶和华必使你在仇敌面前溃败。你从一条路去攻击他们，必从七条路逃跑。地上万国必因你而惊骇。
DEUT|28|26|你的尸首必给空中的飞鸟和地上的走兽作食物，却无人哄赶。
DEUT|28|27|耶和华必用 埃及 人的疮、溃疡、癣和疥攻击你，使你不得医治。
DEUT|28|28|耶和华必用癫狂、眼瞎、心惊攻击你。
DEUT|28|29|你必在午间摸索，好像盲人在黑暗中摸索。你的道路必不亨通，天天受人欺压、抢夺，无人搭救。
DEUT|28|30|你聘了妻子，别人必与她同寝；你建了房屋，却不得住在其内；你栽植了葡萄园，却不得享用所结的果子。
DEUT|28|31|你的牛在你眼前宰了，你吃不到它的肉；你的驴在你眼前被人抢夺，却讨不回来；你的羊被敌人拿走，无人帮助你。
DEUT|28|32|你的儿女被交给别国的民；你的眼目终日切望，甚至失明，你的手却无能为力。
DEUT|28|33|你地所产的和你劳力所得的，必被你所不认识的百姓吃尽。你天天只被欺负，受压制，
DEUT|28|34|甚至你因眼中所见的景象而疯狂。
DEUT|28|35|耶和华必攻击你，使你膝上腿上，从脚掌到头顶，都长满了毒疮，无法医治。
DEUT|28|36|“耶和华必将你和你所立统治你的王，领到你和你列祖不认识的国去；在那里你必事奉别神，就是木头和石头。
DEUT|28|37|你在耶和华赶你到的万民中，要令人惊骇，成为笑柄，被人讥诮。
DEUT|28|38|你撒在田里的种子虽多，收的却少，因为蝗虫把它吃光了。
DEUT|28|39|你栽植修整葡萄园，却没有酒喝，也不得储存，因为虫子把它吃了。
DEUT|28|40|你全境有橄榄树，却得不到油抹身，因为你的橄榄都掉光了。
DEUT|28|41|你生儿育女，却不属于你，因为他们必被掳去。
DEUT|28|42|你所有的树木和你地里的出产必被蝗虫吃尽了。
DEUT|28|43|在你中间寄居的必上升高过你，高而又高；你必下降，低而又低。
DEUT|28|44|他必借给你，你却不能借给他；他必作首，你必作尾。
DEUT|28|45|这一切的诅咒必临到你，追赶你，赶上你，直到把你除灭，因为你不听从耶和华－你上帝的话，不遵守他吩咐的诫命律例。
DEUT|28|46|这些诅咒必在你和你后裔身上成为神迹奇事，直到永远！
DEUT|28|47|因为你富裕的时候，不以欢喜快乐的心事奉耶和华－你的上帝，
DEUT|28|48|所以你必在饥饿、干渴、赤身、缺乏中事奉仇敌，那是耶和华派来攻击你的。他必把铁轭加在你的颈项上，直到把你除灭。
DEUT|28|49|耶和华要从远方、地极之处带一国来，如鹰飞来攻击你；这国的语言，你听不懂。
DEUT|28|50|这国的人面貌凶恶，不给长者面子，也不恩待年轻人。
DEUT|28|51|他们必吃你牲畜所生的和你土地所产的，直到你被除灭。你的五谷、新酒和新的油，以及牛犊、羔羊，他都不给你留下，直到使你灭亡。
DEUT|28|52|他们必在你的各城围困你，直到你在全地所倚靠、高大坚固的城墙都倒塌。他们必在耶和华－你上帝所赐给你全地的各城围困你。
DEUT|28|53|你在仇敌围困的窘迫中，必吃你本身所生的，就是耶和华－你上帝所赐给你的儿女之肉。
DEUT|28|54|你中间，连那温和文雅的人都必冷眼恶待自己的兄弟和怀中的妻子，以及他所剩下其余的儿女，
DEUT|28|55|不把所吃儿女的肉分一点给他们任何一个人，因为在被仇敌围困、陷入窘迫的各城中，他已经一无所剩了。
DEUT|28|56|你中间柔顺娇嫩的妇人，甚至因柔顺娇嫩脚不肯踏地的妇人，也必冷眼恶待她怀中的丈夫和自己的儿女。
DEUT|28|57|在被仇敌围困、陷入窘迫的城镇中，她因缺乏一切，就要暗中把从她两腿中间出来的胞衣和所生下的儿女吃了。
DEUT|28|58|“这书上所写律法的一切话，是叫你敬畏耶和华－你上帝尊荣可畏的名，你若不谨守遵行，
DEUT|28|59|耶和华就必将奇异的灾害，就是严重持久的灾害和长期难治的疾病，加在你和你后裔的身上。
DEUT|28|60|他必使你所畏惧、 埃及 一切的疾病临到你，紧贴着你，
DEUT|28|61|没有写在这律法书上的各样疾病、灾害，耶和华也必降在你身上，直到你被除灭。
DEUT|28|62|你们虽然曾像天上的星那样多，却因不听从耶和华－你上帝的话，所剩的人丁就稀少了。
DEUT|28|63|耶和华先前怎样喜爱善待你们，使你们增多，耶和华也要照样喜爱消灭你们，使你们灭绝。你们必从所要进去得为业的地上被拔除。
DEUT|28|64|耶和华必把你们分散在万民中，从地的这边到地的另一边，在那里你必事奉你和你列祖不认识的神明，就是木头和石头。
DEUT|28|65|在那些国中，你必得不到安宁，脚掌也没有安歇之处；耶和华却要使你在那里心中发颤，眼目失明，精神沮丧。
DEUT|28|66|你的一生悬空不安；你昼夜恐惧，生命没有保障。
DEUT|28|67|你因心中的恐惧，眼睛所见的景象，早晨必说：‘但愿现在是晚上！’晚上必说：‘但愿现在是早晨！’
DEUT|28|68|耶和华要用船把你送回 埃及 去，走那我曾告诉你不再看见的路；在那里你们必卖身给你的仇敌作奴婢，却没有人要买。”
DEUT|29|1|耶和华在 何烈山 与 以色列 人立约以外，这是耶和华在 摩押 地吩咐 摩西 与 以色列 人立约的话。
DEUT|29|2|摩西 召全 以色列 来，对他们说：“耶和华在 埃及 地，在你们眼前向法老和他众臣仆，以及他的全地所做的一切事，你们都看见了，
DEUT|29|3|就是你亲眼看见的大考验，那些神迹和大奇事。
DEUT|29|4|但耶和华到今日还没有使你们心能明白，眼能看见，耳能听见。
DEUT|29|5|我领你们在旷野四十年，你们身上的衣服没有穿破，脚上的鞋也没有穿坏；
DEUT|29|6|你们没有吃饼，也没有喝清酒烈酒，好让你们知道‘我─耶和华是你们的上帝’。
DEUT|29|7|你们来到这地方， 希实本 王 西宏 和 巴珊 王 噩 出来迎击我们，与我们交战，我们击败了他们，
DEUT|29|8|取了他们的地，给 吕便 支派、 迦得 支派和 玛拿西 半支派为业。
DEUT|29|9|所以你们要谨守这约的话，遵行它们，好使你们在一切所做的事上亨通。
DEUT|29|10|“今日你们全都要站在耶和华－你们的上帝面前，就是各领袖、族长 、长老、官长、 以色列 所有的男子、
DEUT|29|11|你们的妻子儿女、你营中寄居的，从为你砍柴到为你挑水的人，
DEUT|29|12|为要使你进入耶和华－你上帝的约，就是耶和华－你上帝今日向你起誓所立的；
DEUT|29|13|这样，他今日要立你作他的子民，他作你的上帝，是照他向你所应许的，又照他向你列祖 亚伯拉罕 、 以撒 、 雅各 所起的誓。
DEUT|29|14|我不单单与你们立这约，起这誓，
DEUT|29|15|就是今日与我们一同站在耶和华－我们上帝面前的，而且也包括今日不在我们这里的人。
DEUT|29|16|“你们知道，我们曾住过 埃及 地，也经过列国，从他们中间穿越。
DEUT|29|17|你们也见过他们的可憎之物，他们木、石、金、银的偶像。
DEUT|29|18|惟恐你们中间有人，或男或女，或宗族或支派，今日心里偏离耶和华－我们的上帝，去事奉那些国的神明，又怕你们中间有根长出苦菜和茵蔯来。
DEUT|29|19|这样的人听见这诅咒的话，心里还庆幸，说：‘我虽然随着顽固的心行事，却还是平安无事。’以致有水的和无水的都消灭了。
DEUT|29|20|耶和华必不愿饶恕他；耶和华的怒气与妒忌必向他如烟冒出，将这书上所写的一切诅咒都加在他身上，耶和华也要从天下涂去他的名。
DEUT|29|21|耶和华又必照着写在律法书上，约中的一切诅咒，将他从 以色列 众支派中分别出来，使他遭受祸害。
DEUT|29|22|你们的后代，就是接续你们兴起的子孙，和远方来的外邦人，看见这地的灾祸，以及耶和华所降于这地的疾病，
DEUT|29|23|遍地都被硫磺和盐所侵蚀，不能耕种，没有出产，连草都长不出来，好像耶和华在怒气和愤怒中所倾覆的 所多玛 、 蛾摩拉 、 押玛 、 洗扁 一样，
DEUT|29|24|万国必说：‘耶和华为什么向此地这样做呢？为什么要大发烈怒呢？’
DEUT|29|25|人必说：‘这是因为这地的人离弃了耶和华─他们列祖的上帝领他们出 埃及 地的时候与他们所立的约，
DEUT|29|26|去事奉别神，敬拜他们所不认识的神明，这是耶和华未曾允许的。
DEUT|29|27|所以耶和华的怒气向这地发作，将这书上所写的一切诅咒都降在这地上。
DEUT|29|28|耶和华在怒气、愤怒、大恼恨中将他们从本地拔出来，扔到别的地上，像今日一样。’
DEUT|29|29|“隐秘的事是属耶和华─我们上帝的，但明显的事是永远属我们和我们子孙的，为要叫我们遵行这律法上的一切话。”
DEUT|30|1|“当这一切的事，就是我摆在你面前的祝福和诅咒临到你的时候，你在耶和华－你上帝赶逐你去的万国中，心里回想这些事，
DEUT|30|2|你和你的子孙若尽心尽性归向耶和华－你的上帝，照我今日一切所吩咐你的，听从他的话，
DEUT|30|3|耶和华－你的上帝就必怜悯你，使你这被掳的子民归回。耶和华－你的上帝必转回，从分散你到的万民中把你召集回来。
DEUT|30|4|你就是被赶逐到天涯，耶和华－你的上帝也必从那里召集你，从那里领你回来。
DEUT|30|5|耶和华－你的上帝必领你进入你列祖所得的地，你必得着这地为业。他必善待你，使你增多，胜过你的列祖。
DEUT|30|6|耶和华－你的上帝要使你的心和你后裔的心受割礼，好叫你尽心尽性爱耶和华－你的上帝，使你可以存活。
DEUT|30|7|耶和华－你的上帝必将这一切诅咒加在你仇敌和恨恶你、迫害你的人身上。
DEUT|30|8|你必回转，听从耶和华的话，遵行他的一切诫命，就是我今日所吩咐你的。
DEUT|30|9|耶和华－你的上帝必使你手里所做的一切，以及你身所生的，牲畜所生的，土地所产的都丰富有余，而且顺利；耶和华必再喜爱善待你，正如他喜爱你的列祖一样，
DEUT|30|10|只要你听从耶和华－你上帝的话，谨守这律法书上所写的诫命律例，尽心尽性归向耶和华－你的上帝。”
DEUT|30|11|“我今日所吩咐你的诫命，对你并不困难，也不太远；
DEUT|30|12|不是在天上，使你说：‘谁为我们上天去取来给我们，使我们听了可以遵行呢？’
DEUT|30|13|也不是在海的那边，使你说：‘谁为我们渡海到另一边，去取来给我们，使我们听了可以遵行呢？’
DEUT|30|14|因这话离你很近，就在你口中，在你心里，使你可以遵行。
DEUT|30|15|“看，我今日将生死祸福摆在你面前。
DEUT|30|16|我今日所吩咐你的 ，就是要爱耶和华－你的上帝，遵行他的道，谨守他的诫命、律例、典章，使你可以存活，增多，而且耶和华－你的上帝必在你所要进去得为业的地上赐福给你。
DEUT|30|17|倘若你的心偏离，不肯听从，却被引诱去敬拜别神，事奉它们，
DEUT|30|18|我今日向你们申明，你们必定灭亡；在你过 约旦河 进去得为业的地上，你的日子必不长久。
DEUT|30|19|我今日呼天唤地向你作见证：我已经将生与死，祝福与诅咒，摆在你面前。所以你要拣选生命，好使你和你的后裔都得存活。
DEUT|30|20|要爱耶和华－你的上帝，听从他的话，紧紧跟随他，因为他是你的生命，必使你的日子得以长久，可以在耶和华向你列祖 亚伯拉罕 、 以撒 、 雅各 起誓要给他们的地上居住。”
DEUT|31|1|摩西 去把这些话吩咐 以色列 众人 ，
DEUT|31|2|对他们说：“我已经一百二十岁了，现在不能照常出入。耶和华曾对我说：‘你不得过这 约旦河 。’
DEUT|31|3|耶和华－你的上帝必在你面前过河，把这些国从你面前除灭，你就必得他们的地。 约书亚 要在你面前过河，是照耶和华所吩咐的。
DEUT|31|4|耶和华必对待他们，如同从前待他所除灭的 亚摩利 人的王 西宏 与 噩 ，以及他们的国一样。
DEUT|31|5|耶和华必将他们交在你们面前，你们要照我所吩咐的一切命令待他们。
DEUT|31|6|你们当刚强壮胆，不要害怕，也不要畏惧他们，因为耶和华－你的上帝必与你同去；他必不撇下你，也不丢弃你。”
DEUT|31|7|摩西 召了 约书亚 来，在 以色列 众人眼前对他说：“你当刚强壮胆！因为你要和这百姓一同进入 耶和华向他们列祖起誓要给他们的地，你也要使他们承受那地为业。
DEUT|31|8|耶和华必在你前面行，他必亲自与你同在，必不撇下你，也不丢弃你。你不要惧怕，也不要惊惶。”
DEUT|31|9|摩西 写下这律法，交给抬耶和华约柜的 利未 人祭司和 以色列 的众长老。
DEUT|31|10|摩西 吩咐他们说：“每逢七年的最后一年，就是定期的豁免年，在住棚节的时候，
DEUT|31|11|当 以色列 众人来到耶和华－你上帝所选择的地方朝见他的时候，你要在 以色列 众人面前念这律法给他们听。
DEUT|31|12|要召集百姓，男人、女人、孩子，和在你城里寄居的，叫他们都得以听见，好学习敬畏耶和华－你们的上帝，谨守遵行这律法的一切话。
DEUT|31|13|他们的儿女，就是那未曾认识的，也可以听，学习敬畏耶和华－你们的上帝；你们一生的日子，在你们过 约旦河 得为业的地上，都要这样做。”
DEUT|31|14|耶和华对 摩西 说：“看哪，你的死期已近了。要召 约书亚 来，和你一起站在会幕里，我好吩咐他。”于是 摩西 和 约书亚 去站在会幕里。
DEUT|31|15|耶和华在会幕里，在云柱中显现，云柱停在会幕门口的上面。
DEUT|31|16|耶和华对 摩西 说：“看哪，你必和你的祖先同睡。这百姓要起来，在他们所要去的地上，在那地的人中，随从外邦的神明行淫，离弃我，违背我与他们所立的约。
DEUT|31|17|那时，我的怒气必向他们发作，我必离弃他们，转脸不顾他们，以致他们被吞灭，并有许多的祸患灾难临到他们。在那日，人必说：‘这些祸患临到我，岂不是因为我的上帝不在我中间吗？’
DEUT|31|18|在那日，因人偏向别神所行的一切恶事，我必定转脸不顾。
DEUT|31|19|现在你们要写下这首歌，教导 以色列 人，放在他们口中，使这首歌成为我指责 以色列 人的见证。
DEUT|31|20|因为我将他们领进我向他们列祖起誓应许那流奶与蜜之地，他们在那里吃得饱足，长得肥胖，就偏向别神，事奉它们，藐视我，背弃我的约。
DEUT|31|21|当许多祸患灾难临到他们的时候，这首歌必在他们面前作见证，因为他们后裔的口必吟诵不忘。我未领他们到我所起誓应许之地以先，他们所怀的意念我都知道了。”
DEUT|31|22|当日 摩西 就写了一首歌，教导 以色列 人。
DEUT|31|23|耶和华吩咐 嫩 的儿子 约书亚 说：“你当刚强壮胆，因为你必领 以色列 人进入我所起誓应许他们的地，我必与你同在。”
DEUT|31|24|当 摩西 把这律法的话写完在书上，到完成的时候，
DEUT|31|25|摩西 吩咐抬耶和华约柜的 利未 人说：
DEUT|31|26|“把这律法书拿来，放在耶和华－你们上帝的约柜旁，可以在那里作指责你们的见证。
DEUT|31|27|因为我知道你们是悖逆的，是硬着颈项的。看哪，我今日还活着与你们同在，你们尚且悖逆耶和华，何况我死后呢？
DEUT|31|28|你们要召集你们支派的众长老和官长到我这里来，我好把这些话说给他们听，并且呼唤天地见证他们的不是。
DEUT|31|29|我知道我死后你们必全然败坏，偏离我所吩咐你们的道。日后必有祸患临到你们，因为你们做了耶和华眼中看为恶的事，以你们手中所做的惹他发怒。”
DEUT|31|30|摩西 把这首歌的话，从头到尾吟诵给 以色列 全会众听。
DEUT|32|1|“诸天哪，要侧耳听我说话； 愿地聆听我口中的言语。
DEUT|32|2|我的教导要淋漓如雨， 我的言语要滴落如露， 如细雨降在嫩草上， 如甘霖降在蔬菜中。
DEUT|32|3|因为我要宣扬耶和华的名， 你们要把伟大归给我们的上帝。
DEUT|32|4|“他是磐石，他的作为完全， 他一切所行的都公平； 他是信实无伪的上帝， 又公义，又正直。
DEUT|32|5|这乖僻弯曲的世代 向他行了败坏的事； 因着他们的弊病， 不再是他的儿女。
DEUT|32|6|愚昧无知的百姓啊， 你们这样报答耶和华吗？ 他岂不是你的父，创造了你吗？ 他造了你，坚立你。
DEUT|32|7|你当回想上古之日， 思念历代之年； 问你的父亲，他必告诉你； 问你的长者，他必向你述说。
DEUT|32|8|至高者将地业赐给列国， 将世人分开， 他按照神明 的数目， 为万民划定疆界。
DEUT|32|9|因为耶和华的份是他的百姓， 他的产业就是 雅各 。
DEUT|32|10|“耶和华在旷野之地， 在空旷，野兽吼叫之荒地遇见他， 就环绕他，看顾他， 保护他，如同保护眼中的瞳人。
DEUT|32|11|鹰怎样搅动巢窝， 在雏鹰上面飞翔， 展开双翅接住雏鹰， 背在两翼之上，
DEUT|32|12|耶和华也照样独自引导他， 并无外邦神明与他同在。
DEUT|32|13|耶和华使他驰骋在地的高处， 他吃田间的出产； 耶和华使他从岩石中吃蜜， 从坚石中吸油，
DEUT|32|14|也吃牛的乳酪、羊的奶、 羔羊的脂肪， 巴珊 所出的公绵羊和山羊， 和上好的麦子。 你要喝葡萄汁酿的美酒。
DEUT|32|15|“ 耶书仑 渐渐肥胖，能踼跳。 你长得肥胖，粗壮，丰润。 他离弃造他的上帝， 轻看救他的磐石。
DEUT|32|16|他们用外邦神明惹上帝妒忌， 以可憎之物惹他发怒。
DEUT|32|17|他们祭祀鬼魔，而非上帝， 是他们不认识的神明， 是近来新兴的， 是你们列祖所不畏惧的。
DEUT|32|18|你轻忽生你的磐石， 忘记生产你的上帝。
DEUT|32|19|“耶和华看见了， 因他儿女惹动他就抛弃他们，
DEUT|32|20|说：‘我要转脸离开他们， 看他们的结局如何。 他们是极乖谬的世代， 是不忠实的儿女。
DEUT|32|21|他们以那不是上帝的激起我妒忌， 以虚无的神明 惹我发怒。 我也要以不成国的激起你们嫉妒， 我要以愚顽的国惹起你们发怒。
DEUT|32|22|因为我的怒火焚烧， 直烧到极深的阴间， 吞噬地和地的出产， 连山的根基也烧着了。
DEUT|32|23|“‘我要把祸患堆在他们身上， 我用尽我的箭射向他们：
DEUT|32|24|饿死人的饥荒、 灼人的热症、 痛苦的灾害。 我要叫野兽用牙齿咬他们， 叫土中爬行的用毒液害他们。
DEUT|32|25|外有刀剑使人丧亡， 内有惊恐， 少男少女是如此， 吃奶的、白发的也是如此。
DEUT|32|26|我曾说，我要粉碎他们， 使他们的名 从人间消失。
DEUT|32|27|惟恐仇敌挑衅， 他们的敌人误解， 说，我们的手得胜了， 这一切并非耶和华做的。’
DEUT|32|28|“因为他们是缺乏智谋的国家， 他们里面毫无聪明。
DEUT|32|29|惟愿他们有智慧，能明白这事， 他们就会想到自己的结局。
DEUT|32|30|若非他们的磐石卖了他们， 若非耶和华交出他们， 一人岂能追赶千人， 二人焉能使万人逃跑呢？
DEUT|32|31|甚至我们的仇敌都承认， 他们的磐石不如我们的磐石。
DEUT|32|32|他们的葡萄树是 所多玛 的葡萄树， 是 蛾摩拉 田园所长的； 他们的葡萄是毒葡萄， 整串都是苦的。
DEUT|32|33|他们的酒是大蛇的毒液， 是毒蛇剧烈的毒汁。
DEUT|32|34|“这岂不都存放在我这里， 封存在我库房中吗？
DEUT|32|35|伸冤报应在我 ， 到了时候他们会失脚。 因为他们遭难的日子近了， 他们的厄运快要临到。
DEUT|32|36|耶和华见他的百姓毫无能力， 无论是为奴的、自由的，都没有存留， 就必为他们伸冤， 为自己的仆人发怜悯。
DEUT|32|37|他必说：‘他们的神明， 他们所投靠的磐石，在哪里呢？
DEUT|32|38|吃了他们祭牲脂肪的， 喝了他们浇酒祭之酒的， 叫那些神明站出来帮助你们， 作为你们的保障吧！
DEUT|32|39|“‘如今，看！我，惟有我是上帝 ； 我以外并无别神。 我使人死，我使人活； 我击伤人，也医治人， 没有人能从我手中救出来。
DEUT|32|40|我向天举手， 我凭我的永生起誓说：
DEUT|32|41|我若磨我闪亮的刀， 我的手掌握审判权， 就必报复我的敌人， 报应那些恨我的人。
DEUT|32|42|我要使我的箭饮血而醉， 就是被杀被掳之人的血； 我的刀也要吃肉， 就是仇敌披发头颅 的肉。’
DEUT|32|43|“列国啊，当与耶和华的子民一同欢呼 ； 因为他要为他仆人 所流的血伸冤， 报应他的敌人 ， 救赎他的土地和他的子民 。”
DEUT|32|44|摩西 和 嫩 的儿子 约书亚 前来把这首歌的一切话吟诵给百姓听。
DEUT|32|45|摩西 向 以色列 众人吟诵完了这一切话，
DEUT|32|46|对他们说：“我今日以这一切话警戒你们，你们都要记在心中，要吩咐你们的子孙谨守遵行这律法上一切的话。
DEUT|32|47|因为这不是与你们无关的空话，而是你们的生命；因遵行这话，你们的日子必在你们过 约旦河 得为业的地上得以长久。”
DEUT|32|48|就在那日，耶和华吩咐 摩西 说：
DEUT|32|49|“你上 摩押 地的 亚巴琳山脉 ，到面对 耶利哥 的 尼波山 去，看我所要赐给 以色列 人为业的 迦南 地。
DEUT|32|50|你必死在你所登的山上，归到你祖先 那里，像你哥哥 亚伦 死在 何珥山 上，归到他祖先 那里一样。
DEUT|32|51|因为你们在 以色列 人中得罪了我，在 寻 的旷野， 加低斯 的 米利巴 水那里，在 以色列 人中没有尊我为圣。
DEUT|32|52|我所赐给 以色列 人的地，你只可从对面观看，却不得进到那里去。”
DEUT|33|1|这是神人 摩西 未死以前为 以色列 人的祝福。
DEUT|33|2|他说： “耶和华从 西奈 来， 从 西珥 向他们显现， 从 巴兰山 发出光辉； 从万万圣者中来临 ， 从他右手向他们发出烈火的律法 。
DEUT|33|3|他实在疼爱万民。 他的众圣徒都在你手中， 他们坐在你的脚下， 领受你的言语。”
DEUT|33|4|摩西 将律法传给我们， 作为 雅各 会众的产业。
DEUT|33|5|“耶和华 在 耶书仑 作王； 百姓的众领袖和 以色列 各支派一同欢聚。
DEUT|33|6|愿 吕便 存活，不致死亡， 虽然他的人丁稀少。
DEUT|33|7|关于 犹大 ，他这么说： ‘耶和华啊，求你垂听 犹大 的声音， 引导他归回他的百姓中。 他曾用手为自己争战， 你必帮助他攻击敌人。’
DEUT|33|8|关于 利未 ，他说： ‘愿你的土明和乌陵都在你的虔诚人那里 。 你在 玛撒 曾考验他， 在 米利巴 水与他争论。
DEUT|33|9|关于自己的父母，他说：我未曾关注。 他的弟兄，他不承认， 他的儿女，他也不认识， 因为 利未 人遵行你的话， 谨守你的约。
DEUT|33|10|他们将你的典章教导 雅各 ， 将你的律法教导 以色列 。 他们奉上香让你闻， 把全牲的燔祭献在你坛上。
DEUT|33|11|求耶和华赐福给他的财物 ， 悦纳他手里的工作。 求你刺透起来攻击他的人的腰， 使那些恨恶他的人不再起来。’
DEUT|33|12|关于 便雅悯 ，他说： ‘耶和华所亲爱的必同耶和华安然居住， 耶和华终日庇护他， 他也住在耶和华两肩之中 。’
DEUT|33|13|关于 约瑟 ，他说： ‘愿他的地蒙耶和华赐福， 得天上的甘露， 地下的泉源；
DEUT|33|14|得太阳下的美果， 月光中的佳谷；
DEUT|33|15|得古老山岳的至宝， 永恒山岭的宝物；
DEUT|33|16|得地的宝物和其中所充满的， 得住在荆棘中者的喜悦。 愿这些福都临到 约瑟 的头上， 临到那与兄弟有分别之人的头顶上。
DEUT|33|17|他是牛群中头生的， 大有威严； 他的双角是野牛的角， 用以抵触万民，直到地极。 这对角是 以法莲 的万万， 这对角是 玛拿西 的千千。’
DEUT|33|18|关于 西布伦 ，他说： ‘ 西布伦 哪，你出外可以欢喜。 以萨迦 啊，你在帐棚里可以快乐。
DEUT|33|19|他们要召集万民到山上， 在那里献公义的祭。 因为他们要吸取海里的财富， 沙中隐藏的珍宝。’
DEUT|33|20|关于 迦得 ，他说： ‘那使 迦得 扩张的，当受称颂！ 迦得 卧如母狮， 撕裂膀臂和头皮。
DEUT|33|21|他为自己看中了最好的， 因为那是为掌权者所存留的一份。 他与百姓的领袖同来 ， 执行耶和华的公义 和耶和华为 以色列 所立的典章。’
DEUT|33|22|关于 但 ，他说： ‘ 但 是小狮子， 从 巴珊 跳出来。’
DEUT|33|23|关于 拿弗他利 ，他说： ‘ 拿弗他利 啊，你享足恩宠， 满得耶和华的福， 可以得西方和南方为业。’
DEUT|33|24|关于 亚设 ，他说： ‘愿 亚设 在众子中蒙福 ， 愿他得他弟兄的喜悦， 可以把脚蘸在油中。
DEUT|33|25|你的门闩是铁的，是铜的。 只要你有多少日子，你就有多少力量 。’
DEUT|33|26|“ 耶书仑 哪，没有谁能比上帝！ 他腾云，大显威荣， 从天空来帮助你。
DEUT|33|27|亘古的上帝是避难所， 下面有永久的膀臂。 他从你面前赶走仇敌， 说：‘毁灭吧！’
DEUT|33|28|因此， 以色列 独自安然居住， 雅各 的泉源在五谷新酒之地， 他的天也滴下露水。
DEUT|33|29|以色列 啊，你有福了！ 蒙耶和华拯救的百姓啊，谁能像你？ 他是帮助你的盾牌， 是你威荣的刀剑。 你的仇敌要屈身就你； 你却要践踏他们的背脊 。”
DEUT|34|1|摩西 从 摩押 平原登上 尼波山 ，到了 耶利哥 对面的 毗斯迦山 顶。耶和华把全地指给他看：从 基列 到 但 ，
DEUT|34|2|拿弗他利 全地， 以法莲 、 玛拿西 的地， 犹大 全地直到西边的海，
DEUT|34|3|尼革夫 ，从棕树城 耶利哥 的平原到 琐珥 。
DEUT|34|4|耶和华对他说：“这就是我向 亚伯拉罕 、 以撒 、 雅各 起誓应许之地，说：‘我必将这地赐给你的后裔。’现在我使你亲眼看见了，你却不得过到那里去。”
DEUT|34|5|于是耶和华的仆人 摩西 死在 摩押 地那里，正如耶和华所说的。
DEUT|34|6|耶和华将他葬在 摩押 地， 伯．毗珥 对面的谷中，只是到今日，没有人知道他的坟墓。
DEUT|34|7|摩西 死的时候一百二十岁，眼目没有昏花，力量没有衰退。
DEUT|34|8|以色列 人在 摩押 平原为 摩西 哀哭了三十天，为 摩西 哀哭居丧的日期才结束。
DEUT|34|9|嫩 的儿子 约书亚 ，因为 摩西 曾为他按手，他就被智慧的灵充满。 以色列 人听从他，照着耶和华所吩咐 摩西 的去做。
DEUT|34|10|以后， 以色列 中再没有兴起一位先知像 摩西 的，他是耶和华面对面所认识的。
DEUT|34|11|耶和华差派他在 埃及 地，向法老和他的一切臣仆，以及他的全地，行了各样神迹奇事，
DEUT|34|12|又在 以色列 众人眼前显出大能的手，行了一切大而可畏的事。
