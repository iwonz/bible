JOEL|1|1|耶和華的話臨到 毗土珥 的兒子 約珥 。
JOEL|1|2|老年人哪，當聽這話； 這地所有的居民哪，要側耳而聽。 在你們的日子， 或你們祖先的日子， 曾發生過這樣的事嗎？
JOEL|1|3|你們要將這事傳與子， 子傳與孫， 孫傳與後代。
JOEL|1|4|剪蟲吃剩的，蝗蟲來吃； 蝗蟲吃剩的，蝻子來吃； 蝻子吃剩的，螞蚱 來吃。
JOEL|1|5|醉酒的人哪，要清醒，要哭泣； 好酒的人哪，都要為甜酒哀號， 因為酒從你們的口中斷絕了。
JOEL|1|6|有一隊蝗蟲 ，強盛且不可數， 上來侵犯我的地； 牠的牙齒如獅子的牙齒， 如母獅的大牙。
JOEL|1|7|牠毀壞我的葡萄樹， 撕裂我的無花果樹， 剝光又丟棄，使枝條露白。
JOEL|1|8|你要像童女腰束麻布， 為她年少時的丈夫哀號。
JOEL|1|9|耶和華的殿中斷絕素祭和澆酒祭， 事奉耶和華的祭司都悲哀。
JOEL|1|10|田荒涼，地悲哀； 因為五穀毀壞， 新酒枯竭， 新的油也缺乏。
JOEL|1|11|農夫啊，要慚愧； 修整葡萄園的啊，你們要哀號； 因為大麥、小麥與田間的莊稼全都毀了。
JOEL|1|12|葡萄樹枯乾， 無花果樹衰殘， 石榴樹、棕樹、蘋果樹， 田野一切的樹木都枯乾； 眾人的喜樂盡都消逝。
JOEL|1|13|祭司啊，當束上麻布痛哭； 事奉祭壇的啊，要哀號； 事奉我上帝的啊，你們要來，披上麻布過夜， 因為在你們上帝的殿中不再有素祭和澆酒祭了。
JOEL|1|14|你們要使禁食的日子分別為聖， 宣告嚴肅會， 召集長老和這地所有的居民 來到耶和華－你們上帝的殿， 向耶和華哀求。
JOEL|1|15|哀哉，這日子！ 因為耶和華的日子臨近， 好像毀滅從全能者來到。
JOEL|1|16|糧食不是在我們眼前斷絕了嗎？ 歡喜快樂不是從我們上帝的殿中止息了嗎？
JOEL|1|17|種子在土塊下朽爛， 倉荒涼，廩破壞， 因為五穀枯乾了。
JOEL|1|18|牲畜哀鳴， 牛群混亂，因無草場， 羊群也受苦。
JOEL|1|19|耶和華啊，我向你求告， 因為有火吞噬野地的草場， 火焰燒盡田野的樹木。
JOEL|1|20|田野的走獸切慕你， 因為溪水乾涸， 火吞噬了野地的草場。
JOEL|2|1|你們要在 錫安 吹角， 在我的聖山發出警報。 這地所有的居民要發顫， 因為耶和華的日子快到， 已經臨近了。
JOEL|2|2|那是黑暗、陰森的日子， 是密雲、烏黑的日子， 如同黎明籠罩山嶺。 有一隊蝗蟲，又大又強， 自古以來沒有像這樣的， 以後直到萬代也必沒有。
JOEL|2|3|牠們前面有火吞噬， 後面有火焰燒盡。 牠們未到以前，地如 伊甸園 ， 過去以後，卻成了荒涼的曠野， 沒有一樣能躲避牠們。
JOEL|2|4|牠們形狀如馬， 奔跑如戰馬。
JOEL|2|5|響聲如戰車在山頂上跳動， 如火焰吞噬碎秸， 好像強大的軍隊擺陣備戰。
JOEL|2|6|在牠們面前，萬民傷慟， 臉都變色。
JOEL|2|7|牠們如勇士奔跑， 如戰士攀登城牆， 各行於自己的道路， 不亂隊伍；
JOEL|2|8|牠們並不彼此推擠， 各行於自己的大道， 衝過防禦 ， 並不停止。
JOEL|2|9|牠們蹦上城， 跳上牆， 爬上房屋， 從窗戶進來，如同盜賊。
JOEL|2|10|在牠們面前， 地動天搖， 日月昏暗， 星宿無光。
JOEL|2|11|耶和華在他的軍旅前出聲， 他的隊伍龐大， 遵行他命令的強盛。 耶和華的日子大而可畏， 誰能當得起呢？
JOEL|2|12|然而你們現在要禁食，哭泣，哀號， 一心歸向我。 這是耶和華說的。
JOEL|2|13|你們要撕裂心腸， 不要撕裂衣服。 歸向耶和華－你們的上帝， 因為他有恩惠，有憐憫， 不輕易發怒， 有豐盛的慈愛， 並且會改變心意， 不降那災難。
JOEL|2|14|誰知道他也許會回心轉意，留下餘福， 就是獻給耶和華－你們上帝的素祭和澆酒祭。
JOEL|2|15|你們要在 錫安 吹角， 使禁食的日子分別為聖， 宣告嚴肅會。
JOEL|2|16|聚集百姓，使會眾自潔； 召集老年人， 聚集孩童和在母懷吃奶的； 使新郎出內室， 新娘離開洞房。
JOEL|2|17|事奉耶和華的祭司 要在走廊和祭壇間哭泣，說： 「耶和華啊，求你顧惜你的百姓， 不要使你的產業受羞辱， 在列國中成為笑柄。 為何讓人在萬民中說 『他們的上帝在哪裏』呢？」
JOEL|2|18|耶和華為自己的地發熱心， 憐憫他的百姓。
JOEL|2|19|耶和華應允他的百姓說： 「看哪，我要賞賜你們五穀、新酒和新的油， 使你們飽足， 我必不再使你們受列國的羞辱。
JOEL|2|20|我要使北方來的隊伍遠離你們， 將他們趕到乾旱荒蕪之地： 前隊趕入東海， 後隊趕入西海； 臭氣上升，惡臭騰空。 耶和華果然行了大事！
JOEL|2|21|「土地啊，不要懼怕， 要歡喜快樂， 因為耶和華行了大事。
JOEL|2|22|田野的走獸啊，不要懼怕， 因為曠野的草已生長， 樹木結果， 無花果樹、葡萄樹也都效力 。
JOEL|2|23|「 錫安 的民哪，你們要歡喜， 要因耶和華－你們的上帝快樂； 因他賞賜你們合宜的秋雨 ， 為你們降下甘霖， 秋雨和春雨，和先前一樣。
JOEL|2|24|「禾場充滿五穀， 池中漫溢新酒和新的油。
JOEL|2|25|我差遣到你們中間的大軍隊， 就是蝗蟲、蝻子、螞蚱、剪蟲， 那些年間所吃的，我要補還給你們。
JOEL|2|26|「你們必吃得飽足， 讚美耶和華－你們上帝的名， 他為你們行了奇妙的事。 我的百姓不致羞愧，直到永遠。
JOEL|2|27|你們必知道我是在 以色列 中， 又知道我是耶和華－你們的上帝，沒有別的。 我的百姓不致羞愧，直到永遠。」
JOEL|2|28|「以後，我要將我的靈澆灌凡有血肉之軀的。 你們的兒女要說預言， 你們的老人要做異夢， 你們的少年要見異象。
JOEL|2|29|在那些日子， 我要將我的靈澆灌我的僕人和婢女。
JOEL|2|30|「我要在天上地下顯出奇事，有血，有火，有煙柱。
JOEL|2|31|太陽要變為黑暗，月亮要變為血，這都在耶和華大而可畏的日子未到以前。
JOEL|2|32|那時，凡求告耶和華名的就必得救；因為照耶和華所說的，在 錫安山 ，在 耶路撒冷 將有逃脫的人。凡耶和華所召的 ，都在餘民之列。」
JOEL|3|1|「看哪，在那些日子，到那個時候，我使 猶大 和 耶路撒冷 被擄之人歸回的時候，
JOEL|3|2|我要聚集萬民，帶他們下到 約沙法谷 去，在那裏我要為我百姓，我產業 以色列 的緣故，向萬民施行審判；因為他們把我的百姓分散到列國，瓜分了我的土地，
JOEL|3|3|為我的百姓抽籤，以男孩換取妓女，為喝酒賣掉女孩。
JOEL|3|4|「 推羅 、 西頓 和 非利士 四境的人哪，你們與我何干？你們要報復我嗎？若要報復我，我必使報應速速歸到你們頭上。
JOEL|3|5|你們奪取我的金銀，把我珍貴的寶物帶入你們的廟宇 ，
JOEL|3|6|並將 猶大 人和 耶路撒冷 人賣給 希臘 人 ，使他們遠離自己的疆土。
JOEL|3|7|看哪，我必激發他們離開你們把他們賣去的地方，又必使報應歸到你們頭上。
JOEL|3|8|我要將你們的兒女賣到 猶大 人手中，他們必轉賣給遠方的國家 示巴 人。這是耶和華說的。」
JOEL|3|9|當在列國中宣告： 預備打仗， 激發勇士， 使所有戰士上前來。
JOEL|3|10|要將犁頭打成刀劍， 鐮刀打成戈矛； 弱者要說：「我是勇士。」
JOEL|3|11|四圍的列國啊， 要速速前來， 一同聚集。 耶和華啊， 求你使你的勇士降臨。
JOEL|3|12|列國都當興起， 上到 約沙法谷 ； 因為我必坐在那裏， 審判四圍的列國。
JOEL|3|13|揮鐮刀吧！因為莊稼熟了； 來踩踏吧！因為醡酒池滿了。 酒池已經滿溢， 因為他們的罪惡甚大。
JOEL|3|14|在 斷定谷 有許多許多的人， 因為耶和華的日子臨近 斷定谷 了。
JOEL|3|15|日月昏暗， 星宿無光。
JOEL|3|16|耶和華必從 錫安 吼叫， 從 耶路撒冷 出聲， 天地就震動。 耶和華卻要作他百姓的避難所， 作 以色列 人的保障。
JOEL|3|17|你們就知道我是耶和華－你們的上帝， 我住在 錫安 －我的聖山。 耶路撒冷 必成為聖； 陌生人不再從其中經過。
JOEL|3|18|在那日，大山要滴甜酒， 小山要流奶， 猶大 的溪河都有水流出； 必有泉源從耶和華的殿中流出， 滋潤 什亭谷 。
JOEL|3|19|埃及 必定荒涼， 以東 成為荒涼的曠野， 因為他們向 猶大 人行殘暴， 又因他們在本地流無辜人的血。
JOEL|3|20|但 猶大 必存到永遠， 耶路撒冷 必存到萬代。
JOEL|3|21|我要免除 流人血的罪， 是先前未曾免除的， 耶和華居住在 錫安 。
