PROV|1|1|parabolae Salomonis filii David regis Israhel
PROV|1|2|ad sciendam sapientiam et disciplinam
PROV|1|3|ad intellegenda verba prudentiae et suscipiendam eruditionem doctrinae iustitiam et iudicium et aequitatem
PROV|1|4|ut detur parvulis astutia adulescenti scientia et intellectus
PROV|1|5|audiens sapiens sapientior erit et intellegens gubernacula possidebit
PROV|1|6|animadvertet parabolam et interpretationem verba sapientium et enigmata eorum
PROV|1|7|timor Domini principium scientiae sapientiam atque doctrinam stulti despiciunt
PROV|1|8|audi fili mi disciplinam patris tui et ne dimittas legem matris tuae
PROV|1|9|ut addatur gratia capiti tuo et torques collo tuo
PROV|1|10|fili mi si te lactaverint peccatores ne adquiescas
PROV|1|11|si dixerint veni nobiscum insidiemur sanguini abscondamus tendiculas contra insontem frustra
PROV|1|12|degluttiamus eum sicut infernus viventem et integrum quasi descendentem in lacum
PROV|1|13|omnem pretiosam substantiam repperiemus implebimus domos nostras spoliis
PROV|1|14|sortem mitte nobiscum marsuppium unum sit omnium nostrum
PROV|1|15|fili mi ne ambules cum eis prohibe pedem tuum a semitis eorum
PROV|1|16|pedes enim illorum ad malum currunt et festinant ut effundant sanguinem
PROV|1|17|frustra autem iacitur rete ante oculos pinnatorum
PROV|1|18|ipsique contra sanguinem suum insidiantur et moliuntur fraudes contra animas suas
PROV|1|19|sic semitae omnis avari animas possidentium rapiunt
PROV|1|20|sapientia foris praedicat in plateis dat vocem suam
PROV|1|21|in capite turbarum clamitat in foribus portarum urbis profert verba sua dicens
PROV|1|22|usquequo parvuli diligitis infantiam et stulti ea quae sibi sunt noxia cupiunt et inprudentes odibunt scientiam
PROV|1|23|convertimini ad correptionem meam en proferam vobis spiritum meum et ostendam verba mea
PROV|1|24|quia vocavi et rennuistis extendi manum meam et non fuit qui aspiceret
PROV|1|25|despexistis omne consilium meum et increpationes meas neglexistis
PROV|1|26|ego quoque in interitu vestro ridebo et subsannabo cum vobis quod timebatis advenerit
PROV|1|27|cum inruerit repentina calamitas et interitus quasi tempestas ingruerit quando venerit super vos tribulatio et angustia
PROV|1|28|tunc invocabunt me et non exaudiam mane consurgent et non invenient me
PROV|1|29|eo quod exosam habuerint disciplinam et timorem Domini non susceperint
PROV|1|30|nec adquieverint consilio meo et detraxerint universae correptioni meae
PROV|1|31|comedent igitur fructus viae suae suisque consiliis saturabuntur
PROV|1|32|aversio parvulorum interficiet eos et prosperitas stultorum perdet illos
PROV|1|33|qui autem me audierit absque terrore requiescet et abundantia perfruetur malorum timore sublato
PROV|2|1|fili mi si susceperis sermones meos et mandata mea absconderis penes te
PROV|2|2|ut audiat sapientiam auris tua inclina cor tuum ad noscendam prudentiam
PROV|2|3|si enim sapientiam invocaveris et inclinaveris cor tuum prudentiae
PROV|2|4|si quaesieris eam quasi pecuniam et sicut thesauros effoderis illam
PROV|2|5|tunc intelleges timorem Domini et scientiam Dei invenies
PROV|2|6|quia Dominus dat sapientiam et ex ore eius scientia et prudentia
PROV|2|7|custodiet rectorum salutem et proteget gradientes simpliciter
PROV|2|8|servans semitas iustitiae et vias sanctorum custodiens
PROV|2|9|tunc intelleges iustitiam et iudicium et aequitatem et omnem semitam bonam
PROV|2|10|si intraverit sapientia cor tuum et scientia animae tuae placuerit
PROV|2|11|consilium custodiet te prudentia servabit te
PROV|2|12|ut eruaris de via mala ab homine qui perversa loquitur
PROV|2|13|qui relinquunt iter rectum et ambulant per vias tenebrosas
PROV|2|14|qui laetantur cum malefecerint et exultant in rebus pessimis
PROV|2|15|quorum viae perversae et infames gressus eorum
PROV|2|16|ut eruaris a muliere aliena et ab extranea quae mollit sermones suos
PROV|2|17|et relinquit ducem pubertatis suae
PROV|2|18|et pacti Dei sui oblita est inclinata est enim ad mortem domus eius et ad impios semitae ipsius
PROV|2|19|omnes qui ingrediuntur ad eam non revertentur nec adprehendent semitas vitae
PROV|2|20|ut ambules in via bona et calles iustorum custodias
PROV|2|21|qui enim recti sunt habitabunt in terra et simplices permanebunt in ea
PROV|2|22|impii vero de terra perdentur et qui inique agunt auferentur ex ea
PROV|3|1|fili mi ne obliviscaris legis meae et praecepta mea custodiat cor tuum
PROV|3|2|longitudinem enim dierum et annos vitae et pacem adponent tibi
PROV|3|3|misericordia et veritas non te deserant circumda eas gutturi tuo et describe in tabulis cordis tui
PROV|3|4|et invenies gratiam et disciplinam bonam coram Deo et hominibus
PROV|3|5|habe fiduciam in Domino ex toto corde tuo et ne innitaris prudentiae tuae
PROV|3|6|in omnibus viis tuis cogita illum et ipse diriget gressus tuos
PROV|3|7|ne sis sapiens apud temet ipsum time Dominum et recede a malo
PROV|3|8|sanitas quippe erit umbilico tuo et inrigatio ossuum tuorum
PROV|3|9|honora Dominum de tua substantia et de primitiis omnium frugum tuarum
PROV|3|10|et implebuntur horrea tua saturitate et vino torcularia redundabunt
PROV|3|11|disciplinam Domini fili mi ne abicias nec deficias cum ab eo corriperis
PROV|3|12|quem enim diligit Dominus corripit et quasi pater in filio conplacet sibi
PROV|3|13|beatus homo qui invenit sapientiam et qui affluit prudentia
PROV|3|14|melior est adquisitio eius negotiatione argenti et auro primo fructus eius
PROV|3|15|pretiosior est cunctis opibus et omnia quae desiderantur huic non valent conparari
PROV|3|16|longitudo dierum in dextera eius in sinistra illius divitiae et gloria
PROV|3|17|viae eius viae pulchrae et omnes semitae illius pacificae
PROV|3|18|lignum vitae est his qui adprehenderint eam et qui tenuerit eam beatus
PROV|3|19|Dominus sapientia fundavit terram stabilivit caelos prudentia
PROV|3|20|sapientia illius eruperunt abyssi et nubes rore concrescunt
PROV|3|21|fili mi ne effluant haec ab oculis tuis custodi legem atque consilium
PROV|3|22|et erit vita animae tuae et gratia faucibus tuis
PROV|3|23|tunc ambulabis fiducialiter in via tua et pes tuus non inpinget
PROV|3|24|si dormieris non timebis quiesces et suavis erit somnus tuus
PROV|3|25|ne paveas repentino terrore et inruentes tibi potentias impiorum
PROV|3|26|Dominus enim erit in latere tuo et custodiet pedem tuum ne capiaris
PROV|3|27|noli prohibere benefacere eum qui potest si vales et ipse benefac
PROV|3|28|ne dicas amico tuo vade et revertere et cras dabo tibi cum statim possis dare
PROV|3|29|ne moliaris amico tuo malum cum ille in te habeat fiduciam
PROV|3|30|ne contendas adversus hominem frustra cum ipse tibi nihil mali fecerit
PROV|3|31|ne aemuleris hominem iniustum nec imiteris vias eius
PROV|3|32|quia abominatio Domini est omnis inlusor et cum simplicibus sermocinatio eius
PROV|3|33|egestas a Domino in domo impii habitacula autem iustorum benedicentur
PROV|3|34|inlusores ipse deludet et mansuetis dabit gratiam
PROV|3|35|gloriam sapientes possidebunt stultorum exaltatio ignominia
PROV|4|1|audite filii disciplinam patris et adtendite ut sciatis prudentiam
PROV|4|2|donum bonum tribuam vobis legem meam ne derelinquatis
PROV|4|3|nam et ego filius fui patris mei tenellus et unigenitus coram matre mea
PROV|4|4|et docebat me atque dicebat suscipiat verba mea cor tuum custodi praecepta mea et vives
PROV|4|5|posside sapientiam posside prudentiam ne obliviscaris neque declines a verbis oris mei
PROV|4|6|ne dimittas eam et custodiet te dilige eam et servabit te
PROV|4|7|principium sapientiae posside sapientiam et in omni possessione tua adquire prudentiam
PROV|4|8|arripe illam et exaltabit te glorificaberis ab ea cum eam fueris amplexatus
PROV|4|9|dabit capiti tuo augmenta gratiarum et corona inclita proteget te
PROV|4|10|audi fili mi et suscipe verba mea ut multiplicentur tibi anni vitae
PROV|4|11|viam sapientiae monstravi tibi duxi te per semitas aequitatis
PROV|4|12|quas cum ingressus fueris non artabuntur gressus tui et currens non habebis offendiculum
PROV|4|13|tene disciplinam ne dimittas eam custodi illam quia ipsa est vita tua
PROV|4|14|ne delecteris semitis impiorum nec tibi placeat malorum via
PROV|4|15|fuge ab ea ne transeas per illam declina et desere eam
PROV|4|16|non enim dormiunt nisi malefecerint et rapitur somnus ab eis nisi subplantaverint
PROV|4|17|comedunt panem impietatis et vinum iniquitatis bibunt
PROV|4|18|iustorum autem semita quasi lux splendens procedit et crescit usque ad perfectam diem
PROV|4|19|via impiorum tenebrosa nesciunt ubi corruant
PROV|4|20|fili mi ausculta sermones meos et ad eloquia mea inclina aurem tuam
PROV|4|21|ne recedant ab oculis tuis custodi ea in medio cordis tui
PROV|4|22|vita enim sunt invenientibus ea et universae carni sanitas
PROV|4|23|omni custodia serva cor tuum quia ex ipso vita procedit
PROV|4|24|remove a te os pravum et detrahentia labia sint procul a te
PROV|4|25|oculi tui recta videant et palpebrae tuae praecedant gressus tuos
PROV|4|26|dirige semitam pedibus tuis et omnes viae tuae stabilientur
PROV|4|27|ne declines ad dexteram et ad sinistram averte pedem tuum a malo
PROV|5|1|fili mi adtende sapientiam meam et prudentiae meae inclina aurem tuam
PROV|5|2|ut custodias cogitationes et disciplinam labia tua conservent
PROV|5|3|favus enim stillans labia meretricis et nitidius oleo guttur eius
PROV|5|4|novissima autem illius amara quasi absinthium et acuta quasi gladius biceps
PROV|5|5|pedes eius descendunt in mortem et ad inferos gressus illius penetrant
PROV|5|6|per semitam vitae non ambulat vagi sunt gressus eius et investigabiles
PROV|5|7|nunc ergo fili audi me et ne recedas a verbis oris mei
PROV|5|8|longe fac ab ea viam tuam et ne adpropinques foribus domus eius
PROV|5|9|ne des alienis honorem tuum et annos tuos crudeli
PROV|5|10|ne forte impleantur extranei viribus tuis et labores tui sint in domo aliena
PROV|5|11|et gemas in novissimis quando consumpseris carnes et corpus tuum et dicas
PROV|5|12|cur detestatus sum disciplinam et increpationibus non adquievit cor meum
PROV|5|13|nec audivi vocem docentium me et magistris non inclinavi aurem meam
PROV|5|14|paene fui in omni malo in medio ecclesiae et synagogae
PROV|5|15|bibe aquam de cisterna tua et fluenta putei tui
PROV|5|16|deriventur fontes tui foras et in plateis aquas tuas divide
PROV|5|17|habeto eas solus nec sint alieni participes tui
PROV|5|18|sit vena tua benedicta et laetare cum muliere adulescentiae tuae
PROV|5|19|cerva carissima et gratissimus hinulus ubera eius inebrient te omni tempore in amore illius delectare iugiter
PROV|5|20|quare seduceris fili mi ab aliena et foveris sinu alterius
PROV|5|21|respicit Dominus vias hominis et omnes gressus illius considerat
PROV|5|22|iniquitates suae capiunt impium et funibus peccatorum suorum constringitur
PROV|5|23|ipse morietur quia non habuit disciplinam et multitudine stultitiae suae decipietur
PROV|6|1|fili mi si spoponderis pro amico tuo defixisti apud extraneum manum tuam
PROV|6|2|inlaqueatus es verbis oris tui et captus propriis sermonibus
PROV|6|3|fac ergo quod dico fili mi et temet ipsum libera quia incidisti in manu proximi tui discurre festina suscita amicum tuum
PROV|6|4|ne dederis somnum oculis tuis nec dormitent palpebrae tuae
PROV|6|5|eruere quasi dammula de manu et quasi avis de insidiis aucupis
PROV|6|6|vade ad formicam o piger et considera vias eius et disce sapientiam
PROV|6|7|quae cum non habeat ducem nec praeceptorem nec principem
PROV|6|8|parat aestate cibum sibi et congregat in messe quod comedat
PROV|6|9|usquequo piger dormis quando consurges ex somno tuo
PROV|6|10|paululum dormies paululum dormitabis paululum conseres manus ut dormias
PROV|6|11|et veniet tibi quasi viator egestas et pauperies quasi vir armatus
PROV|6|12|homo apostata vir inutilis graditur ore perverso
PROV|6|13|annuit oculis terit pede digito loquitur
PROV|6|14|pravo corde machinatur malum et in omni tempore iurgia seminat
PROV|6|15|huic extemplo veniet perditio sua et subito conteretur nec habebit ultra medicinam
PROV|6|16|sex sunt quae odit Dominus et septimum detestatur anima eius
PROV|6|17|oculos sublimes linguam mendacem manus effundentes innoxium sanguinem
PROV|6|18|cor machinans cogitationes pessimas pedes veloces ad currendum in malum
PROV|6|19|proferentem mendacia testem fallacem et eum qui seminat inter fratres discordias
PROV|6|20|conserva fili mi praecepta patris tui et ne dimittas legem matris tuae
PROV|6|21|liga ea in corde tuo iugiter et circumda gutturi tuo
PROV|6|22|cum ambulaveris gradiantur tecum cum dormieris custodiant te et evigilans loquere cum eis
PROV|6|23|quia mandatum lucerna est et lex lux et via vitae increpatio disciplinae
PROV|6|24|ut custodiant te a muliere mala et a blanda lingua extraneae
PROV|6|25|non concupiscat pulchritudinem eius cor tuum nec capiaris nutibus illius
PROV|6|26|pretium enim scorti vix unius est panis mulier autem viri pretiosam animam capit
PROV|6|27|numquid abscondere potest homo ignem in sinu suo ut vestimenta illius non ardeant
PROV|6|28|aut ambulare super prunas et non conburentur plantae eius
PROV|6|29|sic qui ingreditur ad mulierem proximi sui non erit mundus cum tetigerit eam
PROV|6|30|non grandis est culpae cum quis furatus fuerit furatur enim ut esurientem impleat animam
PROV|6|31|deprehensus quoque reddet septuplum et omnem substantiam domus suae tradet
PROV|6|32|qui autem adulter est propter cordis inopiam perdet animam suam
PROV|6|33|turpitudinem et ignominiam congregat sibi et obprobrium illius non delebitur
PROV|6|34|quia zelus et furor viri non parcet in die vindictae
PROV|6|35|nec adquiescet cuiusquam precibus nec suscipiet pro redemptione dona plurima
PROV|7|1|fili mi custodi sermones meos et praecepta mea reconde tibi
PROV|7|2|serva mandata mea et vives et legem meam quasi pupillam oculi tui
PROV|7|3|liga eam in digitis tuis scribe illam in tabulis cordis tui
PROV|7|4|dic sapientiae soror mea es et prudentiam voca amicam tuam
PROV|7|5|ut custodiat te a muliere extranea et ab aliena quae verba sua dulcia facit
PROV|7|6|de fenestra enim domus meae per cancellos prospexi
PROV|7|7|et video parvulos considero vecordem iuvenem
PROV|7|8|qui transit in platea iuxta angulum et propter viam domus illius graditur
PROV|7|9|in obscuro advesperascente die in noctis tenebris et caligine
PROV|7|10|et ecce mulier occurrit illi ornatu meretricio praeparata ad capiendas animas garrula et vaga
PROV|7|11|quietis inpatiens nec valens in domo consistere pedibus suis
PROV|7|12|nunc foris nunc in plateis nunc iuxta angulos insidians
PROV|7|13|adprehensumque deosculatur iuvenem et procaci vultu blanditur dicens
PROV|7|14|victimas pro salute debui hodie reddidi vota mea
PROV|7|15|idcirco egressa sum in occursum tuum desiderans te videre et repperi
PROV|7|16|intexui funibus lectum meum stravi tapetibus pictis ex Aegypto
PROV|7|17|aspersi cubile meum murra et aloe et cinnamomo
PROV|7|18|veni inebriemur uberibus donec inlucescat dies et fruamur cupitis amplexibus
PROV|7|19|non est enim vir in domo sua abiit via longissima
PROV|7|20|sacculum pecuniae secum tulit in die plenae lunae reversurus est domum suam
PROV|7|21|inretivit eum multis sermonibus et blanditiis labiorum protraxit illum
PROV|7|22|statim eam sequitur quasi bos ductus ad victimam et quasi agnus lasciviens et ignorans quod ad vincula stultus trahatur
PROV|7|23|donec transfigat sagitta iecur eius velut si avis festinet ad laqueum et nescit quia de periculo animae illius agitur
PROV|7|24|nunc ergo fili audi me et adtende verba oris mei
PROV|7|25|ne abstrahatur in viis illius mens tua neque decipiaris semitis eius
PROV|7|26|multos enim vulneratos deiecit et fortissimi quique interfecti sunt ab ea
PROV|7|27|viae inferi domus eius penetrantes interiora mortis
PROV|8|1|numquid non sapientia clamitat et prudentia dat vocem suam
PROV|8|2|in summis excelsisque verticibus super viam in mediis semitis stans
PROV|8|3|iuxta portas civitatis in ipsis foribus loquitur dicens
PROV|8|4|o viri ad vos clamito et vox mea ad filios hominum
PROV|8|5|intellegite parvuli astutiam et insipientes animadvertite
PROV|8|6|audite quoniam de rebus magnis locutura sum et aperientur labia mea ut recta praedicent
PROV|8|7|veritatem meditabitur guttur meum et labia mea detestabuntur impium
PROV|8|8|iusti sunt omnes sermones mei non est in eis pravum quid neque perversum
PROV|8|9|recti sunt intellegentibus et aequi invenientibus scientiam
PROV|8|10|accipite disciplinam meam et non pecuniam doctrinam magis quam aurum eligite
PROV|8|11|melior est enim sapientia cunctis pretiosissimis et omne desiderabile ei non potest conparari
PROV|8|12|ego sapientia habito in consilio et eruditis intersum cogitationibus
PROV|8|13|timor Domini odit malum arrogantiam et superbiam et viam pravam et os bilingue detestor
PROV|8|14|meum est consilium et aequitas mea prudentia mea est fortitudo
PROV|8|15|per me reges regnant et legum conditores iusta decernunt
PROV|8|16|per me principes imperant et potentes decernunt iustitiam
PROV|8|17|ego diligentes me diligo et qui mane vigilant ad me invenient me
PROV|8|18|mecum sunt divitiae et gloria opes superbae et iustitia
PROV|8|19|melior est fructus meus auro et pretioso lapide et genimina mea argento electo
PROV|8|20|in viis iustitiae ambulo in medio semitarum iudicii
PROV|8|21|ut ditem diligentes me et thesauros eorum repleam
PROV|8|22|Dominus possedit me initium viarum suarum antequam quicquam faceret a principio
PROV|8|23|ab aeterno ordita sum et ex antiquis antequam terra fieret
PROV|8|24|necdum erant abyssi et ego iam concepta eram necdum fontes aquarum eruperant
PROV|8|25|necdum montes gravi mole constiterant ante colles ego parturiebar
PROV|8|26|adhuc terram non fecerat et flumina et cardines orbis terrae
PROV|8|27|quando praeparabat caelos aderam quando certa lege et gyro vallabat abyssos
PROV|8|28|quando aethera firmabat sursum et librabat fontes aquarum
PROV|8|29|quando circumdabat mari terminum suum et legem ponebat aquis ne transirent fines suos quando adpendebat fundamenta terrae
PROV|8|30|cum eo eram cuncta conponens et delectabar per singulos dies ludens coram eo omni tempore
PROV|8|31|ludens in orbe terrarum et deliciae meae esse cum filiis hominum
PROV|8|32|nunc ergo filii audite me beati qui custodiunt vias meas
PROV|8|33|audite disciplinam et estote sapientes et nolite abicere eam
PROV|8|34|beatus homo qui audit me qui vigilat ad fores meas cotidie et observat ad postes ostii mei
PROV|8|35|qui me invenerit inveniet vitam et hauriet salutem a Domino
PROV|8|36|qui autem in me peccaverit laedet animam suam omnes qui me oderunt diligunt mortem
PROV|9|1|sapientia aedificavit sibi domum excidit columnas septem
PROV|9|2|immolavit victimas suas miscuit vinum et proposuit mensam suam
PROV|9|3|misit ancillas suas ut vocarent ad arcem et ad moenia civitatis
PROV|9|4|si quis est parvulus veniat ad me et insipientibus locuta est
PROV|9|5|venite comedite panem meum et bibite vinum quod miscui vobis
PROV|9|6|relinquite infantiam et vivite et ambulate per vias prudentiae
PROV|9|7|qui erudit derisorem ipse sibi facit iniuriam et qui arguit impium generat maculam sibi
PROV|9|8|noli arguere derisorem ne oderit te argue sapientem et diliget te
PROV|9|9|da sapienti et addetur ei sapientia doce iustum et festinabit accipere
PROV|9|10|principium sapientiae timor Domini et scientia sanctorum prudentia
PROV|9|11|per me enim multiplicabuntur dies tui et addentur tibi anni vitae
PROV|9|12|si sapiens fueris tibimet ipsi eris si inlusor solus portabis malum
PROV|9|13|mulier stulta et clamosa plenaque inlecebris et nihil omnino sciens
PROV|9|14|sedit in foribus domus suae super sellam in excelso urbis loco
PROV|9|15|ut vocaret transeuntes viam et pergentes itinere suo
PROV|9|16|quis est parvulus declinet ad me et vecordi locuta est
PROV|9|17|aquae furtivae dulciores sunt et panis absconditus suavior
PROV|9|18|et ignoravit quod gigantes ibi sint et in profundis inferni convivae eius
PROV|10|1|parabolae Salomonis filius sapiens laetificat patrem filius vero stultus maestitia est matris suae
PROV|10|2|non proderunt thesauri impietatis iustitia vero liberabit a morte
PROV|10|3|non adfliget Dominus fame animam iusti et insidias impiorum subvertet
PROV|10|4|egestatem operata est manus remissa manus autem fortium divitias parat
PROV|10|5|qui congregat in messe filius sapiens est qui autem stertit aestate filius confusionis
PROV|10|6|benedictio super caput iusti os autem impiorum operit iniquitatem
PROV|10|7|memoria iusti cum laudibus et nomen impiorum putrescet
PROV|10|8|sapiens corde praecepta suscipiet stultus caeditur labiis
PROV|10|9|qui ambulat simpliciter ambulat confidenter qui autem depravat vias suas manifestus erit
PROV|10|10|qui annuit oculo dabit dolorem stultus labiis verberabitur
PROV|10|11|vena vitae os iusti et os impiorum operiet iniquitatem
PROV|10|12|odium suscitat rixas et universa delicta operit caritas
PROV|10|13|in labiis sapientis invenietur sapientia et virga in dorso eius qui indiget corde
PROV|10|14|sapientes abscondunt scientiam os autem stulti confusioni proximum est
PROV|10|15|substantia divitis urbs fortitudinis eius pavor pauperum egestas eorum
PROV|10|16|opus iusti ad vitam fructus impii ad peccatum
PROV|10|17|via vitae custodienti disciplinam qui autem increpationes relinquit errat
PROV|10|18|abscondunt odium labia mendacia qui profert contumeliam insipiens est
PROV|10|19|in multiloquio peccatum non deerit qui autem moderatur labia sua prudentissimus est
PROV|10|20|argentum electum lingua iusti cor impiorum pro nihilo
PROV|10|21|labia iusti erudiunt plurimos qui autem indocti sunt in cordis egestate morientur
PROV|10|22|benedictio Domini divites facit nec sociabitur ei adflictio
PROV|10|23|quasi per risum stultus operatur scelus sapientia autem est viro prudentia
PROV|10|24|quod timet impius veniet super eum desiderium suum iustis dabitur
PROV|10|25|quasi tempestas transiens non erit impius iustus autem quasi fundamentum sempiternum
PROV|10|26|sicut acetum dentibus et fumus oculis sic piger his qui miserunt eum
PROV|10|27|timor Domini adponet dies et anni impiorum breviabuntur
PROV|10|28|expectatio iustorum laetitia spes autem impiorum peribit
PROV|10|29|fortitudo simplicis via Domini et pavor his qui operantur malum
PROV|10|30|iustus in aeternum non commovebitur impii autem non habitabunt in terram
PROV|10|31|os iusti parturiet sapientiam lingua pravorum peribit
PROV|10|32|labia iusti considerant placita et os impiorum perversa
PROV|11|1|statera dolosa abominatio apud Dominum et pondus aequum voluntas eius
PROV|11|2|ubi fuerit superbia ibi erit et contumelia ubi autem humilitas ibi et sapientia
PROV|11|3|simplicitas iustorum diriget eos et subplantatio perversorum vastabit illos
PROV|11|4|non proderunt divitiae in die ultionis iustitia autem liberabit a morte
PROV|11|5|iustitia simplicis diriget viam eius et in impietate sua corruet impius
PROV|11|6|iustitia rectorum liberabit eos et in insidiis suis capientur iniqui
PROV|11|7|mortuo homine impio nulla erit ultra spes et expectatio sollicitorum peribit
PROV|11|8|iustus de angustia liberatus est et tradetur impius pro eo
PROV|11|9|simulator ore decipit amicum suum iusti autem liberabuntur scientia
PROV|11|10|in bonis iustorum exultabit civitas et in perditione impiorum erit laudatio
PROV|11|11|benedictione iustorum exaltabitur civitas et ore impiorum subvertetur
PROV|11|12|qui despicit amicum suum indigens corde est vir autem prudens tacebit
PROV|11|13|qui ambulat fraudulenter revelat arcana qui autem fidelis est animi celat commissum
PROV|11|14|ubi non est gubernator populus corruet salus autem ubi multa consilia
PROV|11|15|adfligetur malo qui fidem facit pro extraneo qui autem cavet laqueos securus erit
PROV|11|16|mulier gratiosa inveniet gloriam et robusti habebunt divitias
PROV|11|17|benefacit animae suae vir misericors qui autem crudelis est et propinquos abicit
PROV|11|18|impius facit opus instabile seminanti autem iustitiam merces fidelis
PROV|11|19|clementia praeparat vitam et sectatio malorum mortem
PROV|11|20|abominabile Domino pravum cor et voluntas eius in his qui simpliciter ambulant
PROV|11|21|manus in manu non erit innocens malus semen autem iustorum salvabitur
PROV|11|22|circulus aureus in naribus suis mulier pulchra et fatua
PROV|11|23|desiderium iustorum omne bonum est praestolatio impiorum furor
PROV|11|24|alii dividunt propria et ditiores fiunt alii rapiunt non sua et semper in egestate sunt
PROV|11|25|anima quae benedicit inpinguabitur et qui inebriat ipse quoque inebriabitur
PROV|11|26|qui abscondit frumenta maledicetur in populis benedictio autem super caput vendentium
PROV|11|27|bene consurgit diluculo qui quaerit bona qui autem investigator malorum est opprimetur ab eis
PROV|11|28|qui confidet in divitiis suis corruet iusti autem quasi virens folium germinabunt
PROV|11|29|qui conturbat domum suam possidebit ventos et qui stultus est serviet sapienti
PROV|11|30|fructus iusti lignum vitae et qui suscipit animas sapiens est
PROV|11|31|si iustus in terra recipit quanto magis impius et peccator
PROV|12|1|qui diligit disciplinam diligit scientiam qui autem odit increpationes insipiens est
PROV|12|2|qui bonus est hauriet a Domino gratiam qui autem confidit cogitationibus suis impie agit
PROV|12|3|non roborabitur homo ex impietate et radix iustorum non commovebitur
PROV|12|4|mulier diligens corona viro suo et putredo in ossibus eius quae confusione res dignas gerit
PROV|12|5|cogitationes iustorum iudicia et consilia impiorum fraudulentia
PROV|12|6|verba impiorum insidiantur sanguini os iustorum liberabit eos
PROV|12|7|verte impios et non erunt domus autem iustorum permanebit
PROV|12|8|doctrina sua noscetur vir qui autem vanus et excors est patebit contemptui
PROV|12|9|melior est pauper et sufficiens sibi quam gloriosus et indigens pane
PROV|12|10|novit iustus animas iumentorum suorum viscera autem impiorum crudelia
PROV|12|11|qui operatur terram suam saturabitur panibus qui autem sectatur otium stultissimus est
PROV|12|12|desiderium impii munimentum est pessimorum radix autem iustorum proficiet
PROV|12|13|propter peccata labiorum ruina proximat malo effugiet autem iustus de angustia
PROV|12|14|de fructu oris sui unusquisque replebitur bonis et iuxta opera manuum suarum retribuetur ei
PROV|12|15|via stulti recta in oculis eius qui autem sapiens est audit consilia
PROV|12|16|fatuus statim indicat iram suam qui autem dissimulat iniuriam callidus est
PROV|12|17|qui quod novit loquitur index iustitiae est qui autem mentitur testis est fraudulentus
PROV|12|18|est qui promittit et quasi gladio pungitur conscientiae lingua autem sapientium sanitas est
PROV|12|19|labium veritatis firmum erit in perpetuum qui autem testis est repentinus concinnat linguam mendacii
PROV|12|20|dolus in corde cogitantium mala qui autem ineunt pacis consilia sequitur eos gaudium
PROV|12|21|non contristabit iustum quicquid ei acciderit impii autem replebuntur malo
PROV|12|22|abominatio Domino labia mendacia qui autem fideliter agunt placent ei
PROV|12|23|homo versutus celat scientiam et cor insipientium provocabit stultitiam
PROV|12|24|manus fortium dominabitur quae autem remissa est tributis serviet
PROV|12|25|maeror in corde viri humiliabit illud et sermone bono laetificabitur
PROV|12|26|qui neglegit damnum propter amicum iustus est iter autem impiorum decipiet eos
PROV|12|27|non inveniet fraudulentus lucrum et substantia hominis erit auri pretium
PROV|12|28|in semita iustitiae vita iter autem devium ducit ad mortem
PROV|13|1|filius sapiens doctrina patris qui autem inlusor est non audit cum arguitur
PROV|13|2|de fructu oris homo saturabitur bonis anima autem praevaricatorum iniqua
PROV|13|3|qui custodit os suum custodit animam suam qui autem inconsideratus est ad loquendum sentiet mala
PROV|13|4|vult et non vult piger anima autem operantium inpinguabitur
PROV|13|5|verbum mendax iustus detestabitur impius confundit et confundetur
PROV|13|6|iustitia custodit innocentis viam impietas vero peccato subplantat
PROV|13|7|est quasi dives cum nihil habeat et est quasi pauper cum in multis divitiis sit
PROV|13|8|redemptio animae viri divitiae suae qui autem pauper est increpationem non sustinet
PROV|13|9|lux iustorum laetificat lucerna autem impiorum extinguetur
PROV|13|10|inter superbos semper iurgia sunt qui autem agunt cuncta consilio reguntur sapientia
PROV|13|11|substantia festinata minuetur quae autem paulatim colligitur manu multiplicabitur
PROV|13|12|spes quae differtur adfligit animam lignum vitae desiderium veniens
PROV|13|13|qui detrahit alicui rei ipse se in futurum obligat qui autem timet praeceptum in pace versabitur
PROV|13|14|lex sapientis fons vitae ut declinet a ruina mortis
PROV|13|15|doctrina bona dabit gratiam in itinere contemptorum vorago
PROV|13|16|astutus omnia agit cum consilio qui autem fatuus est aperit stultitiam
PROV|13|17|nuntius impii cadet in malum legatus fidelis sanitas
PROV|13|18|egestas et ignominia ei qui deserit disciplinam qui autem adquiescit arguenti glorificabitur
PROV|13|19|desiderium si conpleatur delectat animam detestantur stulti eos qui fugiunt mala
PROV|13|20|qui cum sapientibus graditur sapiens erit amicus stultorum efficietur similis
PROV|13|21|peccatores persequetur malum et iustis retribuentur bona
PROV|13|22|bonus relinquet heredes filios et nepotes et custoditur iusto substantia peccatoris
PROV|13|23|multi cibi in novalibus patrum et alii congregantur absque iudicio
PROV|13|24|qui parcit virgae suae odit filium suum qui autem diligit illum instanter erudit
PROV|13|25|iustus comedit et replet animam suam venter autem impiorum insaturabilis
PROV|14|1|sapiens mulier aedificavit domum suam insipiens instructam quoque destruet manibus
PROV|14|2|ambulans recto itinere et timens Deum despicitur ab eo qui infami graditur via
PROV|14|3|in ore stulti virga superbiae labia sapientium custodiunt eos
PROV|14|4|ubi non sunt boves praesepe vacuum est ubi autem plurimae segetes ibi manifesta fortitudo bovis
PROV|14|5|testis fidelis non mentietur profert mendacium testis dolosus
PROV|14|6|quaerit derisor sapientiam et non inveniet doctrina prudentium facilis
PROV|14|7|vade contra virum stultum et nescito labia prudentiae
PROV|14|8|sapientia callidi est intellegere viam suam et inprudentia stultorum errans
PROV|14|9|stultis inludet peccatum inter iustos morabitur gratia
PROV|14|10|cor quod novit amaritudinem animae suae in gaudio eius non miscebitur extraneus
PROV|14|11|domus impiorum delebitur tabernacula iustorum germinabunt
PROV|14|12|est via quae videtur homini iusta novissima autem eius deducunt ad mortem
PROV|14|13|risus dolore miscebitur et extrema gaudii luctus occupat
PROV|14|14|viis suis replebitur stultus et super eum erit vir bonus
PROV|14|15|innocens credit omni verbo astutus considerat gressus suos
PROV|14|16|sapiens timet et declinat malum stultus transilit et confidit
PROV|14|17|inpatiens operabitur stultitiam et vir versutus odiosus est
PROV|14|18|possidebunt parvuli stultitiam et astuti expectabunt scientiam
PROV|14|19|iacebunt mali ante bonos et impii ante portas iustorum
PROV|14|20|etiam proximo suo pauper odiosus erit amici vero divitum multi
PROV|14|21|qui despicit proximum suum peccat qui autem miseretur pauperi beatus erit
PROV|14|22|errant qui operantur malum misericordia et veritas praeparant bona
PROV|14|23|in omni opere erit abundantia ubi autem verba sunt plurima frequenter egestas
PROV|14|24|corona sapientium divitiae eorum fatuitas stultorum inprudentia
PROV|14|25|liberat animas testis fidelis et profert mendacia versipellis
PROV|14|26|in timore Domini fiducia fortitudinis et filiis eius erit spes
PROV|14|27|timor Domini fons vitae ut declinet a ruina mortis
PROV|14|28|in multitudine populi dignitas regis et in paucitate plebis ignominia principis
PROV|14|29|qui patiens est multa gubernatur prudentia qui autem inpatiens exaltat stultitiam suam
PROV|14|30|vita carnium sanitas cordis putredo ossuum invidia
PROV|14|31|qui calumniatur egentem exprobrat factori eius honorat autem eum qui miseretur pauperis
PROV|14|32|in malitia sua expelletur impius sperat autem iustus in morte sua
PROV|14|33|in corde prudentis requiescit sapientia et indoctos quoque erudiet
PROV|14|34|iustitia elevat gentem miseros facit populos peccatum
PROV|14|35|acceptus est regi minister intellegens iracundiam eius inutilis sustinebit
PROV|15|1|responsio mollis frangit iram sermo durus suscitat furorem
PROV|15|2|lingua sapientium ornat scientiam os fatuorum ebullit stultitiam
PROV|15|3|in omni loco oculi Domini contemplantur malos et bonos
PROV|15|4|lingua placabilis lignum vitae quae inmoderata est conteret spiritum
PROV|15|5|stultus inridet disciplinam patris sui qui autem custodit increpationes astutior fiet
PROV|15|6|domus iusti plurima fortitudo et in fructibus impii conturbatur
PROV|15|7|labia sapientium disseminabunt scientiam cor stultorum dissimile erit
PROV|15|8|victimae impiorum abominabiles Domino vota iustorum placabilia
PROV|15|9|abominatio est Domino via impii qui sequitur iustitiam diligetur ab eo
PROV|15|10|doctrina mala deserenti viam qui increpationes odit morietur
PROV|15|11|infernus et perditio coram Domino quanto magis corda filiorum hominum
PROV|15|12|non amat pestilens eum qui se corripit nec ad sapientes graditur
PROV|15|13|cor gaudens exhilarat faciem in maerore animi deicitur spiritus
PROV|15|14|cor sapientis quaerit doctrinam et os stultorum pascetur inperitia
PROV|15|15|omnes dies pauperis mali secura mens quasi iuge convivium
PROV|15|16|melius est parum cum timore Domini quam thesauri magni et insatiabiles
PROV|15|17|melius est vocare ad holera cum caritate quam ad vitulum saginatum cum odio
PROV|15|18|vir iracundus provocat rixas qui patiens est mitigat suscitatas
PROV|15|19|iter pigrorum quasi sepes spinarum via iustorum absque offendiculo
PROV|15|20|filius sapiens laetificat patrem et stultus homo despicit matrem suam
PROV|15|21|stultitia gaudium stulto et vir prudens dirigit gressus
PROV|15|22|dissipantur cogitationes ubi non est consilium ubi vero plures sunt consiliarii confirmantur
PROV|15|23|laetatur homo in sententia oris sui et sermo oportunus est optimus
PROV|15|24|semita vitae super eruditum ut declinet de inferno novissimo
PROV|15|25|domum superborum demolietur Dominus et firmos facit terminos viduae
PROV|15|26|abominatio Domini cogitationes malae et purus sermo pulcherrimus
PROV|15|27|conturbat domum suam qui sectatur avaritiam qui autem odit munera vivet
PROV|15|28|mens iusti meditatur oboedientiam os impiorum redundat malis
PROV|15|29|longe est Dominus ab impiis et orationes iustorum exaudiet
PROV|15|30|lux oculorum laetificat animam fama bona inpinguat ossa
PROV|15|31|auris quae audit increpationes vitae in medio sapientium commorabitur
PROV|15|32|qui abicit disciplinam despicit animam suam qui adquiescit increpationibus possessor est cordis
PROV|15|33|timor Domini disciplina sapientiae et gloriam praecedit humilitas
PROV|16|1|hominis est animum praeparare et Dei gubernare linguam
PROV|16|2|omnes viae hominum patent oculis eius spirituum ponderator est Dominus
PROV|16|3|revela Domino opera tua et dirigentur cogitationes tuae
PROV|16|4|universa propter semet ipsum operatus est Dominus impium quoque ad diem malum
PROV|16|5|abominatio Domini omnis arrogans etiam si manus ad manum fuerit non erit innocens
PROV|16|6|misericordia et veritate redimitur iniquitas et in timore Domini declinatur a malo
PROV|16|7|cum placuerint Domino viae hominis inimicos quoque eius convertet ad pacem
PROV|16|8|melius est parum cum iustitia quam multi fructus cum iniquitate
PROV|16|9|cor hominis disponet viam suam sed Domini est dirigere gressus eius
PROV|16|10|divinatio in labiis regis in iudicio non errabit os eius
PROV|16|11|pondus et statera iudicia Domini sunt et opera eius omnes lapides sacculi
PROV|16|12|abominabiles regi qui agunt impie quoniam iustitia firmatur solium
PROV|16|13|voluntas regum labia iusta qui recta loquitur diligetur
PROV|16|14|indignatio regis nuntii mortis et vir sapiens placabit eam
PROV|16|15|in hilaritate vultus regis vita et clementia eius quasi imber serotinus
PROV|16|16|posside sapientiam quia auro melior est et adquire prudentiam quia pretiosior est argento
PROV|16|17|semita iustorum declinat mala custos animae suae servat viam suam
PROV|16|18|contritionem praecedit superbia et ante ruinam exaltatur spiritus
PROV|16|19|melius est humiliari cum mitibus quam dividere spolia cum superbis
PROV|16|20|eruditus in verbo repperiet bona et qui in Domino sperat beatus est
PROV|16|21|qui sapiens corde est appellabitur prudens et qui dulcis eloquio maiora percipiet
PROV|16|22|fons vitae eruditio possidentis doctrina stultorum fatuitas
PROV|16|23|cor sapientis erudiet os eius et labiis illius addet gratiam
PROV|16|24|favus mellis verba conposita dulcedo animae et sanitas ossuum
PROV|16|25|est via quae videtur homini recta et novissimum eius ducit ad mortem
PROV|16|26|anima laborantis laborat sibi quia conpulit eum os suum
PROV|16|27|vir impius fodit malum et in labiis eius ignis ardescit
PROV|16|28|homo perversus suscitat lites et verbosus separat principes
PROV|16|29|vir iniquus lactat amicum suum et ducit eum per viam non bonam
PROV|16|30|qui adtonitis oculis cogitat prava mordens labia sua perficit malum
PROV|16|31|corona dignitatis senectus in viis iustitiae repperietur
PROV|16|32|melior est patiens viro forte et qui dominatur animo suo expugnatore urbium
PROV|16|33|sortes mittuntur in sinu sed a Domino temperantur
PROV|17|1|melior est buccella sicca cum gaudio quam domus plena victimis cum iurgio
PROV|17|2|servus sapiens dominabitur filiis stultis et inter fratres hereditatem dividet
PROV|17|3|sicut igne probatur argentum et aurum camino ita corda probat Dominus
PROV|17|4|malus oboedit linguae iniquae et fallax obtemperat labiis mendacibus
PROV|17|5|qui despicit pauperem exprobrat factori eius et qui in ruina laetatur alterius non erit inpunitus
PROV|17|6|corona senum filii filiorum et gloria filiorum patres sui
PROV|17|7|non decent stultum verba conposita nec principem labium mentiens
PROV|17|8|gemma gratissima expectatio praestolantis quocumque se verterit prudenter intellegit
PROV|17|9|qui celat delictum quaerit amicitias qui altero sermone repetit separat foederatos
PROV|17|10|plus proficit correptio apud prudentem quam centum plagae apud stultum
PROV|17|11|semper iurgia quaerit malus angelus autem crudelis mittetur contra eum
PROV|17|12|expedit magis ursae occurrere raptis fetibus quam fatuo confidenti sibi in stultitia sua
PROV|17|13|qui reddit mala pro bonis non recedet malum de domo eius
PROV|17|14|qui dimittit aquam caput est iurgiorum et antequam patiatur contumeliam iudicium deserit
PROV|17|15|et qui iustificat impium et qui condemnat iustum abominabilis est uterque apud Dominum
PROV|17|16|quid prodest habere divitias stultum cum sapientiam emere non possit
PROV|17|17|omni tempore diligit qui amicus est et frater in angustiis conprobatur
PROV|17|18|homo stultus plaudet manibus cum spoponderit pro amico suo
PROV|17|19|qui meditatur discordiam diligit rixas et qui exaltat ostium quaerit ruinam
PROV|17|20|qui perversi cordis est non inveniet bonum et qui vertit linguam incidet in malum
PROV|17|21|natus est stultus in ignominiam suam sed nec pater in fatuo laetabitur
PROV|17|22|animus gaudens aetatem floridam facit spiritus tristis exsiccat ossa
PROV|17|23|munera de sinu impius accipit ut pervertat semitas iudicii
PROV|17|24|in facie prudentis lucet sapientia oculi stultorum in finibus terrae
PROV|17|25|ira patris filius stultus et dolor matris quae genuit eum
PROV|17|26|non est bonum damnum inferre iusto nec percutere principem qui recta iudicat
PROV|17|27|qui moderatur sermones suos doctus et prudens est et pretiosi spiritus vir eruditus
PROV|17|28|stultus quoque si tacuerit sapiens putabitur et si conpresserit labia sua intellegens
PROV|18|1|occasiones quaerit qui vult recedere ab amico omni tempore erit exprobrabilis
PROV|18|2|non recipit stultus verba prudentiae nisi ea dixeris quae versantur in corde eius
PROV|18|3|impius cum in profundum venerit peccatorum contemnit sed sequitur eum ignominia et obprobrium
PROV|18|4|aqua profunda verba ex ore viri et torrens redundans fons sapientiae
PROV|18|5|accipere personam impii non est bonum ut declines a veritate iudicii
PROV|18|6|labia stulti inmiscunt se rixis et os eius iurgia provocat
PROV|18|7|os stulti contritio eius et labia illius ruina animae eius
PROV|18|8|verba bilinguis quasi simplicia et ipsa perveniunt usque ad interiora ventris
PROV|18|9|qui mollis et dissolutus est in opere suo frater est sua opera dissipantis
PROV|18|10|turris fortissima nomen Domini ad ipsum currit iustus et exaltabitur
PROV|18|11|substantia divitis urbs roboris eius et quasi murus validus circumdans eum
PROV|18|12|antequam conteratur exaltatur cor hominis et antequam glorificetur humiliatur
PROV|18|13|qui prius respondit quam audiat stultum se esse demonstrat et confusione dignum
PROV|18|14|spiritus viri sustentat inbecillitatem suam spiritum vero ad irascendum facilem quis poterit sustinere
PROV|18|15|cor prudens possidebit scientiam et auris sapientium quaerit doctrinam
PROV|18|16|donum hominis dilatat viam eius et ante principes spatium ei facit
PROV|18|17|iustus prior est accusator sui venit amicus eius et investigavit eum
PROV|18|18|contradictiones conprimit sors et inter potentes quoque diiudicat
PROV|18|19|frater qui adiuvatur a fratre quasi civitas firma et iudicia quasi vectes urbium
PROV|18|20|de fructu oris viri replebitur venter eius et genimina labiorum illius saturabunt eum
PROV|18|21|mors et vita in manu linguae qui diligunt eam comedent fructus eius
PROV|18|22|qui invenit mulierem invenit bonum et hauriet iucunditatem a Domino
PROV|18|23|cum obsecrationibus loquetur pauper et dives effabitur rigide
PROV|18|24|vir amicalis ad societatem magis amicus erit quam frater
PROV|19|1|melior est pauper qui ambulat in simplicitate sua quam torquens labia insipiens
PROV|19|2|ubi non est scientia animae non est bonum et qui festinus est pedibus offendit
PROV|19|3|stultitia hominis subplantat gressus eius et contra Deum fervet animo suo
PROV|19|4|divitiae addunt amicos plurimos a paupere autem et hii quos habuit separantur
PROV|19|5|testis falsus non erit inpunitus et qui mendacia loquitur non effugiet
PROV|19|6|multi colunt personam potentis et amici sunt dona tribuenti
PROV|19|7|fratres hominis pauperis oderunt eum insuper et amici procul recesserunt ab eo qui tantum verba sectatur nihil habebit
PROV|19|8|qui autem possessor est mentis diligit animam suam et custos prudentiae inveniet bona
PROV|19|9|testis falsus non erit inpunitus et qui loquitur mendacia peribit
PROV|19|10|non decent stultum deliciae nec servum dominari principibus
PROV|19|11|doctrina viri per patientiam noscitur et gloria eius est iniqua praetergredi
PROV|19|12|sicut fremitus leonis ita et regis ira et sicut ros super herbam ita hilaritas eius
PROV|19|13|dolor patris filius stultus et tecta iugiter perstillantia litigiosa mulier
PROV|19|14|domus et divitiae dantur a patribus a Domino autem proprie uxor prudens
PROV|19|15|pigredo inmittit soporem et anima dissoluta esuriet
PROV|19|16|qui custodit mandatum custodit animam suam qui autem neglegit vias suas mortificabitur
PROV|19|17|feneratur Domino qui miseretur pauperis et vicissitudinem suam reddet ei
PROV|19|18|erudi filium tuum ne desperes ad interfectionem autem eius ne ponas animam tuam
PROV|19|19|qui inpatiens est sustinebit damnum et cum rapuerit aliud adponet
PROV|19|20|audi consilium et suscipe disciplinam ut sis sapiens in novissimis tuis
PROV|19|21|multae cogitationes in corde viri voluntas autem Domini permanebit
PROV|19|22|homo indigens misericors est et melior pauper quam vir mendax
PROV|19|23|timor Domini ad vitam et in plenitudine commorabitur absque visitatione pessimi
PROV|19|24|abscondit piger manum suam sub ascella nec ad os suum adplicat eam
PROV|19|25|pestilente flagellato stultus sapientior erit sin autem corripueris sapientem intelleget disciplinam
PROV|19|26|qui adfligit patrem et fugat matrem ignominiosus est et infelix
PROV|19|27|non cesses fili audire doctrinam nec ignores sermones scientiae
PROV|19|28|testis iniquus deridet iudicium et os impiorum devorat iniquitatem
PROV|19|29|parata sunt derisoribus iudicia et mallei percutientes stultorum corporibus
PROV|20|1|luxuriosa res vinum et tumultuosa ebrietas quicumque his delectatur non erit sapiens
PROV|20|2|sicut rugitus leonis ita terror regis qui provocat eum peccat in animam suam
PROV|20|3|honor est homini qui separat se a contentionibus omnes autem stulti miscentur contumeliis
PROV|20|4|propter frigus piger arare noluit mendicabit ergo aestate et non dabitur ei
PROV|20|5|sicut aqua profunda sic consilium in corde viri sed homo sapiens exhauriet illud
PROV|20|6|multi homines misericordes vocantur virum autem fidelem quis inveniet
PROV|20|7|iustus qui ambulat in simplicitate sua beatos post se filios derelinquet
PROV|20|8|rex qui sedet in solio iudicii dissipat omne malum intuitu suo
PROV|20|9|quis potest dicere mundum est cor meum purus sum a peccato
PROV|20|10|pondus et pondus mensura et mensura utrumque abominabile est apud Deum
PROV|20|11|ex studiis suis intellegitur puer si munda et si recta sint opera eius
PROV|20|12|aurem audientem et oculum videntem Dominus fecit utrumque
PROV|20|13|noli diligere somnum ne te egestas opprimat aperi oculos tuos et saturare panibus
PROV|20|14|malum est malum est dicit omnis emptor et cum recesserit tunc gloriabitur
PROV|20|15|est aurum et multitudo gemmarum vas autem pretiosum labia scientiae
PROV|20|16|tolle vestimentum eius qui fideiussor extitit alieni et pro extraneis aufer pignus ab eo
PROV|20|17|suavis est homini panis mendacii et postea implebitur os eius calculo
PROV|20|18|cogitationes consiliis roborantur et gubernaculis tractanda sunt bella
PROV|20|19|ei qui revelat mysteria et ambulat fraudulenter et dilatat labia sua ne commiscearis
PROV|20|20|qui maledicit patri suo et matri extinguetur lucerna eius in mediis tenebris
PROV|20|21|hereditas ad quam festinatur in principio in novissimo benedictione carebit
PROV|20|22|ne dicas reddam malum expecta Dominum et liberabit te
PROV|20|23|abominatio est apud Deum pondus et pondus statera dolosa non est bona
PROV|20|24|a Domino diriguntur gressus viri quis autem hominum intellegere potest viam suam
PROV|20|25|ruina est hominis devorare sanctos et post vota tractare
PROV|20|26|dissipat impios rex sapiens et curvat super eos fornicem
PROV|20|27|lucerna Domini spiraculum hominis quae investigat omnia secreta ventris
PROV|20|28|misericordia et veritas custodiunt regem et roboratur clementia thronus eius
PROV|20|29|exultatio iuvenum fortitudo eorum et dignitas senum canities
PROV|20|30|livor vulneris absterget mala et plagae in secretioribus ventris
PROV|21|1|sicut divisiones aquarum ita cor regis in manu Domini quocumque voluerit inclinabit illud
PROV|21|2|omnis via viri recta sibi videtur adpendit autem corda Dominus
PROV|21|3|facere misericordiam et iudicium magis placent Domino quam victimae
PROV|21|4|exaltatio oculorum et dilatatio cordis lucerna impiorum peccatum
PROV|21|5|cogitationes robusti semper in abundantia omnis autem piger semper in egestate
PROV|21|6|qui congregat thesauros lingua mendacii vanus est et inpingetur ad laqueos mortis
PROV|21|7|rapinae impiorum detrahent eos quia noluerunt facere iudicium
PROV|21|8|perversa via viri aliena est qui autem mundus est rectum opus eius
PROV|21|9|melius est sedere in angulo domatis quam cum muliere litigiosa et in domo communi
PROV|21|10|anima impii desiderat malum non miserebitur proximo suo
PROV|21|11|multato pestilente sapientior erit parvulus et si sectetur sapientem sumet scientiam
PROV|21|12|excogitat iustus de domo impii ut detrahat impios in malum
PROV|21|13|qui obturat aurem suam ad clamorem pauperis et ipse clamabit et non exaudietur
PROV|21|14|munus absconditum extinguet iras et donum in sinu indignationem maximam
PROV|21|15|gaudium iusto est facere iudicium et pavor operantibus iniquitatem
PROV|21|16|vir qui erraverit a via doctrinae in coetu gigantum commorabitur
PROV|21|17|qui diligit epulas in egestate erit qui amat vinum et pinguia non ditabitur
PROV|21|18|pro iusto datur impius et pro rectis iniquus
PROV|21|19|melius est habitare in terra deserta quam cum muliere rixosa et iracunda
PROV|21|20|thesaurus desiderabilis et oleum in habitaculo iusti et inprudens homo dissipabit illud
PROV|21|21|qui sequitur iustitiam et misericordiam inveniet vitam et iustitiam et gloriam
PROV|21|22|civitatem fortium ascendit sapiens et destruxit robur fiduciae eius
PROV|21|23|qui custodit os suum et linguam suam custodit ab angustiis animam suam
PROV|21|24|superbus et arrogans vocatur indoctus qui in ira operatur superbiam
PROV|21|25|desideria occidunt pigrum noluerunt enim quicquam manus eius operari
PROV|21|26|tota die concupiscit et desiderat qui autem iustus est tribuet et non cessabit
PROV|21|27|hostiae impiorum abominabiles quia offeruntur ex scelere
PROV|21|28|testis mendax peribit vir oboediens loquitur victoriam
PROV|21|29|vir impius procaciter obfirmat vultum suum qui autem rectus est corrigit viam suam
PROV|21|30|non est sapientia non est prudentia non est consilium contra Dominum
PROV|21|31|equus paratur ad diem belli Dominus autem salutem tribuet
PROV|22|1|melius est nomen bonum quam divitiae multae super argentum et aurum gratia bona
PROV|22|2|dives et pauper obviaverunt sibi utriusque operator est Dominus
PROV|22|3|callidus vidit malum et abscondit se innocens pertransiit et adflictus est damno
PROV|22|4|finis modestiae timor Domini divitiae et gloria et vita
PROV|22|5|arma et gladii in via perversi custos animae suae longe recedit ab eis
PROV|22|6|proverbium est adulescens iuxta viam suam etiam cum senuerit non recedet ab ea
PROV|22|7|dives pauperibus imperat et qui accipit mutuum servus est fenerantis
PROV|22|8|qui seminat iniquitatem metet mala et virga irae suae consummabitur
PROV|22|9|qui pronus est ad misericordiam benedicetur de panibus enim suis dedit pauperi
PROV|22|10|eice derisorem et exibit cum eo iurgium cessabuntque causae et contumeliae
PROV|22|11|qui diligit cordis munditiam propter gratiam labiorum suorum habebit amicum regem
PROV|22|12|oculi Domini custodiunt scientiam et subplantantur verba iniqui
PROV|22|13|dicit piger leo foris in medio platearum occidendus sum
PROV|22|14|fovea profunda os alienae cui iratus est Dominus incidet in eam
PROV|22|15|stultitia conligata est in corde pueri et virga disciplinae fugabit eam
PROV|22|16|qui calumniatur pauperem ut augeat divitias suas dabit ipse ditiori et egebit
PROV|22|17|inclina aurem tuam et audi verba sapientium adpone autem cor ad doctrinam meam
PROV|22|18|quae pulchra erit tibi cum servaveris eam in ventre tuo et redundabit in labiis tuis
PROV|22|19|ut sit in Domino fiducia tua unde et ostendi eam tibi hodie
PROV|22|20|ecce descripsi eam tibi tripliciter in cogitationibus et scientia
PROV|22|21|ut ostenderem tibi firmitatem et eloquia veritatis respondere ex his illi qui misit te
PROV|22|22|non facias violentiam pauperi quia pauper est neque conteras egenum in porta
PROV|22|23|quia Dominus iudicabit causam eius et configet eos qui confixerint animam eius
PROV|22|24|noli esse amicus homini iracundo neque ambules cum viro furioso
PROV|22|25|ne forte discas semitas eius et sumas scandalum animae tuae
PROV|22|26|noli esse cum his qui defigunt manus suas et qui vades se offerunt pro debitis
PROV|22|27|si enim non habes unde restituas quid causae est ut tollat operimentum de cubili tuo
PROV|22|28|ne transgrediaris terminos antiquos quos posuerunt patres tui
PROV|22|29|vidisti virum velocem in opere suo coram regibus stabit nec erit ante ignobiles
PROV|23|1|quando sederis ut comedas cum principe diligenter adtende quae posita sunt ante faciem tuam
PROV|23|2|et statue cultrum in gutture tuo si tamen habes in potestate animam tuam
PROV|23|3|ne desideres de cibis eius in quo est panis mendacii
PROV|23|4|noli laborare ut diteris sed prudentiae tuae pone modum
PROV|23|5|ne erigas oculos tuos ad opes quas habere non potes quia facient sibi pinnas quasi aquilae et avolabunt in caelum
PROV|23|6|ne comedas cum homine invido et ne desideres cibos eius
PROV|23|7|quoniam in similitudinem arioli et coniectoris aestimat quod ignorat comede et bibe dicet tibi et mens eius non est tecum
PROV|23|8|cibos quos comederas evomes et perdes pulchros sermones tuos
PROV|23|9|in auribus insipientium ne loquaris quia despicient doctrinam eloquii tui
PROV|23|10|ne adtingas terminos parvulorum et agrum pupillorum ne introeas
PROV|23|11|propinquus enim eorum Fortis est et ipse iudicabit contra te causam illorum
PROV|23|12|ingrediatur ad doctrinam cor tuum et aures tuae ad verba scientiae
PROV|23|13|noli subtrahere a puero disciplinam si enim percusseris eum virga non morietur
PROV|23|14|tu virga percuties eum et animam eius de inferno liberabis
PROV|23|15|fili mi si sapiens fuerit animus tuus gaudebit tecum cor meum
PROV|23|16|et exultabunt renes mei cum locuta fuerint rectum labia tua
PROV|23|17|non aemuletur cor tuum peccatores sed in timore Domini esto tota die
PROV|23|18|quia habebis spem in novissimo et praestolatio tua non auferetur
PROV|23|19|audi fili mi et esto sapiens et dirige in via animum tuum
PROV|23|20|noli esse in conviviis potatorum nec in comesationibus eorum qui carnes ad vescendum conferunt
PROV|23|21|quia vacantes potibus et dantes symbola consumentur et vestietur pannis dormitatio
PROV|23|22|audi patrem tuum qui genuit te et ne contemnas cum senuerit mater tua
PROV|23|23|veritatem eme et noli vendere sapientiam et doctrinam et intellegentiam
PROV|23|24|exultat gaudio pater iusti qui sapientem genuit laetabitur in eo
PROV|23|25|gaudeat pater tuus et mater tua et exultet quae genuit te
PROV|23|26|praebe fili mi cor tuum mihi et oculi tui vias meas custodiant
PROV|23|27|fovea enim profunda est meretrix et puteus angustus aliena
PROV|23|28|insidiatur in via quasi latro et quos incautos viderit interficit
PROV|23|29|cui vae cuius patri vae cui rixae cui foveae cui sine causa vulnera cui suffusio oculorum
PROV|23|30|nonne his qui morantur in vino et student calicibus epotandis
PROV|23|31|ne intuearis vinum quando flavescit cum splenduerit in vitro color eius ingreditur blande
PROV|23|32|sed in novissimo mordebit ut coluber et sicut regulus venena diffundet
PROV|23|33|oculi tui videbunt extraneas et cor tuum loquetur perversa
PROV|23|34|et eris sicut dormiens in medio mari et quasi sopitus gubernator amisso clavo
PROV|23|35|et dices verberaverunt me sed non dolui traxerunt me et ego non sensi quando evigilabo et rursum vina repperiam
PROV|24|1|ne aemuleris viros malos nec desideres esse cum eis
PROV|24|2|quia rapinas meditatur mens eorum et fraudes labia eorum loquuntur
PROV|24|3|sapientia aedificabitur domus et prudentia roborabitur
PROV|24|4|in doctrina replebuntur cellaria universa substantia pretiosa et pulcherrima
PROV|24|5|vir sapiens et fortis est et vir doctus robustus et validus
PROV|24|6|quia cum dispositione initur bellum et erit salus ubi multa consilia sunt
PROV|24|7|excelsa stulto sapientia in porta non aperiet os suum
PROV|24|8|qui cogitat malefacere stultus vocabitur
PROV|24|9|cogitatio stulti peccatum est et abominatio hominum detractor
PROV|24|10|si desperaveris lassus in die angustiae inminuetur fortitudo tua
PROV|24|11|erue eos qui ducuntur ad mortem et qui trahuntur ad interitum liberare ne cesses
PROV|24|12|si dixeris vires non suppetunt qui inspector est cordis ipse intellegit et servatorem animae tuae nihil fallit reddetque homini iuxta opera sua
PROV|24|13|comede fili mi mel quia bonum est et favum dulcissimum gutturi tuo
PROV|24|14|sic et doctrina sapientiae animae tuae quam cum inveneris habebis in novissimis et spes tua non peribit
PROV|24|15|ne insidieris et quaeras impietatem in domo iusti neque vastes requiem eius
PROV|24|16|septies enim cadet iustus et resurget impii autem corruent in malum
PROV|24|17|cum ceciderit inimicus tuus ne gaudeas et in ruina eius ne exultet cor tuum
PROV|24|18|ne forte videat Dominus et displiceat ei et auferat ab eo iram suam
PROV|24|19|ne contendas cum pessimis nec aemuleris impios
PROV|24|20|quoniam non habent futurorum spem mali et lucerna impiorum extinguetur
PROV|24|21|time Dominum fili mi et regem et cum detractoribus non commiscearis
PROV|24|22|quoniam repente consurget perditio eorum et ruinam utriusque quis novit
PROV|24|23|haec quoque sapientibus cognoscere personam in iudicio non est bonum
PROV|24|24|qui dicit impio iustus es maledicent ei populi et detestabuntur eum tribus
PROV|24|25|qui arguunt laudabuntur et super ipsos veniet benedictio
PROV|24|26|labia deosculabitur qui recta verba respondet
PROV|24|27|praepara foris opus tuum et diligenter exerce agrum tuum ut postea aedifices domum tuam
PROV|24|28|ne sis testis frustra contra proximum tuum nec lactes quemquam labiis tuis
PROV|24|29|ne dicas quomodo fecit mihi sic faciam ei reddam unicuique secundum opus suum
PROV|24|30|per agrum hominis pigri transivi et per vineam viri stulti
PROV|24|31|et ecce totum repleverant urticae operuerant superficiem eius spinae et maceria lapidum destructa erat
PROV|24|32|quod cum vidissem posui in corde meo et exemplo didici disciplinam
PROV|24|33|parum inquam dormies modicum dormitabis pauxillum manus conseres ut quiescas
PROV|24|34|et veniet quasi cursor egestas tua et mendicitas quasi vir armatus
PROV|25|1|haec quoque parabolae Salomonis quas transtulerunt viri Ezechiae regis Iuda
PROV|25|2|gloria Dei celare verbum et gloria regum investigare sermonem
PROV|25|3|caelum sursum et terra deorsum et cor regum inscrutabile
PROV|25|4|aufer robiginem de argento et egredietur vas purissimum
PROV|25|5|aufer impietatem de vultu regis et firmabitur iustitia thronus eius
PROV|25|6|ne gloriosus appareas coram rege et in loco magnorum ne steteris
PROV|25|7|melius est enim ut dicatur tibi ascende huc quam ut humilieris coram principe
PROV|25|8|quae viderunt oculi tui ne proferas in iurgio cito ne postea emendare non possis cum dehonestaveris amicum tuum
PROV|25|9|causam tuam tracta cum amico tuo et secretum extraneo non reveles
PROV|25|10|ne forte insultet tibi cum audierit et exprobrare non cesset
PROV|25|11|mala aurea in lectis argenteis qui loquitur verbum in tempore suo
PROV|25|12|inauris aurea et margaritum fulgens qui arguit sapientem et aurem oboedientem
PROV|25|13|sicut frigus nivis in die messis ita legatus fidelis ei qui misit eum animam illius requiescere facit
PROV|25|14|nubes et ventus et pluviae non sequentes vir gloriosus et promissa non conplens
PROV|25|15|patientia lenietur princeps et lingua mollis confringet duritiam
PROV|25|16|mel invenisti comede quod sufficit tibi ne forte saturatus evomas illud
PROV|25|17|subtrahe pedem tuum de domo proximi tui nequando satiatus oderit te
PROV|25|18|iaculum et gladius et sagitta acuta homo qui loquitur contra proximum suum testimonium falsum
PROV|25|19|dens putridus et pes lapsus qui sperat super infideli in die angustiae
PROV|25|20|et amittit pallium in die frigoris acetum in nitro et qui cantat carmina cordi pessimo
PROV|25|21|si esurierit inimicus tuus ciba illum et si sitierit da ei aquam bibere
PROV|25|22|prunam enim congregabis super caput eius et Dominus reddet tibi
PROV|25|23|ventus aquilo dissipat pluvias et facies tristis linguam detrahentem
PROV|25|24|melius est sedere in angulo domatis quam cum muliere litigiosa et in domo communi
PROV|25|25|aqua frigida animae sitienti et nuntius bonus de terra longinqua
PROV|25|26|fons turbatus pede et vena corrupta iustus cadens coram impio
PROV|25|27|sicut qui mel multum comedit non est ei bonum sic qui scrutator est maiestatis opprimitur gloria
PROV|25|28|sicut urbs patens et absque murorum ambitu ita vir qui non potest in loquendo cohibere spiritum suum
PROV|26|1|quomodo nix aestate et pluvia in messe sic indecens est stulto gloria
PROV|26|2|sicut avis ad alia transvolans et passer quolibet vadens sic maledictum frustra prolatum in quempiam superveniet
PROV|26|3|flagellum equo et camus asino et virga dorso inprudentium
PROV|26|4|ne respondeas stulto iuxta stultitiam suam ne efficiaris ei similis
PROV|26|5|responde stulto iuxta stultitiam suam ne sibi sapiens esse videatur
PROV|26|6|claudus pedibus et iniquitatem bibens qui mittit verba per nuntium stultum
PROV|26|7|quomodo pulchras frustra habet claudus tibias sic indecens est in ore stultorum parabola
PROV|26|8|sicut qui mittit lapidem in acervum Mercurii ita qui tribuit insipienti honorem
PROV|26|9|quomodo si spina nascatur in manu temulenti sic parabola in ore stultorum
PROV|26|10|iudicium determinat causas et qui inponit stulto silentium iras mitigat
PROV|26|11|sicut canis qui revertitur ad vomitum suum sic inprudens qui iterat stultitiam suam
PROV|26|12|vidisti hominem sapientem sibi videri magis illo spem habebit stultus
PROV|26|13|dicit piger leaena in via leo in itineribus
PROV|26|14|sicut ostium vertitur in cardine suo ita piger in lectulo suo
PROV|26|15|abscondit piger manus sub ascellas suas et laborat si ad os suum eas converterit
PROV|26|16|sapientior sibi piger videtur septem viris loquentibus sententias
PROV|26|17|sicut qui adprehendit auribus canem sic qui transit et inpatiens commiscetur rixae alterius
PROV|26|18|sicut noxius est qui mittit lanceas et sagittas et mortem
PROV|26|19|sic vir qui fraudulenter nocet amico suo et cum fuerit deprehensus dicit ludens feci
PROV|26|20|cum defecerint ligna extinguetur ignis et susurrone subtracto iurgia conquiescunt
PROV|26|21|sicut carbones ad prunam et ligna ad ignem sic homo iracundus suscitat rixas
PROV|26|22|verba susurronis quasi simplicia et ipsa perveniunt ad intima ventris
PROV|26|23|quomodo si argento sordido ornare velis vas fictile sic labia tumentia cum pessimo corde sociata
PROV|26|24|labiis suis intellegitur inimicus cum in corde tractaverit dolos
PROV|26|25|quando submiserit vocem suam ne credideris ei quoniam septem nequitiae sunt in corde illius
PROV|26|26|qui operit odium fraudulenter revelabitur malitia eius in concilio
PROV|26|27|qui fodit foveam incidet in eam et qui volvit lapidem revertetur ad eum
PROV|26|28|lingua fallax non amat veritatem et os lubricum operatur ruinas
PROV|27|1|ne glorieris in crastinum ignorans quid superventura pariat dies
PROV|27|2|laudet te alienus et non os tuum extraneus et non labia tua
PROV|27|3|grave est saxum et onerosa harena sed ira stulti utroque gravior
PROV|27|4|ira non habet misericordiam nec erumpens furor et impetum concitati ferre quis poterit
PROV|27|5|melior est manifesta correptio quam amor absconditus
PROV|27|6|meliora sunt vulnera diligentis quam fraudulenta odientis oscula
PROV|27|7|anima saturata calcabit favum anima esuriens et amarum pro dulce sumet
PROV|27|8|sicut avis transmigrans de nido suo sic vir qui relinquit locum suum
PROV|27|9|unguento et variis odoribus delectatur cor et bonis amici consiliis anima dulcoratur
PROV|27|10|amicum tuum et amicum patris tui ne dimiseris et domum fratris tui ne ingrediaris in die adflictionis tuae melior est vicinus iuxta quam frater procul
PROV|27|11|stude sapientiae fili mi et laetifica cor meum ut possim exprobranti respondere sermonem
PROV|27|12|astutus videns malum absconditus est parvuli transeuntes sustinuere dispendia
PROV|27|13|tolle vestimentum eius qui spopondit pro extraneo et pro alienis auferto pignus
PROV|27|14|qui benedicit proximo suo voce grandi de nocte consurgens maledicenti similis erit
PROV|27|15|tecta perstillantia in die frigoris et litigiosa mulier conparantur
PROV|27|16|qui retinet eam quasi qui ventum teneat et oleum dexterae suae vocabit
PROV|27|17|ferrum ferro acuitur et homo exacuit faciem amici sui
PROV|27|18|qui servat ficum comedet fructus eius et qui custos est domini sui glorificabitur
PROV|27|19|quomodo in aquis resplendent vultus prospicientium sic corda hominum manifesta sunt prudentibus
PROV|27|20|infernus et perditio non replentur similiter et oculi hominum insatiabiles
PROV|27|21|quomodo probatur in conflatorio argentum et in fornace aurum sic probatur homo ore laudantis
PROV|27|22|si contuderis stultum in pila quasi tisanas feriente desuper pilo non auferetur ab eo stultitia eius
PROV|27|23|diligenter agnosce vultum pecoris tui tuosque greges considera
PROV|27|24|non enim habebis iugiter potestatem sed corona tribuetur in generatione generationum
PROV|27|25|aperta sunt prata et apparuerunt herbae virentes et collecta sunt faena de montibus
PROV|27|26|agni ad vestimentum tuum et hedi agri pretium
PROV|27|27|sufficiat tibi lac caprarum in cibos tuos in necessaria domus tuae et ad victum ancillis tuis
PROV|28|1|fugit impius nemine persequente iustus autem quasi leo confidens absque terrore erit
PROV|28|2|propter peccata terrae multi principes eius et propter hominis sapientiam et horum scientiam quae dicuntur vita ducis longior erit
PROV|28|3|vir pauper calumnians pauperes similis imbri vehementi in quo paratur fames
PROV|28|4|qui derelinquunt legem laudant impium qui custodiunt succenduntur contra eum
PROV|28|5|viri mali non cogitant iudicium qui autem requirunt Dominum animadvertunt omnia
PROV|28|6|melior est pauper ambulans in simplicitate sua quam dives pravis itineribus
PROV|28|7|qui custodit legem filius sapiens est qui pascit comesatores confundit patrem suum
PROV|28|8|qui coacervat divitias usuris et fenore liberali in pauperes congregat eas
PROV|28|9|qui declinat aurem suam ne audiat legem oratio eius erit execrabilis
PROV|28|10|qui decipit iustos in via mala in interitu suo corruet et simplices possidebunt bona
PROV|28|11|sapiens sibi videtur vir dives pauper autem prudens scrutabitur eum
PROV|28|12|in exultatione iustorum multa gloria regnantibus impiis ruinae hominum
PROV|28|13|qui abscondit scelera sua non dirigetur qui confessus fuerit et reliquerit ea misericordiam consequetur
PROV|28|14|beatus homo qui semper est pavidus qui vero mentis est durae corruet in malum
PROV|28|15|leo rugiens et ursus esuriens princeps impius super populum pauperem
PROV|28|16|dux indigens prudentia multos opprimet per calumniam qui autem odit avaritiam longi fient dies eius
PROV|28|17|hominem qui calumniatur animae sanguinem si usque ad lacum fugerit nemo sustentet
PROV|28|18|qui ambulat simpliciter salvus erit qui perversis ingreditur viis concidet semel
PROV|28|19|qui operatur terram suam saturabitur panibus qui sectatur otium replebitur egestate
PROV|28|20|vir fidelis multum laudabitur qui autem festinat ditari non erit innocens
PROV|28|21|qui cognoscit in iudicio faciem non facit bene iste et pro buccella panis deserit veritatem
PROV|28|22|vir qui festinat ditari et aliis invidet ignorat quod egestas superveniat ei
PROV|28|23|qui corripit hominem gratiam postea inveniet apud eum magis quam ille qui per linguae blandimenta decipit
PROV|28|24|qui subtrahit aliquid a patre suo et matre et dicit hoc non est peccatum particeps homicidae est
PROV|28|25|qui se iactat et dilatat iurgia concitat qui sperat in Domino saginabitur
PROV|28|26|qui confidit in corde suo stultus est qui autem graditur sapienter iste salvabitur
PROV|28|27|qui dat pauperi non indigebit qui despicit deprecantem sustinebit penuriam
PROV|28|28|cum surrexerint impii abscondentur homines cum illi perierint multiplicabuntur iusti
PROV|29|1|viro qui corripientem dura cervice contemnit repentinus superveniet interitus et eum sanitas non sequitur
PROV|29|2|in multiplicatione iustorum laetabitur vulgus cum impii sumpserint principatum gemet populus
PROV|29|3|vir qui amat sapientiam laetificat patrem suum qui autem nutrit scorta perdet substantiam
PROV|29|4|rex iustus erigit terram vir avarus destruet eam
PROV|29|5|homo qui blandis fictisque sermonibus loquitur amico suo rete expandit gressibus eius
PROV|29|6|peccantem virum iniquum involvet laqueus et iustus laudabit atque gaudebit
PROV|29|7|novit iustus causam pauperum impius ignorat scientiam
PROV|29|8|homines pestilentes dissipant civitatem sapientes avertunt furorem
PROV|29|9|vir sapiens si cum stulto contenderit sive irascatur sive rideat non inveniet requiem
PROV|29|10|viri sanguinum oderunt simplicem iusti quaerunt animam eius
PROV|29|11|totum spiritum suum profert stultus sapiens differt et reservat in posterum
PROV|29|12|princeps qui libenter audit verba mendacii omnes ministros habebit impios
PROV|29|13|pauper et creditor obviam fuerunt sibi utriusque inluminator est Dominus
PROV|29|14|rex qui iudicat in veritate pauperes thronus eius in aeternum firmabitur
PROV|29|15|virga atque correptio tribuet sapientiam puer autem qui dimittitur voluntati suae confundet matrem suam
PROV|29|16|in multiplicatione impiorum multiplicabuntur scelera et iusti ruinas eorum videbunt
PROV|29|17|erudi filium tuum et refrigerabit te et dabit delicias animae tuae
PROV|29|18|cum prophetia defecerit dissipabitur populus qui custodit legem beatus est
PROV|29|19|servus verbis non potest erudiri quia quod dicis intellegit et respondere contemnit
PROV|29|20|vidisti hominem velocem ad loquendum stulti magis speranda est quam illius correptio
PROV|29|21|qui delicate a pueritia nutrit servum suum postea illum sentiet contumacem
PROV|29|22|vir iracundus provocat rixas et qui ad indignandum facilis est erit ad peccata proclivior
PROV|29|23|superbum sequitur humilitas et humilem spiritu suscipiet gloria
PROV|29|24|qui cum fure partitur odit animam suam adiurantem audit et non indicat
PROV|29|25|qui timet hominem cito corruet qui sperat in Domino sublevabitur
PROV|29|26|multi requirunt faciem principis et a Domino iudicium egreditur singulorum
PROV|29|27|abominantur iusti virum impium et abominantur impii eos qui in recta sunt via
PROV|30|1|verba Congregantis filii Vomentis visio quam locutus est vir cum quo est Deus et qui Deo secum morante confortatus ait
PROV|30|2|stultissimus sum virorum et sapientia hominum non est mecum
PROV|30|3|non didici sapientiam et non novi sanctorum scientiam
PROV|30|4|quis ascendit in caelum atque descendit quis continuit spiritum manibus suis quis conligavit aquas quasi in vestimento quis suscitavit omnes terminos terrae quod nomen eius et quod nomen filii eius si nosti
PROV|30|5|omnis sermo Dei ignitus clypeus est sperantibus in se
PROV|30|6|ne addas quicquam verbis illius et arguaris inveniarisque mendax
PROV|30|7|duo rogavi te ne deneges mihi antequam moriar
PROV|30|8|vanitatem et verba mendacia longe fac a me mendicitatem et divitias ne dederis mihi tribue tantum victui meo necessaria
PROV|30|9|ne forte saturatus inliciar ad negandum et dicam quis est Dominus et egestate conpulsus furer et peierem nomen Dei mei
PROV|30|10|ne accuses servum ad dominum suum ne forte maledicat tibi et corruas
PROV|30|11|generatio quae patri suo maledicit et quae non benedicit matri suae
PROV|30|12|generatio quae sibi munda videtur et tamen non est lota a sordibus suis
PROV|30|13|generatio cuius excelsi sunt oculi et palpebrae eius in alta subrectae
PROV|30|14|generatio quae pro dentibus gladios habet et commandit molaribus suis ut comedat inopes de terra et pauperes ex hominibus
PROV|30|15|sanguisugae duae sunt filiae dicentes adfer adfer tria sunt insaturabilia et quartum quod numquam dicit sufficit
PROV|30|16|infernus et os vulvae et terra quae non satiatur aqua ignis vero numquam dicit sufficit
PROV|30|17|oculum qui subsannat patrem et qui despicit partum matris suae effodiant corvi de torrentibus et comedant illum filii aquilae
PROV|30|18|tria sunt difficilia mihi et quartum penitus ignoro
PROV|30|19|viam aquilae in caelo viam colubri super petram viam navis in medio mari et viam viri in adulescentula
PROV|30|20|talis est via mulieris adulterae quae comedit et tergens os suum dicit non sum operata malum
PROV|30|21|per tria movetur terra et quartum non potest sustinere
PROV|30|22|per servum cum regnaverit per stultum cum saturatus fuerit cibo
PROV|30|23|per odiosam mulierem cum in matrimonio fuerit adsumpta et per ancillam cum heres fuerit dominae suae
PROV|30|24|quattuor sunt minima terrae et ipsa sunt sapientiora sapientibus
PROV|30|25|formicae populus infirmus quae praeparant in messe cibum sibi
PROV|30|26|lepusculus plebs invalida quae conlocat in petra cubile suum
PROV|30|27|regem lucusta non habet et egreditur universa per turmas
PROV|30|28|stilio manibus nititur et moratur in aedibus regis
PROV|30|29|tria sunt quae bene gradiuntur et quartum quod incedit feliciter
PROV|30|30|leo fortissimus bestiarum ad nullius pavebit occursum
PROV|30|31|gallus succinctus lumbos et aries nec est rex qui resistat ei
PROV|30|32|et qui stultus apparuit postquam elatus est in sublime si enim intellexisset ori inposuisset manum
PROV|30|33|qui autem fortiter premit ubera ad eliciendum lac exprimit butyrum et qui vehementer emungitur elicit sanguinem et qui provocat iras producit discordias
PROV|31|1|verba Lamuhel regis visio qua erudivit eum mater sua
PROV|31|2|quid dilecte mi quid dilecte uteri mei quid dilecte votorum meorum
PROV|31|3|ne dederis mulieribus substantiam tuam et vias tuas ad delendos reges
PROV|31|4|noli regibus o Lamuhel noli regibus dare vinum quia nullum secretum est ubi regnat ebrietas
PROV|31|5|ne forte bibat et obliviscatur iudiciorum et mutet causam filiorum pauperis
PROV|31|6|date siceram maerentibus et vinum his qui amaro sunt animo
PROV|31|7|bibant ut obliviscantur egestatis suae et doloris non recordentur amplius
PROV|31|8|aperi os tuum muto et causis omnium filiorum qui pertranseunt
PROV|31|9|aperi os tuum decerne quod iustum est et iudica inopem et pauperem
PROV|31|10|aleph mulierem fortem quis inveniet procul et de ultimis finibus pretium eius
PROV|31|11|beth confidit in ea cor viri sui et spoliis non indigebit
PROV|31|12|gimel reddet ei bonum et non malum omnibus diebus vitae suae
PROV|31|13|deleth quaesivit lanam et linum et operata est consilio manuum suarum
PROV|31|14|he facta est quasi navis institoris de longe portat panem suum
PROV|31|15|vav et de nocte surrexit deditque praedam domesticis suis et cibaria ancillis suis
PROV|31|16|zai consideravit agrum et emit eum de fructu manuum suarum plantavit vineam
PROV|31|17|heth accinxit fortitudine lumbos suos et roboravit brachium suum
PROV|31|18|teth gustavit quia bona est negotiatio eius non extinguetur in nocte lucerna illius
PROV|31|19|ioth manum suam misit ad fortia et digiti eius adprehenderunt fusum
PROV|31|20|caph manum suam aperuit inopi et palmas suas extendit ad pauperem
PROV|31|21|lameth non timebit domui suae a frigoribus nivis omnes enim domestici eius vestiti duplicibus
PROV|31|22|mem stragulam vestem fecit sibi byssus et purpura indumentum eius
PROV|31|23|nun nobilis in portis vir eius quando sederit cum senatoribus terrae
PROV|31|24|samech sindonem fecit et vendidit et cingulum tradidit Chananeo
PROV|31|25|ain fortitudo et decor indumentum eius et ridebit in die novissimo
PROV|31|26|phe os suum aperuit sapientiae et lex clementiae in lingua eius
PROV|31|27|sade considerat semitas domus suae et panem otiosa non comedet
PROV|31|28|coph surrexerunt filii eius et beatissimam praedicaverunt vir eius et laudavit eam
PROV|31|29|res multae filiae congregaverunt divitias tu supergressa es universas
PROV|31|30|sin fallax gratia et vana est pulchritudo mulier timens Dominum ipsa laudabitur
PROV|31|31|thau date ei de fructu manuum suarum et laudent eam in portis opera eius
