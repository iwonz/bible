ISA|1|1|The vision of Isaiah the son of Amoz, which he saw concerning Judah and Jerusalem in the days of Uzziah, Jotham, Ahaz, and Hezekiah, kings of Judah.
ISA|1|2|Hear, O heavens, and give ear, O earth; for the LORD has spoken: "Children have I reared and brought up, but they have rebelled against me.
ISA|1|3|The ox knows its owner, and the donkey its master's crib, but Israel does not know, my people do not understand."
ISA|1|4|Ah, sinful nation, a people laden with iniquity, offspring of evildoers, children who deal corruptly! They have forsaken the LORD, they have despised the Holy One of Israel, they are utterly estranged.
ISA|1|5|Why will you still be struck down? Why will you continue to rebel? The whole head is sick, and the whole heart faint.
ISA|1|6|From the sole of the foot even to the head, there is no soundness in it, but bruises and sores and raw wounds; they are not pressed out or bound up or softened with oil.
ISA|1|7|Your country lies desolate; your cities are burned with fire; in your very presence foreigners devour your land; it is desolate, as overthrown by foreigners.
ISA|1|8|And the daughter of Zion is left like a booth in a vineyard, like a lodge in a cucumber field, like a besieged city.
ISA|1|9|If the LORD of hosts had not left us a few survivors, we should have been like Sodom, and become like Gomorrah.
ISA|1|10|Hear the word of the LORD, you rulers of Sodom! Give ear to the teaching of our God, you people of Gomorrah!
ISA|1|11|"What to me is the multitude of your sacrifices? says the LORD; I have had enough of burnt offerings of rams and the fat of well-fed beasts; I do not delight in the blood of bulls, or of lambs, or of goats.
ISA|1|12|"When you come to appear before me, who has required of you this trampling of my courts?
ISA|1|13|Bring no more vain offerings; incense is an abomination to me. New moon and Sabbath and the calling of convocations- I cannot endure iniquity and solemn assembly.
ISA|1|14|Your new moons and your appointed feasts my soul hates; they have become a burden to me; I am weary of bearing them.
ISA|1|15|When you spread out your hands, I will hide my eyes from you; even though you make many prayers, I will not listen; your hands are full of blood.
ISA|1|16|Wash yourselves; make yourselves clean; remove the evil of your deeds from before my eyes; cease to do evil,
ISA|1|17|learn to do good; seek justice, correct oppression; bring justice to the fatherless, plead the widow's cause.
ISA|1|18|"Come now, let us reason together, says the LORD: though your sins are like scarlet, they shall be as white as snow; though they are red like crimson, they shall become like wool.
ISA|1|19|If you are willing and obedient, you shall eat the good of the land;
ISA|1|20|but if you refuse and rebel, you shall be eaten by the sword; for the mouth of the LORD has spoken."
ISA|1|21|How the faithful city has become a whore, she who was full of justice! Righteousness lodged in her, but now murderers.
ISA|1|22|Your silver has become dross, your best wine mixed with water.
ISA|1|23|Your princes are rebels and companions of thieves. Everyone loves a bribe and runs after gifts. They do not bring justice to the fatherless, and the widow's cause does not come to them.
ISA|1|24|Therefore the Lord declares, the LORD of hosts, the Mighty One of Israel: "Ah, I will get relief from my enemies and avenge myself on my foes.
ISA|1|25|I will turn my hand against you and will smelt away your dross as with lye and remove all your alloy.
ISA|1|26|And I will restore your judges as at the first, and your counselors as at the beginning. Afterward you shall be called the city of righteousness, the faithful city."
ISA|1|27|Zion shall be redeemed by justice, and those in her who repent, by righteousness.
ISA|1|28|But rebels and sinners shall be broken together, and those who forsake the LORD shall be consumed.
ISA|1|29|For they shall be ashamed of the oaks that you desired; and you shall blush for the gardens that you have chosen.
ISA|1|30|For you shall be like an oak whose leaf withers, and like a garden without water.
ISA|1|31|And the strong shall become tinder, and his work a spark, and both of them shall burn together, with none to quench them.
ISA|2|1|The word that Isaiah the son of Amoz saw concerning Judah and Jerusalem.
ISA|2|2|It shall come to pass in the latter days that the mountain of the house of the LORD shall be established as the highest of the mountains, and shall be lifted up above the hills; and all the nations shall flow to it,
ISA|2|3|and many peoples shall come, and say: "Come, let us go up to the mountain of the LORD, to the house of the God of Jacob, that he may teach us his ways and that we may walk in his paths." For out of Zion shall go the law, and the word of the LORD from Jerusalem.
ISA|2|4|He shall judge between the nations, and shall decide disputes for many peoples; and they shall beat their swords into plowshares, and their spears into pruning hooks; nation shall not lift up sword against nation, neither shall they learn war anymore.
ISA|2|5|O house of Jacob, come, let us walk in the light of the LORD.
ISA|2|6|For you have rejected your people, the house of Jacob, because they are full of things from the east and of fortunetellers like the Philistines, and they strike hands with the children of foreigners.
ISA|2|7|Their land is filled with silver and gold, and there is no end to their treasures; their land is filled with horses, and there is no end to their chariots.
ISA|2|8|Their land is filled with idols; they bow down to the work of their hands, to what their own fingers have made.
ISA|2|9|So man is humbled, and each one is brought low- do not forgive them!
ISA|2|10|Enter into the rock and hide in the dust from before the terror of the LORD, and from the splendor of his majesty.
ISA|2|11|The haughty looks of man shall be brought low, and the lofty pride of men shall be humbled, and the LORD alone will be exalted in that day.
ISA|2|12|For the LORD of hosts has a day against all that is proud and lofty, against all that is lifted up- and it shall be brought low;
ISA|2|13|against all the cedars of Lebanon, lofty and lifted up; and against all the oaks of Bashan;
ISA|2|14|against all the lofty mountains, and against all the uplifted hills;
ISA|2|15|against every high tower, and against every fortified wall;
ISA|2|16|against all the ships of Tarshish, and against all the beautiful craft.
ISA|2|17|And the haughtiness of man shall be humbled, and the lofty pride of men shall be brought low, and the LORD alone will be exalted in that day.
ISA|2|18|And the idols shall utterly pass away.
ISA|2|19|And people shall enter the caves of the rocks and the holes of the ground, from before the terror of the LORD, and from the splendor of his majesty, when he rises to terrify the earth.
ISA|2|20|In that day mankind will cast away their idols of silver and their idols of gold, which they made for themselves to worship, to the moles and to the bats,
ISA|2|21|to enter the caverns of the rocks and the clefts of the cliffs, from before the terror of the LORD, and from the splendor of his majesty, when he rises to terrify the earth.
ISA|2|22|Stop regarding man in whose nostrils is breath, for of what account is he?
ISA|3|1|For behold, the Lord GOD of hosts is taking away from Jerusalem and from Judah support and supply, all support of bread, and all support of water;
ISA|3|2|the mighty man and the soldier, the judge and the prophet, the diviner and the elder,
ISA|3|3|the captain of fifty and the man of rank, the counselor and the skillful magician and the expert in charms.
ISA|3|4|And I will make boys their princes, and infants shall rule over them.
ISA|3|5|And the people will oppress one another, every one his fellow and every one his neighbor; the youth will be insolent to the elder, and the despised to the honorable.
ISA|3|6|For a man will take hold of his brother in the house of his father, saying: "You have a cloak; you shall be our leader, and this heap of ruins shall be under your rule";
ISA|3|7|in that day he will speak out, saying: "I will not be a healer; in my house there is neither bread nor cloak; you shall not make me leader of the people."
ISA|3|8|For Jerusalem has stumbled, and Judah has fallen, because their speech and their deeds are against the LORD, defying his glorious presence.
ISA|3|9|For the look on their faces bears witness against them; they proclaim their sin like Sodom; they do not hide it. Woe to them! For they have brought evil on themselves.
ISA|3|10|Tell the righteous that it shall be well with them, for they shall eat the fruit of their deeds.
ISA|3|11|Woe to the wicked! It shall be ill with him, for what his hands have dealt out shall be done to him.
ISA|3|12|My people- infants are their oppressors, and women rule over them. O my people, your guides mislead you and they have swallowed up the course of your paths.
ISA|3|13|The LORD has taken his place to contend; he stands to judge peoples.
ISA|3|14|The LORD will enter into judgment with the elders and princes of his people: "It is you who have devoured the vineyard, the spoil of the poor is in your houses.
ISA|3|15|What do you mean by crushing my people, by grinding the face of the poor?" declares the Lord GOD of hosts.
ISA|3|16|The LORD said: Because the daughters of Zion are haughty and walk with outstretched necks, glancing wantonly with their eyes, mincing along as they go, tinkling with their feet,
ISA|3|17|therefore the Lord will strike with a scab the heads of the daughters of Zion, and the LORD will lay bare their secret parts.
ISA|3|18|In that day the Lord will take away the finery of the anklets, the headbands, and the crescents;
ISA|3|19|the pendants, the bracelets, and the scarves;
ISA|3|20|the headdresses, the armlets, the sashes, the perfume boxes, and the amulets;
ISA|3|21|the signet rings and nose rings;
ISA|3|22|the festal robes, the mantles, the cloaks, and the handbags;
ISA|3|23|the mirrors, the linen garments, the turbans, and the veils.
ISA|3|24|Instead of perfume there will be rottenness; and instead of a belt, a rope; and instead of well-set hair, baldness; and instead of a rich robe, a skirt of sackcloth; and branding instead of beauty.
ISA|3|25|Your men shall fall by the sword and your mighty men in battle.
ISA|3|26|And her gates shall lament and mourn; empty, she shall sit on the ground.
ISA|4|1|And seven women shall take hold of one man in that day, saying, "We will eat our own bread and wear our own clothes, only let us be called by your name; take away our reproach."
ISA|4|2|In that day the branch of the LORD shall be beautiful and glorious, and the fruit of the land shall be the pride and honor of the survivors of Israel.
ISA|4|3|And he who is left in Zion and remains in Jerusalem will be called holy, everyone who has been recorded for life in Jerusalem,
ISA|4|4|when the Lord shall have washed away the filth of the daughters of Zion and cleansed the bloodstains of Jerusalem from its midst by a spirit of judgment and by a spirit of burning.
ISA|4|5|Then the LORD will create over the whole site of Mount Zion and over her assemblies a cloud by day, and smoke and the shining of a flaming fire by night; for over all the glory there will be a canopy.
ISA|4|6|There will be a booth for shade by day from the heat, and for a refuge and a shelter from the storm and rain.
ISA|5|1|Let me sing for my beloved my love song concerning his vineyard: My beloved had a vineyard on a very fertile hill.
ISA|5|2|He dug it and cleared it of stones, and planted it with choice vines; he built a watchtower in the midst of it, and hewed out a wine vat in it; and he looked for it to yield grapes, but it yielded wild grapes.
ISA|5|3|And now, O inhabitants of Jerusalem and men of Judah, judge between me and my vineyard.
ISA|5|4|What more was there to do for my vineyard, that I have not done in it? When I looked for it to yield grapes, why did it yield wild grapes?
ISA|5|5|And now I will tell you what I will do to my vineyard. I will remove its hedge, and it shall be devoured; I will break down its wall, and it shall be trampled down.
ISA|5|6|I will make it a waste; it shall not be pruned or hoed, and briers and thorns shall grow up; I will also command the clouds that they rain no rain upon it.
ISA|5|7|For the vineyard of the LORD of hosts is the house of Israel, and the men of Judah are his pleasant planting; and he looked for justice, but behold, bloodshed; for righteousness, but behold, an outcry!
ISA|5|8|Woe to those who join house to house, who add field to field, until there is no more room, and you are made to dwell alone in the midst of the land.
ISA|5|9|The LORD of hosts has sworn in my hearing: "Surely many houses shall be desolate, large and beautiful houses, without inhabitant.
ISA|5|10|For ten acres of vineyard shall yield but one bath, and a homer of seed shall yield but an ephah."
ISA|5|11|Woe to those who rise early in the morning, that they may run after strong drink, who tarry late into the evening as wine inflames them!
ISA|5|12|They have lyre and harp, tambourine and flute and wine at their feasts, but they do not regard the deeds of the LORD, or see the work of his hands.
ISA|5|13|Therefore my people go into exile for lack of knowledge; their honored men go hungry, and their multitude is parched with thirst.
ISA|5|14|Therefore Sheol has enlarged its appetite and opened its mouth beyond measure, and the nobility of Jerusalem and her multitude will go down, her revelers and he who exults in her.
ISA|5|15|Man is humbled, and each one is brought low, and the eyes of the haughty are brought low.
ISA|5|16|But the LORD of hosts is exalted in justice, and the Holy God shows himself holy in righteousness.
ISA|5|17|Then shall the lambs graze as in their pasture, and nomads shall eat among the ruins of the rich.
ISA|5|18|Woe to those who draw iniquity with cords of falsehood, who draw sin as with cart ropes,
ISA|5|19|who say: "Let him be quick, let him speed his work that we may see it; let the counsel of the Holy One of Israel draw near, and let it come, that we may know it!"
ISA|5|20|Woe to those who call evil good and good evil, who put darkness for light and light for darkness, who put bitter for sweet and sweet for bitter!
ISA|5|21|Woe to those who are wise in their own eyes, and shrewd in their own sight!
ISA|5|22|Woe to those who are heroes at drinking wine, and valiant men in mixing strong drink,
ISA|5|23|who acquit the guilty for a bribe, and deprive the innocent of his right!
ISA|5|24|Therefore, as the tongue of fire devours the stubble, and as dry grass sinks down in the flame, so their root will be as rottenness, and their blossom go up like dust; for they have rejected the law of the LORD of hosts, and have despised the word of the Holy One of Israel.
ISA|5|25|Therefore the anger of the LORD was kindled against his people, and he stretched out his hand against them and struck them, and the mountains quaked; and their corpses were as refuse in the midst of the streets. For all this his anger has not turned away, and his hand is stretched out still.
ISA|5|26|He will raise a signal for nations afar off, and whistle for them from the ends of the earth; and behold, quickly, speedily they come!
ISA|5|27|None is weary, none stumbles, none slumbers or sleeps, not a waistband is loose, not a sandal strap broken;
ISA|5|28|their arrows are sharp, all their bows bent, their horses' hoofs seem like flint, and their wheels like the whirlwind.
ISA|5|29|Their roaring is like a lion, like young lions they roar; they growl and seize their prey; they carry it off, and none can rescue.
ISA|5|30|They will growl over it on that day, like the growling of the sea. And if one looks to the land, behold, darkness and distress; and the light is darkened by its clouds.
ISA|6|1|In the year that King Uzziah died I saw the Lord sitting upon a throne, high and lifted up; and the train of his robe filled the temple.
ISA|6|2|Above him stood the seraphim. Each had six wings: with two he covered his face, and with two he covered his feet, and with two he flew.
ISA|6|3|And one called to another and said: "Holy, holy, holy is the LORD of hosts; the whole earth is full of his glory!"
ISA|6|4|And the foundations of the thresholds shook at the voice of him who called, and the house was filled with smoke.
ISA|6|5|And I said: "Woe is me! For I am lost; for I am a man of unclean lips, and I dwell in the midst of a people of unclean lips; for my eyes have seen the King, the LORD of hosts!"
ISA|6|6|Then one of the seraphim flew to me, having in his hand a burning coal that he had taken with tongs from the altar.
ISA|6|7|And he touched my mouth and said: "Behold, this has touched your lips; your guilt is taken away, and your sin atoned for.
ISA|6|8|And I heard the voice of the Lord saying, "Whom shall I send, and who will go for us?" Then I said, "Here am I! Send me."
ISA|6|9|And he said, "Go, and say to this people: "' Keep on hearing, but do not understand; keep on seeing, but do not perceive.'
ISA|6|10|Make the heart of this people dull, and their ears heavy, and blind their eyes; lest they see with their eyes, and hear with their ears, and understand with their hearts, and turn and be healed."
ISA|6|11|Then I said, "How long, O Lord?" And he said: "Until cities lie waste without inhabitant, and houses without people, and the land is a desolate waste,
ISA|6|12|and the LORD removes people far away, and the forsaken places are many in the midst of the land.
ISA|6|13|And though a tenth remain in it, it will be burned again, like a terebinth or an oak, whose stump remains when it is felled." The holy seed is its stump.
ISA|7|1|In the days of Ahaz the son of Jotham, son of Uzziah, king of Judah, Rezin the king of Syria and Pekah the son of Remaliah the king of Israel came up to Jerusalem to wage war against it, but could not yet mount an attack against it.
ISA|7|2|When the house of David was told, "Syria is in league with Ephraim," the heart of Ahaz and the heart of his people shook as the trees of the forest shake before the wind.
ISA|7|3|And the LORD said to Isaiah, "Go out to meet Ahaz, you and Shear-jashub your son, at the end of the conduit of the upper pool on the highway to the Washer's Field.
ISA|7|4|And say to him, 'Be careful, be quiet, do not fear, and do not let your heart be faint because of these two smoldering stumps of firebrands, at the fierce anger of Rezin and Syria and the son of Remaliah.
ISA|7|5|Because Syria, with Ephraim and the son of Remaliah, has devised evil against you, saying,
ISA|7|6|"Let us go up against Judah and terrify it, and let us conquer it for ourselves, and set up the son of Tabeel as king in the midst of it,"
ISA|7|7|thus says the Lord GOD: "' It shall not stand, and it shall not come to pass.
ISA|7|8|For the head of Syria is Damascus, and the head of Damascus is Rezin. (Within sixty-five years Ephraim will be broken to pieces so that it will no longer be a people.)
ISA|7|9|"'And the head of Ephraim is Samaria, and the head of Samaria is the son of Remaliah. If you are not firm in faith, you will not be firm at all.'"
ISA|7|10|Again the LORD spoke to Ahaz,
ISA|7|11|"Ask a sign of the LORD your God; let it be deep as Sheol or high as heaven."
ISA|7|12|But Ahaz said, "I will not ask, and I will not put the LORD to the test."
ISA|7|13|And he said, "Hear then, O house of David! Is it too little for you to weary men, that you weary my God also?
ISA|7|14|Therefore the Lord himself will give you a sign. Behold, the virgin shall conceive and bear a son, and shall call his name Immanuel.
ISA|7|15|He shall eat curds and honey when he knows how to refuse the evil and choose the good.
ISA|7|16|For before the boy knows how to refuse the evil and choose the good, the land whose two kings you dread will be deserted.
ISA|7|17|The LORD will bring upon you and upon your people and upon your father's house such days as have not come since the day that Ephraim departed from Judah- the king of Assyria."
ISA|7|18|In that day the LORD will whistle for the fly that is at the end of the streams of Egypt, and for the bee that is in the land of Assyria.
ISA|7|19|And they will all come and settle in the steep ravines, and in the clefts of the rocks, and on all the thornbushes, and on all the pastures.
ISA|7|20|In that day the Lord will shave with a razor that is hired beyond the River- with the king of Assyria- the head and the hair of the feet, and it will sweep away the beard also.
ISA|7|21|In that day a man will keep alive a young cow and two sheep,
ISA|7|22|and because of the abundance of milk that they give, he will eat curds, for everyone who is left in the land will eat curds and honey.
ISA|7|23|In that day every place where there used to be a thousand vines, worth a thousand shekels of silver, will become briers and thorns.
ISA|7|24|With bow and arrows a man will come there, for all the land will be briers and thorns.
ISA|7|25|And as for all the hills that used to be hoed with a hoe, you will not come there for fear of briers and thorns, but they will become a place where cattle are let loose and where sheep tread.
ISA|8|1|Then the LORD said to me, "Take a large tablet and write on it in common characters, 'Belonging to Maher-shalal-hashbaz.'
ISA|8|2|And I will get reliable witnesses, Uriah the priest and Zechariah the son of Jeberechiah, to attest for me."
ISA|8|3|And I went to the prophetess, and she conceived and bore a son. Then the LORD said to me, "Call his name Maher-shalal-hashbaz;
ISA|8|4|for before the boy knows how to cry 'My father' or 'My mother,' the wealth of Damascus and the spoil of Samaria will be carried away before the king of Assyria."
ISA|8|5|The LORD spoke to me again:
ISA|8|6|"Because this people have refused the waters of Shiloah that flow gently, and rejoice over Rezin and the son of Remaliah,
ISA|8|7|therefore, behold, the Lord is bringing up against them the waters of the River, mighty and many, the king of Assyria and all his glory. And it will rise over all its channels and go over all its banks,
ISA|8|8|and it will sweep on into Judah, it will overflow and pass on, reaching even to the neck, and its outspread wings will fill the breadth of your land, O Immanuel."
ISA|8|9|Be broken, you peoples, and be shattered; give ear, all you far countries; strap on your armor and be shattered; strap on your armor and be shattered.
ISA|8|10|Take counsel together, but it will come to nothing; speak a word, but it will not stand, for God is with us.
ISA|8|11|For the LORD spoke thus to me with his strong hand upon me, and warned me not to walk in the way of this people, saying:
ISA|8|12|"Do not call conspiracy all that this people calls conspiracy, and do not fear what they fear, nor be in dread.
ISA|8|13|But the LORD of hosts, him you shall regard as holy. Let him be your fear, and let him be your dread.
ISA|8|14|And he will become a sanctuary and a stone of offense and a rock of stumbling to both houses of Israel, a trap and a snare to the inhabitants of Jerusalem.
ISA|8|15|And many shall stumble on it. They shall fall and be broken; they shall be snared and taken."
ISA|8|16|Bind up the testimony; seal the teaching among my disciples.
ISA|8|17|I will wait for the LORD, who is hiding his face from the house of Jacob, and I will hope in him.
ISA|8|18|Behold, I and the children whom the LORD has given me are signs and portents in Israel from the LORD of hosts, who dwells on Mount Zion.
ISA|8|19|And when they say to you, "Inquire of the mediums and the necromancers who chirp and mutter," should not a people inquire of their God? Should they inquire of the dead on behalf of the living?
ISA|8|20|To the teaching and to the testimony! If they will not speak according to this word, it is because they have no dawn.
ISA|8|21|They will pass through the land, greatly distressed and hungry. And when they are hungry, they will be enraged and will speak contemptuously against their king and their God, and turn their faces upward.
ISA|8|22|And they will look to the earth, but behold, distress and darkness, the gloom of anguish. And they will be thrust into thick darkness.
ISA|9|1|But there will be no gloom for her who was in anguish. In the former time he brought into contempt the land of Zebulun and the land of Naphtali, but in the latter time he has made glorious the way of the sea, the land beyond the Jordan, Galilee of the nations.
ISA|9|2|The people who walked in darkness have seen a great light; those who dwelt in a land of deep darkness, on them has light shined.
ISA|9|3|You have multiplied the nation; you have increased its joy; they rejoice before you as with joy at the harvest, as they are glad when they divide the spoil.
ISA|9|4|For the yoke of his burden, and the staff for his shoulder, the rod of his oppressor, you have broken as on the day of Midian.
ISA|9|5|For every boot of the tramping warrior in battle tumult and every garment rolled in blood will be burned as fuel for the fire.
ISA|9|6|For to us a child is born, to us a son is given; and the government shall be upon his shoulder, and his name shall be called Wonderful Counselor, Mighty God, Everlasting Father, Prince of Peace.
ISA|9|7|Of the increase of his government and of peace there will be no end, on the throne of David and over his kingdom, to establish it and to uphold it with justice and with righteousness from this time forth and forevermore. The zeal of the LORD of hosts will do this.
ISA|9|8|The Lord has sent a word against Jacob, and it will fall on Israel;
ISA|9|9|and all the people will know, Ephraim and the inhabitants of Samaria, who say in pride and in arrogance of heart:
ISA|9|10|"The bricks have fallen, but we will build with dressed stones; the sycamores have been cut down, but we will put cedars in their place."
ISA|9|11|But the LORD raises the adversaries of Rezin against him, and stirs up his enemies.
ISA|9|12|The Syrians on the east and the Philistines on the west devour Israel with open mouth. For all this his anger has not turned away, and his hand is stretched out still.
ISA|9|13|The people did not turn to him who struck them, nor inquire of the LORD of hosts.
ISA|9|14|So the LORD cut off from Israel head and tail, palm branch and reed in one day-
ISA|9|15|the elder and honored man is the head, and the prophet who teaches lies is the tail;
ISA|9|16|for those who guide this people have been leading them astray, and those who are guided by them are swallowed up.
ISA|9|17|Therefore the Lord does not rejoice over their young men, and has no compassion on their fatherless and widows; for everyone is godless and an evildoer, and every mouth speaks folly. For all this his anger has not turned away, and his hand is stretched out still.
ISA|9|18|For wickedness burns like a fire; it consumes briers and thorns; it kindles the thickets of the forest, and they roll upward in a column of smoke.
ISA|9|19|Through the wrath of the LORD of hosts the land is scorched, and the people are like fuel for the fire; no one spares another.
ISA|9|20|They slice meat on the right, but are still hungry, and they devour on the left, but are not satisfied; each devours the flesh of his own arm,
ISA|9|21|Manasseh devours Ephraim, and Ephraim devours Manasseh; together they are against Judah. For all this his anger has not turned away, and his hand is stretched out still.
ISA|10|1|Woe to those who decree iniquitous decrees, and the writers who keep writing oppression,
ISA|10|2|to turn aside the needy from justice and to rob the poor of my people of their right, that widows may be their spoil, and that they may make the fatherless their prey!
ISA|10|3|What will you do on the day of punishment, in the ruin that will come from afar? To whom will you flee for help, and where will you leave your wealth?
ISA|10|4|Nothing remains but to crouch among the prisoners or fall among the slain. For all this his anger has not turned away, and his hand is stretched out still.
ISA|10|5|Ah, Assyria, the rod of my anger; the staff in their hands is my fury!
ISA|10|6|Against a godless nation I send him, and against the people of my wrath I command him, to take spoil and seize plunder, and to tread them down like the mire of the streets.
ISA|10|7|But he does not so intend, and his heart does not so think; but it is in his heart to destroy, and to cut off nations not a few;
ISA|10|8|for he says: "Are not my commanders all kings?
ISA|10|9|Is not Calno like Carchemish? Is not Hamath like Arpad? Is not Samaria like Damascus?
ISA|10|10|As my hand has reached to the kingdoms of the idols, whose carved images were greater than those of Jerusalem and Samaria,
ISA|10|11|shall I not do to Jerusalem and her idols as I have done to Samaria and her images?"
ISA|10|12|When the Lord has finished all his work on Mount Zion and on Jerusalem, he will punish the speech of the arrogant heart of the king of Assyria and the boastful look in his eyes.
ISA|10|13|For he says: "By the strength of my hand I have done it, and by my wisdom, for I have understanding; I remove the boundaries of peoples, and plunder their treasures; like a bull I bring down those who sit on thrones.
ISA|10|14|My hand has found like a nest the wealth of the peoples; and as one gathers eggs that have been forsaken, so I have gathered all the earth; and there was none that moved a wing or opened the mouth or chirped."
ISA|10|15|Shall the axe boast over him who hews with it, or the saw magnify itself against him who wields it? As if a rod should wield him who lifts it, or as if a staff should lift him who is not wood!
ISA|10|16|Therefore the Lord GOD of hosts will send wasting sickness among his stout warriors, and under his glory a burning will be kindled, like the burning of fire.
ISA|10|17|The light of Israel will become a fire, and his Holy One a flame, and it will burn and devour his thorns and briers in one day.
ISA|10|18|The glory of his forest and of his fruitful land the LORD will destroy, both soul and body, and it will be as when a sick man wastes away.
ISA|10|19|The remnant of the trees of his forest will be so few that a child can write them down.
ISA|10|20|In that day the remnant of Israel and the survivors of the house of Jacob will no more lean on him who struck them, but will lean on the LORD, the Holy One of Israel, in truth.
ISA|10|21|A remnant will return, the remnant of Jacob, to the mighty God.
ISA|10|22|For though your people Israel be as the sand of the sea, only a remnant of them will return. Destruction is decreed, overflowing with righteousness.
ISA|10|23|For the Lord GOD of hosts will make a full end, as decreed, in the midst of all the earth.
ISA|10|24|Therefore thus says the Lord GOD of hosts: "O my people, who dwell in Zion, be not afraid of the Assyrians when they strike with the rod and lift up their staff against you as the Egyptians did.
ISA|10|25|For in a very little while my fury will come to an end, and my anger will be directed to their destruction.
ISA|10|26|And the LORD of hosts will wield against them a whip, as when he struck Midian at the rock of Oreb. And his staff will be over the sea, and he will lift it as he did in Egypt.
ISA|10|27|And in that day his burden will depart from your shoulder, and his yoke from your neck; and the yoke will be broken because of the fat."
ISA|10|28|He has come to Aiath; he has passed through Migron; at Michmash he stores his baggage;
ISA|10|29|they have crossed over the pass; at Geba they lodge for the night; Ramah trembles; Gibeah of Saul has fled.
ISA|10|30|Cry aloud, O daughter of Gallim! Give attention, O Laishah! O Poor Anathoth!
ISA|10|31|Madmenah is in flight; the inhabitants of Gebim flee for safety.
ISA|10|32|This very day he will halt at Nob; he will shake his fist at the mount of the daughter of Zion, the hill of Jerusalem.
ISA|10|33|Behold, the Lord GOD of hosts will lop the boughs with terrifying power; the great in height will be hewn down, and the lofty will be brought low.
ISA|10|34|He will cut down the thickets of the forest with an axe, and Lebanon will fall by the Majestic One.
ISA|11|1|There shall come forth a shoot from the stump of Jesse, and a branch from his roots shall bear fruit.
ISA|11|2|And the Spirit of the LORD shall rest upon him, the Spirit of wisdom and understanding, the Spirit of counsel and might, the Spirit of knowledge and the fear of the LORD.
ISA|11|3|And his delight shall be in the fear of the LORD. He shall not judge by what his eyes see, or decide disputes by what his ears hear,
ISA|11|4|but with righteousness he shall judge the poor, and decide with equity for the meek of the earth; and he shall strike the earth with the rod of his mouth, and with the breath of his lips he shall kill the wicked.
ISA|11|5|Righteousness shall be the belt of his waist, and faithfulness the belt of his loins.
ISA|11|6|The wolf shall dwell with the lamb, and the leopard shall lie down with the young goat, and the calf and the lion and the fattened calf together; and a little child shall lead them.
ISA|11|7|The cow and the bear shall graze; their young shall lie down together; and the lion shall eat straw like the ox.
ISA|11|8|The nursing child shall play over the hole of the cobra, and the weaned child shall put his hand on the adder's den.
ISA|11|9|They shall not hurt or destroy in all my holy mountain; for the earth shall be full of the knowledge of the LORD as the waters cover the sea.
ISA|11|10|In that day the root of Jesse, who shall stand as a signal for the peoples- of him shall the nations inquire, and his resting place shall be glorious.
ISA|11|11|In that day the Lord will extend his hand yet a second time to recover the remnant that remains of his people, from Assyria, from Egypt, from Pathros, from Cush, from Elam, from Shinar, from Hamath, and from the coastlands of the sea.
ISA|11|12|He will raise a signal for the nations and will assemble the banished of Israel, and gather the dispersed of Judah from the four corners of the earth.
ISA|11|13|The jealousy of Ephraim shall depart, and those who harass Judah shall be cut off; Ephraim shall not be jealous of Judah, and Judah shall not harass Ephraim.
ISA|11|14|But they shall swoop down on the shoulder of the Philistines in the west, and together they shall plunder the people of the east. They shall put out their hand against Edom and Moab, and the Ammonites shall obey them.
ISA|11|15|And the LORD will utterly destroy the tongue of the Sea of Egypt, and will wave his hand over the River with his scorching breath, and strike it into seven channels, and he will lead people across in sandals.
ISA|11|16|And there will be a highway from Assyria for the remnant that remains of his people, as there was for Israel when they came up from the land of Egypt.
ISA|12|1|You will say in that day:"I will give thanks to you, O LORD, for though you were angry with me, your anger turned away, that you might comfort me.
ISA|12|2|"Behold, God is my salvation; I will trust, and will not be afraid; for the LORD GOD is my strength and my song, and he has become my salvation."
ISA|12|3|With joy you will draw water from the wells of salvation.
ISA|12|4|And you will say in that day: "Give thanks to the LORD, call upon his name, make known his deeds among the peoples, proclaim that his name is exalted.
ISA|12|5|"Sing praises to the LORD, for he has done gloriously; let this be made known in all the earth.
ISA|12|6|Shout, and sing for joy, O inhabitant of Zion, for great in your midst is the Holy One of Israel."
ISA|13|1|The oracle concerning Babylon which Isaiah the son of Amoz saw.
ISA|13|2|On a bare hill raise a signal; cry aloud to them; wave the hand for them to enter the gates of the nobles.
ISA|13|3|I myself have commanded my consecrated ones, and have summoned my mighty men to execute my anger, my proudly exulting ones.
ISA|13|4|The sound of a tumult is on the mountains as of a great multitude! The sound of an uproar of kingdoms, of nations gathering together! The LORD of hosts is mustering a host for battle.
ISA|13|5|They come from a distant land, from the end of the heavens, the LORD and the weapons of his indignation, to destroy the whole land.
ISA|13|6|Wail, for the day of the LORD is near; as destruction from the Almighty it will come!
ISA|13|7|Therefore all hands will be feeble, and every human heart will melt.
ISA|13|8|They will be dismayed: pangs and agony will seize them; they will be in anguish like a woman in labor. They will look aghast at one another; their faces will be aflame.
ISA|13|9|Behold, the day of the LORD comes, cruel, with wrath and fierce anger, to make the land a desolation and to destroy its sinners from it.
ISA|13|10|For the stars of the heavens and their constellations will not give their light; the sun will be dark at its rising, and the moon will not shed its light.
ISA|13|11|I will punish the world for its evil, and the wicked for their iniquity; I will put an end to the pomp of the arrogant, and lay low the pompous pride of the ruthless.
ISA|13|12|I will make people more rare than fine gold, and mankind than the gold of Ophir.
ISA|13|13|Therefore I will make the heavens tremble, and the earth will be shaken out of its place, at the wrath of the LORD of hosts in the day of his fierce anger.
ISA|13|14|And like a hunted gazelle, or like sheep with none to gather them, each will turn to his own people, and each will flee to his own land.
ISA|13|15|Whoever is found will be thrust through, and whoever is caught will fall by the sword.
ISA|13|16|Their infants will be dashed in pieces before their eyes; their houses will be plundered and their wives ravished.
ISA|13|17|Behold, I am stirring up the Medes against them, who have no regard for silver and do not delight in gold.
ISA|13|18|Their bows will slaughter the young men; they will have no mercy on the fruit of the womb; their eyes will not pity children.
ISA|13|19|And Babylon, the glory of kingdoms, the splendor and pomp of the Chaldeans, will be like Sodom and Gomorrah when God overthrew them.
ISA|13|20|It will never be inhabited or lived in for all generations; no Arab will pitch his tent there; no shepherds will make their flocks lie down there.
ISA|13|21|But wild animals will lie down there, and their houses will be full of howling creatures; there ostriches will dwell, and there wild goats will dance.
ISA|13|22|Hyenas will cry in its towers, and jackals in the pleasant palaces; its time is close at hand and its days will not be prolonged.
ISA|14|1|For the LORD will have compassion on Jacob and will again choose Israel, and will set them in their own land, and sojourners will join them and will attach themselves to the house of Jacob.
ISA|14|2|And the peoples will take them and bring them to their place, and the house of Israel will possess them in the LORD's land as male and female slaves. They will take captive those who were their captors, and rule over those who oppressed them.
ISA|14|3|When the LORD has given you rest from your pain and turmoil and the hard service with which you were made to serve,
ISA|14|4|you will take up this taunt against the king of Babylon: "How the oppressor has ceased, the insolent fury ceased!
ISA|14|5|The LORD has broken the staff of the wicked, the scepter of rulers,
ISA|14|6|that struck the peoples in wrath with unceasing blows, that ruled the nations in anger with unrelenting persecution.
ISA|14|7|The whole earth is at rest and quiet; they break forth into singing.
ISA|14|8|The cypresses rejoice at you, the cedars of Lebanon, saying, 'Since you were laid low, no woodcutter comes up against us.'
ISA|14|9|Sheol beneath is stirred up to meet you when you come; it rouses the shades to greet you, all who were leaders of the earth; it raises from their thrones all who were kings of the nations.
ISA|14|10|All of them will answer and say to you: 'You too have become as weak as we! You have become like us!'
ISA|14|11|Your pomp is brought down to Sheol, the sound of your harps; maggots are laid as a bed beneath you, and worms are your covers.
ISA|14|12|"How you are fallen from heaven, O Day Star, son of Dawn! How you are cut down to the ground, you who laid the nations low!
ISA|14|13|You said in your heart, 'I will ascend to heaven; above the stars of God I will set my throne on high; I will sit on the mount of assembly in the far reaches of the north;
ISA|14|14|I will ascend above the heights of the clouds; I will make myself like the Most High.'
ISA|14|15|But you are brought down to Sheol, to the far reaches of the pit.
ISA|14|16|Those who see you will stare at you and ponder over you: 'Is this the man who made the earth tremble, who shook kingdoms,
ISA|14|17|who made the world like a desert and overthrew its cities, who did not let his prisoners go home?'
ISA|14|18|All the kings of the nations lie in glory, each in his own tomb;
ISA|14|19|but you are cast out, away from your grave, like a loathed branch, clothed with the slain, those pierced by the sword, who go down to the stones of the pit, like a dead body trampled underfoot.
ISA|14|20|You will not be joined with them in burial, because you have destroyed your land, you have slain your people. "May the offspring of evildoers nevermore be named!
ISA|14|21|Prepare slaughter for his sons because of the guilt of their fathers, lest they rise and possess the earth, and fill the face of the world with cities."
ISA|14|22|"I will rise up against them," declares the LORD of hosts, "and will cut off from Babylon name and remnant, descendants and posterity," says the LORD.
ISA|14|23|"And I will make it a possession of the hedgehog, and pools of water, and I will sweep it with the broom of destruction," declares the LORD of hosts.
ISA|14|24|The LORD of hosts has sworn: "As I have planned, so shall it be, and as I have purposed, so shall it stand,
ISA|14|25|that I will break the Assyrian in my land, and on my mountains trample him underfoot; and his yoke shall depart from them, and his burden from their shoulder."
ISA|14|26|This is the purpose that is purposed concerning the whole earth, and this is the hand that is stretched out over all the nations.
ISA|14|27|For the LORD of hosts has purposed, and who will annul it? His hand is stretched out, and who will turn it back?
ISA|14|28|In the year that King Ahaz died came this oracle:
ISA|14|29|Rejoice not, O Philistia, all of you, that the rod that struck you is broken, for from the serpent's root will come forth an adder, and its fruit will be a flying fiery serpent.
ISA|14|30|And the firstborn of the poor will graze, and the needy lie down in safety; but I will kill your root with famine, and your remnant it will slay.
ISA|14|31|Wail, O gate; cry out, O city; melt in fear, O Philistia, all of you! For smoke comes out of the north, and there is no straggler in his ranks.
ISA|14|32|What will one answer the messengers of the nation? "The LORD has founded Zion, and in her the afflicted of his people find refuge."
ISA|15|1|An oracle concerning Moab. Because Ar of Moab is laid waste in a night, Moab is undone; because Kir of Moab is laid waste in a night, Moab is undone.
ISA|15|2|He has gone up to the temple, and to Dibon, to the high places to weep; over Nebo and over Medeba Moab wails. On every head is baldness; every beard is shorn;
ISA|15|3|in the streets they wear sackcloth; on the housetops and in the squares everyone wails and melts in tears.
ISA|15|4|Heshbon and Elealeh cry out; their voice is heard as far as Jahaz; therefore the armed men of Moab cry aloud; his soul trembles.
ISA|15|5|My heart cries out for Moab; her fugitives flee to Zoar, to Eglath-shelishiyah. For at the ascent of Luhith they go up weeping; on the road to Horonaim they raise a cry of destruction;
ISA|15|6|the waters of Nimrim are a desolation; the grass is withered, the vegetation fails, the greenery is no more.
ISA|15|7|Therefore the abundance they have gained and what they have laid up they carry away over the Brook of the Willows.
ISA|15|8|For a cry has gone around the land of Moab; her wailing reaches to Eglaim; her wailing reaches to Beer-elim.
ISA|15|9|For the waters of Dibon are full of blood; for I will bring upon Dibon even more, a lion for those of Moab who escape, for the remnant of the land.
ISA|16|1|Send the lamb to the ruler of the land, from Sela, by way of the desert, to the mount of the daughter of Zion.
ISA|16|2|Like fleeing birds, like a scattered nest, so are the daughters of Moab at the fords of the Arnon.
ISA|16|3|"Give counsel; grant justice; make your shade like night at the height of noon; shelter the outcasts; do not reveal the fugitive;
ISA|16|4|let the outcasts of Moab sojourn among you; be a shelter to them from the destroyer. When the oppressor is no more and destruction has ceased, and he who tramples underfoot has vanished from the land,
ISA|16|5|then a throne will be established in steadfast love, and on it will sit in faithfulness in the tent of David one who judges and seeks justice and is swift to do righteousness."
ISA|16|6|We have heard of the pride of Moab- how proud he is!- of his arrogance, his pride, and his insolence; in his idle boasting he is not right.
ISA|16|7|Therefore let Moab wail for Moab, let everyone wail. Mourn, utterly stricken, for the raisin cakes of Kir-hareseth.
ISA|16|8|For the fields of Heshbon languish, and the vine of Sibmah; the lords of the nations have struck down its branches, which reached to Jazer and strayed to the desert; its shoots spread abroad and passed over the sea.
ISA|16|9|Therefore I weep with the weeping of Jazer for the vine of Sibmah; I drench you with my tears, O Heshbon and Elealeh; for over your summer fruit and your harvest the shout has ceased.
ISA|16|10|And joy and gladness are taken away from the fruitful field, and in the vineyards no songs are sung, no cheers are raised; no treader treads out wine in the presses; I have put an end to the shouting.
ISA|16|11|Therefore my inner parts moan like a lyre for Moab, and my inmost self for Kir-hareseth.
ISA|16|12|And when Moab presents himself, when he wearies himself on the high place, when he comes to his sanctuary to pray, he will not prevail.
ISA|16|13|This is the word that the LORD spoke concerning Moab in the past.
ISA|16|14|But now the LORD has spoken, saying, "In three years, like the years of a hired worker, the glory of Moab will be brought into contempt, in spite of all his great multitude, and those who remain will be very few and feeble."
ISA|17|1|An oracle concerning Damascus. Behold, Damascus will cease to be a city and will become a heap of ruins.
ISA|17|2|The cities of Aroer are deserted; they will be for flocks, which will lie down, and none will make them afraid.
ISA|17|3|The fortress will disappear from Ephraim, and the kingdom from Damascus; and the remnant of Syria will be like the glory of the children of Israel, declares the LORD of hosts.
ISA|17|4|And in that day the glory of Jacob will be brought low, and the fat of his flesh will grow lean.
ISA|17|5|And it shall be as when the reaper gathers standing grain and his arm harvests the ears, and as when one gleans the ears of grain in the Valley of Rephaim.
ISA|17|6|Gleanings will be left in it, as when an olive tree is beaten- two or three berries in the top of the highest bough, four or five on the branches of a fruit tree, declares the LORD God of Israel.
ISA|17|7|In that day man will look to his Maker, and his eyes will look on the Holy One of Israel.
ISA|17|8|He will not look to the altars, the work of his hands, and he will not look on what his own fingers have made, either the Asherim or the altars of incense.
ISA|17|9|In that day their strong cities will be like the deserted places of the wooded heights and the hilltops, which they deserted because of the children of Israel, and there will be desolation.
ISA|17|10|For you have forgotten the God of your salvation and have not remembered the Rock of your refuge; therefore, though you plant pleasant plants and sow the vine-branch of a stranger,
ISA|17|11|though you make them grow on the day that you plant them, and make them blossom in the morning that you sow, yet the harvest will flee away in a day of grief and incurable pain.
ISA|17|12|Ah, the thunder of many peoples; they thunder like the thundering of the sea! Ah, the roar of nations; they roar like the roaring of mighty waters!
ISA|17|13|The nations roar like the roaring of many waters, but he will rebuke them, and they will flee far away, chased like chaff on the mountains before the wind and whirling dust before the storm.
ISA|17|14|At evening time, behold, terror! Before morning, they are no more! This is the portion of those who loot us, and the lot of those who plunder us.
ISA|18|1|Ah, land of whirring wings that is beyond the rivers of Cush,
ISA|18|2|which sends ambassadors by the sea, in vessels of papyrus on the waters! Go, you swift messengers, to a nation, tall and smooth, to a people feared near and far, a nation mighty and conquering, whose land the rivers divide.
ISA|18|3|All you inhabitants of the world, you who dwell on the earth, when a signal is raised on the mountains, look! When a trumpet is blown, hear!
ISA|18|4|For thus the LORD said to me: "I will quietly look from my dwelling like clear heat in sunshine, like a cloud of dew in the heat of harvest."
ISA|18|5|For before the harvest, when the blossom is over, and the flower becomes a ripening grape, he cuts off the shoots with pruning hooks, and the spreading branches he lops off and clears away.
ISA|18|6|They shall all of them be left to the birds of prey of the mountains and to the beasts of the earth. And the birds of prey will summer on them, and all the beasts of the earth will winter on them.
ISA|18|7|At that time tribute will be brought to the LORD of hosts from a people tall and smooth, from a people feared near and far, a nation mighty and conquering, whose land the rivers divide, to Mount Zion, the place of the name of the LORD of hosts.
ISA|19|1|An oracle concerning Egypt. Behold, the LORD is riding on a swift cloud and comes to Egypt; and the idols of Egypt will tremble at his presence, and the heart of the Egyptians will melt within them.
ISA|19|2|And I will stir up Egyptians against Egyptians, and they will fight, each against another and each against his neighbor, city against city, kingdom against kingdom;
ISA|19|3|and the spirit of the Egyptians within them will be emptied out, and I will confound their counsel; and they will inquire of the idols and the sorcerers, and the mediums and the necromancers;
ISA|19|4|and I will give over the Egyptians into the hand of a hard master, and a fierce king will rule over them, declares the Lord GOD of hosts.
ISA|19|5|And the waters of the sea will be dried up, and the river will be dry and parched,
ISA|19|6|and its canals will become foul, and the branches of Egypt's Nile will diminish and dry up, reeds and rushes will rot away.
ISA|19|7|There will be bare places by the Nile, on the brink of the Nile, and all that is sown by the Nile will be parched, will be driven away, and will be no more.
ISA|19|8|The fishermen will mourn and lament, all who cast a hook in the Nile; and they will languish who spread nets on the water.
ISA|19|9|The workers in combed flax will be in despair, and the weavers of white cotton.
ISA|19|10|Those who are the pillars of the land will be crushed, and all who work for pay will be grieved.
ISA|19|11|The princes of Zoan are utterly foolish; the wisest counselors of Pharaoh give stupid counsel. How can you say to Pharaoh, "I am a son of the wise, a son of ancient kings"?
ISA|19|12|Where then are your wise men? Let them tell you that they might know what the LORD of hosts has purposed against Egypt.
ISA|19|13|The princes of Zoan have become fools, and the princes of Memphis are deluded; those who are the cornerstones of her tribes have made Egypt stagger.
ISA|19|14|The LORD has mingled within her a spirit of confusion, and they will make Egypt stagger in all its deeds, as a drunken man staggers in his vomit.
ISA|19|15|And there will be nothing for Egypt that head or tail, palm branch or reed, may do.
ISA|19|16|In that day the Egyptians will be like women, and tremble with fear before the hand that the LORD of hosts shakes over them.
ISA|19|17|And the land of Judah will become a terror to the Egyptians. Everyone to whom it is mentioned will fear because of the purpose that the LORD of hosts has purposed against them.
ISA|19|18|In that day there will be five cities in the land of Egypt that speak the language of Canaan and swear allegiance to the LORD of hosts. One of these will be called the City of Destruction.
ISA|19|19|In that day there will be an altar to the LORD in the midst of the land of Egypt, and a pillar to the LORD at its border.
ISA|19|20|It will be a sign and a witness to the LORD of hosts in the land of Egypt. When they cry to the LORD because of oppressors, he will send them a savior and defender, and deliver them.
ISA|19|21|And the LORD will make himself known to the Egyptians, and the Egyptians will know the LORD in that day and worship with sacrifice and offering, and they will make vows to the LORD and perform them.
ISA|19|22|And the LORD will strike Egypt, striking and healing, and they will return to the LORD, and he will listen to their pleas for mercy and heal them.
ISA|19|23|In that day there will be a highway from Egypt to Assyria, and Assyria will come into Egypt, and Egypt into Assyria, and the Egyptians will worship with the Assyrians.
ISA|19|24|In that day Israel will be the third with Egypt and Assyria, a blessing in the midst of the earth,
ISA|19|25|whom the LORD of hosts has blessed, saying, "Blessed be Egypt my people, and Assyria the work of my hands, and Israel my inheritance."
ISA|20|1|In the year that the commander in chief, who was sent by Sargon the king of Assyria, came to Ashdod and fought against it and captured it-
ISA|20|2|at that time the LORD spoke by Isaiah the son of Amoz, saying, "Go, and loose the sackcloth from your waist and take off your sandals from your feet," and he did so, walking naked and barefoot.
ISA|20|3|Then the LORD said, "As my servant Isaiah has walked naked and barefoot for three years as a sign and a portent against Egypt and Cush,
ISA|20|4|so shall the king of Assyria lead away the Egyptian captives and the Cushite exiles, both the young and the old, naked and barefoot, with buttocks uncovered, the nakedness of Egypt.
ISA|20|5|Then they shall be dismayed and ashamed because of Cush their hope and of Egypt their boast.
ISA|20|6|And the inhabitants of this coastland will say in that day, 'Behold, this is what has happened to those in whom we hoped and to whom we fled for help to be delivered from the king of Assyria! And we, how shall we escape?'"
ISA|21|1|The oracle concerning the wilderness of the sea. As whirlwinds in the Negeb sweep on, it comes from the wilderness, from a terrible land.
ISA|21|2|A stern vision is told to me; the traitor betrays, and the destroyer destroys. Go up, O Elam; lay siege, O Media; all the sighing she has caused I bring to an end.
ISA|21|3|Therefore my loins are filled with anguish; pangs have seized me, like the pangs of a woman in labor; I am bowed down so that I cannot hear; I am dismayed so that I cannot see.
ISA|21|4|My heart staggers; horror has appalled me; the twilight I longed for has been turned for me into trembling.
ISA|21|5|They prepare the table, they spread the rugs, they eat, they drink. Arise, O princes; oil the shield!
ISA|21|6|For thus the Lord said to me: "Go, set a watchman; let him announce what he sees.
ISA|21|7|When he sees riders, horsemen in pairs, riders on donkeys, riders on camels, let him listen diligently, very diligently."
ISA|21|8|Then he who saw cried out: "Upon a watchtower I stand, O Lord, continually by day, and at my post I am stationed whole nights.
ISA|21|9|And behold, here come riders, horsemen in pairs!" And he answered, "Fallen, fallen is Babylon; and all the carved images of her gods he has shattered to the ground."
ISA|21|10|O my threshed and winnowed one, what I have heard from the LORD of hosts, the God of Israel, I announce to you.
ISA|21|11|The oracle concerning Dumah. One is calling to me from Seir, "Watchman, what time of the night? Watchman, what time of the night?"
ISA|21|12|The watchman says: "Morning comes, and also the night. If you will inquire, inquire; come back again."
ISA|21|13|The oracle concerning Arabia. In the thickets in Arabia you will lodge, O caravans of Dedanites.
ISA|21|14|To the thirsty bring water; meet the fugitive with bread, O inhabitants of the land of Tema.
ISA|21|15|For they have fled from the swords, from the drawn sword, from the bent bow, and from the press of battle.
ISA|21|16|For thus the Lord said to me, "Within a year, according to the years of a hired worker, all the glory of Kedar will come to an end.
ISA|21|17|And the remainder of the archers of the mighty men of the sons of Kedar will be few, for the LORD, the God of Israel, has spoken."
ISA|22|1|The oracle concerning the valley of vision. What do you mean that you have gone up, all of you, to the housetops,
ISA|22|2|you who are full of shoutings, tumultuous city, exultant town? Your slain are not slain with the sword or dead in battle.
ISA|22|3|All your leaders have fled together; without the bow they were captured. All of you who were found were captured, though they had fled far away.
ISA|22|4|Therefore I said: "Look away from me; let me weep bitter tears; do not labor to comfort me concerning the destruction of the daughter of my people."
ISA|22|5|For the Lord GOD of hosts has a day of tumult and trampling and confusion in the valley of vision, a battering down of walls and a shouting to the mountains.
ISA|22|6|And Elam bore the quiver with chariots and horsemen, and Kir uncovered the shield.
ISA|22|7|Your choicest valleys were full of chariots, and the horsemen took their stand at the gates.
ISA|22|8|He has taken away the covering of Judah. In that day you looked to the weapons of the House of the Forest,
ISA|22|9|and you saw that the breaches of the city of David were many. You collected the waters of the lower pool,
ISA|22|10|and you counted the houses of Jerusalem, and you broke down the houses to fortify the wall.
ISA|22|11|You made a reservoir between the two walls for the water of the old pool. But you did not look to him who did it, or see him who planned it long ago.
ISA|22|12|In that day the Lord GOD of hosts called for weeping and mourning, for baldness and wearing sackcloth;
ISA|22|13|and behold, joy and gladness, killing oxen and slaughtering sheep, eating flesh and drinking wine. "Let us eat and drink, for tomorrow we die."
ISA|22|14|The LORD of hosts has revealed himself in my ears: "Surely this iniquity will not be atoned for you until you die," says the Lord GOD of hosts.
ISA|22|15|Thus says the Lord GOD of hosts, "Come, go to this steward, to Shebna, who is over the household, and say to him:
ISA|22|16|What have you to do here, and whom have you here, that you have cut out here a tomb for yourself, you who cut out a tomb on the height and carve a dwelling for yourself in the rock?
ISA|22|17|Behold, the LORD will hurl you away violently, O you strong man. He will seize firm hold on you
ISA|22|18|and whirl you around and around, and throw you like a ball into a wide land. There you shall die, and there shall be your glorious chariots, you shame of your master's house.
ISA|22|19|I will thrust you from your office, and you will be pulled down from your station.
ISA|22|20|In that day I will call my servant Eliakim the son of Hilkiah,
ISA|22|21|and I will clothe him with your robe, and will bind your sash on him, and will commit your authority to his hand. And he shall be a father to the inhabitants of Jerusalem and to the house of Judah.
ISA|22|22|And I will place on his shoulder the key of the house of David. He shall open, and none shall shut; and he shall shut, and none shall open.
ISA|22|23|And I will fasten him like a peg in a secure place, and he will become a throne of honor to his father's house.
ISA|22|24|And they will hang on him the whole honor of his father's house, the offspring and issue, every small vessel, from the cups to all the flagons.
ISA|22|25|In that day, declares the LORD of hosts, the peg that was fastened in a secure place will give way, and it will be cut down and fall, and the load that was on it will be cut off, for the LORD has spoken."
ISA|23|1|The oracle concerning Tyre. Wail, O ships of Tarshish, for Tyre is laid waste, without house or harbor! From the land of Cyprus it is revealed to them.
ISA|23|2|Be still, O inhabitants of the coast; the merchants of Sidon, who cross the sea, have filled you.
ISA|23|3|And on many waters your revenue was the grain of Shihor, the harvest of the Nile; you were the merchant of the nations.
ISA|23|4|Be ashamed, O Sidon, for the sea has spoken, the stronghold of the sea, saying: "I have neither labored nor given birth, I have neither reared young men nor brought up young women."
ISA|23|5|When the report comes to Egypt, they will be in anguish over the report about Tyre.
ISA|23|6|Cross over to Tarshish; wail, O inhabitants of the coast!
ISA|23|7|Is this your exultant city whose origin is from days of old, whose feet carried her to settle far away?
ISA|23|8|Who has purposed this against Tyre, the bestower of crowns, whose merchants were princes, whose traders were the honored of the earth?
ISA|23|9|The LORD of hosts has purposed it, to defile the pompous pride of all glory, to dishonor all the honored of the earth.
ISA|23|10|Cross over your land like the Nile, O daughter of Tarshish; there is no restraint anymore.
ISA|23|11|He has stretched out his hand over the sea; he has shaken the kingdoms; the LORD has given command concerning Canaan to destroy its strongholds.
ISA|23|12|And he said: "You will no more exult, O oppressed virgin daughter of Sidon; arise, cross over to Cyprus, even there you will have no rest."
ISA|23|13|Behold the land of the Chaldeans! This is the people that was not; Assyria destined it for wild beasts. They erected their siege towers, they stripped her palaces bare, they made her a ruin.
ISA|23|14|Wail, O ships of Tarshish, for your stronghold is laid waste.
ISA|23|15|In that day Tyre will be forgotten for seventy years, like the days of one king. At the end of seventy years, it will happen to Tyre as in the song of the prostitute:
ISA|23|16|"Take a harp; go about the city, O forgotten prostitute! Make sweet melody; sing many songs, that you may be remembered."
ISA|23|17|At the end of seventy years, the LORD will visit Tyre, and she will return to her wages and will prostitute herself with all the kingdoms of the world on the face of the earth.
ISA|23|18|Her merchandise and her wages will be holy to the LORD. It will not be stored or hoarded, but her merchandise will supply abundant food and fine clothing for those who dwell before the LORD.
ISA|24|1|Behold, the LORD will empty the earth and make it desolate, and he will twist its surface and scatter its inhabitants.
ISA|24|2|And it shall be, as with the people, so with the priest; as with the slave, so with his master; as with the maid, so with her mistress; as with the buyer, so with the seller; as with the lender, so with the borrower; as with the creditor, so with the debtor.
ISA|24|3|The earth shall be utterly empty and utterly plundered; for the LORD has spoken this word.
ISA|24|4|The earth mourns and withers; the world languishes and withers; the highest people of the earth languish.
ISA|24|5|The earth lies defiled under its inhabitants; for they have transgressed the laws, violated the statutes, broken the everlasting covenant.
ISA|24|6|Therefore a curse devours the earth, and its inhabitants suffer for their guilt; therefore the inhabitants of the earth are scorched, and few men are left.
ISA|24|7|The wine mourns, the vine languishes, all the merry-hearted sigh.
ISA|24|8|The mirth of the tambourines is stilled, the noise of the jubilant has ceased, the mirth of the lyre is stilled.
ISA|24|9|No more do they drink wine with singing; strong drink is bitter to those who drink it.
ISA|24|10|The wasted city is broken down; every house is shut up so that none can enter.
ISA|24|11|There is an outcry in the streets for lack of wine; all joy has grown dark; the gladness of the earth is banished.
ISA|24|12|Desolation is left in the city; the gates are battered into ruins.
ISA|24|13|For thus it shall be in the midst of the earth among the nations, as when an olive tree is beaten, as at the gleaning when the grape harvest is done.
ISA|24|14|They lift up their voices, they sing for joy; over the majesty of the LORD they shout from the west.
ISA|24|15|Therefore in the east give glory to the LORD; in the coastlands of the sea, give glory to the name of the LORD, the God of Israel.
ISA|24|16|From the ends of the earth we hear songs of praise, of glory to the Righteous One. But I say, "I waste away, I waste away. Woe is me! For the traitors have betrayed, with betrayal the traitors have betrayed."
ISA|24|17|Terror and the pit and the snare are upon you, O inhabitant of the earth!
ISA|24|18|He who flees at the sound of the terror shall fall into the pit, and he who climbs out of the pit shall be caught in the snare. For the windows of heaven are opened, and the foundations of the earth tremble.
ISA|24|19|The earth is utterly broken, the earth is split apart, the earth is violently shaken.
ISA|24|20|The earth staggers like a drunken man; it sways like a hut; its transgression lies heavy upon it, and it falls, and will not rise again.
ISA|24|21|On that day the LORD will punish the host of heaven, in heaven, and the kings of the earth, on the earth.
ISA|24|22|They will be gathered together as prisoners in a pit; they will be shut up in a prison, and after many days they will be punished.
ISA|24|23|Then the moon will be confounded and the sun ashamed, for the LORD of hosts reigns on Mount Zion and in Jerusalem, and his glory will be before his elders.
ISA|25|1|O LORD, you are my God; I will exalt you; I will praise your name, for you have done wonderful things, plans formed of old, faithful and sure.
ISA|25|2|For you have made the city a heap, the fortified city a ruin; the foreigners' palace is a city no more; it will never be rebuilt.
ISA|25|3|Therefore strong peoples will glorify you; cities of ruthless nations will fear you.
ISA|25|4|For you have been a stronghold to the poor, a stronghold to the needy in his distress, a shelter from the storm and a shade from the heat; for the breath of the ruthless is like a storm against a wall,
ISA|25|5|like heat in a dry place. You subdue the noise of the foreigners; as heat by the shade of a cloud, so the song of the ruthless is put down.
ISA|25|6|On this mountain the LORD of hosts will make for all peoples a feast of rich food, a feast of well-aged wine, of rich food full of marrow, of aged wine well refined.
ISA|25|7|And he will swallow up on this mountain the covering that is cast over all peoples, the veil that is spread over all nations.
ISA|25|8|He will swallow up death forever; and the Lord GOD will wipe away tears from all faces, and the reproach of his people he will take away from all the earth, for the LORD has spoken.
ISA|25|9|It will be said on that day, "Behold, this is our God; we have waited for him, that he might save us. This is the LORD; we have waited for him; let us be glad and rejoice in his salvation."
ISA|25|10|For the hand of the LORD will rest on this mountain, and Moab shall be trampled down in his place, as straw is trampled down in a dunghill.
ISA|25|11|And he will spread out his hands in the midst of it as a swimmer spreads his hands out to swim, but the LORD will lay low his pompous pride together with the skill of his hands.
ISA|25|12|And the high fortifications of his walls he will bring down, lay low, and cast to the ground, to the dust.
ISA|26|1|In that day this song will be sung in the land of Judah: "We have a strong city; he sets up salvation as walls and bulwarks.
ISA|26|2|Open the gates, that the righteous nation that keeps faith may enter in.
ISA|26|3|You keep him in perfect peace whose mind is stayed on you, because he trusts in you.
ISA|26|4|Trust in the LORD forever, for the LORD GOD is an everlasting rock.
ISA|26|5|For he has humbled the inhabitants of the height, the lofty city. He lays it low, lays it low to the ground, casts it to the dust.
ISA|26|6|The foot tramples it, the feet of the poor, the steps of the needy."
ISA|26|7|The path of the righteous is level; you make level the way of the righteous.
ISA|26|8|In the path of your judgments, O LORD, we wait for you; your name and remembrance are the desire of our soul.
ISA|26|9|My soul yearns for you in the night; my spirit within me earnestly seeks you. For when your judgments are in the earth, the inhabitants of the world learn righteousness.
ISA|26|10|If favor is shown to the wicked, he does not learn righteousness; in the land of uprightness he deals corruptly and does not see the majesty of the LORD.
ISA|26|11|O LORD, your hand is lifted up, but they do not see it. Let them see your zeal for your people, and be ashamed. Let the fire for your adversaries consume them.
ISA|26|12|O LORD, you will ordain peace for us; you have done for us all our works.
ISA|26|13|O LORD our God, other lords besides you have ruled over us, but your name alone we bring to remembrance.
ISA|26|14|They are dead, they will not live; they are shades, they will not arise; to that end you have visited them with destruction and wiped out all remembrance of them.
ISA|26|15|But you have increased the nation, O LORD, you have increased the nation; you are glorified; you have enlarged all the borders of the land.
ISA|26|16|O LORD, in distress they sought you; they poured out a whispered prayer when your discipline was upon them.
ISA|26|17|Like a pregnant woman who writhes and cries out in her pangs when she is near to giving birth, so were we because of you, O LORD;
ISA|26|18|we were pregnant, we writhed, but we have given birth to wind. We have accomplished no deliverance in the earth, and the inhabitants of the world have not fallen.
ISA|26|19|Your dead shall live; their bodies shall rise. You who dwell in the dust, awake and sing for joy! For your dew is a dew of light, and the earth will give birth to the dead.
ISA|26|20|Come, my people, enter your chambers, and shut your doors behind you; hide yourselves for a little while until the fury has passed by.
ISA|26|21|For behold, the LORD is coming out from his place to punish the inhabitants of the earth for their iniquity, and the earth will disclose the blood shed on it, and will no more cover its slain.
ISA|27|1|In that day the LORD with his hard and great and strong sword will punish Leviathan the fleeing serpent, Leviathan the twisting serpent, and he will slay the dragon that is in the sea.
ISA|27|2|In that day, "A pleasant vineyard, sing of it!
ISA|27|3|I, the LORD, am its keeper; every moment I water it. Lest anyone punish it, I keep it night and day;
ISA|27|4|I have no wrath. Would that I had thorns and briers to battle! I would march against them, I would burn them up together.
ISA|27|5|Or let them lay hold of my protection, let them make peace with me, let them make peace with me."
ISA|27|6|In days to come Jacob shall take root, Israel shall blossom and put forth shoots and fill the whole world with fruit.
ISA|27|7|Has he struck them as he struck those who struck them? Or have they been slain as their slayers were slain?
ISA|27|8|Measure by measure, by exile you contended with them; he removed them with his fierce breath in the day of the east wind.
ISA|27|9|Therefore by this the guilt of Jacob will be atoned for, and this will be the full fruit of the removal of his sin: when he makes all the stones of the altars like chalkstones crushed to pieces, no Asherim or incense altars will remain standing.
ISA|27|10|For the fortified city is solitary, a habitation deserted and forsaken, like the wilderness; there the calf grazes; there it lies down and strips its branches.
ISA|27|11|When its boughs are dry, they are broken; women come and make a fire of them. For this is a people without discernment; therefore he who made them will not have compassion on them; he who formed them will show them no favor.
ISA|27|12|In that day from the river Euphrates to the Brook of Egypt the LORD will thresh out the grain, and you will be gleaned one by one, O people of Israel.
ISA|27|13|And in that day a great trumpet will be blown, and those who were lost in the land of Assyria and those who were driven out to the land of Egypt will come and worship the LORD on the holy mountain at Jerusalem.
ISA|28|1|Ah, the proud crown of the drunkards of Ephraim, and the fading flower of its glorious beauty, which is on the head of the rich valley of those overcome with wine!
ISA|28|2|Behold, the Lord has one who is mighty and strong; like a storm of hail, a destroying tempest, like a storm of mighty, overflowing waters, he casts down to the earth with his hand.
ISA|28|3|The proud crown of the drunkards of Ephraim will be trodden underfoot;
ISA|28|4|and the fading flower of its glorious beauty, which is on the head of the rich valley, will be like a first-ripe fig before the summer: when someone sees it, he swallows it as soon as it is in his hand.
ISA|28|5|In that day the LORD of hosts will be a crown of glory, and a diadem of beauty, to the remnant of his people,
ISA|28|6|and a spirit of justice to him who sits in judgment, and strength to those who turn back the battle at the gate.
ISA|28|7|These also reel with wine and stagger with strong drink; the priest and the prophet reel with strong drink, they are swallowed by wine, they stagger with strong drink, they reel in vision, they stumble in giving judgment.
ISA|28|8|For all tables are full of filthy vomit, with no space left.
ISA|28|9|"To whom will he teach knowledge, and to whom will he explain the message? Those who are weaned from the milk, those taken from the breast?
ISA|28|10|For it is precept upon precept, precept upon precept, line upon line, line upon line, here a little, there a little."
ISA|28|11|For by people of strange lips and with a foreign tongue the LORD will speak to this people,
ISA|28|12|to whom he has said, "This is rest; give rest to the weary; and this is repose"; yet they would not hear.
ISA|28|13|And the word of the LORD will be to them precept upon precept, precept upon precept, line upon line, line upon line, here a little, there a little, that they may go, and fall backward, and be broken, and snared, and taken.
ISA|28|14|Therefore hear the word of the LORD, you scoffers, who rule this people in Jerusalem!
ISA|28|15|Because you have said, "We have made a covenant with death, and with Sheol we have an agreement, when the overwhelming whip passes through it will not come to us, for we have made lies our refuge, and in falsehood we have taken shelter";
ISA|28|16|therefore thus says the Lord GOD, "Behold, I am the one who has laid as a foundation in Zion, a stone, a tested stone, a precious cornerstone, of a sure foundation: 'Whoever believes will not be in haste.'
ISA|28|17|And I will make justice the line, and righteousness the plumb line; and hail will sweep away the refuge of lies, and waters will overwhelm the shelter."
ISA|28|18|Then your covenant with death will be annulled, and your agreement with Sheol will not stand; when the overwhelming scourge passes through, you will be beaten down by it.
ISA|28|19|As often as it passes through it will take you; for morning by morning it will pass through, by day and by night; and it will be sheer terror to understand the message.
ISA|28|20|For the bed is too short to stretch oneself on, and the covering too narrow to wrap oneself in.
ISA|28|21|For the LORD will rise up as on Mount Perazim; as in the Valley of Gibeon he will be roused; to do his deed- strange is his deed! and to work his work- alien is his work!
ISA|28|22|Now therefore do not scoff, lest your bonds be made strong; for I have heard a decree of destruction from the Lord GOD of hosts against the whole land.
ISA|28|23|Give ear, and hear my voice; give attention, and hear my speech.
ISA|28|24|Does he who plows for sowing plow continually? does he continually open and harrow his ground?
ISA|28|25|When he has leveled its surface, does he not scatter dill, sow cumin, and put in wheat in rows and barley in its proper place, and emmer as the border?
ISA|28|26|For he is rightly instructed; his God teaches him.
ISA|28|27|Dill is not threshed with a threshing sledge, nor is a cart wheel rolled over cumin, but dill is beaten out with a stick, and cumin with a rod.
ISA|28|28|Does one crush grain for bread? No, he does not thresh it forever; when he drives his cart wheel over it with his horses, he does not crush it.
ISA|28|29|This also comes from the LORD of hosts; he is wonderful in counsel and excellent in wisdom.
ISA|29|1|Ah, Ariel, Ariel, the city where David encamped! Add year to year; let the feasts run their round.
ISA|29|2|Yet I will distress Ariel, and there shall be moaning and lamentation, and she shall be to me like an Ariel.
ISA|29|3|And I will encamp against you all around, and will besiege you with towers and I will raise siegeworks against you.
ISA|29|4|And you will be brought low; from the earth you shall speak, and from the dust your speech will be bowed down; your voice shall come from the ground like the voice of a ghost, and from the dust your speech shall whisper.
ISA|29|5|But the multitude of your foreign foes shall be like small dust, and the multitude of the ruthless like passing chaff. And in an instant, suddenly,
ISA|29|6|you will be visited by the LORD of hosts with thunder and with earthquake and great noise, with whirlwind and tempest, and the flame of a devouring fire.
ISA|29|7|And the multitude of all the nations that fight against Ariel, all that fight against her and her stronghold and distress her, shall be like a dream, a vision of the night.
ISA|29|8|As when a hungry man dreams he is eating and awakes with his hunger not satisfied, or as when a thirsty man dreams he is drinking and awakes faint, with his thirst not quenched, so shall the multitude of all the nations be that fight against Mount Zion.
ISA|29|9|Astonish yourselves and be astonished; blind yourselves and be blind! Be drunk, but not with wine; stagger, but not with strong drink!
ISA|29|10|For the LORD has poured out upon you a spirit of deep sleep, and has closed your eyes (the prophets), and covered your heads (the seers).
ISA|29|11|And the vision of all this has become to you like the words of a book that is sealed. When men give it to one who can read, saying, "Read this," he says, "I cannot, for it is sealed."
ISA|29|12|And when they give the book to one who cannot read, saying, "Read this," he says, "I cannot read."
ISA|29|13|And the Lord said: "Because this people draw near with their mouth and honor me with their lips, while their hearts are far from me, and their fear of me is a commandment taught by men,
ISA|29|14|therefore, behold, I will again do wonderful things with this people, with wonder upon wonder; and the wisdom of their wise men shall perish, and the discernment of their discerning men shall be hidden."
ISA|29|15|Ah, you who hide deep from the LORD your counsel, whose deeds are in the dark, and who say, "Who sees us? Who knows us?"
ISA|29|16|You turn things upside down! Shall the potter be regarded as the clay, that the thing made should say of its maker, "He did not make me"; or the thing formed say of him who formed it, "He has no understanding"?
ISA|29|17|Is it not yet a very little while until Lebanon shall be turned into a fruitful field, and the fruitful field shall be regarded as a forest?
ISA|29|18|In that day the deaf shall hear the words of a book, and out of their gloom and darkness the eyes of the blind shall see.
ISA|29|19|The meek shall obtain fresh joy in the LORD, and the poor among mankind shall exult in the Holy One of Israel.
ISA|29|20|For the ruthless shall come to nothing and the scoffer cease, and all who watch to do evil shall be cut off,
ISA|29|21|who by a word make a man out to be an offender, and lay a snare for him who reproves in the gate, and with an empty plea turn aside him who is in the right.
ISA|29|22|Therefore thus says the LORD, who redeemed Abraham, concerning the house of Jacob: "Jacob shall no more be ashamed, no more shall his face grow pale.
ISA|29|23|For when he sees his children, the work of my hands, in his midst, they will sanctify my name; they will sanctify the Holy One of Jacob and will stand in awe of the God of Israel.
ISA|29|24|And those who go astray in spirit will come to understanding, and those who murmur will accept instruction."
ISA|30|1|"Ah, stubborn children," declares the LORD, "who carry out a plan, but not mine, and who make an alliance, but not of my Spirit, that they may add sin to sin;
ISA|30|2|who set out to go down to Egypt, without asking for my direction, to take refuge in the protection of Pharaoh and to seek shelter in the shadow of Egypt!
ISA|30|3|Therefore shall the protection of Pharaoh turn to your shame, and the shelter in the shadow of Egypt to your humiliation.
ISA|30|4|For though his officials are at Zoan and his envoys reach Hanes,
ISA|30|5|everyone comes to shame through a people that cannot profit them, that brings neither help nor profit, but shame and disgrace."
ISA|30|6|An oracle on the beasts of the Negeb. Through a land of trouble and anguish, from where come the lioness and the lion, the adder and the flying fiery serpent, they carry their riches on the backs of donkeys, and their treasures on the humps of camels, to a people that cannot profit them.
ISA|30|7|Egypt's help is worthless and empty; therefore I have called her "Rahab who sits still."
ISA|30|8|And now, go, write it before them on a tablet and inscribe it in a book, that it may be for the time to come as a witness forever.
ISA|30|9|For they are a rebellious people, lying children, children unwilling to hear the instruction of the LORD;
ISA|30|10|who say to the seers, "Do not see," and to the prophets, "Do not prophesy to us what is right; speak to us smooth things, prophesy illusions,
ISA|30|11|leave the way, turn aside from the path, let us hear no more about the Holy One of Israel."
ISA|30|12|Therefore thus says the Holy One of Israel, "Because you despise this word and trust in oppression and perverseness and rely on them,
ISA|30|13|therefore this iniquity shall be to you like a breach in a high wall, bulging out, and about to collapse, whose breaking comes suddenly, in an instant;
ISA|30|14|and its breaking is like that of a potter's vessel that is smashed so ruthlessly that among its fragments not a shard is found with which to take fire from the hearth, or to dip up water out of the cistern."
ISA|30|15|For thus said the Lord GOD, the Holy One of Israel, "In returning and rest you shall be saved; in quietness and in trust shall be your strength." But you were unwilling,
ISA|30|16|and you said, "No! We will flee upon horses"; therefore you shall flee away; and, "We will ride upon swift steeds"; therefore your pursuers shall be swift.
ISA|30|17|A thousand shall flee at the threat of one; at the threat of five you shall flee, till you are left like a flagstaff on the top of a mountain, like a signal on a hill.
ISA|30|18|Therefore the LORD waits to be gracious to you, and therefore he exalts himself to show mercy to you. For the LORD is a God of justice; blessed are all those who wait for him.
ISA|30|19|For a people shall dwell in Zion, in Jerusalem; you shall weep no more. He will surely be gracious to you at the sound of your cry. As soon as he hears it, he answers you.
ISA|30|20|And though the Lord give you the bread of adversity and the water of affliction, yet your Teacher will not hide himself anymore, but your eyes shall see your Teacher.
ISA|30|21|And your ears shall hear a word behind you, saying, "This is the way, walk in it," when you turn to the right or when you turn to the left.
ISA|30|22|Then you will defile your carved idols overlaid with silver and your gold-plated metal images. You will scatter them as unclean things. You will say to them, "Be gone!"
ISA|30|23|And he will give rain for the seed with which you sow the ground, and bread, the produce of the ground, which will be rich and plenteous. In that day your livestock will graze in large pastures,
ISA|30|24|and the oxen and the donkeys that work the ground will eat seasoned fodder, which has been winnowed with shovel and fork.
ISA|30|25|And on every lofty mountain and every high hill there will be brooks running with water, in the day of the great slaughter, when the towers fall.
ISA|30|26|Moreover, the light of the moon will be as the light of the sun, and the light of the sun will be sevenfold, as the light of seven days, in the day when the LORD binds up the brokenness of his people, and heals the wounds inflicted by his blow.
ISA|30|27|Behold, the name of the LORD comes from far, burning with his anger, and in thick rising smoke; his lips are full of fury, and his tongue is like a devouring fire;
ISA|30|28|his breath is like an overflowing stream that reaches up to the neck; to sift the nations with the sieve of destruction, and to place on the jaws of the peoples a bridle that leads astray.
ISA|30|29|You shall have a song as in the night when a holy feast is kept, and gladness of heart, as when one sets out to the sound of the flute to go to the mountain of the LORD, to the Rock of Israel.
ISA|30|30|And the LORD will cause his majestic voice to be heard and the descending blow of his arm to be seen, in furious anger and a flame of devouring fire, with a cloudburst and storm and hailstones.
ISA|30|31|The Assyrians will be terror-stricken at the voice of the LORD, when he strikes with his rod.
ISA|30|32|And every stroke of the appointed staff that the LORD lays on them will be to the sound of tambourines and lyres. Battling with brandished arm, he will fight with them.
ISA|30|33|For a burning place has long been prepared; indeed, for the king it is made ready, its pyre made deep and wide, with fire and wood in abundance; the breath of the LORD, like a stream of sulfur, kindles it.
ISA|31|1|Woe to those who go down to Egypt for help and rely on horses, who trust in chariots because they are many and in horsemen because they are very strong, but do not look to the Holy One of Israel or consult the LORD!
ISA|31|2|And yet he is wise and brings disaster; he does not call back his words, but will arise against the house of the evildoers and against the helpers of those who work iniquity.
ISA|31|3|The Egyptians are man, and not God, and their horses are flesh, and not spirit. When the LORD stretches out his hand, the helper will stumble, and he who is helped will fall, and they will all perish together.
ISA|31|4|For thus the LORD said to me, "As a lion or a young lion growls over his prey, and when a band of shepherds is called out against him is not terrified by their shouting or daunted at their noise, so the LORD of hosts will come down to fight on Mount Zion and on its hill.
ISA|31|5|Like birds hovering, so the LORD of hosts will protect Jerusalem; he will protect and deliver it; he will spare and rescue it."
ISA|31|6|Turn to him from whom people have deeply revolted, O children of Israel.
ISA|31|7|For in that day everyone shall cast away his idols of silver and his idols of gold, which your hands have sinfully made for you.
ISA|31|8|"And the Assyrian shall fall by a sword, not of man; and a sword, not of man, shall devour him; and he shall flee from the sword, and his young men shall be put to forced labor.
ISA|31|9|His rock shall pass away in terror, and his officers desert the standard in panic," declares the LORD, whose fire is in Zion, and whose furnace is in Jerusalem.
ISA|32|1|Behold, a king will reign in righteousness, and princes will rule in justice.
ISA|32|2|Each will be like a hiding place from the wind, a shelter from the storm, like streams of water in a dry place, like the shade of a great rock in a weary land.
ISA|32|3|Then the eyes of those who see will not be closed, and the ears of those who hear will give attention.
ISA|32|4|The heart of the hasty will understand and know, and the tongue of the stammerers will hasten to speak distinctly.
ISA|32|5|The fool will no more be called noble, nor the scoundrel said to be honorable.
ISA|32|6|For the fool speaks folly, and his heart is busy with iniquity, to practice ungodliness, to utter error concerning the LORD, to leave the craving of the hungry unsatisfied, and to deprive the thirsty of drink.
ISA|32|7|As for the scoundrel- his devices are evil; he plans wicked schemes to ruin the poor with lying words, even when the plea of the needy is right.
ISA|32|8|But he who is noble plans noble things, and on noble things he stands.
ISA|32|9|Rise up, you women who are at ease, hear my voice; you complacent daughters, give ear to my speech.
ISA|32|10|In little more than a year you will shudder, you complacent women; for the grape harvest fails, the fruit harvest will not come.
ISA|32|11|Tremble, you women who are at ease, shudder, you complacent ones; strip, and make yourselves bare, and tie sackcloth around your waist.
ISA|32|12|Beat your breasts for the pleasant fields, for the fruitful vine,
ISA|32|13|for the soil of my people growing up in thorns and briers, yes, for all the joyous houses in the exultant city.
ISA|32|14|For the palace is forsaken, the populous city deserted; the hill and the watchtower will become dens forever, a joy of wild donkeys, a pasture of flocks;
ISA|32|15|until the Spirit is poured upon us from on high, and the wilderness becomes a fruitful field, and the fruitful field is deemed a forest.
ISA|32|16|Then justice will dwell in the wilderness, and righteousness abide in the fruitful field.
ISA|32|17|And the effect of righteousness will be peace, and the result of righteousness, quietness and trust forever.
ISA|32|18|My people will abide in a peaceful habitation, in secure dwellings, and in quiet resting places.
ISA|32|19|And it will hail when the forest falls down, and the city will be utterly laid low.
ISA|32|20|Happy are you who sow beside all waters, who let the feet of the ox and the donkey range free.
ISA|33|1|Ah, you destroyer, who yourself have not been destroyed, you traitor, whom none has betrayed! When you have ceased to destroy, you will be destroyed; and when you have finished betraying, they will betray you.
ISA|33|2|O LORD, be gracious to us; we wait for you. Be our arm every morning, our salvation in the time of trouble.
ISA|33|3|At the tumultuous noise peoples flee; when you lift yourself up, nations are scattered,
ISA|33|4|and your spoil is gathered as the caterpillar gathers; as locusts leap, it is leapt upon.
ISA|33|5|The LORD is exalted, for he dwells on high; he will fill Zion with justice and righteousness,
ISA|33|6|and he will be the stability of your times, abundance of salvation, wisdom, and knowledge; the fear of the LORD is Zion's treasure.
ISA|33|7|Behold, their heroes cry in the streets; the envoys of peace weep bitterly.
ISA|33|8|The highways lie waste; the traveler ceases. Covenants are broken; cities are despised; there is no regard for man.
ISA|33|9|The land mourns and languishes; Lebanon is confounded and withers away; Sharon is like a desert, and Bashan and Carmel shake off their leaves.
ISA|33|10|"Now I will arise," says the LORD, "now I will lift myself up; now I will be exalted.
ISA|33|11|You conceive chaff; you give birth to stubble; your breath is a fire that will consume you.
ISA|33|12|And the peoples will be as if burned to lime, like thorns cut down, that are burned in the fire."
ISA|33|13|Hear, you who are far off, what I have done; and you who are near, acknowledge my might.
ISA|33|14|The sinners in Zion are afraid; trembling has seized the godless: "Who among us can dwell with the consuming fire? Who among us can dwell with everlasting burnings?"
ISA|33|15|He who walks righteously and speaks uprightly, who despises the gain of oppressions, who shakes his hands, lest they hold a bribe, who stops his ears from hearing of bloodshed and shuts his eyes from looking on evil,
ISA|33|16|he will dwell on the heights; his place of defense will be the fortresses of rocks; his bread will be given him; his water will be sure.
ISA|33|17|Your eyes will behold the king in his beauty; they will see a land that stretches afar.
ISA|33|18|Your heart will muse on the terror: "Where is he who counted, where is he who weighed the tribute? Where is he who counted the towers?"
ISA|33|19|You will see no more the insolent people, the people of an obscure speech that you cannot comprehend, stammering in a tongue that you cannot understand.
ISA|33|20|Behold Zion, the city of our appointed feasts! Your eyes will see Jerusalem, an untroubled habitation, an immovable tent, whose stakes will never be plucked up, nor will any of its cords be broken.
ISA|33|21|But there the LORD in majesty will be for us a place of broad rivers and streams, where no galley with oars can go, nor majestic ship can pass.
ISA|33|22|For the LORD is our judge; the LORD is our lawgiver; the LORD is our king; he will save us.
ISA|33|23|Your cords hang loose; they cannot hold the mast firm in its place or keep the sail spread out. Then prey and spoil in abundance will be divided; even the lame will take the prey.
ISA|33|24|And no inhabitant will say, "I am sick"; the people who dwell there will be forgiven their iniquity.
ISA|34|1|Draw near, O nations, to hear, and give attention, O peoples! Let the earth hear, and all that fills it; the world, and all that comes from it.
ISA|34|2|For the LORD is enraged against all the nations, and furious against all their host; he has devoted them to destruction, has given them over for slaughter.
ISA|34|3|Their slain shall be cast out, and the stench of their corpses shall rise; the mountains shall flow with their blood.
ISA|34|4|All the host of heaven shall rot away, and the skies roll up like a scroll. All their host shall fall, as leaves fall from the vine, like leaves falling from the fig tree.
ISA|34|5|For my sword has drunk its fill in the heavens; behold, it descends for judgment upon Edom, upon the people I have devoted to destruction.
ISA|34|6|The LORD has a sword; it is sated with blood; it is gorged with fat, with the blood of lambs and goats, with the fat of the kidneys of rams. For the LORD has a sacrifice in Bozrah, a great slaughter in the land of Edom.
ISA|34|7|Wild oxen shall fall with them, and young steers with the mighty bulls. Their land shall drink its fill of blood, and their soil shall be gorged with fat.
ISA|34|8|For the LORD has a day of vengeance, a year of recompense for the cause of Zion.
ISA|34|9|And the streams of Edom shall be turned into pitch, and her soil into sulfur; her land shall become burning pitch.
ISA|34|10|Night and day it shall not be quenched; its smoke shall go up forever. From generation to generation it shall lie waste; none shall pass through it forever and ever.
ISA|34|11|But the hawk and the porcupine shall possess it, the owl and the raven shall dwell in it. He shall stretch the line of confusion over it, and the plumb line of emptiness.
ISA|34|12|Its nobles- there is no one there to call it a kingdom, and all its princes shall be nothing.
ISA|34|13|Thorns shall grow over its strongholds, nettles and thistles in its fortresses. It shall be the haunt of jackals, an abode for ostriches.
ISA|34|14|And wild animals shall meet with hyenas; the wild goat shall cry to his fellow; indeed, there the night bird settles and finds for herself a resting place.
ISA|34|15|There the owl nests and lays and hatches and gathers her young in her shadow; indeed, there the hawks are gathered, each one with her mate.
ISA|34|16|Seek and read from the book of the LORD: Not one of these shall be missing; none shall be without her mate. For the mouth of the LORD has commanded, and his Spirit has gathered them.
ISA|34|17|He has cast the lot for them; his hand has portioned it out to them with the line; they shall possess it forever; from generation to generation they shall dwell in it.
ISA|35|1|The wilderness and the dry land shall be glad; the desert shall rejoice and blossom like the crocus;
ISA|35|2|it shall blossom abundantly and rejoice with joy and singing. The glory of Lebanon shall be given to it, the majesty of Carmel and Sharon. They shall see the glory of the LORD, the majesty of our God.
ISA|35|3|Strengthen the weak hands, and make firm the feeble knees.
ISA|35|4|Say to those who have an anxious heart, "Be strong; fear not! Behold, your God will come with vengeance, with the recompense of God. He will come and save you."
ISA|35|5|Then the eyes of the blind shall be opened, and the ears of the deaf unstopped;
ISA|35|6|then shall the lame man leap like a deer, and the tongue of the mute sing for joy. For waters break forth in the wilderness, and streams in the desert;
ISA|35|7|the burning sand shall become a pool, and the thirsty ground springs of water; in the haunt of jackals, where they lie down, the grass shall become reeds and rushes.
ISA|35|8|And a highway shall be there, and it shall be called the Way of Holiness; the unclean shall not pass over it. It shall belong to those who walk on the way; even if they are fools, they shall not go astray.
ISA|35|9|No lion shall be there, nor shall any ravenous beast come up on it; they shall not be found there, but the redeemed shall walk there.
ISA|35|10|And the ransomed of the LORD shall return and come to Zion with singing; everlasting joy shall be upon their heads; they shall obtain gladness and joy, and sorrow and sighing shall flee away.
ISA|36|1|In the fourteenth year of King Hezekiah, Sennacherib king of Assyria came up against all the fortified cities of Judah and took them.
ISA|36|2|And the king of Assyria sent the Rabshakeh from Lachish to King Hezekiah at Jerusalem, with a great army. And he stood by the conduit of the upper pool on the highway to the Washer's Field.
ISA|36|3|And there came out to him Eliakim the son of Hilkiah, who was over the household, and Shebna the secretary, and Joah the son of Asaph, the recorder.
ISA|36|4|And the Rabshakeh said to them, "Say to Hezekiah, 'Thus says the great king, the king of Assyria: On what do you rest this trust of yours?
ISA|36|5|Do you think that mere words are strategy and power for war? In whom do you now trust, that you have rebelled against me?
ISA|36|6|Behold, you are trusting in Egypt, that broken reed of a staff, which will pierce the hand of any man who leans on it. Such is Pharaoh king of Egypt to all who trust in him.
ISA|36|7|But if you say to me, "We trust in the LORD our God," is it not he whose high places and altars Hezekiah has removed, saying to Judah and to Jerusalem, "You shall worship before this altar"?
ISA|36|8|Come now, make a wager with my master the king of Assyria: I will give you two thousand horses, if you are able on your part to set riders on them.
ISA|36|9|How then can you repulse a single captain among the least of my master's servants, when you trust in Egypt for chariots and for horsemen?
ISA|36|10|Moreover, is it without the LORD that I have come up against this land to destroy it? The LORD said to me, Go up against this land and destroy it.'"
ISA|36|11|Then Eliakim, Shebna, and Joah said to the Rabshakeh, "Please speak to your servants in Aramaic, for we understand it. Do not speak to us in the language of Judah within the hearing of the people who are on the wall."
ISA|36|12|But the Rabshakeh said, "Has my master sent me to speak these words to your master and to you, and not to the men sitting on the wall, who are doomed with you to eat their own dung and drink their own urine?"
ISA|36|13|Then the Rabshakeh stood and called out in a loud voice in the language of Judah: "Hear the words of the great king, the king of Assyria!
ISA|36|14|Thus says the king: 'Do not let Hezekiah deceive you, for he will not be able to deliver you.
ISA|36|15|Do not let Hezekiah make you trust in the LORD by saying, "The LORD will surely deliver us. This city will not be given into the hand of the king of Assyria."
ISA|36|16|Do not listen to Hezekiah. For thus says the king of Assyria: Make your peace with me and come out to me. Then each one of you will eat of his own vine, and each one of his own fig tree, and each one of you will drink the water of his own cistern,
ISA|36|17|until I come and take you away to a land like your own land, a land of grain and wine, a land of bread and vineyards.
ISA|36|18|Beware lest Hezekiah mislead you by saying, "The LORD will deliver us." Has any of the gods of the nations delivered his land out of the hand of the king of Assyria?
ISA|36|19|Where are the gods of Hamath and Arpad? Where are the gods of Sepharvaim? Have they delivered Samaria out of my hand?
ISA|36|20|Who among all the gods of these lands have delivered their lands out of my hand, that the LORD should deliver Jerusalem out of my hand?'"
ISA|36|21|But they were silent and answered him not a word, for the king's command was, "Do not answer him."
ISA|36|22|Then Eliakim the son of Hilkiah, who was over the household, and Shebna the secretary, and Joah the son of Asaph, the recorder, came to Hezekiah with their clothes torn, and told him the words of the Rabshakeh.
ISA|37|1|As soon as King Hezekiah heard it, he tore his clothes and covered himself with sackcloth and went into the house of the LORD.
ISA|37|2|And he sent Eliakim, who was over the household, and Shebna the secretary, and the senior priests, covered with sackcloth, to the prophet Isaiah the son of Amoz.
ISA|37|3|They said to him, "Thus says Hezekiah, 'This day is a day of distress, of rebuke, and of disgrace; children have come to the point of birth, and there is no strength to bring them forth.
ISA|37|4|It may be that the LORD your God will hear the words of the Rabshakeh, whom his master the king of Assyria has sent to mock the living God, and will rebuke the words that the LORD your God has heard; therefore lift up your prayer for the remnant that is left.'"
ISA|37|5|When the servants of King Hezekiah came to Isaiah,
ISA|37|6|Isaiah said to them, "Say to your master, 'Thus says the LORD: Do not be afraid because of the words that you have heard, with which the young men of the king of Assyria have reviled me.
ISA|37|7|Behold, I will put a spirit in him, so that he shall hear a rumor and return to his own land, and I will make him fall by the sword in his own land.'"
ISA|37|8|The Rabshakeh returned, and found the king of Assyria fighting against Libnah, for he had heard that the king had left Lachish.
ISA|37|9|Now the king heard concerning Tirhakah king of Cush, "He has set out to fight against you." And when he heard it, he sent messengers to Hezekiah, saying,
ISA|37|10|"Thus shall you speak to Hezekiah king of Judah: 'Do not let your God in whom you trust deceive you by promising that Jerusalem will not be given into the hand of the king of Assyria.
ISA|37|11|Behold, you have heard what the kings of Assyria have done to all lands, devoting them to destruction. And shall you be delivered?
ISA|37|12|Have the gods of the nations delivered them, the nations that my fathers destroyed, Gozan, Haran, Rezeph, and the people of Eden who were in Telassar?
ISA|37|13|Where is the king of Hamath, the king of Arpad, the king of the city of Sepharvaim, the king of Hena, or the king of Ivvah?'"
ISA|37|14|Hezekiah received the letter from the hand of the messengers, and read it; and Hezekiah went up to the house of the LORD, and spread it before the LORD.
ISA|37|15|And Hezekiah prayed to the LORD:
ISA|37|16|"O LORD of hosts, God of Israel, who is enthroned above the cherubim, you are the God, you alone, of all the kingdoms of the earth; you have made heaven and earth.
ISA|37|17|Incline your ear, O LORD, and hear; open your eyes, O LORD, and see; and hear all the words of Sennacherib, which he has sent to mock the living God.
ISA|37|18|Truly, O LORD, the kings of Assyria have laid waste all the nations and their lands,
ISA|37|19|and have cast their gods into the fire. For they were no gods, but the work of men's hands, wood and stone. Therefore they were destroyed.
ISA|37|20|So now, O LORD our God, save us from his hand, that all the kingdoms of the earth may know that you alone are the LORD."
ISA|37|21|Then Isaiah the son of Amoz sent to Hezekiah, saying, "Thus says the LORD, the God of Israel: Because you have prayed to me concerning Sennacherib king of Assyria,
ISA|37|22|this is the word that the LORD has spoken concerning him: "' She despises you, she scorns you- the virgin daughter of Zion; she wags her head behind you- the daughter of Jerusalem.
ISA|37|23|"'Whom have you mocked and reviled? Against whom have you raised your voice and lifted your eyes to the heights? Against the Holy One of Israel!
ISA|37|24|By your servants you have mocked the Lord, and you have said, With my many chariots I have gone up the heights of the mountains, to the far recesses of Lebanon, to cut down its tallest cedars, its choicest cypresses, to come to its remotest height, its most fruitful forest.
ISA|37|25|I dug wells and drank waters, to dry up with the sole of my foot all the streams of Egypt.
ISA|37|26|"'Have you not heard that I determined it long ago? I planned from days of old what now I bring to pass, that you should make fortified cities crash into heaps of ruins,
ISA|37|27|while their inhabitants, shorn of strength, are dismayed and confounded, and have become like plants of the field and like tender grass, like grass on the housetops, blighted before it is grown.
ISA|37|28|"'I know your sitting down and your going out and coming in, and your raging against me.
ISA|37|29|Because you have raged against me and your complacency has come to my ears, I will put my hook in your nose and my bit in your mouth, and I will turn you back on the way by which you came.'
ISA|37|30|"And this shall be the sign for you: this year you shall eat what grows of itself, and in the second year what springs from that. Then in the third year sow and reap, and plant vineyards, and eat their fruit.
ISA|37|31|And the surviving remnant of the house of Judah shall again take root downward and bear fruit upward.
ISA|37|32|For out of Jerusalem shall go a remnant, and out of Mount Zion a band of survivors. The zeal of the LORD of hosts will do this.
ISA|37|33|"Therefore thus says the LORD concerning the king of Assyria: He shall not come into this city or shoot an arrow there or come before it with a shield or cast up a siege mound against it.
ISA|37|34|By the way that he came, by the same he shall return, and he shall not come into this city, declares the LORD.
ISA|37|35|For I will defend this city to save it, for my own sake and for the sake of my servant David."
ISA|37|36|And the angel of the LORD went out and struck down a hundred and eighty-five thousand in the camp of the Assyrians. And when people arose early in the morning, behold, these were all dead bodies.
ISA|37|37|Then Sennacherib king of Assyria departed and returned home and lived at Nineveh.
ISA|37|38|And as he was worshiping in the house of Nisroch his god, Adrammelech and Sharezer, his sons, struck him down with the sword. And after they escaped into the land of Ararat, Esarhaddon his son reigned in his place.
ISA|38|1|In those days Hezekiah became sick and was at the point of death. And Isaiah the prophet the son of Amoz came to him, and said to him, "Thus says the LORD: Set your house in order, for you shall die, you shall not recover."
ISA|38|2|Then Hezekiah turned his face to the wall and prayed to the LORD,
ISA|38|3|and said, "Please, O LORD, remember how I have walked before you in faithfulness and with a whole heart, and have done what is good in your sight." And Hezekiah wept bitterly.
ISA|38|4|Then the word of the LORD came to Isaiah:
ISA|38|5|"Go and say to Hezekiah, Thus says the LORD, the God of David your father: I have heard your prayer; I have seen your tears. Behold, I will add fifteen years to your life.
ISA|38|6|I will deliver you and this city out of the hand of the king of Assyria, and will defend this city.
ISA|38|7|"This shall be the sign to you from the LORD, that the LORD will do this thing that he has promised:
ISA|38|8|Behold, I will make the shadow cast by the declining sun on the dial of Ahaz turn back ten steps." So the sun turned back on the dial the ten steps by which it had declined.
ISA|38|9|A writing of Hezekiah king of Judah, after he had been sick and had recovered from his sickness:
ISA|38|10|I said, In the middle of my days I must depart; I am consigned to the gates of Sheol for the rest of my years.
ISA|38|11|I said, I shall not see the LORD, the LORD in the land of the living; I shall look on man no more among the inhabitants of the world.
ISA|38|12|My dwelling is plucked up and removed from me like a shepherd's tent; like a weaver I have rolled up my life; he cuts me off from the loom; from day to night you bring me to an end;
ISA|38|13|I calmed myself until morning; like a lion he breaks all my bones; from day to night you bring me to an end.
ISA|38|14|Like a swallow or a crane I chirp; I moan like a dove. My eyes are weary with looking upward. O Lord, I am oppressed; be my pledge of safety!
ISA|38|15|What shall I say? For he has spoken to me, and he himself has done it. I walk slowly all my years because of the bitterness of my soul.
ISA|38|16|O Lord, by these things men live, and in all these is the life of my spirit. Oh restore me to health and make me live!
ISA|38|17|Behold, it was for my welfare that I had great bitterness; but in love you have delivered my life from the pit of destruction, for you have cast all my sins behind your back.
ISA|38|18|For Sheol does not thank you; death does not praise you; those who go down to the pit do not hope for your faithfulness.
ISA|38|19|The living, the living, he thanks you, as I do this day; the father makes known to the children your faithfulness.
ISA|38|20|The LORD will save me, and we will play my music on stringed instruments all the days of our lives, at the house of the LORD.
ISA|38|21|Now Isaiah had said, "Let them take a cake of figs and apply it to the boil, that he may recover."
ISA|38|22|Hezekiah also had said, "What is the sign that I shall go up to the house of the LORD?"
ISA|39|1|At that time Merodach-baladan the son of Baladan, king of Babylon, sent envoys with letters and a present to Hezekiah, for he heard that he had been sick and had recovered.
ISA|39|2|And Hezekiah welcomed them gladly. And he showed them his treasure house, the silver, the gold, the spices, the precious oil, his whole armory, all that was found in his storehouses. There was nothing in his house or in all his realm that Hezekiah did not show them.
ISA|39|3|Then Isaiah the prophet came to King Hezekiah, and said to him, "What did these men say? And from where did they come to you?" Hezekiah said, "They have come to me from a far country, from Babylon."
ISA|39|4|He said, "What have they seen in your house?" Hezekiah answered, "They have seen all that is in my house. There is nothing in my storehouses that I did not show them."
ISA|39|5|Then Isaiah said to Hezekiah, "Hear the word of the LORD of hosts:
ISA|39|6|Behold, the days are coming, when all that is in your house, and that which your fathers have stored up till this day, shall be carried to Babylon. Nothing shall be left, says the LORD.
ISA|39|7|And some of your own sons, who will come from you, whom you will father, shall be taken away, and they shall be eunuchs in the palace of the king of Babylon."
ISA|39|8|Then said Hezekiah to Isaiah, "The word of the LORD that you have spoken is good." For he thought, "There will be peace and security in my days."
ISA|40|1|Comfort, comfort my people, says your God.
ISA|40|2|Speak tenderly to Jerusalem, and cry to her that her warfare is ended, that her iniquity is pardoned, that she has received from the LORD's hand double for all her sins.
ISA|40|3|A voice cries: "In the wilderness prepare the way of the LORD; make straight in the desert a highway for our God.
ISA|40|4|Every valley shall be lifted up, and every mountain and hill be made low; the uneven ground shall become level, and the rough places a plain.
ISA|40|5|And the glory of the LORD shall be revealed, and all flesh shall see it together, for the mouth of the LORD has spoken."
ISA|40|6|A voice says, "Cry!" And I said, "What shall I cry?" All flesh is grass, and all its beauty is like the flower of the field.
ISA|40|7|The grass withers, the flower fades when the breath of the LORD blows on it; surely the people are grass.
ISA|40|8|The grass withers, the flower fades, but the word of our God will stand forever.
ISA|40|9|Get you up to a high mountain, O Zion, herald of good news; lift up your voice with strength, O Jerusalem, herald of good news; lift it up, fear not; say to the cities of Judah, "Behold your God!"
ISA|40|10|Behold, the Lord GOD comes with might, and his arm rules for him; behold, his reward is with him, and his recompense before him.
ISA|40|11|He will tend his flock like a shepherd; he will gather the lambs in his arms; he will carry them in his bosom, and gently lead those that are with young.
ISA|40|12|Who has measured the waters in the hollow of his hand and marked off the heavens with a span, enclosed the dust of the earth in a measure and weighed the mountains in scales and the hills in a balance?
ISA|40|13|Who has measured the Spirit of the LORD, or what man shows him his counsel?
ISA|40|14|Whom did he consult, and who made him understand? Who taught him the path of justice, and taught him knowledge, and showed him the way of understanding?
ISA|40|15|Behold, the nations are like a drop from a bucket, and are accounted as the dust on the scales; behold, he takes up the coastlands like fine dust.
ISA|40|16|Lebanon would not suffice for fuel, nor are its beasts enough for a burnt offering.
ISA|40|17|All the nations are as nothing before him, they are accounted by him as less than nothing and emptiness.
ISA|40|18|To whom then will you liken God, or what likeness compare with him?
ISA|40|19|An idol! A craftsman casts it, and a goldsmith overlays it with gold and casts for it silver chains.
ISA|40|20|He who is too impoverished for an offering chooses wood that will not rot; he seeks out a skillful craftsman to set up an idol that will not move.
ISA|40|21|Do you not know? Do you not hear? Has it not been told you from the beginning? Have you not understood from the foundations of the earth?
ISA|40|22|It is he who sits above the circle of the earth, and its inhabitants are like grasshoppers; who stretches out the heavens like a curtain, and spreads them like a tent to dwell in;
ISA|40|23|who brings princes to nothing, and makes the rulers of the earth as emptiness.
ISA|40|24|Scarcely are they planted, scarcely sown, scarcely has their stem taken root in the earth, when he blows on them, and they wither, and the tempest carries them off like stubble.
ISA|40|25|To whom then will you compare me, that I should be like him? says the Holy One.
ISA|40|26|Lift up your eyes on high and see: who created these? He who brings out their host by number, calling them all by name, by the greatness of his might, and because he is strong in power not one is missing.
ISA|40|27|Why do you say, O Jacob, and speak, O Israel, "My way is hidden from the LORD, and my right is disregarded by my God"?
ISA|40|28|Have you not known? Have you not heard? The LORD is the everlasting God, the Creator of the ends of the earth. He does not faint or grow weary; his understanding is unsearchable.
ISA|40|29|He gives power to the faint, and to him who has no might he increases strength.
ISA|40|30|Even youths shall faint and be weary, and young men shall fall exhausted;
ISA|40|31|but they who wait for the LORD shall renew their strength; they shall mount up with wings like eagles; they shall run and not be weary; they shall walk and not faint.
ISA|41|1|Listen to me in silence, O coastlands; let the peoples renew their strength; let them approach, then let them speak; let us together draw near for judgment.
ISA|41|2|Who stirred up one from the east whom victory meets at every step? He gives up nations before him, so that he tramples kings underfoot; he makes them like dust with his sword, like driven stubble with his bow.
ISA|41|3|He pursues them and passes on safely, by paths his feet have not trod.
ISA|41|4|Who has performed and done this, calling the generations from the beginning? I, the LORD, the first, and with the last; I am he.
ISA|41|5|The coastlands have seen and are afraid; the ends of the earth tremble; they have drawn near and come.
ISA|41|6|Everyone helps his neighbor and says to his brother, "Be strong!"
ISA|41|7|The craftsman strengthens the goldsmith, and he who smooths with the hammer him who strikes the anvil, saying of the soldering, "It is good"; and they strengthen it with nails so that it cannot be moved.
ISA|41|8|But you, Israel, my servant, Jacob, whom I have chosen, the offspring of Abraham, my friend;
ISA|41|9|you whom I took from the ends of the earth, and called from its farthest corners, saying to you, "You are my servant, I have chosen you and not cast you off";
ISA|41|10|fear not, for I am with you; be not dismayed, for I am your God; I will strengthen you, I will help you, I will uphold you with my righteous right hand.
ISA|41|11|Behold, all who are incensed against you shall be put to shame and confounded; those who strive against you shall be as nothing and shall perish.
ISA|41|12|You shall seek those who contend with you, but you shall not find them; those who war against you shall be as nothing at all.
ISA|41|13|For I, the LORD your God, hold your right hand; it is I who say to you, "Fear not, I am the one who helps you."
ISA|41|14|Fear not, you worm Jacob, you men of Israel! I am the one who helps you, declares the LORD; your Redeemer is the Holy One of Israel.
ISA|41|15|Behold, I make of you a threshing sledge, new, sharp, and having teeth; you shall thresh the mountains and crush them, and you shall make the hills like chaff;
ISA|41|16|you shall winnow them, and the wind shall carry them away, and the tempest shall scatter them. And you shall rejoice in the LORD; in the Holy One of Israel you shall glory.
ISA|41|17|When the poor and needy seek water, and there is none, and their tongue is parched with thirst, I the LORD will answer them; I the God of Israel will not forsake them.
ISA|41|18|I will open rivers on the bare heights, and fountains in the midst of the valleys. I will make the wilderness a pool of water, and the dry land springs of water.
ISA|41|19|I will put in the wilderness the cedar, the acacia, the myrtle, and the olive. I will set in the desert the cypress, the plane and the pine together,
ISA|41|20|that men may see and know, may consider and understand together, that the hand of the LORD has done this, the Holy One of Israel has created it.
ISA|41|21|Set forth your case, says the LORD; bring your proofs, says the King of Jacob.
ISA|41|22|Let them bring them, and tell us what is to happen. Tell us the former things, what they are, that we may consider them, that we may know their outcome; or declare to us the things to come.
ISA|41|23|Tell us what is to come hereafter, that we may know that you are gods; do good, or do harm, that we may be dismayed and terrified.
ISA|41|24|Behold, you are nothing, and your work is less than nothing; an abomination is he who chooses you.
ISA|41|25|I stirred up one from the north, and he has come, from the rising of the sun, and he shall call upon my name; he shall trample on rulers as on mortar, as the potter treads clay.
ISA|41|26|Who declared it from the beginning, that we might know, and beforehand, that we might say, "He is right"? There was none who declared it, none who proclaimed, none who heard your words.
ISA|41|27|I was the first to say to Zion, "Behold, here they are!" and I give to Jerusalem a herald of good news.
ISA|41|28|But when I look there is no one; among these there is no counselor who, when I ask, gives an answer.
ISA|41|29|Behold, they are all a delusion; their works are nothing; their metal images are empty wind.
ISA|42|1|Behold my servant, whom I uphold, my chosen, in whom my soul delights; I have put my Spirit upon him; he will bring forth justice to the nations.
ISA|42|2|He will not cry aloud or lift up his voice, or make it heard in the street;
ISA|42|3|a bruised reed he will not break, and a faintly burning wick he will not quench; he will faithfully bring forth justice.
ISA|42|4|He will not grow faint or be discouraged till he has established justice in the earth; and the coastlands wait for his law.
ISA|42|5|Thus says God, the LORD, who created the heavens and stretched them out, who spread out the earth and what comes from it, who gives breath to the people on it and spirit to those who walk in it:
ISA|42|6|"I am the LORD; I have called you in righteousness; I will take you by the hand and keep you; I will give you as a covenant for the people, a light for the nations,
ISA|42|7|to open the eyes that are blind, to bring out the prisoners from the dungeon, from the prison those who sit in darkness.
ISA|42|8|I am the LORD; that is my name; my glory I give to no other, nor my praise to carved idols.
ISA|42|9|Behold, the former things have come to pass, and new things I now declare; before they spring forth I tell you of them."
ISA|42|10|Sing to the LORD a new song, his praise from the end of the earth, you who go down to the sea, and all that fills it, the coastlands and their inhabitants.
ISA|42|11|Let the desert and its cities lift up their voice, the villages that Kedar inhabits; let the habitants of Sela sing for joy, let them shout from the top of the mountains.
ISA|42|12|Let them give glory to the LORD, and declare his praise in the coastlands.
ISA|42|13|The LORD goes out like a mighty man, like a man of war he stirs up his zeal; he cries out, he shouts aloud, he shows himself mighty against his foes.
ISA|42|14|For a long time I have held my peace; I have kept still and restrained myself; now I will cry out like a woman in labor; I will gasp and pant.
ISA|42|15|I will lay waste mountains and hills, and dry up all their vegetation; I will turn the rivers into islands, and dry up the pools.
ISA|42|16|And I will lead the blind in a way that they do not know, in paths that they have not known I will guide them. I will turn the darkness before them into light, the rough places into level ground. These are the things I do, and I do not forsake them.
ISA|42|17|They are turned back and utterly put to shame, who trust in carved idols, who say to metal images, "You are our gods."
ISA|42|18|Hear, you deaf, and look, you blind, that you may see!
ISA|42|19|Who is blind but my servant, or deaf as my messenger whom I send? Who is blind as my dedicated one, or blind as the servant of the LORD?
ISA|42|20|He sees many things, but does not observe them; his ears are open, but he does not hear.
ISA|42|21|The LORD was pleased, for his righteousness' sake, to magnify his law and make it glorious.
ISA|42|22|But this is a people plundered and looted; they are all of them trapped in holes and hidden in prisons; they have become plunder with none to rescue, spoil with none to say, "Restore!"
ISA|42|23|Who among you will give ear to this, will attend and listen for the time to come?
ISA|42|24|Who gave up Jacob to the looter, and Israel to the plunderers? Was it not the LORD, against whom we have sinned, in whose ways they would not walk, and whose law they would not obey?
ISA|42|25|So he poured on him the heat of his anger and the might of battle; it set him on fire all around, but he did not understand; it burned him up, but he did not take it to heart.
ISA|43|1|But now thus says the LORD, he who created you, O Jacob, he who formed you, O Israel: "Fear not, for I have redeemed you; I have called you by name, you are mine.
ISA|43|2|When you pass through the waters, I will be with you; and through the rivers, they shall not overwhelm you; when you walk through fire you shall not be burned, and the flame shall not consume you.
ISA|43|3|For I am the LORD your God, the Holy One of Israel, your Savior. I give Egypt as your ransom, Cush and Seba in exchange for you.
ISA|43|4|Because you are precious in my eyes, and honored, and I love you, I give men in return for you, peoples in exchange for your life.
ISA|43|5|Fear not, for I am with you; I will bring your offspring from the east, and from the west I will gather you.
ISA|43|6|I will say to the north, Give up, and to the south, Do not withhold; bring my sons from afar and my daughters from the end of the earth,
ISA|43|7|everyone who is called by my name, whom I created for my glory, whom I formed and made."
ISA|43|8|Bring out the people who are blind, yet have eyes, who are deaf, yet have ears!
ISA|43|9|All the nations gather together, and the peoples assemble. Who among them can declare this, and show us the former things? Let them bring their witnesses to prove them right, and let them hear and say, It is true.
ISA|43|10|"You are my witnesses," declares the LORD, "and my servant whom I have chosen, that you may know and believe me and understand that I am he. Before me no god was formed, nor shall there be any after me.
ISA|43|11|I, I am the LORD, and besides me there is no savior.
ISA|43|12|I declared and saved and proclaimed, when there was no strange god among you; and you are my witnesses," declares the LORD, "and I am God.
ISA|43|13|Also henceforth I am he; there is none who can deliver from my hand; I work, and who can turn it back?"
ISA|43|14|Thus says the LORD, your Redeemer, the Holy One of Israel: "For your sake I send to Babylon and bring them all down as fugitives, even the Chaldeans, in the ships in which they rejoice.
ISA|43|15|I am the LORD, your Holy One, the Creator of Israel, your King."
ISA|43|16|Thus says the LORD, who makes a way in the sea, a path in the mighty waters,
ISA|43|17|who brings forth chariot and horse, army and warrior; they lie down, they cannot rise, they are extinguished, quenched like a wick:
ISA|43|18|"Remember not the former things, nor consider the things of old.
ISA|43|19|Behold, I am doing a new thing; now it springs forth, do you not perceive it? I will make a way in the wilderness and rivers in the desert.
ISA|43|20|The wild beasts will honor me, the jackals and the ostriches, for I give water in the wilderness, rivers in the desert, to give drink to my chosen people,
ISA|43|21|the people whom I formed for myself that they might declare my praise.
ISA|43|22|"Yet you did not call upon me, O Jacob; but you have been weary of me, O Israel!
ISA|43|23|You have not brought me your sheep for burnt offerings, or honored me with your sacrifices. I have not burdened you with offerings, or wearied you with frankincense.
ISA|43|24|You have not bought me sweet cane with money, or satisfied me with the fat of your sacrifices. But you have burdened me with your sins; you have wearied me with your iniquities.
ISA|43|25|"I, I am he who blots out your transgressions for my own sake, and I will not remember your sins.
ISA|43|26|Put me in remembrance; let us argue together; set forth your case, that you may be proved right.
ISA|43|27|Your first father sinned, and your mediators transgressed against me.
ISA|43|28|Therefore I will profane the princes of the sanctuary, and deliver Jacob to utter destruction and Israel to reviling.
ISA|44|1|"But now hear, O Jacob my servant, Israel whom I have chosen!
ISA|44|2|Thus says the LORD who made you, who formed you from the womb and will help you: Fear not, O Jacob my servant, Jeshurun whom I have chosen.
ISA|44|3|For I will pour water on the thirsty land, and streams on the dry ground; I will pour my Spirit upon your offspring, and my blessing on your descendants.
ISA|44|4|They shall spring up among the grass like willows by flowing streams.
ISA|44|5|This one will say, 'I am the LORD's,' another will call on the name of Jacob, and another will write on his hand, 'The LORD's,' and name himself by the name of Israel."
ISA|44|6|Thus says the LORD, the King of Israel and his Redeemer, the LORD of hosts: "I am the first and I am the last; besides me there is no god.
ISA|44|7|Who is like me? Let him proclaim it. Let him declare and set it before me, since I appointed an ancient people. Let them declare what is to come, and what will happen.
ISA|44|8|Fear not, nor be afraid; have I not told you from of old and declared it? And you are my witnesses! Is there a God besides me? There is no Rock; I know not any."
ISA|44|9|All who fashion idols are nothing, and the things they delight in do not profit. Their witnesses neither see nor know, that they may be put to shame.
ISA|44|10|Who fashions a god or casts an idol that is profitable for nothing?
ISA|44|11|Behold, all his companions shall be put to shame, and the craftsmen are only human. Let them all assemble, let them stand forth. They shall be terrified; they shall be put to shame together.
ISA|44|12|The ironsmith takes a cutting tool and works it over the coals. He fashions it with hammers and works it with his strong arm. He becomes hungry, and his strength fails; he drinks no water and is faint.
ISA|44|13|The carpenter stretches a line; he marks it out with a pencil. He shapes it with planes and marks it with a compass. He shapes it into the figure of a man, with the beauty of a man, to dwell in a house.
ISA|44|14|He cuts down cedars, or he chooses a cypress tree or an oak and lets it grow strong among the trees of the forest. He plants a cedar and the rain nourishes it.
ISA|44|15|Then it becomes fuel for a man. He takes a part of it and warms himself; he kindles a fire and bakes bread. Also he makes a god and worships it; he makes it an idol and falls down before it.
ISA|44|16|Half of it he burns in the fire. Over the half he eats meat; he roasts it and is satisfied. Also he warms himself and says, "Aha, I am warm, I have seen the fire!"
ISA|44|17|And the rest of it he makes into a god, his idol, and falls down to it and worships it. He prays to it and says, "Deliver me, for you are my god!"
ISA|44|18|They know not, nor do they discern, for he has shut their eyes, so that they cannot see, and their hearts, so that they cannot understand.
ISA|44|19|No one considers, nor is there knowledge or discernment to say, "Half of it I burned in the fire; I also baked bread on its coals; I roasted meat and have eaten. And shall I make the rest of it an abomination? Shall I fall down before a block of wood?"
ISA|44|20|He feeds on ashes; a deluded heart has led him astray, and he cannot deliver himself or say, "Is there not a lie in my right hand?"
ISA|44|21|Remember these things, O Jacob, and Israel, for you are my servant; I formed you; you are my servant; O Israel, you will not be forgotten by me.
ISA|44|22|I have blotted out your transgressions like a cloud and your sins like mist; return to me, for I have redeemed you.
ISA|44|23|Sing, O heavens, for the LORD has done it; shout, O depths of the earth; break forth into singing, O mountains, O forest, and every tree in it! For the LORD has redeemed Jacob, and will be glorified in Israel.
ISA|44|24|Thus says the LORD, your Redeemer, who formed you from the womb: "I am the LORD, who made all things, who alone stretched out the heavens, who spread out the earth by myself,
ISA|44|25|who frustrates the signs of liars and makes fools of diviners, who turns wise men back and makes their knowledge foolish,
ISA|44|26|who confirms the word of his servant and fulfills the counsel of his messengers, who says of Jerusalem, 'She shall be inhabited,' and of the cities of Judah, 'They shall be built, and I will raise up their ruins';
ISA|44|27|who says to the deep, 'Be dry; I will dry up your rivers';
ISA|44|28|who says of Cyrus, 'He is my shepherd, and he shall fulfill all my purpose'; saying of Jerusalem, 'She shall be built,' and of the temple, 'Your foundation shall be laid.'"
ISA|45|1|Thus says the LORD to his anointed, to Cyrus, whose right hand I have grasped, to subdue nations before him and to loose the belts of kings, to open doors before him that gates may not be closed:
ISA|45|2|"I will go before you and level the exalted places, I will break in pieces the doors of bronze and cut through the bars of iron,
ISA|45|3|I will give you the treasures of darkness and the hoards in secret places, that you may know that it is I, the LORD, the God of Israel, who call you by your name.
ISA|45|4|For the sake of my servant Jacob, and Israel my chosen, I call you by your name, I name you, though you do not know me.
ISA|45|5|I am the LORD, and there is no other, besides me there is no God; I equip you, though you do not know me,
ISA|45|6|that people may know, from the rising of the sun and from the west, that there is none besides me; I am the LORD, and there is no other.
ISA|45|7|I form light and create darkness, I make well-being and create calamity, I am the LORD, who does all these things.
ISA|45|8|"Shower, O heavens, from above, and let the clouds rain down righteousness; let the earth open, that salvation and righteousness may bear fruit; let the earth cause them both to sprout; I the LORD have created it.
ISA|45|9|"Woe to him who strives with him who formed him, a pot among earthen pots! Does the clay say to him who forms it, 'What are you making?' or 'Your work has no handles'?
ISA|45|10|Woe to him who says to a father, 'What are you begetting?' or to a woman, 'With what are you in labor?'"
ISA|45|11|Thus says the LORD, the Holy One of Israel, and the one who formed him: "Ask me of things to come; will you command me concerning my children and the work of my hands?
ISA|45|12|I made the earth and created man on it; it was my hands that stretched out the heavens, and I commanded all their host.
ISA|45|13|I have stirred him up in righteousness, and I will make all his ways level; he shall build my city and set my exiles free, not for price or reward," says the LORD of hosts.
ISA|45|14|Thus says the LORD: "The wealth of Egypt and the merchandise of Cush, and the Sabeans, men of stature, shall come over to you and be yours; they shall follow you; they shall come over in chains and bow down to you. They will plead with you, saying: 'Surely God is in you, and there is no other, no god besides him.'"
ISA|45|15|Truly, you are a God who hides yourself, O God of Israel, the Savior.
ISA|45|16|All of them are put to shame and confounded; the makers of idols go in confusion together.
ISA|45|17|But Israel is saved by the LORD with everlasting salvation; you shall not be put to shame or confounded to all eternity.
ISA|45|18|For thus says the LORD, who created the heavens (he is God!), who formed the earth and made it (he established it; he did not create it empty, he formed it to be inhabited!): "I am the LORD, and there is no other.
ISA|45|19|I did not speak in secret, in a land of darkness; I did not say to the offspring of Jacob, 'Seek me in vain.' I the LORD speak the truth; I declare what is right.
ISA|45|20|"Assemble yourselves and come; draw near together, you survivors of the nations! They have no knowledge who carry about their wooden idols, and keep on praying to a god that cannot save.
ISA|45|21|Declare and present your case; let them take counsel together! Who told this long ago? Who declared it of old? Was it not I, the LORD? And there is no other god besides me, a righteous God and a Savior; there is none besides me.
ISA|45|22|"Turn to me and be saved, all the ends of the earth! For I am God, and there is no other.
ISA|45|23|By myself I have sworn; from my mouth has gone out in righteousness a word that shall not return: 'To me every knee shall bow, every tongue shall swear allegiance.'
ISA|45|24|"Only in the LORD, it shall be said of me, are righteousness and strength; to him shall come and be ashamed all who were incensed against him.
ISA|45|25|In the LORD all the offspring of Israel shall be justified and shall glory."
ISA|46|1|Bel bows down; Nebo stoops; their idols are on beasts and livestock; these things you carry are borne as burdens on weary beasts.
ISA|46|2|They stoop; they bow down together; they cannot save the burden, but themselves go into captivity.
ISA|46|3|"Listen to me, O house of Jacob, all the remnant of the house of Israel, who have been borne by me from before your birth, carried from the womb;
ISA|46|4|even to your old age I am he, and to gray hairs I will carry you. I have made, and I will bear; I will carry and will save.
ISA|46|5|"To whom will you liken me and make me equal, and compare me, that we may be alike?
ISA|46|6|Those who lavish gold from the purse, and weigh out silver in the scales, hire a goldsmith, and he makes it into a god; then they fall down and worship!
ISA|46|7|They lift it to their shoulders, they carry it, they set it in its place, and it stands there; it cannot move from its place. If one cries to it, it does not answer or save him from his trouble.
ISA|46|8|"Remember this and stand firm, recall it to mind, you transgressors,
ISA|46|9|remember the former things of old; for I am God, and there is no other; I am God, and there is none like me,
ISA|46|10|declaring the end from the beginning and from ancient times things not yet done, saying, 'My counsel shall stand, and I will accomplish all my purpose,'
ISA|46|11|calling a bird of prey from the east, the man of my counsel from a far country. I have spoken, and I will bring it to pass; I have purposed, and I will do it.
ISA|46|12|"Listen to me, you stubborn of heart, you who are far from righteousness:
ISA|46|13|I bring near my righteousness; it is not far off, and my salvation will not delay; I will put salvation in Zion, for Israel my glory."
ISA|47|1|Come down and sit in the dust, O virgin daughter of Babylon; sit on the ground without a throne, O daughter of the Chaldeans! For you shall no more be called tender and delicate.
ISA|47|2|Take the millstones and grind flour, put off your veil, strip off your robe, uncover your legs, pass through the rivers.
ISA|47|3|Your nakedness shall be uncovered, and your disgrace shall be seen. I will take vengeance, and I will spare no one.
ISA|47|4|Our Redeemer- the LORD of hosts is his name- is the Holy One of Israel.
ISA|47|5|Sit in silence, and go into darkness, O daughter of the Chaldeans; for you shall no more be called the mistress of kingdoms.
ISA|47|6|I was angry with my people; I profaned my heritage; I gave them into your hand; you showed them no mercy; on the aged you made your yoke exceedingly heavy.
ISA|47|7|You said, "I shall be mistress forever," so that you did not lay these things to heart or remember their end.
ISA|47|8|Now therefore hear this, you lover of pleasures, who sit securely, who say in your heart, "I am, and there is no one besides me; I shall not sit as a widow or know the loss of children":
ISA|47|9|These two things shall come to you in a moment, in one day; the loss of children and widowhood shall come upon you in full measure, in spite of your many sorceries and the great power of your enchantments.
ISA|47|10|You felt secure in your wickedness, you said, "No one sees me"; your wisdom and your knowledge led you astray, and you said in your heart, "I am, and there is no one besides me."
ISA|47|11|But evil shall come upon you, which you will not know how to charm away; disaster shall fall upon you, for which you will not be able to atone; and ruin shall come upon you suddenly, of which you know nothing.
ISA|47|12|Stand fast in your enchantments and your many sorceries, with which you have labored from your youth; perhaps you may be able to succeed; perhaps you may inspire terror.
ISA|47|13|You are wearied with your many counsels; let them stand forth and save you, those who divide the heavens, who gaze at the stars, who at the new moons make known what shall come upon you.
ISA|47|14|Behold, they are like stubble; the fire consumes them; they cannot deliver themselves from the power of the flame. No coal for warming oneself is this, no fire to sit before!
ISA|47|15|Such to you are those with whom you have labored, who have done business with you from your youth; they wander about each in his own direction; there is no one to save you.
ISA|48|1|Hear this, O house of Jacob, who are called by the name of Israel, and who came from the waters of Judah, who swear by the name of the LORD and confess the God of Israel, but not in truth or right.
ISA|48|2|For they call themselves after the holy city, and stay themselves on the God of Israel; the LORD of hosts is his name.
ISA|48|3|"The former things I declared of old; they went out from my mouth and I announced them; then suddenly I did them and they came to pass.
ISA|48|4|Because I know that you are obstinate, and your neck is an iron sinew and your forehead brass,
ISA|48|5|I declared them to you from of old, before they came to pass I announced them to you, lest you should say, 'My idol did them, my carved image and my metal image commanded them.'
ISA|48|6|"You have heard; now see all this; and will you not declare it? From this time forth I announce to you new things, hidden things that you have not known.
ISA|48|7|They are created now, not long ago; before today you have never heard of them, lest you should say, 'Behold, I knew them.'
ISA|48|8|You have never heard, you have never known, from of old your ear has not been opened. For I knew that you would surely deal treacherously, and that from before birth you were called a rebel.
ISA|48|9|"For my name's sake I defer my anger, for the sake of my praise I restrain it for you, that I may not cut you off.
ISA|48|10|Behold, I have refined you, but not as silver; I have tried you in the furnace of affliction.
ISA|48|11|For my own sake, for my own sake, I do it, for how should my name be profaned? My glory I will not give to another.
ISA|48|12|"Listen to me, O Jacob, and Israel, whom I called! I am he; I am the first, and I am the last.
ISA|48|13|My hand laid the foundation of the earth, and my right hand spread out the heavens; when I call to them, they stand forth together.
ISA|48|14|"Assemble, all of you, and listen! who among them has declared these things? The LORD loves him; he shall perform his purpose on Babylon, and his arm shall be against the Chaldeans.
ISA|48|15|I, even I, have spoken and called him; I have brought him, and he will prosper in his way.
ISA|48|16|Draw near to me, hear this: from the beginning I have not spoken in secret, from the time it came to be I have been there." And now the Lord GOD has sent me, and his Spirit.
ISA|48|17|Thus says the LORD, your Redeemer, the Holy One of Israel: "I am the LORD your God, who teaches you to profit, who leads you in the way you should go.
ISA|48|18|Oh that you had paid attention to my commandments! Then your peace would have been like a river, and your righteousness like the waves of the sea;
ISA|48|19|your offspring would have been like the sand, and your descendants like its grains; their name would never be cut off or destroyed from before me."
ISA|48|20|Go out from Babylon, flee from Chaldea, declare this with a shout of joy, proclaim it, send it out to the end of the earth; say, "The LORD has redeemed his servant Jacob!"
ISA|48|21|They did not thirst when he led them through the deserts; he made water flow for them from the rock; he split the rock and the water gushed out.
ISA|48|22|"There is no peace," says the LORD, "for the wicked."
ISA|49|1|Listen to me, O coastlands, and give attention, you peoples from afar. The LORD called me from the womb, from the body of my mother he named my name.
ISA|49|2|He made my mouth like a sharp sword; in the shadow of his hand he hid me; he made me a polished arrow; in his quiver he hid me away.
ISA|49|3|And he said to me, "You are my servant, Israel, in whom I will be glorified."
ISA|49|4|But I said, "I have labored in vain; I have spent my strength for nothing and vanity; yet surely my right is with the LORD, and my recompense with my God."
ISA|49|5|And now the LORD says, he who formed me from the womb to be his servant, to bring Jacob back to him; and that Israel might be gathered to him- for I am honored in the eyes of the LORD, and my God has become my strength-
ISA|49|6|he says: "It is too light a thing that you should be my servant to raise up the tribes of Jacob and to bring back the preserved of Israel; I will make you as a light for the nations, that my salvation may reach to the end of the earth."
ISA|49|7|Thus says the LORD, the Redeemer of Israel and his Holy One, to one deeply despised, abhorred by the nation, the servant of rulers: "Kings shall see and arise; princes, and they shall prostrate themselves; because of the LORD, who is faithful, the Holy One of Israel, who has chosen you."
ISA|49|8|Thus says the LORD: "In a time of favor I have answered you; in a day of salvation I have helped you; I will keep you and give you as a covenant to the people, to establish the land, to apportion the desolate heritages,
ISA|49|9|saying to the prisoners, 'Come out,' to those who are in darkness, 'Appear.' They shall feed along the ways; on all bare heights shall be their pasture;
ISA|49|10|they shall not hunger or thirst, neither scorching wind nor sun shall strike them, for he who has pity on them will lead them, and by springs of water will guide them.
ISA|49|11|And I will make all my mountains a road, and my highways shall be raised up.
ISA|49|12|Behold, these shall come from afar, and behold, these from the north and from the west, and these from the land of Syene."
ISA|49|13|Sing for joy, O heavens, and exult, O earth; break forth, O mountains, into singing! for the LORD has comforted his people and will have compassion on his afflicted.
ISA|49|14|But Zion said, "The LORD has forsaken me; my Lord has forgotten me."
ISA|49|15|"Can a woman forget her nursing child, that she should have no compassion on the son of her womb? Even these may forget, yet I will not forget you.
ISA|49|16|Behold, I have engraved you on the palms of my hands; your walls are continually before me.
ISA|49|17|Your builders make haste; your destroyers and those who laid you waste go out from you.
ISA|49|18|Lift up your eyes around and see; they all gather, they come to you. As I live, declares the LORD, you shall put them all on as an ornament; you shall bind them on as a bride does.
ISA|49|19|"Surely your waste and your desolate places and your devastated land- surely now you will be too narrow for your inhabitants, and those who swallowed you up will be far away.
ISA|49|20|The children of your bereavement will yet say in your ears: 'The place is too narrow for me; make room for me to dwell in.'
ISA|49|21|Then you will say in your heart: 'Who has borne me these? I was bereaved and barren, exiled and put away, but who has brought up these? Behold, I was left alone; from where have these come?'"
ISA|49|22|Thus says the Lord GOD: "Behold, I will lift up my hand to the nations, and raise my signal to the peoples; and they shall bring your sons in their bosom, and your daughters shall be carried on their shoulders.
ISA|49|23|Kings shall be your foster fathers, and their queens your nursing mothers. With their faces to the ground they shall bow down to you, and lick the dust of your feet. Then you will know that I am the LORD; those who wait for me shall not be put to shame."
ISA|49|24|Can the prey be taken from the mighty, or the captives of a tyrant be rescued?
ISA|49|25|For thus says the LORD: "Even the captives of the mighty shall be taken, and the prey of the tyrant be rescued, for I will contend with those who contend with you, and I will save your children.
ISA|49|26|I will make your oppressors eat their own flesh, and they shall be drunk with their own blood as with wine. Then all flesh shall know that I am the LORD your Savior, and your Redeemer, the Mighty One of Jacob."
ISA|50|1|Thus says the LORD:"Where is your mother's certificate of divorce, with which I sent her away? Or which of my creditors is it to whom I have sold you? Behold, for your iniquities you were sold, and for your transgressions your mother was sent away.
ISA|50|2|Why, when I came, was there no man; why, when I called, was there no one to answer? Is my hand shortened, that it cannot redeem? Or have I no power to deliver? Behold, by my rebuke I dry up the sea, I make the rivers a desert; their fish stink for lack of water and die of thirst.
ISA|50|3|I clothe the heavens with blackness and make sackcloth their covering."
ISA|50|4|The Lord GOD has given me the tongue of those who are taught, that I may know how to sustain with a word him who is weary. Morning by morning he awakens; he awakens my ear to hear as those who are taught.
ISA|50|5|The Lord GOD has opened my ear, and I was not rebellious; I turned not backward.
ISA|50|6|I gave my back to those who strike, and my cheeks to those who pull out the beard; I hid not my face from disgrace and spitting.
ISA|50|7|But the Lord GOD helps me; therefore I have not been disgraced; therefore I have set my face like a flint, and I know that I shall not be put to shame.
ISA|50|8|He who vindicates me is near. Who will contend with me? Let us stand up together. Who is my adversary? Let him come near to me.
ISA|50|9|Behold, the Lord GOD helps me; who will declare me guilty? Behold, all of them will wear out like a garment; the moth will eat them up.
ISA|50|10|Who among you fears the LORD and obeys the voice of his servant? Let him who walks in darkness and has no light trust in the name of the LORD and rely on his God.
ISA|50|11|Behold, all you who kindle a fire, who equip yourselves with burning torches! Walk by the light of your fire, and by the torches that you have kindled! This you have from my hand: you shall lie down in torment.
ISA|51|1|"Listen to me, you who pursue righteousness, you who seek the LORD: look to the rock from which you were hewn, and to the quarry from which you were dug.
ISA|51|2|Look to Abraham your father and to Sarah who bore you; for he was but one when I called him, that I might bless him and multiply him.
ISA|51|3|For the LORD comforts Zion; he comforts all her waste places and makes her wilderness like Eden, her desert like the garden of the LORD; joy and gladness will be found in her, thanksgiving and the voice of song.
ISA|51|4|"Give attention to me, my people, and give ear to me, my nation; for a law will go out from me, and I will set my justice for a light to the peoples.
ISA|51|5|My righteousness draws near, my salvation has gone out, and my arms will judge the peoples; the coastlands hope for me, and for my arm they wait.
ISA|51|6|Lift up your eyes to the heavens, and look at the earth beneath; for the heavens vanish like smoke, the earth will wear out like a garment, and they who dwell in it will die in like manner; but my salvation will be forever, and my righteousness will never be dismayed.
ISA|51|7|"Listen to me, you who know righteousness, the people in whose heart is my law; fear not the reproach of man, nor be dismayed at their revilings.
ISA|51|8|For the moth will eat them up like a garment, and the worm will eat them like wool; but my righteousness will be forever, and my salvation to all generations."
ISA|51|9|Awake, awake, put on strength, O arm of the LORD; awake, as in days of old, the generations of long ago. Was it not you who cut Rahab in pieces, that pierced the dragon?
ISA|51|10|Was it not you who dried up the sea, the waters of the great deep, who made the depths of the sea a way for the redeemed to pass over?
ISA|51|11|And the ransomed of the LORD shall return and come to Zion with singing; everlasting joy shall be upon their heads; they shall obtain gladness and joy, and sorrow and sighing shall flee away.
ISA|51|12|"I, I am he who comforts you; who are you that you are afraid of man who dies, of the son of man who is made like grass,
ISA|51|13|and have forgotten the LORD, your Maker, who stretched out the heavens and laid the foundations of the earth, and you fear continually all the day because of the wrath of the oppressor, when he sets himself to destroy? And where is the wrath of the oppressor?
ISA|51|14|He who is bowed down shall speedily be released; he shall not die and go down to the pit, neither shall his bread be lacking.
ISA|51|15|I am the LORD your God, who stirs up the sea so that its waves roar- the LORD of hosts is his name.
ISA|51|16|And I have put my words in your mouth and covered you in the shadow of my hand, establishing the heavens and laying the foundations of the earth, and saying to Zion, 'You are my people.'"
ISA|51|17|Wake yourself, wake yourself, stand up, O Jerusalem, you who have drunk from the hand of the LORD the cup of his wrath, who have drunk to the dregs the bowl, the cup of staggering.
ISA|51|18|There is none to guide her among all the sons she has borne; there is none to take her by the hand among all the sons she has brought up.
ISA|51|19|These two things have happened to you- who will console you?- devastation and destruction, famine and sword; who will comfort you?
ISA|51|20|Your sons have fainted; they lie at the head of every street like an antelope in a net; they are full of the wrath of the LORD, the rebuke of your God.
ISA|51|21|Therefore hear this, you who are afflicted, who are drunk, but not with wine:
ISA|51|22|Thus says your Lord, the LORD, your God who pleads the cause of his people: "Behold, I have taken from your hand the cup of staggering; the bowl of my wrath you shall drink no more;
ISA|51|23|and I will put it into the hand of your tormentors, who have said to you, 'Bow down, that we may pass over'; and you have made your back like the ground and like the street for them to pass over."
ISA|52|1|Awake, awake, put on your strength, O Zion; put on your beautiful garments, O Jerusalem, the holy city; for there shall no more come into you the uncircumcised and the unclean.
ISA|52|2|Shake yourself from the dust and arise; be seated, O Jerusalem; loose the bonds from your neck, O captive daughter of Zion.
ISA|52|3|For thus says the LORD: "You were sold for nothing, and you shall be redeemed without money."
ISA|52|4|For thus says the Lord GOD: "My people went down at the first into Egypt to sojourn there, and the Assyrian oppressed them for nothing.
ISA|52|5|Now therefore what have I here," declares the LORD, "seeing that my people are taken away for nothing? Their rulers wail," declares the LORD, "and continually all the day my name is despised.
ISA|52|6|Therefore my people shall know my name. Therefore in that day they shall know that it is I who speak; here am I."
ISA|52|7|How beautiful upon the mountains are the feet of him who brings good news, who publishes peace, who brings good news of happiness, who publishes salvation, who says to Zion, "Your God reigns."
ISA|52|8|The voice of your watchmen- they lift up their voice; together they sing for joy; for eye to eye they see the return of the LORD to Zion.
ISA|52|9|Break forth together into singing, you waste places of Jerusalem, for the LORD has comforted his people; he has redeemed Jerusalem.
ISA|52|10|The LORD has bared his holy arm before the eyes of all the nations, and all the ends of the earth shall see the salvation of our God.
ISA|52|11|Depart, depart, go out from there; touch no unclean thing; go out from the midst of her; purify yourselves, you who bear the vessels of the LORD.
ISA|52|12|For you shall not go out in haste, and you shall not go in flight, for the LORD will go before you, and the God of Israel will be your rear guard.
ISA|52|13|Behold, my servant shall act wisely; he shall be high and lifted up, and shall be exalted.
ISA|52|14|As many were astonished at you- his appearance was so marred, beyond human semblance, and his form beyond that of the children of mankind-
ISA|52|15|so shall he sprinkle many nations; kings shall shut their mouths because of him; for that which has not been told them they see, and that which they have not heard they understand.
ISA|53|1|Who has believed what they heard from us? And to whom has the arm of the LORD been revealed?
ISA|53|2|For he grew up before him like a young plant, and like a root out of dry ground; he had no form or majesty that we should look at him, and no beauty that we should desire him.
ISA|53|3|He was despised and rejected by men; a man of sorrows, and acquainted with grief; and as one from whom men hide their faces he was despised, and we esteemed him not.
ISA|53|4|Surely he has borne our griefs and carried our sorrows; yet we esteemed him stricken, smitten by God, and afflicted.
ISA|53|5|But he was wounded for our transgressions; he was crushed for our iniquities; upon him was the chastisement that brought us peace, and with his stripes we are healed.
ISA|53|6|All we like sheep have gone astray; we have turned every one to his own way; and the LORD has laid on him the iniquity of us all.
ISA|53|7|He was oppressed, and he was afflicted, yet he opened not his mouth; like a lamb that is led to the slaughter, and like a sheep that before its shearers is silent, so he opened not his mouth.
ISA|53|8|By oppression and judgment he was taken away; and as for his generation, who considered that he was cut off out of the land of the living, stricken for the transgression of my people?
ISA|53|9|And they made his grave with the wicked and with a rich man in his death, although he had done no violence, and there was no deceit in his mouth.
ISA|53|10|Yet it was the will of the LORD to crush him; he has put him to grief; when his soul makes an offering for sin, he shall see his offspring; he shall prolong his days; the will of the LORD shall prosper in his hand.
ISA|53|11|Out of the anguish of his soul he shall see and be satisfied; by his knowledge shall the righteous one, my servant, make many to be accounted righteous, and he shall bear their iniquities.
ISA|53|12|Therefore I will divide him a portion with the many, and he shall divide the spoil with the strong, because he poured out his soul to death and was numbered with the transgressors; yet he bore the sin of many, and makes intercession for the transgressors.
ISA|54|1|"Sing, O barren one, who did not bear; break forth into singing and cry aloud, you who have not been in labor! For the children of the desolate one will be more than the children of her who is married," says the LORD.
ISA|54|2|"Enlarge the place of your tent, and let the curtains of your habitations be stretched out; do not hold back; lengthen your cords and strengthen your stakes.
ISA|54|3|For you will spread abroad to the right and to the left, and your offspring will possess the nations and will people the desolate cities.
ISA|54|4|"Fear not, for you will not be ashamed; be not confounded, for you will not be disgraced; for you will forget the shame of your youth, and the reproach of your widowhood you will remember no more.
ISA|54|5|For your Maker is your husband, the LORD of hosts is his name; and the Holy One of Israel is your Redeemer, the God of the whole earth he is called.
ISA|54|6|For the LORD has called you like a wife deserted and grieved in spirit, like a wife of youth when she is cast off, says your God.
ISA|54|7|For a brief moment I deserted you, but with great compassion I will gather you.
ISA|54|8|In overflowing anger for a moment I hid my face from you, but with everlasting love I will have compassion on you," says the LORD, your Redeemer.
ISA|54|9|"This is like the days of Noah to me: as I swore that the waters of Noah should no more go over the earth, so I have sworn that I will not be angry with you, and will not rebuke you.
ISA|54|10|For the mountains may depart and the hills be removed, but my steadfast love shall not depart from you, and my covenant of peace shall not be removed," says the LORD, who has compassion on you.
ISA|54|11|"O afflicted one, storm-tossed and not comforted, behold, I will set your stones in antimony, and lay your foundations with sapphires.
ISA|54|12|I will make your pinnacles of agate, your gates of carbuncles, and all your wall of precious stones.
ISA|54|13|All your children shall be taught by the LORD, and great shall be the peace of your children.
ISA|54|14|In righteousness you shall be established; you shall be far from oppression, for you shall not fear; and from terror, for it shall not come near you.
ISA|54|15|If anyone stirs up strife, it is not from me; whoever stirs up strife with you shall fall because of you.
ISA|54|16|Behold, I have created the smith who blows the fire of coals and produces a weapon for its purpose. I have also created the ravager to destroy;
ISA|54|17|no weapon that is fashioned against you shall succeed, and you shall confute every tongue that rises against you in judgment. This is the heritage of the servants of the LORD and their vindication from me, declares the LORD."
ISA|55|1|"Come, everyone who thirsts, come to the waters; and he who has no money, come, buy and eat! Come, buy wine and milk without money and without price.
ISA|55|2|Why do you spend your money for that which is not bread, and your labor for that which does not satisfy? Listen diligently to me, and eat what is good, and delight yourselves in rich food.
ISA|55|3|Incline your ear, and come to me; hear, that your soul may live; and I will make with you an everlasting covenant, my steadfast, sure love for David.
ISA|55|4|Behold, I made him a witness to the peoples, a leader and commander for the peoples.
ISA|55|5|Behold, you shall call a nation that you do not know, and a nation that did not know you shall run to you, because of the LORD your God, and of the Holy One of Israel, for he has glorified you.
ISA|55|6|"Seek the LORD while he may be found; call upon him while he is near;
ISA|55|7|let the wicked forsake his way, and the unrighteous man his thoughts; let him return to the LORD, that he may have compassion on him, and to our God, for he will abundantly pardon.
ISA|55|8|For my thoughts are not your thoughts, neither are your ways my ways, declares the LORD.
ISA|55|9|For as the heavens are higher than the earth, so are my ways higher than your ways and my thoughts than your thoughts.
ISA|55|10|"For as the rain and the snow come down from heaven and do not return there but water the earth, making it bring forth and sprout, giving seed to the sower and bread to the eater,
ISA|55|11|so shall my word be that goes out from my mouth; it shall not return to me empty, but it shall accomplish that which I purpose, and shall succeed in the thing for which I sent it.
ISA|55|12|"For you shall go out in joy and be led forth in peace; the mountains and the hills before you shall break forth into singing, and all the trees of the field shall clap their hands.
ISA|55|13|Instead of the thorn shall come up the cypress; instead of the brier shall come up the myrtle; and it shall make a name for the LORD, an everlasting sign that shall not be cut off."
ISA|56|1|Thus says the LORD:"Keep justice, and do righteousness, for soon my salvation will come, and my deliverance be revealed.
ISA|56|2|Blessed is the man who does this, and the son of man who holds it fast, who keeps the Sabbath, not profaning it, and keeps his hand from doing any evil."
ISA|56|3|Let not the foreigner who has joined himself to the LORD say, "The LORD will surely separate me from his people"; and let not the eunuch say, "Behold, I am a dry tree."
ISA|56|4|For thus says the LORD: "To the eunuchs who keep my Sabbaths, who choose the things that please me and hold fast my covenant,
ISA|56|5|I will give in my house and within my walls a monument and a name better than sons and daughters; I will give them an everlasting name that shall not be cut off.
ISA|56|6|"And the foreigners who join themselves to the LORD, to minister to him, to love the name of the LORD, and to be his servants, everyone who keeps the Sabbath and does not profane it, and holds fast my covenant-
ISA|56|7|these I will bring to my holy mountain, and make them joyful in my house of prayer; their burnt offerings and their sacrifices will be accepted on my altar; for my house shall be called a house of prayer for all peoples."
ISA|56|8|The Lord GOD, who gathers the outcasts of Israel, declares, "I will gather yet others to him besides those already gathered."
ISA|56|9|All you beasts of the field, come to devour- all you beasts in the forest.
ISA|56|10|His watchmen are blind; they are all without knowledge; they are all silent dogs; they cannot bark, dreaming, lying down, loving to slumber.
ISA|56|11|The dogs have a mighty appetite; they never have enough. But they are shepherds who have no understanding; they have all turned to their own way, each to his own gain, one and all.
ISA|56|12|"Come," they say, "let me get wine; let us fill ourselves with strong drink; and tomorrow will be like this day, great beyond measure."
ISA|57|1|The righteous man perishes, and no one lays it to heart; devout men are taken away, while no one understands. For the righteous man is taken away from calamity;
ISA|57|2|he enters into peace; they rest in their beds who walk in their uprightness.
ISA|57|3|But you, draw near, sons of the sorceress, offspring of the adulterer and the loose woman.
ISA|57|4|Whom are you mocking? Against whom do you open your mouth wide and stick out your tongue? Are you not children of transgression, the offspring of deceit,
ISA|57|5|you who burn with lust among the oaks, under every green tree, who slaughter your children in the valleys, under the clefts of the rocks?
ISA|57|6|Among the smooth stones of the valley is your portion; they, they, are your lot; to them you have poured out a drink offering, you have brought a grain offering. Shall I relent for these things?
ISA|57|7|On a high and lofty mountain you have set your bed, and there you went up to offer sacrifice.
ISA|57|8|Behind the door and the doorpost you have set up your memorial; for, deserting me, you have uncovered your bed, you have gone up to it, you have made it wide; and you have made a covenant for yourself with them, you have loved their bed, you have looked on nakedness.
ISA|57|9|You journeyed to the king with oil and multiplied your perfumes; you sent your envoys far off, and sent down even to Sheol.
ISA|57|10|You were wearied with the length of your way, but you did not say, "It is hopeless"; you found new life for your strength, and so you were not faint.
ISA|57|11|Whom did you dread and fear, so that you lied, and did not remember me, did not lay it to heart? Have I not held my peace, even for a long time, and you do not fear me?
ISA|57|12|I will declare your righteousness and your deeds, but they will not profit you.
ISA|57|13|When you cry out, let your collection of idols deliver you! The wind will carry them off, a breath will take them away. But he who takes refuge in me shall possess the land and shall inherit my holy mountain.
ISA|57|14|And it shall be said, "Build up, build up, prepare the way, remove every obstruction from my people's way."
ISA|57|15|For thus says the One who is high and lifted up, who inhabits eternity, whose name is Holy: "I dwell in the high and holy place, and also with him who is of a contrite and lowly spirit, to revive the spirit of the lowly, and to revive the heart of the contrite.
ISA|57|16|For I will not contend forever, nor will I always be angry; for the spirit would grow faint before me, and the breath of life that I made.
ISA|57|17|Because of the iniquity of his unjust gain I was angry, I struck him; I hid my face and was angry, but he went on backsliding in the way of his own heart.
ISA|57|18|I have seen his ways, but I will heal him; I will lead him and restore comfort to him and his mourners,
ISA|57|19|creating the fruit of the lips. Peace, peace, to the far and to the near," says the LORD, "and I will heal him.
ISA|57|20|But the wicked are like the tossing sea; for it cannot be quiet, and its waters toss up mire and dirt.
ISA|57|21|There is no peace," says my God, "for the wicked."
ISA|58|1|"Cry aloud; do not hold back; lift up your voice like a trumpet; declare to my people their transgression, to the house of Jacob their sins.
ISA|58|2|Yet they seek me daily and delight to know my ways, as if they were a nation that did righteousness and did not forsake the judgment of their God; they ask of me righteous judgments; they delight to draw near to God.
ISA|58|3|'Why have we fasted, and you see it not? Why have we humbled ourselves, and you take no knowledge of it?' Behold, in the day of your fast you seek your own pleasure, and oppress all your workers.
ISA|58|4|Behold, you fast only to quarrel and to fight and to hit with a wicked fist. Fasting like yours this day will not make your voice to be heard on high.
ISA|58|5|Is such the fast that I choose, a day for a person to humble himself? Is it to bow down his head like a reed, and to spread sackcloth and ashes under him? Will you call this a fast, and a day acceptable to the LORD?
ISA|58|6|"Is not this the fast that I choose: to loose the bonds of wickedness, to undo the straps of the yoke, to let the oppressed go free, and to break every yoke?
ISA|58|7|Is it not to share your bread with the hungry and bring the homeless poor into your house; when you see the naked, to cover him, and not to hide yourself from your own flesh?
ISA|58|8|Then shall your light break forth like the dawn, and your healing shall spring up speedily; your righteousness shall go before you; the glory of the LORD shall be your rear guard.
ISA|58|9|Then you shall call, and the LORD will answer; you shall cry, and he will say, 'Here I am.' If you take away the yoke from your midst, the pointing of the finger, and speaking wickedness,
ISA|58|10|if you pour yourself out for the hungry and satisfy the desire of the afflicted, then shall your light rise in the darkness and your gloom be as the noonday.
ISA|58|11|And the LORD will guide you continually and satisfy your desire in scorched places and make your bones strong; and you shall be like a watered garden, like a spring of water, whose waters do not fail.
ISA|58|12|And your ancient ruins shall be rebuilt; you shall raise up the foundations of many generations; you shall be called the repairer of the breach, the restorer of streets to dwell in.
ISA|58|13|"If you turn back your foot from the Sabbath, from doing your pleasure on my holy day, and call the Sabbath a delight and the holy day of the LORD honorable; if you honor it, not going your own ways, or seeking your own pleasure, or talking idly;
ISA|58|14|then you shall take delight in the LORD, and I will make you ride on the heights of the earth; I will feed you with the heritage of Jacob your father, for the mouth of the LORD has spoken."
ISA|59|1|Behold, the LORD's hand is not shortened, that it cannot save, or his ear dull, that it cannot hear;
ISA|59|2|but your iniquities have made a separation between you and your God, and your sins have hidden his face from you so that he does not hear.
ISA|59|3|For your hands are defiled with blood and your fingers with iniquity; your lips have spoken lies; your tongue mutters wickedness.
ISA|59|4|No one enters suit justly; no one goes to law honestly; they rely on empty pleas, they speak lies, they conceive mischief and give birth to iniquity.
ISA|59|5|They hatch adders' eggs; they weave the spider's web; he who eats their eggs dies, and from one that is crushed a viper is hatched.
ISA|59|6|Their webs will not serve as clothing; men will not cover themselves with what they make. Their works are works of iniquity, and deeds of violence are in their hands.
ISA|59|7|Their feet run to evil, and they are swift to shed innocent blood; their thoughts are thoughts of iniquity; desolation and destruction are in their highways.
ISA|59|8|The way of peace they do not know, and there is no justice in their paths; they have made their roads crooked; no one who treads on them knows peace.
ISA|59|9|Therefore justice is far from us, and righteousness does not overtake us; we hope for light, and behold, darkness, and for brightness, but we walk in gloom.
ISA|59|10|We grope for the wall like the blind; we grope like those who have no eyes; we stumble at noon as in the twilight, among those in full vigor we are like dead men.
ISA|59|11|We all growl like bears; we moan and moan like doves; we hope for justice, but there is none; for salvation, but it is far from us.
ISA|59|12|For our transgressions are multiplied before you, and our sins testify against us; for our transgressions are with us, and we know our iniquities:
ISA|59|13|transgressing, and denying the LORD, and turning back from following our God, speaking oppression and revolt, conceiving and uttering from the heart lying words.
ISA|59|14|Justice is turned back, and righteousness stands afar off; for truth has stumbled in the public squares, and uprightness cannot enter.
ISA|59|15|Truth is lacking, and he who departs from evil makes himself a prey. The LORD saw it, and it displeased him that there was no justice.
ISA|59|16|He saw that there was no man, and wondered that there was no one to intercede; then his own arm brought him salvation, and his righteousness upheld him.
ISA|59|17|He put on righteousness as a breastplate, and a helmet of salvation on his head; he put on garments of vengeance for clothing, and wrapped himself in zeal as a cloak.
ISA|59|18|According to their deeds, so will he repay, wrath to his adversaries, repayment to his enemies; to the coastlands he will render repayment.
ISA|59|19|So they shall fear the name of the LORD from the west, and his glory from the rising of the sun; for he will come like a rushing stream, which the wind of the LORD drives.
ISA|59|20|"And a Redeemer will come to Zion, to those in Jacob who turn from transgression," declares the LORD.
ISA|59|21|"And as for me, this is my covenant with them," says the LORD: "My Spirit that is upon you, and my words that I have put in your mouth, shall not depart out of your mouth, or out of the mouth of your offspring, or out of the mouth of your children's offspring," says the LORD, "from this time forth and forevermore."
ISA|60|1|Arise, shine, for your light has come, and the glory of the LORD has risen upon you.
ISA|60|2|For behold, darkness shall cover the earth, and thick darkness the peoples; but the LORD will arise upon you, and his glory will be seen upon you.
ISA|60|3|And nations shall come to your light, and kings to the brightness of your rising.
ISA|60|4|Lift up your eyes all around, and see; they all gather together, they come to you; your sons shall come from far, and your daughters shall be carried on the hip.
ISA|60|5|Then you shall see and be radiant; your heart shall thrill and exult, because the abundance of the sea shall be turned to you, the wealth of the nations shall come to you.
ISA|60|6|A multitude of camels shall cover you, the young camels of Midian and Ephah; all those from Sheba shall come. They shall bring gold and frankincense, and shall bring good news, the praises of the LORD.
ISA|60|7|All the flocks of Kedar shall be gathered to you; the rams of Nebaioth shall minister to you; they shall come up with acceptance on my altar, and I will beautify my beautiful house.
ISA|60|8|Who are these that fly like a cloud, and like doves to their windows?
ISA|60|9|For the coastlands shall hope for me, the ships of Tarshish first, to bring your children from afar, their silver and gold with them, for the name of the LORD your God, and for the Holy One of Israel, because he has made you beautiful.
ISA|60|10|Foreigners shall build up your walls, and their kings shall minister to you; for in my wrath I struck you, but in my favor I have had mercy on you.
ISA|60|11|Your gates shall be open continually; day and night they shall not be shut, that people may bring to you the wealth of the nations, with their kings led in procession.
ISA|60|12|For the nation and kingdom that will not serve you shall perish; those nations shall be utterly laid waste.
ISA|60|13|The glory of Lebanon shall come to you, the cypress, the plane, and the pine, to beautify the place of my sanctuary, and I will make the place of my feet glorious.
ISA|60|14|The sons of those who afflicted you shall come bending low to you, and all who despised you shall bow down at your feet; they shall call you the City of the LORD, the Zion of the Holy One of Israel.
ISA|60|15|Whereas you have been forsaken and hated, with no one passing through, I will make you majestic forever, a joy from age to age.
ISA|60|16|You shall suck the milk of nations; you shall nurse at the breast of kings; and you shall know that I, the LORD, am your Savior and your Redeemer, the Mighty One of Jacob.
ISA|60|17|Instead of bronze I will bring gold, and instead of iron I will bring silver; instead of wood, bronze, instead of stones, iron. I will make your overseers peace and your taskmasters righteousness.
ISA|60|18|Violence shall no more be heard in your land, devastation or destruction within your borders; you shall call your walls Salvation, and your gates Praise.
ISA|60|19|The sun shall be no more your light by day, nor for brightness shall the moon give you light; but the LORD will be your everlasting light, and your God will be your glory.
ISA|60|20|Your sun shall no more go down, nor your moon withdraw itself; for the LORD will be your everlasting light, and your days of mourning shall be ended.
ISA|60|21|Your people shall all be righteous; they shall possess the land forever, the branch of my planting, the work of my hands, that I might be glorified.
ISA|60|22|The least one shall become a clan, and the smallest one a mighty nation; I am the LORD; in its time I will hasten it.
ISA|61|1|The Spirit of the Lord GOD is upon me, because the LORD has anointed me to bring good news to the poor; he has sent me to bind up the brokenhearted, to proclaim liberty to the captives, and the opening of the prison to those who are bound;
ISA|61|2|to proclaim the year of the LORD's favor, and the day of vengeance of our God; to comfort all who mourn;
ISA|61|3|to grant to those who mourn in Zion- to give them a beautiful headdress instead of ashes, the oil of gladness instead of mourning, the garment of praise instead of a faint spirit; that they may be called oaks of righteousness, the planting of the LORD, that he may be glorified.
ISA|61|4|They shall build up the ancient ruins; they shall raise up the former devastations; they shall repair the ruined cities, the devastations of many generations.
ISA|61|5|Strangers shall stand and tend your flocks; foreigners shall be your plowmen and vinedressers;
ISA|61|6|but you shall be called the priests of the LORD; they shall speak of you as the ministers of our God; you shall eat the wealth of the nations, and in their glory you shall boast.
ISA|61|7|Instead of your shame there shall be a double portion; instead of dishonor they shall rejoice in their lot; therefore in their land they shall possess a double portion; they shall have everlasting joy.
ISA|61|8|For I the LORD love justice; I hate robbery and wrong; I will faithfully give them their recompense, and I will make an everlasting covenant with them.
ISA|61|9|Their offspring shall be known among the nations, and their descendants in the midst of the peoples; all who see them shall acknowledge them, that they are an offspring the LORD has blessed.
ISA|61|10|I will greatly rejoice in the LORD; my soul shall exult in my God, for he has clothed me with the garments of salvation; he has covered me with the robe of righteousness, as a bridegroom decks himself like a priest with a beautiful headdress, and as a bride adorns herself with her jewels.
ISA|61|11|For as the earth brings forth its sprouts, and as a garden causes what is sown in it to sprout up, so the Lord GOD will cause righteousness and praise to sprout up before all the nations.
ISA|62|1|For Zion's sake I will not keep silent, and for Jerusalem's sake I will not be quiet, until her righteousness goes forth as brightness, and her salvation as a burning torch.
ISA|62|2|The nations shall see your righteousness, and all the kings your glory, and you shall be called by a new name that the mouth of the LORD will give.
ISA|62|3|You shall be a crown of beauty in the hand of the LORD, and a royal diadem in the hand of your God.
ISA|62|4|You shall no more be termed Forsaken, and your land shall no more be termed Desolate, but you shall be called My Delight Is in Her, and your land Married; for the LORD delights in you, and your land shall be married.
ISA|62|5|For as a young man marries a young woman, so shall your sons marry you, and as the bridegroom rejoices over the bride, so shall your God rejoice over you.
ISA|62|6|On your walls, O Jerusalem, I have set watchmen; all the day and all the night they shall never be silent. You who put the LORD in remembrance, take no rest,
ISA|62|7|and give him no rest until he establishes Jerusalem and makes it a praise in the earth.
ISA|62|8|The LORD has sworn by his right hand and by his mighty arm: "I will not again give your grain to be food for your enemies, and foreigners shall not drink your wine for which you have labored;
ISA|62|9|but those who garner it shall eat it and praise the LORD, and those who gather it shall drink it in the courts of my sanctuary."
ISA|62|10|Go through, go through the gates; prepare the way for the people; build up, build up the highway; clear it of stones; lift up a signal over the peoples.
ISA|62|11|Behold, the LORD has proclaimed to the end of the earth: Say to the daughter of Zion, "Behold, your salvation comes; behold, his reward is with him, and his recompense before him."
ISA|62|12|And they shall be called The Holy People, The Redeemed of the LORD; and you shall be called Sought Out, A City Not Forsaken.
ISA|63|1|Who is this who comes from Edom, in crimsoned garments from Bozrah, he who is splendid in his apparel, marching in the greatness of his strength? "It is I, speaking in righteousness, mighty to save."
ISA|63|2|Why is your apparel red, and your garments like his who treads in the winepress?
ISA|63|3|"I have trodden the winepress alone, and from the peoples no one was with me; I trod them in my anger and trampled them in my wrath; their lifeblood spattered on my garments, and stained all my apparel.
ISA|63|4|For the day of vengeance was in my heart, and my year of redemption had come.
ISA|63|5|I looked, but there was no one to help; I was appalled, but there was no one to uphold; so my own arm brought me salvation, and my wrath upheld me.
ISA|63|6|I trampled down the peoples in my anger; I made them drunk in my wrath, and I poured out their lifeblood on the earth."
ISA|63|7|I will recount the steadfast love of the LORD, the praises of the LORD, according to all that the LORD has granted us, and the great goodness to the house of Israel that he has granted them according to his compassion, according to the abundance of his steadfast love.
ISA|63|8|For he said, "Surely they are my people, children who will not deal falsely." And he became their Savior.
ISA|63|9|In all their affliction he was afflicted, and the angel of his presence saved them; in his love and in his pity he redeemed them; he lifted them up and carried them all the days of old.
ISA|63|10|But they rebelled and grieved his Holy Spirit; therefore he turned to be their enemy, and himself fought against them.
ISA|63|11|Then he remembered the days of old, of Moses and his people. Where is he who brought them up out of the sea with the shepherds of his flock? Where is he who put in the midst of them his Holy Spirit,
ISA|63|12|who caused his glorious arm to go at the right hand of Moses, who divided the waters before them to make for himself an everlasting name,
ISA|63|13|who led them through the depths? Like a horse in the desert, they did not stumble.
ISA|63|14|Like livestock that go down into the valley, the Spirit of the LORD gave them rest. So you led your people, to make for yourself a glorious name.
ISA|63|15|Look down from heaven and see, from your holy and beautiful habitation. Where are your zeal and your might? The stirring of your inner parts and your compassion are held back from me.
ISA|63|16|For you are our Father, though Abraham does not know us, and Israel does not acknowledge us; you, O LORD, are our Father, our Redeemer from of old is your name.
ISA|63|17|O LORD, why do you make us wander from your ways and harden our heart, so that we fear you not? Return for the sake of your servants, the tribes of your heritage.
ISA|63|18|Your holy people held possession for a little while; our adversaries have trampled down your sanctuary.
ISA|63|19|We have become like those over whom you have never ruled, like those who are not called by your name.
ISA|64|1|Oh that you would rend the heavens and come down, that the mountains might quake at your presence-
ISA|64|2|as when fire kindles brushwood and the fire causes water to boil- to make your name known to your adversaries, and that the nations might tremble at your presence!
ISA|64|3|When you did awesome things that we did not look for, you came down, the mountains quaked at your presence.
ISA|64|4|From of old no one has heard or perceived by the ear, no eye has seen a God besides you, who acts for those who wait for him.
ISA|64|5|You meet him who joyfully works righteousness, those who remember you in your ways. Behold, you were angry, and we sinned; in our sins we have been a long time, and shall we be saved?
ISA|64|6|We have all become like one who is unclean, and all our righteous deeds are like a polluted garment. We all fade like a leaf, and our iniquities, like the wind, take us away.
ISA|64|7|There is no one who calls upon your name, who rouses himself to take hold of you; for you have hidden your face from us, and have made us melt in the hand of our iniquities.
ISA|64|8|But now, O LORD, you are our Father; we are the clay, and you are our potter; we are all the work of your hand.
ISA|64|9|Be not so terribly angry, O LORD, and remember not iniquity forever. Behold, please look, we are all your people.
ISA|64|10|Your holy cities have become a wilderness; Zion has become a wilderness, Jerusalem a desolation.
ISA|64|11|Our holy and beautiful house, where our fathers praised you, has been burned by fire, and all our pleasant places have become ruins.
ISA|64|12|Will you restrain yourself at these things, O LORD? Will you keep silent, and afflict us so terribly?
ISA|65|1|I was ready to be sought by those who did not ask for me; I was ready to be found by those who did not seek me. I said, "Here am I, here am I," to a nation that was not called by my name.
ISA|65|2|I spread out my hands all the day to a rebellious people, who walk in a way that is not good, following their own devices;
ISA|65|3|a people who provoke me to my face continually, sacrificing in gardens and making offerings on bricks;
ISA|65|4|who sit in tombs, and spend the night in secret places; who eat pig's flesh, and broth of tainted meat is in their vessels;
ISA|65|5|who say, "Keep to yourself, do not come near me, for I am too holy for you." These are a smoke in my nostrils, a fire that burns all the day.
ISA|65|6|Behold, it is written before me: "I will not keep silent, but I will repay; I will indeed repay into their bosom
ISA|65|7|both your iniquities and your fathers' iniquities together, says the LORD; because they made offerings on the mountains and insulted me on the hills, I will measure into their bosom payment for their former deeds."
ISA|65|8|Thus says the LORD: "As the new wine is found in the cluster, and they say, 'Do not destroy it, for there is a blessing in it,' so I will do for my servants' sake, and not destroy them all.
ISA|65|9|I will bring forth offspring from Jacob, and from Judah possessors of my mountains; my chosen shall possess it, and my servants shall dwell there.
ISA|65|10|Sharon shall become a pasture for flocks, and the Valley of Achor a place for herds to lie down, for my people who have sought me.
ISA|65|11|But you who forsake the LORD, who forget my holy mountain, who set a table for Fortune and fill cups of mixed wine for Destiny,
ISA|65|12|I will destine you to the sword, and all of you shall bow down to the slaughter, because, when I called, you did not answer; when I spoke, you did not listen, but you did what was evil in my eyes and chose what I did not delight in."
ISA|65|13|Therefore thus says the Lord GOD: "Behold, my servants shall eat, but you shall be hungry; behold, my servants shall drink, but you shall be thirsty; behold, my servants shall rejoice, but you shall be put to shame;
ISA|65|14|behold, my servants shall sing for gladness of heart, but you shall cry out for pain of heart and shall wail for breaking of spirit.
ISA|65|15|You shall leave your name to my chosen for a curse, and the Lord GOD will put you to death, but his servants he will call by another name.
ISA|65|16|So that he who blesses himself in the land shall bless himself by the God of truth, and he who takes an oath in the land shall swear by the God of truth; because the former troubles are forgotten and are hidden from my eyes.
ISA|65|17|"For behold, I create new heavens and a new earth, and the former things shall not be remembered or come into mind.
ISA|65|18|But be glad and rejoice forever in that which I create; for behold, I create Jerusalem to be a joy, and her people to be a gladness.
ISA|65|19|I will rejoice in Jerusalem and be glad in my people; no more shall be heard in it the sound of weeping and the cry of distress.
ISA|65|20|No more shall there be in it an infant who lives but a few days, or an old man who does not fill out his days, for the young man shall die a hundred years old, and the sinner a hundred years old shall be accursed.
ISA|65|21|They shall build houses and inhabit them; they shall plant vineyards and eat their fruit.
ISA|65|22|They shall not build and another inhabit; they shall not plant and another eat; for like the days of a tree shall the days of my people be, and my chosen shall long enjoy the work of their hands.
ISA|65|23|They shall not labor in vain or bear children for calamity, for they shall be the offspring of the blessed of the LORD, and their descendants with them.
ISA|65|24|Before they call I will answer; while they are yet speaking I will hear.
ISA|65|25|The wolf and the lamb shall graze together; the lion shall eat straw like the ox, and dust shall be the serpent's food. They shall not hurt or destroy in all my holy mountain," says the LORD.
ISA|66|1|Thus says the LORD: "Heaven is my throne, and the earth is my footstool; what is the house that you would build for me, and what is the place of my rest?
ISA|66|2|All these things my hand has made, and so all these things came to be, declares the LORD. But this is the one to whom I will look: he who is humble and contrite in spirit and trembles at my word.
ISA|66|3|"He who slaughters an ox is like one who kills a man; he who sacrifices a lamb, like one who breaks a dog's neck; he who presents a grain offering, like one who offers pig's blood; he who makes a memorial offering of frankincense, like one who blesses an idol. These have chosen their own ways, and their soul delights in their abominations;
ISA|66|4|I also will choose harsh treatment for them and bring their fears upon them, because when I called, no one answered, when I spoke they did not listen; but they did what was evil in my eyes and chose that in which I did not delight."
ISA|66|5|Hear the word of the LORD, you who tremble at his word: "Your brothers who hate you and cast you out for my name's sake have said, 'Let the LORD be glorified, that we may see your joy'; but it is they who shall be put to shame.
ISA|66|6|"The sound of an uproar from the city! A sound from the temple! The sound of the LORD, rendering recompense to his enemies!
ISA|66|7|"Before she was in labor she gave birth; before her pain came upon her she delivered a son.
ISA|66|8|Who has heard such a thing? Who has seen such things? Shall a land be born in one day? Shall a nation be brought forth in one moment? For as soon as Zion was in labor she brought forth her children.
ISA|66|9|Shall I bring to the point of birth and not cause to bring forth?" says the LORD; "shall I, who cause to bring forth, shut the womb?" says your God.
ISA|66|10|"Rejoice with Jerusalem, and be glad for her, all you who love her; rejoice with her in joy, all you who mourn over her;
ISA|66|11|that you may nurse and be satisfied from her consoling breast; that you may drink deeply with delight from her glorious abundance."
ISA|66|12|For thus says the LORD: "Behold, I will extend peace to her like a river, and the glory of the nations like an overflowing stream; and you shall nurse, you shall be carried upon her hip, and bounced upon her knees.
ISA|66|13|As one whom his mother comforts, so I will comfort you; you shall be comforted in Jerusalem.
ISA|66|14|You shall see, and your heart shall rejoice; your bones shall flourish like the grass; and the hand of the LORD shall be known to his servants, and he shall show his indignation against his enemies.
ISA|66|15|"For behold, the LORD will come in fire, and his chariots like the whirlwind, to render his anger in fury, and his rebuke with flames of fire.
ISA|66|16|For by fire will the LORD enter into judgment, and by his sword, with all flesh; and those slain by the LORD shall be many.
ISA|66|17|"Those who sanctify and purify themselves to go into the gardens, following one in the midst, eating pig's flesh and the abomination and mice, shall come to an end together, declares the LORD.
ISA|66|18|"For I know their works and their thoughts, and the time is coming to gather all nations and tongues. And they shall come and shall see my glory,
ISA|66|19|and I will set a sign among them. And from them I will send survivors to the nations, to Tarshish, Pul, and Lud, who draw the bow, to Tubal and Javan, to the coastlands afar off, that have not heard my fame or seen my glory. And they shall declare my glory among the nations.
ISA|66|20|And they shall bring all your brothers from all the nations as an offering to the LORD, on horses and in chariots and in litters and on mules and on dromedaries, to my holy mountain Jerusalem, says the LORD, just as the Israelites bring their grain offering in a clean vessel to the house of the LORD.
ISA|66|21|And some of them also I will take for priests and for Levites, says the LORD.
ISA|66|22|"For as the new heavens and the new earth that I make shall remain before me, says the LORD, so shall your offspring and your name remain.
ISA|66|23|From new moon to new moon, and from Sabbath to Sabbath, all flesh shall come to worship before me, declares the LORD.
ISA|66|24|"And they shall go out and look on the dead bodies of the men who have rebelled against me. For their worm shall not die, their fire shall not be quenched, and they shall be an abhorrence to all flesh."
