1KGS|1|1|When King David was old and well advanced in years, he could not keep warm even when they put covers over him.
1KGS|1|2|So his servants said to him, "Let us look for a young virgin to attend the king and take care of him. She can lie beside him so that our lord the king may keep warm."
1KGS|1|3|Then they searched throughout Israel for a beautiful girl and found Abishag, a Shunammite, and brought her to the king.
1KGS|1|4|The girl was very beautiful; she took care of the king and waited on him, but the king had no intimate relations with her.
1KGS|1|5|Now Adonijah, whose mother was Haggith, put himself forward and said, "I will be king." So he got chariots and horses ready, with fifty men to run ahead of him.
1KGS|1|6|(His father had never interfered with him by asking, "Why do you behave as you do?" He was also very handsome and was born next after Absalom.)
1KGS|1|7|Adonijah conferred with Joab son of Zeruiah and with Abiathar the priest, and they gave him their support.
1KGS|1|8|But Zadok the priest, Benaiah son of Jehoiada, Nathan the prophet, Shimei and Rei and David's special guard did not join Adonijah.
1KGS|1|9|Adonijah then sacrificed sheep, cattle and fattened calves at the Stone of Zoheleth near En Rogel. He invited all his brothers, the king's sons, and all the men of Judah who were royal officials,
1KGS|1|10|but he did not invite Nathan the prophet or Benaiah or the special guard or his brother Solomon.
1KGS|1|11|Then Nathan asked Bathsheba, Solomon's mother, "Have you not heard that Adonijah, the son of Haggith, has become king without our lord David's knowing it?
1KGS|1|12|Now then, let me advise you how you can save your own life and the life of your son Solomon.
1KGS|1|13|Go in to King David and say to him, 'My lord the king, did you not swear to me your servant: "Surely Solomon your son shall be king after me, and he will sit on my throne"? Why then has Adonijah become king?'
1KGS|1|14|While you are still there talking to the king, I will come in and confirm what you have said."
1KGS|1|15|So Bathsheba went to see the aged king in his room, where Abishag the Shunammite was attending him.
1KGS|1|16|Bathsheba bowed low and knelt before the king. "What is it you want?" the king asked.
1KGS|1|17|She said to him, "My lord, you yourself swore to me your servant by the LORD your God: 'Solomon your son shall be king after me, and he will sit on my throne.'
1KGS|1|18|But now Adonijah has become king, and you, my lord the king, do not know about it.
1KGS|1|19|He has sacrificed great numbers of cattle, fattened calves, and sheep, and has invited all the king's sons, Abiathar the priest and Joab the commander of the army, but he has not invited Solomon your servant.
1KGS|1|20|My lord the king, the eyes of all Israel are on you, to learn from you who will sit on the throne of my lord the king after him.
1KGS|1|21|Otherwise, as soon as my lord the king is laid to rest with his fathers, I and my son Solomon will be treated as criminals."
1KGS|1|22|While she was still speaking with the king, Nathan the prophet arrived.
1KGS|1|23|And they told the king, "Nathan the prophet is here." So he went before the king and bowed with his face to the ground.
1KGS|1|24|Nathan said, "Have you, my lord the king, declared that Adonijah shall be king after you, and that he will sit on your throne?
1KGS|1|25|Today he has gone down and sacrificed great numbers of cattle, fattened calves, and sheep. He has invited all the king's sons, the commanders of the army and Abiathar the priest. Right now they are eating and drinking with him and saying, 'Long live King Adonijah!'
1KGS|1|26|But me your servant, and Zadok the priest, and Benaiah son of Jehoiada, and your servant Solomon he did not invite.
1KGS|1|27|Is this something my lord the king has done without letting his servants know who should sit on the throne of my lord the king after him?"
1KGS|1|28|Then King David said, "Call in Bathsheba." So she came into the king's presence and stood before him.
1KGS|1|29|The king then took an oath: "As surely as the LORD lives, who has delivered me out of every trouble,
1KGS|1|30|I will surely carry out today what I swore to you by the LORD, the God of Israel: Solomon your son shall be king after me, and he will sit on my throne in my place."
1KGS|1|31|Then Bathsheba bowed low with her face to the ground and, kneeling before the king, said, "May my lord King David live forever!"
1KGS|1|32|King David said, "Call in Zadok the priest, Nathan the prophet and Benaiah son of Jehoiada." When they came before the king,
1KGS|1|33|he said to them: "Take your lord's servants with you and set Solomon my son on my own mule and take him down to Gihon.
1KGS|1|34|There have Zadok the priest and Nathan the prophet anoint him king over Israel. Blow the trumpet and shout, 'Long live King Solomon!'
1KGS|1|35|Then you are to go up with him, and he is to come and sit on my throne and reign in my place. I have appointed him ruler over Israel and Judah."
1KGS|1|36|Benaiah son of Jehoiada answered the king, "Amen! May the LORD, the God of my lord the king, so declare it.
1KGS|1|37|As the LORD was with my lord the king, so may he be with Solomon to make his throne even greater than the throne of my lord King David!"
1KGS|1|38|So Zadok the priest, Nathan the prophet, Benaiah son of Jehoiada, the Kerethites and the Pelethites went down and put Solomon on King David's mule and escorted him to Gihon.
1KGS|1|39|Zadok the priest took the horn of oil from the sacred tent and anointed Solomon. Then they sounded the trumpet and all the people shouted, "Long live King Solomon!"
1KGS|1|40|And all the people went up after him, playing flutes and rejoicing greatly, so that the ground shook with the sound.
1KGS|1|41|Adonijah and all the guests who were with him heard it as they were finishing their feast. On hearing the sound of the trumpet, Joab asked, "What's the meaning of all the noise in the city?"
1KGS|1|42|Even as he was speaking, Jonathan son of Abiathar the priest arrived. Adonijah said, "Come in. A worthy man like you must be bringing good news."
1KGS|1|43|"Not at all!" Jonathan answered. "Our lord King David has made Solomon king.
1KGS|1|44|The king has sent with him Zadok the priest, Nathan the prophet, Benaiah son of Jehoiada, the Kerethites and the Pelethites, and they have put him on the king's mule,
1KGS|1|45|and Zadok the priest and Nathan the prophet have anointed him king at Gihon. From there they have gone up cheering, and the city resounds with it. That's the noise you hear.
1KGS|1|46|Moreover, Solomon has taken his seat on the royal throne.
1KGS|1|47|Also, the royal officials have come to congratulate our lord King David, saying, 'May your God make Solomon's name more famous than yours and his throne greater than yours!' And the king bowed in worship on his bed
1KGS|1|48|and said, 'Praise be to the LORD, the God of Israel, who has allowed my eyes to see a successor on my throne today.'"
1KGS|1|49|At this, all Adonijah's guests rose in alarm and dispersed.
1KGS|1|50|But Adonijah, in fear of Solomon, went and took hold of the horns of the altar.
1KGS|1|51|Then Solomon was told, "Adonijah is afraid of King Solomon and is clinging to the horns of the altar. He says, 'Let King Solomon swear to me today that he will not put his servant to death with the sword.'"
1KGS|1|52|Solomon replied, "If he shows himself to be a worthy man, not a hair of his head will fall to the ground; but if evil is found in him, he will die."
1KGS|1|53|Then King Solomon sent men, and they brought him down from the altar. And Adonijah came and bowed down to King Solomon, and Solomon said, "Go to your home."
1KGS|2|1|When the time drew near for David to die, he gave a charge to Solomon his son.
1KGS|2|2|"I am about to go the way of all the earth," he said. "So be strong, show yourself a man,
1KGS|2|3|and observe what the LORD your God requires: Walk in his ways, and keep his decrees and commands, his laws and requirements, as written in the Law of Moses, so that you may prosper in all you do and wherever you go,
1KGS|2|4|and that the LORD may keep his promise to me: 'If your descendants watch how they live, and if they walk faithfully before me with all their heart and soul, you will never fail to have a man on the throne of Israel.'
1KGS|2|5|"Now you yourself know what Joab son of Zeruiah did to me-what he did to the two commanders of Israel's armies, Abner son of Ner and Amasa son of Jether. He killed them, shedding their blood in peacetime as if in battle, and with that blood stained the belt around his waist and the sandals on his feet.
1KGS|2|6|Deal with him according to your wisdom, but do not let his gray head go down to the grave in peace.
1KGS|2|7|"But show kindness to the sons of Barzillai of Gilead and let them be among those who eat at your table. They stood by me when I fled from your brother Absalom.
1KGS|2|8|"And remember, you have with you Shimei son of Gera, the Benjamite from Bahurim, who called down bitter curses on me the day I went to Mahanaim. When he came down to meet me at the Jordan, I swore to him by the LORD: 'I will not put you to death by the sword.'
1KGS|2|9|But now, do not consider him innocent. You are a man of wisdom; you will know what to do to him. Bring his gray head down to the grave in blood."
1KGS|2|10|Then David rested with his fathers and was buried in the City of David.
1KGS|2|11|He had reigned forty years over Israel-seven years in Hebron and thirty-three in Jerusalem.
1KGS|2|12|So Solomon sat on the throne of his father David, and his rule was firmly established.
1KGS|2|13|Now Adonijah, the son of Haggith, went to Bathsheba, Solomon's mother. Bathsheba asked him, "Do you come peacefully?" He answered, "Yes, peacefully."
1KGS|2|14|Then he added, "I have something to say to you.You may say it," she replied.
1KGS|2|15|"As you know," he said, "the kingdom was mine. All Israel looked to me as their king. But things changed, and the kingdom has gone to my brother; for it has come to him from the LORD.
1KGS|2|16|Now I have one request to make of you. Do not refuse me.You may make it," she said.
1KGS|2|17|So he continued, "Please ask King Solomon-he will not refuse you-to give me Abishag the Shunammite as my wife."
1KGS|2|18|"Very well," Bathsheba replied, "I will speak to the king for you."
1KGS|2|19|When Bathsheba went to King Solomon to speak to him for Adonijah, the king stood up to meet her, bowed down to her and sat down on his throne. He had a throne brought for the king's mother, and she sat down at his right hand.
1KGS|2|20|"I have one small request to make of you," she said. "Do not refuse me." The king replied, "Make it, my mother; I will not refuse you."
1KGS|2|21|So she said, "Let Abishag the Shunammite be given in marriage to your brother Adonijah."
1KGS|2|22|King Solomon answered his mother, "Why do you request Abishag the Shunammite for Adonijah? You might as well request the kingdom for him-after all, he is my older brother-yes, for him and for Abiathar the priest and Joab son of Zeruiah!"
1KGS|2|23|Then King Solomon swore by the LORD: "May God deal with me, be it ever so severely, if Adonijah does not pay with his life for this request!
1KGS|2|24|And now, as surely as the LORD lives-he who has established me securely on the throne of my father David and has founded a dynasty for me as he promised-Adonijah shall be put to death today!"
1KGS|2|25|So King Solomon gave orders to Benaiah son of Jehoiada, and he struck down Adonijah and he died.
1KGS|2|26|To Abiathar the priest the king said, "Go back to your fields in Anathoth. You deserve to die, but I will not put you to death now, because you carried the ark of the Sovereign LORD before my father David and shared all my father's hardships."
1KGS|2|27|So Solomon removed Abiathar from the priesthood of the LORD, fulfilling the word the LORD had spoken at Shiloh about the house of Eli.
1KGS|2|28|When the news reached Joab, who had conspired with Adonijah though not with Absalom, he fled to the tent of the LORD and took hold of the horns of the altar.
1KGS|2|29|King Solomon was told that Joab had fled to the tent of the LORD and was beside the altar. Then Solomon ordered Benaiah son of Jehoiada, "Go, strike him down!"
1KGS|2|30|So Benaiah entered the tent of the LORD and said to Joab, "The king says, 'Come out!'" But he answered, "No, I will die here." Benaiah reported to the king, "This is how Joab answered me."
1KGS|2|31|Then the king commanded Benaiah, "Do as he says. Strike him down and bury him, and so clear me and my father's house of the guilt of the innocent blood that Joab shed.
1KGS|2|32|The LORD will repay him for the blood he shed, because without the knowledge of my father David he attacked two men and killed them with the sword. Both of them-Abner son of Ner, commander of Israel's army, and Amasa son of Jether, commander of Judah's army-were better men and more upright than he.
1KGS|2|33|May the guilt of their blood rest on the head of Joab and his descendants forever. But on David and his descendants, his house and his throne, may there be the LORD's peace forever."
1KGS|2|34|So Benaiah son of Jehoiada went up and struck down Joab and killed him, and he was buried on his own land in the desert.
1KGS|2|35|The king put Benaiah son of Jehoiada over the army in Joab's position and replaced Abiathar with Zadok the priest.
1KGS|2|36|Then the king sent for Shimei and said to him, "Build yourself a house in Jerusalem and live there, but do not go anywhere else.
1KGS|2|37|The day you leave and cross the Kidron Valley, you can be sure you will die; your blood will be on your own head."
1KGS|2|38|Shimei answered the king, "What you say is good. Your servant will do as my lord the king has said." And Shimei stayed in Jerusalem for a long time.
1KGS|2|39|But three years later, two of Shimei's slaves ran off to Achish son of Maacah, king of Gath, and Shimei was told, "Your slaves are in Gath."
1KGS|2|40|At this, he saddled his donkey and went to Achish at Gath in search of his slaves. So Shimei went away and brought the slaves back from Gath.
1KGS|2|41|When Solomon was told that Shimei had gone from Jerusalem to Gath and had returned,
1KGS|2|42|the king summoned Shimei and said to him, "Did I not make you swear by the LORD and warn you, 'On the day you leave to go anywhere else, you can be sure you will die'? At that time you said to me, 'What you say is good. I will obey.'
1KGS|2|43|Why then did you not keep your oath to the LORD and obey the command I gave you?"
1KGS|2|44|The king also said to Shimei, "You know in your heart all the wrong you did to my father David. Now the LORD will repay you for your wrongdoing.
1KGS|2|45|But King Solomon will be blessed, and David's throne will remain secure before the LORD forever."
1KGS|2|46|Then the king gave the order to Benaiah son of Jehoiada, and he went out and struck Shimei down and killed him. The kingdom was now firmly established in Solomon's hands.
1KGS|3|1|Solomon made an alliance with Pharaoh king of Egypt and married his daughter. He brought her to the City of David until he finished building his palace and the temple of the LORD, and the wall around Jerusalem.
1KGS|3|2|The people, however, were still sacrificing at the high places, because a temple had not yet been built for the Name of the LORD.
1KGS|3|3|Solomon showed his love for the LORD by walking according to the statutes of his father David, except that he offered sacrifices and burned incense on the high places.
1KGS|3|4|The king went to Gibeon to offer sacrifices, for that was the most important high place, and Solomon offered a thousand burnt offerings on that altar.
1KGS|3|5|At Gibeon the LORD appeared to Solomon during the night in a dream, and God said, "Ask for whatever you want me to give you."
1KGS|3|6|Solomon answered, "You have shown great kindness to your servant, my father David, because he was faithful to you and righteous and upright in heart. You have continued this great kindness to him and have given him a son to sit on his throne this very day.
1KGS|3|7|"Now, O LORD my God, you have made your servant king in place of my father David. But I am only a little child and do not know how to carry out my duties.
1KGS|3|8|Your servant is here among the people you have chosen, a great people, too numerous to count or number.
1KGS|3|9|So give your servant a discerning heart to govern your people and to distinguish between right and wrong. For who is able to govern this great people of yours?"
1KGS|3|10|The Lord was pleased that Solomon had asked for this.
1KGS|3|11|So God said to him, "Since you have asked for this and not for long life or wealth for yourself, nor have asked for the death of your enemies but for discernment in administering justice,
1KGS|3|12|I will do what you have asked. I will give you a wise and discerning heart, so that there will never have been anyone like you, nor will there ever be.
1KGS|3|13|Moreover, I will give you what you have not asked for-both riches and honor-so that in your lifetime you will have no equal among kings.
1KGS|3|14|And if you walk in my ways and obey my statutes and commands as David your father did, I will give you a long life."
1KGS|3|15|Then Solomon awoke-and he realized it had been a dream. He returned to Jerusalem, stood before the ark of the Lord's covenant and sacrificed burnt offerings and fellowship offerings. Then he gave a feast for all his court.
1KGS|3|16|Now two prostitutes came to the king and stood before him.
1KGS|3|17|One of them said, "My lord, this woman and I live in the same house. I had a baby while she was there with me.
1KGS|3|18|The third day after my child was born, this woman also had a baby. We were alone; there was no one in the house but the two of us.
1KGS|3|19|"During the night this woman's son died because she lay on him.
1KGS|3|20|So she got up in the middle of the night and took my son from my side while I your servant was asleep. She put him by her breast and put her dead son by my breast.
1KGS|3|21|The next morning, I got up to nurse my son-and he was dead! But when I looked at him closely in the morning light, I saw that it wasn't the son I had borne."
1KGS|3|22|The other woman said, "No! The living one is my son; the dead one is yours." But the first one insisted, "No! The dead one is yours; the living one is mine." And so they argued before the king.
1KGS|3|23|The king said, "This one says, 'My son is alive and your son is dead,' while that one says, 'No! Your son is dead and mine is alive.'"
1KGS|3|24|Then the king said, "Bring me a sword." So they brought a sword for the king.
1KGS|3|25|He then gave an order: "Cut the living child in two and give half to one and half to the other."
1KGS|3|26|The woman whose son was alive was filled with compassion for her son and said to the king, "Please, my lord, give her the living baby! Don't kill him!" But the other said, "Neither I nor you shall have him. Cut him in two!"
1KGS|3|27|Then the king gave his ruling: "Give the living baby to the first woman. Do not kill him; she is his mother."
1KGS|3|28|When all Israel heard the verdict the king had given, they held the king in awe, because they saw that he had wisdom from God to administer justice.
1KGS|4|1|So King Solomon ruled over all Israel.
1KGS|4|2|And these were his chief officials: Azariah son of Zadok-the priest;
1KGS|4|3|Elihoreph and Ahijah, sons of Shisha-secretaries; Jehoshaphat son of Ahilud-recorder;
1KGS|4|4|Benaiah son of Jehoiada-commander in chief; Zadok and Abiathar-priests;
1KGS|4|5|Azariah son of Nathan-in charge of the district officers; Zabud son of Nathan-a priest and personal adviser to the king;
1KGS|4|6|Ahishar-in charge of the palace; Adoniram son of Abda-in charge of forced labor.
1KGS|4|7|Solomon also had twelve district governors over all Israel, who supplied provisions for the king and the royal household. Each one had to provide supplies for one month in the year.
1KGS|4|8|These are their names: Ben-Hur-in the hill country of Ephraim;
1KGS|4|9|Ben-Deker-in Makaz, Shaalbim, Beth Shemesh and Elon Bethhanan;
1KGS|4|10|Ben-Hesed-in Arubboth (Socoh and all the land of Hepher were his);
1KGS|4|11|Ben-Abinadab-in Naphoth Dor (he was married to Taphath daughter of Solomon);
1KGS|4|12|Baana son of Ahilud-in Taanach and Megiddo, and in all of Beth Shan next to Zarethan below Jezreel, from Beth Shan to Abel Meholah across to Jokmeam;
1KGS|4|13|Ben-Geber-in Ramoth Gilead (the settlements of Jair son of Manasseh in Gilead were his, as well as the district of Argob in Bashan and its sixty large walled cities with bronze gate bars);
1KGS|4|14|Ahinadab son of Iddo-in Mahanaim;
1KGS|4|15|Ahimaaz-in Naphtali (he had married Basemath daughter of Solomon);
1KGS|4|16|Baana son of Hushai-in Asher and in Aloth;
1KGS|4|17|Jehoshaphat son of Paruah-in Issachar;
1KGS|4|18|Shimei son of Ela-in Benjamin;
1KGS|4|19|Geber son of Uri-in Gilead (the country of Sihon king of the Amorites and the country of Og king of Bashan). He was the only governor over the district.
1KGS|4|20|The people of Judah and Israel were as numerous as the sand on the seashore; they ate, they drank and they were happy.
1KGS|4|21|And Solomon ruled over all the kingdoms from the River to the land of the Philistines, as far as the border of Egypt. These countries brought tribute and were Solomon's subjects all his life.
1KGS|4|22|Solomon's daily provisions were thirty cors of fine flour and sixty cors of meal,
1KGS|4|23|ten head of stall-fed cattle, twenty of pasture-fed cattle and a hundred sheep and goats, as well as deer, gazelles, roebucks and choice fowl.
1KGS|4|24|For he ruled over all the kingdoms west of the River, from Tiphsah to Gaza, and had peace on all sides.
1KGS|4|25|During Solomon's lifetime Judah and Israel, from Dan to Beersheba, lived in safety, each man under his own vine and fig tree.
1KGS|4|26|Solomon had four thousand stalls for chariot horses, and twelve thousand horses.
1KGS|4|27|The district officers, each in his month, supplied provisions for King Solomon and all who came to the king's table. They saw to it that nothing was lacking.
1KGS|4|28|They also brought to the proper place their quotas of barley and straw for the chariot horses and the other horses.
1KGS|4|29|God gave Solomon wisdom and very great insight, and a breadth of understanding as measureless as the sand on the seashore.
1KGS|4|30|Solomon's wisdom was greater than the wisdom of all the men of the East, and greater than all the wisdom of Egypt.
1KGS|4|31|He was wiser than any other man, including Ethan the Ezrahite-wiser than Heman, Calcol and Darda, the sons of Mahol. And his fame spread to all the surrounding nations.
1KGS|4|32|He spoke three thousand proverbs and his songs numbered a thousand and five.
1KGS|4|33|He described plant life, from the cedar of Lebanon to the hyssop that grows out of walls. He also taught about animals and birds, reptiles and fish.
1KGS|4|34|Men of all nations came to listen to Solomon's wisdom, sent by all the kings of the world, who had heard of his wisdom.
1KGS|5|1|When Hiram king of Tyre heard that Solomon had been anointed king to succeed his father David, he sent his envoys to Solomon, because he had always been on friendly terms with David.
1KGS|5|2|Solomon sent back this message to Hiram:
1KGS|5|3|"You know that because of the wars waged against my father David from all sides, he could not build a temple for the Name of the LORD his God until the LORD put his enemies under his feet.
1KGS|5|4|But now the LORD my God has given me rest on every side, and there is no adversary or disaster.
1KGS|5|5|I intend, therefore, to build a temple for the Name of the LORD my God, as the LORD told my father David, when he said, 'Your son whom I will put on the throne in your place will build the temple for my Name.'
1KGS|5|6|"So give orders that cedars of Lebanon be cut for me. My men will work with yours, and I will pay you for your men whatever wages you set. You know that we have no one so skilled in felling timber as the Sidonians."
1KGS|5|7|When Hiram heard Solomon's message, he was greatly pleased and said, "Praise be to the LORD today, for he has given David a wise son to rule over this great nation."
1KGS|5|8|So Hiram sent word to Solomon: "I have received the message you sent me and will do all you want in providing the cedar and pine logs.
1KGS|5|9|My men will haul them down from Lebanon to the sea, and I will float them in rafts by sea to the place you specify. There I will separate them and you can take them away. And you are to grant my wish by providing food for my royal household."
1KGS|5|10|In this way Hiram kept Solomon supplied with all the cedar and pine logs he wanted,
1KGS|5|11|and Solomon gave Hiram twenty thousand cors of wheat as food for his household, in addition to twenty thousand baths, of pressed olive oil. Solomon continued to do this for Hiram year after year.
1KGS|5|12|The LORD gave Solomon wisdom, just as he had promised him. There were peaceful relations between Hiram and Solomon, and the two of them made a treaty.
1KGS|5|13|King Solomon conscripted laborers from all Israel-thirty thousand men.
1KGS|5|14|He sent them off to Lebanon in shifts of ten thousand a month, so that they spent one month in Lebanon and two months at home. Adoniram was in charge of the forced labor.
1KGS|5|15|Solomon had seventy thousand carriers and eighty thousand stonecutters in the hills,
1KGS|5|16|as well as thirty-three hundred foremen who supervised the project and directed the workmen.
1KGS|5|17|At the king's command they removed from the quarry large blocks of quality stone to provide a foundation of dressed stone for the temple.
1KGS|5|18|The craftsmen of Solomon and Hiram and the men of Gebal cut and prepared the timber and stone for the building of the temple.
1KGS|6|1|In the four hundred and eightieth year after the Israelites had come out of Egypt, in the fourth year of Solomon's reign over Israel, in the month of Ziv, the second month, he began to build the temple of the LORD.
1KGS|6|2|The temple that King Solomon built for the LORD was sixty cubits long, twenty wide and thirty high.
1KGS|6|3|The portico at the front of the main hall of the temple extended the width of the temple, that is twenty cubits, and projected ten cubits from the front of the temple.
1KGS|6|4|He made narrow clerestory windows in the temple.
1KGS|6|5|Against the walls of the main hall and inner sanctuary he built a structure around the building, in which there were side rooms.
1KGS|6|6|The lowest floor was five cubits wide, the middle floor six cubits and the third floor seven. He made offset ledges around the outside of the temple so that nothing would be inserted into the temple walls.
1KGS|6|7|In building the temple, only blocks dressed at the quarry were used, and no hammer, chisel or any other iron tool was heard at the temple site while it was being built.
1KGS|6|8|The entrance to the lowest floor was on the south side of the temple; a stairway led up to the middle level and from there to the third.
1KGS|6|9|So he built the temple and completed it, roofing it with beams and cedar planks.
1KGS|6|10|And he built the side rooms all along the temple. The height of each was five cubits, and they were attached to the temple by beams of cedar.
1KGS|6|11|The word of the LORD came to Solomon:
1KGS|6|12|"As for this temple you are building, if you follow my decrees, carry out my regulations and keep all my commands and obey them, I will fulfill through you the promise I gave to David your father.
1KGS|6|13|And I will live among the Israelites and will not abandon my people Israel."
1KGS|6|14|So Solomon built the temple and completed it.
1KGS|6|15|He lined its interior walls with cedar boards, paneling them from the floor of the temple to the ceiling, and covered the floor of the temple with planks of pine.
1KGS|6|16|He partitioned off twenty cubits at the rear of the temple with cedar boards from floor to ceiling to form within the temple an inner sanctuary, the Most Holy Place.
1KGS|6|17|The main hall in front of this room was forty cubits long.
1KGS|6|18|The inside of the temple was cedar, carved with gourds and open flowers. Everything was cedar; no stone was to be seen.
1KGS|6|19|He prepared the inner sanctuary within the temple to set the ark of the covenant of the LORD there.
1KGS|6|20|The inner sanctuary was twenty cubits long, twenty wide and twenty high. He overlaid the inside with pure gold, and he also overlaid the altar of cedar.
1KGS|6|21|Solomon covered the inside of the temple with pure gold, and he extended gold chains across the front of the inner sanctuary, which was overlaid with gold.
1KGS|6|22|So he overlaid the whole interior with gold. He also overlaid with gold the altar that belonged to the inner sanctuary.
1KGS|6|23|In the inner sanctuary he made a pair of cherubim of olive wood, each ten cubits high.
1KGS|6|24|One wing of the first cherub was five cubits long, and the other wing five cubits-ten cubits from wing tip to wing tip.
1KGS|6|25|The second cherub also measured ten cubits, for the two cherubim were identical in size and shape.
1KGS|6|26|The height of each cherub was ten cubits.
1KGS|6|27|He placed the cherubim inside the innermost room of the temple, with their wings spread out. The wing of one cherub touched one wall, while the wing of the other touched the other wall, and their wings touched each other in the middle of the room.
1KGS|6|28|He overlaid the cherubim with gold.
1KGS|6|29|On the walls all around the temple, in both the inner and outer rooms, he carved cherubim, palm trees and open flowers.
1KGS|6|30|He also covered the floors of both the inner and outer rooms of the temple with gold.
1KGS|6|31|For the entrance of the inner sanctuary he made doors of olive wood with five-sided jambs.
1KGS|6|32|And on the two olive wood doors he carved cherubim, palm trees and open flowers, and overlaid the cherubim and palm trees with beaten gold.
1KGS|6|33|In the same way he made four-sided jambs of olive wood for the entrance to the main hall.
1KGS|6|34|He also made two pine doors, each having two leaves that turned in sockets.
1KGS|6|35|He carved cherubim, palm trees and open flowers on them and overlaid them with gold hammered evenly over the carvings.
1KGS|6|36|And he built the inner courtyard of three courses of dressed stone and one course of trimmed cedar beams.
1KGS|6|37|The foundation of the temple of the LORD was laid in the fourth year, in the month of Ziv.
1KGS|6|38|In the eleventh year in the month of Bul, the eighth month, the temple was finished in all its details according to its specifications. He had spent seven years building it.
1KGS|7|1|It took Solomon thirteen years, however, to complete the construction of his palace.
1KGS|7|2|He built the Palace of the Forest of Lebanon a hundred cubits long, fifty wide and thirty high, with four rows of cedar columns supporting trimmed cedar beams.
1KGS|7|3|It was roofed with cedar above the beams that rested on the columns-forty-five beams, fifteen to a row.
1KGS|7|4|Its windows were placed high in sets of three, facing each other.
1KGS|7|5|All the doorways had rectangular frames; they were in the front part in sets of three, facing each other.
1KGS|7|6|He made a colonnade fifty cubits long and thirty wide. In front of it was a portico, and in front of that were pillars and an overhanging roof.
1KGS|7|7|He built the throne hall, the Hall of Justice, where he was to judge, and he covered it with cedar from floor to ceiling.
1KGS|7|8|And the palace in which he was to live, set farther back, was similar in design. Solomon also made a palace like this hall for Pharaoh's daughter, whom he had married.
1KGS|7|9|All these structures, from the outside to the great courtyard and from foundation to eaves, were made of blocks of high-grade stone cut to size and trimmed with a saw on their inner and outer faces.
1KGS|7|10|The foundations were laid with large stones of good quality, some measuring ten cubits and some eight.
1KGS|7|11|Above were high-grade stones, cut to size, and cedar beams.
1KGS|7|12|The great courtyard was surrounded by a wall of three courses of dressed stone and one course of trimmed cedar beams, as was the inner courtyard of the temple of the LORD with its portico.
1KGS|7|13|King Solomon sent to Tyre and brought Huram,
1KGS|7|14|whose mother was a widow from the tribe of Naphtali and whose father was a man of Tyre and a craftsman in bronze. Huram was highly skilled and experienced in all kinds of bronze work. He came to King Solomon and did all the work assigned to him.
1KGS|7|15|He cast two bronze pillars, each eighteen cubits high and twelve cubits around, by line.
1KGS|7|16|He also made two capitals of cast bronze to set on the tops of the pillars; each capital was five cubits high.
1KGS|7|17|A network of interwoven chains festooned the capitals on top of the pillars, seven for each capital.
1KGS|7|18|He made pomegranates in two rows encircling each network to decorate the capitals on top of the pillars. He did the same for each capital.
1KGS|7|19|The capitals on top of the pillars in the portico were in the shape of lilies, four cubits high.
1KGS|7|20|On the capitals of both pillars, above the bowl-shaped part next to the network, were the two hundred pomegranates in rows all around.
1KGS|7|21|He erected the pillars at the portico of the temple. The pillar to the south he named Jakin and the one to the north Boaz.
1KGS|7|22|The capitals on top were in the shape of lilies. And so the work on the pillars was completed.
1KGS|7|23|He made the Sea of cast metal, circular in shape, measuring ten cubits from rim to rim and five cubits high. It took a line of thirty cubits to measure around it.
1KGS|7|24|Below the rim, gourds encircled it-ten to a cubit. The gourds were cast in two rows in one piece with the Sea.
1KGS|7|25|The Sea stood on twelve bulls, three facing north, three facing west, three facing south and three facing east. The Sea rested on top of them, and their hindquarters were toward the center.
1KGS|7|26|It was a handbreadth in thickness, and its rim was like the rim of a cup, like a lily blossom. It held two thousand baths.
1KGS|7|27|He also made ten movable stands of bronze; each was four cubits long, four wide and three high.
1KGS|7|28|This is how the stands were made: They had side panels attached to uprights.
1KGS|7|29|On the panels between the uprights were lions, bulls and cherubim-and on the uprights as well. Above and below the lions and bulls were wreaths of hammered work.
1KGS|7|30|Each stand had four bronze wheels with bronze axles, and each had a basin resting on four supports, cast with wreaths on each side.
1KGS|7|31|On the inside of the stand there was an opening that had a circular frame one cubit deep. This opening was round, and with its basework it measured a cubit and a half. Around its opening there was engraving. The panels of the stands were square, not round.
1KGS|7|32|The four wheels were under the panels, and the axles of the wheels were attached to the stand. The diameter of each wheel was a cubit and a half.
1KGS|7|33|The wheels were made like chariot wheels; the axles, rims, spokes and hubs were all of cast metal.
1KGS|7|34|Each stand had four handles, one on each corner, projecting from the stand.
1KGS|7|35|At the top of the stand there was a circular band half a cubit deep. The supports and panels were attached to the top of the stand.
1KGS|7|36|He engraved cherubim, lions and palm trees on the surfaces of the supports and on the panels, in every available space, with wreaths all around.
1KGS|7|37|This is the way he made the ten stands. They were all cast in the same molds and were identical in size and shape.
1KGS|7|38|He then made ten bronze basins, each holding forty baths and measuring four cubits across, one basin to go on each of the ten stands.
1KGS|7|39|He placed five of the stands on the south side of the temple and five on the north. He placed the Sea on the south side, at the southeast corner of the temple.
1KGS|7|40|He also made the basins and shovels and sprinkling bowls. So Huram finished all the work he had undertaken for King Solomon in the temple of the LORD:
1KGS|7|41|the two pillars; the two bowl-shaped capitals on top of the pillars; the two sets of network decorating the two bowl-shaped capitals on top of the pillars;
1KGS|7|42|the four hundred pomegranates for the two sets of network (two rows of pomegranates for each network, decorating the bowl-shaped capitals on top of the pillars);
1KGS|7|43|the ten stands with their ten basins;
1KGS|7|44|the Sea and the twelve bulls under it;
1KGS|7|45|the pots, shovels and sprinkling bowls. All these objects that Huram made for King Solomon for the temple of the LORD were of burnished bronze.
1KGS|7|46|The king had them cast in clay molds in the plain of the Jordan between Succoth and Zarethan.
1KGS|7|47|Solomon left all these things unweighed, because there were so many; the weight of the bronze was not determined.
1KGS|7|48|Solomon also made all the furnishings that were in the LORD's temple: the golden altar; the golden table on which was the bread of the Presence;
1KGS|7|49|the lampstands of pure gold (five on the right and five on the left, in front of the inner sanctuary); the gold floral work and lamps and tongs;
1KGS|7|50|the pure gold basins, wick trimmers, sprinkling bowls, dishes and censers; and the gold sockets for the doors of the innermost room, the Most Holy Place, and also for the doors of the main hall of the temple.
1KGS|7|51|When all the work King Solomon had done for the temple of the LORD was finished, he brought in the things his father David had dedicated-the silver and gold and the furnishings-and he placed them in the treasuries of the LORD's temple.
1KGS|8|1|Then King Solomon summoned into his presence at Jerusalem the elders of Israel, all the heads of the tribes and the chiefs of the Israelite families, to bring up the ark of the LORD's covenant from Zion, the City of David.
1KGS|8|2|All the men of Israel came together to King Solomon at the time of the festival in the month of Ethanim, the seventh month.
1KGS|8|3|When all the elders of Israel had arrived, the priests took up the ark,
1KGS|8|4|and they brought up the ark of the LORD and the Tent of Meeting and all the sacred furnishings in it. The priests and Levites carried them up,
1KGS|8|5|and King Solomon and the entire assembly of Israel that had gathered about him were before the ark, sacrificing so many sheep and cattle that they could not be recorded or counted.
1KGS|8|6|The priests then brought the ark of the LORD's covenant to its place in the inner sanctuary of the temple, the Most Holy Place, and put it beneath the wings of the cherubim.
1KGS|8|7|The cherubim spread their wings over the place of the ark and overshadowed the ark and its carrying poles.
1KGS|8|8|These poles were so long that their ends could be seen from the Holy Place in front of the inner sanctuary, but not from outside the Holy Place; and they are still there today.
1KGS|8|9|There was nothing in the ark except the two stone tablets that Moses had placed in it at Horeb, where the LORD made a covenant with the Israelites after they came out of Egypt.
1KGS|8|10|When the priests withdrew from the Holy Place, the cloud filled the temple of the LORD.
1KGS|8|11|And the priests could not perform their service because of the cloud, for the glory of the LORD filled his temple.
1KGS|8|12|Then Solomon said, "The LORD has said that he would dwell in a dark cloud;
1KGS|8|13|I have indeed built a magnificent temple for you, a place for you to dwell forever."
1KGS|8|14|While the whole assembly of Israel was standing there, the king turned around and blessed them.
1KGS|8|15|Then he said: "Praise be to the LORD, the God of Israel, who with his own hand has fulfilled what he promised with his own mouth to my father David. For he said,
1KGS|8|16|'Since the day I brought my people Israel out of Egypt, I have not chosen a city in any tribe of Israel to have a temple built for my Name to be there, but I have chosen David to rule my people Israel.'
1KGS|8|17|"My father David had it in his heart to build a temple for the Name of the LORD, the God of Israel.
1KGS|8|18|But the LORD said to my father David, 'Because it was in your heart to build a temple for my Name, you did well to have this in your heart.
1KGS|8|19|Nevertheless, you are not the one to build the temple, but your son, who is your own flesh and blood-he is the one who will build the temple for my Name.'
1KGS|8|20|"The LORD has kept the promise he made: I have succeeded David my father and now I sit on the throne of Israel, just as the LORD promised, and I have built the temple for the Name of the LORD, the God of Israel.
1KGS|8|21|I have provided a place there for the ark, in which is the covenant of the LORD that he made with our fathers when he brought them out of Egypt."
1KGS|8|22|Then Solomon stood before the altar of the LORD in front of the whole assembly of Israel, spread out his hands toward heaven
1KGS|8|23|and said: "O LORD, God of Israel, there is no God like you in heaven above or on earth below-you who keep your covenant of love with your servants who continue wholeheartedly in your way.
1KGS|8|24|You have kept your promise to your servant David my father; with your mouth you have promised and with your hand you have fulfilled it-as it is today.
1KGS|8|25|"Now LORD, God of Israel, keep for your servant David my father the promises you made to him when you said, 'You shall never fail to have a man to sit before me on the throne of Israel, if only your sons are careful in all they do to walk before me as you have done.'
1KGS|8|26|And now, O God of Israel, let your word that you promised your servant David my father come true.
1KGS|8|27|"But will God really dwell on earth? The heavens, even the highest heaven, cannot contain you. How much less this temple I have built!
1KGS|8|28|Yet give attention to your servant's prayer and his plea for mercy, O LORD my God. Hear the cry and the prayer that your servant is praying in your presence this day.
1KGS|8|29|May your eyes be open toward this temple night and day, this place of which you said, 'My Name shall be there,' so that you will hear the prayer your servant prays toward this place.
1KGS|8|30|Hear the supplication of your servant and of your people Israel when they pray toward this place. Hear from heaven, your dwelling place, and when you hear, forgive.
1KGS|8|31|"When a man wrongs his neighbor and is required to take an oath and he comes and swears the oath before your altar in this temple,
1KGS|8|32|then hear from heaven and act. Judge between your servants, condemning the guilty and bringing down on his own head what he has done. Declare the innocent not guilty, and so establish his innocence.
1KGS|8|33|"When your people Israel have been defeated by an enemy because they have sinned against you, and when they turn back to you and confess your name, praying and making supplication to you in this temple,
1KGS|8|34|then hear from heaven and forgive the sin of your people Israel and bring them back to the land you gave to their fathers.
1KGS|8|35|"When the heavens are shut up and there is no rain because your people have sinned against you, and when they pray toward this place and confess your name and turn from their sin because you have afflicted them,
1KGS|8|36|then hear from heaven and forgive the sin of your servants, your people Israel. Teach them the right way to live, and send rain on the land you gave your people for an inheritance.
1KGS|8|37|"When famine or plague comes to the land, or blight or mildew, locusts or grasshoppers, or when an enemy besieges them in any of their cities, whatever disaster or disease may come,
1KGS|8|38|and when a prayer or plea is made by any of your people Israel-each one aware of the afflictions of his own heart, and spreading out his hands toward this temple-
1KGS|8|39|then hear from heaven, your dwelling place. Forgive and act; deal with each man according to all he does, since you know his heart (for you alone know the hearts of all men),
1KGS|8|40|so that they will fear you all the time they live in the land you gave our fathers.
1KGS|8|41|"As for the foreigner who does not belong to your people Israel but has come from a distant land because of your name-
1KGS|8|42|for men will hear of your great name and your mighty hand and your outstretched arm-when he comes and prays toward this temple,
1KGS|8|43|then hear from heaven, your dwelling place, and do whatever the foreigner asks of you, so that all the peoples of the earth may know your name and fear you, as do your own people Israel, and may know that this house I have built bears your Name.
1KGS|8|44|"When your people go to war against their enemies, wherever you send them, and when they pray to the LORD toward the city you have chosen and the temple I have built for your Name,
1KGS|8|45|then hear from heaven their prayer and their plea, and uphold their cause.
1KGS|8|46|"When they sin against you-for there is no one who does not sin-and you become angry with them and give them over to the enemy, who takes them captive to his own land, far away or near;
1KGS|8|47|and if they have a change of heart in the land where they are held captive, and repent and plead with you in the land of their conquerors and say, 'We have sinned, we have done wrong, we have acted wickedly';
1KGS|8|48|and if they turn back to you with all their heart and soul in the land of their enemies who took them captive, and pray to you toward the land you gave their fathers, toward the city you have chosen and the temple I have built for your Name;
1KGS|8|49|then from heaven, your dwelling place, hear their prayer and their plea, and uphold their cause.
1KGS|8|50|And forgive your people, who have sinned against you; forgive all the offenses they have committed against you, and cause their conquerors to show them mercy;
1KGS|8|51|for they are your people and your inheritance, whom you brought out of Egypt, out of that iron-smelting furnace.
1KGS|8|52|"May your eyes be open to your servant's plea and to the plea of your people Israel, and may you listen to them whenever they cry out to you.
1KGS|8|53|For you singled them out from all the nations of the world to be your own inheritance, just as you declared through your servant Moses when you, O Sovereign LORD, brought our fathers out of Egypt."
1KGS|8|54|When Solomon had finished all these prayers and supplications to the LORD, he rose from before the altar of the LORD, where he had been kneeling with his hands spread out toward heaven.
1KGS|8|55|He stood and blessed the whole assembly of Israel in a loud voice, saying:
1KGS|8|56|"Praise be to the LORD, who has given rest to his people Israel just as he promised. Not one word has failed of all the good promises he gave through his servant Moses.
1KGS|8|57|May the LORD our God be with us as he was with our fathers; may he never leave us nor forsake us.
1KGS|8|58|May he turn our hearts to him, to walk in all his ways and to keep the commands, decrees and regulations he gave our fathers.
1KGS|8|59|And may these words of mine, which I have prayed before the LORD, be near to the LORD our God day and night, that he may uphold the cause of his servant and the cause of his people Israel according to each day's need,
1KGS|8|60|so that all the peoples of the earth may know that the LORD is God and that there is no other.
1KGS|8|61|But your hearts must be fully committed to the LORD our God, to live by his decrees and obey his commands, as at this time."
1KGS|8|62|Then the king and all Israel with him offered sacrifices before the LORD.
1KGS|8|63|Solomon offered a sacrifice of fellowship offerings to the LORD: twenty-two thousand cattle and a hundred and twenty thousand sheep and goats. So the king and all the Israelites dedicated the temple of the LORD.
1KGS|8|64|On that same day the king consecrated the middle part of the courtyard in front of the temple of the LORD, and there he offered burnt offerings, grain offerings and the fat of the fellowship offerings, because the bronze altar before the LORD was too small to hold the burnt offerings, the grain offerings and the fat of the fellowship offerings.
1KGS|8|65|So Solomon observed the festival at that time, and all Israel with him-a vast assembly, people from Lebo Hamath to the Wadi of Egypt. They celebrated it before the LORD our God for seven days and seven days more, fourteen days in all.
1KGS|8|66|On the following day he sent the people away. They blessed the king and then went home, joyful and glad in heart for all the good things the LORD had done for his servant David and his people Israel.
1KGS|9|1|When Solomon had finished building the temple of the LORD and the royal palace, and had achieved all he had desired to do,
1KGS|9|2|the LORD appeared to him a second time, as he had appeared to him at Gibeon.
1KGS|9|3|The LORD said to him: "I have heard the prayer and plea you have made before me; I have consecrated this temple, which you have built, by putting my Name there forever. My eyes and my heart will always be there.
1KGS|9|4|"As for you, if you walk before me in integrity of heart and uprightness, as David your father did, and do all I command and observe my decrees and laws,
1KGS|9|5|I will establish your royal throne over Israel forever, as I promised David your father when I said, 'You shall never fail to have a man on the throne of Israel.'
1KGS|9|6|"But if you or your sons turn away from me and do not observe the commands and decrees I have given you and go off to serve other gods and worship them,
1KGS|9|7|then I will cut off Israel from the land I have given them and will reject this temple I have consecrated for my Name. Israel will then become a byword and an object of ridicule among all peoples.
1KGS|9|8|And though this temple is now imposing, all who pass by will be appalled and will scoff and say, 'Why has the LORD done such a thing to this land and to this temple?'
1KGS|9|9|People will answer, 'Because they have forsaken the LORD their God, who brought their fathers out of Egypt, and have embraced other gods, worshiping and serving them-that is why the LORD brought all this disaster on them.'"
1KGS|9|10|At the end of twenty years, during which Solomon built these two buildings-the temple of the LORD and the royal palace-
1KGS|9|11|King Solomon gave twenty towns in Galilee to Hiram king of Tyre, because Hiram had supplied him with all the cedar and pine and gold he wanted.
1KGS|9|12|But when Hiram went from Tyre to see the towns that Solomon had given him, he was not pleased with them.
1KGS|9|13|"What kind of towns are these you have given me, my brother?" he asked. And he called them the Land of Cabul, a name they have to this day.
1KGS|9|14|Now Hiram had sent to the king 120 talents of gold.
1KGS|9|15|Here is the account of the forced labor King Solomon conscripted to build the LORD's temple, his own palace, the supporting terraces, the wall of Jerusalem, and Hazor, Megiddo and Gezer.
1KGS|9|16|(Pharaoh king of Egypt had attacked and captured Gezer. He had set it on fire. He killed its Canaanite inhabitants and then gave it as a wedding gift to his daughter, Solomon's wife.
1KGS|9|17|And Solomon rebuilt Gezer.) He built up Lower Beth Horon,
1KGS|9|18|Baalath, and Tadmor in the desert, within his land,
1KGS|9|19|as well as all his store cities and the towns for his chariots and for his horses -whatever he desired to build in Jerusalem, in Lebanon and throughout all the territory he ruled.
1KGS|9|20|All the people left from the Amorites, Hittites, Perizzites, Hivites and Jebusites (these peoples were not Israelites),
1KGS|9|21|that is, their descendants remaining in the land, whom the Israelites could not exterminate -these Solomon conscripted for his slave labor force, as it is to this day.
1KGS|9|22|But Solomon did not make slaves of any of the Israelites; they were his fighting men, his government officials, his officers, his captains, and the commanders of his chariots and charioteers.
1KGS|9|23|They were also the chief officials in charge of Solomon's projects-550 officials supervising the men who did the work.
1KGS|9|24|After Pharaoh's daughter had come up from the City of David to the palace Solomon had built for her, he constructed the supporting terraces.
1KGS|9|25|Three times a year Solomon sacrificed burnt offerings and fellowship offerings on the altar he had built for the LORD, burning incense before the LORD along with them, and so fulfilled the temple obligations.
1KGS|9|26|King Solomon also built ships at Ezion Geber, which is near Elath in Edom, on the shore of the Red Sea.
1KGS|9|27|And Hiram sent his men-sailors who knew the sea-to serve in the fleet with Solomon's men.
1KGS|9|28|They sailed to Ophir and brought back 420 talents of gold, which they delivered to King Solomon.
1KGS|10|1|When the queen of Sheba heard about the fame of Solomon and his relation to the name of the LORD, she came to test him with hard questions.
1KGS|10|2|Arriving at Jerusalem with a very great caravan-with camels carrying spices, large quantities of gold, and precious stones-she came to Solomon and talked with him about all that she had on her mind.
1KGS|10|3|Solomon answered all her questions; nothing was too hard for the king to explain to her.
1KGS|10|4|When the queen of Sheba saw all the wisdom of Solomon and the palace he had built,
1KGS|10|5|the food on his table, the seating of his officials, the attending servants in their robes, his cupbearers, and the burnt offerings he made at the temple of the LORD, she was overwhelmed.
1KGS|10|6|She said to the king, "The report I heard in my own country about your achievements and your wisdom is true.
1KGS|10|7|But I did not believe these things until I came and saw with my own eyes. Indeed, not even half was told me; in wisdom and wealth you have far exceeded the report I heard.
1KGS|10|8|How happy your men must be! How happy your officials, who continually stand before you and hear your wisdom!
1KGS|10|9|Praise be to the LORD your God, who has delighted in you and placed you on the throne of Israel. Because of the LORD's eternal love for Israel, he has made you king, to maintain justice and righteousness."
1KGS|10|10|And she gave the king 120 talents of gold, large quantities of spices, and precious stones. Never again were so many spices brought in as those the queen of Sheba gave to King Solomon.
1KGS|10|11|(Hiram's ships brought gold from Ophir; and from there they brought great cargoes of almugwood and precious stones.
1KGS|10|12|The king used the almugwood to make supports for the temple of the LORD and for the royal palace, and to make harps and lyres for the musicians. So much almugwood has never been imported or seen since that day.)
1KGS|10|13|King Solomon gave the queen of Sheba all she desired and asked for, besides what he had given her out of his royal bounty. Then she left and returned with her retinue to her own country.
1KGS|10|14|The weight of the gold that Solomon received yearly was 666 talents,
1KGS|10|15|not including the revenues from merchants and traders and from all the Arabian kings and the governors of the land.
1KGS|10|16|King Solomon made two hundred large shields of hammered gold; six hundred bekas of gold went into each shield.
1KGS|10|17|He also made three hundred small shields of hammered gold, with three minas of gold in each shield. The king put them in the Palace of the Forest of Lebanon.
1KGS|10|18|Then the king made a great throne inlaid with ivory and overlaid with fine gold.
1KGS|10|19|The throne had six steps, and its back had a rounded top. On both sides of the seat were armrests, with a lion standing beside each of them.
1KGS|10|20|Twelve lions stood on the six steps, one at either end of each step. Nothing like it had ever been made for any other kingdom.
1KGS|10|21|All King Solomon's goblets were gold, and all the household articles in the Palace of the Forest of Lebanon were pure gold. Nothing was made of silver, because silver was considered of little value in Solomon's days.
1KGS|10|22|The king had a fleet of trading ships at sea along with the ships of Hiram. Once every three years it returned, carrying gold, silver and ivory, and apes and baboons.
1KGS|10|23|King Solomon was greater in riches and wisdom than all the other kings of the earth.
1KGS|10|24|The whole world sought audience with Solomon to hear the wisdom God had put in his heart.
1KGS|10|25|Year after year, everyone who came brought a gift-articles of silver and gold, robes, weapons and spices, and horses and mules.
1KGS|10|26|Solomon accumulated chariots and horses; he had fourteen hundred chariots and twelve thousand horses, which he kept in the chariot cities and also with him in Jerusalem.
1KGS|10|27|The king made silver as common in Jerusalem as stones, and cedar as plentiful as sycamore-fig trees in the foothills.
1KGS|10|28|Solomon's horses were imported from Egypt and from Kue - the royal merchants purchased them from Kue.
1KGS|10|29|They imported a chariot from Egypt for six hundred shekels of silver, and a horse for a hundred and fifty. They also exported them to all the kings of the Hittites and of the Arameans.
1KGS|11|1|King Solomon, however, loved many foreign women besides Pharaoh's daughter-Moabites, Ammonites, Edomites, Sidonians and Hittites.
1KGS|11|2|They were from nations about which the LORD had told the Israelites, "You must not intermarry with them, because they will surely turn your hearts after their gods." Nevertheless, Solomon held fast to them in love.
1KGS|11|3|He had seven hundred wives of royal birth and three hundred concubines, and his wives led him astray.
1KGS|11|4|As Solomon grew old, his wives turned his heart after other gods, and his heart was not fully devoted to the LORD his God, as the heart of David his father had been.
1KGS|11|5|He followed Ashtoreth the goddess of the Sidonians, and Molech the detestable god of the Ammonites.
1KGS|11|6|So Solomon did evil in the eyes of the LORD; he did not follow the LORD completely, as David his father had done.
1KGS|11|7|On a hill east of Jerusalem, Solomon built a high place for Chemosh the detestable god of Moab, and for Molech the detestable god of the Ammonites.
1KGS|11|8|He did the same for all his foreign wives, who burned incense and offered sacrifices to their gods.
1KGS|11|9|The LORD became angry with Solomon because his heart had turned away from the LORD, the God of Israel, who had appeared to him twice.
1KGS|11|10|Although he had forbidden Solomon to follow other gods, Solomon did not keep the LORD's command.
1KGS|11|11|So the LORD said to Solomon, "Since this is your attitude and you have not kept my covenant and my decrees, which I commanded you, I will most certainly tear the kingdom away from you and give it to one of your subordinates.
1KGS|11|12|Nevertheless, for the sake of David your father, I will not do it during your lifetime. I will tear it out of the hand of your son.
1KGS|11|13|Yet I will not tear the whole kingdom from him, but will give him one tribe for the sake of David my servant and for the sake of Jerusalem, which I have chosen."
1KGS|11|14|Then the LORD raised up against Solomon an adversary, Hadad the Edomite, from the royal line of Edom.
1KGS|11|15|Earlier when David was fighting with Edom, Joab the commander of the army, who had gone up to bury the dead, had struck down all the men in Edom.
1KGS|11|16|Joab and all the Israelites stayed there for six months, until they had destroyed all the men in Edom.
1KGS|11|17|But Hadad, still only a boy, fled to Egypt with some Edomite officials who had served his father.
1KGS|11|18|They set out from Midian and went to Paran. Then taking men from Paran with them, they went to Egypt, to Pharaoh king of Egypt, who gave Hadad a house and land and provided him with food.
1KGS|11|19|Pharaoh was so pleased with Hadad that he gave him a sister of his own wife, Queen Tahpenes, in marriage.
1KGS|11|20|The sister of Tahpenes bore him a son named Genubath, whom Tahpenes brought up in the royal palace. There Genubath lived with Pharaoh's own children.
1KGS|11|21|While he was in Egypt, Hadad heard that David rested with his fathers and that Joab the commander of the army was also dead. Then Hadad said to Pharaoh, "Let me go, that I may return to my own country."
1KGS|11|22|"What have you lacked here that you want to go back to your own country?" Pharaoh asked. "Nothing," Hadad replied, "but do let me go!"
1KGS|11|23|And God raised up against Solomon another adversary, Rezon son of Eliada, who had fled from his master, Hadadezer king of Zobah.
1KGS|11|24|He gathered men around him and became the leader of a band of rebels when David destroyed the forces of Zobah; the rebels went to Damascus, where they settled and took control.
1KGS|11|25|Rezon was Israel's adversary as long as Solomon lived, adding to the trouble caused by Hadad. So Rezon ruled in Aram and was hostile toward Israel.
1KGS|11|26|Also, Jeroboam son of Nebat rebelled against the king. He was one of Solomon's officials, an Ephraimite from Zeredah, and his mother was a widow named Zeruah.
1KGS|11|27|Here is the account of how he rebelled against the king: Solomon had built the supporting terraces and had filled in the gap in the wall of the city of David his father.
1KGS|11|28|Now Jeroboam was a man of standing, and when Solomon saw how well the young man did his work, he put him in charge of the whole labor force of the house of Joseph.
1KGS|11|29|About that time Jeroboam was going out of Jerusalem, and Ahijah the prophet of Shiloh met him on the way, wearing a new cloak. The two of them were alone out in the country,
1KGS|11|30|and Ahijah took hold of the new cloak he was wearing and tore it into twelve pieces.
1KGS|11|31|Then he said to Jeroboam, "Take ten pieces for yourself, for this is what the LORD, the God of Israel, says: 'See, I am going to tear the kingdom out of Solomon's hand and give you ten tribes.
1KGS|11|32|But for the sake of my servant David and the city of Jerusalem, which I have chosen out of all the tribes of Israel, he will have one tribe.
1KGS|11|33|I will do this because they have forsaken me and worshiped Ashtoreth the goddess of the Sidonians, Chemosh the god of the Moabites, and Molech the god of the Ammonites, and have not walked in my ways, nor done what is right in my eyes, nor kept my statutes and laws as David, Solomon's father, did.
1KGS|11|34|"'But I will not take the whole kingdom out of Solomon's hand; I have made him ruler all the days of his life for the sake of David my servant, whom I chose and who observed my commands and statutes.
1KGS|11|35|I will take the kingdom from his son's hands and give you ten tribes.
1KGS|11|36|I will give one tribe to his son so that David my servant may always have a lamp before me in Jerusalem, the city where I chose to put my Name.
1KGS|11|37|However, as for you, I will take you, and you will rule over all that your heart desires; you will be king over Israel.
1KGS|11|38|If you do whatever I command you and walk in my ways and do what is right in my eyes by keeping my statutes and commands, as David my servant did, I will be with you. I will build you a dynasty as enduring as the one I built for David and will give Israel to you.
1KGS|11|39|I will humble David's descendants because of this, but not forever.'"
1KGS|11|40|Solomon tried to kill Jeroboam, but Jeroboam fled to Egypt, to Shishak the king, and stayed there until Solomon's death.
1KGS|11|41|As for the other events of Solomon's reign-all he did and the wisdom he displayed-are they not written in the book of the annals of Solomon?
1KGS|11|42|Solomon reigned in Jerusalem over all Israel forty years.
1KGS|11|43|Then he rested with his fathers and was buried in the city of David his father. And Rehoboam his son succeeded him as king.
1KGS|12|1|Rehoboam went to Shechem, for all the Israelites had gone there to make him king.
1KGS|12|2|When Jeroboam son of Nebat heard this (he was still in Egypt, where he had fled from King Solomon), he returned from Egypt.
1KGS|12|3|So they sent for Jeroboam, and he and the whole assembly of Israel went to Rehoboam and said to him:
1KGS|12|4|"Your father put a heavy yoke on us, but now lighten the harsh labor and the heavy yoke he put on us, and we will serve you."
1KGS|12|5|Rehoboam answered, "Go away for three days and then come back to me." So the people went away.
1KGS|12|6|Then King Rehoboam consulted the elders who had served his father Solomon during his lifetime. "How would you advise me to answer these people?" he asked.
1KGS|12|7|They replied, "If today you will be a servant to these people and serve them and give them a favorable answer, they will always be your servants."
1KGS|12|8|But Rehoboam rejected the advice the elders gave him and consulted the young men who had grown up with him and were serving him.
1KGS|12|9|He asked them, "What is your advice? How should we answer these people who say to me, 'Lighten the yoke your father put on us'?"
1KGS|12|10|The young men who had grown up with him replied, "Tell these people who have said to you, 'Your father put a heavy yoke on us, but make our yoke lighter'-tell them, 'My little finger is thicker than my father's waist.
1KGS|12|11|My father laid on you a heavy yoke; I will make it even heavier. My father scourged you with whips; I will scourge you with scorpions.'"
1KGS|12|12|Three days later Jeroboam and all the people returned to Rehoboam, as the king had said, "Come back to me in three days."
1KGS|12|13|The king answered the people harshly. Rejecting the advice given him by the elders,
1KGS|12|14|he followed the advice of the young men and said, "My father made your yoke heavy; I will make it even heavier. My father scourged you with whips; I will scourge you with scorpions."
1KGS|12|15|So the king did not listen to the people, for this turn of events was from the LORD, to fulfill the word the LORD had spoken to Jeroboam son of Nebat through Ahijah the Shilonite.
1KGS|12|16|When all Israel saw that the king refused to listen to them, they answered the king: "What share do we have in David, what part in Jesse's son? To your tents, O Israel! Look after your own house, O David!" So the Israelites went home.
1KGS|12|17|But as for the Israelites who were living in the towns of Judah, Rehoboam still ruled over them.
1KGS|12|18|King Rehoboam sent out Adoniram, who was in charge of forced labor, but all Israel stoned him to death. King Rehoboam, however, managed to get into his chariot and escape to Jerusalem.
1KGS|12|19|So Israel has been in rebellion against the house of David to this day.
1KGS|12|20|When all the Israelites heard that Jeroboam had returned, they sent and called him to the assembly and made him king over all Israel. Only the tribe of Judah remained loyal to the house of David.
1KGS|12|21|When Rehoboam arrived in Jerusalem, he mustered the whole house of Judah and the tribe of Benjamin-a hundred and eighty thousand fighting men-to make war against the house of Israel and to regain the kingdom for Rehoboam son of Solomon.
1KGS|12|22|But this word of God came to Shemaiah the man of God:
1KGS|12|23|"Say to Rehoboam son of Solomon king of Judah, to the whole house of Judah and Benjamin, and to the rest of the people,
1KGS|12|24|'This is what the LORD says: Do not go up to fight against your brothers, the Israelites. Go home, every one of you, for this is my doing.'" So they obeyed the word of the LORD and went home again, as the LORD had ordered.
1KGS|12|25|Then Jeroboam fortified Shechem in the hill country of Ephraim and lived there. From there he went out and built up Peniel.
1KGS|12|26|Jeroboam thought to himself, "The kingdom will now likely revert to the house of David.
1KGS|12|27|If these people go up to offer sacrifices at the temple of the LORD in Jerusalem, they will again give their allegiance to their lord, Rehoboam king of Judah. They will kill me and return to King Rehoboam."
1KGS|12|28|After seeking advice, the king made two golden calves. He said to the people, "It is too much for you to go up to Jerusalem. Here are your gods, O Israel, who brought you up out of Egypt."
1KGS|12|29|One he set up in Bethel, and the other in Dan.
1KGS|12|30|And this thing became a sin; the people went even as far as Dan to worship the one there.
1KGS|12|31|Jeroboam built shrines on high places and appointed priests from all sorts of people, even though they were not Levites.
1KGS|12|32|He instituted a festival on the fifteenth day of the eighth month, like the festival held in Judah, and offered sacrifices on the altar. This he did in Bethel, sacrificing to the calves he had made. And at Bethel he also installed priests at the high places he had made.
1KGS|12|33|On the fifteenth day of the eighth month, a month of his own choosing, he offered sacrifices on the altar he had built at Bethel. So he instituted the festival for the Israelites and went up to the altar to make offerings.
1KGS|13|1|By the word of the LORD a man of God came from Judah to Bethel, as Jeroboam was standing by the altar to make an offering.
1KGS|13|2|He cried out against the altar by the word of the LORD: "O altar, altar! This is what the LORD says: 'A son named Josiah will be born to the house of David. On you he will sacrifice the priests of the high places who now make offerings here, and human bones will be burned on you.'"
1KGS|13|3|That same day the man of God gave a sign: "This is the sign the LORD has declared: The altar will be split apart and the ashes on it will be poured out."
1KGS|13|4|When King Jeroboam heard what the man of God cried out against the altar at Bethel, he stretched out his hand from the altar and said, "Seize him!" But the hand he stretched out toward the man shriveled up, so that he could not pull it back.
1KGS|13|5|Also, the altar was split apart and its ashes poured out according to the sign given by the man of God by the word of the LORD.
1KGS|13|6|Then the king said to the man of God, "Intercede with the LORD your God and pray for me that my hand may be restored." So the man of God interceded with the LORD, and the king's hand was restored and became as it was before.
1KGS|13|7|The king said to the man of God, "Come home with me and have something to eat, and I will give you a gift."
1KGS|13|8|But the man of God answered the king, "Even if you were to give me half your possessions, I would not go with you, nor would I eat bread or drink water here.
1KGS|13|9|For I was commanded by the word of the LORD: 'You must not eat bread or drink water or return by the way you came.'"
1KGS|13|10|So he took another road and did not return by the way he had come to Bethel.
1KGS|13|11|Now there was a certain old prophet living in Bethel, whose sons came and told him all that the man of God had done there that day. They also told their father what he had said to the king.
1KGS|13|12|Their father asked them, "Which way did he go?" And his sons showed him which road the man of God from Judah had taken.
1KGS|13|13|So he said to his sons, "Saddle the donkey for me." And when they had saddled the donkey for him, he mounted it
1KGS|13|14|and rode after the man of God. He found him sitting under an oak tree and asked, "Are you the man of God who came from Judah?I am," he replied.
1KGS|13|15|So the prophet said to him, "Come home with me and eat."
1KGS|13|16|The man of God said, "I cannot turn back and go with you, nor can I eat bread or drink water with you in this place.
1KGS|13|17|I have been told by the word of the LORD: 'You must not eat bread or drink water there or return by the way you came.'"
1KGS|13|18|The old prophet answered, "I too am a prophet, as you are. And an angel said to me by the word of the LORD: 'Bring him back with you to your house so that he may eat bread and drink water.'" (But he was lying to him.)
1KGS|13|19|So the man of God returned with him and ate and drank in his house.
1KGS|13|20|While they were sitting at the table, the word of the LORD came to the old prophet who had brought him back.
1KGS|13|21|He cried out to the man of God who had come from Judah, "This is what the LORD says: 'You have defied the word of the LORD and have not kept the command the LORD your God gave you.
1KGS|13|22|You came back and ate bread and drank water in the place where he told you not to eat or drink. Therefore your body will not be buried in the tomb of your fathers.'"
1KGS|13|23|When the man of God had finished eating and drinking, the prophet who had brought him back saddled his donkey for him.
1KGS|13|24|As he went on his way, a lion met him on the road and killed him, and his body was thrown down on the road, with both the donkey and the lion standing beside it.
1KGS|13|25|Some people who passed by saw the body thrown down there, with the lion standing beside the body, and they went and reported it in the city where the old prophet lived.
1KGS|13|26|When the prophet who had brought him back from his journey heard of it, he said, "It is the man of God who defied the word of the LORD. The LORD has given him over to the lion, which has mauled him and killed him, as the word of the LORD had warned him."
1KGS|13|27|The prophet said to his sons, "Saddle the donkey for me," and they did so.
1KGS|13|28|Then he went out and found the body thrown down on the road, with the donkey and the lion standing beside it. The lion had neither eaten the body nor mauled the donkey.
1KGS|13|29|So the prophet picked up the body of the man of God, laid it on the donkey, and brought it back to his own city to mourn for him and bury him.
1KGS|13|30|Then he laid the body in his own tomb, and they mourned over him and said, "Oh, my brother!"
1KGS|13|31|After burying him, he said to his sons, "When I die, bury me in the grave where the man of God is buried; lay my bones beside his bones.
1KGS|13|32|For the message he declared by the word of the LORD against the altar in Bethel and against all the shrines on the high places in the towns of Samaria will certainly come true."
1KGS|13|33|Even after this, Jeroboam did not change his evil ways, but once more appointed priests for the high places from all sorts of people. Anyone who wanted to become a priest he consecrated for the high places.
1KGS|13|34|This was the sin of the house of Jeroboam that led to its downfall and to its destruction from the face of the earth.
1KGS|14|1|At that time Abijah son of Jeroboam became ill,
1KGS|14|2|and Jeroboam said to his wife, "Go, disguise yourself, so you won't be recognized as the wife of Jeroboam. Then go to Shiloh. Ahijah the prophet is there-the one who told me I would be king over this people.
1KGS|14|3|Take ten loaves of bread with you, some cakes and a jar of honey, and go to him. He will tell you what will happen to the boy."
1KGS|14|4|So Jeroboam's wife did what he said and went to Ahijah's house in Shiloh. Now Ahijah could not see; his sight was gone because of his age.
1KGS|14|5|But the LORD had told Ahijah, "Jeroboam's wife is coming to ask you about her son, for he is ill, and you are to give her such and such an answer. When she arrives, she will pretend to be someone else."
1KGS|14|6|So when Ahijah heard the sound of her footsteps at the door, he said, "Come in, wife of Jeroboam. Why this pretense? I have been sent to you with bad news.
1KGS|14|7|Go, tell Jeroboam that this is what the LORD, the God of Israel, says: 'I raised you up from among the people and made you a leader over my people Israel.
1KGS|14|8|I tore the kingdom away from the house of David and gave it to you, but you have not been like my servant David, who kept my commands and followed me with all his heart, doing only what was right in my eyes.
1KGS|14|9|You have done more evil than all who lived before you. You have made for yourself other gods, idols made of metal; you have provoked me to anger and thrust me behind your back.
1KGS|14|10|"'Because of this, I am going to bring disaster on the house of Jeroboam. I will cut off from Jeroboam every last male in Israel-slave or free. I will burn up the house of Jeroboam as one burns dung, until it is all gone.
1KGS|14|11|Dogs will eat those belonging to Jeroboam who die in the city, and the birds of the air will feed on those who die in the country. The LORD has spoken!'
1KGS|14|12|"As for you, go back home. When you set foot in your city, the boy will die.
1KGS|14|13|All Israel will mourn for him and bury him. He is the only one belonging to Jeroboam who will be buried, because he is the only one in the house of Jeroboam in whom the LORD, the God of Israel, has found anything good.
1KGS|14|14|"The LORD will raise up for himself a king over Israel who will cut off the family of Jeroboam. This is the day! What? Yes, even now.
1KGS|14|15|And the LORD will strike Israel, so that it will be like a reed swaying in the water. He will uproot Israel from this good land that he gave to their forefathers and scatter them beyond the River, because they provoked the LORD to anger by making Asherah poles.
1KGS|14|16|And he will give Israel up because of the sins Jeroboam has committed and has caused Israel to commit."
1KGS|14|17|Then Jeroboam's wife got up and left and went to Tirzah. As soon as she stepped over the threshold of the house, the boy died.
1KGS|14|18|They buried him, and all Israel mourned for him, as the LORD had said through his servant the prophet Ahijah.
1KGS|14|19|The other events of Jeroboam's reign, his wars and how he ruled, are written in the book of the annals of the kings of Israel.
1KGS|14|20|He reigned for twenty-two years and then rested with his fathers. And Nadab his son succeeded him as king.
1KGS|14|21|Rehoboam son of Solomon was king in Judah. He was forty-one years old when he became king, and he reigned seventeen years in Jerusalem, the city the LORD had chosen out of all the tribes of Israel in which to put his Name. His mother's name was Naamah; she was an Ammonite.
1KGS|14|22|Judah did evil in the eyes of the LORD. By the sins they committed they stirred up his jealous anger more than their fathers had done.
1KGS|14|23|They also set up for themselves high places, sacred stones and Asherah poles on every high hill and under every spreading tree.
1KGS|14|24|There were even male shrine prostitutes in the land; the people engaged in all the detestable practices of the nations the LORD had driven out before the Israelites.
1KGS|14|25|In the fifth year of King Rehoboam, Shishak king of Egypt attacked Jerusalem.
1KGS|14|26|He carried off the treasures of the temple of the LORD and the treasures of the royal palace. He took everything, including all the gold shields Solomon had made.
1KGS|14|27|So King Rehoboam made bronze shields to replace them and assigned these to the commanders of the guard on duty at the entrance to the royal palace.
1KGS|14|28|Whenever the king went to the LORD's temple, the guards bore the shields, and afterward they returned them to the guardroom.
1KGS|14|29|As for the other events of Rehoboam's reign, and all he did, are they not written in the book of the annals of the kings of Judah?
1KGS|14|30|There was continual warfare between Rehoboam and Jeroboam.
1KGS|14|31|And Rehoboam rested with his fathers and was buried with them in the City of David. His mother's name was Naamah; she was an Ammonite. And Abijah his son succeeded him as king.
1KGS|15|1|In the eighteenth year of the reign of Jeroboam son of Nebat, Abijah became king of Judah,
1KGS|15|2|and he reigned in Jerusalem three years. His mother's name was Maacah daughter of Abishalom.
1KGS|15|3|He committed all the sins his father had done before him; his heart was not fully devoted to the LORD his God, as the heart of David his forefather had been.
1KGS|15|4|Nevertheless, for David's sake the LORD his God gave him a lamp in Jerusalem by raising up a son to succeed him and by making Jerusalem strong.
1KGS|15|5|For David had done what was right in the eyes of the LORD and had not failed to keep any of the LORD's commands all the days of his life-except in the case of Uriah the Hittite.
1KGS|15|6|There was war between Rehoboam and Jeroboam throughout Abijah's lifetime.
1KGS|15|7|As for the other events of Abijah's reign, and all he did, are they not written in the book of the annals of the kings of Judah? There was war between Abijah and Jeroboam.
1KGS|15|8|And Abijah rested with his fathers and was buried in the City of David. And Asa his son succeeded him as king.
1KGS|15|9|In the twentieth year of Jeroboam king of Israel, Asa became king of Judah,
1KGS|15|10|and he reigned in Jerusalem forty-one years. His grandmother's name was Maacah daughter of Abishalom.
1KGS|15|11|Asa did what was right in the eyes of the LORD, as his father David had done.
1KGS|15|12|He expelled the male shrine prostitutes from the land and got rid of all the idols his fathers had made.
1KGS|15|13|He even deposed his grandmother Maacah from her position as queen mother, because she had made a repulsive Asherah pole. Asa cut the pole down and burned it in the Kidron Valley.
1KGS|15|14|Although he did not remove the high places, Asa's heart was fully committed to the LORD all his life.
1KGS|15|15|He brought into the temple of the LORD the silver and gold and the articles that he and his father had dedicated.
1KGS|15|16|There was war between Asa and Baasha king of Israel throughout their reigns.
1KGS|15|17|Baasha king of Israel went up against Judah and fortified Ramah to prevent anyone from leaving or entering the territory of Asa king of Judah.
1KGS|15|18|Asa then took all the silver and gold that was left in the treasuries of the LORD's temple and of his own palace. He entrusted it to his officials and sent them to Ben-Hadad son of Tabrimmon, the son of Hezion, the king of Aram, who was ruling in Damascus.
1KGS|15|19|"Let there be a treaty between me and you," he said, "as there was between my father and your father. See, I am sending you a gift of silver and gold. Now break your treaty with Baasha king of Israel so he will withdraw from me."
1KGS|15|20|Ben-Hadad agreed with King Asa and sent the commanders of his forces against the towns of Israel. He conquered Ijon, Dan, Abel Beth Maacah and all Kinnereth in addition to Naphtali.
1KGS|15|21|When Baasha heard this, he stopped building Ramah and withdrew to Tirzah.
1KGS|15|22|Then King Asa issued an order to all Judah-no one was exempt-and they carried away from Ramah the stones and timber Baasha had been using there. With them King Asa built up Geba in Benjamin, and also Mizpah.
1KGS|15|23|As for all the other events of Asa's reign, all his achievements, all he did and the cities he built, are they not written in the book of the annals of the kings of Judah? In his old age, however, his feet became diseased.
1KGS|15|24|Then Asa rested with his fathers and was buried with them in the city of his father David. And Jehoshaphat his son succeeded him as king.
1KGS|15|25|Nadab son of Jeroboam became king of Israel in the second year of Asa king of Judah, and he reigned over Israel two years.
1KGS|15|26|He did evil in the eyes of the LORD, walking in the ways of his father and in his sin, which he had caused Israel to commit.
1KGS|15|27|Baasha son of Ahijah of the house of Issachar plotted against him, and he struck him down at Gibbethon, a Philistine town, while Nadab and all Israel were besieging it.
1KGS|15|28|Baasha killed Nadab in the third year of Asa king of Judah and succeeded him as king.
1KGS|15|29|As soon as he began to reign, he killed Jeroboam's whole family. He did not leave Jeroboam anyone that breathed, but destroyed them all, according to the word of the LORD given through his servant Ahijah the Shilonite-
1KGS|15|30|because of the sins Jeroboam had committed and had caused Israel to commit, and because he provoked the LORD, the God of Israel, to anger.
1KGS|15|31|As for the other events of Nadab's reign, and all he did, are they not written in the book of the annals of the kings of Israel?
1KGS|15|32|There was war between Asa and Baasha king of Israel throughout their reigns.
1KGS|15|33|In the third year of Asa king of Judah, Baasha son of Ahijah became king of all Israel in Tirzah, and he reigned twenty-four years.
1KGS|15|34|He did evil in the eyes of the LORD, walking in the ways of Jeroboam and in his sin, which he had caused Israel to commit.
1KGS|16|1|Then the word of the LORD came to Jehu son of Hanani against Baasha:
1KGS|16|2|"I lifted you up from the dust and made you leader of my people Israel, but you walked in the ways of Jeroboam and caused my people Israel to sin and to provoke me to anger by their sins.
1KGS|16|3|So I am about to consume Baasha and his house, and I will make your house like that of Jeroboam son of Nebat.
1KGS|16|4|Dogs will eat those belonging to Baasha who die in the city, and the birds of the air will feed on those who die in the country."
1KGS|16|5|As for the other events of Baasha's reign, what he did and his achievements, are they not written in the book of the annals of the kings of Israel?
1KGS|16|6|Baasha rested with his fathers and was buried in Tirzah. And Elah his son succeeded him as king.
1KGS|16|7|Moreover, the word of the LORD came through the prophet Jehu son of Hanani to Baasha and his house, because of all the evil he had done in the eyes of the LORD, provoking him to anger by the things he did, and becoming like the house of Jeroboam-and also because he destroyed it.
1KGS|16|8|In the twenty-sixth year of Asa king of Judah, Elah son of Baasha became king of Israel, and he reigned in Tirzah two years.
1KGS|16|9|Zimri, one of his officials, who had command of half his chariots, plotted against him. Elah was in Tirzah at the time, getting drunk in the home of Arza, the man in charge of the palace at Tirzah.
1KGS|16|10|Zimri came in, struck him down and killed him in the twenty-seventh year of Asa king of Judah. Then he succeeded him as king.
1KGS|16|11|As soon as he began to reign and was seated on the throne, he killed off Baasha's whole family. He did not spare a single male, whether relative or friend.
1KGS|16|12|So Zimri destroyed the whole family of Baasha, in accordance with the word of the LORD spoken against Baasha through the prophet Jehu-
1KGS|16|13|because of all the sins Baasha and his son Elah had committed and had caused Israel to commit, so that they provoked the LORD, the God of Israel, to anger by their worthless idols.
1KGS|16|14|As for the other events of Elah's reign, and all he did, are they not written in the book of the annals of the kings of Israel?
1KGS|16|15|In the twenty-seventh year of Asa king of Judah, Zimri reigned in Tirzah seven days. The army was encamped near Gibbethon, a Philistine town.
1KGS|16|16|When the Israelites in the camp heard that Zimri had plotted against the king and murdered him, they proclaimed Omri, the commander of the army, king over Israel that very day there in the camp.
1KGS|16|17|Then Omri and all the Israelites with him withdrew from Gibbethon and laid siege to Tirzah.
1KGS|16|18|When Zimri saw that the city was taken, he went into the citadel of the royal palace and set the palace on fire around him. So he died,
1KGS|16|19|because of the sins he had committed, doing evil in the eyes of the LORD and walking in the ways of Jeroboam and in the sin he had committed and had caused Israel to commit.
1KGS|16|20|As for the other events of Zimri's reign, and the rebellion he carried out, are they not written in the book of the annals of the kings of Israel?
1KGS|16|21|Then the people of Israel were split into two factions; half supported Tibni son of Ginath for king, and the other half supported Omri.
1KGS|16|22|But Omri's followers proved stronger than those of Tibni son of Ginath. So Tibni died and Omri became king.
1KGS|16|23|In the thirty-first year of Asa king of Judah, Omri became king of Israel, and he reigned twelve years, six of them in Tirzah.
1KGS|16|24|He bought the hill of Samaria from Shemer for two talents of silver and built a city on the hill, calling it Samaria, after Shemer, the name of the former owner of the hill.
1KGS|16|25|But Omri did evil in the eyes of the LORD and sinned more than all those before him.
1KGS|16|26|He walked in all the ways of Jeroboam son of Nebat and in his sin, which he had caused Israel to commit, so that they provoked the LORD, the God of Israel, to anger by their worthless idols.
1KGS|16|27|As for the other events of Omri's reign, what he did and the things he achieved, are they not written in the book of the annals of the kings of Israel?
1KGS|16|28|Omri rested with his fathers and was buried in Samaria. And Ahab his son succeeded him as king.
1KGS|16|29|In the thirty-eighth year of Asa king of Judah, Ahab son of Omri became king of Israel, and he reigned in Samaria over Israel twenty-two years.
1KGS|16|30|Ahab son of Omri did more evil in the eyes of the LORD than any of those before him.
1KGS|16|31|He not only considered it trivial to commit the sins of Jeroboam son of Nebat, but he also married Jezebel daughter of Ethbaal king of the Sidonians, and began to serve Baal and worship him.
1KGS|16|32|He set up an altar for Baal in the temple of Baal that he built in Samaria.
1KGS|16|33|Ahab also made an Asherah pole and did more to provoke the LORD, the God of Israel, to anger than did all the kings of Israel before him.
1KGS|16|34|In Ahab's time, Hiel of Bethel rebuilt Jericho. He laid its foundations at the cost of his firstborn son Abiram, and he set up its gates at the cost of his youngest son Segub, in accordance with the word of the LORD spoken by Joshua son of Nun.
1KGS|17|1|Now Elijah the Tishbite, from Tishbe in Gilead, said to Ahab, "As the LORD, the God of Israel, lives, whom I serve, there will be neither dew nor rain in the next few years except at my word."
1KGS|17|2|Then the word of the LORD came to Elijah:
1KGS|17|3|"Leave here, turn eastward and hide in the Kerith Ravine, east of the Jordan.
1KGS|17|4|You will drink from the brook, and I have ordered the ravens to feed you there."
1KGS|17|5|So he did what the LORD had told him. He went to the Kerith Ravine, east of the Jordan, and stayed there.
1KGS|17|6|The ravens brought him bread and meat in the morning and bread and meat in the evening, and he drank from the brook.
1KGS|17|7|Some time later the brook dried up because there had been no rain in the land.
1KGS|17|8|Then the word of the LORD came to him:
1KGS|17|9|"Go at once to Zarephath of Sidon and stay there. I have commanded a widow in that place to supply you with food."
1KGS|17|10|So he went to Zarephath. When he came to the town gate, a widow was there gathering sticks. He called to her and asked, "Would you bring me a little water in a jar so I may have a drink?"
1KGS|17|11|As she was going to get it, he called, "And bring me, please, a piece of bread."
1KGS|17|12|"As surely as the LORD your God lives," she replied, "I don't have any bread-only a handful of flour in a jar and a little oil in a jug. I am gathering a few sticks to take home and make a meal for myself and my son, that we may eat it-and die."
1KGS|17|13|Elijah said to her, "Don't be afraid. Go home and do as you have said. But first make a small cake of bread for me from what you have and bring it to me, and then make something for yourself and your son.
1KGS|17|14|For this is what the LORD, the God of Israel, says: 'The jar of flour will not be used up and the jug of oil will not run dry until the day the LORD gives rain on the land.'"
1KGS|17|15|She went away and did as Elijah had told her. So there was food every day for Elijah and for the woman and her family.
1KGS|17|16|For the jar of flour was not used up and the jug of oil did not run dry, in keeping with the word of the LORD spoken by Elijah.
1KGS|17|17|Some time later the son of the woman who owned the house became ill. He grew worse and worse, and finally stopped breathing.
1KGS|17|18|She said to Elijah, "What do you have against me, man of God? Did you come to remind me of my sin and kill my son?"
1KGS|17|19|"Give me your son," Elijah replied. He took him from her arms, carried him to the upper room where he was staying, and laid him on his bed.
1KGS|17|20|Then he cried out to the LORD, "O LORD my God, have you brought tragedy also upon this widow I am staying with, by causing her son to die?"
1KGS|17|21|Then he stretched himself out on the boy three times and cried to the LORD, "O LORD my God, let this boy's life return to him!"
1KGS|17|22|The LORD heard Elijah's cry, and the boy's life returned to him, and he lived.
1KGS|17|23|Elijah picked up the child and carried him down from the room into the house. He gave him to his mother and said, "Look, your son is alive!"
1KGS|17|24|Then the woman said to Elijah, "Now I know that you are a man of God and that the word of the LORD from your mouth is the truth."
1KGS|18|1|After a long time, in the third year, the word of the LORD came to Elijah: "Go and present yourself to Ahab, and I will send rain on the land."
1KGS|18|2|So Elijah went to present himself to Ahab. Now the famine was severe in Samaria,
1KGS|18|3|and Ahab had summoned Obadiah, who was in charge of his palace. (Obadiah was a devout believer in the LORD.
1KGS|18|4|While Jezebel was killing off the LORD's prophets, Obadiah had taken a hundred prophets and hidden them in two caves, fifty in each, and had supplied them with food and water.)
1KGS|18|5|Ahab had said to Obadiah, "Go through the land to all the springs and valleys. Maybe we can find some grass to keep the horses and mules alive so we will not have to kill any of our animals."
1KGS|18|6|So they divided the land they were to cover, Ahab going in one direction and Obadiah in another.
1KGS|18|7|As Obadiah was walking along, Elijah met him. Obadiah recognized him, bowed down to the ground, and said, "Is it really you, my lord Elijah?"
1KGS|18|8|"Yes," he replied. "Go tell your master, 'Elijah is here.'"
1KGS|18|9|"What have I done wrong," asked Obadiah, "that you are handing your servant over to Ahab to be put to death?
1KGS|18|10|As surely as the LORD your God lives, there is not a nation or kingdom where my master has not sent someone to look for you. And whenever a nation or kingdom claimed you were not there, he made them swear they could not find you.
1KGS|18|11|But now you tell me to go to my master and say, 'Elijah is here.'
1KGS|18|12|I don't know where the Spirit of the LORD may carry you when I leave you. If I go and tell Ahab and he doesn't find you, he will kill me. Yet I your servant have worshiped the LORD since my youth.
1KGS|18|13|Haven't you heard, my lord, what I did while Jezebel was killing the prophets of the LORD? I hid a hundred of the LORD's prophets in two caves, fifty in each, and supplied them with food and water.
1KGS|18|14|And now you tell me to go to my master and say, 'Elijah is here.' He will kill me!"
1KGS|18|15|Elijah said, "As the LORD Almighty lives, whom I serve, I will surely present myself to Ahab today."
1KGS|18|16|So Obadiah went to meet Ahab and told him, and Ahab went to meet Elijah.
1KGS|18|17|When he saw Elijah, he said to him, "Is that you, you troubler of Israel?"
1KGS|18|18|"I have not made trouble for Israel," Elijah replied. "But you and your father's family have. You have abandoned the LORD's commands and have followed the Baals.
1KGS|18|19|Now summon the people from all over Israel to meet me on Mount Carmel. And bring the four hundred and fifty prophets of Baal and the four hundred prophets of Asherah, who eat at Jezebel's table."
1KGS|18|20|So Ahab sent word throughout all Israel and assembled the prophets on Mount Carmel.
1KGS|18|21|Elijah went before the people and said, "How long will you waver between two opinions? If the LORD is God, follow him; but if Baal is God, follow him." But the people said nothing.
1KGS|18|22|Then Elijah said to them, "I am the only one of the LORD's prophets left, but Baal has four hundred and fifty prophets.
1KGS|18|23|Get two bulls for us. Let them choose one for themselves, and let them cut it into pieces and put it on the wood but not set fire to it. I will prepare the other bull and put it on the wood but not set fire to it.
1KGS|18|24|Then you call on the name of your god, and I will call on the name of the LORD. The god who answers by fire-he is God." Then all the people said, "What you say is good."
1KGS|18|25|Elijah said to the prophets of Baal, "Choose one of the bulls and prepare it first, since there are so many of you. Call on the name of your god, but do not light the fire."
1KGS|18|26|So they took the bull given them and prepared it. Then they called on the name of Baal from morning till noon. "O Baal, answer us!" they shouted. But there was no response; no one answered. And they danced around the altar they had made.
1KGS|18|27|At noon Elijah began to taunt them. "Shout louder!" he said. "Surely he is a god! Perhaps he is deep in thought, or busy, or traveling. Maybe he is sleeping and must be awakened."
1KGS|18|28|So they shouted louder and slashed themselves with swords and spears, as was their custom, until their blood flowed.
1KGS|18|29|Midday passed, and they continued their frantic prophesying until the time for the evening sacrifice. But there was no response, no one answered, no one paid attention.
1KGS|18|30|Then Elijah said to all the people, "Come here to me." They came to him, and he repaired the altar of the LORD, which was in ruins.
1KGS|18|31|Elijah took twelve stones, one for each of the tribes descended from Jacob, to whom the word of the LORD had come, saying, "Your name shall be Israel."
1KGS|18|32|With the stones he built an altar in the name of the LORD, and he dug a trench around it large enough to hold two seahs of seed.
1KGS|18|33|He arranged the wood, cut the bull into pieces and laid it on the wood. Then he said to them, "Fill four large jars with water and pour it on the offering and on the wood."
1KGS|18|34|"Do it again," he said, and they did it again. "Do it a third time," he ordered, and they did it the third time.
1KGS|18|35|The water ran down around the altar and even filled the trench.
1KGS|18|36|At the time of sacrifice, the prophet Elijah stepped forward and prayed: "O LORD, God of Abraham, Isaac and Israel, let it be known today that you are God in Israel and that I am your servant and have done all these things at your command.
1KGS|18|37|Answer me, O LORD, answer me, so these people will know that you, O LORD, are God, and that you are turning their hearts back again."
1KGS|18|38|Then the fire of the LORD fell and burned up the sacrifice, the wood, the stones and the soil, and also licked up the water in the trench.
1KGS|18|39|When all the people saw this, they fell prostrate and cried, "The LORD -he is God! The LORD -he is God!"
1KGS|18|40|Then Elijah commanded them, "Seize the prophets of Baal. Don't let anyone get away!" They seized them, and Elijah had them brought down to the Kishon Valley and slaughtered there.
1KGS|18|41|And Elijah said to Ahab, "Go, eat and drink, for there is the sound of a heavy rain."
1KGS|18|42|So Ahab went off to eat and drink, but Elijah climbed to the top of Carmel, bent down to the ground and put his face between his knees.
1KGS|18|43|"Go and look toward the sea," he told his servant. And he went up and looked. "There is nothing there," he said. Seven times Elijah said, "Go back."
1KGS|18|44|The seventh time the servant reported, "A cloud as small as a man's hand is rising from the sea." So Elijah said, "Go and tell Ahab, 'Hitch up your chariot and go down before the rain stops you.'"
1KGS|18|45|Meanwhile, the sky grew black with clouds, the wind rose, a heavy rain came on and Ahab rode off to Jezreel.
1KGS|18|46|The power of the LORD came upon Elijah and, tucking his cloak into his belt, he ran ahead of Ahab all the way to Jezreel.
1KGS|19|1|Now Ahab told Jezebel everything Elijah had done and how he had killed all the prophets with the sword.
1KGS|19|2|So Jezebel sent a messenger to Elijah to say, "May the gods deal with me, be it ever so severely, if by this time tomorrow I do not make your life like that of one of them."
1KGS|19|3|Elijah was afraid and ran for his life. When he came to Beersheba in Judah, he left his servant there,
1KGS|19|4|while he himself went a day's journey into the desert. He came to a broom tree, sat down under it and prayed that he might die. "I have had enough, LORD," he said. "Take my life; I am no better than my ancestors."
1KGS|19|5|Then he lay down under the tree and fell asleep. All at once an angel touched him and said, "Get up and eat."
1KGS|19|6|He looked around, and there by his head was a cake of bread baked over hot coals, and a jar of water. He ate and drank and then lay down again.
1KGS|19|7|The angel of the LORD came back a second time and touched him and said, "Get up and eat, for the journey is too much for you."
1KGS|19|8|So he got up and ate and drank. Strengthened by that food, he traveled forty days and forty nights until he reached Horeb, the mountain of God.
1KGS|19|9|There he went into a cave and spent the night. And the word of the LORD came to him: "What are you doing here, Elijah?"
1KGS|19|10|He replied, "I have been very zealous for the LORD God Almighty. The Israelites have rejected your covenant, broken down your altars, and put your prophets to death with the sword. I am the only one left, and now they are trying to kill me too."
1KGS|19|11|The LORD said, "Go out and stand on the mountain in the presence of the LORD, for the LORD is about to pass by." Then a great and powerful wind tore the mountains apart and shattered the rocks before the LORD, but the LORD was not in the wind. After the wind there was an earthquake, but the LORD was not in the earthquake.
1KGS|19|12|After the earthquake came a fire, but the LORD was not in the fire. And after the fire came a gentle whisper.
1KGS|19|13|When Elijah heard it, he pulled his cloak over his face and went out and stood at the mouth of the cave. Then a voice said to him, "What are you doing here, Elijah?"
1KGS|19|14|He replied, "I have been very zealous for the LORD God Almighty. The Israelites have rejected your covenant, broken down your altars, and put your prophets to death with the sword. I am the only one left, and now they are trying to kill me too."
1KGS|19|15|The LORD said to him, "Go back the way you came, and go to the Desert of Damascus. When you get there, anoint Hazael king over Aram.
1KGS|19|16|Also, anoint Jehu son of Nimshi king over Israel, and anoint Elisha son of Shaphat from Abel Meholah to succeed you as prophet.
1KGS|19|17|Jehu will put to death any who escape the sword of Hazael, and Elisha will put to death any who escape the sword of Jehu.
1KGS|19|18|Yet I reserve seven thousand in Israel-all whose knees have not bowed down to Baal and all whose mouths have not kissed him."
1KGS|19|19|So Elijah went from there and found Elisha son of Shaphat. He was plowing with twelve yoke of oxen, and he himself was driving the twelfth pair. Elijah went up to him and threw his cloak around him.
1KGS|19|20|Elisha then left his oxen and ran after Elijah. "Let me kiss my father and mother good-by," he said, "and then I will come with you.Go back," Elijah replied. "What have I done to you?"
1KGS|19|21|So Elisha left him and went back. He took his yoke of oxen and slaughtered them. He burned the plowing equipment to cook the meat and gave it to the people, and they ate. Then he set out to follow Elijah and became his attendant.
1KGS|20|1|Now Ben-Hadad king of Aram mustered his entire army. Accompanied by thirty-two kings with their horses and chariots, he went up and besieged Samaria and attacked it.
1KGS|20|2|He sent messengers into the city to Ahab king of Israel, saying, "This is what Ben-Hadad says:
1KGS|20|3|'Your silver and gold are mine, and the best of your wives and children are mine.'"
1KGS|20|4|The king of Israel answered, "Just as you say, my lord the king. I and all I have are yours."
1KGS|20|5|The messengers came again and said, "This is what Ben-Hadad says: 'I sent to demand your silver and gold, your wives and your children.
1KGS|20|6|But about this time tomorrow I am going to send my officials to search your palace and the houses of your officials. They will seize everything you value and carry it away.'"
1KGS|20|7|The king of Israel summoned all the elders of the land and said to them, "See how this man is looking for trouble! When he sent for my wives and my children, my silver and my gold, I did not refuse him."
1KGS|20|8|The elders and the people all answered, "Don't listen to him or agree to his demands."
1KGS|20|9|So he replied to Ben-Hadad's messengers, "Tell my lord the king, 'Your servant will do all you demanded the first time, but this demand I cannot meet.'" They left and took the answer back to Ben-Hadad.
1KGS|20|10|Then Ben-Hadad sent another message to Ahab: "May the gods deal with me, be it ever so severely, if enough dust remains in Samaria to give each of my men a handful."
1KGS|20|11|The king of Israel answered, "Tell him: 'One who puts on his armor should not boast like one who takes it off.'"
1KGS|20|12|Ben-Hadad heard this message while he and the kings were drinking in their tents, and he ordered his men: "Prepare to attack." So they prepared to attack the city.
1KGS|20|13|Meanwhile a prophet came to Ahab king of Israel and announced, "This is what the LORD says: 'Do you see this vast army? I will give it into your hand today, and then you will know that I am the LORD.'"
1KGS|20|14|"But who will do this?" asked Ahab. The prophet replied, "This is what the LORD says: 'The young officers of the provincial commanders will do it.' And who will start the battle?" he asked. The prophet answered, "You will."
1KGS|20|15|So Ahab summoned the young officers of the provincial commanders, 232 men. Then he assembled the rest of the Israelites, 7,000 in all.
1KGS|20|16|They set out at noon while Ben-Hadad and the 32 kings allied with him were in their tents getting drunk.
1KGS|20|17|The young officers of the provincial commanders went out first. Now Ben-Hadad had dispatched scouts, who reported, "Men are advancing from Samaria."
1KGS|20|18|He said, "If they have come out for peace, take them alive; if they have come out for war, take them alive."
1KGS|20|19|The young officers of the provincial commanders marched out of the city with the army behind them
1KGS|20|20|and each one struck down his opponent. At that, the Arameans fled, with the Israelites in pursuit. But Ben-Hadad king of Aram escaped on horseback with some of his horsemen.
1KGS|20|21|The king of Israel advanced and overpowered the horses and chariots and inflicted heavy losses on the Arameans.
1KGS|20|22|Afterward, the prophet came to the king of Israel and said, "Strengthen your position and see what must be done, because next spring the king of Aram will attack you again."
1KGS|20|23|Meanwhile, the officials of the king of Aram advised him, "Their gods are gods of the hills. That is why they were too strong for us. But if we fight them on the plains, surely we will be stronger than they.
1KGS|20|24|Do this: Remove all the kings from their commands and replace them with other officers.
1KGS|20|25|You must also raise an army like the one you lost-horse for horse and chariot for chariot-so we can fight Israel on the plains. Then surely we will be stronger than they." He agreed with them and acted accordingly.
1KGS|20|26|The next spring Ben-Hadad mustered the Arameans and went up to Aphek to fight against Israel.
1KGS|20|27|When the Israelites were also mustered and given provisions, they marched out to meet them. The Israelites camped opposite them like two small flocks of goats, while the Arameans covered the countryside.
1KGS|20|28|The man of God came up and told the king of Israel, "This is what the LORD says: 'Because the Arameans think the LORD is a god of the hills and not a god of the valleys, I will deliver this vast army into your hands, and you will know that I am the LORD.'"
1KGS|20|29|For seven days they camped opposite each other, and on the seventh day the battle was joined. The Israelites inflicted a hundred thousand casualties on the Aramean foot soldiers in one day.
1KGS|20|30|The rest of them escaped to the city of Aphek, where the wall collapsed on twenty-seven thousand of them. And Ben-Hadad fled to the city and hid in an inner room.
1KGS|20|31|His officials said to him, "Look, we have heard that the kings of the house of Israel are merciful. Let us go to the king of Israel with sackcloth around our waists and ropes around our heads. Perhaps he will spare your life."
1KGS|20|32|Wearing sackcloth around their waists and ropes around their heads, they went to the king of Israel and said, "Your servant Ben-Hadad says: 'Please let me live.'" The king answered, "Is he still alive? He is my brother."
1KGS|20|33|The men took this as a good sign and were quick to pick up his word. "Yes, your brother Ben-Hadad!" they said. "Go and get him," the king said. When Ben-Hadad came out, Ahab had him come up into his chariot.
1KGS|20|34|"I will return the cities my father took from your father," Ben-Hadad offered. "You may set up your own market areas in Damascus, as my father did in Samaria." Ahab said, "On the basis of a treaty I will set you free." So he made a treaty with him, and let him go.
1KGS|20|35|By the word of the LORD one of the sons of the prophets said to his companion, "Strike me with your weapon," but the man refused.
1KGS|20|36|So the prophet said, "Because you have not obeyed the LORD, as soon as you leave me a lion will kill you." And after the man went away, a lion found him and killed him.
1KGS|20|37|The prophet found another man and said, "Strike me, please." So the man struck him and wounded him.
1KGS|20|38|Then the prophet went and stood by the road waiting for the king. He disguised himself with his headband down over his eyes.
1KGS|20|39|As the king passed by, the prophet called out to him, "Your servant went into the thick of the battle, and someone came to me with a captive and said, 'Guard this man. If he is missing, it will be your life for his life, or you must pay a talent of silver.'
1KGS|20|40|While your servant was busy here and there, the man disappeared.That is your sentence," the king of Israel said. "You have pronounced it yourself."
1KGS|20|41|Then the prophet quickly removed the headband from his eyes, and the king of Israel recognized him as one of the prophets.
1KGS|20|42|He said to the king, "This is what the LORD says: 'You have set free a man I had determined should die. Therefore it is your life for his life, your people for his people.'"
1KGS|20|43|Sullen and angry, the king of Israel went to his palace in Samaria.
1KGS|21|1|Some time later there was an incident involving a vineyard belonging to Naboth the Jezreelite. The vineyard was in Jezreel, close to the palace of Ahab king of Samaria.
1KGS|21|2|Ahab said to Naboth, "Let me have your vineyard to use for a vegetable garden, since it is close to my palace. In exchange I will give you a better vineyard or, if you prefer, I will pay you whatever it is worth."
1KGS|21|3|But Naboth replied, "The LORD forbid that I should give you the inheritance of my fathers."
1KGS|21|4|So Ahab went home, sullen and angry because Naboth the Jezreelite had said, "I will not give you the inheritance of my fathers." He lay on his bed sulking and refused to eat.
1KGS|21|5|His wife Jezebel came in and asked him, "Why are you so sullen? Why won't you eat?"
1KGS|21|6|He answered her, "Because I said to Naboth the Jezreelite, 'Sell me your vineyard; or if you prefer, I will give you another vineyard in its place.' But he said, 'I will not give you my vineyard.'"
1KGS|21|7|Jezebel his wife said, "Is this how you act as king over Israel? Get up and eat! Cheer up. I'll get you the vineyard of Naboth the Jezreelite."
1KGS|21|8|So she wrote letters in Ahab's name, placed his seal on them, and sent them to the elders and nobles who lived in Naboth's city with him.
1KGS|21|9|In those letters she wrote: "Proclaim a day of fasting and seat Naboth in a prominent place among the people.
1KGS|21|10|But seat two scoundrels opposite him and have them testify that he has cursed both God and the king. Then take him out and stone him to death."
1KGS|21|11|So the elders and nobles who lived in Naboth's city did as Jezebel directed in the letters she had written to them.
1KGS|21|12|They proclaimed a fast and seated Naboth in a prominent place among the people.
1KGS|21|13|Then two scoundrels came and sat opposite him and brought charges against Naboth before the people, saying, "Naboth has cursed both God and the king." So they took him outside the city and stoned him to death.
1KGS|21|14|Then they sent word to Jezebel: "Naboth has been stoned and is dead."
1KGS|21|15|As soon as Jezebel heard that Naboth had been stoned to death, she said to Ahab, "Get up and take possession of the vineyard of Naboth the Jezreelite that he refused to sell you. He is no longer alive, but dead."
1KGS|21|16|When Ahab heard that Naboth was dead, he got up and went down to take possession of Naboth's vineyard.
1KGS|21|17|Then the word of the LORD came to Elijah the Tishbite:
1KGS|21|18|"Go down to meet Ahab king of Israel, who rules in Samaria. He is now in Naboth's vineyard, where he has gone to take possession of it.
1KGS|21|19|Say to him, 'This is what the LORD says: Have you not murdered a man and seized his property?' Then say to him, 'This is what the LORD says: In the place where dogs licked up Naboth's blood, dogs will lick up your blood-yes, yours!'"
1KGS|21|20|Ahab said to Elijah, "So you have found me, my enemy!I have found you," he answered, "because you have sold yourself to do evil in the eyes of the LORD.
1KGS|21|21|'I am going to bring disaster on you. I will consume your descendants and cut off from Ahab every last male in Israel-slave or free.
1KGS|21|22|I will make your house like that of Jeroboam son of Nebat and that of Baasha son of Ahijah, because you have provoked me to anger and have caused Israel to sin.'
1KGS|21|23|"And also concerning Jezebel the LORD says: 'Dogs will devour Jezebel by the wall of Jezreel.'
1KGS|21|24|"Dogs will eat those belonging to Ahab who die in the city, and the birds of the air will feed on those who die in the country."
1KGS|21|25|(There was never a man like Ahab, who sold himself to do evil in the eyes of the LORD, urged on by Jezebel his wife.
1KGS|21|26|He behaved in the vilest manner by going after idols, like the Amorites the LORD drove out before Israel.)
1KGS|21|27|When Ahab heard these words, he tore his clothes, put on sackcloth and fasted. He lay in sackcloth and went around meekly.
1KGS|21|28|Then the word of the LORD came to Elijah the Tishbite:
1KGS|21|29|"Have you noticed how Ahab has humbled himself before me? Because he has humbled himself, I will not bring this disaster in his day, but I will bring it on his house in the days of his son."
1KGS|22|1|For three years there was no war between Aram and Israel.
1KGS|22|2|But in the third year Jehoshaphat king of Judah went down to see the king of Israel.
1KGS|22|3|The king of Israel had said to his officials, "Don't you know that Ramoth Gilead belongs to us and yet we are doing nothing to retake it from the king of Aram?"
1KGS|22|4|So he asked Jehoshaphat, "Will you go with me to fight against Ramoth Gilead?" Jehoshaphat replied to the king of Israel, "I am as you are, my people as your people, my horses as your horses."
1KGS|22|5|But Jehoshaphat also said to the king of Israel, "First seek the counsel of the LORD."
1KGS|22|6|So the king of Israel brought together the prophets-about four hundred men-and asked them, "Shall I go to war against Ramoth Gilead, or shall I refrain?Go," they answered, "for the Lord will give it into the king's hand."
1KGS|22|7|But Jehoshaphat asked, "Is there not a prophet of the LORD here whom we can inquire of?"
1KGS|22|8|The king of Israel answered Jehoshaphat, "There is still one man through whom we can inquire of the LORD, but I hate him because he never prophesies anything good about me, but always bad. He is Micaiah son of Imlah.The king should not say that," Jehoshaphat replied.
1KGS|22|9|So the king of Israel called one of his officials and said, "Bring Micaiah son of Imlah at once."
1KGS|22|10|Dressed in their royal robes, the king of Israel and Jehoshaphat king of Judah were sitting on their thrones at the threshing floor by the entrance of the gate of Samaria, with all the prophets prophesying before them.
1KGS|22|11|Now Zedekiah son of Kenaanah had made iron horns and he declared, "This is what the LORD says: 'With these you will gore the Arameans until they are destroyed.'"
1KGS|22|12|All the other prophets were prophesying the same thing. "Attack Ramoth Gilead and be victorious," they said, "for the LORD will give it into the king's hand."
1KGS|22|13|The messenger who had gone to summon Micaiah said to him, "Look, as one man the other prophets are predicting success for the king. Let your word agree with theirs, and speak favorably."
1KGS|22|14|But Micaiah said, "As surely as the LORD lives, I can tell him only what the LORD tells me."
1KGS|22|15|When he arrived, the king asked him, "Micaiah, shall we go to war against Ramoth Gilead, or shall I refrain?Attack and be victorious," he answered, "for the LORD will give it into the king's hand."
1KGS|22|16|The king said to him, "How many times must I make you swear to tell me nothing but the truth in the name of the LORD?"
1KGS|22|17|Then Micaiah answered, "I saw all Israel scattered on the hills like sheep without a shepherd, and the LORD said, 'These people have no master. Let each one go home in peace.'"
1KGS|22|18|The king of Israel said to Jehoshaphat, "Didn't I tell you that he never prophesies anything good about me, but only bad?"
1KGS|22|19|Micaiah continued, "Therefore hear the word of the LORD: I saw the LORD sitting on his throne with all the host of heaven standing around him on his right and on his left.
1KGS|22|20|And the LORD said, 'Who will entice Ahab into attacking Ramoth Gilead and going to his death there?'"One suggested this, and another that.
1KGS|22|21|Finally, a spirit came forward, stood before the LORD and said, 'I will entice him.'
1KGS|22|22|"'By what means?' the LORD asked. "'I will go out and be a lying spirit in the mouths of all his prophets,' he said. "'You will succeed in enticing him,' said the LORD. 'Go and do it.'
1KGS|22|23|"So now the LORD has put a lying spirit in the mouths of all these prophets of yours. The LORD has decreed disaster for you."
1KGS|22|24|Then Zedekiah son of Kenaanah went up and slapped Micaiah in the face. "Which way did the spirit from the LORD go when he went from me to speak to you?" he asked.
1KGS|22|25|Micaiah replied, "You will find out on the day you go to hide in an inner room."
1KGS|22|26|The king of Israel then ordered, "Take Micaiah and send him back to Amon the ruler of the city and to Joash the king's son
1KGS|22|27|and say, 'This is what the king says: Put this fellow in prison and give him nothing but bread and water until I return safely.'"
1KGS|22|28|Micaiah declared, "If you ever return safely, the LORD has not spoken through me." Then he added, "Mark my words, all you people!"
1KGS|22|29|So the king of Israel and Jehoshaphat king of Judah went up to Ramoth Gilead.
1KGS|22|30|The king of Israel said to Jehoshaphat, "I will enter the battle in disguise, but you wear your royal robes." So the king of Israel disguised himself and went into battle.
1KGS|22|31|Now the king of Aram had ordered his thirty-two chariot commanders, "Do not fight with anyone, small or great, except the king of Israel."
1KGS|22|32|When the chariot commanders saw Jehoshaphat, they thought, "Surely this is the king of Israel." So they turned to attack him, but when Jehoshaphat cried out,
1KGS|22|33|the chariot commanders saw that he was not the king of Israel and stopped pursuing him.
1KGS|22|34|But someone drew his bow at random and hit the king of Israel between the sections of his armor. The king told his chariot driver, "Wheel around and get me out of the fighting. I've been wounded."
1KGS|22|35|All day long the battle raged, and the king was propped up in his chariot facing the Arameans. The blood from his wound ran onto the floor of the chariot, and that evening he died.
1KGS|22|36|As the sun was setting, a cry spread through the army: "Every man to his town; everyone to his land!"
1KGS|22|37|So the king died and was brought to Samaria, and they buried him there.
1KGS|22|38|They washed the chariot at a pool in Samaria (where the prostitutes bathed), and the dogs licked up his blood, as the word of the LORD had declared.
1KGS|22|39|As for the other events of Ahab's reign, including all he did, the palace he built and inlaid with ivory, and the cities he fortified, are they not written in the book of the annals of the kings of Israel?
1KGS|22|40|Ahab rested with his fathers. And Ahaziah his son succeeded him as king.
1KGS|22|41|Jehoshaphat son of Asa became king of Judah in the fourth year of Ahab king of Israel.
1KGS|22|42|Jehoshaphat was thirty-five years old when he became king, and he reigned in Jerusalem twenty-five years. His mother's name was Azubah daughter of Shilhi.
1KGS|22|43|In everything he walked in the ways of his father Asa and did not stray from them; he did what was right in the eyes of the LORD. The high places, however, were not removed, and the people continued to offer sacrifices and burn incense there.
1KGS|22|44|Jehoshaphat was also at peace with the king of Israel.
1KGS|22|45|As for the other events of Jehoshaphat's reign, the things he achieved and his military exploits, are they not written in the book of the annals of the kings of Judah?
1KGS|22|46|He rid the land of the rest of the male shrine prostitutes who remained there even after the reign of his father Asa.
1KGS|22|47|There was then no king in Edom; a deputy ruled.
1KGS|22|48|Now Jehoshaphat built a fleet of trading ships to go to Ophir for gold, but they never set sail-they were wrecked at Ezion Geber.
1KGS|22|49|At that time Ahaziah son of Ahab said to Jehoshaphat, "Let my men sail with your men," but Jehoshaphat refused.
1KGS|22|50|Then Jehoshaphat rested with his fathers and was buried with them in the city of David his father. And Jehoram his son succeeded him.
1KGS|22|51|Ahaziah son of Ahab became king of Israel in Samaria in the seventeenth year of Jehoshaphat king of Judah, and he reigned over Israel two years.
1KGS|22|52|He did evil in the eyes of the LORD, because he walked in the ways of his father and mother and in the ways of Jeroboam son of Nebat, who caused Israel to sin.
1KGS|22|53|He served and worshiped Baal and provoked the LORD, the God of Israel, to anger, just as his father had done.
