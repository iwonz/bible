2COR|1|1|Paulus, apostolus Christi Iesu per voluntatem Dei, et Timo theus frater ecclesiae Dei, quae est Corinthi, cum sanctis omnibus, qui sunt in universa Achaia:
2COR|1|2|gratia vobis et pax a Deo Patre nostro et Domino Iesu Christo.
2COR|1|3|Benedictus Deus et Pater Domini nostri Iesu Christi, Pater misericordiarum et Deus totius consolationis,
2COR|1|4|qui consolatur nos in omni tribulatione nostra, ut possimus et ipsi consolari eos, qui in omni pressura sunt, per exhortationem, qua exhortamur et ipsi a Deo;
2COR|1|5|quoniam, sicut abundant passiones Christi in nobis, ita per Christum abundat et consolatio nostra.
2COR|1|6|Sive autem tribulamur, pro vestra exhortatione et salute; sive exhortamur, pro vestra exhortatione, quae operatur in tolerantia earundem passionum, quas et nos patimur.
2COR|1|7|Et spes nostra firma pro vobis, scientes quoniam, sicut socii passionum estis, sic eritis et consolationis.
2COR|1|8|Non enim volumus ignorare vos, fratres, de tribulatione nostra, quae facta est in Asia, quoniam supra modum gravati sumus supra virtutem, ita ut taederet nos etiam vivere;
2COR|1|9|sed ipsi in nobis ipsis responsum mortis habuimus, ut non simus fidentes in nobis sed in Deo, qui suscitat mortuos:
2COR|1|10|qui de tanta morte eripuit nos et eruet, in quem speramus, et adhuc eripiet;
2COR|1|11|adiuvantibus et vobis in oratione pro nobis, ut propter eam, quae ex multis personis in nos est, donationem, per multos gratiae agantur pro nobis.
2COR|1|12|Nam gloria nostra haec est, testimonium conscientiae nostrae, quod in simplicitate et sinceritate Dei et non in sapientia carnali, sed in gratia Dei conversati sumus in mundo, abundantius autem ad vos.
2COR|1|13|Non enim alia scribimus vobis quam quae legitis aut etiam cognoscitis; spero autem quod usque in finem cognoscetis,
2COR|1|14|sicut et cognovistis nos ex parte, quia gloria vestra sumus, sicut et vos nostra in die Domini nostri Iesu.
2COR|1|15|Et hac confidentia volui prius venire ad vos, ut secundam gratiam haberetis,
2COR|1|16|et per vos transire in Macedoniam et iterum a Macedonia venire ad vos et a vobis deduci in Iudaeam.
2COR|1|17|Cum hoc ergo voluissem, numquid levitate usus sum? Aut, quae cogito, secundum carnem cogito, ut sit apud me " Est, est " et " Non, non "?
2COR|1|18|Fidelis autem Deus, quia sermo noster, qui fit apud vos, non est " Est et " Non "!
2COR|1|19|Dei enim Filius Iesus Christus, qui in vobis per nos praedicatus est, per me et Silvanum et Timotheum, non fuit " Est " et " Non ", sed " Est " in illo fuit.
2COR|1|20|Quotquot enim promissiones Dei sunt, in illo " Est "; ideo et per ipsum Amen " Deo ad gloriam per nos.
2COR|1|21|Qui autem confirmat nos vobiscum in Christum et qui unxit nos, Deus,
2COR|1|22|et qui signavit nos et dedit arrabonem Spiritus in cordibus nostris.
2COR|1|23|Ego autem testem Deum invoco in animam meam, quod parcens vobis non veni ultra Corinthum.
2COR|1|24|Non quia dominamur fidei vestrae, sed adiutores sumus gaudii vestri, nam fide stetistis.
2COR|2|1|Statui autem hoc ipse apud me, ne iterum in tristitia venirem ad vos;
2COR|2|2|si enim ego contristo vos, et quis est qui me laetificet, nisi qui contristatur ex me?
2COR|2|3|Et hoc ipsum scripsi, ut non, cum venero, tristitiam habeam de quibus oportebat me gaudere, confidens in omnibus vobis, quia meum gaudium omnium vestrum est.
2COR|2|4|Nam ex multa tribulatione et angustia cordis scripsi vobis per multas lacrimas, non ut contristemini, sed ut sciatis quam carita tem habeo abundantius in vos.
2COR|2|5|Si quis autem contristavit, non me contristavit, sed ex parte, ut non onerem, omnes vos.
2COR|2|6|Sufficit illi, qui eiusmodi est, obiurgatio haec, quae fit a pluribus,
2COR|2|7|ita ut e contra magis donetis et consolemini, ne forte abundantiore tristitia absorbeatur, qui eiusmodi est.
2COR|2|8|Propter quod obsecro vos, ut confirmetis in illum caritatem;
2COR|2|9|ideo enim et scripsi, ut cognoscam probationem vestram, an in omnibus oboedientes sitis.
2COR|2|10|Cui autem aliquid donatis, et ego; nam et ego, quod donavi, si quid donavi, propter vos in persona Christi,
2COR|2|11|ut non circumveniamur a Satana; non enim ignoramus cogitationes eius.
2COR|2|12|Cum venissem autem Troadem ob evangelium Christi, et ostium mihi apertum esset in Domino,
2COR|2|13|non habui requiem spiritui meo, eo quod non invenerim Titum fratrem meum, sed valefaciens eis profectus sum in Macedoniam.
2COR|2|14|Deo autem gratias, qui semper triumphat nos in Christo et odorem notitiae suae manifestat per nos in omni loco.
2COR|2|15|Quia Christi bonus odor sumus Deo in his, qui salvi fiunt, et in his, qui pereunt:
2COR|2|16|aliis quidem odor ex morte in mortem, aliis autem odor ex vita in vitam. Et ad haec quis idoneus?
2COR|2|17|Non enim sumus sicut plurimi adulterantes verbum Dei, sed sicut ex sinceritate, sed sicut ex Deo coram Deo in Christo loquimur.
2COR|3|1|Incipimus iterum nosmetipsos commendare? Aut numquid egemus, sicut quidam, commendaticiis epistulis ad vos aut ex vobis?
2COR|3|2|Epistula nostra vos estis, scripta in cordibus nostris, quae scitur et legitur ab omnibus hominibus;
2COR|3|3|manifestati quoniam epistula estis Christi ministrata a nobis, scripta non atramento sed Spiritu Dei vivi, non in tabulis lapideis sed in tabulis cordis carnalibus.
2COR|3|4|Fiduciam autem talem habemus per Christum ad Deum.
2COR|3|5|Non quod sufficientes simus cogitare aliquid a nobis quasi ex nobis, sed sufficientia nostra ex Deo est,
2COR|3|6|qui et idoneos nos fecit ministros Novi Testamenti, non litterae sed Spiritus: littera enim occidit, Spiritus autem vivificat.
2COR|3|7|Quod si ministratio mortis, litteris deformata in lapidibus, fuit in gloria, ita ut non possent intendere filii Israel in faciem Moysis propter gloriam vultus eius, quae evacuatur,
2COR|3|8|quomodo non magis ministratio Spiritus erit in gloria?
2COR|3|9|Nam si ministerium damnationis gloria est, multo magis abundat ministerium iustitiae in gloria.
2COR|3|10|Nam nec glorificatum est, quod claruit in hac parte, propter excellentem gloriam;
2COR|3|11|si enim, quod evacuatur, per gloriam est, multo magis, quod manet, in gloria est.
2COR|3|12|Habentes igitur talem spem multa fiducia utimur,
2COR|3|13|et non sicut Moyses: ponebat velamen super faciem suam, ut non intenderent filii Israel in finem illius quod evacuatur.
2COR|3|14|Sed obtusi sunt sensus eorum. Usque in hodiernum enim diem idipsum velamen in lectione Veteris Testamenti manet non revelatum, quoniam in Christo evacuatur;
2COR|3|15|sed usque in hodiernum diem, cum legitur Moyses, velamen est positum super cor eorum.
2COR|3|16|Quando autem conversus fuerit ad Dominum, aufertur velamen.
2COR|3|17|Dominus autem Spiritus est; ubi autem Spiritus Domini, ibi libertas.
2COR|3|18|Nos vero omnes revelata facie gloriam Domini speculantes, in eandem imaginem transformamur a claritate in clarita tem tamquam a Domini Spiritu.
2COR|4|1|Ideo habentes hanc ministra tionem, iuxta quod misericor diam consecuti sumus, non deficimus,
2COR|4|2|sed abdicavimus occulta dedecoris non ambulantes in astutia neque adulterantes verbum Dei, sed in manifestatione veritatis commendantes nosmetipsos ad omnem conscientiam hominum coram Deo.
2COR|4|3|Quod si etiam velatum est evangelium nostrum, in his, qui pereunt, est velatum;
2COR|4|4|in quibus deus huius saeculi excaecavit mentes infidelium, ut non fulgeat illuminatio evangelii gloriae Christi, qui est imago Dei.
2COR|4|5|Non enim nosmetipsos praedicamus sed Iesum Christum Dominum; nos autem servos vestros per Iesum.
2COR|4|6|Quoniam Deus, qui dixit: " De tenebris lux splendescat ", ipse illuxit in cordibus nostris ad illuminationem scientiae claritatis Dei in facie Iesu Christi.
2COR|4|7|Habemus autem thesaurum istum in vasis fictilibus, ut sublimitas sit virtutis Dei et non ex nobis.
2COR|4|8|In omnibus tribulationem patimur, sed non angustiamur; aporiamur, sed non destituimur;
2COR|4|9|persecutionem patimur, sed non derelinquimur; deicimur, sed non perimus;
2COR|4|10|semper mortificationem Iesu in corpore circumferentes, ut et vita Iesu in corpore nostro manifestetur.
2COR|4|11|Semper enim nos, qui vivimus, in mortem tradimur propter Iesum, ut et vita Iesu manifestetur in carne nostra mortali.
2COR|4|12|Ergo mors in nobis operatur, vita autem in vobis.
2COR|4|13|Habentes autem eundem spiritum fidei, sicut scriptum est: " Credidi, propter quod locutus sum ", et nos credimus, propter quod et loquimur,
2COR|4|14|scientes quoniam, qui suscitavit Dominum Iesum, et nos cum Iesu suscitabit et constituet vobiscum.
2COR|4|15|Omnia enim propter vos, ut gratia abundans per multos gratiarum actionem abundare faciat in gloriam Dei.
2COR|4|16|Propter quod non deficimus, sed licet is, qui foris est, noster homo corrumpitur, tamen is, qui intus est, noster renovatur de die in diem.
2COR|4|17|Id enim, quod in praesenti est, leve tribulationis nostrae supra modum in sublimitatem aeternum gloriae pondus operatur nobis,
2COR|4|18|non contemplantibus nobis, quae videntur, sed quae non videntur; quae enim videntur, temporalia sunt, quae autem non videntur, aeterna sunt.
2COR|5|1|Scimus enim quoniam, si terre stris domus nostra huius taber naculi dissolvatur, aedificationem ex Deo habemus domum non manufactam, aeternam in caelis.
2COR|5|2|Nam et in hoc ingemiscimus, habitationem nostram, quae de caelo est, superindui cupientes,
2COR|5|3|si tamen et exspoliati, non nudi inveniamur.
2COR|5|4|Nam et, qui sumus in tabernaculo, ingemiscimus gravati, eo quod nolumus exspoliari, sed supervestiri, ut absorbeatur, quod mortale est, a vita.
2COR|5|5|Qui autem effecit nos in hoc ipsum, Deus, qui dedit nobis arrabonem Spiritus.
2COR|5|6|Audentes igitur semper et scientes quoniam, dum praesentes sumus in corpore, peregrinamur a Domino;
2COR|5|7|per fidem enim ambulamus et non per speciem.
2COR|5|8|Audemus autem et bonam voluntatem habemus magis peregrinari a corpore et praesentes esse ad Dominum.
2COR|5|9|Et ideo contendimus sive praesentes sive absentes placere illi.
2COR|5|10|Omnes enim nos manifestari oportet ante tribunal Christi, ut referat unusquisque pro eis, quae per corpus gessit, sive bonum sive malum.
2COR|5|11|Scientes ergo timorem Domini hominibus suademus, Deo autem manifesti sumus; spero autem et in conscientiis vestris manifestos nos esse.
2COR|5|12|Non iterum nos commendamus vobis, sed occasionem damus vobis gloriandi pro nobis, ut habeatis ad eos, qui in facie gloriantur et non in corde.
2COR|5|13|Sive enim mente excedimus, Deo; sive sobrii sumus, vobis.
2COR|5|14|Caritas enim Christi urget nos, aestimantes, hoc, quoniam, si unus pro omnibus mortuus est, ergo omnes mortui sunt;
2COR|5|15|et pro omnibus mortuus est, ut et, qui vivunt, iam non sibi vivant, sed ei, qui pro ipsis mortuus est et resurrexit.
2COR|5|16|Itaque nos ex hoc neminem novimus secundum carnem; et si cognovimus secundum carnem Christum, sed nunc iam non novimus.
2COR|5|17|Si quis ergo in Christo, nova creatura; vetera transierunt, ecce, facta sunt nova.
2COR|5|18|Omnia autem ex Deo, qui reconciliavit nos sibi per Christum et dedit nobis ministerium reconciliationis,
2COR|5|19|quoniam quidem Deus erat in Christo mundum reconcilians sibi, non reputans illis delicta ipsorum; et posuit in nobis verbum reconciliationis.
2COR|5|20|Pro Christo ergo legatione fungimur, tamquam Deo exhortante per nos. Obsecramus pro Christo, reconciliamini Deo.
2COR|5|21|Eum, qui non noverat peccatum, pro nobis peccatum fecit, ut nos efficeremur iustitia Dei in ipso.
2COR|6|1|Adiuvantes autem et exhor tamur, ne in vacuum gratiam Dei recipiatis
2COR|6|2|- ait enim: Tempore accepto exaudivi teet in die salutis adiuvi te ";ecce nunc tempus acceptabile, ecce nunc dies salutis -
2COR|6|3|nemini dantes ullam offensionem, ut non vituperetur ministerium,
2COR|6|4|sed in omnibus exhibentes nosmetipsos sicut Dei ministros in multa patientia, in tribulationibus, in necessitatibus, in angustiis,
2COR|6|5|in plagis, in carceribus, in seditionibus, in laboribus, in vigiliis, in ieiuniis,
2COR|6|6|in castitate, in scientia, in longanimitate, in suavitate, in Spiritu Sancto, in caritate non ficta,
2COR|6|7|in verbo veritatis, in virtute Dei; per arma iustitiae a dextris et sinistris,
2COR|6|8|per gloriam et ignobilitatem, per infamiam et bonam famam; ut seductores, et veraces;
2COR|6|9|sicut qui ignoti, et cogniti; quasi morientes, et ecce vivimus; ut castigati, et non mortificati;
2COR|6|10|quasi tristes, semper autem gaudentes; sicut egentes, multos autem locupletantes; tamquam nihil habentes, et omnia possidentes.
2COR|6|11|Os nostrum patet ad vos, o Corinthii, cor nostrum dilatatum est.
2COR|6|12|Non angustiamini in nobis, sed angustiamini in visceribus vestris;
2COR|6|13|eandem autem habentes remunerationem, tamquam filiis dico, dilatamini et vos.
2COR|6|14|Nolite iugum ducere cum infidelibus! Quae enim participatio iustitiae cum iniquitate? Aut quae societas luci ad tenebras?
2COR|6|15|Quae autem conventio Christi cum Beliar, aut quae pars fideli cum infideli?
2COR|6|16|Qui autem consensus templo Dei cum idolis? Vos enim estis templum Dei vivi; sicut dicit Deus: Inhabitabo in illis et inambulaboet ero illorum Deus, et ipsi erunt mihi populus.
2COR|6|17|Propter quod exite de medio eorumet separamini, dicit Dominus,et immundum ne tetigeritis;et ego recipiam vos
2COR|6|18|et ero vobis in Patrem,et vos eritis mihi in filios et filias,dicit Dominus omnipotens ".
2COR|7|1|Has igitur habentes promissio nes, carissimi, mundemus nos ab omni inquinamento carnis et spiritus, perficientes sanctificationem in timore Dei.
2COR|7|2|Capite nos! Neminem laesimus, neminem corrupimus, neminem circumvenimus.
2COR|7|3|Non ad condemnationem dico; praedixi enim quod in cordibus nostris estis ad commoriendum et ad convivendum.
2COR|7|4|Multa mihi fiducia est apud vos, multa mihi gloriatio pro vobis; repletus sum consolatione, superabundo gaudio in omni tribulatione nostra.
2COR|7|5|Nam et cum venissemus Macedoniam, nullam requiem habuit caro nostra, sed omnem tribulationem passi: foris pugnae, intus timores.
2COR|7|6|Sed qui consolatur humiles, consolatus est nos Deus in adventu Titi;
2COR|7|7|non solum autem in adventu eius sed etiam in solacio, quo consolatus est in vobis, referens nobis vestrum desiderium, vestrum fletum, vestram aemulationem pro me, ita ut magis gauderem.
2COR|7|8|Quoniam etsi contristavi vos in epistula, non me paenitet; etsi paeniteret - video quod epistula illa, etsi ad horam, vos contristavit -
2COR|7|9|nunc gaudeo, non quia contristati estis, sed quia contristati estis ad paenitentiam; contristati enim estis secundum Deum, ut in nullo detrimentum patiamini ex nobis.
2COR|7|10|Quae enim secundum Deum tristitia, paenitentiam in salutem stabilem operatur; saeculi autem tristitia mortem operatur.
2COR|7|11|Ecce enim hoc ipsum secundum Deum contristari: quantam in vobis operatum est sollicitudinem, sed defensionem, sed indignationem, sed timorem, sed desiderium, sed aemulationem, sed vindictam! In omnibus exhibuistis vos incontaminatos esse negotio.
2COR|7|12|Igitur etsi scripsi vobis, non propter eum, qui fecit iniuriam, nec propter eum, qui passus est, sed ad manifestandam sollicitudinem vestram, quam pro nobis habetis, ad vos coram Deo.
2COR|7|13|Ideo consolati sumus.In consolatione autem nostra abundantius magis gavisi sumus super gaudium Titi, quia refectus est spiritus eius ab omnibus vobis;
2COR|7|14|et si quid apud illum de vobis gloriatus sum, non sum confusus, sed sicut omnia vobis in veritate locuti sumus, ita et gloriatio nostra, quae fuit ad Titum, veritas facta est.
2COR|7|15|Et viscera eius abundantius in vos sunt, reminiscentis omnium vestrum oboedientiam, quomodo cum timore et tremore excepistis eum.
2COR|7|16|Gaudeo quod in omnibus confido in vobis.
2COR|8|1|Notam autem facimus vobis, fratres, gratiam Dei, quae data est in ecclesiis Macedoniae,
2COR|8|2|quod in multo experimento tribulationis abundantia gaudii ipsorum et altissima paupertas eorum abundavit in divitias simplicitatis eorum;
2COR|8|3|quia secundum virtutem, testimonium reddo, et supra virtutem voluntarii fuerunt
2COR|8|4|cum multa exhortatione obsecrantes nos gratiam et communicationem ministerii, quod fit in sanctos.
2COR|8|5|Et non sicut speravimus, sed semetipsos dederunt primum Domino, deinde nobis per voluntatem Dei,
2COR|8|6|ita ut rogaremus Titum, ut, quemadmodum coepit, ita et perficiat in vos etiam gratiam istam.
2COR|8|7|Sed sicut in omnibus abundatis, fide et sermone et scientia et omni sollicitudine et caritate ex nobis in vobis, ut et in hac gratia abundetis.
2COR|8|8|Non quasi imperans dico, sed per aliorum sollicitudinem etiam vestrae caritatis ingenitum bonum comprobans;
2COR|8|9|scitis enim gratiam Domini nostri Iesu Christi, quoniam propter vos egenus factus est, cum esset dives, ut illius inopia vos divites essetis.
2COR|8|10|Et consilium in hoc do. Hoc enim vobis utile est, qui non solum facere, sed et velle coepistis ab anno priore;
2COR|8|11|nunc vero et facto perficite, ut, quemadmodum promptus est animus velle, ita sit et perficere ex eo, quod habetis.
2COR|8|12|Si enim voluntas prompta est, secundum id quod habet, accepta est, non secundum quod non habet.
2COR|8|13|Non enim, ut aliis sit remissio, vobis autem tribulatio; sed ex aequalitate
2COR|8|14|in praesenti tempore vestra abundantia illorum inopiam suppleat, ut et illorum abundantia vestram inopiam suppleat, ut fiat aequalitas, sicut scriptum est:
2COR|8|15|" Qui multum, non abundavit; et, qui modicum, non minoravit ".
2COR|8|16|Gratias autem Deo, qui dedit eandem sollicitudinem pro vobis in corde Titi,
2COR|8|17|quoniam exhortationem quidem suscepit, sed, cum sollicitior esset, sua voluntate profectus est ad vos.
2COR|8|18|Misimus etiam cum illo fratrem, cuius laus est in evangelio per omnes ecclesias
2COR|8|19|- non solum autem, sed et ordinatus ab ecclesiis comes noster cum hac gratia, quae ministratur a nobis ad Domini gloriam et destinatam voluntatem nostram -
2COR|8|20|devitantes hoc, ne quis nos vituperet in hac plenitudine, quae ministratur a nobis;
2COR|8|21|providemus enim bona non solum coram Domino sed etiam coram hominibus.
2COR|8|22|Misimus autem cum illis et fratrem nostrum, quem probavimus in multis saepe sollicitum esse, nunc autem multo sollicitiorem, confidentia multa in vos.
2COR|8|23|Sive pro Tito, est socius meus et in vos adiutor; sive fratres nostri, apostoli ecclesiarum, gloria Christi.
2COR|8|24|Ostensionem ergo, quae est caritatis vestrae et nostrae gloriationis pro vobis, in illos ostendite in faciem ecclesiarum.
2COR|9|1|Nam de ministerio, quod fit in sanctos, superfluum est mihi scribere vobis;
2COR|9|2|scio enim promptum animum vestrum, pro quo de vobis glorior apud Macedonas, quoniam Achaia parata est ab anno praeterito, et vestra aemulatio provocavit plurimos.
2COR|9|3|Misi autem fratres, ut ne, quod gloriamur de vobis, evacuetur in hac parte, ut, quemadmodum dixi, parati sitis,
2COR|9|4|ne, cum venerint mecum Macedones et invenerint vos imparatos, erubescamus nos, ut non dicam vos, in hac substantia.
2COR|9|5|Necessarium ergo existimavi rogare fratres, ut praeveniant ad vos et praeparent repromissam benedictionem vestram, ut haec sit parata sic quasi benedictio, non quasi avaritia.
2COR|9|6|Hoc autem: qui parce seminat, parce et metet; et, qui seminat in benedictionibus, in benedictionibus et metet.
2COR|9|7|Unusquisque prout destinavit corde suo, non ex tristitia aut ex necessitate; hilarem enim datorem diligit Deus.
2COR|9|8|Potens est autem Deus omnem gratiam abundare facere in vobis, ut, in omnibus semper omnem sufficientiam habentes, abundetis in omne opus bonum,
2COR|9|9|sicut scriptum est: Dispersit, dedit pauperibus;iustitia eius manet in aeternum ".
2COR|9|10|Qui autem administrat semen seminanti, et panem ad manducandum praestabit et multiplicabit semen vestrum et augebit incrementa frugum iustitiae vestrae.
2COR|9|11|In omnibus locupletati in omnem simplicitatem, quae operatur per nos gratiarum actionem Deo
2COR|9|12|- quoniam ministerium huius officii non solum supplet ea, quae desunt sanctis, sed etiam abundat per multas gratiarum actiones Deo -
2COR|9|13|per probationem ministerii huius glorificantes Deum in oboedientia confessionis vestrae in evangelium Christi et simplicitate communionis in illos et in omnes,
2COR|9|14|et ipsorum obsecratione pro vobis, desiderantium vos propter eminentem gratiam Dei in vobis.
2COR|9|15|Gratias Deo super inenarrabili dono eius.
2COR|10|1|Ipse autem ego Paulus obse cro vos per mansuetudinem et modestiam Christi, qui in facie quidem humilis inter vos, absens autem confido in vobis;
2COR|10|2|rogo autem, ne praesens audeam per eam confidentiam, quae existimo audere in quosdam, qui arbitrantur nos tamquam secundum carnem ambulemus.
2COR|10|3|In carne enim ambulantes, non secundum carnem militamus
2COR|10|4|- nam arma militiae nostrae non carnalia sed potentia Deo ad destructionem munitionum - consilia destruentes
2COR|10|5|et omnem altitudinem extollentem se adversus scientiam Dei, et in captivitatem redigentes omnem intellectum in obsequium Christi,
2COR|10|6|et in promptu habentes ulcisci omnem inoboedientiam, cum impleta fuerit vestra oboedientia.
2COR|10|7|Quae secundum faciem sunt, videte. Si quis confidit sibi Christi se esse, hoc cogitet iterum apud se, quia sicut ipse Christi est, ita et nos.
2COR|10|8|Nam et si amplius aliquid gloriatus fuero de potestate nostra, quam dedit Dominus in aedificationem et non in destructionem vestram, non erubescam,
2COR|10|9|ut non existimer tamquam terrere vos per epistulas;
2COR|10|10|quoniam quidem " Epistulae - inquiunt - graves sunt et fortes, praesentia autem corporis infirma, et sermo contemptibilis ".
2COR|10|11|Hoc cogitet, qui eiusmodi est, quia quales sumus verbo per epistulas absentes, tales et praesentes in facto.
2COR|10|12|Non enim audemus inserere aut comparare nos quibusdam, qui seipsos commendant; sed ipsi se in semetipsis metientes et comparantes semetipsos sibi, non intellegunt.
2COR|10|13|Nos autem non ultra mensuram gloriabimur sed secundum mensuram regulae, quam impertitus est nobis Deus, mensuram pertingendi usque ad vos.
2COR|10|14|Non enim quasi non pertingentes ad vos superextendimus nosmetipsos, usque ad vos enim pervenimus in evangelio Christi;
2COR|10|15|non ultra mensuram gloriantes in alienis laboribus, spem autem habentes, crescente fide vestra, in vobis magnificari secundum regulam nostram in abundantiam,
2COR|10|16|ad evangelizandum in iis, quae ultra vos sunt, et non in aliena regula gloriari in his, quae praeparata sunt.
2COR|10|17|Qui autem gloriatur, in Domino glorietur;
2COR|10|18|non enim qui seipsum commendat, ille probatus est, sed quem Dominus commendat.
2COR|11|1|Utinam sustineretis modi cum quid insipientiae meae; sed et supportate me!
2COR|11|2|Aemulor enim vos Dei aemulatione; despondi enim vos uni viro virginem castam exhibere Christo.
2COR|11|3|Timeo autem, ne, sicut serpens Evam seduxit astutia sua, ita corrumpantur sensus vestri a simplicitate et castitate, quae est in Christum.
2COR|11|4|Nam si is qui venit, alium Christum praedicat, quem non praedicavimus, aut alium Spiritum accipitis, quem non accepistis, aut aliud evangelium, quod non recepistis, recte pateremini.
2COR|11|5|Existimo enim nihil me minus fecisse magnis apostolis;
2COR|11|6|nam etsi imperitus sermone, sed non scientia, in omni autem manifestantes in omnibus ad vos.
2COR|11|7|Aut numquid peccatum feci meipsum humilians, ut vos exaltemini, quoniam gratis evangelium Dei evangelizavi vobis?
2COR|11|8|Alias ecclesias exspoliavi accipiens stipendium ad ministerium vestrum
2COR|11|9|et, cum essem apud vos et egerem, nulli onerosus fui; nam, quod mihi deerat, suppleverunt fratres, qui venerunt a Macedonia; et in omnibus sine onere me vobis servavi et servabo.
2COR|11|10|Est veritas Christi in me, quoniam haec gloria non infringetur in me in regionibus Achaiae.
2COR|11|11|Quare? Quia non diligo vos? Deus scit!
2COR|11|12|Quod autem facio et faciam, ut amputem occasionem eorum, qui volunt occasionem, ut in quo gloriantur, inveniantur sicut et nos.
2COR|11|13|Nam eiusmodi pseudoapostoli, operarii subdoli, transfigurantes se in apostolos Christi.
2COR|11|14|Et non mirum, ipse enim Satanas transfigurat se in angelum lucis;
2COR|11|15|non est ergo magnum, si et ministri eius transfigurentur velut ministri iustitiae, quorum finis erit secundum opera ipsorum.
2COR|11|16|Iterum dico, ne quis me putet insipientem esse; alioquin velut insipientem accipite me, ut et ego modicum quid glorier.
2COR|11|17|Quod loquor, non loquor secundum Dominum, sed quasi in insipientia, in hac substantia gloriationis.
2COR|11|18|Quoniam multi gloriantur secundum carnem, et ego gloriabor.
2COR|11|19|Libenter enim suffertis insipientes, cum sitis ipsi sapientes;
2COR|11|20|sustinetis enim, si quis vos in servitutem redigit, si quis devorat, si quis accipit, si quis extollitur, si quis in faciem vos caedit.
2COR|11|21|Secundum ignobilitatem dico, quasi nos infirmi fuerimus; in quo quis audet, in insipientia dico, audeo et ego.
2COR|11|22|Hebraei sunt? Et ego. Israelitae sunt? Et ego. Semen Abrahae sunt? Et ego.
2COR|11|23|Ministri Christi sunt? Minus sapiens dico, plus ego: in laboribus plurimis, in carceribus abundantius, in plagis supra modum, in mortibus frequenter;
2COR|11|24|a Iudaeis quinquies quadragenas una minus accepi,
2COR|11|25|ter virgis caesus sum, semel lapidatus sum, ter naufragium feci, nocte et die in profundo maris fui;
2COR|11|26|in itineribus saepe, periculis fluminum, periculis latronum, periculis ex genere, periculis ex gentibus, periculis in civitate, periculis in solitudine, periculis in mari, periculis in falsis fratribus;
2COR|11|27|in labore et aerumna, in vigiliis saepe, in fame et siti, in ieiuniis frequenter, in frigore et nuditate;
2COR|11|28|praeter illa, quae extrinsecus sunt, instantia mea cotidiana, sollicitudo omnium ecclesiarum.
2COR|11|29|Quis infirmatur, et non infirmor? Quis scandalizatur, et ego non uror?
2COR|11|30|Si gloriari oportet, quae infirmitatis meae sunt, gloriabor.
2COR|11|31|Deus et Pater Domini Iesu scit, qui est benedictus in saecula, quod non mentior.
2COR|11|32|Damasci praepositus gentis Aretae regis custodiebat civitatem Damascenorum, ut me comprehenderet;
2COR|11|33|et per fenestram in sporta dimissus sum per murum et effugi manus eius.
2COR|12|1|Gloriari oportet; non expedit quidem, veniam autem ad visiones et revelationes Domini.
2COR|12|2|Scio hominem in Christo ante annos quattuordecim - sive in corpore nescio, sive extra corpus nescio, Deus scit - raptum eiusmodi usque ad tertium caelum.
2COR|12|3|Et scio huiusmodi hominem - sive in corpore sive extra corpus nescio, Deus scit -
2COR|12|4|quoniam raptus est in paradisum et audivit arcana verba, quae non licet homini loqui.
2COR|12|5|Pro eiusmodi gloriabor; pro me autem nihil gloriabor nisi in infirmitatibus meis.
2COR|12|6|Nam, et si voluero gloriari, non ero insipiens, veritatem enim dicam; parco autem, ne quis in me existimet supra id, quod videt me aut audit ex me,
2COR|12|7|et ex magnitudine revelationum. Propter quod, ne extollar, datus est mihi stimulus carni, angelus Satanae, ut me colaphizet, ne extollar.
2COR|12|8|Propter quod ter Dominum rogavi, ut discederet a me;
2COR|12|9|et dixit mihi: " Sufficit tibi gratia mea, nam virtus in infirmitate perficitur ". Libentissime igitur potius gloriabor in infirmitatibus meis, ut inhabitet in me virtus Christi.
2COR|12|10|Propter quod placeo mihi in infirmitatibus, in contumeliis, in necessitatibus, in persecutionibus et in angustiis, pro Christo; cum enim infirmor, tunc potens sum.
2COR|12|11|Factus sum insipiens. Vos me coegistis; ego enim debui a vobis commendari. Nihil enim minus fui ab his, qui sunt supra modum apostoli, tametsi nihil sum;
2COR|12|12|signa tamen apostoli facta sunt super vos in omni patientia, signis quoque et prodigiis et virtutibus.
2COR|12|13|Quid est enim quod minus habuistis prae ceteris ecclesiis, nisi quod ego ipse non gravavi vos? Donate mihi hanc iniuriam.
2COR|12|14|Ecce tertio hoc paratus sum venire ad vos et non ero gravis vobis; non enim quaero, quae vestra sunt, sed vos; nec enim debent filii parentibus thesaurizare, sed parentes filiis.
2COR|12|15|Ego autem libentissime impendam et superimpendar ipse pro animabus vestris. Si plus vos diligo, minus diligar?
2COR|12|16|Esto quidem, ego vos non gravavi; sed cum essem astutus, dolo vos cepi.
2COR|12|17|Numquid per aliquem eorum, quos misi ad vos, circumveni vos?
2COR|12|18|Rogavi Titum et misi cum illo fratrem; numquid Titus vos circumvenit? Nonne eodem spiritu ambulavimus? Nonne iisdem vestigiis?
2COR|12|19|Olim putatis quod excusemus nos apud vos? Coram Deo in Christo loquimur; omnia autem, carissimi, propter vestram aedificationem.
2COR|12|20|Timeo enim, ne forte, cum venero, non quales volo, inveniam vos, et ego inveniar a vobis, qualem non vultis; ne forte contentiones, aemulationes, animositates, dissensiones, detractiones, susurrationes, inflationes, seditiones sint;
2COR|12|21|ne iterum, cum venero, humiliet me Deus meus apud vos, et lugeam multos ex his, qui ante peccaverunt et non egerunt paenitentiam super immunditia et fornicatione et impudicitia, quam gesserunt.
2COR|13|1|Ecce tertio hoc venio ad vos; in ore duorum vel trium testium stabit omne verbum.
2COR|13|2|Praedixi et praedico, ut praesens bis et nunc absens his, qui ante peccaverunt, et ceteris omnibus, quoniam, si venero iterum, non parcam,
2COR|13|3|quoniam experimentum quaeritis eius, qui in me loquitur, Christi, qui in vos non infirmatur, sed potens est in vobis.
2COR|13|4|Nam etsi crucifixus est ex infirmitate, sed vivit ex virtute Dei. Nam et nos infirmi sumus in illo, sed vivemus cum eo ex virtute Dei in vos.
2COR|13|5|Vosmetipsos tentate, si estis in fide; ipsi vos probate. An non cognoscitis vos ipsos, quia Iesus Christus in vobis est? Nisi forte reprobi estis.
2COR|13|6|Spero autem quod cognoscetis quia nos non sumus reprobi.
2COR|13|7|Oramus autem Deum, ut nihil mali faciatis, non ut nos probati pareamus, sed ut vos, quod bonum est, faciatis, nos autem ut reprobi simus.
2COR|13|8|Non enim possumus aliquid adversus veritatem, sed pro veritate.
2COR|13|9|Gaudemus enim, quando nos infirmi sumus, vos autem potentes estis; hoc et oramus, vestram consummationem.
2COR|13|10|Ideo haec absens scribo, ut non praesens durius agam secundum potestatem, quam Dominus dedit mihi in aedificationem et non in destructionem.
2COR|13|11|De cetero, fratres, gaudete, perfecti estote, exhortamini invicem, idem sapite, pacem habete, et Deus dilectionis et pacis erit vobiscum.
2COR|13|12|Salutate invicem in osculo sancto. Salutant vos sancti omnes.
2COR|13|13|Gratia Domini Iesu Christi et caritas Dei et communicatio Sancti Spiritus cum omnibus vobis.
