LUKE|1|1|提阿非罗 大人哪，有好些人提笔作书，述说在我们中间所实现的事，是照传道的人从起初亲眼看见又传给我们的。这些事我从起头都详细考察了，我也想按着次序写给你，
LUKE|1|2|
LUKE|1|3|
LUKE|1|4|要让你知道所学的道都是确实的。
LUKE|1|5|在 希律 作 犹太 王的时候， 亚比雅 班里有一个祭司，名叫 撒迦利亚 ；他妻子是 亚伦 的后代，名叫 伊利莎白 。
LUKE|1|6|他们两人在上帝面前都是义人，遵行主的一切诫命和条例，没有可指责的。
LUKE|1|7|只是他们没有孩子，因为 伊利莎白 不生育，两个人又年纪老迈了。
LUKE|1|8|撒迦利亚 按班次在上帝面前执行祭司的职务，
LUKE|1|9|照祭司的规矩抽签，进到主的殿里烧香。
LUKE|1|10|烧香的时候，众百姓在外面祷告。
LUKE|1|11|有主的一个使者站在香坛的右边，向他显现。
LUKE|1|12|撒迦利亚 看见，就惊慌害怕。
LUKE|1|13|天使对他说：“ 撒迦利亚 ，不要害怕，因为你的祈祷已经被听见了。你的妻子 伊利莎白 要给你生一个儿子，你要给他起名叫 约翰 。
LUKE|1|14|你必欢喜快乐；有许多人因他出世也必喜乐。
LUKE|1|15|他在主面前将要为大，淡酒烈酒都不喝，从母腹里就被圣灵充满。
LUKE|1|16|他要使许多 以色列 人回转，归于主—他们的上帝。
LUKE|1|17|他将有 以利亚 的精神和能力，走在主的前面，叫父亲的心转向儿女，叫悖逆的人转向义人的智慧，又为主预备迎接他的百姓。”
LUKE|1|18|撒迦利亚 对天使说：“我怎么能知道这事呢？我已经老了，我的妻子也年纪老迈了。”
LUKE|1|19|天使回答他说：“我是站在上帝面前的 加百列 ，奉差遣来对你说话，把这好信息报给你。
LUKE|1|20|到了时候，这些话必然应验；只因你不信我的话，你会成为哑巴，不能说话，直到这些事实现的日子。”
LUKE|1|21|百姓等候 撒迦利亚 ，诧异他在圣所里迟延那么久。
LUKE|1|22|到他出来，却不能和他们说话，他们就知道他在圣所里见了异象；他直向他们打手势，因为他成了哑巴。
LUKE|1|23|他供职的日子一满，就回家去了。
LUKE|1|24|这些日子以后，他的妻子 伊利莎白 就怀孕，隐藏了五个月；
LUKE|1|25|她说：“主在眷顾我的日子，这样看顾我，要除掉我在人前的羞耻。”
LUKE|1|26|到了第六个月，天使 加百列 奉上帝的差遣往 加利利 的一座城去，这城名叫 拿撒勒 ，
LUKE|1|27|到一个童女那里，她已经许配 大卫 家的一个人，名叫 约瑟 ；童女的名字叫 马利亚 。
LUKE|1|28|天使进去，对她说：“蒙大恩的女子，你好，主和你同在！”
LUKE|1|29|马利亚 因这话就很惊慌，又反覆思考这样问候是什么意思。
LUKE|1|30|天使对她说： “ 马利亚 ，不要怕，你在上帝面前已经蒙恩了。
LUKE|1|31|你要怀孕生子，要给他起名叫耶稣。
LUKE|1|32|他将要为大，称为至高者的儿子； 主上帝要把他祖先 大卫 的王位给他。
LUKE|1|33|他要作 雅各 家的王，直到永远； 他的国没有穷尽。”
LUKE|1|34|马利亚 对天使说：“我没有出嫁，怎么会有这事呢？”
LUKE|1|35|天使回答她说： “圣灵要临到你身上； 至高者的能力要庇荫你， 因此，那要出生的圣者要称为上帝的儿子 。
LUKE|1|36|况且，你的亲戚 伊利莎白 ，就是那素来称为不生育的，在年老的时候也怀了男胎，现在怀孕六个月了。
LUKE|1|37|因为，出于上帝的话，没有一句不带能力的。”
LUKE|1|38|马利亚 说：“我是主的使女，愿意照你的话实现在我身上。”于是天使离开她去了。
LUKE|1|39|在那些日子， 马利亚 起身，急忙前往山区，来到 犹大 的一座城，
LUKE|1|40|进了 撒迦利亚 的家，向 伊利莎白 问安。
LUKE|1|41|伊利莎白 一听到 马利亚 问安，所怀的胎就在腹里跳动。 伊利莎白 被圣灵充满，
LUKE|1|42|高声喊着说： “你在妇女中是有福的！ 你所怀的胎也是有福的！
LUKE|1|43|我主的母亲到我这里来，为何这事临到我呢？
LUKE|1|44|因为你问安的声音一入我耳，我腹里的胎就欢喜跳动。
LUKE|1|45|这相信的女子是有福的！因为主对她所说的话都要应验。”
LUKE|1|46|马利亚 说： “我心尊主为大；
LUKE|1|47|我灵以上帝我的救主为乐；
LUKE|1|48|因为他顾念他使女的卑微； 从今以后，万代要称我有福。
LUKE|1|49|因为那有权能的为我做了大事； 他的名是圣的。
LUKE|1|50|他怜悯敬畏他的人， 直到世世代代。
LUKE|1|51|他用膀臂施展大能； 他赶散心里妄想的狂傲人。
LUKE|1|52|他叫有权柄的失位， 叫卑贱的升高。
LUKE|1|53|他叫饥饿的饱餐美食， 叫富足的空手回去。
LUKE|1|54|他扶助了他的仆人 以色列 ，不忘记施怜悯，
LUKE|1|55|正如他对我们的列祖说过， ‘怜悯 亚伯拉罕 和他的后裔，直到永远。’”
LUKE|1|56|马利亚 和 伊利莎白 同住，约有三个月，然后回家去了。
LUKE|1|57|伊利莎白 的产期到了，生了一个儿子。
LUKE|1|58|邻里亲属听见主向她大施怜悯，就和她一同欢乐。
LUKE|1|59|到了第八日，他们来给孩子行割礼，并要照他父亲的名字叫他 撒迦利亚 。
LUKE|1|60|他母亲回应说：“不！要叫他 约翰 。”
LUKE|1|61|他们对她说：“你亲族中没有叫这名字的。”
LUKE|1|62|他们就向他父亲打手势，问他这孩子要叫什么名字。
LUKE|1|63|他要了一块写字的板，写上：“他的名字是 约翰 。”他们就都惊讶。
LUKE|1|64|撒迦利亚 的口立刻开了，舌头也松了，就开始说话称颂上帝。
LUKE|1|65|周围居住的人都惧怕；这一切的事就传遍了 犹太 山区。
LUKE|1|66|凡听见的人都把这事放在心里，他们说：“这个孩子将来会怎么样呢？”因为有主的手与他同在。
LUKE|1|67|他父亲 撒迦利亚 被圣灵充满，就预言说：
LUKE|1|68|“主— 以色列 的上帝是应当称颂的！ 因他眷顾他的百姓，为他们施行救赎，
LUKE|1|69|在他仆人 大卫 家中， 为我们兴起了拯救的角，
LUKE|1|70|正如主藉着古时候圣先知的口所说的，
LUKE|1|71|‘他拯救我们脱离仇敌， 脱离一切恨我们之人的手。
LUKE|1|72|他向我们列祖施怜悯， 记得他的圣约，
LUKE|1|73|就是他对我们祖宗 亚伯拉罕 所起的誓，
LUKE|1|74|叫我们既从仇敌手中被救出来， 就可以终身在他面前， 无所惧怕地用圣洁和公义事奉他。
LUKE|1|75|
LUKE|1|76|孩子啊，你要称为至高者的先知； 因为你要走在主的前面，为他预备道路，
LUKE|1|77|叫他的百姓因罪得赦， 认识救恩；
LUKE|1|78|因我们上帝怜悯的心肠， 叫清晨的日光从高天临到我们，
LUKE|1|79|要照亮坐在黑暗中死荫里的人， 把我们的脚引到和平的路上。’”
LUKE|1|80|这孩子渐渐长大，心灵坚强，住在旷野，直到他在 以色列 人面前公开出现的日子。
LUKE|2|1|在那些日子，凯撒 奥古斯都 降旨，叫全国人民都登记户籍。
LUKE|2|2|这第一次登记户籍是在 居里扭 作 叙利亚 总督的时候行的。
LUKE|2|3|众人各归各城，办理登记。
LUKE|2|4|约瑟 也从 加利利 的 拿撒勒城 上 犹太 去，到了 大卫 的城名叫 伯利恒 ，因为他是 大卫 家族的人，
LUKE|2|5|要和他所聘之妻 马利亚 一同登记户籍。那时 马利亚 已经怀孕。
LUKE|2|6|他们在那里的时候， 马利亚 的产期到了，
LUKE|2|7|就生了头胎的儿子，用布包起来，放在马槽里，因为客店里没有地方。
LUKE|2|8|在 伯利恒 的野外有牧羊人，夜间值班看守羊群。
LUKE|2|9|有主的一个使者站在他们旁边，主的荣光四面照着他们，牧羊人就很惧怕。
LUKE|2|10|那天使对他们说：“不要惧怕！看哪！因为我报给你们大喜的信息，是关乎万民的：
LUKE|2|11|因今天在 大卫 的城里，为你们生了救主，就是主基督。
LUKE|2|12|你们要看见一个婴孩，包着布，卧在马槽里，那就是给你们的记号。”
LUKE|2|13|忽然，有一大队天兵同那天使赞美上帝说：
LUKE|2|14|“在至高之处荣耀归与上帝！ 在地上平安归与他所喜悦的人！”
LUKE|2|15|众天使离开他们，升天去了。牧羊人彼此说：“我们往 伯利恒 去，看看所成的事，就是主所告诉我们的。”
LUKE|2|16|他们急忙去了，找到 马利亚 和 约瑟 ，还有那婴孩卧在马槽里。
LUKE|2|17|他们看见，就把天使论这孩子的话传开了。
LUKE|2|18|听见的人都诧异牧羊人对他们所说的话。
LUKE|2|19|马利亚 却把这一切的事存在心里，反覆思考。
LUKE|2|20|牧羊人回去了，因所听见所看见的一切事，正如天使向他们所说的，就归荣耀于上帝，赞美他。
LUKE|2|21|满了八天，他们就给孩子行割礼，又给他起名叫耶稣；这是他还没有在母腹里成胎以前天使所起的名。
LUKE|2|22|按 摩西 律法满了洁净的日子，他们就带着孩子上 耶路撒冷 去，要把他献给主。
LUKE|2|23|正如主的律法上所记：“凡头生的男子必归主为圣”；
LUKE|2|24|又要照主的律法上所说，用一对斑鸠，或用两只雏鸽献祭。
LUKE|2|25|那时，在 耶路撒冷 有一个人，名叫 西面 ；这人又公义又虔诚，素常盼望 以色列 的安慰者来到，又有圣灵在他身上。
LUKE|2|26|他得了圣灵的启示，知道自己未死以前必看见主所立的基督。
LUKE|2|27|他受了圣灵的感动，进入圣殿，正遇见耶稣的父母抱着孩子进来，要照律法的规矩而行。
LUKE|2|28|西面 就把他抱过来，称颂上帝说：
LUKE|2|29|“主啊，如今可以照你的话， 容你的仆人安然去世；
LUKE|2|30|因为我的眼睛已经看见你的救恩，
LUKE|2|31|就是你在万民面前所预备的：
LUKE|2|32|是启示外邦人的光， 是你民 以色列 的荣耀。”
LUKE|2|33|孩子的父母因论耶稣的这些话就惊讶。
LUKE|2|34|西面 给他们祝福，又对孩子的母亲 马利亚 说：“这孩子被立，是要叫 以色列 中许多人跌倒，许多人兴起；又要成为毁谤的对象，
LUKE|2|35|叫许多人心里的意念显露出来；你自己的心也要被剑刺透。”
LUKE|2|36|又有位女先知，名叫 亚拿 ，是 亚设 支派 法内力 的女儿，年纪已经老迈，从童女出嫁，同丈夫住了七年，
LUKE|2|37|就寡居了，现在已经八十四岁 。她不离开圣殿，禁食祈求，昼夜事奉上帝。
LUKE|2|38|正当那时，她进前来感谢上帝，对一切盼望 耶路撒冷 得救赎的人讲论这孩子的事。
LUKE|2|39|约瑟 和 马利亚 照主的律法办完了一切的事，就回 加利利 ，到自己的城 拿撒勒 去了。
LUKE|2|40|孩子渐渐长大，强健起来，充满智慧，又有上帝的恩典在他身上。
LUKE|2|41|每年逾越节，他父母都上 耶路撒冷 去。
LUKE|2|42|当他十二岁的时候，他们按着过节的规矩上去。
LUKE|2|43|守满了节期，他们回去，孩童耶稣仍旧在 耶路撒冷 。他的父母并不知道，
LUKE|2|44|以为他在同行的人中间，走了一天的路程才在亲属和熟悉的人中找他，
LUKE|2|45|既找不着，就回 耶路撒冷 去找他。
LUKE|2|46|过了三天，他们发现他在圣殿里，坐在教师中间，一面听，一面问。
LUKE|2|47|凡听见他的人都对他的聪明和应对感到惊奇。
LUKE|2|48|他父母看见就很惊奇。他母亲对他说：“我儿啊，为什么对我们这样做呢？看哪，你父亲和我很焦急，到处找你！”
LUKE|2|49|耶稣对他们说：“为什么找我呢？难道你们不知道我应当在我父的家里吗？ ”
LUKE|2|50|他所说的这话，他们不明白。
LUKE|2|51|他就同他们下去，回到 拿撒勒 ，并且顺从他们。他母亲把这一切的事都存在心里。
LUKE|2|52|耶稣的智慧和身量 ，并上帝和人喜爱他的心，都一齐增长。
LUKE|3|1|凯撒 提庇留 在位第十五年， 本丢．彼拉多 作 犹太 总督， 希律 作 加利利 分封的王，他兄弟 腓力 作 以土利亚 和 特拉可尼 地区分封的王， 吕撒聂 作 亚比利尼 分封的王，
LUKE|3|2|亚那 和 该亚法 作大祭司。那时， 撒迦利亚 的儿子 约翰 在旷野里，上帝的话临到他。
LUKE|3|3|他就走遍 约旦河 一带地方，宣讲悔改的洗礼，使罪得赦。
LUKE|3|4|正如 以赛亚 先知书上所记的话： “在旷野有声音呼喊着： 预备主的道， 修直他的路！
LUKE|3|5|一切山洼都要填满； 大小山冈都要削平！ 弯弯曲曲的地方要改为笔直； 高高低低的道路要改为平坦！
LUKE|3|6|凡血肉之躯的，都要看见上帝的救恩！”
LUKE|3|7|约翰 对那出来要受他洗的众人说：“毒蛇的孽种啊，谁指示你们逃避那将要来的愤怒呢？
LUKE|3|8|你们要结出果子来，和悔改的心相称。不要自己心里说：‘我们有 亚伯拉罕 为祖宗。’我告诉你们，上帝能从这些石头中给 亚伯拉罕 兴起子孙来。
LUKE|3|9|现在斧子已经放在树根上，凡不结好果子的树就砍下来，丢在火里。”
LUKE|3|10|众人问他：“这样，我们该做什么呢？”
LUKE|3|11|约翰 回答：“有两件衣裳的，就分给那没有的；有食物的，也该这样做。”
LUKE|3|12|也有税吏来要受洗，对他说：“老师，我们该做什么呢？”
LUKE|3|13|约翰 对他们说：“除了规定的数目，不要多收。”
LUKE|3|14|也有士兵问他说：“我们该做什么呢？” 约翰 说：“不要勒索任何人，也不要敲诈人；自己有粮饷就该知足。”
LUKE|3|15|百姓期待基督的来临；他们心里猜测，或许 约翰 是基督。
LUKE|3|16|约翰 对众人说：“我是用水给你们施洗，但有一位能力比我更大的要来，我就是给他解鞋带也不配。他要用圣灵与火给你们施洗。
LUKE|3|17|他手里拿着簸箕，要扬净他的谷物，把麦子收在仓里，把糠用不灭的火烧尽。”
LUKE|3|18|约翰 又用许多别的话劝百姓，向他们传福音。
LUKE|3|19|希律 分封王，因他兄弟之妻 希罗底 的缘故，并因他所做的一切恶事，受了 约翰 的责备。
LUKE|3|20|希律 在一切事上又添了这一件，就是把 约翰 收在监里。
LUKE|3|21|众百姓都受了洗，耶稣也受了洗。他正祷告的时候，天开了，
LUKE|3|22|圣灵降在他身上，形状仿佛鸽子；又有声音从天上来，说：“你是我的爱子，我喜爱你。”
LUKE|3|23|耶稣开始传道，年纪约有三十岁。依人看来，他是 约瑟 的儿子， 约瑟 是 希里 的儿子，
LUKE|3|24|希里 是 玛塔 的儿子， 玛塔 是 利未 的儿子， 利未 是 麦基 的儿子， 麦基 是 雅拿 的儿子， 雅拿 是 约瑟 的儿子，
LUKE|3|25|约瑟 是 玛他提亚 的儿子， 玛他提亚 是 亚摩斯 的儿子， 亚摩斯 是 拿鸿 的儿子， 拿鸿 是 以斯利 的儿子， 以斯利 是 拿该 的儿子，
LUKE|3|26|拿该 是 玛押 的儿子， 玛押 是 玛他提亚 的儿子， 玛他提亚 是 西美 的儿子， 西美 是 约瑟 的儿子， 约瑟 是 犹大 的儿子， 犹大 是 约亚拿 的儿子，
LUKE|3|27|约亚拿 是 利撒 的儿子， 利撒 是 所罗巴伯 的儿子， 所罗巴伯 是 撒拉铁 的儿子， 撒拉铁 是 尼利 的儿子， 尼利 是 麦基 的儿子，
LUKE|3|28|麦基 是 亚底 的儿子， 亚底 是 哥桑 的儿子， 哥桑 是 以摩当 的儿子， 以摩当 是 珥 的儿子， 珥 是 约细 的儿子，
LUKE|3|29|约细 是 以利以谢 的儿子， 以利以谢 是 约令 的儿子， 约令 是 玛塔 的儿子， 玛塔 是 利未 的儿子，
LUKE|3|30|利未 是 西缅 的儿子， 西缅 是 犹大 的儿子， 犹大 是 约瑟 的儿子， 约瑟 是 约南 的儿子， 约南 是 以利亚敬 的儿子，
LUKE|3|31|以利亚敬 是 米利亚 的儿子， 米利亚 是 买南 的儿子， 买南 是 玛达他 的儿子， 玛达他 是 拿单 的儿子， 拿单 是 大卫 的儿子，
LUKE|3|32|大卫 是 耶西 的儿子， 耶西 是 俄备得 的儿子， 俄备得 是 波阿斯 的儿子， 波阿斯 是 沙拉 的儿子， 沙拉 是 拿顺 的儿子 ，
LUKE|3|33|拿顺 是 亚米拿达 的儿子， 亚米拿达 是 亚民 的儿子， 亚民 是 亚尼 的儿子， 亚尼 是 希斯仑 的儿子 ， 希斯仑 是 法勒斯 的儿子， 法勒斯 是 犹大 的儿子，
LUKE|3|34|犹大 是 雅各 的儿子， 雅各 是 以撒 的儿子， 以撒 是 亚伯拉罕 的儿子， 亚伯拉罕 是 他拉 的儿子， 他拉 是 拿鹤 的儿子，
LUKE|3|35|拿鹤 是 西鹿 的儿子， 西鹿 是 拉吴 的儿子， 拉吴 是 法勒 的儿子， 法勒 是 希伯 的儿子， 希伯 是 沙拉 的儿子，
LUKE|3|36|沙拉 是 该南 的儿子， 该南 是 亚法撒 的儿子， 亚法撒 是 闪 的儿子， 闪 是 挪亚 的儿子， 挪亚 是 拉麦 的儿子，
LUKE|3|37|拉麦 是 玛土撒拉 的儿子， 玛土撒拉 是 以诺 的儿子， 以诺 是 雅列 的儿子， 雅列 是 玛勒列 的儿子， 玛勒列 是 该南 的儿子， 该南 是 以挪士 的儿子，
LUKE|3|38|以挪士 是 塞特 的儿子， 塞特 是 亚当 的儿子， 亚当 是上帝的儿子。
LUKE|4|1|耶稣满有圣灵，从 约旦河 回来，圣灵把他引到旷野，
LUKE|4|2|四十天受魔鬼的试探。在那些日子，他没有吃什么，日子满了，他饿了。
LUKE|4|3|魔鬼对他说：“你若是上帝的儿子，叫这块石头变成食物吧。”
LUKE|4|4|耶稣回答：“经上记着： ‘人活着，不是单靠食物。 ’”
LUKE|4|5|魔鬼又领他上了高山，霎时间把天下万国都指给他看，
LUKE|4|6|对他说：“这一切权柄和荣华我都要给你，因为这原是交给我的，我愿意给谁就给谁。
LUKE|4|7|你若在我面前下拜，这一切都归你。”
LUKE|4|8|耶稣回答他说：“经上记着： ‘要拜主—你的上帝， 惟独事奉他。’”
LUKE|4|9|魔鬼又领他到 耶路撒冷 去，叫他站在圣殿顶上，对他说：“你若是上帝的儿子，从这里跳下去！
LUKE|4|10|因为经上记着： ‘主要为你命令他的使者保护你；
LUKE|4|11|他们要用手托住你， 免得你的脚碰在石头上。’”
LUKE|4|12|耶稣回答他说：“经上说：‘不可试探主—你的上帝。’”
LUKE|4|13|魔鬼用完了各样的试探，就离开耶稣，再等时机。
LUKE|4|14|耶稣带着圣灵的能力回到 加利利 ，他的名声传遍了四方。
LUKE|4|15|他在各会堂里教导人，众人都称赞他。
LUKE|4|16|耶稣来到 拿撒勒 ，就是他长大的地方。在安息日，照他素常的规矩进了会堂，站起来要念圣经。
LUKE|4|17|有人把 以赛亚 先知的书交给他，他就打开，找到一处写着：
LUKE|4|18|“主的灵在我身上， 因为他用膏膏我， 叫我传福音给贫穷的人； 差遣我宣告： 被掳的得释放， 失明的得看见， 受压迫的得自由，
LUKE|4|19|宣告上帝悦纳人的禧年。”
LUKE|4|20|于是他把书卷起来，交还给管理人，就坐下。会堂里的人都定睛看他。
LUKE|4|21|耶稣对他们说：“你们听见的这段经文，今天已经应验了。”
LUKE|4|22|众人都称赞他，并对他口中所出的恩言感到惊讶；他们说：“这不是 约瑟 的儿子吗？”
LUKE|4|23|耶稣对他们说：“你们一定会用这俗语向我说：‘医生，你医治自己吧！我们听见你在 迦百农 所做的事，也该在你自己的家乡做吧。’”
LUKE|4|24|他又说：“我实在告诉你们，没有先知在自己家乡被人接纳的。
LUKE|4|25|我对你们说实话，在 以利亚 的时候，天闭塞了三年六个月，遍地有大饥荒，那时， 以色列 中有许多寡妇，
LUKE|4|26|以利亚 并没有奉差往她们中任何一个人那里去，只奉差往 西顿 的 撒勒法 一个寡妇那里去。
LUKE|4|27|在 以利沙 先知的时候， 以色列 中有许多痲疯病人，但除了 叙利亚 的 乃缦 ，没有一个得洁净的。”
LUKE|4|28|会堂里的人听见这些话，都怒气填胸，
LUKE|4|29|就起来赶他出城。他们的城造在山上；他们带他到山崖，要把他推下去。
LUKE|4|30|他却从他们中间穿过去，走了。
LUKE|4|31|耶稣下到 迦百农 ，就是 加利利 的一座城，在安息日教导众人。
LUKE|4|32|他们对他的教导感到很惊奇，因为他的话里有权柄。
LUKE|4|33|在会堂里有一个人，被污鬼的灵附着，大声喊叫说：
LUKE|4|34|“唉！ 拿撒勒 人耶稣，你为什么干扰我们？你来消灭我们吗？我知道你是谁，你是上帝的圣者。”
LUKE|4|35|耶稣斥责他说：“不要作声，从这人身上出来吧！”鬼把那人摔倒在众人中间，就出来了，却没有伤害他。
LUKE|4|36|众人都惊讶，彼此对问：“这是什么道理呢？因为他用权柄能力命令污灵，污灵就出来。”
LUKE|4|37|于是耶稣的名声传遍了周围各地。
LUKE|4|38|耶稣出了会堂，进了 西门 的家。 西门 的岳母在发高烧，有些人为她求耶稣。
LUKE|4|39|耶稣站在她旁边，斥责那高烧，烧就退了。她立刻起来服事他们。
LUKE|4|40|日落的时候，凡有病人的，不论害什么病，都带到耶稣那里。耶稣给他们每一个人按手，治好他们。
LUKE|4|41|又有鬼从好些人身上出来，喊着说：“你是上帝的儿子！”耶稣斥责他们，不许他们说话，因为他们知道他是基督。
LUKE|4|42|天亮的时候，耶稣出来，走到荒野的地方。众人去找他，到了他那里，要留住他，不让他离开他们。
LUKE|4|43|但耶稣对他们说：“我也必须在别的城传上帝国的福音，因我奉差原是为此。”
LUKE|4|44|于是耶稣在 犹太 的各会堂传道。
LUKE|5|1|耶稣站在 革尼撒勒 湖边，众人拥挤他，要听上帝的道。
LUKE|5|2|他见有两只船靠在湖边，打鱼的人却离开船，洗网去了。
LUKE|5|3|有一只船是 西门 的，耶稣就上去，请他把船撑开，稍微离岸，就坐下，在船上教导众人。
LUKE|5|4|他讲完了，对 西门 说：“把船开到水深的地方下网打鱼。”
LUKE|5|5|西门 说：“老师，我们整夜劳累，并没有打着什么。但依从你的话，我就下网。”
LUKE|5|6|他们下了网，圈住许多鱼，网险些裂开，
LUKE|5|7|就招手叫另一只船上的同伴来帮助。他们就来，把鱼装满了两只船，船甚至要沉下去。
LUKE|5|8|西门．彼得 看见，就俯伏在耶稣膝前，说：“主啊，离开我，我是个罪人。”
LUKE|5|9|他和一切跟他一起的人对打到了这一网的鱼都很惊讶。
LUKE|5|10|他的伙伴 西庇太 的儿子 雅各 、 约翰 ，也是这样。耶稣对 西门 说：“不要怕！从今以后，你要得人了。”
LUKE|5|11|他们把两只船靠了岸，就撇下所有的，跟从了耶稣。
LUKE|5|12|有一回，耶稣在一个城里，有人满身长了痲疯，看见他，就俯伏在地，求他说：“主啊，你若肯，你能使我洁净。”
LUKE|5|13|耶稣伸手摸他，说：“我肯，你洁净了吧！”痲疯病立刻离开了他。
LUKE|5|14|耶稣吩咐他：“你不可告诉任何人，只要去，把自己给祭司察看，又因为你已经洁净，要照 摩西 所吩咐的献上祭物，作为证据给众人看。”
LUKE|5|15|但耶稣的名声越发传扬出去。有一大群人聚集来听道，也希望耶稣医治他们的病。
LUKE|5|16|耶稣却退到旷野去祷告。
LUKE|5|17|有一天，耶稣教导人，有法利赛人和律法教师在旁边坐着；他们是从 加利利 各乡村、 犹太 和 耶路撒冷 来的。主的能力与耶稣同在，使他能治好病人。
LUKE|5|18|这时，有些人用褥子抬着一个瘫子，要把他抬进去放在耶稣面前，
LUKE|5|19|却因人多，找不出法子抬进去，就上了房顶，从瓦间把他连褥子缒到当中，在耶稣面前。
LUKE|5|20|耶稣见他们的信心，就说：“朋友，你的罪赦了。”
LUKE|5|21|文士和法利赛人就开始议论说：“这个人是谁，竟说亵渎的话？除了上帝一位之外，谁能赦罪呢？”
LUKE|5|22|耶稣知道他们所议论的，就回答他们说：“你们心里为什么议论呢？
LUKE|5|23|说‘你的罪赦了’，或说‘你起来行走’，哪一样容易呢？
LUKE|5|24|但要让你们知道，人子在地上有赦罪的权柄。”他就对瘫子说：“我吩咐你，起来！拿你的褥子回家去吧。”
LUKE|5|25|那人当着众人面前立刻起来，拿了他所躺卧的褥子回家去，归荣耀给上帝。
LUKE|5|26|众人都惊奇，也归荣耀给上帝，并且满心惧怕，说：“我们今日看见不寻常的事了！”
LUKE|5|27|这些事以后，耶稣出去，看见一个税吏，名叫 利未 ，在税关坐着，就对他说：“来跟从我！”
LUKE|5|28|他就撇下所有的，起来跟从耶稣。
LUKE|5|29|利未 在自己家里为耶稣大摆宴席，有一大群税吏和别的人与他们一同坐席。
LUKE|5|30|法利赛人和文士就向耶稣的门徒发怨言说：“你们为什么跟税吏和罪人一同吃喝呢？”
LUKE|5|31|耶稣回答他们：“健康的人用不着医生；有病的人才用得着。
LUKE|5|32|我不是来召义人悔改，而是召罪人悔改。”
LUKE|5|33|他们对耶稣说：“ 约翰 的门徒常常禁食祈祷，法利赛人的门徒也是这样，惟独跟你在一起的又吃又喝。”
LUKE|5|34|耶稣对他们说：“新郎和宾客在一起的时候，你们怎么能叫宾客禁食呢？
LUKE|5|35|但日子将到，新郎要被带走，那些日子他们就要禁食了。”
LUKE|5|36|耶稣又讲一个比喻，对他们说：“没有人把新衣服撕下一块来补在旧衣服上，若是这样，会把新的撕裂了，并且所撕下来的那块新的和旧的也不相称。
LUKE|5|37|也没有人把新酒装在旧皮袋里；若是这样，新酒会胀破皮袋，酒就漏出来，皮袋也糟蹋了。
LUKE|5|38|相反地，新酒必须装在新皮袋里。
LUKE|5|39|没有人喝了陈酒又想喝新的；他总说陈的好。”
LUKE|6|1|有一个安息日 ，耶稣从麦田经过。他的门徒摘了麦穗，用手搓着吃。
LUKE|6|2|有几个法利赛人说：“你们为什么做安息日不合法的事呢？”
LUKE|6|3|耶稣回答他们：“ 大卫 和跟从他的人饥饿时所做的事，你们没有念过吗？
LUKE|6|4|他怎么进了上帝的居所，拿供饼吃，又给跟从的人吃呢？这饼惟独祭司可以吃，别人都不可以吃。”
LUKE|6|5|他又对他们说：“人子是安息日的主。”
LUKE|6|6|又有一个安息日，耶稣进了会堂教导人，在那里有一个人，他的右手萎缩了。
LUKE|6|7|文士和法利赛人窥探耶稣会不会在安息日治病，为要找把柄告他。
LUKE|6|8|耶稣却知道他们的意念，就对那萎缩了手的人说：“起来，站在当中！”那人就起来，站着。
LUKE|6|9|耶稣对他们说：“我问你们，在安息日行善行恶，救命害命，哪样是合法的呢？”
LUKE|6|10|他就环视众人，对那人说：“伸出手来！”他照着做，他的手就复原了。
LUKE|6|11|他们怒气填胸，彼此商议怎样对付耶稣。
LUKE|6|12|在那些日子，耶稣出去，上山祈祷，整夜向上帝祷告。
LUKE|6|13|到了天亮，他叫门徒来，就从他们中间挑选十二个人，称他们为使徒。
LUKE|6|14|这十二个人有 西门 （耶稣又给他起名叫 彼得 ），还有他弟弟 安得烈 ，又有 雅各 和 约翰 ， 腓力 和 巴多罗买 ，
LUKE|6|15|马太 和 多马 ， 亚勒腓 的儿子 雅各 和激进党的 西门 ，
LUKE|6|16|雅各 的儿子 犹大 和后来成为出卖者的 加略 人 犹大 。
LUKE|6|17|耶稣和他们下了山，站在一块平地上；在一起的有许多门徒，又有许多百姓从全 犹太 和 耶路撒冷 ，并 推罗 、 西顿 的海边来，
LUKE|6|18|都要听他讲道，又希望耶稣医治他们的病；还有被污灵缠磨的，也得了医治。
LUKE|6|19|众人都想要摸他，因为有能力从他身上发出来，治好了他们。
LUKE|6|20|耶稣举目看着门徒，说： “贫穷的人有福了！ 因为上帝的国是你们的。
LUKE|6|21|现在饥饿的人有福了！ 因为你们将得饱足。 现在哭泣的人有福了！ 因为你们将要欢笑。
LUKE|6|22|人为人子的缘故憎恨你们，拒绝你们，辱骂你们，把你们当恶人除掉你们的名，你们就有福了！
LUKE|6|23|在那日，你们要欢欣雀跃，因为你们在天上的赏赐是很多的；他们的祖宗也是这样待先知的。
LUKE|6|24|但你们富足的人有祸了！ 因为你们已经受过安慰。
LUKE|6|25|你们现在饱足的人有祸了！ 因为你们将要饥饿。 你们现在欢笑的人有祸了！ 因为你们将要哀恸哭泣。
LUKE|6|26|人都说你们好的时候，你们有祸了！因为他们的祖宗也是这样待假先知的。”
LUKE|6|27|“可是我告诉你们这些听的人，要爱你们的仇敌！要善待恨你们的人！
LUKE|6|28|要祝福诅咒你们的人！要为凌辱你们的人祷告！
LUKE|6|29|有人打你的脸，连另一边也由他打。有人拿你的外衣，连内衣也由他拿去。
LUKE|6|30|凡求你的，就给他；有人拿走你的东西，不要讨回来。
LUKE|6|31|“你们想要人怎样待你们，你们也要怎样待人。
LUKE|6|32|你们若只爱那爱你们的人，有什么可感谢的呢？就是罪人也爱那爱他们的人。
LUKE|6|33|你们若善待那善待你们的人，有什么可感谢的呢？就是罪人也是这样做。
LUKE|6|34|你们若借给人，希望从他收回，有什么可感谢的呢？就是罪人也借给罪人，再如数收回。
LUKE|6|35|你们倒要爱仇敌，要善待他们，并要借给人不指望偿还，你们的赏赐就很多了，你们必作至高者的儿子，因为他恩待那忘恩的和作恶的。
LUKE|6|36|你们要仁慈，像你们的父是仁慈的。”
LUKE|6|37|“你们不要评断别人，就不被审判；你们不要定人的罪，就不被定罪；你们要饶恕人，就必蒙饶恕。
LUKE|6|38|你们要给人，就必有给你们的，并且用十足的升斗，连摇带按，上尖下流地倒在你们怀里；因为你们用什么量器量给人，也必用什么量器量给你们。”
LUKE|6|39|耶稣又用比喻对他们说：“瞎子岂能领瞎子，两个人不是都要掉在坑里吗？
LUKE|6|40|学生不高过老师，凡学成了的会和老师一样。
LUKE|6|41|为什么看见你弟兄眼中有刺，却不想自己眼中有梁木呢？
LUKE|6|42|你不见自己眼中有梁木，怎能对你弟兄说：‘让我去掉你眼中的刺’呢？你这假冒为善的人！先去掉自己眼中的梁木，然后才能看得清楚，好去掉你弟兄眼中的刺。”
LUKE|6|43|“没有好树结坏果子，也没有坏树结好果子。
LUKE|6|44|每一种树木可以从其果子看出来。人不是从荆棘上摘无花果的，也不是从蒺藜里摘葡萄的。
LUKE|6|45|善人从他心里所存的善发出善来，恶人从他所存的恶发出恶来；因为心里所充满的，口里就说出来。”
LUKE|6|46|“你们为什么称呼我‘主啊，主啊’，却不照我的话做呢？
LUKE|6|47|凡到我这里来，听了我的话又去做的，我要告诉你们他像什么人：
LUKE|6|48|他像一个人盖房子，把地挖深，将根基立在磐石上，到发大水的时候，水冲那房子，房子总不动摇，因为盖造得好。
LUKE|6|49|但听了不去做的，就像一个人在土地上盖房子，没有根基，水一冲，立刻倒塌了，并且那房子损坏得很厉害。”
LUKE|7|1|耶稣对百姓讲完了这一切的话，就进了 迦百农 。
LUKE|7|2|有一个百夫长所器重的仆人害病，快要死了。
LUKE|7|3|百夫长风闻耶稣的事，就托 犹太 人的几个长老去求耶稣来救他的仆人。
LUKE|7|4|他们到了耶稣那里，切切地求他说：“你为他做这事是他配得的；
LUKE|7|5|因为他爱我们的民族，为我们建造会堂。”
LUKE|7|6|耶稣就和他们同去。离那家不远，百夫长托几个朋友去见耶稣，对他说：“主啊，不必劳驾，因你到舍下来，我不敢当。
LUKE|7|7|我也自以为不配去见你，只要你说一句话，就会让我的僮仆得痊愈。
LUKE|7|8|因为我被派在人的权下，也有兵在我之下。我对这个说：‘去！’他就去；对那个说：‘来！’他就来；对我的仆人说：‘做这事！’他就去做。”
LUKE|7|9|耶稣听到这些话，就很惊讶，转身对跟随的众人说：“我告诉你们，这么大的信心，就是在 以色列 ，我也没有见过。”
LUKE|7|10|那差来的人回到百夫长家里，发现仆人已经好了。
LUKE|7|11|过了不久 ，耶稣往一座城去，这城名叫 拿因 ，他的门徒和一大群人与他同行。
LUKE|7|12|当他走近城门时，有一个死人被抬出来。这人是他母亲独生的儿子，而他母亲又是寡妇。城里的许多人与她一同送殡。
LUKE|7|13|主看见那寡妇就怜悯她，对她说：“不要哭。”
LUKE|7|14|于是耶稣进前来，按着杠，抬的人就站住了。耶稣说：“年轻人，我吩咐你，起来！”
LUKE|7|15|那死人就坐了起来，开始说话，耶稣就把他交给他的母亲。
LUKE|7|16|众人都惊奇，归荣耀给上帝，说：“有大先知在我们当中兴起了！”又说：“上帝眷顾了他的百姓！”
LUKE|7|17|关于耶稣的这事就传遍了 犹太 和周围地区。
LUKE|7|18|约翰 的门徒把这些事都告诉 约翰 。于是 约翰 叫了两个门徒来，
LUKE|7|19|差他们到主 那里去，说：“将要来的那位就是你吗？还是我们要等候别人呢？”
LUKE|7|20|那两个人来到耶稣那里，说：“施洗的 约翰 差我们来问你：‘将要来的那位就是你吗？还是我们要等候别人呢？’”
LUKE|7|21|就在那时，耶稣治好了许多患疾病的，得瘟疫的，被邪灵附身的，又开恩使好些盲人能看见。
LUKE|7|22|耶稣回答他们：“你们去，把所看见、所听见的告诉 约翰 ：就是盲人看见，瘸子行走，痲疯病人得洁净，聋子听见，死人复活，穷人听到福音。
LUKE|7|23|凡不因我跌倒的有福了！”
LUKE|7|24|约翰 所差来的人一走，耶稣就对众人谈到 约翰 ，说：“你们从前到旷野去，是要看什么呢？被吹动的芦苇吗？
LUKE|7|25|你们出去到底是要看什么？穿细软衣服的人吗？看哪，那穿华丽衣服、宴乐度日的人是在王宫里。
LUKE|7|26|你们出去究竟是要看什么？是先知吗？是的，我告诉你们，他比先知大多了。
LUKE|7|27|这个人就是经上所说的： ‘看哪，我要差遣我的使者在你面前， 他要在你前面为你预备道路。’
LUKE|7|28|我告诉你们，凡女子所生的，没有比 约翰 大的；但在上帝国里，最小的比他还大。”
LUKE|7|29|众百姓和税吏已受过 约翰 的洗，听见这话，就以上帝为义；
LUKE|7|30|但法利赛人和律法师没有受过 约翰 的洗，竟废弃了上帝为他们所定的旨意。
LUKE|7|31|主又说：“这样，我该用什么来比这世代的人呢？他们好像什么呢？
LUKE|7|32|这正像孩童坐在街市上，彼此喊叫： ‘我们为你们吹笛，你们不跳舞； 我们唱哀歌，你们不啼哭。’
LUKE|7|33|施洗的 约翰 来，不吃饼，不喝酒，你们说他是被鬼附的。
LUKE|7|34|人子来，也吃也喝，你们又说这人贪食好酒，是税吏和罪人的朋友。
LUKE|7|35|而智慧是由所有智慧的人来证实的。”
LUKE|7|36|有一个法利赛人请耶稣和他吃饭，耶稣就到那法利赛人家里去坐席。
LUKE|7|37|那城里有一个女人，是个罪人，知道耶稣在法利赛人家里坐席，就拿着盛满香膏的玉瓶，
LUKE|7|38|站在耶稣背后，挨着他的脚哭，眼泪滴湿了耶稣的脚，就用自己的头发擦干，又用嘴连连亲他的脚，把香膏抹上。
LUKE|7|39|请耶稣的法利赛人看见这事，心里说：“这人若是先知，一定知道摸他的是谁，是个怎样的女人；她是个罪人哪！”
LUKE|7|40|耶稣回应他说：“ 西门 ，我有话要对你说。” 西门 说：“老师，请说。”
LUKE|7|41|耶稣说：“有两个人欠了某一个债主的钱，一个欠五百个银币，一个欠五十个银币。
LUKE|7|42|因为他们无力偿还，债主就开恩赦免了他们两个人的债。那么，这两个人哪一个更爱他呢？”
LUKE|7|43|西门 回答：“我想是那多得赦免的人。”耶稣对他说：“你的判断不错。”
LUKE|7|44|于是他转过来向着那女人，对 西门 说：“你看见这女人吗？我进了你的家，你没有给我水洗脚，但这女人用眼泪滴湿了我的脚，又用头发擦干。
LUKE|7|45|你没有亲我，但这女人从我进来就不住地亲我的脚。
LUKE|7|46|你没有用油抹我的头，但这女人用香膏抹我的脚。
LUKE|7|47|所以我告诉你，她许多的罪都赦免了，因为她爱的多；而那少得赦免的，爱的就少。”
LUKE|7|48|于是耶稣对那女人说：“你的罪都赦免了。”
LUKE|7|49|同席的人心里说：“这是什么人，竟赦免人的罪呢？”
LUKE|7|50|耶稣对那女人说：“你的信救了你，平安地回去吧！”
LUKE|8|1|过了不久，耶稣周游各城各乡传道，宣讲上帝国的福音。和他同去的有十二个使徒，
LUKE|8|2|还有曾被邪灵所附，被疾病所缠，而已经治好的几个妇女，其中有称为 抹大拉 的 马利亚 ，曾有七个鬼从她身上赶出来，
LUKE|8|3|又有 希律 的管家 苦撒 的妻子 约亚拿 ，和 苏撒拿 以及好些别的妇女，她们都是用自己的财物供给耶稣和使徒。
LUKE|8|4|当一大群人聚集，又有人从各城里出来见耶稣的时候，耶稣用比喻说：
LUKE|8|5|“有一个撒种的出去撒种。他撒的时候，有的落在路旁，被人践踏，天上的飞鸟又来把它吃掉了。
LUKE|8|6|有的落在磐石上，一出来就枯干了，因为得不着滋润。
LUKE|8|7|有的落在荆棘里，荆棘跟它一同生长，把它挤住了。
LUKE|8|8|又有的落在好土里，生长起来，结实百倍。”耶稣说完这些话，大声说：“有耳可听的，就应当听！”
LUKE|8|9|门徒问耶稣这比喻是什么意思。
LUKE|8|10|他说：“上帝国的奥秘只让你们知道，至于别人，就用比喻，要 他们看也看不见， 听也不明白。”
LUKE|8|11|“这比喻是这样的：种子就是上帝的道。
LUKE|8|12|那些在路旁的，就是人听了道，随后魔鬼来，从他们心里把道夺去，以免他们信了得救。
LUKE|8|13|那些在磐石上的，就是人听道，欢喜领受，但没有根，不过暂时相信，等到碰上试炼就退后了。
LUKE|8|14|那落在荆棘里的，就是人听了道，走开以后，被今生的忧虑、钱财、宴乐挤住了，结不出成熟的子粒来。
LUKE|8|15|那落在好土里的，就是人听了道，并用纯真善良的心持守它，耐心等候结果实。”
LUKE|8|16|“没有人点灯用器皿盖上，或放在床底下，而是放在灯台上，让进来的人看见亮光。
LUKE|8|17|因为掩藏的事没有不显出来的，隐瞒的事也没有不露出来被人知道的。
LUKE|8|18|所以，你们应当小心怎样听。因为凡有的，还要给他；凡没有的，连他自以为有的也要夺去。”
LUKE|8|19|耶稣的母亲和他兄弟来看他，因为人多，不能到他跟前。
LUKE|8|20|有人告诉他说：“你母亲和你兄弟站在外边，要见你。”
LUKE|8|21|耶稣回答他们：“听了上帝的道而遵行的人，就是我的母亲，我的兄弟了。”
LUKE|8|22|有一天，耶稣和门徒上了船，他对门徒说：“我们渡到湖的对岸去吧。”他们就开了船。
LUKE|8|23|船行的时候，耶稣睡着了。湖上忽然起了狂风，船将灌满了水，很危险。
LUKE|8|24|门徒去叫醒他，说：“老师！老师！我们快没命啦！”耶稣醒了，斥责那狂风大浪，风浪就止住，平静了。
LUKE|8|25|耶稣对他们说：“你们的信心在哪里呢？”他们又惧怕又惊讶，彼此说：“这到底是谁？他吩咐风和水，连风和水都听从他。”
LUKE|8|26|他们到了 格拉森 人的地区，就在 加利利 的对面。
LUKE|8|27|耶稣上了岸，就有城里一个被鬼附的人迎着他走来。这个人好久不穿衣服，不住在屋子里，而住在坟墓里。
LUKE|8|28|他看见耶稣，就喊叫着俯伏在他面前，大声说：“至高上帝的儿子耶稣，你为什么干扰我？我求你，不要叫我受苦！”
LUKE|8|29|这是因耶稣曾吩咐污灵从这人身上出来。原来这污灵屡次抓住他；他常被人看守，又被铁链和脚镣捆锁，他竟把锁链挣断，被鬼赶到旷野去。
LUKE|8|30|耶稣问他：“你的名字叫什么？”他说：“ 群 ”；这是因为附着他的鬼多。
LUKE|8|31|鬼就央求耶稣不要命令他们到无底坑里去。
LUKE|8|32|那里有一大群猪正在山坡上吃食，鬼央求耶稣准他们进入猪里；耶稣准了他们。
LUKE|8|33|于是鬼从那人出来，进入猪里，那群猪就闯下山崖，投进湖里，淹死了。
LUKE|8|34|放猪的看见这事就逃跑了，去告诉城里和乡下的人。
LUKE|8|35|众人出来，要看发生了什么事；到了耶稣那里，发现那人坐在耶稣脚前，鬼已离开了他，穿着衣服，神智清醒，他们就害怕。
LUKE|8|36|看见这事的人把被鬼附的人怎么得医治的事告诉他们。
LUKE|8|37|格拉森 周围地区的人，因为害怕得很，都求耶稣离开他们；耶稣就上船回去了。
LUKE|8|38|鬼已从身上出去的那人恳求要和耶稣在一起，耶稣却打发他回去，说：
LUKE|8|39|“你回家去，传讲上帝为你做了多么大的事。”他就走遍全城，传扬耶稣为他做了多么大的事。
LUKE|8|40|耶稣回来的时候，众人迎接他，因为他们都等候着他。
LUKE|8|41|有一个会堂主管，名叫 叶鲁 ，来俯伏在耶稣脚前，求耶稣到他家里去，
LUKE|8|42|因为他有一个独生女，约十二岁，快要死了。 耶稣去的时候，众人簇拥着他。
LUKE|8|43|有一个女人，患了经血不止的病有十二年，在医生手里花尽了一生所有的 ，但没有人能治好她。
LUKE|8|44|她来到耶稣背后，摸他的衣裳繸子，经血立刻止住了。
LUKE|8|45|耶稣说：“摸我的是谁？”众人都不承认。 彼得 说：“老师，众人拥拥挤挤紧靠着你。”
LUKE|8|46|耶稣说：“有人摸了我，因为我觉得有能力从我身上出去。”
LUKE|8|47|那女人知道瞒不住了，就战战兢兢地俯伏在耶稣跟前，把摸他的缘故和怎样立刻痊愈的事，当着众人都说出来。
LUKE|8|48|耶稣对她说：“女儿，你的信救了你。平安地回去吧！”
LUKE|8|49|耶稣还在说话的时候，有人从会堂主管的家里来，说：“你的女儿死了，不要劳驾老师了。”
LUKE|8|50|耶稣听见就对他说：“不要怕，只要信！她必得痊愈。”
LUKE|8|51|耶稣到了他的家，除了 彼得 、 约翰 、 雅各 ，和女儿的父母，不许别人同他进去。
LUKE|8|52|众人都在为这女孩哀哭捶胸。耶稣说：“不要哭，她不是死了，是睡着了。”
LUKE|8|53|他们知道她已经死了，就嘲笑耶稣。
LUKE|8|54|耶稣拉着她的手，呼叫着：“孩子，起来吧！”
LUKE|8|55|她的灵魂就回来了，她立刻起来。耶稣吩咐给她东西吃。
LUKE|8|56|她的父母非常惊奇；耶稣吩咐他们不要把所发生的事告诉任何人。
LUKE|9|1|耶稣叫齐了十二使徒，给他们能力和权柄制伏一切的鬼，医治疾病，
LUKE|9|2|又差遣他们宣讲上帝的国，医治病人，
LUKE|9|3|对他们说：“途中什么都不要带；不要带手杖和行囊，不要带食物和银钱，也不要带两件内衣 。
LUKE|9|4|你们无论进哪一家，就住在哪里，也从那里离开。
LUKE|9|5|凡不接待你们的，你们离开那城的时候，要跺掉你们脚上的尘土，证明他们的不是。”
LUKE|9|6|于是使徒出去，走遍各乡传福音，到处治病。
LUKE|9|7|希律 分封王听见耶稣所做的一切事，就困惑起来，因为有人说：“ 约翰 从死人中复活了。”
LUKE|9|8|又有人说：“ 以利亚 显现了。”还有人说：“古时的一个先知又活了。”
LUKE|9|9|希律 说：“ 约翰 我已经斩了，但这是什么人？关于他，我竟听到这样的事！”于是 希律 想要见他。
LUKE|9|10|使徒们回来，把所做的事告诉耶稣，耶稣就私下带他们离开那里，往一座叫 伯赛大 的城去。
LUKE|9|11|众人知道了，就跟着他去；耶稣接待他们，对他们讲论上帝国的事，治好那些需要医治的人。
LUKE|9|12|太阳快要下山，十二使徒进前来对他说：“请叫众人散去，他们好往四面村庄乡镇里去借宿和找吃的，因为我们这里地方偏僻。”
LUKE|9|13|耶稣对他们说：“你们给他们吃吧！”他们说：“我们不过有五个饼、两条鱼，若不去为这许多人买食物就不够。”
LUKE|9|14|那时，男人约有五千。耶稣对门徒说：“叫他们分组坐下，每组大约五十个人。”
LUKE|9|15|门徒就这样做了，叫众人都坐下。
LUKE|9|16|耶稣拿着这五个饼和两条鱼，望着天祝福，擘开，递给门徒，摆在众人面前。
LUKE|9|17|所有的人都吃，并且吃饱了。他们把剩下的碎屑收拾起来，装满了十二个篮子。
LUKE|9|18|耶稣独自祷告的时候，门徒也同他在那里。耶稣问他们：“众人说我是谁？”
LUKE|9|19|他们回答：“是施洗的 约翰 ；有人说是 以利亚 ；还有人说是古时的一个先知又活了。”
LUKE|9|20|耶稣问他们：“你们说我是谁？” 彼得 回答：“是上帝所立的基督。”
LUKE|9|21|耶稣切切吩咐他们，命令他们不可把这事告诉任何人；
LUKE|9|22|又说：“人子必须受许多的苦，被长老、祭司长和文士弃绝，并且被杀，第三天复活。”
LUKE|9|23|耶稣又对众人说：“若有人要跟从我，就当舍己，天天背起自己的十字架来跟从我。
LUKE|9|24|因为凡要救自己生命的，必丧失生命；凡为我丧失生命的，他必救自己的生命。
LUKE|9|25|人就是赚得全世界，却丧失了自己，或赔上自己，有什么益处呢？
LUKE|9|26|凡把我和我的道当作可耻的，人子在自己的荣耀里，和天父与圣天使的荣耀里来临的时候，也要把那人当作可耻的。
LUKE|9|27|我实在告诉你们，站在这里的，有人在没经历死亡以前，必定看见上帝的国。”
LUKE|9|28|说了这些话以后约有八天，耶稣带着 彼得 、 约翰 、 雅各 上山去祷告。
LUKE|9|29|正祷告的时候，他的面貌改变了，衣服洁白放光。
LUKE|9|30|忽然有 摩西 和 以利亚 两个人同耶稣说话；
LUKE|9|31|他们在荣光里显现，谈论耶稣去世的事，就是他在 耶路撒冷 将要完成的事。
LUKE|9|32|彼得 和他的同伴都打盹，但一清醒，就看见耶稣的荣光和与他一起站着的那两个人。
LUKE|9|33|二人正要和耶稣分离的时候， 彼得 对耶稣说：“老师，我们在这里真好！我们来搭三座棚，一座为你，一座为 摩西 ，一座为 以利亚 。”他却不知道自己在说些什么。
LUKE|9|34|说这些话的时候，有一朵云彩来遮盖他们；他们一进入云彩就很惧怕。
LUKE|9|35|有声音从云彩里出来，说：“这是我的儿子，我所拣选的 。你们要听从他！”
LUKE|9|36|声音停止后，只见耶稣独自一人。当那些日子，门徒保持沉默，不把所看见的事告诉任何人。
LUKE|9|37|第二天，他们下了山，有一大群人来迎见耶稣。
LUKE|9|38|其中有一人喊着说：“老师！求你看看我的儿子，因为他是我的独子。
LUKE|9|39|他被灵拿住就突然喊叫，那灵又使他抽风，口吐白沫，并且重重地伤害他，不轻易放过他。
LUKE|9|40|我求过你的门徒把那灵赶出去，他们却不能。”
LUKE|9|41|耶稣回答：“唉！这又不信又悖谬的世代啊，我和你们在一起，忍耐你们，要到几时呢？把你的儿子带到这里来！”
LUKE|9|42|他正来的时候，那鬼把他摔倒，使他重重地抽风。耶稣斥责那污灵，把孩子治好了，交给他父亲。
LUKE|9|43|众人都诧异上帝的大能 。 众人正惊讶于耶稣所做的一切事的时候，耶稣对门徒说：
LUKE|9|44|“你们要把这些话听进去，因为人子将要被交在人手里。”
LUKE|9|45|门徒却不明白这话，其中的意思对他们隐藏着，使他们不能明白，他们也不敢问这话的意思。
LUKE|9|46|门徒互相议论，他们中间谁最大。
LUKE|9|47|耶稣看出他们心中的议论，就领一个小孩子来，叫他站在自己旁边，
LUKE|9|48|对他们说：“凡为我的名接纳这小孩子的，就是接纳我；凡接纳我的，就是接纳那差我来的。你们中间最小的，他就是最大的。”
LUKE|9|49|约翰 回应说：“老师，我们看见一个人奉你的名赶鬼，我们就阻止他，因为他不与我们一同跟从你。”
LUKE|9|50|耶稣对他说：“不要阻止他，因为不抵挡你们的，就是帮助你们的。”
LUKE|9|51|耶稣被接上升的日子将到，他决定面向 耶路撒冷 走去。
LUKE|9|52|他打发使者在他前头走；他们进了 撒玛利亚 的一个村庄，要为他作准备。
LUKE|9|53|那里的人不接待他，因为他面向着 耶路撒冷 去。
LUKE|9|54|他的门徒 雅各 和 约翰 看见了，就说：“主啊！你要我们吩咐火从天上降下来，烧灭他们 吗？”
LUKE|9|55|耶稣转身责备两个门徒。
LUKE|9|56|于是他们就往别的村庄去了。
LUKE|9|57|他们在路上走的时候，有一个人对耶稣说：“你无论往哪里去，我都要跟从你。”
LUKE|9|58|耶稣对他说：“狐狸有洞，天空的飞鸟有窝，人子却没有枕头的地方。”
LUKE|9|59|他又对另一个人说：“来跟从我！”那人说：“主啊 ，容许我先回去埋葬我的父亲。”
LUKE|9|60|耶稣对他说：“让死人埋葬他们的死人，你只管去传讲上帝的国。”
LUKE|9|61|又有一人说：“主啊，我要跟从你，但容许我先去辞别我家里的人。”
LUKE|9|62|耶稣对他说：“手扶着犁向后看的人，不配进上帝的国。”
LUKE|10|1|这些事以后，主另外指定七十二个人 ，差遣他们两个两个地在他前面，往自己所要到的各城各地去。
LUKE|10|2|他对他们说：“要收的庄稼多，做工的人少。所以，你们要求庄稼的主差遣做工的人出去收他的庄稼。
LUKE|10|3|你们去吧！看！我差你们出去，如同羔羊进入狼群。
LUKE|10|4|不要带钱囊，不要带行囊，不要带鞋子；在路上也不要向人问安。
LUKE|10|5|无论进哪一家，先要说：‘愿这一家平安。’
LUKE|10|6|那里若有当得平安的人，你们所求的平安就必临到那家，不然，将归还你们。
LUKE|10|7|你们要住在那家，吃喝他们所供给的，因为工人得工钱是应当的；不要从这家搬到那家。
LUKE|10|8|无论进哪一城，人若接待你们，给你们摆上什么食物，你们就吃什么。
LUKE|10|9|要医治那城里的病人，对他们说：‘上帝的国临近你们了。’
LUKE|10|10|无论进哪一城，人若不接待你们，你们就到大街上去，说：
LUKE|10|11|‘就是你们城里的尘土粘在我们的脚上，我们也当着你们擦去。但是，你们该知道上帝的国临近了。’
LUKE|10|12|我告诉你们，在那日子， 所多玛 所受的，比那城还容易受呢！”
LUKE|10|13|“ 哥拉汛 哪，你有祸了！ 伯赛大 啊，你有祸了！因为在你们中间所行的异能，若行在 推罗 、 西顿 ，他们早已披麻蒙灰，坐在地上悔改了。
LUKE|10|14|在审判的时候， 推罗 和 西顿 所受的，比你们还容易受呢！
LUKE|10|15|迦百农 啊， 你以为要被举到天上吗？ 你要被推下阴间！”
LUKE|10|16|耶稣又对门徒说：“听从你们的就是听从我；弃绝你们的就是弃绝我；弃绝我的就是弃绝差遣我来的那位。”
LUKE|10|17|那七十二个人欢欢喜喜地回来，说：“主啊，因你的名，就是鬼也服了我们。”
LUKE|10|18|耶稣对他们说：“我看见撒但从天上坠落，像闪电一样。
LUKE|10|19|我已经给你们权柄可以践踏蛇和蝎子，又胜过仇敌一切的能力，绝没有什么能害你们。
LUKE|10|20|然而，不要因灵服了你们就欢喜，而要因你们的名记录在天上欢喜。”
LUKE|10|21|正当那时，耶稣被圣灵感动而欢喜快乐，说：“父啊，天地的主，我感谢你！因为你把这些事向聪明智慧的人隐藏起来，而向婴孩启示出来。父啊，是的，因为你的美意本是如此。
LUKE|10|22|一切都是我父交给我的。除了父，没有人知道子是谁；除了子和子所愿意启示的人，没有人知道父是谁。”
LUKE|10|23|耶稣转身私下对门徒说：“看见你们所看见的，那眼睛有福了。
LUKE|10|24|我告诉你们，从前有许多先知和君王要看你们所看的，却没有看见，要听你们所听的，却没有听见。”
LUKE|10|25|有一个律法师起来试探耶稣，说：“老师！我该做什么才可以承受永生？”
LUKE|10|26|耶稣对他说：“律法上写的是什么？你是怎样念的呢？”
LUKE|10|27|他回答说：“你要尽心、尽性、尽力、尽意爱主—你的上帝，又要爱邻 如己。”
LUKE|10|28|耶稣对他说：“你回答得正确，你这样做就会得永生。”
LUKE|10|29|那人要证明自己有理，就对耶稣说：“谁是我的邻舍呢？”
LUKE|10|30|耶稣回答：“有一个人从 耶路撒冷 下 耶利哥 去，落在强盗手中。他们剥去他的衣裳，把他打个半死，丢下他走了。
LUKE|10|31|偶然有一个祭司从那条路下来，看见他就从另一边过去了。
LUKE|10|32|又有一个 利未 人来到那里，看见他，也照样从另一边过去了。
LUKE|10|33|可是，有一个 撒玛利亚 人路过那里，看见他就动了慈心，
LUKE|10|34|上前用油和酒倒在他的伤处，包裹好了，扶他骑上自己的牲口，带他到旅店里去，照应他。
LUKE|10|35|第二天，他拿出两个银币来，交给店主，说：‘请你照应他，额外的费用，我回来时会还你。’
LUKE|10|36|你想，这三个人哪一个是落在强盗手中那人的邻舍呢？”
LUKE|10|37|他说：“是怜悯他的。”耶稣对他说：“你去，照样做吧！”
LUKE|10|38|他们继续前行，耶稣进了一个村庄。有一个女人，名叫 马大 ，接他到自己家里。
LUKE|10|39|她有一个妹妹，名叫 马利亚 ，在主的脚前坐着听他的道。
LUKE|10|40|马大 伺候的事多，心里忙乱，进前来，说：“主啊，我的妹妹留下我一个人伺候，你不在意吗？请吩咐她来帮助我。”
LUKE|10|41|主回答说：“ 马大 ， 马大 ，你为许多的事操心烦恼，
LUKE|10|42|但是不可少的只有一件 。 马利亚 已经选择了那上好的福分，是没有人能从她夺去的。”
LUKE|11|1|耶稣在一个地方祷告。祷告完了，有个门徒对他说：“主啊，求你教导我们祷告，像 约翰 教导他的门徒一样。”
LUKE|11|2|耶稣对他们说：“你们祷告的时候，要说： ‘父啊， 愿人都尊你的名为圣； 愿你的国降临；
LUKE|11|3|我们日用的饮食，天天赐给我们。
LUKE|11|4|赦免我们的罪， 因为我们也赦免凡亏欠我们的人。 不叫我们陷入试探。 ’”
LUKE|11|5|耶稣又对他们说：“你们中间谁有一个朋友半夜到他那里去，对他说：‘朋友！请借给我三个饼；
LUKE|11|6|因为我有一个朋友旅途中来到我这里，我没有东西招待他。’
LUKE|11|7|那人在里面回答：‘不要打扰我，门已经关了，孩子们也同我在床上了，我不能起来给你。’
LUKE|11|8|我告诉你们，虽不因他是朋友起来给他，也会因他不顾面子地直求，起来照他所需要的给他。
LUKE|11|9|我又告诉你们，祈求，就给你们；寻找，就找到；叩门，就给你们开门。
LUKE|11|10|因为凡祈求的，就得着；寻找的，就找到；叩门的，就给他开门。
LUKE|11|11|你们中间作父亲的，谁有儿子 求鱼，反拿蛇当鱼给他呢？
LUKE|11|12|求鸡蛋，反给他蝎子呢？
LUKE|11|13|你们虽然不好，尚且知道拿好东西给儿女，何况 天父，他岂不更要把圣灵赐给求他的人吗？”
LUKE|11|14|耶稣赶出一个使人成为哑巴的鬼 ，鬼出去了，哑巴就说出话来；众人都很惊讶。
LUKE|11|15|其中却有人说：“他是靠着鬼王 别西卜 赶鬼。”
LUKE|11|16|又有人试探耶稣，要他显个来自天上的神迹。
LUKE|11|17|他知道他们的意念，就对他们说：“一国自相纷争，必定荒芜；一家自相纷争，就必败落。
LUKE|11|18|撒但若自相纷争，他的国怎能立得住呢？因为你们说我是靠着 别西卜 赶鬼。
LUKE|11|19|我若靠着 别西卜 赶鬼，你们的子弟赶鬼又靠着谁呢？这样，他们要作你们的判官。
LUKE|11|20|我若靠着上帝的能力赶鬼，那么，上帝的国就已临到你们了。
LUKE|11|21|壮士全副武装，看守自己的住宅，他所有的都很安全；
LUKE|11|22|但有一个比他更强的来攻击他，并且战胜了他，就夺去他所倚靠的盔甲兵器，又分了他的掠物。
LUKE|11|23|不跟我一起的，就是反对我；不与我一起收聚的，就是在拆散。”
LUKE|11|24|“污灵离了人身，走遍无水之地寻找安歇之处，却找不到。就说：‘我要回到我原来的屋里去。’
LUKE|11|25|他到了，看见里面打扫干净，修饰好了，
LUKE|11|26|就去另带了七个比自己更恶的灵来，都进去住在那里。那人后来的景况比先前更坏了。”
LUKE|11|27|耶稣正说这些话的时候，众人中间有一个女人高声对他说：“怀你胎乳养你的有福了！”
LUKE|11|28|耶稣却说：“更有福的是听上帝的道而遵守的人！”
LUKE|11|29|当众人越来越拥挤的时候，耶稣说：“这世代是一个邪恶的世代。他们求看神迹，除了 约拿 的神迹以外，再没有神迹给他们看了。
LUKE|11|30|约拿 怎样为 尼尼微 人成了神迹，人子也要照样为这世代的人成为神迹。
LUKE|11|31|在审判的时候，南方的女王要起来定这世代的人的罪，因为她从地极而来，要听 所罗门 智慧的话。看哪，比 所罗门 更大的在这里！
LUKE|11|32|在审判的时候， 尼尼微 人要起来定这世代的罪，因为 尼尼微 人听了 约拿 所传的就悔改了。看哪，比 约拿 更大的在这里！”
LUKE|11|33|“没有人点灯放在地窖里，或是斗底下 ，总是放在灯台上，让进来的人看见亮光。
LUKE|11|34|你的眼睛就是身体的灯。当你的眼睛明亮，全身就光明，当眼睛昏花，全身就黑暗。
LUKE|11|35|所以，你要注意，免得你里面的光暗了。
LUKE|11|36|若是你全身光明，毫无黑暗，就必全然光明，如同灯的明光照亮你。”
LUKE|11|37|耶稣正说话的时候，有一个法利赛人请他吃饭，耶稣就进去坐席。
LUKE|11|38|这法利赛人看见耶稣饭前不先洗手就很诧异。
LUKE|11|39|主对他说：“如今你们法利赛人洗净杯盘的外面，你们里面却满了贪婪和邪恶。
LUKE|11|40|无知的人哪！造外面的，不也造了里面吗？
LUKE|11|41|只要把杯盘里面的施舍给人，对你们来说一切就都洁净了。
LUKE|11|42|“但是你们法利赛人有祸了！因为你们将薄荷、芸香，和各样蔬菜献上十分之一，疏忽了公义和爱上帝的事；这原是你们该做的—至于其他也不可忽略。
LUKE|11|43|你们法利赛人有祸了！因为你们喜爱会堂里的高位，又喜欢人们在街市上向你们问安。
LUKE|11|44|你们有祸了！因为你们如同不显露的坟墓，走在上面的人并不知道。”
LUKE|11|45|律法师中有一个回答耶稣，说：“老师，你这样说也把我们侮辱了。”
LUKE|11|46|耶稣说：“你们律法师也有祸了！因为你们把难挑的担子放在别人身上，自己却不肯动一个指头去减轻这些担子。
LUKE|11|47|你们有祸了！因为你们建造先知的坟墓，那些先知正是你们的祖宗所杀的。
LUKE|11|48|可见你们祖宗所做的事，你们是证人，你们也赞同，因为他们杀了先知，你们建造先知的坟墓。
LUKE|11|49|所以，上帝的智慧也曾说：‘我要差遣先知和使徒到他们那里去，有的他们要残杀，有的他们要迫害’，
LUKE|11|50|为使创世以来所流众先知的血的罪都归在这世代的人身上，
LUKE|11|51|就是从 亚伯 的血起，直到被杀在祭坛和圣所中间的 撒迦利亚 的血为止。是的，我告诉你们，这都要向这世代的人追讨。
LUKE|11|52|你们律法师有祸了！因为你们把知识的钥匙夺了去，自己不进去，要进去的人，你们也阻挡他们。”
LUKE|11|53|耶稣从那里出来，文士和法利赛人就开始极力地催逼他，盘问他许多事，
LUKE|11|54|伺机要抓他的话柄。
LUKE|12|1|这时，有几万人聚集，甚至彼此践踏。耶稣就先对门徒说：“你们要防备法利赛人的酵，就是假冒为善。
LUKE|12|2|掩盖的事没有不显露出来的，隐藏的事也没有不被人知道的。
LUKE|12|3|因此，你们在暗中所说的，将要在明处被人听见；在密室附耳所说的，将要在屋顶上被人宣扬。”
LUKE|12|4|“我的朋友，我对你们说，那最多只能杀人身体而不能再做什么的，不要怕他们。
LUKE|12|5|我提醒你们该怕的是谁：该怕那杀了以后又有权柄把人扔在地狱里的。是的，我告诉你们，正要怕他。
LUKE|12|6|五只麻雀不是卖二铜钱 吗？但在上帝面前，一只也不被忘记；
LUKE|12|7|就是你们的头发也都数过了。不要惧怕，你们比许多的麻雀还贵重！”
LUKE|12|8|“我又告诉你们，凡在人面前认我的，人子在上帝的使者面前也必认他；
LUKE|12|9|在人面前不认我的，人子在上帝的使者面前也必不认他。
LUKE|12|10|凡说话干犯人子的，还可得赦免；但是亵渎圣灵的，总不得赦免。
LUKE|12|11|有人带你们到会堂、官长和掌权的人面前，不要担心怎么答辩，说什么话；
LUKE|12|12|因为就在那时候，圣灵要指教你们该说的话。”
LUKE|12|13|人群中有一个人对耶稣说：“老师！请你吩咐我的兄弟和我分家产。”
LUKE|12|14|耶稣对他说：“你这个人！谁立我作你们的判官，或给你们分家产的呢？”
LUKE|12|15|于是他对他们说：“你们要谨慎自守，躲避一切的贪心，因为人的生命不在于家道丰富。”
LUKE|12|16|然后他用比喻对他们说：“有一个财主，田地出产丰富。
LUKE|12|17|他自己心里想：‘我的出产没有地方储藏，怎么办呢？’
LUKE|12|18|就说：‘我要这么办：要把我的仓库拆了，另盖更大的，在那里好储藏我一切的粮食和财物，
LUKE|12|19|然后要对我自己说：你这个人哪，你有许多财物积存，可供多年享用，只管安安逸逸吃喝快乐吧！’
LUKE|12|20|上帝却对他说：‘无知的人哪！今夜就要你的性命，你所预备的要归谁呢？’
LUKE|12|21|凡为自己积财，在上帝面前却不富足的，也是这样。”
LUKE|12|22|耶稣又对门徒说：“所以，我告诉你们，不要为生命忧虑吃什么，为身体忧虑穿什么。
LUKE|12|23|因为生命胜于饮食，身体胜于衣裳。
LUKE|12|24|你们想一想乌鸦：它们既不种也不收，既没有仓又没有库，上帝尚且养活它们。你们比飞鸟要贵重得多呢！
LUKE|12|25|你们哪一个能藉着忧虑使寿数多加一刻呢 ？
LUKE|12|26|这最小的事你们尚且不能做，何必忧虑其余的事呢？
LUKE|12|27|你们想一想百合花是怎么长起来的：它也不劳动，也不纺线。然而我告诉你们，就是 所罗门 极荣华的时候，他所穿戴的还不如这些花的一朵呢！
LUKE|12|28|你们这小信的人哪！野地里的草今天还在，明天就丢在炉里，上帝还给它这样的妆饰，何况你们呢？
LUKE|12|29|你们不要求吃什么，喝什么，也不要挂虑。
LUKE|12|30|这都是世上的外邦人所求的；你们需要这些东西，你们的父都知道。
LUKE|12|31|你们只要求他的国，这些东西就必加给你们了。
LUKE|12|32|你们这小群，不要惧怕，因为你们的父乐意把国赐给你们。
LUKE|12|33|你们要变卖财产周济人，为自己预备永不坏的钱囊和用不尽的财宝在天上，就是贼不能近，虫不能蛀的地方。
LUKE|12|34|因为你们的财宝在哪里，你们的心也在哪里。”
LUKE|12|35|“你们要束紧腰带，灯也要点着，
LUKE|12|36|好像仆人等候自己的主人从婚宴上回来。他来叩门，就立刻给他开门。
LUKE|12|37|主人来了，看见仆人警醒，那些仆人就有福了。我实在告诉你们，主人会叫他们坐席，自己束上腰带，前来伺候他们。
LUKE|12|38|他或是半夜来，或是天亮之前来，看见仆人这样，那些仆人就有福了。
LUKE|12|39|你们要知道，一家的主人若知道贼什么时候来，就 不容贼挖穿房屋。
LUKE|12|40|你们也要预备，因为在你们想不到的时候，人子就来了。”
LUKE|12|41|彼得 说：“主啊，这比喻是对我们说的呢？还是也对众人呢？”
LUKE|12|42|主说：“那么，谁是那忠心又精明的管家，主人要派他管理自己的家仆，按时定量分粮给他们的呢？
LUKE|12|43|主人来到，看见仆人这样做，那仆人就有福了。
LUKE|12|44|我实在告诉你们，主人要派他管理所有的财产。
LUKE|12|45|如果那仆人心里说‘我的主人会来得迟’，就动手打僮仆和使女，并且吃喝醉酒，
LUKE|12|46|在想不到的日子，不知道的时候，那仆人的主人要来，重重地惩罚他 ，定他和不忠心的人同罪。
LUKE|12|47|仆人知道主人的意思，却没预备，又未顺他的意思做，那仆人要多受责打；
LUKE|12|48|至于那不知道而做了当受责打的事的，要少受责打。多给谁，就向谁多取；多托谁，就向谁多要。”
LUKE|12|49|“我来是要把火丢在地上，假如已经烧起来，不也是我所希望的吗？
LUKE|12|50|我有当受的洗还没有受，在这事完成之前，我是多么地焦急！
LUKE|12|51|你们以为我来是要使地上太平吗？不！我告诉你们，是使人纷争。
LUKE|12|52|从今以后，一家五个人将要纷争，三个和两个相争，两个和三个相争：
LUKE|12|53|父亲和儿子相争， 儿子和父亲相争； 母亲和女儿相争， 女儿和母亲相争； 婆婆和媳妇相争， 媳妇和婆婆相争。”
LUKE|12|54|耶稣又对众人说：“你们看见西边起了云彩，就说：‘要下大雨了’，果然就有；
LUKE|12|55|起了南风，你们就说：‘要燥热了’，也就有了。
LUKE|12|56|假冒为善的人哪，你们知道分辨天地的气象，怎么不知道分辨这是什么时代呢？”
LUKE|12|57|“你们又为何不自己判断什么是合理的呢？
LUKE|12|58|你同告你的冤家去见官，还在路上，要尽力跟他和解，免得他拉你到法官面前，法官把你交给法警，法警把你下在监里。
LUKE|12|59|我告诉你，就是最后一小文钱 还没有还清，你也绝不能从那里出来。”
LUKE|13|1|正当那时，有些在场的人把 彼拉多 使 加利利 人的血搀杂在他们祭物中的事，告诉耶稣。
LUKE|13|2|耶稣对他们说：“你们以为这些 加利利 人比其他的 加利利 人更有罪，所以受这害吗？
LUKE|13|3|我告诉你们，不是的！你们若不悔改，都同样要灭亡！
LUKE|13|4|从前 西罗亚 楼倒塌，压死了十八个人，你们以为那些人比一切住在 耶路撒冷 的人更有罪吗？
LUKE|13|5|我告诉你们，不是的！你们若不悔改，都照样要灭亡！”
LUKE|13|6|于是，耶稣用比喻说：“有一个人在葡萄园里栽了一棵无花果树。他前来在树上找果子，却找不到，
LUKE|13|7|就对园丁说：‘看哪，我这三年来到这棵无花果树前找果子，竟找不到。把它砍了吧，何必白占土地呢？’
LUKE|13|8|园丁回答：‘主啊，今年且留着，等我在树周围掘开土，加上肥料，
LUKE|13|9|以后若结果子便罢，不然再把它砍了。’”
LUKE|13|10|安息日，耶稣在一个会堂里教导人。
LUKE|13|11|有一个女人被灵附身，病了十八年，腰弯得一点都直不起来。
LUKE|13|12|耶稣看见，就叫她过来，对她说：“妇人，你的病好了！”
LUKE|13|13|于是用双手按着她，她立刻直起腰来，就归荣耀给上帝。
LUKE|13|14|会堂的主管因为耶稣在安息日治病，就很生气，对众人说：“有六天应当做工，那六天之内可以来求医，在安息日却不可。”
LUKE|13|15|主回答他：“假冒为善的人哪，难道你们各人在安息日不解开槽上的牛和驴，牵去喝水吗？
LUKE|13|16|何况她本是 亚伯拉罕 的后裔，被撒但捆绑了十八年，不该在安息日这天解开她的绑吗？”
LUKE|13|17|耶稣说这些话，他的敌人都惭愧了；所有的人因他所做一切荣耀的事都很欢喜。
LUKE|13|18|耶稣说：“上帝的国像什么？我拿什么来比拟呢？
LUKE|13|19|它好比一粒芥菜种，有人拿去种在园子里，长大成树，天上的飞鸟在它的枝上筑巢。”
LUKE|13|20|他又说：“我拿什么来比拟上帝的国呢？
LUKE|13|21|它好比面酵，有妇人拿来放进三斗面里，直到全团都发起来。”
LUKE|13|22|耶稣往 耶路撒冷 去，在所经过的各城各乡教导人。
LUKE|13|23|有一个人问他：“主啊，得救的人很少吧？” 耶稣对众人说：
LUKE|13|24|“你们要努力进窄门。我告诉你们，将来有许多人想要进去，却不能。
LUKE|13|25|等到一家之主起来关了门，你们才站在外面敲门，说：‘主啊，给我们开门！’他要回答你们说：‘我不认识你们，不知道你们是哪里来的。’
LUKE|13|26|那时，你们要说：‘我们在你面前吃过喝过，你也在我们的街上教导过人。’
LUKE|13|27|他要对你们说：‘我 告诉你们，我不知道你们是哪里来的。你们这一切不义的人，给我走开！’
LUKE|13|28|你们要看见 亚伯拉罕 、 以撒 、 雅各 和众先知都在上帝的国里，你们却被赶到外面，在那里要哀哭切齿了。
LUKE|13|29|从东从西，从南从北，将有人来，在上帝的国里坐席。
LUKE|13|30|看吧，在后的，将要在前；在前的，将要在后。”
LUKE|13|31|就在那时，有几个法利赛人来对耶稣说：“离开这里到别处去吧，因为 希律 想要杀你。”
LUKE|13|32|耶稣对他们说：“你们去告诉那个狐狸：‘你看吧，今天明天我赶鬼治病，第三天我的事就成了。’
LUKE|13|33|虽然这样，今天明天后天我必须向前走，因为先知是不可能在 耶路撒冷 之外被害的。
LUKE|13|34|耶路撒冷 啊， 耶路撒冷 啊，你常杀害先知，又用石头打死那奉差遣到你这里来的人。我多少次想聚集你的儿女，好像母鸡把小鸡聚集在翅膀底下，可是你们不愿意。
LUKE|13|35|看吧，你们的家要被废弃。我告诉你们，你们绝不会再见到我，直到你们说：‘奉主名来的是应当称颂的！’”
LUKE|14|1|安息日，耶稣到一个法利赛人的领袖家里去吃饭，他们就窥探他。
LUKE|14|2|这时在他面前有一个患水肿病的人。
LUKE|14|3|耶稣回答律法师和法利赛人，说：“安息日治病合不合法？”
LUKE|14|4|他们却不说话。耶稣扶着那人，治好了他，叫他走了。
LUKE|14|5|耶稣对他们说：“你们中间谁有儿子 或有牛在安息日掉在井里，不立刻拉他上来呢？”
LUKE|14|6|他们对这些事不能反驳。
LUKE|14|7|耶稣见所请的客人选择首位，就用比喻对他们说：
LUKE|14|8|“你被人请去赴婚宴，不要坐在首位上，恐怕主人请了比你尊贵的客人，
LUKE|14|9|请了你和他的那人前来，对你说：‘请让座给这一位吧。’你就羞羞惭惭地退到末位去了。
LUKE|14|10|你被请的时候，去坐在末位上，好让主人来对你说：‘朋友，请上座。’那时，你在同席的人面前就有光彩了。
LUKE|14|11|因为凡自高的，必降为卑；自甘卑微的，必升为高。”
LUKE|14|12|耶稣又对请他的人说：“你准备午饭或晚餐，不要请你的朋友、弟兄、亲属和富足的邻舍，免得他们回请你，你就得了报答。
LUKE|14|13|你摆设宴席，倒要请那贫穷的、残疾的、瘸腿的、失明的，
LUKE|14|14|你就有福了！因为他们没有什么可报答你。到义人复活的时候，你要得到报答。”
LUKE|14|15|同席的有一人听见这些话，就对耶稣说：“在上帝国里吃饭的有福了！”
LUKE|14|16|耶稣对他说：“有人摆设大宴席，请了许多客人。
LUKE|14|17|到了坐席的时候，他打发仆人去对所请的人说：‘请来吧！样样都已齐备了。’
LUKE|14|18|众人异口同声地推辞。头一个对他说：‘我买了一块地，必须去看看。请你准我辞了。’
LUKE|14|19|另一个说：‘我买了五对牛，要去试一试。请你准我辞了。’
LUKE|14|20|又有一个说：‘我才娶了妻子，所以不能去。’
LUKE|14|21|那仆人回来，把这些事都告诉了主人。这家的主人就发怒，对仆人说：‘快出去，到城里大街小巷，领那贫穷的、残疾的、失明的、瘸腿的来。’
LUKE|14|22|仆人说：‘主啊，你所吩咐的已经办了，还有空位。’
LUKE|14|23|主人对仆人说：‘你出去，到大街小巷强拉人进来，坐满我的屋子。
LUKE|14|24|我告诉你们，先前所请的人没有一个可以尝到我的宴席。’”
LUKE|14|25|有一大群人和耶稣同行。他转过来对他们说：
LUKE|14|26|“无论什么人到我这里来，若不爱我胜过爱 自己的父母、妻子、儿女、兄弟、姊妹，甚至自己的性命，就不能作我的门徒。
LUKE|14|27|凡不背着自己的十字架来跟从我的，也不能作我的门徒。
LUKE|14|28|你们哪一个要盖一座楼，不先坐下来计算费用，看能不能盖成？
LUKE|14|29|免得安了地基，不能盖成，看见的人都笑话他，说：
LUKE|14|30|‘这个人开了工，却不能完工。’
LUKE|14|31|或是一个王出去和别的王打仗，岂不先坐下来酌量，他能不能用一万兵去抵抗那领二万兵来攻打他的吗？
LUKE|14|32|若是不能，他就趁敌人还远的时候，派使者去谈和平的条件。
LUKE|14|33|这样，你们无论什么人，若不撇下一切所有的，就不能作我的门徒。”
LUKE|14|34|“盐本是好的；盐若失了味，怎能叫它再咸呢？
LUKE|14|35|或用在田里，或堆在粪里，都不合适，只好丢在外面。有耳可听的，就应当听！”
LUKE|15|1|许多税吏和罪人都挨近耶稣，要听他讲道。
LUKE|15|2|法利赛人和文士私下议论说：“这个人接纳罪人，又同他们吃饭。”
LUKE|15|3|耶稣就用比喻对他们说：
LUKE|15|4|“你们中间谁有一百只羊，失去其中的一只，不把这九十九只留在旷野，去找那失去的羊，直到找着呢？
LUKE|15|5|找到了，他就欢欢喜喜地把羊扛在肩上。
LUKE|15|6|他回到家里，请朋友和邻舍来，对他们说：‘你们和我一同欢喜吧，我失去的羊已经找到了！’
LUKE|15|7|我告诉你们，一个罪人悔改，在天上也要这样为他欢喜，比为九十九个不用悔改的义人欢喜还大呢！”
LUKE|15|8|“同样，哪一个妇人有十块钱 ，若失落一块，不点上灯，打扫屋子，细细地找，直到找着呢？
LUKE|15|9|找到了，她就请朋友和邻舍来，对她们说：‘你们和我一同欢喜吧，我失落的那块钱已经找到了！’
LUKE|15|10|我告诉你们，一个罪人悔改，上帝的使者也是这样为他欢喜。”
LUKE|15|11|耶稣又说：“一个人有两个儿子。
LUKE|15|12|小儿子对父亲说：‘父亲，请你把我应得的家业分给我。’他父亲就把财产分给他们。
LUKE|15|13|过了不多几天，小儿子把他一切所有的都收拾起来，往远方去了。在那里，他任意放荡，浪费钱财。
LUKE|15|14|他耗尽了一切所有的，又恰逢那地方有大饥荒，就穷困起来。
LUKE|15|15|于是他去投靠当地的一个居民，那人打发他到田里去放猪。
LUKE|15|16|他恨不得拿猪所吃的豆荚充饥，也没有人给他什么吃的。
LUKE|15|17|他醒悟过来，就说：‘我父亲有多少雇工，粮食有余，我倒在这里饿死吗？
LUKE|15|18|我要起来，到我父亲那里去，对他说：父亲！我得罪了天，又得罪了你，
LUKE|15|19|从今以后，我不配称为你的儿子，把我当作一个雇工吧。’
LUKE|15|20|于是他起来，往他父亲那里去。相离还远，他父亲看见，就动了慈心，跑去拥抱着他，连连亲他。
LUKE|15|21|儿子对他说：‘父亲！我得罪了天，又得罪了你，从今以后，我不配称为你的儿子。’
LUKE|15|22|父亲却吩咐仆人：‘快把那上好的袍子拿出来给他穿，把戒指戴在他指头上，把鞋穿在他脚上，
LUKE|15|23|把那肥牛犊牵来宰了，我们来吃喝庆祝；
LUKE|15|24|因为我这个儿子是死而复活，失而复得的。’他们就开始庆祝。
LUKE|15|25|“那时，大儿子正在田里。他回来，离家不远时，听见奏乐跳舞的声音，
LUKE|15|26|就叫一个僮仆来，问是什么事。
LUKE|15|27|僮仆对他说：‘你弟弟回来了，你父亲因为他无灾无病地回来，把肥牛犊宰了。’
LUKE|15|28|大儿子就生气，不肯进去，他父亲出来劝他。
LUKE|15|29|他对父亲说：‘你看，我服侍你这么多年，从来没有违背过你的命令，而你从来没有给我一只小山羊，叫我和朋友们一同快乐。
LUKE|15|30|但你这个儿子和娼妓吃光了你的财产，他一回来，你倒为他宰了肥牛犊。’
LUKE|15|31|父亲对他说：‘儿啊！你常和我同在，我所有的一切都是你的；
LUKE|15|32|可是你这个弟弟是死而复活，失而复得的，所以我们理当欢喜庆祝。’”
LUKE|16|1|耶稣又对门徒说：“某财主有一个管家，有人向主人告管家浪费他的财物。
LUKE|16|2|主人叫他来，对他说：‘我听到了，你做的是什么事？把你所经管的交代清楚，你不能再作我的管家了。’
LUKE|16|3|那管家心里说：‘主人辞我，不用我再作管家，我将来做什么呢？锄地嘛，没有力气；讨饭嘛，怕羞。
LUKE|16|4|我知道怎么做，好叫人们在我不作管家之后，接我到他们家里去。’
LUKE|16|5|于是他把欠他主人债的，一个一个地叫了来，问头一个说：‘你欠我主人多少？’
LUKE|16|6|他说：‘一百篓 油。’管家对他说：‘拿你的账，快坐下，写五十。’
LUKE|16|7|他问另一个说：‘你欠多少？’他说：‘一百石麦子。’管家对他说：‘拿你的账，写八十。’
LUKE|16|8|主人就夸奖这不义的管家做事精明，因为今世之子应付自己的世代比光明之子更加精明。
LUKE|16|9|我又告诉你们，要藉着那不义的钱财结交朋友，到了钱财无用的时候，他们可以接你们到永远的住处 去。
LUKE|16|10|人在最小的事上忠心，在大事上也忠心；在最小的事上不义，在大事上也不义。
LUKE|16|11|若是你们在不义的钱财上不忠心，谁还把那真实的钱财托付你们呢？
LUKE|16|12|如果你们在别人的东西上不忠心，谁还把你们自己的东西给你们呢？
LUKE|16|13|一个仆人不能服侍两个主；他不是恨这个爱那个，就是重这个轻那个。你们不能又服侍上帝，又服侍 玛门 。”
LUKE|16|14|法利赛人是贪爱钱财的；他们听见这一切话，就嘲笑耶稣。
LUKE|16|15|耶稣对他们说：“你们是在人面前自称为义的，你们的心，上帝却知道；因为人以为尊贵的，是上帝看为可憎恶的。
LUKE|16|16|律法和先知到 约翰 为止，从此上帝国的福音传开了，人人努力要进去。
LUKE|16|17|天地废去比律法的一点一画落空还要容易。
LUKE|16|18|凡休妻另娶的，就是犯奸淫；娶被丈夫休了的妇人的，也是犯奸淫。”
LUKE|16|19|“有一个财主穿着紫色袍和细麻布衣服，天天奢华宴乐。
LUKE|16|20|又有一个讨饭的，名叫 拉撒路 ，浑身长疮，被人放在财主门口，
LUKE|16|21|想得财主桌子上掉下来的碎食充饥，甚至还有狗来舔他的疮。
LUKE|16|22|后来那讨饭的死了，被天使带去放在 亚伯拉罕 的怀里。财主也死了，并且埋葬了。
LUKE|16|23|他在阴间受苦，举目远远地望见 亚伯拉罕 ，又望见 拉撒路 在他怀里，
LUKE|16|24|他就喊着说：‘我祖 亚伯拉罕 哪，可怜我吧！请打发 拉撒路 来，用指头尖蘸点水，凉凉我的舌头，因为我在这火焰里，极其痛苦。’
LUKE|16|25|亚伯拉罕 说：‘孩子啊，你该回想你生前享过福， 拉撒路 也同样受过苦，如今他在这里得安慰，你却受痛苦。
LUKE|16|26|除此之外，在你们和我们之间，有深渊隔开，以致人要从这边过到你们那边是不可能的；要从那边过到这边也是不可能的。’
LUKE|16|27|财主说：‘我祖啊，既然这样，求你打发 拉撒路 到我父家去，
LUKE|16|28|因为我还有五个兄弟，他可以警告他们，免得他们也来到这痛苦的地方。’
LUKE|16|29|亚伯拉罕 说：‘他们有 摩西 和先知的话可以听从。’
LUKE|16|30|他说：‘不！我祖 亚伯拉罕 哪，假如有一个人从死人中到他们那里去，他们一定会悔改。’
LUKE|16|31|亚伯拉罕 对他说：‘如果他们不听从 摩西 和先知的话，就是有人从死人中复活，他们也不会信服的。’”
LUKE|17|1|耶稣又对门徒说：“绊倒人的事是免不了的，但那绊倒人的有祸了！
LUKE|17|2|人若把这些小子中的一个绊倒的，还不如把磨石拴在他的颈项上，丢在海里。
LUKE|17|3|你们要谨慎！若是你的弟兄犯罪，就劝戒他；他若懊悔，就饶恕他。
LUKE|17|4|如果他一天七次得罪你，又七次回头，说：‘我懊悔了’，你总要饶恕他。”
LUKE|17|5|使徒对主说：“请加增我们的信心。”
LUKE|17|6|主说：“你们若有信心像一粒芥菜种，就是对这棵桑树说：‘你要连根拔起，栽在海里’，它也会听从你们。”
LUKE|17|7|“你们当中谁有仆人耕地或是放羊，从田里回来，就对他说‘你快来坐下吃饭’呢？
LUKE|17|8|他岂不对仆人说‘你给我预备晚饭，束上带子伺候我，等我吃喝完了，你才可以吃喝’吗？
LUKE|17|9|仆人照所吩咐的去做，主人还谢谢他吗？
LUKE|17|10|这样，你们做完了一切所吩咐的，要说：‘我们是无用的仆人，所做的本是我们该做的。’”
LUKE|17|11|耶稣往 耶路撒冷 去，经过 撒玛利亚 和 加利利 中间的地区。
LUKE|17|12|他进入一个村子，有十个痲疯病人迎面而来，远远地站着，
LUKE|17|13|高声说：“耶稣，老师啊，可怜我们吧！”
LUKE|17|14|耶稣看见，就对他们说：“你们去，把身体给祭司检查。”他们正去的时候就洁净了。
LUKE|17|15|其中有一个见自己已经好了，就回来大声归荣耀给上帝，
LUKE|17|16|又俯伏在耶稣脚前感谢他。这人是 撒玛利亚 人。
LUKE|17|17|耶稣回答说：“洁净了的不是十个人吗？那九个在哪里呢？
LUKE|17|18|除了这外族人，再没有别人回来归荣耀给上帝吗？”
LUKE|17|19|于是他对那人说：“起来，走吧，你的信救了你！”
LUKE|17|20|法利赛人问：“上帝的国几时来到？”耶稣回答：“上帝的国来到，不是眼睛看得见的。
LUKE|17|21|人也不能说：‘看哪，在这里！’或说：‘在那里！’因为上帝的国就在你们心里 。”
LUKE|17|22|他又对门徒说：“那些日子将到，你们渴望能看见人子的一个日子，却看不见。
LUKE|17|23|有人要对你们说：‘看哪，在那里！’或说：‘看哪，在这里！’你们不要出去，也不要追随他们。
LUKE|17|24|好像闪电从天这边一闪直照到天那边，人子在他的日子 也要这样。
LUKE|17|25|可是他必须先受许多苦，又被这世代所弃绝。
LUKE|17|26|挪亚 的日子怎样，人子的日子也要怎样。
LUKE|17|27|那时，人又吃又喝，又娶又嫁，直到 挪亚 进方舟的那日，洪水就来，把他们全都灭了。
LUKE|17|28|同样，就像在 罗得 的日子，人又吃又喝，又买又卖，又耕种又建造，
LUKE|17|29|到 罗得 离开 所多玛 的那日，有火与硫磺从天上降下来，把他们全都灭了。
LUKE|17|30|人子显现的日子也要这样。
LUKE|17|31|在那日，人在屋顶上，东西在屋里，不要下来拿；人在田里，也不要回家。
LUKE|17|32|你们想想 罗得 的妻子吧！
LUKE|17|33|凡想保全性命的，要丧失性命；凡丧失性命的，要保存性命。
LUKE|17|34|我告诉你们，在那一夜，两个人在一张床上，一个被接去，一个被撇下。
LUKE|17|35|两个女人一同推磨，一个被接去，一个被撇下。 ”
LUKE|17|36|
LUKE|17|37|门徒回答他说：“主啊，在哪里呢？”耶稣对他们说：“尸首在哪里，鹰也会聚在哪里。”
LUKE|18|1|耶稣对门徒讲了一个比喻，为了要他们常常祷告，不可灰心。
LUKE|18|2|他说：“某城有一个官，不惧怕上帝，也不尊重人。
LUKE|18|3|那城里有个寡妇，常到他那里，说：‘我有一个冤家，求你给我伸冤。’
LUKE|18|4|他很久不受理，后来心里说：‘我虽不惧怕上帝，也不尊重人，
LUKE|18|5|只因这寡妇烦扰我，我就给她伸冤吧，免得她常来纠缠我。’”
LUKE|18|6|主说：“你们听这不义的官所说的话。
LUKE|18|7|上帝的选民昼夜呼吁他，他岂会延迟不给他们伸冤吗？
LUKE|18|8|我告诉你们，他很快就要给他们伸冤。然而，人子来的时候，能在世上找到这样的信德吗？”
LUKE|18|9|耶稣向那些自以为义而藐视别人的人讲了这比喻：
LUKE|18|10|“有两个人上圣殿去祷告，一个是法利赛人，一个是税吏。
LUKE|18|11|法利赛人独自站着，自言自语地祷告说：‘上帝啊，我感谢你，我不像别人勒索、不义、奸淫，也不像这个税吏。
LUKE|18|12|我每周禁食两次，凡我所得的都献上十分之一。’
LUKE|18|13|那税吏远远地站着，连举目望天也不敢，只捶着胸，说：‘上帝啊，开恩可怜我这个罪人！’
LUKE|18|14|我告诉你们，这人回家去比那人倒算为义了。因为凡自高的，必降为卑；自甘卑微的，必升为高。”
LUKE|18|15|有人甚至连婴孩也带来见耶稣，要他摸他们，门徒看见就责备那些人。
LUKE|18|16|耶稣却叫他们来，说：“让小孩子到我这里来，不要阻止他们，因为在上帝国的正是这样的人。
LUKE|18|17|我实在告诉你们，凡要接受上帝国的，若不像小孩子，绝不能进去。”
LUKE|18|18|有一个官问耶稣说：“善良的老师，我该做什么事才能承受永生？”
LUKE|18|19|耶稣对他说：“你为什么称我是善良的？除了上帝一位之外，再没有善良的。
LUKE|18|20|诫命你是知道的：‘不可奸淫；不可杀人；不可偷盗；不可作假见证；当孝敬父母。’”
LUKE|18|21|那人说：“这一切我从小都遵守了。”
LUKE|18|22|耶稣听见了，就对他说：“你还缺少一件：要变卖你一切所有的，分给穷人，就必有财宝在天上；你还要来跟从我。”
LUKE|18|23|他听见这些话，就很忧愁，因为他很富有。
LUKE|18|24|耶稣见他变得很忧愁 ，就说：“有钱财的人进上帝的国是何等的难哪！
LUKE|18|25|骆驼穿过针眼比财主进上帝的国还容易呢！”
LUKE|18|26|听见的人说：“这样，谁能得救呢？”
LUKE|18|27|耶稣说：“在人所不能的事，在上帝都能。”
LUKE|18|28|彼得 说：“看哪，我们已经撇下自己所有的跟从你了。”
LUKE|18|29|耶稣对他们说：“我实在告诉你们，凡是为上帝的国撇下房屋，或是妻子、兄弟、父母、儿女的，
LUKE|18|30|没有不在今世得更多倍，而在来世得永生的。”
LUKE|18|31|耶稣把十二使徒带到一边，对他们说：“看哪，我们上 耶路撒冷 去，先知所写的一切事都要成就在人子身上。
LUKE|18|32|他将被交给外邦人；他们要戏弄他，凌辱他，向他吐唾沫，
LUKE|18|33|并要鞭打他，杀害他；第三天他要复活。”
LUKE|18|34|这些事门徒一点也不明白，这话的意思对他们是隐藏的；他们不知道所说的是什么。
LUKE|18|35|耶稣将近 耶利哥 的时候，有一个盲人坐在路旁讨饭。
LUKE|18|36|他听见许多人经过，就问是什么事。
LUKE|18|37|他们告诉他，是 拿撒勒 人耶稣经过。
LUKE|18|38|他就呼叫说：“ 大卫 之子耶稣啊，可怜我吧！”
LUKE|18|39|在前头走的人就责备他，不许他作声，他却越发喊叫：“ 大卫 之子啊，可怜我吧！”
LUKE|18|40|耶稣就站住，吩咐把他领过来，他到了跟前，就问他：
LUKE|18|41|“你要我为你做什么？”他说：“主啊，我要能看见。”
LUKE|18|42|耶稣对他说：“你看见吧！你的信救了你。”
LUKE|18|43|那盲人立刻看得见了，就跟随耶稣，一路归荣耀给上帝。众人看见这事，也都赞美上帝。
LUKE|19|1|耶稣进了 耶利哥 ，要从那里经过。
LUKE|19|2|有一个人名叫 撒该 ，作税吏长，是个财主。
LUKE|19|3|他要看看耶稣是怎样的人，只因人多，他的身材又矮，所以看不见。
LUKE|19|4|于是他跑到前头，爬上桑树，要看耶稣，因为耶稣要从那里经过。
LUKE|19|5|耶稣到了那里，抬头一看，对他说：“ 撒该 ，快下来！今天我必须住在你家里。”
LUKE|19|6|他就急忙下来，欢欢喜喜地接待耶稣。
LUKE|19|7|众人看见，都私下议论说：“他竟然到罪人家里去住宿。”
LUKE|19|8|撒该 站着对主说：“主啊，我把所有的一半给穷人；我若勒索了谁，就还他四倍。”
LUKE|19|9|耶稣对他说：“今天救恩到了这家，因为他也是 亚伯拉罕 的子孙。
LUKE|19|10|人子来是要寻找和拯救失丧的人。”
LUKE|19|11|众人正听见这些话的时候，耶稣因为将近 耶路撒冷 ，又因他们以为上帝的国快要显现，就接着讲了一个比喻，
LUKE|19|12|说：“有一个贵族往远方去，为要取得王位，然后回来。
LUKE|19|13|他叫了自己的十个仆人来，交给他们十锭银子，说：‘你们去做生意，直到我回来。’
LUKE|19|14|他本国的百姓却恨他，打发使者随后去，说：‘我们不愿意这个人作我们的王。’
LUKE|19|15|他得了王位回来，就吩咐叫那领了银子的仆人来，要知道他们做生意赚了多少。
LUKE|19|16|头一个上来，说：‘主啊，你的一锭银子已经赚了十锭。’
LUKE|19|17|主人对他说：‘好，我善良的仆人，你既在最小的事上忠心，你有权柄管十座城。’
LUKE|19|18|第二个来，说：‘主啊，你的一锭银子已经赚了五锭。’
LUKE|19|19|主人也对这个说：‘你管五座城。’
LUKE|19|20|又有一个来说：‘主啊！看哪，你的一锭银子在这里，我把它包在手巾里存着。
LUKE|19|21|我向来怕你，因为你是严厉的人：没有放的，也要去拿；没有种的，也要去收。’
LUKE|19|22|主人对他说：‘你这恶仆，我要凭你的话定你的罪。你既知道我是严厉的人，没有放的也去拿，没有种的也去收，
LUKE|19|23|为什么不把我的银子存在银行，等我来的时候，连本带利都取回来呢？’
LUKE|19|24|于是他对那些站在旁边的人说：‘把他这一锭夺过来，给那有十锭的。’
LUKE|19|25|他们对他说：‘主啊，他已经有十锭了。’
LUKE|19|26|主人说：‘我告诉你们，凡有的，还要给他；没有的，连他所有的也要夺过来。
LUKE|19|27|至于我那些仇敌，不要我作他们王的，把他们拉来，在我面前杀了！’”
LUKE|19|28|耶稣说完了这些话，就走在前面，上 耶路撒冷 去。
LUKE|19|29|快到 伯法其 和 伯大尼 ，在名叫 橄榄山 的地方，他打发两个门徒，
LUKE|19|30|说：“你们往对面村子里去，进去的时候会看见一匹驴驹拴在那里，是从来没有人骑过的，把它解开，牵来。
LUKE|19|31|若有人问为什么解开它，你们就这样说：‘主要用它。’”
LUKE|19|32|被打发的人去了，所遇见的正如耶稣对他们所说的。
LUKE|19|33|他们解开驴驹的时候，主人问他们：“为什么解开驴驹？”
LUKE|19|34|他们说：“主要用它。”
LUKE|19|35|他们把驴驹牵到耶稣那里，把自己的衣服搭在上面，扶耶稣骑上。
LUKE|19|36|他前进的时候，众人把衣服铺在路上。
LUKE|19|37|他将近 耶路撒冷 ，正下 橄榄山 的时候，一大群门徒因所见过的一切异能，都欢呼起来，大声赞美上帝，
LUKE|19|38|说： “奉主名来的王 是应当称颂的！ 在天上有和平； 在至高之处有荣光。”
LUKE|19|39|人群中有几个法利赛人对耶稣说：“老师，责备你的门徒吧！”
LUKE|19|40|耶稣回答：“我告诉你们，若是这些人闭口不说，石头也要呼叫起来。”
LUKE|19|41|耶稣快到 耶路撒冷 ，看见那城，就为它哀哭，
LUKE|19|42|说：“但愿你在这日子知道有关你平安的事，不过这事现在是隐藏的，你的眼睛看不出来。
LUKE|19|43|因为日子将到，你的仇敌要筑起土垒包围你，四面困住你，
LUKE|19|44|并要消灭你和你里头的儿女，连一块石头也不留在另一块石头上，因为你不知道你蒙眷顾的时候。”
LUKE|19|45|耶稣一进圣殿就赶出在里面做买卖的人，
LUKE|19|46|对他们说：“经上说： ‘我的殿是祷告的殿， 你们倒使它成为贼窝了。’”
LUKE|19|47|耶稣天天在圣殿里教导人。祭司长、文士和百姓的领袖都想杀他，
LUKE|19|48|但找不出方法来，因为百姓都侧耳听他。
LUKE|20|1|有一天，耶稣在圣殿里教导百姓，宣讲福音的时候，祭司长、文士和长老上前来，
LUKE|20|2|问他说：“你告诉我们，你仗着什么权柄做这些事？给你这权柄的是谁呢？”
LUKE|20|3|耶稣回答他们：“我也要问你们一句话，你们告诉我。
LUKE|20|4|约翰 的洗礼是从天上来的，还是从人间来的呢？”
LUKE|20|5|他们彼此商量说：“我们若说‘从天上来的’，他会说‘这样，你们为什么不信他呢？’
LUKE|20|6|我们若说‘从人间来的’，所有的百姓都会用石头打死我们，因为他们信 约翰 是先知。”
LUKE|20|7|于是他们回答：“我们不知道是从哪里来的。”
LUKE|20|8|耶稣对他们说：“我也不告诉你们，我仗着什么权柄做这些事。”
LUKE|20|9|耶稣用这个比喻对百姓说：“有人开垦了一个葡萄园，租给园户，就出外远行，去了许久。
LUKE|20|10|到了时候，他打发一个仆人到园户那里去，叫他们把园中当纳的果子交给他；园户竟打了他，叫他空手回去。
LUKE|20|11|园主又打发另一个仆人去，他们也打了他，并且侮辱他，叫他空手回去。
LUKE|20|12|园主又打发第三个仆人去，他们也打伤了他，把他推出去了。
LUKE|20|13|葡萄园主说：‘我要怎么做呢？我要打发我的爱子去，或许他们会尊敬他。’
LUKE|20|14|可是，园户看见他，彼此说：‘这是承受产业的。我们杀了他，产业就归我们了！’
LUKE|20|15|于是他们把他扔出葡萄园外，杀了。这样，葡萄园主要怎么处置他们呢？
LUKE|20|16|他要来除灭那些园户，将葡萄园转给别人。”听见的人说：“绝对不可！”
LUKE|20|17|耶稣看着他们，说：“那么，经上记着： ‘匠人所丢弃的石头 已作了房角的头块石头。’ 这是什么意思呢？
LUKE|20|18|凡跌在那石头上的，一定会跌得粉碎；那石头掉在谁的身上，就要把谁压得稀烂。”
LUKE|20|19|文士和祭司长看出这比喻是指着他们说的，当时就想要下手拿他，只是惧怕百姓。
LUKE|20|20|于是他们窥探耶稣，打发奸细装作好人，要在他的话上抓把柄，好把他交给总督处置。
LUKE|20|21|奸细就问耶稣：“老师，我们知道你所讲所教的都很正确，也不看人的面子，而是诚诚实实传上帝的道。
LUKE|20|22|我们纳税给凯撒合不合法？”
LUKE|20|23|耶稣看出他们的诡诈，就对他们说：
LUKE|20|24|“拿一个银币来给我看。这像和这名号是谁的？”他们说：“是凯撒的。”
LUKE|20|25|耶稣对他们说：“这样，凯撒的归凯撒，上帝的归上帝。”
LUKE|20|26|他们无法当着百姓在他的话上抓到把柄，又因他的对答而惊讶，就闭口不言了。
LUKE|20|27|有些撒都该人来见耶稣。他们说没有复活这回事，于是问耶稣：
LUKE|20|28|“老师， 摩西 为我们写下这话：‘某人的哥哥若死了，有妻无子，他该娶哥哥的妻子，为哥哥生子立后。’
LUKE|20|29|那么，有兄弟七人，第一个娶了妻，没有孩子死了。
LUKE|20|30|第二个、
LUKE|20|31|第三个也娶过她；同样地，七个人都娶过她，没有留下孩子就死了。
LUKE|20|32|后来，那妇人也死了。
LUKE|20|33|那么，在复活的时候，那妇人是哪一个的妻子呢？因为他们七个人都娶过她。”
LUKE|20|34|耶稣对他们说：“这世代的人有娶有嫁，
LUKE|20|35|惟有配得那要来的世代和从死人中复活的人不娶也不嫁。
LUKE|20|36|因为他们不能再死，和天使一样；既然是复活的人，他们就是上帝的儿子。
LUKE|20|37|至于死人复活， 摩西 在《荆棘篇》上就指明了，他称主是 亚伯拉罕 的上帝， 以撒 的上帝， 雅各 的上帝。
LUKE|20|38|上帝不是死人的上帝，而是活人的上帝，因为对他来说，人都是活的。”
LUKE|20|39|有几个文士说：“老师，你说得好。”
LUKE|20|40|以后，他们不敢再问他什么了。
LUKE|20|41|耶稣对他们说：“人们怎么说基督是 大卫 的后裔呢？
LUKE|20|42|《诗篇》 上 大卫 自己说： “主对我主说： ‘你坐在我的右边，
LUKE|20|43|等我使你的仇敌作你的脚凳。’
LUKE|20|44|大卫 既称他为主，他怎么又是 大卫 的后裔呢？”
LUKE|20|45|众百姓听的时候，耶稣对他的门徒说：
LUKE|20|46|“你们要防备文士。他们好穿长袍走来走去，喜欢人们在街市上向他们问安，又喜爱会堂里的高位，宴席上的首座。
LUKE|20|47|他们侵吞寡妇的家产，假意作很长的祷告。这些人要受更重的惩罚！”
LUKE|21|1|耶稣抬头观看，见财主把捐项投入圣殿银库，
LUKE|21|2|又见一个穷寡妇投了两个小文钱 ，
LUKE|21|3|就说：“我实在告诉你们，这穷寡妇所投的比众人更多。
LUKE|21|4|因为众人都是拿有余的捐献，但这寡妇，虽然自己不足，却把一生所有的都投进去了。”
LUKE|21|5|有人谈论圣殿是用美石和供物装饰的，耶稣就说：
LUKE|21|6|“你们所看见的这一切，日子将到，没有一块石头会留在另一块石头上而不被拆毁的。”
LUKE|21|7|他们问他：“老师，什么时候有这些事呢？这些事将临到的时候有什么预兆呢？”
LUKE|21|8|耶稣说：“你们要谨慎，不要受迷惑，因为将有好些人冒我的名来，说‘我是基督’，又说‘时候近了’，你们不要跟从他们！
LUKE|21|9|当你们听见打仗和动乱的事，不要惊惶；因为这些事必须先发生，但终结不会立刻就到。”
LUKE|21|10|于是耶稣对他们说：“民要攻打民，国要攻打国，
LUKE|21|11|将有大地震，多处必有饥荒、瘟疫，又有可怕的异象和大神迹从天上显现。
LUKE|21|12|但这一切的事以前，有人要下手拿你们，迫害你们，把你们交给会堂，并且关在监里，又为我名的缘故拉你们到君王和统治者面前。
LUKE|21|13|但这些事终必成为你们作见证的机会。
LUKE|21|14|所以，你们要立定心意，不要预先考虑怎样申辩；
LUKE|21|15|因为我必赐你们口才和智慧，是你们一切敌人所敌不住、驳不倒的。
LUKE|21|16|连你们的父母、兄弟、亲族、朋友也要把你们交给官府；你们中间也将有被他们害死的。
LUKE|21|17|你们要为我的名被众人憎恨。
LUKE|21|18|然而，你们连一根头发也不会损失。
LUKE|21|19|你们凭着坚忍，就必保全性命。”
LUKE|21|20|“当你们看见 耶路撒冷 被兵围困，就可知道它成为荒芜的日子近了。
LUKE|21|21|那时，在 犹太 的，应当逃到山上；在城里的，应当出来；在乡下的，不要进城。
LUKE|21|22|因为这是报应的日子，要使经上所写的都得应验。
LUKE|21|23|在那些日子，怀孕的和奶孩子的就苦了。因为将有大灾难降在这地方，也有愤怒临到这百姓。
LUKE|21|24|他们要倒在刀下，又被掳到各国去。 耶路撒冷 要被外邦人践踏，直到外邦人的日子满了。”
LUKE|21|25|“日月星辰要显出预兆，地上的邦国也有困苦，因海中波浪的响声而惶惶不安。
LUKE|21|26|人想到那要临到世界的事，就都吓得魂不附体，因为天上的万象都要震动。
LUKE|21|27|那时，他们要看见人子带着能力和大荣耀驾云来临。
LUKE|21|28|一有这些事，你们就当挺身昂首，因为你们得救赎的日子近了。”
LUKE|21|29|耶稣对他们讲了一个比喻说：“你们看无花果树和各样的树，
LUKE|21|30|树叶一长出来，你们看了自然就知道夏天近了。
LUKE|21|31|同样，当你们看见这些事发生，就知道上帝的国近了。
LUKE|21|32|我实在告诉你们，这世代还没有过去，一切都要发生。
LUKE|21|33|天地要废去，我的话却绝不废去。”
LUKE|21|34|“你们要谨慎，免得被贪食、醉酒和今生的忧虑压住你们的心，那日子就忽然临到你们，
LUKE|21|35|如同罗网一样，因为那日子要临到所有居住在地面上的人。
LUKE|21|36|你们要时时警醒，常常祈求，使你们能逃避这一切要来的事，得以站立在人子面前。”
LUKE|21|37|耶稣每日在圣殿里教导人，每夜出城到 橄榄山 住宿。
LUKE|21|38|众百姓清早上圣殿，到耶稣那里听他讲道。
LUKE|22|1|除酵节，又叫逾越节，近了。
LUKE|22|2|祭司长和文士在想法子怎样杀害耶稣，因他们惧怕百姓。
LUKE|22|3|这时，撒但入了那称为 加略 人 犹大 的心。他本是十二使徒里的一个。
LUKE|22|4|他去跟祭司长和守殿官商量怎样把耶稣交给他们。
LUKE|22|5|他们很高兴，就约定给他银子。
LUKE|22|6|他应允了，就找机会，要趁众人不在跟前的时候把耶稣交给他们。
LUKE|22|7|除酵节到了，这一天必须宰逾越节的羔羊。
LUKE|22|8|耶稣打发 彼得 和 约翰 ，说：“你们去为我们预备逾越节的宴席，好让我们吃。”
LUKE|22|9|他们问他：“你要我们在哪里预备？”
LUKE|22|10|耶稣对他们说：“你们进了城，会有人拿着一罐水迎面而来，你们就跟着他，到他所进的房子里去，
LUKE|22|11|对那家的主人说：‘老师问：客房在哪里？我和我的门徒要在那里吃逾越节的宴席。’
LUKE|22|12|他会带你们看一间摆设齐全的楼上大厅，你们就在那里预备。”
LUKE|22|13|他们去了，所看到的正如耶稣所说的。他们就预备了逾越节的宴席。
LUKE|22|14|时候到了，耶稣坐席，使徒们也和他同坐。
LUKE|22|15|耶稣对他们说：“我非常渴望在受害以前和你们吃这逾越节的宴席。
LUKE|22|16|我告诉你们，我不再吃这宴席，直到它实现在上帝的国里。”
LUKE|22|17|耶稣接过杯来，祝谢了，说：“你们拿这杯，大家分着喝。
LUKE|22|18|我告诉你们，从今以后，我不再喝这葡萄汁，直等上帝的国来到。”
LUKE|22|19|他又拿起饼来，祝谢了，就擘开，递给他们，说：“这是我的身体，为你们舍的，你们要如此行，为的是记念我。”
LUKE|22|20|饭后他照样拿起杯来，说：“这杯是用我的血所立的新约，为你们流出来的。
LUKE|22|21|但是，看哪，那出卖我的人的手跟我一同在桌子上。
LUKE|22|22|人子固然要照所预定的离去，但那出卖人子的人有祸了！”
LUKE|22|23|于是他们开始互相追问他们中间哪一个会做这事。
LUKE|22|24|门徒中间也起了争论：他们中哪一个可算为大。
LUKE|22|25|耶稣对他们说：“外邦人有君王为主治理他们，那掌权管他们的称为恩主。
LUKE|22|26|但你们不可这样。你们中间最大的，倒要成为最小的；为领袖的，倒要像服事人的。
LUKE|22|27|是谁为大？是坐席的还是服事人的呢？不是坐席的大吗？然而，我在你们中间是如同服事人的。
LUKE|22|28|“我在试炼之中，常和我同在的就是你们。
LUKE|22|29|我把国赐给你们，正如我父赐给我一样，
LUKE|22|30|使你们在我的国里坐在我的席上吃喝，并且坐在宝座上审判 以色列 十二个支派。”
LUKE|22|31|主又说：“ 西门 ， 西门 ！撒但要得着你们，好筛你们像筛麦子一样；
LUKE|22|32|但我已经为你祈求，使你不至于失了信心。你回头以后，要坚固你的弟兄。”
LUKE|22|33|彼得 对他说：“主啊，我已准备好要同你坐牢，与你同死。”
LUKE|22|34|耶稣说：“ 彼得 ，我告诉你，今日鸡还没有叫，你要三次说不认得我。”
LUKE|22|35|耶稣又对他们说：“我差你们出去的时候，没有钱囊，没有行囊，没有鞋子，你们缺少什么没有？”他们说：“没有。”
LUKE|22|36|耶稣对他们说：“但如今，有钱囊的要带着，有行囊的也一样；没有刀的要卖衣服买刀。
LUKE|22|37|我告诉你们，经上写着说：‘他被列在罪犯之中。’这话必须应验在我身上，因为那关于我的事必然成就。”
LUKE|22|38|他们说：“主啊，请看！这里有两把刀。”耶稣对他们说：“够了。”
LUKE|22|39|耶稣出来，照常往 橄榄山 去，门徒也跟随他。
LUKE|22|40|到了那地方，他就对他们说：“你们要祷告，免得陷入试探。”
LUKE|22|41|于是他离开他们约有一块石头扔出去那么远，跪下祷告，
LUKE|22|42|说：“父啊！你若愿意，求你将这杯撤去；然而，不是照我的意愿，而是要成全你的旨意。” 〔
LUKE|22|43|有一位天使从天上显现，加添他的力量。
LUKE|22|44|耶稣非常痛苦焦虑，祷告更加恳切，汗如大血点滴在地上。 〕
LUKE|22|45|祷告完了，他起来，到门徒那里，见他们因为忧愁都睡着了，
LUKE|22|46|就对他们说：“你们为什么睡觉呢？起来祷告，免得陷入试探！”
LUKE|22|47|耶稣还在说话的时候，来了一群人。十二使徒之一名叫 犹大 的，走在前头，接近耶稣，要亲他。
LUKE|22|48|耶稣对他说：“ 犹大 ，你用亲吻来出卖人子吗？”
LUKE|22|49|左右的人见了要发生的事，就说：“主啊，我们拿刀砍好不好？”
LUKE|22|50|其中有一个人把大祭司的仆人砍了一刀，削掉了他的右耳。
LUKE|22|51|耶稣回答说：“算了，住手吧！”就摸那人的耳朵，把他治好了。
LUKE|22|52|耶稣对那些来抓他的祭司长、守殿官和长老说：“你们带着刀棒出来，如同对付强盗吗？
LUKE|22|53|我天天同你们在圣殿里，你们不下手抓我。现在却是你们的时候，黑暗掌权了。”
LUKE|22|54|他们拿住耶稣，把他带走，进入大祭司的住宅。 彼得 远远地跟着。
LUKE|22|55|他们在院子中间生了火，一同坐着， 彼得 也坐在他们当中。
LUKE|22|56|有一个使女看见 彼得 面向火光坐着，就定睛看他，说：“这个人素来也是同那人一起的。”
LUKE|22|57|彼得 却不承认，说：“你这个女人，我不认得他！”
LUKE|22|58|过了一会儿，又有一个人看见他，说：“你也是他们一伙的。” 彼得 说：“你这个人，我不是！”
LUKE|22|59|约过了一小时，又有一个人坚持说：“他实在是同那人一起的，因为他也是 加利利 人。”
LUKE|22|60|彼得 说：“你这个人，我不知道你在说什么！”正说话之间，鸡就叫了。
LUKE|22|61|主转过身来看 彼得 ， 彼得 就想起主对他所说的话：“今日鸡叫以前，你要三次不认我。”
LUKE|22|62|他就出去痛哭。
LUKE|22|63|看守耶稣的人戏弄他，打他，
LUKE|22|64|又蒙着他的眼，问他：“你说预言吧！打你的是谁？”
LUKE|22|65|他们还用许多别的话辱骂他。
LUKE|22|66|天一亮，民间的众长老、祭司长和文士都聚集，把耶稣带到他们的议会里，
LUKE|22|67|说：“如果你是基督，就告诉我们。”耶稣对他们说：“我若告诉你们，你们也不信；
LUKE|22|68|我若问你们，你们也不回答。
LUKE|22|69|从今以后，人子要坐在权能者上帝的右边。”
LUKE|22|70|他们都说：“那么，你是上帝的儿子了？”耶稣对他们说：“你们说我是。”
LUKE|22|71|他们说：“我们何必再要见证呢？他亲口所说的，我们都亲耳听见了。”
LUKE|23|1|众人都起来，把耶稣解到 彼拉多 面前。
LUKE|23|2|他们开始控告他说：“我们见这人煽惑我们的国民，禁止我们纳税给凯撒，并说自己是基督，是王。”
LUKE|23|3|彼拉多 问耶稣：“你是 犹太 人的王吗？”耶稣回答：“是你说的。”
LUKE|23|4|彼拉多 对祭司长们和众人说：“我查不出这人有什么罪来。”
LUKE|23|5|但他们越发竭力地说：“他煽动百姓，在 犹太 全地传道，从 加利利 起，直到这里了。”
LUKE|23|6|彼拉多 一听见，就问：“这人是 加利利 人吗？”
LUKE|23|7|既知道耶稣属 希律 所管， 彼拉多 就把他送到 希律 那里去。那时 希律 正在 耶路撒冷 。
LUKE|23|8|希律 看见耶稣就非常高兴；因为听见过他的事，早就想要见他，并且指望看他行些神迹，
LUKE|23|9|于是问他许多的话，耶稣却一言不答。
LUKE|23|10|那些祭司长和文士都站着，竭力控告他。
LUKE|23|11|希律 和他的士兵就藐视耶稣，戏弄他，给他穿上华丽的衣服，把他送回 彼拉多 那里去。
LUKE|23|12|从前 希律 和 彼拉多 彼此有仇，在那一天竟成了朋友。
LUKE|23|13|彼拉多 传齐了众祭司长、官长和百姓，
LUKE|23|14|对他们说：“你们解这人到我这里，说他是煽惑百姓的。看哪，我也曾在你们面前审问他，并没有查出这人犯过你们控告他的任何罪；
LUKE|23|15|就是 希律 也是如此，所以把他送回来。可见他没有做什么该死的事。
LUKE|23|16|所以，我要责打他，把他释放。”
LUKE|23|17|
LUKE|23|18|众人却一齐喊着说：“除掉这个人！释放 巴拉巴 给我们！”
LUKE|23|19|这 巴拉巴 是因在城里作乱和杀人而下在监里的。
LUKE|23|20|彼拉多 愿意释放耶稣，就再次向他们讲话。
LUKE|23|21|无奈他们喊着说：“把他钉十字架！把他钉十字架！”
LUKE|23|22|彼拉多 第三次对他们说：“为什么呢？这人做了什么恶事呢？我并没有查出他有什么该死的罪来。所以，我要责打他，把他释放。”
LUKE|23|23|他们大声催逼 彼拉多 ，要求他把耶稣钉十字架；他们的声音终于得胜。
LUKE|23|24|彼拉多 这才照他们的要求定案；
LUKE|23|25|又把他们所要求的那因作乱和杀人而下在监里的人释放了，而把耶稣交给他们，随他们的意思处置。
LUKE|23|26|他们把耶稣带去的时候，有一个 古利奈 人 西门 从乡下来，他们就拿住他，把十字架搁在他身上，叫他背着跟在耶稣后面。
LUKE|23|27|有许多百姓跟随耶稣，其中有好些妇女为他号啕痛哭。
LUKE|23|28|耶稣转身对她们说：“ 耶路撒冷 的女子，不要为我哭，要为你们自己和你们的儿女哭。
LUKE|23|29|因为日子将到，人要说：‘不生育的、未曾怀孕的，和未曾哺乳孩子的有福了！’
LUKE|23|30|那时，人要向大山说： ‘倒在我们身上！’ 向小山说： ‘遮盖我们！’
LUKE|23|31|他们若在树木青绿的时候做这些事，那么在枯干的时候将会怎么样呢？”
LUKE|23|32|另外有两个犯人也被带来和耶稣一同处死。
LUKE|23|33|到了一个地方，名叫髑髅地，他们就在那里把耶稣钉在十字架上，又钉了两个犯人：一个在右边，一个在左边。 〔
LUKE|23|34|这时，耶稣说：“父啊！赦免他们，因为他们所做的，他们不知道。” 〕士兵就抽签分他的衣服。
LUKE|23|35|百姓站在那里观看。官长也嘲笑他，说：“他救了别人，他若是基督，是上帝所拣选的，救救他自己吧！”
LUKE|23|36|士兵也戏弄他，上前拿醋送给他喝，
LUKE|23|37|说：“你若是 犹太 人的王，救救你自己吧！”
LUKE|23|38|在耶稣上方有一个牌子写着：“这是 犹太 人的王。”
LUKE|23|39|同钉的犯人中有一个讥笑他，说：“你不是基督吗？救救你自己和我们吧！”
LUKE|23|40|另一个就应声责备他，说：“你是一样受刑的，还不怕上帝吗？
LUKE|23|41|我们是应得的，因为我们是自作自受，但这个人没有做过一件不对的事。”
LUKE|23|42|他对耶稣说：“耶稣啊，你进入你国的时候，求你记念我。”
LUKE|23|43|耶稣对他说：“我实在告诉你，今日你要同我在乐园里了。”
LUKE|23|44|那时大约是正午，全地都黑暗了，直到下午三点钟，
LUKE|23|45|太阳变黑了，殿的幔子从当中裂为两半。
LUKE|23|46|耶稣大声喊着说：“父啊，我将我的灵交在你手里！”他说了这话，气就断了。
LUKE|23|47|百夫长看见所发生的事，就归荣耀给上帝，说：“这人真是个义人！”
LUKE|23|48|聚集观看这事的众人，见了所发生的事，都捶着胸回去了。
LUKE|23|49|所有与耶稣熟悉的人，和从 加利利 跟着他来的妇女们，都远远地站着，看这些事。
LUKE|23|50|有一个人名叫 约瑟 ，是个议员，为人善良正直，
LUKE|23|51|却没有附从别人的所谋所为。他是 犹太 的 亚利马太城 人，素常盼望着上帝的国。
LUKE|23|52|这人去见 彼拉多 ，请求要耶稣的身体。
LUKE|23|53|他把耶稣的身体取下来，用细麻布裹好，安放在凿岩而成的坟墓里；那坟墓从来没有葬过人。
LUKE|23|54|那日是预备日，安息日快到了。
LUKE|23|55|那些从 加利利 和耶稣同来的妇女跟在后面，看见了坟墓和他的身体怎样安放。
LUKE|23|56|她们就回去，预备了香料香膏。在安息日，她们遵照诫命安息了。
LUKE|24|1|七日的第一日，黎明的时候，那些妇女带着所预备的香料来到坟墓那里，
LUKE|24|2|发现石头已经从坟墓滚开了，
LUKE|24|3|她们就进去，只是不见主耶稣的身体。
LUKE|24|4|正在为这事困惑的时候，忽然有两个人站在旁边，衣服放光。
LUKE|24|5|妇女们非常害怕，就俯伏在地上。那两个人对她们说：“为什么在死人中找活人呢？
LUKE|24|6|他不在这里，已经复活了。要记得他还在 加利利 的时候怎样告诉你们的，
LUKE|24|7|他说：‘人子必须被交在罪人手里，钉在十字架上，第三天复活。’”
LUKE|24|8|她们就想起耶稣的话来。
LUKE|24|9|于是她们从坟墓那里回去，把这一切事告诉十一个使徒和其余的人。
LUKE|24|10|把这些事告诉使徒的有 抹大拉 的 马利亚 、 约亚拿 ，和 雅各 的母亲 马利亚 ，还有跟她们在一起的妇女。
LUKE|24|11|她们这些话，使徒以为是胡言，就不相信。
LUKE|24|12|彼得 起来，跑到坟墓前，俯身往里看，只见细麻布，就回去了，因所发生的事而心里惊讶。
LUKE|24|13|同一天，门徒中有两个人往一个村子去；这村子名叫 以马忤斯 ，离 耶路撒冷 约有二十五里 。
LUKE|24|14|他们彼此谈论所发生的这一切事。
LUKE|24|15|正交谈议论的时候，耶稣亲自走近他们，和他们同行，
LUKE|24|16|可是他们的眼睛模糊了，没认出他。
LUKE|24|17|耶稣对他们说：“你们一边走一边谈，彼此谈论的是什么事呢？”他们就站住，脸上带着愁容。
LUKE|24|18|两人中有一个名叫 革流巴 的回答：“你是在 耶路撒冷 的旅客中，惟一还不知道这几天在那里发生了什么事的人吗？”
LUKE|24|19|耶稣对他们说：“什么事呢？”他们对他说：“就是 拿撒勒 人耶稣的事。他是个先知，在上帝和众百姓面前，说话行事都大有能力。
LUKE|24|20|祭司长们和我们的官长竟把他解去，定了死罪，钉在十字架上。
LUKE|24|21|但我们素来所盼望要救赎 以色列 民的就是他。不但如此，这些事发生到现在已经三天了。
LUKE|24|22|还有，我们中间的几个妇女使我们惊奇：她们清早去了坟墓，
LUKE|24|23|不见他的身体，就回来告诉我们，说她们看见了天使显现，说他活了。
LUKE|24|24|又有我们的几个人往坟墓那里去，所发现的正如妇女们所说的，只是没有看见他。”
LUKE|24|25|耶稣对他们说：“无知的人哪，先知所说的一切话，你们的心信得太迟钝了。
LUKE|24|26|基督不是必须受这些苦难，然后进入他的荣耀吗？”
LUKE|24|27|于是，他从 摩西 和众先知起，凡经上所指着自己的话都给他们作了解释。
LUKE|24|28|他们走近所要去的村子，耶稣好像还要往前走，
LUKE|24|29|他们却强留他说：“时候晚了，天快黑了，请你同我们住下吧。”耶稣就进去，要同他们住下。
LUKE|24|30|坐下来和他们用餐的时候，耶稣拿起饼来，祝福了，擘开，递给他们。
LUKE|24|31|他们的眼睛开了，这才认出他来。耶稣却从他们眼前消失了。
LUKE|24|32|他们彼此说：“在路上他和我们说话，给我们讲解圣经的时候，我们的心在我们里面 岂不是火热的吗？”
LUKE|24|33|于是他们立刻起身，回 耶路撒冷 去，看见十一个使徒和与他们正在一起的人聚集在一处，
LUKE|24|34|说：“主果然复活了，已经显现给 西门 看了。”
LUKE|24|35|于是，两个人把路上所遇到，和耶稣擘饼的时候怎么被他们认出来的事，都述说了一遍。
LUKE|24|36|正说这些话的时候，耶稣亲自站在他们当中，说：“愿你们平安！”
LUKE|24|37|他们却惊慌害怕，以为所看见的是魂。
LUKE|24|38|耶稣对他们说：“你们为什么惊恐不安？为什么心里起疑惑呢？
LUKE|24|39|你们看我的手和我的脚，就知道实在是我了。摸摸我，看，因为魂无骨无肉，你们看，我是有的。”
LUKE|24|40|说了这话，他就把手和脚给他们看。
LUKE|24|41|他们还在又惊又喜、不敢相信的时候，耶稣对他们说：“你们这里有什么吃的没有？”
LUKE|24|42|他们给了他一片烤鱼，
LUKE|24|43|他接过来，在他们面前吃了。
LUKE|24|44|耶稣对他们说：“这就是我从前和你们同在时所告诉你们的话： 摩西 的律法、先知的书，和《 诗篇》 上所记一切指着我的话都必须应验。”
LUKE|24|45|于是耶稣开他们的心窍，使他们能明白圣经，
LUKE|24|46|又对他们说：“照经上所写的，基督必受害，第三天从死人中复活，
LUKE|24|47|并且人们要奉他的名传悔改、使罪得赦的道，从 耶路撒冷 起直传到万邦。
LUKE|24|48|你们就是这些事的见证。
LUKE|24|49|我要将我父所应许的降在你们身上，你们要在城里等候，直到你们领受从上面来的能力。”
LUKE|24|50|耶稣领他们出来，直到 伯大尼 附近，就举手给他们祝福。
LUKE|24|51|正祝福的时候，他离开他们，被带到天上去了。
LUKE|24|52|他们就拜他，带着极大的喜乐回 耶路撒冷 去，
LUKE|24|53|常在圣殿里称颂上帝。
