JUDE|1|1|Jude, a servant of Jesus Christ and a brother of James, To those who have been called, who are loved by God the Father and kept by Jesus Christ:
JUDE|1|2|Mercy, peace and love be yours in abundance.
JUDE|1|3|Dear friends, although I was very eager to write to you about the salvation we share, I felt I had to write and urge you to contend for the faith that was once for all entrusted to the saints.
JUDE|1|4|For certain men whose condemnation was written about long ago have secretly slipped in among you. They are godless men, who change the grace of our God into a license for immorality and deny Jesus Christ our only Sovereign and Lord.
JUDE|1|5|Though you already know all this, I want to remind you that the Lord delivered his people out of Egypt, but later destroyed those who did not believe.
JUDE|1|6|And the angels who did not keep their positions of authority but abandoned their own home--these he has kept in darkness, bound with everlasting chains for judgment on the great Day.
JUDE|1|7|In a similar way, Sodom and Gomorrah and the surrounding towns gave themselves up to sexual immorality and perversion. They serve as an example of those who suffer the punishment of eternal fire.
JUDE|1|8|In the very same way, these dreamers pollute their own bodies, reject authority and slander celestial beings.
JUDE|1|9|But even the archangel Michael, when he was disputing with the devil about the body of Moses, did not dare to bring a slanderous accusation against him, but said, "The Lord rebuke you!"
JUDE|1|10|Yet these men speak abusively against whatever they do not understand; and what things they do understand by instinct, like unreasoning animals--these are the very things that destroy them.
JUDE|1|11|Woe to them! They have taken the way of Cain; they have rushed for profit into Balaam's error; they have been destroyed in Korah's rebellion.
JUDE|1|12|These men are blemishes at your love feasts, eating with you without the slightest qualm--shepherds who feed only themselves. They are clouds without rain, blown along by the wind; autumn trees, without fruit and uprooted--twice dead.
JUDE|1|13|They are wild waves of the sea, foaming up their shame; wandering stars, for whom blackest darkness has been reserved forever.
JUDE|1|14|Enoch, the seventh from Adam, prophesied about these men: "See, the Lord is coming with thousands upon thousands of his holy ones
JUDE|1|15|to judge everyone, and to convict all the ungodly of all the ungodly acts they have done in the ungodly way, and of all the harsh words ungodly sinners have spoken against him."
JUDE|1|16|These men are grumblers and faultfinders; they follow their own evil desires; they boast about themselves and flatter others for their own advantage.
JUDE|1|17|But, dear friends, remember what the apostles of our Lord Jesus Christ foretold.
JUDE|1|18|They said to you, "In the last times there will be scoffers who will follow their own ungodly desires."
JUDE|1|19|These are the men who divide you, who follow mere natural instincts and do not have the Spirit.
JUDE|1|20|But you, dear friends, build yourselves up in your most holy faith and pray in the Holy Spirit.
JUDE|1|21|Keep yourselves in God's love as you wait for the mercy of our Lord Jesus Christ to bring you to eternal life.
JUDE|1|22|Be merciful to those who doubt;
JUDE|1|23|snatch others from the fire and save them; to others show mercy, mixed with fear--hating even the clothing stained by corrupted flesh.
JUDE|1|24|To him who is able to keep you from falling and to present you before his glorious presence without fault and with great joy--
JUDE|1|25|to the only God our Savior be glory, majesty, power and authority, through Jesus Christ our Lord, before all ages, now and forevermore! Amen.
