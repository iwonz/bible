TITUS|1|1|Paul, a servant of God and an apostle of Jesus Christ for the faith of God's elect and the knowledge of the truth that leads to godliness--
TITUS|1|2|a faith and knowledge resting on the hope of eternal life, which God, who does not lie, promised before the beginning of time,
TITUS|1|3|and at his appointed season he brought his word to light through the preaching entrusted to me by the command of God our Savior,
TITUS|1|4|To Titus, my true son in our common faith: Grace and peace from God the Father and Christ Jesus our Savior.
TITUS|1|5|The reason I left you in Crete was that you might straighten out what was left unfinished and appoint elders in every town, as I directed you.
TITUS|1|6|An elder must be blameless, the husband of but one wife, a man whose children believe and are not open to the charge of being wild and disobedient.
TITUS|1|7|Since an overseer is entrusted with God's work, he must be blameless--not overbearing, not quick-tempered, not given to drunkenness, not violent, not pursuing dishonest gain.
TITUS|1|8|Rather he must be hospitable, one who loves what is good, who is self-controlled, upright, holy and disciplined.
TITUS|1|9|He must hold firmly to the trustworthy message as it has been taught, so that he can encourage others by sound doctrine and refute those who oppose it.
TITUS|1|10|For there are many rebellious people, mere talkers and deceivers, especially those of the circumcision group.
TITUS|1|11|They must be silenced, because they are ruining whole households by teaching things they ought not to teach--and that for the sake of dishonest gain.
TITUS|1|12|Even one of their own prophets has said, "Cretans are always liars, evil brutes, lazy gluttons."
TITUS|1|13|This testimony is true. Therefore, rebuke them sharply, so that they will be sound in the faith
TITUS|1|14|and will pay no attention to Jewish myths or to the commands of those who reject the truth.
TITUS|1|15|To the pure, all things are pure, but to those who are corrupted and do not believe, nothing is pure. In fact, both their minds and consciences are corrupted.
TITUS|1|16|They claim to know God, but by their actions they deny him. They are detestable, disobedient and unfit for doing anything good.
TITUS|2|1|You must teach what is in accord with sound doctrine.
TITUS|2|2|Teach the older men to be temperate, worthy of respect, self-controlled, and sound in faith, in love and in endurance.
TITUS|2|3|Likewise, teach the older women to be reverent in the way they live, not to be slanderers or addicted to much wine, but to teach what is good.
TITUS|2|4|Then they can train the younger women to love their husbands and children,
TITUS|2|5|to be self-controlled and pure, to be busy at home, to be kind, and to be subject to their husbands, so that no one will malign the word of God.
TITUS|2|6|Similarly, encourage the young men to be self-controlled.
TITUS|2|7|In everything set them an example by doing what is good. In your teaching show integrity, seriousness
TITUS|2|8|and soundness of speech that cannot be condemned, so that those who oppose you may be ashamed because they have nothing bad to say about us.
TITUS|2|9|Teach slaves to be subject to their masters in everything, to try to please them, not to talk back to them,
TITUS|2|10|and not to steal from them, but to show that they can be fully trusted, so that in every way they will make the teaching about God our Savior attractive.
TITUS|2|11|For the grace of God that brings salvation has appeared to all men.
TITUS|2|12|It teaches us to say "No" to ungodliness and worldly passions, and to live self-controlled, upright and godly lives in this present age,
TITUS|2|13|while we wait for the blessed hope--the glorious appearing of our great God and Savior, Jesus Christ,
TITUS|2|14|who gave himself for us to redeem us from all wickedness and to purify for himself a people that are his very own, eager to do what is good.
TITUS|2|15|These, then, are the things you should teach. Encourage and rebuke with all authority. Do not let anyone despise you.
TITUS|3|1|Remind the people to be subject to rulers and authorities, to be obedient, to be ready to do whatever is good,
TITUS|3|2|to slander no one, to be peaceable and considerate, and to show true humility toward all men.
TITUS|3|3|At one time we too were foolish, disobedient, deceived and enslaved by all kinds of passions and pleasures. We lived in malice and envy, being hated and hating one another.
TITUS|3|4|But when the kindness and love of God our Savior appeared,
TITUS|3|5|he saved us, not because of righteous things we had done, but because of his mercy. He saved us through the washing of rebirth and renewal by the Holy Spirit,
TITUS|3|6|whom he poured out on us generously through Jesus Christ our Savior,
TITUS|3|7|so that, having been justified by his grace, we might become heirs having the hope of eternal life.
TITUS|3|8|This is a trustworthy saying. And I want you to stress these things, so that those who have trusted in God may be careful to devote themselves to doing what is good. These things are excellent and profitable for everyone.
TITUS|3|9|But avoid foolish controversies and genealogies and arguments and quarrels about the law, because these are unprofitable and useless.
TITUS|3|10|Warn a divisive person once, and then warn him a second time. After that, have nothing to do with him.
TITUS|3|11|You may be sure that such a man is warped and sinful; he is self-condemned.
TITUS|3|12|As soon as I send Artemas or Tychicus to you, do your best to come to me at Nicopolis, because I have decided to winter there.
TITUS|3|13|Do everything you can to help Zenas the lawyer and Apollos on their way and see that they have everything they need.
TITUS|3|14|Our people must learn to devote themselves to doing what is good, in order that they may provide for daily necessities and not live unproductive lives.
TITUS|3|15|Everyone with me sends you greetings. Greet those who love us in the faith. Grace be with you all.
