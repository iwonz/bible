JOB|1|1|vir erat in terra Hus nomine Iob et erat vir ille simplex et rectus ac timens Deum et recedens a malo
JOB|1|2|natique sunt ei septem filii et tres filiae
JOB|1|3|et fuit possessio eius septem milia ovium et tria milia camelorum quingenta quoque iuga boum et quingentae asinae ac familia multa nimis eratque vir ille magnus inter omnes Orientales
JOB|1|4|et ibant filii eius et faciebant convivium per domos unusquisque in die suo et mittentes vocabant tres sorores suas ut comederent et biberent cum eis
JOB|1|5|cumque in orbem transissent dies convivii mittebat ad eos Iob et sanctificabat illos consurgensque diluculo offerebat holocausta per singulos dicebat enim ne forte peccaverint filii mei et benedixerint Deo in cordibus suis sic faciebat Iob cunctis diebus
JOB|1|6|quadam autem die cum venissent filii Dei ut adsisterent coram Domino adfuit inter eos etiam Satan
JOB|1|7|cui dixit Dominus unde venis qui respondens ait circuivi terram et perambulavi eam
JOB|1|8|dixitque Dominus ad eum numquid considerasti servum meum Iob quod non sit ei similis in terra homo simplex et rectus et timens Deum ac recedens a malo
JOB|1|9|cui respondens Satan ait numquid frustra timet Iob Deum
JOB|1|10|nonne tu vallasti eum ac domum eius universamque substantiam per circuitum operibus manuum eius benedixisti et possessio illius crevit in terra
JOB|1|11|sed extende paululum manum tuam et tange cuncta quae possidet nisi in facie tua benedixerit tibi
JOB|1|12|dixit ergo Dominus ad Satan ecce universa quae habet in manu tua sunt tantum in eum ne extendas manum tuam egressusque est Satan a facie Domini
JOB|1|13|cum autem quadam die filii et filiae eius comederent et biberent vinum in domo fratris sui primogeniti
JOB|1|14|nuntius venit ad Iob qui diceret boves arabant et asinae pascebantur iuxta eos
JOB|1|15|et inruerunt Sabei tuleruntque omnia et pueros percusserunt gladio et evasi ego solus ut nuntiarem tibi
JOB|1|16|cumque adhuc ille loqueretur venit alter et dixit ignis Dei cecidit e caelo et tactas oves puerosque consumpsit et effugi ego solus ut nuntiarem tibi
JOB|1|17|sed et illo adhuc loquente venit alius et dixit Chaldei fecerunt tres turmas et invaserunt camelos et tulerunt eos necnon et pueros percusserunt gladio et ego fugi solus ut nuntiarem tibi
JOB|1|18|loquebatur ille et ecce alius intravit et dixit filiis tuis et filiabus vescentibus et bibentibus vinum in domo fratris sui primogeniti
JOB|1|19|repente ventus vehemens inruit a regione deserti et concussit quattuor angulos domus quae corruens oppressit liberos tuos et mortui sunt et effugi ego solus ut nuntiarem tibi
JOB|1|20|tunc surrexit Iob et scidit tunicam suam et tonso capite corruens in terram adoravit
JOB|1|21|et dixit nudus egressus sum de utero matris meae et nudus revertar illuc Dominus dedit Dominus abstulit sit nomen Domini benedictum
JOB|1|22|in omnibus his non peccavit Iob neque stultum quid contra Deum locutus est
JOB|2|1|factum est autem cum quadam die venissent filii Dei et starent coram Domino venisset quoque Satan inter eos et staret in conspectu eius
JOB|2|2|ut diceret Dominus ad Satan unde venis qui respondens ait circuivi terram et perambulavi eam
JOB|2|3|et dixit Dominus ad Satan numquid considerasti servum meum Iob quod non sit ei similis in terra vir simplex et rectus timens Deum ac recedens a malo et adhuc retinens innocentiam tu autem commovisti me adversus eum ut adfligerem illum frustra
JOB|2|4|cui respondens Satan ait pellem pro pelle et cuncta quae habet homo dabit pro anima sua
JOB|2|5|alioquin mitte manum tuam et tange os eius et carnem et tunc videbis quod in facie benedicat tibi
JOB|2|6|dixit ergo Dominus ad Satan ecce in manu tua est verumtamen animam illius serva
JOB|2|7|egressus igitur Satan a facie Domini percussit Iob ulcere pessimo a planta pedis usque ad verticem eius
JOB|2|8|qui testa saniem deradebat sedens in sterquilinio
JOB|2|9|dixit autem illi uxor sua adhuc tu permanes in simplicitate tua benedic Deo et morere
JOB|2|10|qui ait ad illam quasi una de stultis locuta es si bona suscepimus de manu Domini quare mala non suscipiamus in omnibus his non peccavit Iob labiis suis
JOB|2|11|igitur audientes tres amici Iob omne malum quod accidisset ei venerunt singuli de loco suo Eliphaz Themanites et Baldad Suites et Sophar Naamathites condixerant enim ut pariter venientes visitarent eum et consolarentur
JOB|2|12|cumque levassent procul oculos suos non cognoverunt eum et exclamantes ploraverunt scissisque vestibus sparserunt pulverem super caput suum in caelum
JOB|2|13|et sederunt cum eo in terram septem diebus et septem noctibus et nemo loquebatur ei verbum videbant enim dolorem esse vehementem
JOB|3|1|post haec aperuit Iob os suum et maledixit diei suo
JOB|3|2|et locutus est
JOB|3|3|pereat dies in qua natus sum et nox in qua dictum est conceptus est homo
JOB|3|4|dies ille vertatur in tenebras non requirat eum Deus desuper et non inlustret lumine
JOB|3|5|obscurent eum tenebrae et umbra mortis occupet eum caligo et involvatur amaritudine
JOB|3|6|noctem illam tenebrosus turbo possideat non conputetur in diebus anni nec numeretur in mensibus
JOB|3|7|sit nox illa solitaria nec laude digna
JOB|3|8|maledicant ei qui maledicunt diei qui parati sunt suscitare Leviathan
JOB|3|9|obtenebrentur stellae caligine eius expectet lucem et non videat nec ortum surgentis aurorae
JOB|3|10|quia non conclusit ostia ventris qui portavit me nec abstulit mala ab oculis meis
JOB|3|11|quare non in vulva mortuus sum egressus ex utero non statim perii
JOB|3|12|quare exceptus genibus cur lactatus uberibus
JOB|3|13|nunc enim dormiens silerem et somno meo requiescerem
JOB|3|14|cum regibus et consulibus terrae qui aedificant sibi solitudines
JOB|3|15|aut cum principibus qui possident aurum et replent domos suas argento
JOB|3|16|aut sicut abortivum absconditum non subsisterem vel qui concepti non viderunt lucem
JOB|3|17|ibi impii cessaverunt a tumultu et ibi requieverunt fessi robore
JOB|3|18|et quondam vincti pariter sine molestia non audierunt vocem exactoris
JOB|3|19|parvus et magnus ibi sunt et servus liber a domino suo
JOB|3|20|quare data est misero lux et vita his qui in amaritudine animae sunt
JOB|3|21|qui expectant mortem et non venit quasi effodientes thesaurum
JOB|3|22|gaudentque vehementer cum invenerint sepulchrum
JOB|3|23|viro cuius abscondita est via et circumdedit eum Deus tenebris
JOB|3|24|antequam comedam suspiro et quasi inundantes aquae sic rugitus meus
JOB|3|25|quia timor quem timebam evenit mihi et quod verebar accidit
JOB|3|26|nonne dissimulavi nonne silui nonne quievi et venit super me indignatio
JOB|4|1|respondens autem Eliphaz Themanites dixit
JOB|4|2|si coeperimus loqui tibi forsitan moleste accipias sed conceptum sermonem tenere quis possit
JOB|4|3|ecce docuisti multos et manus lassas roborasti
JOB|4|4|vacillantes confirmaverunt sermones tui et genua trementia confortasti
JOB|4|5|nunc autem venit super te plaga et defecisti tetigit te et conturbatus es
JOB|4|6|timor tuus fortitudo tua patientia tua et perfectio viarum tuarum
JOB|4|7|recordare obsecro te quis umquam innocens perierit aut quando recti deleti sint
JOB|4|8|quin potius vidi eos qui operantur iniquitatem et seminant dolores et metunt eos
JOB|4|9|flante Deo perisse et spiritu irae eius esse consumptos
JOB|4|10|rugitus leonis et vox leaenae et dentes catulorum leonum contriti sunt
JOB|4|11|tigris periit eo quod non haberet praedam et catuli leonis dissipati sunt
JOB|4|12|porro ad me dictum est verbum absconditum et quasi furtive suscepit auris mea venas susurri eius
JOB|4|13|in horrore visionis nocturnae quando solet sopor occupare homines
JOB|4|14|pavor tenuit me et tremor et omnia ossa mea perterrita sunt
JOB|4|15|et cum spiritus me praesente transiret inhorruerunt pili carnis meae
JOB|4|16|stetit quidam cuius non agnoscebam vultum imago coram oculis meis et vocem quasi aurae lenis audivi
JOB|4|17|numquid homo Dei conparatione iustificabitur aut factore suo purior erit vir
JOB|4|18|ecce qui serviunt ei non sunt stabiles et in angelis suis repperit pravitatem
JOB|4|19|quanto magis hii qui habitant domos luteas qui terrenum habent fundamentum consumentur velut a tinea
JOB|4|20|de mane usque ad vesperum succidentur et quia nullus intellegit in aeternum peribunt
JOB|4|21|qui autem reliqui fuerint auferentur ex eis morientur et non in sapientia
JOB|5|1|voca ergo si est qui tibi respondeat et ad aliquem sanctorum convertere
JOB|5|2|vere stultum interficit iracundia et parvulum occidit invidia
JOB|5|3|ego vidi stultum firma radice et maledixi pulchritudini eius statim
JOB|5|4|longe fient filii eius a salute et conterentur in porta et non erit qui eruat
JOB|5|5|cuius messem famelicus comedet et ipsum rapiet armatus et ebibent sitientes divitias eius
JOB|5|6|nihil in terra sine causa fit et de humo non orietur dolor
JOB|5|7|homo ad laborem nascitur et avis ad volatum
JOB|5|8|quam ob rem ego deprecabor Dominum et ad Deum ponam eloquium meum
JOB|5|9|qui facit magna et inscrutabilia et mirabilia absque numero
JOB|5|10|qui dat pluviam super faciem terrae et inrigat aquis universa
JOB|5|11|qui ponit humiles in sublimi et maerentes erigit sospitate
JOB|5|12|qui dissipat cogitationes malignorum ne possint implere manus eorum quod coeperant
JOB|5|13|qui adprehendit sapientes in astutia eorum et consilium pravorum dissipat
JOB|5|14|per diem incurrent tenebras et quasi in nocte sic palpabunt in meridie
JOB|5|15|porro salvum faciet a gladio oris eorum et de manu violenti pauperem
JOB|5|16|et erit egeno spes iniquitas autem contrahet os suum
JOB|5|17|beatus homo qui corripitur a Domino increpationem ergo Domini ne reprobes
JOB|5|18|quia ipse vulnerat et medetur percutit et manus eius sanabunt
JOB|5|19|in sex tribulationibus liberabit te et in septima non tanget te malum
JOB|5|20|in fame eruet te de morte et in bello de manu gladii
JOB|5|21|a flagello linguae absconderis et non timebis calamitatem cum venerit
JOB|5|22|in vastitate et fame ridebis et bestiam terrae non formidabis
JOB|5|23|sed cum lapidibus regionum pactum tuum et bestiae terrae pacificae erunt tibi
JOB|5|24|et scies quod pacem habeat tabernaculum tuum et visitans speciem tuam non peccabis
JOB|5|25|scies quoque quoniam multiplex erit semen tuum et progenies tua quasi herba terrae
JOB|5|26|ingredieris in abundantia sepulchrum sicut infertur acervus in tempore suo
JOB|5|27|ecce hoc ut investigavimus ita est quod auditum mente pertracta
JOB|6|1|respondens autem Iob dixit
JOB|6|2|utinam adpenderentur peccata mea quibus iram merui et calamitas quam patior in statera
JOB|6|3|quasi harena maris haec gravior appareret unde et verba mea dolore sunt plena
JOB|6|4|quia sagittae Domini in me sunt quarum indignatio ebibit spiritum meum et terrores Domini militant contra me
JOB|6|5|numquid rugiet onager cum habuerit herbam aut mugiet bos cum ante praesepe plenum steterit
JOB|6|6|aut poterit comedi insulsum quod non est sale conditum aut potest aliquis gustare quod gustatum adfert mortem
JOB|6|7|quae prius tangere nolebat anima mea nunc prae angustia cibi mei sunt
JOB|6|8|quis det ut veniat petitio mea et quod expecto tribuat mihi Deus
JOB|6|9|et qui coepit ipse me conterat solvat manum suam et succidat me
JOB|6|10|et haec mihi sit consolatio ut adfligens me dolore non parcat nec contradicam sermonibus Sancti
JOB|6|11|quae est enim fortitudo mea ut sustineam aut quis finis meus ut patienter agam
JOB|6|12|nec fortitudo lapidum fortitudo mea nec caro mea aerea est
JOB|6|13|ecce non est auxilium mihi in me et necessarii quoque mei recesserunt a me
JOB|6|14|qui tollit ab amico suo misericordiam timorem Domini derelinquit
JOB|6|15|fratres mei praeterierunt me sicut torrens qui raptim transit in convallibus
JOB|6|16|qui timent pruinam inruet super eos nix
JOB|6|17|tempore quo fuerint dissipati peribunt et ut incaluerit solventur de loco suo
JOB|6|18|involutae sunt semitae gressuum eorum ambulabunt in vacuum et peribunt
JOB|6|19|considerate semitas Theman itinera Saba et expectate paulisper
JOB|6|20|confusi sunt quia speravi venerunt quoque usque ad me et pudore cooperti sunt
JOB|6|21|nunc venistis et modo videntes plagam meam timetis
JOB|6|22|numquid dixi adferte mihi et de substantia vestra donate mihi
JOB|6|23|vel liberate me de manu hostis et de manu robustorum eruite me
JOB|6|24|docete me et ego tacebo et si quid forte ignoravi instruite me
JOB|6|25|quare detraxistis sermonibus veritatis cum e vobis nullus sit qui possit arguere
JOB|6|26|ad increpandum tantum eloquia concinnatis et in ventum verba profertis
JOB|6|27|super pupillum inruitis et subvertere nitimini amicum vestrum
JOB|6|28|verumtamen quod coepistis explete praebete aurem et videte an mentiar
JOB|6|29|respondete obsecro absque contentione et loquentes id quod iustum est iudicate
JOB|6|30|et non invenietis in lingua mea iniquitatem nec in faucibus meis stultitia personabit
JOB|7|1|militia est vita hominis super terram et sicut dies mercennarii dies eius
JOB|7|2|sicut servus desiderat umbram et sicut mercennarius praestolatur finem operis sui
JOB|7|3|sic et ego habui menses vacuos et noctes laboriosas enumeravi mihi
JOB|7|4|si dormiero dico quando consurgam et rursum expectabo vesperam et replebor doloribus usque ad tenebras
JOB|7|5|induta est caro mea putredine et sordibus pulveris cutis mea aruit et contracta est
JOB|7|6|dies mei velocius transierunt quam a texente tela succiditur et consumpti sunt absque ulla spe
JOB|7|7|memento quia ventus est vita mea et non revertetur oculus meus ut videat bona
JOB|7|8|nec aspiciet me visus hominis oculi tui in me et non subsistam
JOB|7|9|sicut consumitur nubes et pertransit sic qui descenderit ad inferos non ascendet
JOB|7|10|nec revertetur ultra in domum suam neque cognoscet eum amplius locus eius
JOB|7|11|quapropter et ego non parcam ori meo loquar in tribulatione spiritus mei confabulabor cum amaritudine animae meae
JOB|7|12|numquid mare sum ego aut cetus quia circumdedisti me carcere
JOB|7|13|si dixero consolabitur me lectulus meus et relevabor loquens mecum in strato meo
JOB|7|14|terrebis me per somnia et per visiones horrore concuties
JOB|7|15|quam ob rem elegit suspendium anima mea et mortem ossa mea
JOB|7|16|desperavi nequaquam ultra iam vivam parce mihi nihil enim sunt dies mei
JOB|7|17|quid est homo quia magnificas eum aut quia ponis erga eum cor tuum
JOB|7|18|visitas eum diluculo et subito probas illum
JOB|7|19|usquequo non parces mihi nec dimittis me ut gluttiam salivam meam
JOB|7|20|peccavi quid faciam tibi o custos hominum quare posuisti me contrarium tibi et factus sum mihimet ipsi gravis
JOB|7|21|cur non tolles peccatum meum et quare non auferes iniquitatem meam ecce nunc in pulvere dormiam et si mane me quaesieris non subsistam
JOB|8|1|respondens autem Baldad Suites dixit
JOB|8|2|usquequo loqueris talia et spiritus multiplex sermones oris tui
JOB|8|3|numquid Deus subplantat iudicium et Omnipotens subvertit quod iustum est
JOB|8|4|etiam si filii tui peccaverunt ei et dimisit eos in manu iniquitatis suae
JOB|8|5|tu tamen si diluculo consurrexeris ad Deum et Omnipotentem fueris deprecatus
JOB|8|6|si mundus et rectus incesseris statim evigilabit ad te et pacatum reddet habitaculum iustitiae tuae
JOB|8|7|in tantum ut priora tua fuerint parva et novissima tua multiplicentur nimis
JOB|8|8|interroga enim generationem pristinam et diligenter investiga patrum memoriam
JOB|8|9|hesterni quippe sumus et ignoramus quoniam sicut umbra dies nostri sunt super terram
JOB|8|10|et ipsi docebunt te loquentur tibi et de corde suo proferent eloquia
JOB|8|11|numquid vivere potest scirpus absque humore aut crescet carectum sine aqua
JOB|8|12|cum adhuc sit in flore nec carpatur manu ante omnes herbas arescit
JOB|8|13|sic viae omnium qui obliviscuntur Deum et spes hypocritae peribit
JOB|8|14|non ei placebit vecordia sua et sicut tela aranearum fiducia eius
JOB|8|15|innitetur super domum suam et non stabit fulciet eam et non consurget
JOB|8|16|humectus videtur antequam veniat sol et in horto suo germen eius egreditur
JOB|8|17|super acervum petrarum radices eius densabuntur et inter lapides commorabitur
JOB|8|18|si absorbuerit eum de loco suo negabit eum et dicet non novi te
JOB|8|19|haec est enim laetitia viae eius ut rursum de terra alii germinentur
JOB|8|20|Deus non proiciet simplicem nec porriget manum malignis
JOB|8|21|donec impleatur risu os tuum et labia tua iubilo
JOB|8|22|qui oderunt te induentur confusione et tabernaculum impiorum non subsistet
JOB|9|1|et respondens Iob ait
JOB|9|2|vere scio quod ita sit et quod non iustificetur homo conpositus Deo
JOB|9|3|si voluerit contendere cum eo non poterit ei respondere unum pro mille
JOB|9|4|sapiens corde est et fortis robore quis restitit ei et pacem habuit
JOB|9|5|qui transtulit montes et nescierunt hii quos subvertit in furore suo
JOB|9|6|qui commovet terram de loco suo et columnae eius concutiuntur
JOB|9|7|qui praecipit soli et non oritur et stellas claudit quasi sub signaculo
JOB|9|8|qui extendit caelos solus et graditur super fluctus maris
JOB|9|9|qui facit Arcturum et Oriona et Hyadas et interiora austri
JOB|9|10|qui facit magna et inconprehensibilia et mirabilia quorum non est numerus
JOB|9|11|si venerit ad me non videbo si abierit non intellegam eum
JOB|9|12|si repente interroget quis respondebit ei vel quis dicere potest cur facis
JOB|9|13|Deus cuius resistere irae nemo potest et sub quo curvantur qui portant orbem
JOB|9|14|quantus ergo sum ego qui respondeam ei et loquar verbis meis cum eo
JOB|9|15|qui etiam si habuero quippiam iustum non respondebo sed meum iudicem deprecabor
JOB|9|16|et cum invocantem exaudierit me non credo quod audierit vocem meam
JOB|9|17|in turbine enim conteret me et multiplicabit vulnera mea etiam sine causa
JOB|9|18|non concedit requiescere spiritum meum et implet me amaritudinibus
JOB|9|19|si fortitudo quaeritur robustissimus est si aequitas iudicii nemo pro me audet testimonium dicere
JOB|9|20|si iustificare me voluero os meum condemnabit me si innocentem ostendere pravum me conprobabit
JOB|9|21|etiam si simplex fuero hoc ipsum ignorabit anima mea et taedebit me vitae meae
JOB|9|22|unum est quod locutus sum et innocentem et impium ipse consumit
JOB|9|23|si flagellat occidat semel et non de poenis innocentum rideat
JOB|9|24|terra data est in manu impii vultum iudicum eius operit quod si non ille est quis ergo est
JOB|9|25|dies mei velociores fuerunt cursore fugerunt et non viderunt bonum
JOB|9|26|pertransierunt quasi naves poma portantes sicut aquila volans ad escam
JOB|9|27|cum dixero nequaquam ita loquar commuto faciem meam et dolore torqueor
JOB|9|28|verebar omnia opera mea sciens quod non parceres delinquenti
JOB|9|29|si autem et sic impius sum quare frustra laboravi
JOB|9|30|si lotus fuero quasi aquis nivis et fulserint velut mundissimae manus meae
JOB|9|31|tamen sordibus intingues me et abominabuntur me vestimenta mea
JOB|9|32|neque enim viro qui similis mei est respondebo nec qui mecum in iudicio ex aequo possit audiri
JOB|9|33|non est qui utrumque valeat arguere et ponere manum suam in ambobus
JOB|9|34|auferat a me virgam suam et pavor eius non me terreat
JOB|9|35|loquar et non timebo eum neque enim possum metuens respondere
JOB|10|1|taedet animam meam vitae meae dimittam adversum me eloquium meum loquar in amaritudine animae meae
JOB|10|2|dicam Deo noli me condemnare indica mihi cur me ita iudices
JOB|10|3|numquid bonum tibi videtur si calumnieris et opprimas me opus manuum tuarum et consilium impiorum adiuves
JOB|10|4|numquid oculi carnei tibi sunt aut sicut videt homo et tu videbis
JOB|10|5|numquid sicut dies hominis dies tui et anni tui sicut humana sunt tempora
JOB|10|6|ut quaeras iniquitatem meam et peccatum meum scruteris
JOB|10|7|et scias quia nihil impium fecerim cum sit nemo qui de manu tua possit eruere
JOB|10|8|manus tuae plasmaverunt me et fecerunt me totum in circuitu et sic repente praecipitas me
JOB|10|9|memento quaeso quod sicut lutum feceris me et in pulverem reduces me
JOB|10|10|nonne sicut lac mulsisti me et sicut caseum me coagulasti
JOB|10|11|pelle et carnibus vestisti me et ossibus et nervis conpegisti me
JOB|10|12|vitam et misericordiam tribuisti mihi et visitatio tua custodivit spiritum meum
JOB|10|13|licet haec celes in corde tuo tamen scio quia universorum memineris
JOB|10|14|si peccavi et ad horam pepercisti mihi cur ab iniquitate mea mundum me esse non pateris
JOB|10|15|et si impius fuero vae mihi est et si iustus non levabo caput saturatus adflictione et miseria
JOB|10|16|et propter superbiam quasi leaenam capies me reversusque mirabiliter me crucias
JOB|10|17|instauras testes tuos contra me et multiplicas iram tuam adversum me et poenae militant in me
JOB|10|18|quare de vulva eduxisti me qui utinam consumptus essem ne oculus me videret
JOB|10|19|fuissem quasi qui non essem de utero translatus ad tumulum
JOB|10|20|numquid non paucitas dierum meorum finietur brevi dimitte ergo me ut plangam paululum dolorem meum
JOB|10|21|antequam vadam et non revertar ad terram tenebrosam et opertam mortis caligine
JOB|10|22|terram miseriae et tenebrarum ubi umbra mortis et nullus ordo et sempiternus horror inhabitans
JOB|11|1|respondens autem Sophar Naamathites dixit
JOB|11|2|numquid qui multa loquitur non et audiet aut vir verbosus iustificabitur
JOB|11|3|tibi soli tacebunt homines et cum ceteros inriseris a nullo confutaberis
JOB|11|4|dixisti enim purus est sermo meus et mundus sum in conspectu tuo
JOB|11|5|atque utinam Deus loqueretur tecum et aperiret labia sua tibi
JOB|11|6|ut ostenderet tibi secreta sapientiae et quod multiplex esset lex eius et intellegeres quod multo minora exigaris a Deo quam meretur iniquitas tua
JOB|11|7|forsitan vestigia Dei conprehendes et usque ad perfectum Omnipotentem repperies
JOB|11|8|excelsior caelo est et quid facies profundior inferno et unde cognosces
JOB|11|9|longior terrae mensura eius et latior mari
JOB|11|10|si subverterit omnia vel in unum coartaverit quis contradicet ei
JOB|11|11|ipse enim novit hominum vanitatem et videns iniquitatem nonne considerat
JOB|11|12|vir vanus in superbiam erigitur et tamquam pullum onagri se liberum natum putat
JOB|11|13|tu autem firmasti cor tuum et expandisti ad eum manus tuas
JOB|11|14|si iniquitatem quod est in manu tua abstuleris a te et non manserit in tabernaculo tuo iniustitia
JOB|11|15|tum levare poteris faciem tuam absque macula et eris stabilis et non timebis
JOB|11|16|miseriae quoque oblivisceris et quasi aquarum quae praeterierint recordaberis
JOB|11|17|et quasi meridianus fulgor consurget tibi ad vesperam et cum te consumptum putaveris orieris ut lucifer
JOB|11|18|et habebis fiduciam proposita tibi spe et defossus securus dormies
JOB|11|19|requiesces et non erit qui te exterreat et deprecabuntur faciem tuam plurimi
JOB|11|20|oculi autem impiorum deficient et effugium peribit ab eis et spes eorum abominatio animae
JOB|12|1|respondens autem Iob dixit
JOB|12|2|ergo vos estis soli homines et vobiscum morietur sapientia
JOB|12|3|et mihi est cor sicut et vobis nec inferior vestri sum quis enim haec quae nostis ignorat
JOB|12|4|qui deridetur ab amico suo sicut ego invocabit Deum et exaudiet eum deridetur enim iusti simplicitas
JOB|12|5|lampas contempta apud cogitationes divitum parata ad tempus statutum
JOB|12|6|abundant tabernacula praedonum et audacter provocant Deum cum ipse dederit omnia in manibus eorum
JOB|12|7|nimirum interroga iumenta et docebunt te et volatilia caeli et indicabunt tibi
JOB|12|8|loquere terrae et respondebit tibi et narrabunt pisces maris
JOB|12|9|quis ignorat quod omnia haec manus Domini fecerit
JOB|12|10|in cuius manu anima omnis viventis et spiritus universae carnis hominis
JOB|12|11|nonne auris verba diiudicat et fauces comedentis saporem
JOB|12|12|in antiquis est sapientia et in multo tempore prudentia
JOB|12|13|apud ipsum est sapientia et fortitudo ipse habet consilium et intellegentiam
JOB|12|14|si destruxerit nemo est qui aedificet et si incluserit hominem nullus est qui aperiat
JOB|12|15|si continuerit aquas omnia siccabuntur et si emiserit eas subvertent terram
JOB|12|16|apud ipsum est fortitudo et sapientia ipse novit et decipientem et eum qui decipitur
JOB|12|17|adducit consiliarios in stultum finem et iudices in stuporem
JOB|12|18|balteum regum dissolvit et praecingit fune renes eorum
JOB|12|19|ducit sacerdotes inglorios et optimates subplantat
JOB|12|20|commutans labium veracium et doctrinam senum auferens
JOB|12|21|effundit despectionem super principes et eos qui oppressi fuerant relevans
JOB|12|22|qui revelat profunda de tenebris et producit in lucem umbram mortis
JOB|12|23|qui multiplicat gentes et perdet eas et subversas in integrum restituet
JOB|12|24|qui inmutat cor principum populi terrae et decipit eos ut frustra incedant per invium
JOB|12|25|palpabunt quasi in tenebris et non in luce et errare eos faciet quasi ebrios
JOB|13|1|ecce omnia et vidit oculus meus et audivit auris mea et intellexi singula
JOB|13|2|secundum scientiam vestram et ego novi nec inferior vestri sum
JOB|13|3|sed tamen ad Omnipotentem loquar et disputare cum Deo cupio
JOB|13|4|prius vos ostendens fabricatores mendacii et cultores perversorum dogmatum
JOB|13|5|atque utinam taceretis ut putaremini esse sapientes
JOB|13|6|audite ergo correptiones meas et iudicium labiorum meorum adtendite
JOB|13|7|numquid Deus indiget vestro mendacio ut pro illo loquamini dolos
JOB|13|8|numquid faciem eius accipitis et pro Deo iudicare nitimini
JOB|13|9|aut placebit ei quem celare nihil potest aut decipietur ut homo vestris fraudulentiis
JOB|13|10|ipse vos arguet quoniam in abscondito faciem eius accipitis
JOB|13|11|statim ut se commoverit turbabit vos et terror eius inruet super vos
JOB|13|12|memoria vestra conparabitur cineri et redigentur in lutum cervices vestrae
JOB|13|13|tacete paulisper ut loquar quodcumque mihi mens suggesserit
JOB|13|14|quare lacero carnes meas dentibus meis et animam meam porto in manibus meis
JOB|13|15|etiam si occiderit me in ipso sperabo verumtamen vias meas in conspectu eius arguam
JOB|13|16|et ipse erit salvator meus non enim veniet in conspectu eius omnis hypocrita
JOB|13|17|audite sermonem meum et enigmata percipite auribus vestris
JOB|13|18|si fuero iudicatus scio quod iustus inveniar
JOB|13|19|quis est qui iudicetur mecum veniat quare tacens consumor
JOB|13|20|duo tantum ne facias mihi et tunc a facie tua non abscondar
JOB|13|21|manum tuam longe fac a me et formido tua non me terreat
JOB|13|22|et voca me et respondebo tibi aut certe loquar et tu responde mihi
JOB|13|23|quantas habeo iniquitates et peccata scelera mea et delicta ostende mihi
JOB|13|24|cur faciem tuam abscondis et arbitraris me inimicum tuum
JOB|13|25|contra folium quod vento rapitur ostendis potentiam tuam et stipulam siccam persequeris
JOB|13|26|scribis enim contra me amaritudines et consumere me vis peccatis adulescentiae meae
JOB|13|27|posuisti in nervo pedem meum et observasti omnes semitas meas et vestigia pedum meorum considerasti
JOB|13|28|qui quasi putredo consumendus sum et quasi vestimentum quod comeditur a tinea
JOB|14|1|homo natus de muliere brevi vivens tempore repletus multis miseriis
JOB|14|2|quasi flos egreditur et conteritur et fugit velut umbra et numquam in eodem statu permanet
JOB|14|3|et dignum ducis super huiuscemodi aperire oculos tuos et adducere eum tecum in iudicium
JOB|14|4|quis potest facere mundum de inmundo conceptum semine nonne tu qui solus es
JOB|14|5|breves dies hominis sunt numerus mensuum eius apud te est constituisti terminos eius qui praeterire non poterunt
JOB|14|6|recede paululum ab eo ut quiescat donec optata veniat sicut mercennarii dies eius
JOB|14|7|lignum habet spem si praecisum fuerit rursum virescit et rami eius pullulant
JOB|14|8|si senuerit in terra radix eius et in pulvere emortuus fuerit truncus illius
JOB|14|9|ad odorem aquae germinabit et faciet comam quasi cum primum plantatum est
JOB|14|10|homo vero cum mortuus fuerit et nudatus atque consumptus ubi quaeso est
JOB|14|11|quomodo si recedant aquae de mari et fluvius vacuefactus arescat
JOB|14|12|sic homo cum dormierit non resurget donec adteratur caelum non evigilabit nec consurget de somno suo
JOB|14|13|quis mihi hoc tribuat ut in inferno protegas me ut abscondas me donec pertranseat furor tuus et constituas mihi tempus in quo recorderis mei
JOB|14|14|putasne mortuus homo rursum vivet cunctis diebus quibus nunc milito expecto donec veniat inmutatio mea
JOB|14|15|vocabis et ego respondebo tibi operi manuum tuarum porriges dexteram
JOB|14|16|tu quidem gressus meos dinumerasti sed parces peccatis meis
JOB|14|17|signasti quasi in sacculo delicta mea sed curasti iniquitatem meam
JOB|14|18|mons cadens defluet et saxum transfertur de loco suo
JOB|14|19|lapides excavant aquae et adluvione paulatim terra consumitur et homines ergo similiter perdes
JOB|14|20|roborasti eum paululum ut in perpetuum pertransiret inmutabis faciem eius et emittes eum
JOB|14|21|sive nobiles fuerint filii eius sive ignobiles non intelleget
JOB|14|22|attamen caro eius dum vivet dolebit et anima illius super semet ipso lugebit
JOB|15|1|respondens autem Eliphaz Themanites dixit
JOB|15|2|numquid sapiens respondebit quasi in ventum loquens et implebit ardore stomachum suum
JOB|15|3|arguis verbis eum qui non est aequalis tui et loqueris quod tibi non expedit
JOB|15|4|quantum in te est evacuasti timorem et tulisti preces coram Deo
JOB|15|5|docuit enim iniquitas tua os tuum et imitaris linguam blasphemantium
JOB|15|6|condemnabit te os tuum et non ego et labia tua respondebunt tibi
JOB|15|7|numquid primus homo tu natus es et ante colles formatus
JOB|15|8|numquid consilium Dei audisti et inferior te erit eius sapientia
JOB|15|9|quid nosti quod ignoremus quid intellegis quod nesciamus
JOB|15|10|et senes et antiqui sunt in nobis multo vetustiores quam patres tui
JOB|15|11|numquid grande est ut consoletur te Deus sed verba tua prava hoc prohibent
JOB|15|12|quid te elevat cor tuum et quasi magna cogitans adtonitos habes oculos
JOB|15|13|quid tumet contra Deum spiritus tuus ut proferas de ore huiuscemodi sermones
JOB|15|14|quid est homo ut inmaculatus sit et ut iustus appareat natus de muliere
JOB|15|15|ecce inter sanctos eius nemo inmutabilis et caeli non sunt mundi in conspectu eius
JOB|15|16|quanto magis abominabilis et inutilis homo qui bibit quasi aquas iniquitatem
JOB|15|17|ostendam tibi audi me quod vidi narrabo tibi
JOB|15|18|sapientes confitentur et non abscondunt patres suos
JOB|15|19|quibus solis data est terra et non transibit alienus per eos
JOB|15|20|cunctis diebus suis impius superbit et numerus annorum incertus est tyrannidis eius
JOB|15|21|sonitus terroris semper in auribus illius et cum pax sit ille insidias suspicatur
JOB|15|22|non credit quod reverti possit de tenebris circumspectans undique gladium
JOB|15|23|cum se moverit ad quaerendum panem novit quod paratus sit in manu eius tenebrarum dies
JOB|15|24|terrebit eum tribulatio et angustia vallabit eum sicut regem qui praeparatur ad proelium
JOB|15|25|tetendit enim adversus Deum manum suam et contra Omnipotentem roboratus est
JOB|15|26|cucurrit adversus eum erecto collo et pingui cervice armatus est
JOB|15|27|operuit faciem eius crassitudo et de lateribus eius arvina dependet
JOB|15|28|habitavit in civitatibus desolatis et in domibus desertis quae in tumulos sunt redactae
JOB|15|29|non ditabitur nec perseverabit substantia eius nec mittet in terra radicem suam
JOB|15|30|non recedet de tenebris ramos eius arefaciet flamma et auferetur spiritu oris sui
JOB|15|31|non credat frustra errore deceptus quod aliquo pretio redimendus sit
JOB|15|32|antequam dies eius impleantur peribit et manus eius arescet
JOB|15|33|laedetur quasi vinea in primo flore botrus eius et quasi oliva proiciens florem suum
JOB|15|34|congregatio enim hypocritae sterilis et ignis devorabit tabernacula eorum qui munera libenter accipiunt
JOB|15|35|concepit dolorem et peperit iniquitatem et uterus eius praeparat dolos
JOB|16|1|respondens autem Iob dixit
JOB|16|2|audivi frequenter talia consolatores onerosi omnes vos estis
JOB|16|3|numquid habebunt finem verba ventosa aut aliquid tibi molestum est si loquaris
JOB|16|4|poteram et ego similia vestri loqui atque utinam esset anima vestra pro anima mea
JOB|16|5|consolarer et ego vos sermonibus et moverem caput meum super vos
JOB|16|6|roborarem vos ore meo et moverem labia quasi parcens vobis
JOB|16|7|sed quid agam si locutus fuero non quiescet dolor meus et si tacuero non recedet a me
JOB|16|8|nunc autem oppressit me dolor meus et in nihili redacti sunt omnes artus mei
JOB|16|9|rugae meae testimonium dicunt contra me et suscitatur falsiloquus adversus faciem meam contradicens mihi
JOB|16|10|collegit furorem suum in me et comminans mihi infremuit contra me dentibus suis hostis meus terribilibus oculis me intuitus est
JOB|16|11|aperuerunt super me ora sua exprobrantes percusserunt maxillam meam satiati sunt poenis meis
JOB|16|12|conclusit me Deus apud iniquum et manibus impiorum me tradidit
JOB|16|13|ego ille quondam opulentus repente contritus sum tenuit cervicem meam confregit me et posuit sibi quasi in signum
JOB|16|14|circumdedit me lanceis suis convulneravit lumbos meos non pepercit et effudit in terra viscera mea
JOB|16|15|concidit me vulnere super vulnus inruit in me quasi gigans
JOB|16|16|saccum consui super cutem meam et operui cinere cornu meum
JOB|16|17|facies mea intumuit a fletu et palpebrae meae caligaverunt
JOB|16|18|haec passus sum absque iniquitate manus meae cum haberem mundas ad Deum preces
JOB|16|19|terra ne operias sanguinem meum neque inveniat locum in te latendi clamor meus
JOB|16|20|ecce enim in caelo testis meus et conscius meus in excelsis
JOB|16|21|verbosi mei amici mei ad Deum stillat oculus meus
JOB|16|22|atque utinam sic iudicaretur vir cum Deo quomodo iudicatur filius hominis cum collega suo
JOB|16|23|ecce enim breves anni transeunt et semitam per quam non revertar ambulo
JOB|17|1|spiritus meus adtenuabitur dies mei breviabuntur et solum mihi superest sepulchrum
JOB|17|2|non peccavi et in amaritudinibus moratur oculus meus
JOB|17|3|libera me et pone iuxta te et cuiusvis manus pugnet contra me
JOB|17|4|cor eorum longe fecisti a disciplina et propterea non exaltabuntur
JOB|17|5|praedam pollicetur sociis et oculi filiorum eius deficient
JOB|17|6|posuit me quasi in proverbium vulgi et exemplum sum coram eis
JOB|17|7|caligavit ab indignatione oculus meus et membra mea quasi in nihili redacta sunt
JOB|17|8|stupebunt iusti super hoc et innocens contra hypocritam suscitabitur
JOB|17|9|et tenebit iustus viam suam et mundis manibus addet fortitudinem
JOB|17|10|igitur vos omnes convertimini et venite et non inveniam in vobis ullum sapientem
JOB|17|11|dies mei transierunt cogitationes meae dissipatae sunt torquentes cor meum
JOB|17|12|noctem verterunt in diem et rursum post tenebras spero lucem
JOB|17|13|si sustinuero infernus domus mea est in tenebris stravi lectulum meum
JOB|17|14|putredini dixi pater meus es mater mea et soror mea vermibus
JOB|17|15|ubi est ergo nunc praestolatio mea et patientiam meam quis considerat
JOB|17|16|in profundissimum infernum descendent omnia mea putasne saltim ibi erit requies mihi
JOB|18|1|respondens autem Baldad Suites dixit
JOB|18|2|usque ad quem finem verba iactabitis intellegite prius et sic loquamur
JOB|18|3|quare reputati sumus ut iumenta et sorduimus coram vobis
JOB|18|4|qui perdis animam tuam in furore tuo numquid propter te derelinquetur terra et transferentur rupes de loco suo
JOB|18|5|nonne lux impii extinguetur nec splendebit flamma ignis eius
JOB|18|6|lux obtenebrescet in tabernaculo illius et lucerna quae super eum est extinguetur
JOB|18|7|artabuntur gressus virtutis eius et praecipitabit eum consilium suum
JOB|18|8|inmisit enim in rete pedes suos et in maculis eius ambulat
JOB|18|9|tenebitur planta illius laqueo et exardescet contra eum sitis
JOB|18|10|abscondita est in terra pedica eius et decipula illius super semitam
JOB|18|11|undique terrebunt eum formidines et involvent pedes eius
JOB|18|12|adtenuetur fame robur eius et inedia invadat costas illius
JOB|18|13|devoret pulchritudinem cutis eius consumat brachia illius primogenita mors
JOB|18|14|avellatur de tabernaculo suo fiducia eius et calcet super eum quasi rex interitus
JOB|18|15|habitent in tabernaculo illius socii eius qui non est aspergatur in tabernaculo eius sulphur
JOB|18|16|deorsum radices eius siccentur sursum autem adteratur messis eius
JOB|18|17|memoria illius pereat de terra et non celebretur nomen eius in plateis
JOB|18|18|expellet eum de luce in tenebras et de orbe transferet eum
JOB|18|19|non erit semen eius neque progenies in populo suo nec ullae reliquiae in regionibus eius
JOB|18|20|in die eius stupebunt novissimi et primos invadet horror
JOB|18|21|haec sunt ergo tabernacula iniqui et iste locus eius qui ignorat Deum
JOB|19|1|respondens autem Iob dixit
JOB|19|2|usquequo adfligitis animam meam et adteritis me sermonibus
JOB|19|3|en decies confunditis me et non erubescitis opprimentes me
JOB|19|4|nempe et si ignoravi mecum erit ignorantia mea
JOB|19|5|at vos contra me erigimini et arguitis me obprobriis meis
JOB|19|6|saltim nunc intellegite quia Deus non aequo iudicio adflixerit me et flagellis suis me cinxerit
JOB|19|7|ecce clamabo vim patiens et nemo audiet vociferabor et non est qui iudicet
JOB|19|8|semitam meam circumsepsit et transire non possum et in calle meo tenebras posuit
JOB|19|9|spoliavit me gloria mea et abstulit coronam de capite meo
JOB|19|10|destruxit me undique et pereo et quasi evulsae arbori abstulit spem meam
JOB|19|11|iratus est contra me furor eius et sic me habuit quasi hostem suum
JOB|19|12|simul venerunt latrones eius et fecerunt sibi viam per me et obsederunt in gyro tabernaculum meum
JOB|19|13|fratres meos longe fecit a me et noti mei quasi alieni recesserunt a me
JOB|19|14|dereliquerunt me propinqui mei et qui me noverant obliti sunt mei
JOB|19|15|inquilini domus meae et ancillae meae sicut alienum habuerunt me et quasi peregrinus fui in oculis eorum
JOB|19|16|servum meum vocavi et non respondit ore proprio deprecabar illum
JOB|19|17|halitum meum exhorruit uxor mea et orabam filios uteri mei
JOB|19|18|stulti quoque despiciebant me et cum ab eis recessissem detrahebant mihi
JOB|19|19|abominati sunt me quondam consiliarii mei et quem maxime diligebam aversatus est me
JOB|19|20|pelli meae consumptis carnibus adhesit os meum et derelicta sunt tantummodo labia circa dentes meos
JOB|19|21|miseremini mei miseremini mei saltim vos amici mei quia manus Domini tetigit me
JOB|19|22|quare persequimini me sicut Deus et carnibus meis saturamini
JOB|19|23|quis mihi tribuat ut scribantur sermones mei quis mihi det ut exarentur in libro
JOB|19|24|stilo ferreo et plumbi lammina vel certe sculpantur in silice
JOB|19|25|scio enim quod redemptor meus vivat et in novissimo de terra surrecturus sim
JOB|19|26|et rursum circumdabor pelle mea et in carne mea videbo Deum
JOB|19|27|quem visurus sum ego ipse et oculi mei conspecturi sunt et non alius reposita est haec spes mea in sinu meo
JOB|19|28|quare ergo nunc dicitis persequamur eum et radicem verbi inveniamus contra eum
JOB|19|29|fugite ergo a facie gladii quoniam ultor iniquitatum gladius est et scitote esse iudicium
JOB|20|1|respondens autem Sophar Naamathites dixit
JOB|20|2|idcirco cogitationes meae variae succedunt sibi et mens in diversa rapitur
JOB|20|3|doctrinam qua me arguis audiam et spiritus intellegentiae meae respondebit mihi
JOB|20|4|hoc scio a principio ex quo positus est homo super terram
JOB|20|5|quod laus impiorum brevis sit et gaudium hypocritae ad instar puncti
JOB|20|6|si ascenderit usque ad caelum superbia eius et caput eius nubes tetigerit
JOB|20|7|quasi sterquilinium in fine perdetur et qui eum viderant dicent ubi est
JOB|20|8|velut somnium avolans non invenietur transiet sicut visio nocturna
JOB|20|9|oculus qui eum viderat non videbit neque ultra intuebitur eum locus suus
JOB|20|10|filii eius adterentur egestate et manus illius reddent ei dolorem suum
JOB|20|11|ossa eius implebuntur vitiis adulescentiae eius et cum eo in pulverem dormient
JOB|20|12|cum enim dulce fuerit in ore eius malum abscondet illud sub lingua sua
JOB|20|13|parcet illi et non derelinquet illud et celabit in gutture suo
JOB|20|14|panis eius in utero illius vertetur in fel aspidum intrinsecus
JOB|20|15|divitias quas devoravit evomet et de ventre illius extrahet eas Deus
JOB|20|16|caput aspidum suget occidet eum lingua viperae
JOB|20|17|non videat rivulos fluminis torrentes mellis et butyri
JOB|20|18|luet quae fecit omnia nec tamen consumetur iuxta multitudinem adinventionum suarum sic et sustinebit
JOB|20|19|quoniam confringens nudavit pauperes domum rapuit et non aedificavit eam
JOB|20|20|nec est satiatus venter eius et cum habuerit quae cupierat possidere non poterit
JOB|20|21|non remansit de cibo eius et propterea nihil permanebit de bonis eius
JOB|20|22|cum satiatus fuerit artabitur aestuabit et omnis dolor inruet in eum
JOB|20|23|utinam impleatur venter eius ut emittat in eum iram furoris sui et pluat super illum bellum suum
JOB|20|24|fugiet arma ferrea et inruet in arcum aereum
JOB|20|25|eductus et egrediens de vagina sua et fulgurans in amaritudine sua vadent et venient super eum horribiles
JOB|20|26|omnes tenebrae absconditae sunt in occultis eius devorabit eum ignis qui non succenditur adfligetur relictus in tabernaculo suo
JOB|20|27|revelabunt caeli iniquitatem eius et terra consurget adversus eum
JOB|20|28|apertum erit germen domus illius detrahetur in die furoris Dei
JOB|20|29|haec est pars hominis impii a Deo et hereditas verborum eius a Domino
JOB|21|1|respondens autem Iob dixit
JOB|21|2|audite quaeso sermones meos et agetis paenitentiam
JOB|21|3|sustinete me ut et ego loquar et post mea si videbitur verba ridete
JOB|21|4|numquid contra hominem disputatio mea est ut merito non debeam contristari
JOB|21|5|adtendite me et obstupescite et superponite digitum ori vestro
JOB|21|6|et ego quando recordatus fuero pertimesco et concutit carnem meam tremor
JOB|21|7|quare ergo impii vivunt sublevati sunt confortatique divitiis
JOB|21|8|semen eorum permanet coram eis propinquorum turba et nepotum in conspectu eorum
JOB|21|9|domus eorum securae sunt et pacatae et non est virga Dei super illos
JOB|21|10|bos eorum concepit et non abortit vacca peperit et non est privata fetu suo
JOB|21|11|egrediuntur quasi greges parvuli eorum et infantes eorum exultant lusibus
JOB|21|12|tenent tympanum et citharam et gaudent ad sonitum organi
JOB|21|13|ducunt in bonis dies suos et in puncto ad inferna descendunt
JOB|21|14|qui dixerunt Deo recede a nobis et scientiam viarum tuarum nolumus
JOB|21|15|quid est Omnipotens ut serviamus ei et quid nobis prodest si oraverimus illum
JOB|21|16|verumtamen quia non sunt in manu eorum bona sua consilium impiorum longe sit a me
JOB|21|17|quotiens lucerna impiorum extinguetur et superveniet eis inundatio et dolores dividet furoris sui
JOB|21|18|erunt sicut paleae ante faciem venti et sicut favilla quam turbo dispergit
JOB|21|19|Deus servabit filiis illius dolorem patris et cum reddiderit tunc sciet
JOB|21|20|videbunt oculi eius interfectionem suam et de furore Omnipotentis bibet
JOB|21|21|quid enim ad eum pertinet de domo sua post se et si numerus mensuum eius dimidietur
JOB|21|22|numquid Deum quispiam docebit scientiam qui excelsos iudicat
JOB|21|23|iste moritur robustus et sanus dives et felix
JOB|21|24|viscera eius plena sunt adipe et medullis ossa illius inrigantur
JOB|21|25|alius vero moritur in amaritudine animae absque ullis opibus
JOB|21|26|et tamen simul in pulverem dormient et vermes operient eos
JOB|21|27|certe novi cogitationes vestras et sententias contra me iniquas
JOB|21|28|dicitis enim ubi est domus principis et ubi tabernacula impiorum
JOB|21|29|interrogate quemlibet de viatoribus et haec eadem eum intellegere cognoscetis
JOB|21|30|quia in diem perditionis servabitur malus et ad diem furoris ducitur
JOB|21|31|quis arguet coram eo viam eius et quae fecit quis reddet illi
JOB|21|32|ipse ad sepulchra ducetur et in congerie mortuorum vigilabit
JOB|21|33|dulcis fuit glareis Cocyti et post se omnem hominem trahet et ante se innumerabiles
JOB|21|34|quomodo igitur consolamini me frustra cum responsio vestra repugnare ostensa sit veritati
JOB|22|1|respondens autem Eliphaz Themanites dixit
JOB|22|2|numquid Deo conparari potest homo etiam cum perfectae fuerit scientiae
JOB|22|3|quid prodest Deo si iustus fueris aut quid ei confers si inmaculata fuerit via tua
JOB|22|4|numquid timens arguet te et veniet tecum in iudicium
JOB|22|5|et non propter malitiam tuam plurimam et infinitas iniquitates tuas
JOB|22|6|abstulisti enim pignus fratrum tuorum sine causa et nudos spoliasti vestibus
JOB|22|7|aquam lasso non dedisti et esurienti subtraxisti panem
JOB|22|8|in fortitudine brachii tui possidebas terram et potentissimus obtinebas eam
JOB|22|9|viduas dimisisti vacuas et lacertos pupillorum comminuisti
JOB|22|10|propterea circumdatus es laqueis et conturbat te formido subita
JOB|22|11|et putabas te tenebras non visurum et impetu aquarum inundantium non oppressurum
JOB|22|12|an cogitas quod Deus excelsior caelo et super stellarum vertices sublimetur
JOB|22|13|et dicis quid enim novit Deus et quasi per caliginem iudicat
JOB|22|14|nubes latibulum eius nec nostra considerat et circa cardines caeli perambulat
JOB|22|15|numquid semitam saeculorum custodire cupis quam calcaverunt viri iniqui
JOB|22|16|qui sublati sunt ante tempus suum et fluvius subvertit fundamentum eorum
JOB|22|17|qui dicebant Deo recede a nobis et quasi nihil possit facere Omnipotens aestimabant eum
JOB|22|18|cum ille implesset domos eorum bonis quorum sententia procul sit a me
JOB|22|19|videbunt iusti et laetabuntur et innocens subsannabit eos
JOB|22|20|nonne succisa est erectio eorum et reliquias eorum devoravit ignis
JOB|22|21|adquiesce igitur ei et habeto pacem et per haec habebis fructus optimos
JOB|22|22|suscipe ex ore illius legem et pone sermones eius in corde tuo
JOB|22|23|si reversus fueris ad Omnipotentem aedificaberis et longe facies iniquitatem a tabernaculo tuo
JOB|22|24|dabit pro terra silicem et pro silice torrentes aureos
JOB|22|25|eritque Omnipotens contra hostes tuos et argentum coacervabitur tibi
JOB|22|26|tunc super Omnipotentem deliciis afflues et elevabis ad Deum faciem tuam
JOB|22|27|rogabis eum et exaudiet te et vota tua reddes
JOB|22|28|decernes rem et veniet tibi et in viis tuis splendebit lumen
JOB|22|29|qui enim humiliatus fuerit erit in gloria et qui inclinaverit oculos suos ipse salvabitur
JOB|22|30|salvabitur innocens salvabitur autem munditia manuum suarum
JOB|23|1|respondens autem Iob dixit
JOB|23|2|nunc quoque in amaritudine est sermo meus et manus plagae meae adgravata est super gemitum meum
JOB|23|3|quis mihi tribuat ut cognoscam et inveniam illum et veniam usque ad solium eius
JOB|23|4|ponam coram eo iudicium et os meum replebo increpationibus
JOB|23|5|ut sciam verba quae mihi respondeat et intellegam quid loquatur mihi
JOB|23|6|nolo multa fortitudine contendat mecum nec magnitudinis suae mole me premat
JOB|23|7|proponat aequitatem contra me et perveniat ad victoriam iudicium meum
JOB|23|8|si ad orientem iero non apparet si ad occidentem non intellegam eum
JOB|23|9|si ad sinistram quid agat non adprehendam eum si me vertam ad dextram non videbo illum
JOB|23|10|ipse vero scit viam meam et probavit me quasi aurum quod per ignem transit
JOB|23|11|vestigia eius secutus est pes meus viam eius custodivi et non declinavi ex ea
JOB|23|12|a mandatis labiorum eius non recessi et in sinu meo abscondi verba oris eius
JOB|23|13|ipse enim solus est et nemo avertere potest cogitationem eius et anima eius quodcumque voluerit hoc facit
JOB|23|14|cum expleverit in me voluntatem suam et alia multa similia praesto sunt ei
JOB|23|15|et idcirco a facie eius turbatus sum et considerans eum timore sollicitor
JOB|23|16|Deus mollivit cor meum et Omnipotens conturbavit me
JOB|23|17|non enim perii propter inminentes tenebras nec faciem meam operuit caligo
JOB|24|1|ab Omnipotente non sunt abscondita tempora qui autem noverunt eum ignorant dies illius
JOB|24|2|alii terminos transtulerunt diripuerunt greges et paverunt eos
JOB|24|3|asinum pupillorum abigerunt et abstulerunt pro pignore bovem viduae
JOB|24|4|subverterunt pauperum viam et oppresserunt pariter mansuetos terrae
JOB|24|5|alii quasi onagri in deserto egrediuntur ad opus suum vigilantesque ad praedam praeparant panem liberis
JOB|24|6|agrum non suum demetunt et vineam eius quem vi oppresserunt vindemiant
JOB|24|7|nudos dimittunt homines indumenta tollentes quibus non est operimentum in frigore
JOB|24|8|quos imbres montium rigant et non habentes velamen amplexantur lapides
JOB|24|9|vim fecerunt depraedantes pupillos et vulgum pauperem spoliaverunt
JOB|24|10|nudis et incedentibus absque vestitu et esurientibus tulerunt spicas
JOB|24|11|inter acervos eorum meridiati sunt qui calcatis torcularibus sitiunt
JOB|24|12|de civitatibus fecerunt viros gemere et anima vulneratorum clamavit et Deus inultum abire non patitur
JOB|24|13|ipsi fuerunt rebelles luminis nescierunt vias eius nec reversi sunt per semitas illius
JOB|24|14|mane primo consurgit homicida interficit egenum et pauperem per noctem vero erit quasi fur
JOB|24|15|oculus adulteri observat caliginem dicens non me videbit oculus et operiet vultum suum
JOB|24|16|perfodit in tenebris domos sicut in die condixerant sibi et ignoraverunt lucem
JOB|24|17|si subito apparuerit aurora arbitrantur umbram mortis et sic in tenebris quasi in luce ambulant
JOB|24|18|levis est super faciem aquae maledicta sit pars eius in terra nec ambulet per viam vinearum
JOB|24|19|ad nimium calorem transeat ab aquis nivium et usque ad inferos peccatum illius
JOB|24|20|obliviscatur eius misericordia dulcedo illius vermes non sit in recordatione sed conteratur quasi lignum infructuosum
JOB|24|21|pavit enim sterilem et quae non parit et viduae bene non fecit
JOB|24|22|detraxit fortes in fortitudine sua et cum steterit non credet vitae suae
JOB|24|23|dedit ei Deus locum paenitentiae et ille abutitur eo in superbiam oculi autem eius sunt in viis illius
JOB|24|24|elevati sunt ad modicum et non subsistent et humiliabuntur sicut omnia et auferentur et sicut summitates spicarum conterentur
JOB|24|25|quod si non est ita quis me potest arguere esse mentitum et ponere ante Deum verba mea
JOB|25|1|respondens autem Baldad Suites dixit
JOB|25|2|potestas et terror apud eum est qui facit concordiam in sublimibus suis
JOB|25|3|numquid est numerus militum eius et super quem non surget lumen illius
JOB|25|4|numquid iustificari potest homo conparatus Deo aut apparere mundus natus de muliere
JOB|25|5|ecce etiam luna non splendet et stellae non sunt mundae in conspectu eius
JOB|25|6|quanto magis homo putredo et filius hominis vermis
JOB|26|1|respondens autem Iob dixit
JOB|26|2|cuius adiutor es numquid inbecilli et sustentas brachium eius qui non est fortis
JOB|26|3|cui dedisti consilium forsitan illi qui non habet sapientiam et prudentiam tuam ostendisti plurimam
JOB|26|4|quem docere voluisti nonne eum qui fecit spiramen tuum
JOB|26|5|ecce gigantes gemunt sub aquis et qui habitant cum eis
JOB|26|6|nudus est inferus coram illo et nullum est operimentum perditioni
JOB|26|7|qui extendit aquilonem super vacuum et adpendit terram super nihili
JOB|26|8|qui ligat aquas in nubibus suis ut non erumpant pariter deorsum
JOB|26|9|qui tenet vultum solii sui et expandit super illud nebulam suam
JOB|26|10|terminum circumdedit aquis usque dum finiantur lux et tenebrae
JOB|26|11|columnae caeli contremescunt et pavent ad nutum eius
JOB|26|12|in fortitudine illius repente maria congregata sunt et prudentia eius percussit superbum
JOB|26|13|spiritus eius ornavit caelos et obsetricante manu eius eductus est coluber tortuosus
JOB|26|14|ecce haec ex parte dicta sunt viarum eius et cum vix parvam stillam sermonis eius audierimus quis poterit tonitruum magnitudinis illius intueri
JOB|27|1|addidit quoque Iob adsumens parabolam suam et dixit
JOB|27|2|vivit Deus qui abstulit iudicium meum et Omnipotens qui ad amaritudinem adduxit animam meam
JOB|27|3|quia donec superest halitus in me et spiritus Dei in naribus meis
JOB|27|4|non loquentur labia mea iniquitatem nec lingua mea meditabitur mendacium
JOB|27|5|absit a me ut iustos vos esse iudicem donec deficiam non recedam ab innocentia mea
JOB|27|6|iustificationem meam quam coepi tenere non deseram nec enim reprehendit me cor meum in omni vita mea
JOB|27|7|sit ut impius inimicus meus et adversarius meus quasi iniquus
JOB|27|8|quae enim spes est hypocritae si avare rapiat et non liberet Deus animam eius
JOB|27|9|numquid clamorem eius Deus audiet cum venerit super illum angustia
JOB|27|10|aut poterit in Omnipotente delectari et invocare Deum in omni tempore
JOB|27|11|docebo vos per manum Dei quae Omnipotens habeat nec abscondam
JOB|27|12|ecce vos omnes nostis et quid sine causa vana loquimini
JOB|27|13|haec est pars hominis impii apud Deum et hereditas violentorum quam ab Omnipotente suscipient
JOB|27|14|si multiplicati fuerint filii eius in gladio erunt et nepotes eius non saturabuntur pane
JOB|27|15|qui reliqui fuerint ex eo sepelientur in interitu et viduae illius non plorabunt
JOB|27|16|si conportaverit quasi terram argentum et sicut lutum praeparaverit vestimenta
JOB|27|17|praeparabit quidem sed iustus vestietur illis et argentum innocens dividet
JOB|27|18|aedificavit sicut tinea domum suam et sicut custos fecit umbraculum
JOB|27|19|dives cum dormierit nihil secum auferet aperit oculos suos et nihil inveniet
JOB|27|20|adprehendit eum quasi aqua inopia nocte opprimet eum tempestas
JOB|27|21|tollet eum ventus urens et auferet et velut turbo rapiet eum de loco suo
JOB|27|22|et mittet super eum et non parcet de manu eius fugiens fugiet
JOB|27|23|stringet super eum manus suas et sibilabit super illum intuens locum eius
JOB|28|1|habet argentum venarum suarum principia et auro locus est in quo conflatur
JOB|28|2|ferrum de terra tollitur et lapis solutus calore in aes vertitur
JOB|28|3|tempus posuit tenebris et universorum finem ipse considerat lapidem quoque caliginis et umbram mortis
JOB|28|4|dividit torrens a populo peregrinante eos quos oblitus est pes egentis hominum et invios
JOB|28|5|terra de qua oriebatur panis in loco suo igne subversa est
JOB|28|6|locus sapphyri lapides eius et glebae illius aurum
JOB|28|7|semitam ignoravit avis nec intuitus est oculus vulturis
JOB|28|8|non calcaverunt eam filii institorum nec pertransivit per eam leaena
JOB|28|9|ad silicem extendit manum suam subvertit a radicibus montes
JOB|28|10|in petris rivos excidit et omne pretiosum vidit oculus eius
JOB|28|11|profunda quoque fluviorum scrutatus est et abscondita produxit in lucem
JOB|28|12|sapientia vero ubi invenitur et quis est locus intellegentiae
JOB|28|13|nescit homo pretium eius nec invenitur in terra suaviter viventium
JOB|28|14|abyssus dicit non est in me et mare loquitur non est mecum
JOB|28|15|non dabitur aurum obrizum pro ea nec adpendetur argentum in commutatione eius
JOB|28|16|non conferetur tinctis Indiae coloribus nec lapidi sardonico pretiosissimo vel sapphyro
JOB|28|17|non adaequabitur ei aurum vel vitrum nec commutabuntur pro ea vasa auri
JOB|28|18|excelsa et eminentia non memorabuntur conparatione eius trahitur autem sapientia de occultis
JOB|28|19|non adaequabitur ei topazium de Aethiopia nec tincturae mundissimae conponetur
JOB|28|20|unde ergo sapientia veniet et quis est locus intellegentiae
JOB|28|21|abscondita est ab oculis omnium viventium volucres quoque caeli latet
JOB|28|22|perditio et mors dixerunt auribus nostris audivimus famam eius
JOB|28|23|Deus intellegit viam eius et ipse novit locum illius
JOB|28|24|ipse enim fines mundi intuetur et omnia quae sub caelo sunt respicit
JOB|28|25|qui fecit ventis pondus et aquas adpendit mensura
JOB|28|26|quando ponebat pluviis legem et viam procellis sonantibus
JOB|28|27|tunc vidit illam et enarravit et praeparavit et investigavit
JOB|28|28|et dixit homini ecce timor Domini ipsa est sapientia et recedere a malo intellegentia
JOB|29|1|addidit quoque Iob adsumens parabolam suam et dixit
JOB|29|2|quis mihi tribuat ut sim iuxta menses pristinos secundum dies quibus Deus custodiebat me
JOB|29|3|quando splendebat lucerna eius super caput meum et ad lumen eius ambulabam in tenebris
JOB|29|4|sicut fui in diebus adulescentiae meae quando secreto Deus erat in tabernaculo meo
JOB|29|5|quando erat Omnipotens mecum et in circuitu meo pueri mei
JOB|29|6|quando lavabam pedes meos butyro et petra fundebat mihi rivos olei
JOB|29|7|quando procedebam ad portam civitatis et in platea parabant cathedram mihi
JOB|29|8|videbant me iuvenes et abscondebantur et senes adsurgentes stabant
JOB|29|9|principes cessabant loqui et digitum superponebant ori suo
JOB|29|10|vocem suam cohibebant duces et lingua eorum gutturi suo adherebat
JOB|29|11|auris audiens beatificabat me et oculus videns testimonium reddebat mihi
JOB|29|12|quod liberassem pauperem vociferantem et pupillum cui non esset adiutor
JOB|29|13|benedictio perituri super me veniebat et cor viduae consolatus sum
JOB|29|14|iustitia indutus sum et vestivit me sicut vestimento et diademate iudicio meo
JOB|29|15|oculus fui caeco et pes claudo
JOB|29|16|pater eram pauperum et causam quam nesciebam diligentissime investigabam
JOB|29|17|conterebam molas iniqui et de dentibus illius auferebam praedam
JOB|29|18|dicebamque in nidulo meo moriar et sicut palma multiplicabo dies
JOB|29|19|radix mea aperta est secus aquas et ros morabitur in messione mea
JOB|29|20|gloria mea semper innovabitur et arcus meus in manu mea instaurabitur
JOB|29|21|qui me audiebant expectabant sententiam et intenti tacebant ad consilium meum
JOB|29|22|verbis meis addere nihil audebant et super illos stillabat eloquium meum
JOB|29|23|expectabant me sicut pluviam et os suum aperiebant quasi ad imbrem serotinum
JOB|29|24|si quando ridebam ad eos non credebant et lux vultus mei non cadebat in terram
JOB|29|25|si voluissem ire ad eos sedebam primus cumque sederem quasi rex circumstante exercitu eram tamen maerentium consolator
JOB|30|1|nunc autem derident me iuniores tempore quorum non dignabar patres ponere cum canibus gregis mei
JOB|30|2|quorum virtus manuum erat mihi pro nihilo et vita ipsa putabantur indigni
JOB|30|3|egestate et fame steriles qui rodebant in solitudine squalentes calamitate et miseria
JOB|30|4|et mandebant herbas et arborum cortices et radix iuniperorum erat cibus eorum
JOB|30|5|qui de convallibus ista rapientes cum singula repperissent ad ea cum clamore currebant
JOB|30|6|in desertis habitabant torrentium et in cavernis terrae vel super glaream
JOB|30|7|qui inter huiuscemodi laetabantur et esse sub sentibus delicias conputabant
JOB|30|8|filii stultorum et ignobilium et in terra penitus non parentes
JOB|30|9|nunc in eorum canticum versus sum et factus sum eis proverbium
JOB|30|10|abominantur me et longe fugiunt a me et faciem meam conspuere non verentur
JOB|30|11|faretram enim suam aperuit et adflixit me et frenum posuit in os meum
JOB|30|12|ad dexteram orientis calamitatis meae ilico surrexerunt pedes meos subverterunt et oppresserunt quasi fluctibus semitis suis
JOB|30|13|dissipaverunt itinera mea insidiati sunt mihi et praevaluerunt et non fuit qui ferret auxilium
JOB|30|14|quasi rupto muro et aperta ianua inruerunt super me et ad meas miserias devoluti sunt
JOB|30|15|redactus sum in nihili abstulisti quasi ventus desiderium meum et velut nubes pertransiit salus mea
JOB|30|16|nunc autem in memet ipso marcescit anima mea et possident me dies adflictionis
JOB|30|17|nocte os meum perforatur doloribus et qui me comedunt non dormiunt
JOB|30|18|in multitudine eorum consumitur vestimentum meum et quasi capitio tunicae sic cinxerunt me
JOB|30|19|conparatus sum luto et adsimilatus favillae et cineri
JOB|30|20|clamo ad te et non exaudis me sto et non respicis me
JOB|30|21|mutatus es mihi in crudelem et in duritia manus tuae adversaris mihi
JOB|30|22|elevasti me et quasi super ventum ponens elisisti me valide
JOB|30|23|scio quia morti tradas me ubi constituta domus est omni viventi
JOB|30|24|verumtamen non ad consumptionem eorum emittis manum tuam et si corruerint ipse salvabis
JOB|30|25|flebam quondam super eum qui adflictus erat et conpatiebatur anima mea pauperi
JOB|30|26|expectabam bona et venerunt mihi mala praestolabar lucem et eruperunt tenebrae
JOB|30|27|interiora mea efferbuerunt absque ulla requie praevenerunt me dies adflictionis
JOB|30|28|maerens incedebam sine furore consurgens in turba clamavi
JOB|30|29|frater fui draconum et socius strutionum
JOB|30|30|cutis mea denigrata est super me et ossa mea aruerunt prae caumate
JOB|30|31|versa est in luctum cithara mea et organum meum in vocem flentium
JOB|31|1|pepigi foedus cum oculis meis ut ne cogitarem quidem de virgine
JOB|31|2|quam enim partem haberet Deus in me desuper et hereditatem Omnipotens de excelsis
JOB|31|3|numquid non perditio est iniquo et alienatio operantibus iniustitiam
JOB|31|4|nonne ipse considerat vias meas et cunctos gressus meos dinumerat
JOB|31|5|si ambulavi in vanitate et festinavit in dolo pes meus
JOB|31|6|adpendat me in statera iusta et sciat Deus simplicitatem meam
JOB|31|7|si declinavit gressus meus de via et si secutum est oculos meos cor meum et in manibus meis adhesit macula
JOB|31|8|seram et alius comedat et progenies mea eradicetur
JOB|31|9|si deceptum est cor meum super mulierem et si ad ostium amici mei insidiatus sum
JOB|31|10|scortum sit alteri uxor mea et super illam incurventur alii
JOB|31|11|hoc enim nefas est et iniquitas maxima
JOB|31|12|ignis est usque ad perditionem devorans et omnia eradicans genimina
JOB|31|13|si contempsi subire iudicium cum servo meo et ancillae meae cum disceptarent adversum me
JOB|31|14|quid enim faciam cum surrexerit ad iudicandum Deus et cum quaesierit quid respondebo illi
JOB|31|15|numquid non in utero fecit me qui et illum operatus est et formavit in vulva unus
JOB|31|16|si negavi quod volebant pauperibus et oculos viduae expectare feci
JOB|31|17|si comedi buccellam meam solus et non comedit pupillus ex ea
JOB|31|18|quia ab infantia mea crevit mecum miseratio et de utero matris meae egressa est mecum
JOB|31|19|si despexi pereuntem eo quod non habuerit indumentum et absque operimento pauperem
JOB|31|20|si non benedixerunt mihi latera eius et de velleribus ovium mearum calefactus est
JOB|31|21|si levavi super pupillum manum meam etiam cum viderem me in porta superiorem
JOB|31|22|umerus meus a iunctura sua cadat et brachium meum cum suis ossibus confringatur
JOB|31|23|semper enim quasi tumentes super me fluctus timui Deum et pondus eius ferre non potui
JOB|31|24|si putavi aurum robur meum et obrizae dixi fiducia mea
JOB|31|25|si laetatus sum super multis divitiis meis et quia plurima repperit manus mea
JOB|31|26|si vidi solem cum fulgeret et lunam incedentem clare
JOB|31|27|et lactatum est in abscondito cor meum et osculatus sum manum meam ore meo
JOB|31|28|quae est iniquitas maxima et negatio contra Deum altissimum
JOB|31|29|si gavisus sum ad ruinam eius qui me oderat et exultavi quod invenisset eum malum
JOB|31|30|non enim dedi ad peccandum guttur meum ut expeterem maledicens animam eius
JOB|31|31|si non dixerunt viri tabernaculi mei quis det de carnibus eius ut saturemur
JOB|31|32|foris non mansit peregrinus ostium meum viatori patuit
JOB|31|33|si abscondi quasi homo peccatum meum et celavi in sinu meo iniquitatem meam
JOB|31|34|si expavi ad multitudinem nimiam et despectio propinquorum terruit me et non magis tacui nec egressus sum ostium
JOB|31|35|quis mihi tribuat auditorem ut desiderium meum Omnipotens audiat et librum scribat ipse qui iudicat
JOB|31|36|ut in umero meo portem illum et circumdem illum quasi coronam mihi
JOB|31|37|per singulos gradus meos pronuntiabo illum et quasi principi offeram eum
JOB|31|38|si adversum me terra mea clamat et cum ipsa sulci eius deflent
JOB|31|39|si fructus eius comedi absque pecunia et animam agricolarum eius adflixi
JOB|31|40|pro frumento oriatur mihi tribulus et pro hordeo spina finita sunt verba Iob
JOB|32|1|omiserunt autem tres viri isti respondere Iob eo quod iustus sibi videretur
JOB|32|2|et iratus indignatusque Heliu filius Barachel Buzites de cognatione Ram iratus est autem adversus Iob eo quod iustum se esse diceret coram Deo
JOB|32|3|porro adversum amicos eius indignatus est eo quod non invenissent responsionem rationabilem sed tantummodo condemnassent Iob
JOB|32|4|igitur Heliu expectavit Iob loquentem eo quod seniores se essent qui loquebantur
JOB|32|5|cum autem vidisset quod tres respondere non potuissent iratus est vehementer
JOB|32|6|respondensque Heliu filius Barachel Buzites dixit iunior sum tempore vos autem antiquiores idcirco dimisso capite veritus sum indicare vobis meam sententiam
JOB|32|7|sperabam enim quod aetas prolixior loqueretur et annorum multitudo doceret sapientiam
JOB|32|8|sed ut video spiritus est in hominibus et inspiratio Omnipotentis dat intellegentiam
JOB|32|9|non sunt longevi sapientes nec senes intellegunt iudicium
JOB|32|10|ideo dicam audite me ostendam vobis etiam ego meam scientiam
JOB|32|11|expectavi enim sermones vestros audivi prudentiam vestram donec disceptaremini sermonibus
JOB|32|12|et donec putabam vos aliquid dicere considerabam sed ut video non est qui arguere possit Iob et respondere ex vobis sermonibus eius
JOB|32|13|ne forte dicatis invenimus sapientiam Deus proiecit eum non homo
JOB|32|14|nihil locutus est mihi et ego non secundum vestros sermones respondebo illi
JOB|32|15|extimuerunt non responderunt ultra abstuleruntque a se eloquia
JOB|32|16|quoniam igitur expectavi et non sunt locuti steterunt nec responderunt ultra
JOB|32|17|respondebo et ego partem meam et ostendam scientiam meam
JOB|32|18|plenus sum enim sermonibus et coartat me spiritus uteri mei
JOB|32|19|en venter meus quasi mustum absque spiraculo quod lagunculas novas disrumpit
JOB|32|20|loquar et respirabo paululum aperiam labia mea et respondebo
JOB|32|21|non accipiam personam viri et Deum homini non aequabo
JOB|32|22|nescio enim quamdiu subsistam et si post modicum tollat me factor meus
JOB|33|1|audi igitur Iob eloquia mea et omnes sermones meos ausculta
JOB|33|2|ecce aperui os meum loquatur lingua mea in faucibus meis
JOB|33|3|simplici corde meo sermones mei et sententiam labia mea puram loquentur
JOB|33|4|spiritus Dei fecit me et spiraculum Omnipotentis vivificavit me
JOB|33|5|si potes responde mihi et adversus faciem meam consiste
JOB|33|6|ecce et me sicut et te fecit Deus et de eodem luto ego quoque formatus sum
JOB|33|7|verumtamen miraculum meum non te terreat et eloquentia mea non sit tibi gravis
JOB|33|8|dixisti ergo in auribus meis et vocem verborum audivi
JOB|33|9|mundus sum ego absque delicto inmaculatus et non est iniquitas in me
JOB|33|10|quia querellas in me repperit ideo arbitratus est me inimicum sibi
JOB|33|11|posuit in nervo pedes meos custodivit omnes semitas meas
JOB|33|12|hoc est ergo in quo non es iustificatus respondebo tibi quia maior sit Deus homine
JOB|33|13|adversum eum contendis quod non ad omnia verba responderit tibi
JOB|33|14|semel loquitur Deus et secundo id ipsum non repetit
JOB|33|15|per somnium in visione nocturna quando inruit sopor super homines et dormiunt in lectulo
JOB|33|16|tunc aperit aures virorum et erudiens eos instruit disciplinam
JOB|33|17|ut avertat hominem ab his quae facit et liberet eum de superbia
JOB|33|18|eruens animam eius a corruptione et vitam illius ut non transeat in gladium
JOB|33|19|increpat quoque per dolorem in lectulo et omnia ossa eius marcescere facit
JOB|33|20|abominabilis ei fit in vita sua panis et animae illius cibus ante desiderabilis
JOB|33|21|tabescet caro eius et ossa quae tecta fuerant nudabuntur
JOB|33|22|adpropinquabit corruptioni anima eius et vita illius mortiferis
JOB|33|23|si fuerit pro eo angelus loquens unum de milibus ut adnuntiet hominis aequitatem
JOB|33|24|miserebitur eius et dicet libera eum et non descendat in corruptionem inveni in quo ei propitier
JOB|33|25|consumpta est caro eius a suppliciis revertatur ad dies adulescentiae suae
JOB|33|26|deprecabitur Deum et placabilis ei erit et videbit faciem eius in iubilo et reddet homini iustitiam suam
JOB|33|27|respiciet homines et dicet peccavi et vere deliqui et ut eram dignus non recepi
JOB|33|28|liberavit animam suam ne pergeret in interitum sed vivens lucem videret
JOB|33|29|ecce haec omnia operatur Deus tribus vicibus per singulos
JOB|33|30|ut revocet animas eorum a corruptione et inluminet luce viventium
JOB|33|31|adtende Iob et audi me et tace dum ego loquar
JOB|33|32|si autem habes quod loquaris responde mihi loquere volo enim te apparere iustum
JOB|33|33|quod si non habes audi me tace et docebo te sapientiam
JOB|34|1|pronuntians itaque Heliu etiam haec locutus est
JOB|34|2|audite sapientes verba mea et eruditi auscultate me
JOB|34|3|auris enim verba probat et guttur escas gustu diiudicat
JOB|34|4|iudicium eligamus nobis et inter nos videamus quid sit melius
JOB|34|5|quia dixit Iob iustus sum et Deus subvertit iudicium meum
JOB|34|6|in iudicando enim me mendacium est violenta sagitta mea absque ullo peccato
JOB|34|7|quis est vir ut est Iob qui bibit subsannationem quasi aquam
JOB|34|8|qui graditur cum operantibus iniquitatem et ambulat cum viris impiis
JOB|34|9|dixit enim non placebit vir Deo etiam si cucurrerit cum eo
JOB|34|10|ideo viri cordati audite me absit a Deo impietas et ab Omnipotente iniquitas
JOB|34|11|opus enim hominis reddet ei et iuxta vias singulorum restituet
JOB|34|12|vere enim Deus non condemnabit frustra nec Omnipotens subvertet iudicium
JOB|34|13|quem constituit alium super terram aut quem posuit super orbem quem fabricatus est
JOB|34|14|si direxerit ad eum cor suum spiritum illius et flatum ad se trahet
JOB|34|15|deficiet omnis caro simul et homo in cinerem revertetur
JOB|34|16|si habes ergo intellectum audi quod dicitur et ausculta vocem eloquii mei
JOB|34|17|numquid qui non amat iudicium sanare potest et quomodo tu eum qui iustus est in tantum condemnas
JOB|34|18|qui dicit regi apostata qui vocat duces impios
JOB|34|19|qui non accipit personas principum nec cognovit tyrannum cum disceptaret contra pauperem opus enim manuum eius sunt universi
JOB|34|20|subito morientur et in media nocte turbabuntur populi et pertransibunt et auferent violentum absque manu
JOB|34|21|oculi enim eius super vias hominum et omnes gressus eorum considerat
JOB|34|22|non sunt tenebrae et non est umbra mortis ut abscondantur ibi qui operantur iniquitatem
JOB|34|23|neque enim ultra in hominis potestate est ut veniat ad Deum in iudicium
JOB|34|24|conteret multos innumerabiles et stare faciet alios pro eis
JOB|34|25|novit enim opera eorum et idcirco inducet noctem et conterentur
JOB|34|26|quasi impios percussit eos in loco videntium
JOB|34|27|qui quasi de industria recesserunt ab eo et omnes vias eius intellegere noluerunt
JOB|34|28|ut pervenire facerent ad eum clamorem egeni et audiret vocem pauperum
JOB|34|29|ipso enim concedente pacem quis est qui condemnet ex quo absconderit vultum quis est qui contempletur eum et super gentem et super omnes homines
JOB|34|30|qui regnare facit hominem hypocritam propter peccata populi
JOB|34|31|quia ergo ego locutus sum ad Deum te quoque non prohibeo
JOB|34|32|si erravi tu doce me si iniquitatem locutus sum ultra non addam
JOB|34|33|numquid a te Deus expetit eam quia displicuit tibi tu enim coepisti loqui et non ego quod si quid nosti melius loquere
JOB|34|34|viri intellegentes loquantur mihi et vir sapiens audiat me
JOB|34|35|Iob autem stulte locutus est et verba illius non sonant disciplinam
JOB|34|36|pater mi probetur Iob usque ad finem ne desinas in hominibus iniquitatis
JOB|34|37|quia addit super peccata sua blasphemiam inter nos interim constringatur et tunc ad iudicium provocet sermonibus suis Deum
JOB|35|1|igitur Heliu haec rursum locutus est
JOB|35|2|numquid aequa tibi videtur tua cogitatio ut diceres iustior Deo sum
JOB|35|3|dixisti enim non tibi placet quod rectum est vel quid tibi proderit si ego peccavero
JOB|35|4|itaque ego respondebo sermonibus tuis et amicis tuis tecum
JOB|35|5|suspice caelum et intuere et contemplare aethera quod altior te sit
JOB|35|6|si peccaveris quid ei nocebis et si multiplicatae fuerint iniquitates tuae quid facies contra eum
JOB|35|7|porro si iuste egeris quid donabis ei aut quid de manu tua accipiet
JOB|35|8|homini qui similis tui est nocebit impietas tua et filium hominis adiuvabit iustitia tua
JOB|35|9|propter multitudinem calumniatorum clamabunt et heiulabunt propter vim brachii tyrannorum
JOB|35|10|et non dixit ubi est Deus qui fecit me qui dedit carmina in nocte
JOB|35|11|qui docet nos super iumenta terrae et super volucres caeli erudit nos
JOB|35|12|ibi clamabunt et non exaudiet propter superbiam malorum
JOB|35|13|non ergo frustra audiet Deus et Omnipotens singulorum causas intuebitur
JOB|35|14|etiam cum dixeris non considerat iudicare coram eo et expecta eum
JOB|35|15|nunc enim non infert furorem suum nec ulciscitur scelus valde
JOB|35|16|ergo Iob frustra aperit os suum et absque scientia verba multiplicat
JOB|36|1|addens quoque Heliu haec locutus est
JOB|36|2|sustine me paululum et indicabo tibi adhuc enim habeo quod pro Deo loquar
JOB|36|3|repetam scientiam meam a principio et operatorem meum probabo iustum
JOB|36|4|vere enim absque mendacio sermones mei et perfecta scientia probabitur tibi
JOB|36|5|Deus potentes non abicit cum et ipse sit potens
JOB|36|6|sed non salvat impios et iudicium pauperibus tribuit
JOB|36|7|non aufert a iusto oculos suos et reges in solio conlocat in perpetuum et illi eriguntur
JOB|36|8|et si fuerint in catenis et vinciantur funibus paupertatis
JOB|36|9|indicabit eis opera eorum et scelera eorum quia violenti fuerint
JOB|36|10|revelabit quoque aurem eorum ut corripiat et loquetur ut revertantur ab iniquitate
JOB|36|11|si audierint et observaverint conplebunt dies suos in bono et annos suos in gloria
JOB|36|12|si autem non audierint transibunt per gladium et consumentur in stultitia
JOB|36|13|simulatores et callidi provocant iram Dei neque clamabunt cum vincti fuerint
JOB|36|14|morietur in tempestate anima eorum et vita eorum inter effeminatos
JOB|36|15|eripiet pauperem de angustia sua et revelabit in tribulatione aurem eius
JOB|36|16|igitur salvabit te de ore angusto latissime et non habentis fundamentum subter se requies autem mensae tuae erit plena pinguedine
JOB|36|17|causa tua quasi impii iudicata est causam iudiciumque recipies
JOB|36|18|non te ergo superet ira ut aliquem opprimas nec multitudo donorum inclinet te
JOB|36|19|depone magnitudinem tuam absque tribulatione et omnes robustos fortitudine
JOB|36|20|ne protrahas noctem ut ascendant populi pro eis
JOB|36|21|cave ne declines ad iniquitatem hanc enim coepisti sequi post miseriam
JOB|36|22|ecce Deus excelsus in fortitudine sua et nullus ei similis in legislatoribus
JOB|36|23|quis poterit scrutari vias eius aut quis ei dicere operatus es iniquitatem
JOB|36|24|memento quod ignores opus eius de quo cecinerunt viri
JOB|36|25|omnes homines vident eum unusquisque intuetur procul
JOB|36|26|ecce Deus magnus vincens scientiam nostram numerus annorum eius inaestimabilis
JOB|36|27|qui aufert stillas pluviae et effundit imbres ad instar gurgitum
JOB|36|28|qui de nubibus fluunt quae praetexunt cuncta desuper
JOB|36|29|si voluerit extendere nubes quasi tentorium suum
JOB|36|30|et fulgurare lumine suo desuper cardines quoque maris operiet
JOB|36|31|per haec enim iudicat populos et dat escas multis mortalibus
JOB|36|32|in manibus abscondit lucem et praecipit ei ut rursus adveniat
JOB|36|33|adnuntiat de ea amico suo quod possessio eius sit et ad eam possit ascendere
JOB|37|1|super hoc expavit cor meum et emotum est de loco suo
JOB|37|2|audite auditionem in terrore vocis eius et sonum de ore illius procedentem
JOB|37|3|subter omnes caelos ipse considerat et lumen illius super terminos terrae
JOB|37|4|post eum rugiet sonitus tonabit voce magnitudinis suae et non investigabitur cum audita fuerit vox eius
JOB|37|5|tonabit Deus in voce sua mirabiliter qui facit magna et inscrutabilia
JOB|37|6|qui praecipit nivi ut descendat in terram et hiemis pluviis et imbri fortitudinis suae
JOB|37|7|qui in manu omnium hominum signat ut noverint singuli opera sua
JOB|37|8|ingredietur bestia latibulum et in antro suo morabitur
JOB|37|9|ab interioribus egreditur tempestas et ab Arcturo frigus
JOB|37|10|flante Deo concrescit gelu et rursum latissimae funduntur aquae
JOB|37|11|frumentum desiderat nubes et nubes spargunt lumen suum
JOB|37|12|quae lustrant per circuitum quocumque eas voluntas gubernantis duxerit ad omne quod praeceperit illis super faciem orbis terrarum
JOB|37|13|sive in una tribu sive in terra sua sive in quocumque loco misericordiae suae eas iusserit inveniri
JOB|37|14|ausculta haec Iob sta et considera miracula Dei
JOB|37|15|numquid scis quando praeceperit Deus pluviis ut ostenderent lucem nubium eius
JOB|37|16|numquid nosti semitas nubium magnas et perfectas scientias
JOB|37|17|nonne vestimenta tua calida sunt cum perflata fuerit terra austro
JOB|37|18|tu forsitan cum eo fabricatus es caelos qui solidissimi quasi aere fusi sunt
JOB|37|19|ostende nobis quid dicamus illi nos quippe involvimur tenebris
JOB|37|20|quis narrabit ei quae loquor etiam si locutus fuerit homo devorabitur
JOB|37|21|at nunc non vident lucem subito aer cogitur in nubes et ventus transiens fugabit eas
JOB|37|22|ab aquilone aurum venit et ad Deum formidolosa laudatio
JOB|37|23|digne eum invenire non possumus magnus fortitudine et iudicio et iustitia et enarrari non potest
JOB|37|24|ideo timebunt eum viri et non audebunt contemplari omnes qui sibi videntur esse sapientes
JOB|38|1|respondens autem Dominus Iob de turbine dixit
JOB|38|2|quis est iste involvens sententias sermonibus inperitis
JOB|38|3|accinge sicut vir lumbos tuos interrogabo te et responde mihi
JOB|38|4|ubi eras quando ponebam fundamenta terrae indica mihi si habes intellegentiam
JOB|38|5|quis posuit mensuras eius si nosti vel quis tetendit super eam lineam
JOB|38|6|super quo bases illius solidatae sunt aut quis dimisit lapidem angularem eius
JOB|38|7|cum me laudarent simul astra matutina et iubilarent omnes filii Dei
JOB|38|8|quis conclusit ostiis mare quando erumpebat quasi de vulva procedens
JOB|38|9|cum ponerem nubem vestimentum eius et caligine illud quasi pannis infantiae obvolverem
JOB|38|10|circumdedi illud terminis meis et posui vectem et ostia
JOB|38|11|et dixi usque huc venies et non procedes amplius et hic confringes tumentes fluctus tuos
JOB|38|12|numquid post ortum tuum praecepisti diluculo et ostendisti aurorae locum suum
JOB|38|13|et tenuisti concutiens extrema terrae et excussisti impios ex ea
JOB|38|14|restituetur ut lutum signaculum et stabit sicut vestimentum
JOB|38|15|auferetur ab impiis lux sua et brachium excelsum confringetur
JOB|38|16|numquid ingressus es profunda maris et in novissimis abyssis deambulasti
JOB|38|17|numquid apertae tibi sunt portae mortis et ostia tenebrosa vidisti
JOB|38|18|numquid considerasti latitudines terrae indica mihi si nosti omnia
JOB|38|19|in qua via habitet lux et tenebrarum quis locus sit
JOB|38|20|ut ducas unumquodque ad terminos suos et intellegas semitas domus eius
JOB|38|21|sciebas tunc quod nasciturus esses et numerum dierum tuorum noveras
JOB|38|22|numquid ingressus es thesauros nivis aut thesauros grandinis aspexisti
JOB|38|23|quae praeparavi in tempus hostis in diem pugnae et belli
JOB|38|24|per quam viam spargitur lux dividitur aestus super terram
JOB|38|25|quis dedit vehementissimo imbri cursum et viam sonantis tonitrui
JOB|38|26|ut plueret super terram absque homine in deserto ubi nullus mortalium commoratur
JOB|38|27|ut impleret inviam et desolatam et produceret herbas virentes
JOB|38|28|quis est pluviae pater vel quis genuit stillas roris
JOB|38|29|de cuius utero egressa est glacies et gelu de caelo quis genuit
JOB|38|30|in similitudinem lapidis aquae durantur et superficies abyssi constringitur
JOB|38|31|numquid coniungere valebis micantes stellas Pliadis aut gyrum Arcturi poteris dissipare
JOB|38|32|numquid producis luciferum in tempore suo et vesperum super filios terrae consurgere facis
JOB|38|33|numquid nosti ordinem caeli et pones rationem eius in terra
JOB|38|34|numquid elevabis in nebula vocem tuam et impetus aquarum operiet te
JOB|38|35|numquid mittes fulgura et ibunt et revertentia dicent tibi adsumus
JOB|38|36|quis posuit in visceribus hominis sapientiam vel quis dedit gallo intellegentiam
JOB|38|37|quis enarravit caelorum rationem et concentum caeli quis dormire faciet
JOB|38|38|quando fundebatur pulvis in terram et glebae conpingebantur
JOB|38|39|numquid capies leaenae praedam et animam catulorum eius implebis
JOB|38|40|quando cubant in antris et in specubus insidiantur
JOB|38|41|quis praeparat corvo escam suam quando pulli eius ad Deum clamant vagantes eo quod non habeant cibos
JOB|39|1|numquid nosti tempus partus hibicum in petris vel parturientes cervas observasti
JOB|39|2|dinumerasti menses conceptus earum et scisti tempus partus earum
JOB|39|3|incurvantur ad fetum et pariunt et rugitus emittunt
JOB|39|4|separantur filii earum pergunt ad pastum egrediuntur et non revertuntur ad eas
JOB|39|5|quis dimisit onagrum liberum et vincula eius quis solvit
JOB|39|6|cui dedi in solitudine domum et tabernacula eius in terra salsuginis
JOB|39|7|contemnit multitudinem civitatis clamorem exactoris non audit
JOB|39|8|circumspicit montes pascuae suae et virentia quaeque perquirit
JOB|39|9|numquid volet rinoceros servire tibi aut morabitur ad praesepe tuum
JOB|39|10|numquid alligabis rinocerota ad arandum loro tuo aut confringet glebas vallium post te
JOB|39|11|numquid fiduciam habebis in magna fortitudine eius et derelinques ei labores tuos
JOB|39|12|numquid credes ei quoniam reddat sementem tibi et aream tuam congreget
JOB|39|13|pinna strutionum similis est pinnis herodii et accipitris
JOB|39|14|quando derelinquit in terra ova sua tu forsitan in pulvere calefacis ea
JOB|39|15|obliviscitur quod pes conculcet ea aut bestiae agri conterant
JOB|39|16|duratur ad filios suos quasi non sint sui frustra laboravit nullo timore cogente
JOB|39|17|privavit enim eam Deus sapientia nec dedit illi intellegentiam
JOB|39|18|cum tempus fuerit in altum alas erigit deridet equitem et ascensorem eius
JOB|39|19|numquid praebebis equo fortitudinem aut circumdabis collo eius hinnitum
JOB|39|20|numquid suscitabis eum quasi lucustas gloria narium eius terror
JOB|39|21|terram ungula fodit exultat audacter in occursum pergit armatis
JOB|39|22|contemnit pavorem nec cedit gladio
JOB|39|23|super ipsum sonabit faretra vibrabit hasta et clypeus
JOB|39|24|fervens et fremens sorbet terram nec reputat tubae sonare clangorem
JOB|39|25|ubi audierit bucinam dicet va procul odoratur bellum exhortationem ducum et ululatum exercitus
JOB|39|26|numquid per sapientiam tuam plumescit accipiter expandens alas suas ad austrum
JOB|39|27|aut ad praeceptum tuum elevabitur aquila et in arduis ponet nidum suum
JOB|39|28|in petris manet et in praeruptis silicibus commoratur atque inaccessis rupibus
JOB|39|29|inde contemplatur escam et de longe oculi eius prospiciunt
JOB|39|30|pulli eius lambent sanguinem et ubicumque cadaver fuerit statim adest
JOB|39|31|et adiecit Dominus et locutus est ad Iob
JOB|39|32|numquid qui contendit cum Deo tam facile conquiescit utique qui arguit Deum debet respondere ei
JOB|39|33|respondens autem Iob Domino dixit
JOB|39|34|qui leviter locutus sum respondere quid possum manum meam ponam super os meum
JOB|39|35|unum locutus sum quod utinam non dixissem et alterum quibus ultra non addam
JOB|40|1|respondens autem Dominus Iob de turbine ait
JOB|40|2|accinge sicut vir lumbos tuos interrogabo te et indica mihi
JOB|40|3|numquid irritum facies iudicium meum et condemnabis me ut tu iustificeris
JOB|40|4|et si habes brachium sicut Deus et si voce simili tonas
JOB|40|5|circumda tibi decorem et in sublime erigere et esto gloriosus et speciosis induere vestibus
JOB|40|6|disperge superbos furore tuo et respiciens omnem arrogantem humilia
JOB|40|7|respice cunctos superbos et confunde eos et contere impios in loco suo
JOB|40|8|absconde eos in pulvere simul et facies eorum demerge in foveam
JOB|40|9|et ego confitebor quod salvare te possit dextera tua
JOB|40|10|ecce Behemoth quem feci tecum faenum quasi bos comedet
JOB|40|11|fortitudo eius in lumbis eius et virtus illius in umbilicis ventris eius
JOB|40|12|constringit caudam suam quasi cedrum nervi testiculorum eius perplexi sunt
JOB|40|13|ossa eius velut fistulae aeris cartilago illius quasi lamminae ferreae
JOB|40|14|ipse principium est viarum Dei qui fecit eum adplicabit gladium eius
JOB|40|15|huic montes herbas ferunt omnes bestiae agri ludent ibi
JOB|40|16|sub umbra dormit in secreto calami et locis humentibus
JOB|40|17|protegunt umbrae umbram eius circumdabunt eum salices torrentis
JOB|40|18|ecce absorbebit fluvium et non mirabitur habet fiduciam quod influat Iordanis in os eius
JOB|40|19|in oculis eius quasi hamo capiet eum et in sudibus perforabit nares eius
JOB|40|20|an extrahere poteris Leviathan hamo et fune ligabis linguam eius
JOB|40|21|numquid pones circulum in naribus eius et armilla perforabis maxillam eius
JOB|40|22|numquid multiplicabit ad te preces aut loquetur tibi mollia
JOB|40|23|numquid feriet tecum pactum et accipies eum servum sempiternum
JOB|40|24|numquid inludes ei quasi avi aut ligabis illum ancillis tuis
JOB|40|25|concident eum amici divident illum negotiatores
JOB|40|26|numquid implebis sagenas pelle eius et gurgustium piscium capite illius
JOB|40|27|pone super eum manum tuam memento belli nec ultra addas loqui
JOB|40|28|ecce spes eius frustrabitur eum et videntibus cunctis praecipitabitur
JOB|41|1|non quasi crudelis suscitabo eum quis enim resistere potest vultui meo
JOB|41|2|quis ante dedit mihi ut reddam ei omnia quae sub caelo sunt mea sunt
JOB|41|3|non parcam ei et verbis potentibus et ad deprecandum conpositis
JOB|41|4|quis revelavit faciem indumenti eius et in medium oris eius quis intrabit
JOB|41|5|portas vultus eius quis aperiet per gyrum dentium eius formido
JOB|41|6|corpus illius quasi scuta fusilia et conpactum squamis se prementibus
JOB|41|7|una uni coniungitur et ne spiraculum quidem incedit per eas
JOB|41|8|una alteri adherebunt et tenentes se nequaquam separabuntur
JOB|41|9|sternutatio eius splendor ignis et oculi eius ut palpebrae diluculi
JOB|41|10|de ore eius lampades procedunt sicut taedae ignis accensae
JOB|41|11|de naribus eius procedit fumus sicut ollae succensae atque ferventis
JOB|41|12|halitus eius prunas ardere facit et flamma de ore eius egreditur
JOB|41|13|in collo eius morabitur fortitudo et faciem eius praecedet egestas
JOB|41|14|membra carnium eius coherentia sibi mittet contra eum fulmina et ad locum alium non ferentur
JOB|41|15|cor eius indurabitur quasi lapis et stringetur quasi malleatoris incus
JOB|41|16|cum sublatus fuerit timebunt angeli et territi purgabuntur
JOB|41|17|cum adprehenderit eum gladius subsistere non poterit neque hasta neque torax
JOB|41|18|reputabit enim quasi paleas ferrum et quasi lignum putridum aes
JOB|41|19|non fugabit eum vir sagittarius in stipulam versi sunt ei lapides fundae
JOB|41|20|quasi stipulam aestimabit malleum et deridebit vibrantem hastam
JOB|41|21|sub ipso erunt radii solis sternet sibi aurum quasi lutum
JOB|41|22|fervescere faciet quasi ollam profundum mare ponet quasi cum unguenta bulliunt
JOB|41|23|post eum lucebit semita aestimabit abyssum quasi senescentem
JOB|41|24|non est super terram potestas quae conparetur ei qui factus est ut nullum timeret
JOB|41|25|omne sublime videt ipse est rex super universos filios superbiae
JOB|42|1|respondens autem Iob Domino dixit
JOB|42|2|scio quia omnia potes et nulla te latet cogitatio
JOB|42|3|quis est iste qui celat consilium absque scientia ideo insipienter locutus sum et quae ultra modum excederent scientiam meam
JOB|42|4|audi et ego loquar interrogabo et ostende mihi
JOB|42|5|auditu auris audivi te nunc autem oculus meus videt te
JOB|42|6|idcirco ipse me reprehendo et ago paenitentiam in favilla et cinere
JOB|42|7|postquam autem locutus est Dominus verba haec ad Iob dixit ad Eliphaz Themaniten iratus est furor meus in te et in duos amicos tuos quoniam non estis locuti coram me rectum sicut servus meus Iob
JOB|42|8|sumite igitur vobis septem tauros et septem arietes et ite ad servum meum Iob et offerte holocaustum pro vobis Iob autem servus meus orabit pro vobis faciem eius suscipiam ut non vobis inputetur stultitia neque enim locuti estis ad me recta sicut servus meus Iob
JOB|42|9|abierunt ergo Eliphaz Themanites et Baldad Suites et Sophar Naamathites et fecerunt sicut locutus fuerat ad eos Dominus et suscepit Dominus faciem Iob
JOB|42|10|Dominus quoque conversus est ad paenitentiam Iob cum oraret ille pro amicis suis et addidit Dominus omnia quaecumque fuerant Iob duplicia
JOB|42|11|venerunt autem ad eum omnes fratres sui et universae sorores suae et cuncti qui noverant eum prius et comederunt cum eo panem in domo eius et moverunt super eum caput et consolati sunt eum super omni malo quod intulerat Dominus super eum et dederunt ei unusquisque ovem unam et inaurem auream unam
JOB|42|12|Dominus autem benedixit novissimis Iob magis quam principio eius et facta sunt ei quattuordecim milia ovium et sex milia camelorum et mille iuga boum et mille asinae
JOB|42|13|et fuerunt ei septem filii et filiae tres
JOB|42|14|et vocavit nomen unius Diem et nomen secundae Cassia et nomen tertiae Cornu stibii
JOB|42|15|non sunt autem inventae mulieres speciosae sicut filiae Iob in universa terra deditque eis pater suus hereditatem inter fratres earum
JOB|42|16|vixit autem Iob post haec centum quadraginta annis et vidit filios suos et filios filiorum suorum usque ad quartam generationem et mortuus est senex et plenus dierum
