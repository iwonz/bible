3JOHN|1|1|senior Gaio carissimo quem ego diligo in veritate
3JOHN|1|2|carissime de omnibus orationem facio prospere te ingredi et valere sicut prospere agit anima tua
3JOHN|1|3|gavisus sum valde venientibus fratribus et testimonium perhibentibus veritati tuae sicut tu in veritate ambulas
3JOHN|1|4|maiorem horum non habeo gratiam quam ut audiam filios meos in veritate ambulantes
3JOHN|1|5|carissime fideliter facis quicquid operaris in fratres et hoc in peregrinos
3JOHN|1|6|qui testimonium reddiderunt caritati tuae in conspectu ecclesiae quos bene facies deducens digne Deo
3JOHN|1|7|pro nomine enim profecti sunt nihil accipientes a gentibus
3JOHN|1|8|nos ergo debemus suscipere huiusmodi ut cooperatores simus veritatis
3JOHN|1|9|scripsissem forsitan ecclesiae sed is qui amat primatum gerere in eis Diotrepes non recipit nos
3JOHN|1|10|propter hoc si venero commoneam eius opera quae facit verbis malignis garriens in nos et quasi non ei ista sufficiant nec ipse suscipit fratres et eos qui cupiunt prohibet et de ecclesia eicit
3JOHN|1|11|carissime noli imitari malum sed quod bonum est qui benefacit ex Deo est qui malefacit non vidit Deum
3JOHN|1|12|Demetrio testimonium redditur ab omnibus et ab ipsa veritate et nos autem testimonium perhibemus et nosti quoniam testimonium nostrum verum est
3JOHN|1|13|multa habui scribere tibi sed nolui per atramentum et calamum scribere tibi
3JOHN|1|14|spero autem protinus te videre et os ad os loquemur
3JOHN|1|15|pax tibi salutant te amici saluta amicos per nomen
