LEV|1|1|The LORD called Moses and spoke to him from the tent of meeting, saying,
LEV|1|2|"Speak to the people of Israel and say to them, When any one of you brings an offering to the LORD, you shall bring your offering of livestock from the herd or from the flock.
LEV|1|3|"If his offering is a burnt offering from the herd, he shall offer a male without blemish. He shall bring it to the entrance of the tent of meeting, that he may be accepted before the LORD.
LEV|1|4|He shall lay his hand on the head of the burnt offering, and it shall be accepted for him to make atonement for him.
LEV|1|5|Then he shall kill the bull before the LORD, and Aaron's sons the priests shall bring the blood and throw the blood against the sides of the altar that is at the entrance of the tent of meeting.
LEV|1|6|Then he shall flay the burnt offering and cut it into pieces,
LEV|1|7|and the sons of Aaron the priest shall put fire on the altar and arrange wood on the fire.
LEV|1|8|And Aaron's sons the priests shall arrange the pieces, the head, and the fat, on the wood that is on the fire on the altar;
LEV|1|9|but its entrails and its legs he shall wash with water. And the priest shall burn all of it on the altar, as a burnt offering, a food offering with a pleasing aroma to the LORD.
LEV|1|10|"If his gift for a burnt offering is from the flock, from the sheep or goats, he shall bring a male without blemish,
LEV|1|11|and he shall kill it on the north side of the altar before the LORD, and Aaron's sons the priests shall throw its blood against the sides of the altar.
LEV|1|12|And he shall cut it into pieces, with its head and its fat, and the priest shall arrange them on the wood that is on the fire on the altar,
LEV|1|13|but the entrails and the legs he shall wash with water. And the priest shall offer all of it and burn it on the altar; it is a burnt offering, a food offering with a pleasing aroma to the LORD.
LEV|1|14|"If his offering to the LORD is a burnt offering of birds, then he shall bring his offering of turtledoves or pigeons.
LEV|1|15|And the priest shall bring it to the altar and wring off its head and burn it on the altar. Its blood shall be drained out on the side of the altar.
LEV|1|16|He shall remove its crop with its contents and cast it beside the altar on the east side, in the place for ashes.
LEV|1|17|He shall tear it open by its wings, but shall not sever it completely. And the priest shall burn it on the altar, on the wood that is on the fire. It is a burnt offering, a food offering with a pleasing aroma to the LORD.
LEV|2|1|"When anyone brings a grain offering as an offering to the LORD, his offering shall be of fine flour. He shall pour oil on it and put frankincense on it
LEV|2|2|and bring it to Aaron's sons the priests. And he shall take from it a handful of the fine flour and oil, with all of its frankincense, and the priest shall burn this as its memorial portion on the altar, a food offering with a pleasing aroma to the LORD.
LEV|2|3|But the rest of the grain offering shall be for Aaron and his sons; it is a most holy part of the LORD's food offerings.
LEV|2|4|"When you bring a grain offering baked in the oven as an offering, it shall be unleavened loaves of fine flour mixed with oil or unleavened wafers smeared with oil.
LEV|2|5|And if your offering is a grain offering baked on a griddle, it shall be of fine flour unleavened, mixed with oil.
LEV|2|6|You shall break it in pieces and pour oil on it; it is a grain offering.
LEV|2|7|And if your offering is a grain offering cooked in a pan, it shall be made of fine flour with oil.
LEV|2|8|And you shall bring the grain offering that is made of these things to the LORD, and when it is presented to the priest, he shall bring it to the altar.
LEV|2|9|And the priest shall take from the grain offering its memorial portion and burn this on the altar, a food offering with a pleasing aroma to the LORD.
LEV|2|10|But the rest of the grain offering shall be for Aaron and his sons; it is a most holy part of the LORD's food offerings.
LEV|2|11|"No grain offering that you bring to the LORD shall be made with leaven, for you shall burn no leaven nor any honey as a food offering to the LORD.
LEV|2|12|As an offering of firstfruits you may bring them to the LORD, but they shall not be offered on the altar for a pleasing aroma.
LEV|2|13|You shall season all your grain offerings with salt. You shall not let the salt of the covenant with your God be missing from your grain offering; with all your offerings you shall offer salt.
LEV|2|14|"If you offer a grain offering of firstfruits to the LORD, you shall offer for the grain offering of your firstfruits fresh ears, roasted with fire, crushed new grain.
LEV|2|15|And you shall put oil on it and lay frankincense on it; it is a grain offering.
LEV|2|16|And the priest shall burn as its memorial portion some of the crushed grain and some of the oil with all of its frankincense; it is a food offering to the LORD.
LEV|3|1|"If his offering is a sacrifice of peace offering, if he offers an animal from the herd, male or female, he shall offer it without blemish before the LORD.
LEV|3|2|And he shall lay his hand on the head of his offering and kill it at the entrance of the tent of meeting, and Aaron's sons the priests shall throw the blood against the sides of the altar.
LEV|3|3|And from the sacrifice of the peace offering, as a food offering to the LORD, he shall offer the fat covering the entrails and all the fat that is on the entrails,
LEV|3|4|and the two kidneys with the fat that is on them at the loins, and the long lobe of the liver that he shall remove with the kidneys.
LEV|3|5|Then Aaron's sons shall burn it on the altar on top of the burnt offering, which is on the wood on the fire; it is a food offering with a pleasing aroma to the LORD.
LEV|3|6|"If his offering for a sacrifice of peace offering to the LORD is an animal from the flock, male or female, he shall offer it without blemish.
LEV|3|7|If he offers a lamb for his offering, then he shall offer it before the LORD,
LEV|3|8|lay his hand on the head of his offering, and kill it in front of the tent of meeting; and Aaron's sons shall throw its blood against the sides of the altar.
LEV|3|9|Then from the sacrifice of the peace offering he shall offer as a food offering to the LORD its fat; he shall remove the whole fat tail, cut off close to the backbone, and the fat that covers the entrails and all the fat that is on the entrails
LEV|3|10|and the two kidneys with the fat that is on them at the loins and the long lobe of the liver that he shall remove with the kidneys.
LEV|3|11|And the priest shall burn it on the altar as a food offering to the LORD.
LEV|3|12|"If his offering is a goat, then he shall offer it before the LORD
LEV|3|13|and lay his hand on its head and kill it in front of the tent of meeting, and the sons of Aaron shall throw its blood against the sides of the altar.
LEV|3|14|Then he shall offer from it, as his offering for a food offering to the LORD, the fat covering the entrails and all the fat that is on the entrails
LEV|3|15|and the two kidneys with the fat that is on them at the loins and the long lobe of the liver that he shall remove with the kidneys.
LEV|3|16|And the priest shall burn them on the altar as a food offering with a pleasing aroma. All fat is the LORD's.
LEV|3|17|It shall be a statute forever throughout your generations, in all your dwelling places, that you eat neither fat nor blood."
LEV|4|1|And the LORD spoke to Moses, saying,
LEV|4|2|"Speak to the people of Israel, saying, If anyone sins unintentionally in any of the LORD's commandments about things not to be done, and does any one of them,
LEV|4|3|if it is the anointed priest who sins, thus bringing guilt on the people, then he shall offer for the sin that he has committed a bull from the herd without blemish to the LORD for a sin offering.
LEV|4|4|He shall bring the bull to the entrance of the tent of meeting before the LORD and lay his hand on the head of the bull and kill the bull before the LORD.
LEV|4|5|And the anointed priest shall take some of the blood of the bull and bring it into the tent of meeting,
LEV|4|6|and the priest shall dip his finger in the blood and sprinkle part of the blood seven times before the LORD in front of the veil of the sanctuary.
LEV|4|7|And the priest shall put some of the blood on the horns of the altar of fragrant incense before the LORD that is in the tent of meeting, and all the rest of the blood of the bull he shall pour out at the base of the altar of burnt offering that is at the entrance of the tent of meeting.
LEV|4|8|And all the fat of the bull of the sin offering he shall remove from it, the fat that covers the entrails and all the fat that is on the entrails
LEV|4|9|and the two kidneys with the fat that is on them at the loins and the long lobe of the liver that he shall remove with the kidneys
LEV|4|10|(just as these are taken from the ox of the sacrifice of the peace offerings); and the priest shall burn them on the altar of burnt offering.
LEV|4|11|But the skin of the bull and all its flesh, with its head, its legs, its entrails, and its dung-
LEV|4|12|all the rest of the bull- he shall carry outside the camp to a clean place, to the ash heap, and shall burn it up on a fire of wood. On the ash heap it shall be burned up.
LEV|4|13|"If the whole congregation of Israel sins unintentionally and the thing is hidden from the eyes of the assembly, and they do any one of the things that by the LORD's commandments ought not to be done, and they realize their guilt,
LEV|4|14|when the sin which they have committed becomes known, the assembly shall offer a bull from the herd for a sin offering and bring it in front of the tent of meeting.
LEV|4|15|And the elders of the congregation shall lay their hands on the head of the bull before the LORD, and the bull shall be killed before the LORD.
LEV|4|16|Then the anointed priest shall bring some of the blood of the bull into the tent of meeting,
LEV|4|17|and the priest shall dip his finger in the blood and sprinkle it seven times before the LORD in front of the veil.
LEV|4|18|And he shall put some of the blood on the horns of the altar that is in the tent of meeting before the LORD, and the rest of the blood he shall pour out at the base of the altar of burnt offering that is at the entrance of the tent of meeting.
LEV|4|19|And all its fat he shall take from it and burn on the altar.
LEV|4|20|Thus shall he do with the bull. As he did with the bull of the sin offering, so shall he do with this. And the priest shall make atonement for them, and they shall be forgiven.
LEV|4|21|And he shall carry the bull outside the camp and burn it up as he burned the first bull; it is the sin offering for the assembly.
LEV|4|22|"When a leader sins, doing unintentionally any one of all the things that by the commandments of the LORD his God ought not to be done, and realizes his guilt,
LEV|4|23|or the sin which he has committed is made known to him, he shall bring as his offering a goat, a male without blemish,
LEV|4|24|and shall lay his hand on the head of the goat and kill it in the place where they kill the burnt offering before the LORD; it is a sin offering.
LEV|4|25|Then the priest shall take some of the blood of the sin offering with his finger and put it on the horns of the altar of burnt offering and pour out the rest of its blood at the base of the altar of burnt offering.
LEV|4|26|And all its fat he shall burn on the altar, like the fat of the sacrifice of peace offerings. So the priest shall make atonement for him for his sin, and he shall be forgiven.
LEV|4|27|"If anyone of the common people sins unintentionally in doing any one of the things that by the LORD's commandments ought not to be done, and realizes his guilt,
LEV|4|28|or the sin which he has committed is made known to him, he shall bring for his offering a goat, a female without blemish, for his sin which he has committed.
LEV|4|29|And he shall lay his hand on the head of the sin offering and kill the sin offering in the place of burnt offering.
LEV|4|30|And the priest shall take some of its blood with his finger and put it on the horns of the altar of burnt offering and pour out all the rest of its blood at the base of the altar.
LEV|4|31|And all its fat he shall remove, as the fat is removed from the peace offerings, and the priest shall burn it on the altar for a pleasing aroma to the LORD. And the priest shall make atonement for him, and he shall be forgiven.
LEV|4|32|"If he brings a lamb as his offering for a sin offering, he shall bring a female without blemish
LEV|4|33|and lay his hand on the head of the sin offering and kill it for a sin offering in the place where they kill the burnt offering.
LEV|4|34|Then the priest shall take some of the blood of the sin offering with his finger and put it on the horns of the altar of burnt offering and pour out all the rest of its blood at the base of the altar.
LEV|4|35|And all its fat he shall remove as the fat of the lamb is removed from the sacrifice of peace offerings, and the priest shall burn it on the altar, on top of the LORD's food offerings. And the priest shall make atonement for him for the sin which he has committed, and he shall be forgiven.
LEV|5|1|"If anyone sins in that he hears a public adjuration to testify, and though he is a witness, whether he has seen or come to know the matter, yet does not speak, he shall bear his iniquity;
LEV|5|2|or if anyone touches an unclean thing, whether a carcass of an unclean wild animal or a carcass of unclean livestock or a carcass of unclean swarming things, and it is hidden from him and he has become unclean, and he realizes his guilt;
LEV|5|3|or if he touches human uncleanness, of whatever sort the uncleanness may be with which one becomes unclean, and it is hidden from him, when he comes to know it, and realizes his guilt;
LEV|5|4|or if anyone utters with his lips a rash oath to do evil or to do good, any sort of rash oath that people swear, and it is hidden from him, when he comes to know it, and he realizes his guilt in any of these;
LEV|5|5|when he realizes his guilt in any of these and confesses the sin he has committed,
LEV|5|6|he shall bring to the LORD as his compensation for the sin that he has committed, a female from the flock, a lamb or a goat, for a sin offering. And the priest shall make atonement for him for his sin.
LEV|5|7|"But if he cannot afford a lamb, then he shall bring to the LORD as his compensation for the sin that he has committed two turtledoves or two pigeons, one for a sin offering and the other for a burnt offering.
LEV|5|8|He shall bring them to the priest, who shall offer first the one for the sin offering. He shall wring its head from its neck but shall not sever it completely,
LEV|5|9|and he shall sprinkle some of the blood of the sin offering on the side of the altar, while the rest of the blood shall be drained out at the base of the altar; it is a sin offering.
LEV|5|10|Then he shall offer the second for a burnt offering according to the rule. And the priest shall make atonement for him for the sin that he has committed, and he shall be forgiven.
LEV|5|11|"But if he cannot afford two turtledoves or two pigeons, then he shall bring as his offering for the sin that he has committed a tenth of an ephah of fine flour for a sin offering. He shall put no oil on it and shall put no frankincense on it, for it is a sin offering.
LEV|5|12|And he shall bring it to the priest, and the priest shall take a handful of it as its memorial portion and burn this on the altar, on the LORD's food offerings; it is a sin offering.
LEV|5|13|Thus the priest shall make atonement for him for the sin which he has committed in any one of these things, and he shall be forgiven. And the remainder shall be for the priest, as in the grain offering."
LEV|5|14|The LORD spoke to Moses, saying,
LEV|5|15|"If anyone commits a breach of faith and sins unintentionally in any of the holy things of the LORD, he shall bring to the LORD as his compensation, a ram without blemish out of the flock, valued in silver shekels, according to the shekel of the sanctuary, for a guilt offering.
LEV|5|16|He shall also make restitution for what he has done amiss in the holy thing and shall add a fifth to it and give it to the priest. And the priest shall make atonement for him with the ram of the guilt offering, and he shall be forgiven.
LEV|5|17|"If anyone sins, doing any of the things that by the LORD's commandments ought not to be done, though he did not know it, then realizes his guilt, he shall bear his iniquity.
LEV|5|18|He shall bring to the priest a ram without blemish out of the flock, or its equivalent for a guilt offering, and the priest shall make atonement for him for the mistake that he made unintentionally, and he shall be forgiven.
LEV|5|19|It is a guilt offering; he has indeed incurred guilt before the LORD."
LEV|6|1|The LORD spoke to Moses, saying,
LEV|6|2|"If anyone sins and commits a breach of faith against the LORD by deceiving his neighbor in a matter of deposit or security, or through robbery, or if he has oppressed his neighbor
LEV|6|3|or has found something lost and lied about it, swearing falsely- in any of all the things that people do and sin thereby-
LEV|6|4|if he has sinned and has realized his guilt and will restore what he took by robbery or what he got by oppression or the deposit that was committed to him or the lost thing that he found
LEV|6|5|or anything about which he has sworn falsely, he shall restore it in full and shall add a fifth to it, and give it to him to whom it belongs on the day he realizes his guilt.
LEV|6|6|And he shall bring to the priest as his compensation to the LORD a ram without blemish out of the flock, or its equivalent for a guilt offering.
LEV|6|7|And the priest shall make atonement for him before the LORD, and he shall be forgiven for any of the things that one may do and thereby become guilty."
LEV|6|8|The LORD spoke to Moses, saying,
LEV|6|9|"Command Aaron and his sons, saying, This is the law of the burnt offering. The burnt offering shall be on the hearth on the altar all night until the morning, and the fire of the altar shall be kept burning on it.
LEV|6|10|And the priest shall put on his linen garment and put his linen undergarment on his body, and he shall take up the ashes to which the fire has reduced the burnt offering on the altar and put them beside the altar.
LEV|6|11|Then he shall take off his garments and put on other garments and carry the ashes outside the camp to a clean place.
LEV|6|12|The fire on the altar shall be kept burning on it; it shall not go out. The priest shall burn wood on it every morning, and he shall arrange the burnt offering on it and shall burn on it the fat of the peace offerings.
LEV|6|13|Fire shall be kept burning on the altar continually; it shall not go out.
LEV|6|14|"And this is the law of the grain offering. The sons of Aaron shall offer it before the LORD in front of the altar.
LEV|6|15|And one shall take from it a handful of the fine flour of the grain offering and its oil and all the frankincense that is on the grain offering and burn this as its memorial portion on the altar, a pleasing aroma to the LORD.
LEV|6|16|And the rest of it Aaron and his sons shall eat. It shall be eaten unleavened in a holy place. In the court of the tent of meeting they shall eat it.
LEV|6|17|It shall not be baked with leaven. I have given it as their portion of my food offerings. It is a thing most holy, like the sin offering and the guilt offering.
LEV|6|18|Every male among the children of Aaron may eat of it, as decreed forever throughout your generations, from the LORD's food offerings. Whatever touches them shall become holy."
LEV|6|19|The LORD spoke to Moses, saying,
LEV|6|20|"This is the offering that Aaron and his sons shall offer to the LORD on the day when he is anointed: a tenth of an ephah of fine flour as a regular grain offering, half of it in the morning and half in the evening.
LEV|6|21|It shall be made with oil on a griddle. You shall bring it well mixed, in baked pieces like a grain offering, and offer it for a pleasing aroma to the LORD.
LEV|6|22|The priest from among Aaron's sons, who is anointed to succeed him, shall offer it to the LORD as decreed forever. The whole of it shall be burned.
LEV|6|23|Every grain offering of a priest shall be wholly burned. It shall not be eaten."
LEV|6|24|The LORD spoke to Moses, saying,
LEV|6|25|"Speak to Aaron and his sons, saying, This is the law of the sin offering. In the place where the burnt offering is killed shall the sin offering be killed before the LORD; it is most holy.
LEV|6|26|The priest who offers it for sin shall eat it. In a holy place it shall be eaten, in the court of the tent of meeting.
LEV|6|27|Whatever touches its flesh shall be holy, and when any of its blood is splashed on a garment, you shall wash that on which it was splashed in a holy place.
LEV|6|28|And the earthenware vessel in which it is boiled shall be broken. But if it is boiled in a bronze vessel, that shall be scoured and rinsed in water.
LEV|6|29|Every male among the priests may eat of it; it is most holy.
LEV|6|30|But no sin offering shall be eaten from which any blood is brought into the tent of meeting to make atonement in the Holy Place; it shall be burned up with fire.
LEV|7|1|"This is the law of the guilt offering. It is most holy.
LEV|7|2|In the place where they kill the burnt offering they shall kill the guilt offering, and its blood shall be thrown against the sides of the altar.
LEV|7|3|And all its fat shall be offered, the fat tail, the fat that covers the entrails,
LEV|7|4|the two kidneys with the fat that is on them at the loins, and the long lobe of the liver that he shall remove with the kidneys.
LEV|7|5|The priest shall burn them on the altar as a food offering to the LORD; it is a guilt offering.
LEV|7|6|Every male among the priests may eat of it. It shall be eaten in a holy place. It is most holy.
LEV|7|7|The guilt offering is just like the sin offering; there is one law for them. The priest who makes atonement with it shall have it.
LEV|7|8|And the priest who offers any man's burnt offering shall have for himself the skin of the burnt offering that he has offered.
LEV|7|9|And every grain offering baked in the oven and all that is prepared on a pan or a griddle shall belong to the priest who offers it.
LEV|7|10|And every grain offering, mixed with oil or dry, shall be shared equally among all the sons of Aaron.
LEV|7|11|"And this is the law of the sacrifice of peace offerings that one may offer to the LORD.
LEV|7|12|If he offers it for a thanksgiving, then he shall offer with the thanksgiving sacrifice unleavened loaves mixed with oil, unleavened wafers smeared with oil, and loaves of fine flour well mixed with oil.
LEV|7|13|With the sacrifice of his peace offerings for thanksgiving he shall bring his offering with loaves of leavened bread.
LEV|7|14|And from it he shall offer one loaf from each offering, as a gift to the LORD. It shall belong to the priest who throws the blood of the peace offerings.
LEV|7|15|And the flesh of the sacrifice of his peace offerings for thanksgiving shall be eaten on the day of his offering. He shall not leave any of it until the morning.
LEV|7|16|But if the sacrifice of his offering is a vow offering or a freewill offering, it shall be eaten on the day that he offers his sacrifice, and on the next day what remains of it shall be eaten.
LEV|7|17|But what remains of the flesh of the sacrifice on the third day shall be burned up with fire.
LEV|7|18|If any of the flesh of the sacrifice of his peace offering is eaten on the third day, he who offers it shall not be accepted, neither shall it be credited to him. It is tainted, and he who eats of it shall bear his iniquity.
LEV|7|19|"Flesh that touches any unclean thing shall not be eaten. It shall be burned up with fire. All who are clean may eat flesh,
LEV|7|20|but the person who eats of the flesh of the sacrifice of the LORD's peace offerings while an uncleanness is on him, that person shall be cut off from his people.
LEV|7|21|And if anyone touches an unclean thing, whether human uncleanness or an unclean beast or any unclean detestable creature, and then eats some flesh from the sacrifice of the LORD's peace offerings, that person shall be cut off from his people."
LEV|7|22|The LORD spoke to Moses, saying,
LEV|7|23|"Speak to the people of Israel, saying, You shall eat no fat, of ox or sheep or goat.
LEV|7|24|The fat of an animal that dies of itself and the fat of one that is torn by beasts may be put to any other use, but on no account shall you eat it.
LEV|7|25|For every person who eats of the fat of an animal of which a food offering may be made to the LORD shall be cut off from his people.
LEV|7|26|Moreover, you shall eat no blood whatever, whether of fowl or of animal, in any of your dwelling places.
LEV|7|27|Whoever eats any blood, that person shall be cut off from his people."
LEV|7|28|The LORD spoke to Moses, saying,
LEV|7|29|"Speak to the people of Israel, saying, Whoever offers the sacrifice of his peace offerings to the LORD shall bring his offering to the LORD from the sacrifice of his peace offerings.
LEV|7|30|His own hands shall bring the LORD's food offerings. He shall bring the fat with the breast, that the breast may be waved as a wave offering before the LORD.
LEV|7|31|The priest shall burn the fat on the altar, but the breast shall be for Aaron and his sons.
LEV|7|32|And the right thigh you shall give to the priest as a contribution from the sacrifice of your peace offerings.
LEV|7|33|Whoever among the sons of Aaron offers the blood of the peace offerings and the fat shall have the right thigh for a portion.
LEV|7|34|For the breast that is waved and the thigh that is contributed I have taken from the people of Israel, out of the sacrifices of their peace offerings, and have given them to Aaron the priest and to his sons, as a perpetual due from the people of Israel.
LEV|7|35|This is the portion of Aaron and of his sons from the LORD's food offerings, from the day they were presented to serve as priests of the LORD.
LEV|7|36|The LORD commanded this to be given them by the people of Israel, from the day that he anointed them. It is a perpetual due throughout their generations."
LEV|7|37|This is the law of the burnt offering, of the grain offering, of the sin offering, of the guilt offering, of the ordination offering, and of the peace offering,
LEV|7|38|which the LORD commanded Moses on Mount Sinai, on the day that he commanded the people of Israel to bring their offerings to the LORD, in the wilderness of Sinai.
LEV|8|1|The LORD spoke to Moses, saying,
LEV|8|2|"Take Aaron and his sons with him, and the garments and the anointing oil and the bull of the sin offering and the two rams and the basket of unleavened bread.
LEV|8|3|And assemble all the congregation at the entrance of the tent of meeting."
LEV|8|4|And Moses did as the LORD commanded him, and the congregation was assembled at the entrance of the tent of meeting.
LEV|8|5|And Moses said to the congregation, "This is the thing that the LORD has commanded to be done."
LEV|8|6|And Moses brought Aaron and his sons and washed them with water.
LEV|8|7|And he put the coat on him and tied the sash around his waist and clothed him with the robe and put the ephod on him and tied the skillfully woven band of the ephod around him, binding it to him with the band.
LEV|8|8|And he placed the breastpiece on him, and in the breastpiece he put the Urim and the Thummim.
LEV|8|9|And he set the turban on his head, and on the turban, in front, he set the golden plate, the holy crown, as the LORD commanded Moses.
LEV|8|10|Then Moses took the anointing oil and anointed the tabernacle and all that was in it, and consecrated them.
LEV|8|11|And he sprinkled some of it on the altar seven times, and anointed the altar and all its utensils and the basin and its stand, to consecrate them.
LEV|8|12|And he poured some of the anointing oil on Aaron's head and anointed him to consecrate him.
LEV|8|13|And Moses brought Aaron's sons and clothed them with coats and tied sashes around their waists and bound caps on them, as the LORD commanded Moses.
LEV|8|14|Then he brought the bull of the sin offering, and Aaron and his sons laid their hands on the head of the bull of the sin offering.
LEV|8|15|And he killed it, and Moses took the blood, and with his finger put it on the horns of the altar around it and purified the altar and poured out the blood at the base of the altar and consecrated it to make atonement for it.
LEV|8|16|And he took all the fat that was on the entrails and the long lobe of the liver and the two kidneys with their fat, and Moses burned them on the altar.
LEV|8|17|But the bull and its skin and its flesh and its dung he burned up with fire outside the camp, as the LORD commanded Moses.
LEV|8|18|Then he presented the ram of the burnt offering, and Aaron and his sons laid their hands on the head of the ram.
LEV|8|19|And he killed it, and Moses threw the blood against the sides of the altar.
LEV|8|20|He cut the ram into pieces, and Moses burned the head and the pieces and the fat.
LEV|8|21|He washed the entrails and the legs with water, and Moses burned the whole ram on the altar. It was a burnt offering with a pleasing aroma, a food offering for the LORD, as the LORD commanded Moses.
LEV|8|22|Then he presented the other ram, the ram of ordination, and Aaron and his sons laid their hands on the head of the ram.
LEV|8|23|And he killed it, and Moses took some of its blood and put it on the lobe of Aaron's right ear and on the thumb of his right hand and on the big toe of his right foot.
LEV|8|24|Then he presented Aaron's sons, and Moses put some of the blood on the lobes of their right ears and on the thumbs of their right hands and on the big toes of their right feet. And Moses threw the blood against the sides of the altar.
LEV|8|25|Then he took the fat and the fat tail and all the fat that was on the entrails and the long lobe of the liver and the two kidneys with their fat and the right thigh,
LEV|8|26|and out of the basket of unleavened bread that was before the LORD he took one unleavened loaf and one loaf of bread with oil and one wafer and placed them on the pieces of fat and on the right thigh.
LEV|8|27|And he put all these in the hands of Aaron and in the hands of his sons and waved them as a wave offering before the LORD.
LEV|8|28|Then Moses took them from their hands and burned them on the altar with the burnt offering. This was an ordination offering with a pleasing aroma, a food offering to the LORD.
LEV|8|29|And Moses took the breast and waved it for a wave offering before the LORD. It was Moses' portion of the ram of ordination, as the LORD commanded Moses.
LEV|8|30|Then Moses took some of the anointing oil and of the blood that was on the altar and sprinkled it on Aaron and his garments, and also on his sons and his sons' garments. So he consecrated Aaron and his garments, and his sons and his sons' garments with him.
LEV|8|31|And Moses said to Aaron and his sons, "Boil the flesh at the entrance of the tent of meeting, and there eat it and the bread that is in the basket of ordination offerings, as I commanded, saying, 'Aaron and his sons shall eat it.'
LEV|8|32|And what remains of the flesh and the bread you shall burn up with fire.
LEV|8|33|And you shall not go outside the entrance of the tent of meeting for seven days, until the days of your ordination are completed, for it will take seven days to ordain you.
LEV|8|34|As has been done today, the LORD has commanded to be done to make atonement for you.
LEV|8|35|At the entrance of the tent of meeting you shall remain day and night for seven days, performing what the LORD has charged, so that you do not die, for so I have been commanded."
LEV|8|36|And Aaron and his sons did all the things that the LORD commanded by Moses.
LEV|9|1|On the eighth day Moses called Aaron and his sons and the elders of Israel,
LEV|9|2|and he said to Aaron, "Take for yourself a bull calf for a sin offering and a ram for a burnt offering, both without blemish, and offer them before the LORD.
LEV|9|3|And say to the people of Israel, 'Take a male goat for a sin offering, and a calf and a lamb, both a year old without blemish, for a burnt offering,
LEV|9|4|and an ox and a ram for peace offerings, to sacrifice before the LORD, and a grain offering mixed with oil, for today the LORD will appear to you.'"
LEV|9|5|And they brought what Moses commanded in front of the tent of meeting, and all the congregation drew near and stood before the LORD.
LEV|9|6|And Moses said, "This is the thing that the LORD commanded you to do, that the glory of the LORD may appear to you."
LEV|9|7|Then Moses said to Aaron, "Draw near to the altar and offer your sin offering and your burnt offering and make atonement for yourself and for the people, and bring the offering of the people and make atonement for them, as the LORD has commanded."
LEV|9|8|So Aaron drew near to the altar and killed the calf of the sin offering, which was for himself.
LEV|9|9|And the sons of Aaron presented the blood to him, and he dipped his finger in the blood and put it on the horns of the altar and poured out the blood at the base of the altar.
LEV|9|10|But the fat and the kidneys and the long lobe of the liver from the sin offering he burned on the altar, as the LORD commanded Moses.
LEV|9|11|The flesh and the skin he burned up with fire outside the camp.
LEV|9|12|Then he killed the burnt offering, and Aaron's sons handed him the blood, and he threw it against the sides of the altar.
LEV|9|13|And they handed the burnt offering to him, piece by piece, and the head, and he burned them on the altar.
LEV|9|14|And he washed the entrails and the legs and burned them with the burnt offering on the altar.
LEV|9|15|Then he presented the people's offering and took the goat of the sin offering that was for the people and killed it and offered it as a sin offering, like the first one.
LEV|9|16|And he presented the burnt offering and offered it according to the rule.
LEV|9|17|And he presented the grain offering, took a handful of it, and burned it on the altar, besides the burnt offering of the morning.
LEV|9|18|Then he killed the ox and the ram, the sacrifice of peace offerings for the people. And Aaron's sons handed him the blood, and he threw it against the sides of the altar.
LEV|9|19|But the fat pieces of the ox and of the ram, the fat tail and that which covers the entrails and the kidneys and the long lobe of the liver-
LEV|9|20|they put the fat pieces on the breasts, and he burned the fat pieces on the altar,
LEV|9|21|but the breasts and the right thigh Aaron waved for a wave offering before the LORD, as Moses commanded.
LEV|9|22|Then Aaron lifted up his hands toward the people and blessed them, and he came down from offering the sin offering and the burnt offering and the peace offerings.
LEV|9|23|And Moses and Aaron went into the tent of meeting, and when they came out they blessed the people, and the glory of the LORD appeared to all the people.
LEV|9|24|And fire came out from before the LORD and consumed the burnt offering and the pieces of fat on the altar, and when all the people saw it, they shouted and fell on their faces.
LEV|10|1|Now Nadab and Abihu, the sons of Aaron, each took his censer and put fire in it and laid incense on it and offered unauthorized fire before the LORD, which he had not commanded them.
LEV|10|2|And fire came out from before the LORD and consumed them, and they died before the LORD.
LEV|10|3|Then Moses said to Aaron, "This is what the LORD has said, 'Among those who are near me I will be sanctified, and before all the people I will be glorified.'"And Aaron held his peace.
LEV|10|4|And Moses called Mishael and Elzaphan, the sons of Uzziel the uncle of Aaron, and said to them, "Come near; carry your brothers away from the front of the sanctuary and out of the camp."
LEV|10|5|So they came near and carried them in their coats out of the camp, as Moses had said.
LEV|10|6|And Moses said to Aaron and to Eleazar and Ithamar his sons, "Do not let the hair of your heads hang loose, and do not tear your clothes, lest you die, and wrath come upon all the congregation; but let your brothers, the whole house of Israel, bewail the burning that the LORD has kindled.
LEV|10|7|And do not go outside the entrance of the tent of meeting, lest you die, for the anointing oil of the LORD is upon you." And they did according to the word of Moses.
LEV|10|8|And the LORD spoke to Aaron, saying,
LEV|10|9|"Drink no wine or strong drink, you or your sons with you, when you go into the tent of meeting, lest you die. It shall be a statute forever throughout your generations.
LEV|10|10|You are to distinguish between the holy and the common, and between the unclean and the clean,
LEV|10|11|and you are to teach the people of Israel all the statutes that the LORD has spoken to them by Moses."
LEV|10|12|Moses spoke to Aaron and to Eleazar and Ithamar, his surviving sons: "Take the grain offering that is left of the LORD's food offerings, and eat it unleavened beside the altar, for it is most holy.
LEV|10|13|You shall eat it in a holy place, because it is your due and your sons' due, from the LORD's food offerings, for so I am commanded.
LEV|10|14|But the breast that is waved and the thigh that is contributed you shall eat in a clean place, you and your sons and your daughters with you, for they are given as your due and your sons' due from the sacrifices of the peace offerings of the people of Israel.
LEV|10|15|The thigh that is contributed and the breast that is waved they shall bring with the food offerings of the fat pieces to wave for a wave offering before the LORD, and it shall be yours and your sons' with you as a due forever, as the LORD has commanded."
LEV|10|16|Now Moses diligently inquired about the goat of the sin offering, and behold, it was burned up! And he was angry with Eleazar and Ithamar, the surviving sons of Aaron, saying,
LEV|10|17|"Why have you not eaten the sin offering in the place of the sanctuary, since it is a thing most holy and has been given to you that you may bear the iniquity of the congregation, to make atonement for them before the LORD?
LEV|10|18|Behold, its blood was not brought into the inner part of the sanctuary. You certainly ought to have eaten it in the sanctuary, as I commanded."
LEV|10|19|And Aaron said to Moses, "Behold, today they have offered their sin offering and their burnt offering before the LORD, and yet such things as these have happened to me! If I had eaten the sin offering today, would the LORD have approved?"
LEV|10|20|And when Moses heard that, he approved.
LEV|11|1|And the LORD spoke to Moses and Aaron, saying to them,
LEV|11|2|"Speak to the people of Israel, saying, These are the living things that you may eat among all the animals that are on the earth.
LEV|11|3|Whatever parts the hoof and is cloven-footed and chews the cud, among the animals, you may eat.
LEV|11|4|Nevertheless, among those that chew the cud or part the hoof, you shall not eat these: The camel, because it chews the cud but does not part the hoof, is unclean to you.
LEV|11|5|And the rock badger, because it chews the cud but does not part the hoof, is unclean to you.
LEV|11|6|And the hare, because it chews the cud but does not part the hoof, is unclean to you.
LEV|11|7|And the pig, because it parts the hoof and is cloven-footed but does not chew the cud, is unclean to you.
LEV|11|8|You shall not eat any of their flesh, and you shall not touch their carcasses; they are unclean to you.
LEV|11|9|"These you may eat, of all that are in the waters. Everything in the waters that has fins and scales, whether in the seas or in the rivers, you may eat.
LEV|11|10|But anything in the seas or the rivers that has not fins and scales, of the swarming creatures in the waters and of the living creatures that are in the waters, is detestable to you.
LEV|11|11|You shall regard them as detestable; you shall not eat any of their flesh, and you shall detest their carcasses.
LEV|11|12|Everything in the waters that has not fins and scales is detestable to you.
LEV|11|13|"And these you shall detest among the birds; they shall not be eaten; they are detestable: the eagle, the bearded vulture, the black vulture,
LEV|11|14|the kite, the falcon of any kind,
LEV|11|15|every raven of any kind,
LEV|11|16|the ostrich, the nighthawk, the sea gull, the hawk of any kind,
LEV|11|17|the little owl, the cormorant, the short-eared owl,
LEV|11|18|the barn owl, the tawny owl, the carrion vulture,
LEV|11|19|the stork, the heron of any kind, the hoopoe, and the bat.
LEV|11|20|"All winged insects that go on all fours are detestable to you.
LEV|11|21|Yet among the winged insects that go on all fours you may eat those that have jointed legs above their feet, with which to hop on the ground.
LEV|11|22|Of them you may eat: the locust of any kind, the bald locust of any kind, the cricket of any kind, and the grasshopper of any kind.
LEV|11|23|But all other winged insects that have four feet are detestable to you.
LEV|11|24|"And by these you shall become unclean. Whoever touches their carcass shall be unclean until the evening,
LEV|11|25|and whoever carries any part of their carcass shall wash his clothes and be unclean until the evening.
LEV|11|26|Every animal that parts the hoof but is not cloven-footed or does not chew the cud is unclean to you. Everyone who touches them shall be unclean.
LEV|11|27|And all that walk on their paws, among the animals that go on all fours, are unclean to you. Whoever touches their carcass shall be unclean until the evening,
LEV|11|28|and he who carries their carcass shall wash his clothes and be unclean until the evening; they are unclean to you.
LEV|11|29|"And these are unclean to you among the swarming things that swarm on the ground: the mole rat, the mouse, the great lizard of any kind,
LEV|11|30|the gecko, the monitor lizard, the lizard, the sand lizard, and the chameleon.
LEV|11|31|These are unclean to you among all that swarm. Whoever touches them when they are dead shall be unclean until the evening.
LEV|11|32|And anything on which any of them falls when they are dead shall be unclean, whether it is an article of wood or a garment or a skin or a sack, any article that is used for any purpose. It must be put into water, and it shall be unclean until the evening; then it shall be clean.
LEV|11|33|And if any of them falls into any earthenware vessel, all that is in it shall be unclean, and you shall break it.
LEV|11|34|Any food in it that could be eaten, on which water comes, shall be unclean. And all drink that could be drunk from every such vessel shall be unclean.
LEV|11|35|And everything on which any part of their carcass falls shall be unclean. Whether oven or stove, it shall be broken in pieces. They are unclean and shall remain unclean for you.
LEV|11|36|Nevertheless, a spring or a cistern holding water shall be clean, but whoever touches a carcass in them shall be unclean.
LEV|11|37|And if any part of their carcass falls upon any seed grain that is to be sown, it is clean,
LEV|11|38|but if water is put on the seed and any part of their carcass falls on it, it is unclean to you.
LEV|11|39|"And if any animal which you may eat dies, whoever touches its carcass shall be unclean until the evening,
LEV|11|40|and whoever eats of its carcass shall wash his clothes and be unclean until the evening. And whoever carries the carcass shall wash his clothes and be unclean until the evening.
LEV|11|41|"Every swarming thing that swarms on the ground is detestable; it shall not be eaten.
LEV|11|42|Whatever goes on its belly, and whatever goes on all fours, or whatever has many feet, any swarming thing that swarms on the ground, you shall not eat, for they are detestable.
LEV|11|43|You shall not make yourselves detestable with any swarming thing that swarms, and you shall not defile yourselves with them, and become unclean through them.
LEV|11|44|For I am the LORD your God. Consecrate yourselves therefore, and be holy, for I am holy. You shall not defile yourselves with any swarming thing that crawls on the ground.
LEV|11|45|For I am the LORD who brought you up out of the land of Egypt to be your God. You shall therefore be holy, for I am holy."
LEV|11|46|This is the law about beast and bird and every living creature that moves through the waters and every creature that swarms on the ground,
LEV|11|47|to make a distinction between the unclean and the clean and between the living creature that may be eaten and the living creature that may not be eaten.
LEV|12|1|The LORD spoke to Moses, saying,
LEV|12|2|"Speak to the people of Israel, saying, 'If a woman conceives and bears a male child, then she shall be unclean seven days. As at the time of her menstruation, she shall be unclean.
LEV|12|3|And on the eighth day the flesh of his foreskin shall be circumcised.
LEV|12|4|Then she shall continue for thirty-three days in the blood of her purifying. She shall not touch anything holy, nor come into the sanctuary, until the days of her purifying are completed.
LEV|12|5|But if she bears a female child, then she shall be unclean two weeks, as in her menstruation. And she shall continue in the blood of her purifying for sixty-six days.
LEV|12|6|"'And when the days of her purifying are completed, whether for a son or for a daughter, she shall bring to the priest at the entrance of the tent of meeting a lamb a year old for a burnt offering, and a pigeon or a turtledove for a sin offering,
LEV|12|7|and he shall offer it before the LORD and make atonement for her. Then she shall be clean from the flow of her blood. This is the law for her who bears a child, either male or female.
LEV|12|8|And if she cannot afford a lamb, then she shall take two turtledoves or two pigeons, one for a burnt offering and the other for a sin offering. And the priest shall make atonement for her, and she shall be clean.'"
LEV|13|1|The LORD spoke to Moses and Aaron, saying,
LEV|13|2|"When a person has on the skin of his body a swelling or an eruption or a spot, and it turns into a case of leprous disease on the skin of his body, then he shall be brought to Aaron the priest or to one of his sons the priests,
LEV|13|3|and the priest shall examine the diseased area on the skin of his body. And if the hair in the diseased area has turned white and the disease appears to be deeper than the skin of his body, it is a case of leprous disease. When the priest has examined him, he shall pronounce him unclean.
LEV|13|4|But if the spot is white in the skin of his body and appears no deeper than the skin, and the hair in it has not turned white, the priest shall shut up the diseased person for seven days.
LEV|13|5|And the priest shall examine him on the seventh day, and if in his eyes the disease is checked and the disease has not spread in the skin, then the priest shall shut him up for another seven days.
LEV|13|6|And the priest shall examine him again on the seventh day, and if the diseased area has faded and the disease has not spread in the skin, then the priest shall pronounce him clean; it is only an eruption. And he shall wash his clothes and be clean.
LEV|13|7|But if the eruption spreads in the skin, after he has shown himself to the priest for his cleansing, he shall appear again before the priest.
LEV|13|8|And the priest shall look, and if the eruption has spread in the skin, then the priest shall pronounce him unclean; it is a leprous disease.
LEV|13|9|"When a man is afflicted with a leprous disease, he shall be brought to the priest,
LEV|13|10|and the priest shall look. And if there is a white swelling in the skin that has turned the hair white, and there is raw flesh in the swelling,
LEV|13|11|it is a chronic leprous disease in the skin of his body, and the priest shall pronounce him unclean. He shall not shut him up, for he is unclean.
LEV|13|12|And if the leprous disease breaks out in the skin, so that the leprous disease covers all the skin of the diseased person from head to foot, so far as the priest can see,
LEV|13|13|then the priest shall look, and if the leprous disease has covered all his body, he shall pronounce him clean of the disease; it has all turned white, and he is clean.
LEV|13|14|But when raw flesh appears on him, he shall be unclean.
LEV|13|15|And the priest shall examine the raw flesh and pronounce him unclean. Raw flesh is unclean, for it is a leprous disease.
LEV|13|16|But if the raw flesh recovers and turns white again, then he shall come to the priest,
LEV|13|17|and the priest shall examine him, and if the disease has turned white, then the priest shall pronounce the diseased person clean; he is clean.
LEV|13|18|"If there is in the skin of one's body a boil and it heals,
LEV|13|19|and in the place of the boil there comes a white swelling or a reddish-white spot, then it shall be shown to the priest.
LEV|13|20|And the priest shall look, and if it appears deeper than the skin and its hair has turned white, then the priest shall pronounce him unclean. It is a case of leprous disease that has broken out in the boil.
LEV|13|21|But if the priest examines it and there is no white hair in it and it is not deeper than the skin, but has faded, then the priest shall shut him up seven days.
LEV|13|22|And if it spreads in the skin, then the priest shall pronounce him unclean; it is a disease.
LEV|13|23|But if the spot remains in one place and does not spread, it is the scar of the boil, and the priest shall pronounce him clean.
LEV|13|24|"Or, when the body has a burn on its skin and the raw flesh of the burn becomes a spot, reddish-white or white,
LEV|13|25|the priest shall examine it, and if the hair in the spot has turned white and it appears deeper than the skin, then it is a leprous disease. It has broken out in the burn, and the priest shall pronounce him unclean; it is a case of leprous disease.
LEV|13|26|But if the priest examines it and there is no white hair in the spot and it is no deeper than the skin, but has faded, the priest shall shut him up seven days,
LEV|13|27|and the priest shall examine him the seventh day. If it is spreading in the skin, then the priest shall pronounce him unclean; it is a case of leprous disease.
LEV|13|28|But if the spot remains in one place and does not spread in the skin, but has faded, it is a swelling from the burn, and the priest shall pronounce him clean, for it is the scar of the burn.
LEV|13|29|"When a man or woman has a disease on the head or the beard,
LEV|13|30|the priest shall examine the disease. And if it appears deeper than the skin, and the hair in it is yellow and thin, then the priest shall pronounce him unclean. It is an itch, a leprous disease of the head or the beard.
LEV|13|31|And if the priest examines the itching disease and it appears no deeper than the skin and there is no black hair in it, then the priest shall shut up the person with the itching disease for seven days,
LEV|13|32|and on the seventh day the priest shall examine the disease. If the itch has not spread, and there is in it no yellow hair, and the itch appears to be no deeper than the skin,
LEV|13|33|then he shall shave himself, but the itch he shall not shave; and the priest shall shut up the person with the itching disease for another seven days.
LEV|13|34|And on the seventh day the priest shall examine the itch, and if the itch has not spread in the skin and it appears to be no deeper than the skin, then the priest shall pronounce him clean. And he shall wash his clothes and be clean.
LEV|13|35|But if the itch spreads in the skin after his cleansing,
LEV|13|36|then the priest shall examine him, and if the itch has spread in the skin, the priest need not seek for the yellow hair; he is unclean.
LEV|13|37|But if in his eyes the itch is unchanged and black hair has grown in it, the itch is healed and he is clean, and the priest shall pronounce him clean.
LEV|13|38|"When a man or a woman has spots on the skin of the body, white spots,
LEV|13|39|the priest shall look, and if the spots on the skin of the body are of a dull white, it is leukoderma that has broken out in the skin; he is clean.
LEV|13|40|"If a man's hair falls out from his head, he is bald; he is clean.
LEV|13|41|And if a man's hair falls out from his forehead, he has baldness of the forehead; he is clean.
LEV|13|42|But if there is on the bald head or the bald forehead a reddish-white diseased area, it is a leprous disease breaking out on his bald head or his bald forehead.
LEV|13|43|Then the priest shall examine him, and if the diseased swelling is reddish-white on his bald head or on his bald forehead, like the appearance of leprous disease in the skin of the body,
LEV|13|44|he is a leprous man, he is unclean. The priest must pronounce him unclean; his disease is on his head.
LEV|13|45|"The leprous person who has the disease shall wear torn clothes and let the hair of his head hang loose, and he shall cover his upper lip and cry out, 'Unclean, unclean.'
LEV|13|46|He shall remain unclean as long as he has the disease. He is unclean. He shall live alone. His dwelling shall be outside the camp.
LEV|13|47|"When there is a case of leprous disease in a garment, whether a woolen or a linen garment,
LEV|13|48|in warp or woof of linen or wool, or in a skin or in anything made of skin,
LEV|13|49|if the disease is greenish or reddish in the garment, or in the skin or in the warp or the woof or in any article made of skin, it is a case of leprous disease, and it shall be shown to the priest.
LEV|13|50|And the priest shall examine the disease and shut up that which has the disease for seven days.
LEV|13|51|Then he shall examine the disease on the seventh day. If the disease has spread in the garment, in the warp or the woof, or in the skin, whatever be the use of the skin, the disease is a persistent leprous disease; it is unclean.
LEV|13|52|And he shall burn the garment, or the warp or the woof, the wool or the linen, or any article made of skin that is diseased, for it is a persistent leprous disease. It shall be burned in the fire.
LEV|13|53|"And if the priest examines, and if the disease has not spread in the garment, in the warp or the woof or in any article made of skin,
LEV|13|54|then the priest shall command that they wash the thing in which is the disease, and he shall shut it up for another seven days.
LEV|13|55|And the priest shall examine the diseased thing after it has been washed. And if the appearance of the diseased area has not changed, though the disease has not spread, it is unclean. You shall burn it in the fire, whether the rot is on the back or on the front.
LEV|13|56|"But if the priest examines, and if the diseased area has faded after it has been washed, he shall tear it out of the garment or the skin or the warp or the woof.
LEV|13|57|Then if it appears again in the garment, in the warp or the woof, or in any article made of skin, it is spreading. You shall burn with fire whatever has the disease.
LEV|13|58|But the garment, or the warp or the woof, or any article made of skin from which the disease departs when you have washed it, shall then be washed a second time, and be clean."
LEV|13|59|This is the law for a case of leprous disease in a garment of wool or linen, either in the warp or the woof, or in any article made of skin, to determine whether it is clean or unclean.
LEV|14|1|The LORD spoke to Moses, saying,
LEV|14|2|"This shall be the law of the leprous person for the day of his cleansing. He shall be brought to the priest,
LEV|14|3|and the priest shall go out of the camp, and the priest shall look. Then, if the case of leprous disease is healed in the leprous person,
LEV|14|4|the priest shall command them to take for him who is to be cleansed two live clean birds and cedarwood and scarlet yarn and hyssop.
LEV|14|5|And the priest shall command them to kill one of the birds in an earthenware vessel over fresh water.
LEV|14|6|He shall take the live bird with the cedarwood and the scarlet yarn and the hyssop, and dip them and the live bird in the blood of the bird that was killed over the fresh water.
LEV|14|7|And he shall sprinkle it seven times on him who is to be cleansed of the leprous disease. Then he shall pronounce him clean and shall let the living bird go into the open field.
LEV|14|8|And he who is to be cleansed shall wash his clothes and shave off all his hair and bathe himself in water, and he shall be clean. And after that he may come into the camp, but live outside his tent seven days.
LEV|14|9|And on the seventh day he shall shave off all his hair from his head, his beard, and his eyebrows. He shall shave off all his hair, and then he shall wash his clothes and bathe his body in water, and he shall be clean.
LEV|14|10|"And on the eighth day he shall take two male lambs without blemish, and one ewe lamb a year old without blemish, and a grain offering of three tenths of an ephah of fine flour mixed with oil, and one log of oil.
LEV|14|11|And the priest who cleanses him shall set the man who is to be cleansed and these things before the LORD, at the entrance of the tent of meeting.
LEV|14|12|And the priest shall take one of the male lambs and offer it for a guilt offering, along with the log of oil, and wave them for a wave offering before the LORD.
LEV|14|13|And he shall kill the lamb in the place where they kill the sin offering and the burnt offering, in the place of the sanctuary. For the guilt offering, like the sin offering, belongs to the priest; it is most holy.
LEV|14|14|The priest shall take some of the blood of the guilt offering, and the priest shall put it on the lobe of the right ear of him who is to be cleansed and on the thumb of his right hand and on the big toe of his right foot.
LEV|14|15|Then the priest shall take some of the log of oil and pour it into the palm of his own left hand
LEV|14|16|and dip his right finger in the oil that is in his left hand and sprinkle some oil with his finger seven times before the LORD.
LEV|14|17|And some of the oil that remains in his hand the priest shall put on the lobe of the right ear of him who is to be cleansed and on the thumb of his right hand and on the big toe of his right foot, on top of the blood of the guilt offering.
LEV|14|18|And the rest of the oil that is in the priest's hand he shall put on the head of him who is to be cleansed. Then the priest shall make atonement for him before the LORD.
LEV|14|19|The priest shall offer the sin offering, to make atonement for him who is to be cleansed from his uncleanness. And afterward he shall kill the burnt offering.
LEV|14|20|And the priest shall offer the burnt offering and the grain offering on the altar. Thus the priest shall make atonement for him, and he shall be clean.
LEV|14|21|"But if he is poor and cannot afford so much, then he shall take one male lamb for a guilt offering to be waved, to make atonement for him, and a tenth of an ephah of fine flour mixed with oil for a grain offering, and a log of oil;
LEV|14|22|also two turtledoves or two pigeons, whichever he can afford. The one shall be a sin offering and the other a burnt offering.
LEV|14|23|And on the eighth day he shall bring them for his cleansing to the priest, to the entrance of the tent of meeting, before the LORD.
LEV|14|24|And the priest shall take the lamb of the guilt offering and the log of oil, and the priest shall wave them for a wave offering before the LORD.
LEV|14|25|And he shall kill the lamb of the guilt offering. And the priest shall take some of the blood of the guilt offering and put it on the lobe of the right ear of him who is to be cleansed, and on the thumb of his right hand and on the big toe of his right foot.
LEV|14|26|And the priest shall pour some of the oil into the palm of his own left hand,
LEV|14|27|and shall sprinkle with his right finger some of the oil that is in his left hand seven times before the LORD.
LEV|14|28|And the priest shall put some of the oil that is in his hand on the lobe of the right ear of him who is to be cleansed and on the thumb of his right hand and on the big toe of his right foot, in the place where the blood of the guilt offering was put.
LEV|14|29|And the rest of the oil that is in the priest's hand he shall put on the head of him who is to be cleansed, to make atonement for him before the LORD.
LEV|14|30|And he shall offer, of the turtledoves or pigeons, whichever he can afford,
LEV|14|31|one for a sin offering and the other for a burnt offering, along with a grain offering. And the priest shall make atonement before the LORD for him who is being cleansed.
LEV|14|32|This is the law for him in whom is a case of leprous disease, who cannot afford the offerings for his cleansing."
LEV|14|33|The LORD spoke to Moses and Aaron, saying,
LEV|14|34|"When you come into the land of Canaan, which I give you for a possession, and I put a case of leprous disease in a house in the land of your possession,
LEV|14|35|then he who owns the house shall come and tell the priest, 'There seems to me to be some case of disease in my house.'
LEV|14|36|Then the priest shall command that they empty the house before the priest goes to examine the disease, lest all that is in the house be declared unclean. And afterward the priest shall go in to see the house.
LEV|14|37|And he shall examine the disease. And if the disease is in the walls of the house with greenish or reddish spots, and if it appears to be deeper than the surface,
LEV|14|38|then the priest shall go out of the house to the door of the house and shut up the house seven days.
LEV|14|39|And the priest shall come again on the seventh day, and look. If the disease has spread in the walls of the house,
LEV|14|40|then the priest shall command that they take out the stones in which is the disease and throw them into an unclean place outside the city.
LEV|14|41|And he shall have the inside of the house scraped all around, and the plaster that they scrape off they shall pour out in an unclean place outside the city.
LEV|14|42|Then they shall take other stones and put them in the place of those stones, and he shall take other plaster and plaster the house.
LEV|14|43|"If the disease breaks out again in the house, after he has taken out the stones and scraped the house and plastered it,
LEV|14|44|then the priest shall go and look. And if the disease has spread in the house, it is a persistent leprous disease in the house; it is unclean.
LEV|14|45|And he shall break down the house, its stones and timber and all the plaster of the house, and he shall carry them out of the city to an unclean place.
LEV|14|46|Moreover, whoever enters the house while it is shut up shall be unclean until the evening,
LEV|14|47|and whoever sleeps in the house shall wash his clothes, and whoever eats in the house shall wash his clothes.
LEV|14|48|"But if the priest comes and looks, and if the disease has not spread in the house after the house was plastered, then the priest shall pronounce the house clean, for the disease is healed.
LEV|14|49|And for the cleansing of the house he shall take two small birds, with cedarwood and scarlet yarn and hyssop,
LEV|14|50|and shall kill one of the birds in an earthenware vessel over fresh water
LEV|14|51|and shall take the cedarwood and the hyssop and the scarlet yarn, along with the live bird, and dip them in the blood of the bird that was killed and in the fresh water and sprinkle the house seven times.
LEV|14|52|Thus he shall cleanse the house with the blood of the bird and with the fresh water and with the live bird and with the cedarwood and hyssop and scarlet yarn.
LEV|14|53|And he shall let the live bird go out of the city into the open country. So he shall make atonement for the house, and it shall be clean."
LEV|14|54|This is the law for any case of leprous disease: for an itch,
LEV|14|55|for leprous disease in a garment or in a house,
LEV|14|56|and for a swelling or an eruption or a spot,
LEV|14|57|to show when it is unclean and when it is clean. This is the law for leprous disease.
LEV|15|1|The LORD spoke to Moses and Aaron, saying,
LEV|15|2|"Speak to the people of Israel and say to them, When any man has a discharge from his body, his discharge is unclean.
LEV|15|3|And this is the law of his uncleanness for a discharge: whether his body runs with his discharge, or his body is blocked up by his discharge, it is his uncleanness.
LEV|15|4|Every bed on which the one with the discharge lies shall be unclean, and everything on which he sits shall be unclean.
LEV|15|5|And anyone who touches his bed shall wash his clothes and bathe himself in water and be unclean until the evening.
LEV|15|6|And whoever sits on anything on which the one with the discharge has sat shall wash his clothes and bathe himself in water and be unclean until the evening.
LEV|15|7|And whoever touches the body of the one with the discharge shall wash his clothes and bathe himself in water and be unclean until the evening.
LEV|15|8|And if the one with the discharge spits on someone who is clean, then he shall wash his clothes and bathe himself in water and be unclean until the evening.
LEV|15|9|And any saddle on which the one with the discharge rides shall be unclean.
LEV|15|10|And whoever touches anything that was under him shall be unclean until the evening. And whoever carries such things shall wash his clothes and bathe himself in water and be unclean until the evening.
LEV|15|11|Anyone whom the one with the discharge touches without having rinsed his hands in water shall wash his clothes and bathe himself in water and be unclean until the evening.
LEV|15|12|And an earthenware vessel that the one with the discharge touches shall be broken, and every vessel of wood shall be rinsed in water.
LEV|15|13|"And when the one with a discharge is cleansed of his discharge, then he shall count for himself seven days for his cleansing, and wash his clothes. And he shall bathe his body in fresh water and shall be clean.
LEV|15|14|And on the eighth day he shall take two turtledoves or two pigeons and come before the LORD to the entrance of the tent of meeting and give them to the priest.
LEV|15|15|And the priest shall use them, one for a sin offering and the other for a burnt offering. And the priest shall make atonement for him before the LORD for his discharge.
LEV|15|16|"If a man has an emission of semen, he shall bathe his whole body in water and be unclean until the evening.
LEV|15|17|And every garment and every skin on which the semen comes shall be washed with water and be unclean until the evening.
LEV|15|18|If a man lies with a woman and has an emission of semen, both of them shall bathe themselves in water and be unclean until the evening.
LEV|15|19|"When a woman has a discharge, and the discharge in her body is blood, she shall be in her menstrual impurity for seven days, and whoever touches her shall be unclean until the evening.
LEV|15|20|And everything on which she lies during her menstrual impurity shall be unclean. Everything also on which she sits shall be unclean.
LEV|15|21|And whoever touches her bed shall wash his clothes and bathe himself in water and be unclean until the evening.
LEV|15|22|And whoever touches anything on which she sits shall wash his clothes and bathe himself in water and be unclean until the evening.
LEV|15|23|Whether it is the bed or anything on which she sits, when he touches it he shall be unclean until the evening.
LEV|15|24|And if any man lies with her and her menstrual impurity comes upon him, he shall be unclean seven days, and every bed on which he lies shall be unclean.
LEV|15|25|"If a woman has a discharge of blood for many days, not at the time of her menstrual impurity, or if she has a discharge beyond the time of her impurity, all the days of the discharge she shall continue in uncleanness. As in the days of her impurity, she shall be unclean.
LEV|15|26|Every bed on which she lies, all the days of her discharge, shall be to her as the bed of her impurity. And everything on which she sits shall be unclean, as in the uncleanness of her menstrual impurity.
LEV|15|27|And whoever touches these things shall be unclean, and shall wash his clothes and bathe himself in water and be unclean until the evening.
LEV|15|28|But if she is cleansed of her discharge, she shall count for herself seven days, and after that she shall be clean.
LEV|15|29|And on the eighth day she shall take two turtledoves or two pigeons and bring them to the priest, to the entrance of the tent of meeting.
LEV|15|30|And the priest shall use one for a sin offering and the other for a burnt offering. And the priest shall make atonement for her before the LORD for her unclean discharge.
LEV|15|31|"Thus you shall keep the people of Israel separate from their uncleanness, lest they die in their uncleanness by defiling my tabernacle that is in their midst."
LEV|15|32|This is the law for him who has a discharge and for him who has an emission of semen, becoming unclean thereby;
LEV|15|33|also for her who is unwell with her menstrual impurity, that is, for anyone, male or female, who has a discharge, and for the man who lies with a woman who is unclean.
LEV|16|1|The LORD spoke to Moses after the death of the two sons of Aaron, when they drew near before the LORD and died,
LEV|16|2|and the LORD said to Moses, "Tell Aaron your brother not to come at any time into the Holy Place inside the veil, before the mercy seat that is on the ark, so that he may not die. For I will appear in the cloud over the mercy seat.
LEV|16|3|But in this way Aaron shall come into the Holy Place: with a bull from the herd for a sin offering and a ram for a burnt offering.
LEV|16|4|He shall put on the holy linen coat and shall have the linen undergarment on his body, and he shall tie the linen sash around his waist, and wear the linen turban; these are the holy garments. He shall bathe his body in water and then put them on.
LEV|16|5|And he shall take from the congregation of the people of Israel two male goats for a sin offering, and one ram for a burnt offering.
LEV|16|6|"Aaron shall offer the bull as a sin offering for himself and shall make atonement for himself and for his house.
LEV|16|7|Then he shall take the two goats and set them before the LORD at the entrance of the tent of meeting.
LEV|16|8|And Aaron shall cast lots over the two goats, one lot for the LORD and the other lot for Azazel.
LEV|16|9|And Aaron shall present the goat on which the lot fell for the LORD and use it as a sin offering,
LEV|16|10|but the goat on which the lot fell for Azazel shall be presented alive before the LORD to make atonement over it, that it may be sent away into the wilderness to Azazel.
LEV|16|11|"Aaron shall present the bull as a sin offering for himself, and shall make atonement for himself and for his house. He shall kill the bull as a sin offering for himself.
LEV|16|12|And he shall take a censer full of coals of fire from the altar before the LORD, and two handfuls of sweet incense beaten small, and he shall bring it inside the veil
LEV|16|13|and put the incense on the fire before the LORD, that the cloud of the incense may cover the mercy seat that is over the testimony, so that he does not die.
LEV|16|14|And he shall take some of the blood of the bull and sprinkle it with his finger on the front of the mercy seat on the east side, and in front of the mercy seat he shall sprinkle some of the blood with his finger seven times.
LEV|16|15|"Then he shall kill the goat of the sin offering that is for the people and bring its blood inside the veil and do with its blood as he did with the blood of the bull, sprinkling it over the mercy seat and in front of the mercy seat.
LEV|16|16|Thus he shall make atonement for the Holy Place, because of the uncleannesses of the people of Israel and because of their transgressions, all their sins. And so he shall do for the tent of meeting, which dwells with them in the midst of their uncleannesses.
LEV|16|17|No one may be in the tent of meeting from the time he enters to make atonement in the Holy Place until he comes out and has made atonement for himself and for his house and for all the assembly of Israel.
LEV|16|18|Then he shall go out to the altar that is before the LORD and make atonement for it, and shall take some of the blood of the bull and some of the blood of the goat, and put it on the horns of the altar all around.
LEV|16|19|And he shall sprinkle some of the blood on it with his finger seven times, and cleanse it and consecrate it from the uncleannesses of the people of Israel.
LEV|16|20|"And when he has made an end of atoning for the Holy Place and the tent of meeting and the altar, he shall present the live goat.
LEV|16|21|And Aaron shall lay both his hands on the head of the live goat, and confess over it all the iniquities of the people of Israel, and all their transgressions, all their sins. And he shall put them on the head of the goat and send it away into the wilderness by the hand of a man who is in readiness.
LEV|16|22|The goat shall bear all their iniquities on itself to a remote area, and he shall let the goat go free in the wilderness.
LEV|16|23|"Then Aaron shall come into the tent of meeting and shall take off the linen garments that he put on when he went into the Holy Place and shall leave them there.
LEV|16|24|And he shall bathe his body in water in a holy place and put on his garments and come out and offer his burnt offering and the burnt offering of the people and make atonement for himself and for the people.
LEV|16|25|And the fat of the sin offering he shall burn on the altar.
LEV|16|26|And he who lets the goat go to Azazel shall wash his clothes and bathe his body in water, and afterward he may come into the camp.
LEV|16|27|And the bull for the sin offering and the goat for the sin offering, whose blood was brought in to make atonement in the Holy Place, shall be carried outside the camp. Their skin and their flesh and their dung shall be burned up with fire.
LEV|16|28|And he who burns them shall wash his clothes and bathe his body in water, and afterward he may come into the camp.
LEV|16|29|"And it shall be a statute to you forever that in the seventh month, on the tenth day of the month, you shall afflict yourselves and shall do no work, either the native or the stranger who sojourns among you.
LEV|16|30|For on this day shall atonement be made for you to cleanse you. You shall be clean before the LORD from all your sins.
LEV|16|31|It is a Sabbath of solemn rest to you, and you shall afflict yourselves; it is a statute forever.
LEV|16|32|And the priest who is anointed and consecrated as priest in his father's place shall make atonement, wearing the holy linen garments.
LEV|16|33|He shall make atonement for the holy sanctuary, and he shall make atonement for the tent of meeting and for the altar, and he shall make atonement for the priests and for all the people of the assembly.
LEV|16|34|And this shall be a statute forever for you, that atonement may be made for the people of Israel once in the year because of all their sins." And Moses did as the LORD commanded him.
LEV|17|1|And the LORD spoke to Moses, saying,
LEV|17|2|"Speak to Aaron and his sons and to all the people of Israel and say to them, This is the thing that the LORD has commanded.
LEV|17|3|If any one of the house of Israel kills an ox or a lamb or a goat in the camp, or kills it outside the camp,
LEV|17|4|and does not bring it to the entrance of the tent of meeting to offer it as a gift to the LORD in front of the tabernacle of the LORD, bloodguilt shall be imputed to that man. He has shed blood, and that man shall be cut off from among his people.
LEV|17|5|This is to the end that the people of Israel may bring their sacrifices that they sacrifice in the open field, that they may bring them to the LORD, to the priest at the entrance of the tent of meeting, and sacrifice them as sacrifices of peace offerings to the LORD.
LEV|17|6|And the priest shall throw the blood on the altar of the LORD at the entrance of the tent of meeting and burn the fat for a pleasing aroma to the LORD.
LEV|17|7|So they shall no more sacrifice their sacrifices to goat demons, after whom they whore. This shall be a statute forever for them throughout their generations.
LEV|17|8|"And you shall say to them, Any one of the house of Israel, or of the strangers who sojourn among them, who offers a burnt offering or sacrifice
LEV|17|9|and does not bring it to the entrance of the tent of meeting to offer it to the LORD, that man shall be cut off from his people.
LEV|17|10|"If any one of the house of Israel or of the strangers who sojourn among them eats any blood, I will set my face against that person who eats blood and will cut him off from among his people.
LEV|17|11|For the life of the flesh is in the blood, and I have given it for you on the altar to make atonement for your souls, for it is the blood that makes atonement by the life.
LEV|17|12|Therefore I have said to the people of Israel, No person among you shall eat blood, neither shall any stranger who sojourns among you eat blood.
LEV|17|13|"Any one also of the people of Israel, or of the strangers who sojourn among them, who takes in hunting any beast or bird that may be eaten shall pour out its blood and cover it with earth.
LEV|17|14|For the life of every creature is its blood: its blood is its life. Therefore I have said to the people of Israel, You shall not eat the blood of any creature, for the life of every creature is its blood. Whoever eats it shall be cut off.
LEV|17|15|And every person who eats what dies of itself or what is torn by beasts, whether he is a native or a sojourner, shall wash his clothes and bathe himself in water and be unclean until the evening; then he shall be clean.
LEV|17|16|But if he does not wash them or bathe his flesh, he shall bear his iniquity."
LEV|18|1|And the LORD spoke to Moses, saying,
LEV|18|2|"Speak to the people of Israel and say to them, I am the LORD your God.
LEV|18|3|You shall not do as they do in the land of Egypt, where you lived, and you shall not do as they do in the land of Canaan, to which I am bringing you. You shall not walk in their statutes.
LEV|18|4|You shall follow my rules and keep my statutes and walk in them. I am the LORD your God.
LEV|18|5|You shall therefore keep my statutes and my rules; if a person does them, he shall live by them: I am the LORD.
LEV|18|6|"None of you shall approach any one of his close relatives to uncover nakedness. I am the LORD.
LEV|18|7|You shall not uncover the nakedness of your father, which is the nakedness of your mother; she is your mother, you shall not uncover her nakedness.
LEV|18|8|You shall not uncover the nakedness of your father's wife; it is your father's nakedness.
LEV|18|9|You shall not uncover the nakedness of your sister, your father's daughter or your mother's daughter, whether brought up in the family or in another home.
LEV|18|10|You shall not uncover the nakedness of your son's daughter or of your daughter's daughter, for their nakedness is your own nakedness.
LEV|18|11|You shall not uncover the nakedness of your father's wife's daughter, brought up in your father's family, since she is your sister.
LEV|18|12|You shall not uncover the nakedness of your father's sister; she is your father's relative.
LEV|18|13|You shall not uncover the nakedness of your mother's sister, for she is your mother's relative.
LEV|18|14|You shall not uncover the nakedness of your father's brother, that is, you shall not approach his wife; she is your aunt.
LEV|18|15|You shall not uncover the nakedness of your daughter-in-law; she is your son's wife, you shall not uncover her nakedness.
LEV|18|16|You shall not uncover the nakedness of your brother's wife; it is your brother's nakedness.
LEV|18|17|You shall not uncover the nakedness of a woman and of her daughter, and you shall not take her son's daughter or her daughter's daughter to uncover her nakedness; they are relatives; it is depravity.
LEV|18|18|And you shall not take a woman as a rival wife to her sister, uncovering her nakedness while her sister is still alive.
LEV|18|19|"You shall not approach a woman to uncover her nakedness while she is in her menstrual uncleanness.
LEV|18|20|And you shall not lie sexually with your neighbor's wife and so make yourself unclean with her.
LEV|18|21|You shall not give any of your children to offer them to Molech, and so profane the name of your God: I am the LORD.
LEV|18|22|You shall not lie with a male as with a woman; it is an abomination.
LEV|18|23|And you shall not lie with any animal and so make yourself unclean with it, neither shall any woman give herself to an animal to lie with it: it is perversion.
LEV|18|24|"Do not make yourselves unclean by any of these things, for by all these the nations I am driving out before you have become unclean,
LEV|18|25|and the land became unclean, so that I punished its iniquity, and the land vomited out its inhabitants.
LEV|18|26|But you shall keep my statutes and my rules and do none of these abominations, either the native or the stranger who sojourns among you
LEV|18|27|(for the people of the land, who were before you, did all of these abominations, so that the land became unclean),
LEV|18|28|lest the land vomit you out when you make it unclean, as it vomited out the nation that was before you.
LEV|18|29|For everyone who does any of these abominations, the persons who do them shall be cut off from among their people.
LEV|18|30|So keep my charge never to practice any of these abominable customs that were practiced before you, and never to make yourselves unclean by them: I am the LORD your God."
LEV|19|1|And the LORD spoke to Moses, saying,
LEV|19|2|"Speak to all the congregation of the people of Israel and say to them, You shall be holy, for I the LORD your God am holy.
LEV|19|3|Every one of you shall revere his mother and his father, and you shall keep my Sabbaths: I am the LORD your God.
LEV|19|4|Do not turn to idols or make for yourselves any gods of cast metal: I am the LORD your God.
LEV|19|5|"When you offer a sacrifice of peace offerings to the LORD, you shall offer it so that you may be accepted.
LEV|19|6|It shall be eaten the same day you offer it or on the day after, and anything left over until the third day shall be burned up with fire.
LEV|19|7|If it is eaten at all on the third day, it is tainted; it will not be accepted,
LEV|19|8|and everyone who eats it shall bear his iniquity, because he has profaned what is holy to the LORD, and that person shall be cut off from his people.
LEV|19|9|"When you reap the harvest of your land, you shall not reap your field right up to its edge, neither shall you gather the gleanings after your harvest.
LEV|19|10|And you shall not strip your vineyard bare, neither shall you gather the fallen grapes of your vineyard. You shall leave them for the poor and for the sojourner: I am the LORD your God.
LEV|19|11|"You shall not steal; you shall not deal falsely; you shall not lie to one another.
LEV|19|12|You shall not swear by my name falsely, and so profane the name of your God: I am the LORD.
LEV|19|13|"You shall not oppress your neighbor or rob him. The wages of a hired servant shall not remain with you all night until the morning.
LEV|19|14|You shall not curse the deaf or put a stumbling block before the blind, but you shall fear your God: I am the LORD.
LEV|19|15|"You shall do no injustice in court. You shall not be partial to the poor or defer to the great, but in righteousness shall you judge your neighbor.
LEV|19|16|You shall not go around as a slanderer among your people, and you shall not stand up against the life of your neighbor: I am the LORD.
LEV|19|17|"You shall not hate your brother in your heart, but you shall reason frankly with your neighbor, lest you incur sin because of him.
LEV|19|18|You shall not take vengeance or bear a grudge against the sons of your own people, but you shall love your neighbor as yourself: I am the LORD.
LEV|19|19|"You shall keep my statutes. You shall not let your cattle breed with a different kind. You shall not sow your field with two kinds of seed, nor shall you wear a garment of cloth made of two kinds of material.
LEV|19|20|"If a man lies sexually with a woman who is a slave, assigned to another man and not yet ransomed or given her freedom, a distinction shall be made. They shall not be put to death, because she was not free;
LEV|19|21|but he shall bring his compensation to the LORD, to the entrance of the tent of meeting, a ram for a guilt offering.
LEV|19|22|And the priest shall make atonement for him with the ram of the guilt offering before the LORD for his sin that he has committed, and he shall be forgiven for the sin that he has committed.
LEV|19|23|"When you come into the land and plant any kind of tree for food, then you shall regard its fruit as forbidden. Three years it shall be forbidden to you; it must not be eaten.
LEV|19|24|And in the fourth year all its fruit shall be holy, an offering of praise to the LORD.
LEV|19|25|But in the fifth year you may eat of its fruit, to increase its yield for you: I am the LORD your God.
LEV|19|26|"You shall not eat any flesh with the blood in it. You shall not interpret omens or tell fortunes.
LEV|19|27|You shall not round off the hair on your temples or mar the edges of your beard.
LEV|19|28|You shall not make any cuts on your body for the dead or tattoo yourselves: I am the LORD.
LEV|19|29|"Do not profane your daughter by making her a prostitute, lest the land fall into prostitution and the land become full of depravity.
LEV|19|30|You shall keep my Sabbaths and reverence my sanctuary: I am the LORD.
LEV|19|31|"Do not turn to mediums or wizards; do not seek them out, and so make yourselves unclean by them: I am the LORD your God.
LEV|19|32|"You shall stand up before the gray head and honor the face of an old man, and you shall fear your God: I am the LORD.
LEV|19|33|"When a stranger sojourns with you in your land, you shall not do him wrong.
LEV|19|34|You shall treat the stranger who sojourns with you as the native among you, and you shall love him as yourself, for you were strangers in the land of Egypt: I am the LORD your God.
LEV|19|35|"You shall do no wrong in judgment, in measures of length or weight or quantity.
LEV|19|36|You shall have just balances, just weights, a just ephah, and a just hin: I am the LORD your God, who brought you out of the land of Egypt.
LEV|19|37|And you shall observe all my statutes and all my rules, and do them: I am the LORD."
LEV|20|1|The LORD spoke to Moses, saying,
LEV|20|2|"Say to the people of Israel, Any one of the people of Israel or of the strangers who sojourn in Israel who gives any of his children to Molech shall surely be put to death. The people of the land shall stone him with stones.
LEV|20|3|I myself will set my face against that man and will cut him off from among his people, because he has given one of his children to Molech, to make my sanctuary unclean and to profane my holy name.
LEV|20|4|And if the people of the land do at all close their eyes to that man when he gives one of his children to Molech, and do not put him to death,
LEV|20|5|then I will set my face against that man and against his clan and will cut them off from among their people, him and all who follow him in whoring after Molech.
LEV|20|6|"If a person turns to mediums and wizards, whoring after them, I will set my face against that person and will cut him off from among his people.
LEV|20|7|Consecrate yourselves, therefore, and be holy, for I am the LORD your God.
LEV|20|8|Keep my statutes and do them; I am the LORD who sanctifies you.
LEV|20|9|For anyone who curses his father or his mother shall surely be put to death; he has cursed his father or his mother; his blood is upon him.
LEV|20|10|"If a man commits adultery with the wife of his neighbor, both the adulterer and the adulteress shall surely be put to death.
LEV|20|11|If a man lies with his father's wife, he has uncovered his father's nakedness; both of them shall surely be put to death; their blood is upon them.
LEV|20|12|If a man lies with his daughter-in-law, both of them shall surely be put to death; they have committed perversion; their blood is upon them.
LEV|20|13|If a man lies with a male as with a woman, both of them have committed an abomination; they shall surely be put to death; their blood is upon them.
LEV|20|14|If a man takes a woman and her mother also, it is depravity; he and they shall be burned with fire, that there may be no depravity among you.
LEV|20|15|If a man lies with an animal, he shall surely be put to death, and you shall kill the animal.
LEV|20|16|If a woman approaches any animal and lies with it, you shall kill the woman and the animal; they shall surely be put to death; their blood is upon them.
LEV|20|17|"If a man takes his sister, a daughter of his father or a daughter of his mother, and sees her nakedness, and she sees his nakedness, it is a disgrace, and they shall be cut off in the sight of the children of their people. He has uncovered his sister's nakedness, and he shall bear his iniquity.
LEV|20|18|If a man lies with a woman during her menstrual period and uncovers her nakedness, he has made naked her fountain, and she has uncovered the fountain of her blood. Both of them shall be cut off from among their people.
LEV|20|19|You shall not uncover the nakedness of your mother's sister or of your father's sister, for that is to make naked one's relative; they shall bear their iniquity.
LEV|20|20|If a man lies with his uncle's wife, he has uncovered his uncle's nakedness; they shall bear their sin; they shall die childless.
LEV|20|21|If a man takes his brother's wife, it is impurity. He has uncovered his brother's nakedness; they shall be childless.
LEV|20|22|"You shall therefore keep all my statutes and all my rules and do them, that the land where I am bringing you to live may not vomit you out.
LEV|20|23|And you shall not walk in the customs of the nation that I am driving out before you, for they did all these things, and therefore I detested them.
LEV|20|24|But I have said to you, 'You shall inherit their land, and I will give it to you to possess, a land flowing with milk and honey.' I am the LORD your God, who have separated you from the peoples.
LEV|20|25|You shall therefore separate the clean beast from the unclean, and the unclean bird from the clean. You shall not make yourselves detestable by beast or by bird or by anything with which the ground crawls, which I have set apart for you to hold unclean.
LEV|20|26|You shall be holy to me, for I the LORD am holy and have separated you from the peoples, that you should be mine.
LEV|20|27|"A man or a woman who is a medium or a wizard shall surely be put to death. They shall be stoned with stones; their blood shall be upon them."
LEV|21|1|And the LORD said to Moses, "Speak to the priests, the sons of Aaron, and say to them: 'No one shall make himself unclean for the dead among his people,
LEV|21|2|except for his closest relatives, his mother, his father, his son, his daughter, his brother,
LEV|21|3|or his virgin sister (who is near to him because she has had no husband; for her he may make himself unclean).
LEV|21|4|He shall not make himself unclean as a husband among his people and so profane himself.
LEV|21|5|They shall not make bald patches on their heads, nor shave off the edges of their beards, nor make any cuts on their body.
LEV|21|6|They shall be holy to their God and not profane the name of their God. For they offer the LORD's food offerings, the bread of their God; therefore they shall be holy.
LEV|21|7|They shall not marry a prostitute or a woman who has been defiled, neither shall they marry a woman divorced from her husband, for the priest is holy to his God.
LEV|21|8|You shall sanctify him, for he offers the bread of your God. He shall be holy to you, for I, the LORD, who sanctify you, am holy.
LEV|21|9|And the daughter of any priest, if she profanes herself by whoring, profanes her father; she shall be burned with fire.
LEV|21|10|"The priest who is chief among his brothers, on whose head the anointing oil is poured and who has been consecrated to wear the garments, shall not let the hair of his head hang loose nor tear his clothes.
LEV|21|11|He shall not go in to any dead bodies nor make himself unclean, even for his father or for his mother.
LEV|21|12|He shall not go out of the sanctuary, lest he profane the sanctuary of his God, for the consecration of the anointing oil of his God is on him: I am the LORD.
LEV|21|13|And he shall take a wife in her virginity.
LEV|21|14|A widow, or a divorced woman, or a woman who has been defiled, or a prostitute, these he shall not marry. But he shall take as his wife a virgin of his own people,
LEV|21|15|that he may not profane his offspring among his people, for I am the LORD who sanctifies him."
LEV|21|16|And the LORD spoke to Moses, saying,
LEV|21|17|"Speak to Aaron, saying, None of your offspring throughout their generations who has a blemish may approach to offer the bread of his God.
LEV|21|18|For no one who has a blemish shall draw near, a man blind or lame, or one who has a mutilated face or a limb too long,
LEV|21|19|or a man who has an injured foot or an injured hand,
LEV|21|20|or a hunchback or a dwarf or a man with a defect in his sight or an itching disease or scabs or crushed testicles.
LEV|21|21|No man of the offspring of Aaron the priest who has a blemish shall come near to offer the LORD's food offerings; since he has a blemish, he shall not come near to offer the bread of his God.
LEV|21|22|He may eat the bread of his God, both of the most holy and of the holy things,
LEV|21|23|but he shall not go through the veil or approach the altar, because he has a blemish, that he may not profane my sanctuaries, for I am the LORD who sanctifies them."
LEV|21|24|So Moses spoke to Aaron and to his sons and to all the people of Israel.
LEV|22|1|And the LORD spoke to Moses, saying,
LEV|22|2|"Speak to Aaron and his sons so that they abstain from the holy things of the people of Israel, which they dedicate to me, so that they do not profane my holy name: I am the LORD.
LEV|22|3|Say to them, 'If any one of all your offspring throughout your generations approaches the holy things that the people of Israel dedicate to the LORD, while he has an uncleanness, that person shall be cut off from my presence: I am the LORD.
LEV|22|4|None of the offspring of Aaron who has a leprous disease or a discharge may eat of the holy things until he is clean. Whoever touches anything that is unclean through contact with the dead or a man who has had an emission of semen,
LEV|22|5|and whoever touches a swarming thing by which he may be made unclean or a person from whom he may take uncleanness, whatever his uncleanness may be-
LEV|22|6|the person who touches such a thing shall be unclean until the evening and shall not eat of the holy things unless he has bathed his body in water.
LEV|22|7|When the sun goes down he shall be clean, and afterward he may eat of the holy things, because they are his food.
LEV|22|8|He shall not eat what dies of itself or is torn by beasts, and so make himself unclean by it: I am the LORD.'
LEV|22|9|They shall therefore keep my charge, lest they bear sin for it and die thereby when they profane it: I am the LORD who sanctifies them.
LEV|22|10|"A lay person shall not eat of a holy thing; no foreign guest of the priest or hired servant shall eat of a holy thing,
LEV|22|11|but if a priest buys a slave as his property for money, the slave may eat of it, and anyone born in his house may eat of his food.
LEV|22|12|If a priest's daughter marries a layman, she shall not eat of the contribution of the holy things.
LEV|22|13|But if a priest's daughter is widowed or divorced and has no child and returns to her father's house, as in her youth, she may eat of her father's food; yet no lay person shall eat of it.
LEV|22|14|And if anyone eats of a holy thing unintentionally, he shall add the fifth of its value to it and give the holy thing to the priest.
LEV|22|15|They shall not profane the holy things of the people of Israel, which they contribute to the LORD,
LEV|22|16|and so cause them to bear iniquity and guilt, by eating their holy things: for I am the LORD who sanctifies them."
LEV|22|17|And the LORD spoke to Moses, saying,
LEV|22|18|"Speak to Aaron and his sons and all the people of Israel and say to them, When any one of the house of Israel or of the sojourners in Israel presents a burnt offering as his offering, for any of their vows or freewill offerings that they offer to the LORD,
LEV|22|19|if it is to be accepted for you it shall be a male without blemish, of the bulls or the sheep or the goats.
LEV|22|20|You shall not offer anything that has a blemish, for it will not be acceptable for you.
LEV|22|21|And when anyone offers a sacrifice of peace offerings to the LORD to fulfill a vow or as a freewill offering from the herd or from the flock, to be accepted it must be perfect; there shall be no blemish in it.
LEV|22|22|Animals blind or disabled or mutilated or having a discharge or an itch or scabs you shall not offer to the LORD or give them to the LORD as a food offering on the altar.
LEV|22|23|You may present a bull or a lamb that has a part too long or too short for a freewill offering, but for a vow offering it cannot be accepted.
LEV|22|24|Any animal that has its testicles bruised or crushed or torn or cut you shall not offer to the LORD; you shall not do it within your land,
LEV|22|25|neither shall you offer as the bread of your God any such animals gotten from a foreigner. Since there is a blemish in them, because of their mutilation, they will not be accepted for you."
LEV|22|26|And the LORD spoke to Moses, saying,
LEV|22|27|"When an ox or sheep or goat is born, it shall remain seven days with its mother, and from the eighth day on it shall be acceptable as a food offering to the LORD.
LEV|22|28|But you shall not kill an ox or a sheep and her young in one day.
LEV|22|29|And when you sacrifice a sacrifice of thanksgiving to the LORD, you shall sacrifice it so that you may be accepted.
LEV|22|30|It shall be eaten on the same day; you shall leave none of it until morning: I am the LORD.
LEV|22|31|"So you shall keep my commandments and do them: I am the LORD.
LEV|22|32|And you shall not profane my holy name, that I may be sanctified among the people of Israel. I am the LORD who sanctifies you,
LEV|22|33|who brought you out of the land of Egypt to be your God: I am the LORD."
LEV|23|1|The LORD spoke to Moses, saying,
LEV|23|2|"Speak to the people of Israel and say to them, These are the appointed feasts of the LORD that you shall proclaim as holy convocations; they are my appointed feasts.
LEV|23|3|"Six days shall work be done, but on the seventh day is a Sabbath of solemn rest, a holy convocation. You shall do no work. It is a Sabbath to the LORD in all your dwelling places.
LEV|23|4|"These are the appointed feasts of the LORD, the holy convocations, which you shall proclaim at the time appointed for them.
LEV|23|5|In the first month, on the fourteenth day of the month at twilight, is the LORD's Passover.
LEV|23|6|And on the fifteenth day of the same month is the Feast of Unleavened bread to the LORD; for seven days you shall eat unleavened bread.
LEV|23|7|On the first day you shall have a holy convocation; you shall not do any ordinary work.
LEV|23|8|But you shall present a food offering to the LORD for seven days. On the seventh day is a holy convocation; you shall not do any ordinary work."
LEV|23|9|And the LORD spoke to Moses, saying,
LEV|23|10|"Speak to the people of Israel and say to them, When you come into the land that I give you and reap its harvest, you shall bring the sheaf of the firstfruits of your harvest to the priest,
LEV|23|11|and he shall wave the sheaf before the LORD, so that you may be accepted. On the day after the Sabbath the priest shall wave it.
LEV|23|12|And on the day when you wave the sheaf, you shall offer a male lamb a year old without blemish as a burnt offering to the LORD.
LEV|23|13|And the grain offering with it shall be two tenths of an ephah of fine flour mixed with oil, a food offering to the LORD with a pleasing aroma, and the drink offering with it shall be of wine, a fourth of a hin.
LEV|23|14|And you shall eat neither bread nor grain parched or fresh until this same day, until you have brought the offering of your God: it is a statute forever throughout your generations in all your dwellings.
LEV|23|15|"You shall count seven full weeks from the day after the Sabbath, from the day that you brought the sheaf of the wave offering.
LEV|23|16|You shall count fifty days to the day after the seventh Sabbath. Then you shall present a grain offering of new grain to the LORD.
LEV|23|17|You shall bring from your dwelling places two loaves of bread to be waved, made of two tenths of an ephah. They shall be of fine flour, and they shall be baked with leaven, as firstfruits to the LORD.
LEV|23|18|And you shall present with the bread seven lambs a year old without blemish, and one bull from the herd and two rams. They shall be a burnt offering to the LORD, with their grain offering and their drink offerings, a food offering with a pleasing aroma to the LORD.
LEV|23|19|And you shall offer one male goat for a sin offering, and two male lambs a year old as a sacrifice of peace offerings.
LEV|23|20|And the priest shall wave them with the bread of the firstfruits as a wave offering before the LORD, with the two lambs. They shall be holy to the LORD for the priest.
LEV|23|21|And you shall make proclamation on the same day. You shall hold a holy convocation. You shall not do any ordinary work. It is a statute forever in all your dwelling places throughout your generations.
LEV|23|22|"And when you reap the harvest of your land, you shall not reap your field right up to its edge, nor shall you gather the gleanings after your harvest. You shall leave them for the poor and for the sojourner: I am the LORD your God."
LEV|23|23|And the LORD spoke to Moses, saying,
LEV|23|24|"Speak to the people of Israel, saying, In the seventh month, on the first day of the month, you shall observe a day of solemn rest, a memorial proclaimed with blast of trumpets, a holy convocation.
LEV|23|25|You shall not do any ordinary work, and you shall present a food offering to the LORD."
LEV|23|26|And the LORD spoke to Moses, saying,
LEV|23|27|"Now on the tenth day of this seventh month is the Day of Atonement. It shall be for you a time of holy convocation, and you shall afflict yourselves and present a food offering to the LORD.
LEV|23|28|And you shall not do any work on that very day, for it is a Day of Atonement, to make atonement for you before the LORD your God.
LEV|23|29|For whoever is not afflicted on that very day shall be cut off from his people.
LEV|23|30|And whoever does any work on that very day, that person I will destroy from among his people.
LEV|23|31|You shall not do any work. It is a statute forever throughout your generations in all your dwelling places.
LEV|23|32|It shall be to you a Sabbath of solemn rest, and you shall afflict yourselves. On the ninth day of the month beginning at evening, from evening to evening shall you keep your Sabbath."
LEV|23|33|And the LORD spoke to Moses, saying,
LEV|23|34|"Speak to the people of Israel, saying, On the fifteenth day of this seventh month and for seven days is the Feast of Booths to the LORD.
LEV|23|35|On the first day shall be a holy convocation; you shall not do any ordinary work.
LEV|23|36|For seven days you shall present food offerings to the LORD. On the eighth day you shall hold a holy convocation and present a food offering to the LORD. It is a solemn assembly; you shall not do any ordinary work.
LEV|23|37|"These are the appointed feasts of the LORD, which you shall proclaim as times of holy convocation, for presenting to the LORD food offerings, burnt offerings and grain offerings, sacrifices and drink offerings, each on its proper day,
LEV|23|38|besides the LORD's Sabbaths and besides your gifts and besides all your vow offerings and besides all your freewill offerings, which you give to the LORD.
LEV|23|39|"On the fifteenth day of the seventh month, when you have gathered in the produce of the land, you shall celebrate the feast of the LORD seven days. On the first day shall be a solemn rest, and on the eighth day shall be a solemn rest.
LEV|23|40|And you shall take on the first day the fruit of splendid trees, branches of palm trees and boughs of leafy trees and willows of the brook, and you shall rejoice before the LORD your God seven days.
LEV|23|41|You shall celebrate it as a feast to the LORD for seven days in the year. It is a statute forever throughout your generations; you shall celebrate it in the seventh month.
LEV|23|42|You shall dwell in booths for seven days. All native Israelites shall dwell in booths,
LEV|23|43|that your generations may know that I made the people of Israel dwell in booths when I brought them out of the land of Egypt: I am the LORD your God."
LEV|23|44|Thus Moses declared to the people of Israel the appointed feasts of the LORD.
LEV|24|1|The LORD spoke to Moses, saying,
LEV|24|2|"Command the people of Israel to bring you pure oil from beaten olives for the lamp, that a light may be kept burning regularly.
LEV|24|3|Outside the veil of the testimony, in the tent of meeting, Aaron shall arrange it from evening to morning before the LORD regularly. It shall be a statute forever throughout your generations.
LEV|24|4|He shall arrange the lamps on the lampstand of pure gold before the LORD regularly.
LEV|24|5|"You shall take fine flour and bake twelve loaves from it; two tenths of an ephah shall be in each loaf.
LEV|24|6|And you shall set them in two piles, six in a pile, on the table of pure gold before the LORD.
LEV|24|7|And you shall put pure frankincense on each pile, that it may go with the bread as a memorial portion as a food offering to the LORD.
LEV|24|8|Every Sabbath day Aaron shall arrange it before the LORD regularly; it is from the people of Israel as a covenant forever.
LEV|24|9|And it shall be for Aaron and his sons, and they shall eat it in a holy place, since it is for him a most holy portion out of the LORD's food offerings, a perpetual due."
LEV|24|10|Now an Israelite woman's son, whose father was an Egyptian, went out among the people of Israel. And the Israelite woman's son and a man of Israel fought in the camp,
LEV|24|11|and the Israelite woman's son blasphemed the Name, and cursed. Then they brought him to Moses. His mother's name was Shelomith, the daughter of Dibri, of the tribe of Dan.
LEV|24|12|And they put him in custody, till the will of the LORD should be clear to them.
LEV|24|13|Then the LORD spoke to Moses, saying,
LEV|24|14|"Bring out of the camp the one who cursed, and let all who heard him lay their hands on his head, and let all the congregation stone him.
LEV|24|15|And speak to the people of Israel, saying, Whoever curses his God shall bear his sin.
LEV|24|16|Whoever blasphemes the name of the LORD shall surely be put to death. All the congregation shall stone him. The sojourner as well as the native, when he blasphemes the Name, shall be put to death.
LEV|24|17|"Whoever takes a human life shall surely be put to death.
LEV|24|18|Whoever takes an animal's life shall make it good, life for life.
LEV|24|19|If anyone injures his neighbor, as he has done it shall be done to him,
LEV|24|20|fracture for fracture, eye for eye, tooth for tooth; whatever injury he has given a person shall be given to him.
LEV|24|21|Whoever kills an animal shall make it good, and whoever kills a person shall be put to death.
LEV|24|22|You shall have the same rule for the sojourner and for the native, for I am the LORD your God."
LEV|24|23|So Moses spoke to the people of Israel, and they brought out of the camp the one who had cursed and stoned him with stones. Thus the people of Israel did as the LORD commanded Moses.
LEV|25|1|The LORD spoke to Moses on Mount Sinai, saying,
LEV|25|2|"Speak to the people of Israel and say to them, When you come into the land that I give you, the land shall keep a Sabbath to the LORD.
LEV|25|3|For six years you shall sow your field, and for six years you shall prune your vineyard and gather in its fruits,
LEV|25|4|but in the seventh year there shall be a Sabbath of solemn rest for the land, a Sabbath to the LORD. You shall not sow your field or prune your vineyard.
LEV|25|5|You shall not reap what grows of itself in your harvest, or gather the grapes of your undressed vine. It shall be a year of solemn rest for the land.
LEV|25|6|The Sabbath of the land shall provide food for you, for yourself and for your male and female slaves and for your hired servant and the sojourner who lives with you,
LEV|25|7|and for your cattle and for the wild animals that are in your land: all its yield shall be for food.
LEV|25|8|"You shall count seven weeks of years, seven times seven years, so that the time of the seven weeks of years shall give you forty-nine years.
LEV|25|9|Then you shall sound the loud trumpet on the tenth day of the seventh month. On the Day of Atonement you shall sound the trumpet throughout all your land.
LEV|25|10|And you shall consecrate the fiftieth year, and proclaim liberty throughout the land to all its inhabitants. It shall be a jubilee for you, when each of you shall return to his property and each of you shall return to his clan.
LEV|25|11|That fiftieth year shall be a jubilee for you; in it you shall neither sow nor reap what grows of itself nor gather the grapes from the undressed vines.
LEV|25|12|For it is a jubilee. It shall be holy to you. You may eat the produce of the field.
LEV|25|13|"In this year of jubilee each of you shall return to his property.
LEV|25|14|And if you make a sale to your neighbor or buy from your neighbor, you shall not wrong one another.
LEV|25|15|You shall pay your neighbor according to the number of years after the jubilee, and he shall sell to you according to the number of years for crops.
LEV|25|16|If the years are many, you shall increase the price, and if the years are few, you shall reduce the price, for it is the number of the crops that he is selling to you.
LEV|25|17|You shall not wrong one another, but you shall fear your God, for I am the LORD your God.
LEV|25|18|"Therefore you shall do my statutes and keep my rules and perform them, and then you will dwell in the land securely.
LEV|25|19|The land will yield its fruit, and you will eat your fill and dwell in it securely.
LEV|25|20|And if you say, 'What shall we eat in the seventh year, if we may not sow or gather in our crop?'
LEV|25|21|I will command my blessing on you in the sixth year, so that it will produce a crop sufficient for three years.
LEV|25|22|When you sow in the eighth year, you will be eating some of the old crop; you shall eat the old until the ninth year, when its crop arrives.
LEV|25|23|"The land shall not be sold in perpetuity, for the land is mine. For you are strangers and sojourners with me.
LEV|25|24|And in all the country you possess, you shall allow a redemption of the land.
LEV|25|25|"If your brother becomes poor and sells part of his property, then his nearest redeemer shall come and redeem what his brother has sold.
LEV|25|26|If a man has no one to redeem it and then himself becomes prosperous and finds sufficient means to redeem it,
LEV|25|27|let him calculate the years since he sold it and pay back the balance to the man to whom he sold it, and then return to his property.
LEV|25|28|But if he has not sufficient means to recover it, then what he sold shall remain in the hand of the buyer until the year of jubilee. In the jubilee it shall be released, and he shall return to his property.
LEV|25|29|"If a man sells a dwelling house in a walled city, he may redeem it within a year of its sale. For a full year he shall have the right of redemption.
LEV|25|30|If it is not redeemed within a full year, then the house in the walled city shall belong in perpetuity to the buyer, throughout his generations; it shall not be released in the jubilee.
LEV|25|31|But the houses of the villages that have no wall around them shall be classified with the fields of the land. They may be redeemed, and they shall be released in the jubilee.
LEV|25|32|As for the cities of the Levites, the Levites may redeem at any time the houses in the cities they possess.
LEV|25|33|And if one of the Levites exercises his right of redemption, then the house that was sold in a city they possess shall be released in the jubilee. For the houses in the cities of the Levites are their possession among the people of Israel.
LEV|25|34|But the fields of pastureland belonging to their cities may not be sold, for that is their possession forever.
LEV|25|35|"If your brother becomes poor and cannot maintain himself with you, you shall support him as though he were a stranger and a sojourner, and he shall live with you.
LEV|25|36|Take no interest from him or profit, but fear your God, that your brother may live beside you.
LEV|25|37|You shall not lend him your money at interest, nor give him your food for profit.
LEV|25|38|I am the LORD your God, who brought you out of the land of Egypt to give you the land of Canaan, and to be your God.
LEV|25|39|"If your brother becomes poor beside you and sells himself to you, you shall not make him serve as a slave:
LEV|25|40|he shall be with you as a hired servant and as a sojourner. He shall serve with you until the year of the jubilee.
LEV|25|41|Then he shall go out from you, he and his children with him, and go back to his own clan and return to the possession of his fathers.
LEV|25|42|For they are my servants, whom I brought out of the land of Egypt; they shall not be sold as slaves.
LEV|25|43|You shall not rule over him ruthlessly but shall fear your God.
LEV|25|44|As for your male and female slaves whom you may have: you may buy male and female slaves from among the nations that are around you.
LEV|25|45|You may also buy from among the strangers who sojourn with you and their clans that are with you, who have been born in your land, and they may be your property.
LEV|25|46|You may bequeath them to your sons after you to inherit as a possession forever. You may make slaves of them, but over your brothers the people of Israel you shall not rule, one over another ruthlessly.
LEV|25|47|"If a stranger or sojourner with you becomes rich, and your brother beside him becomes poor and sells himself to the stranger or sojourner with you or to a member of the stranger's clan,
LEV|25|48|then after he is sold he may be redeemed. One of his brothers may redeem him,
LEV|25|49|or his uncle or his cousin may redeem him, or a close relative from his clan may redeem him. Or if he grows rich he may redeem himself.
LEV|25|50|He shall calculate with his buyer from the year when he sold himself to him until the year of jubilee, and the price of his sale shall vary with the number of years. The time he was with his owner shall be rated as the time of a hired servant.
LEV|25|51|If there are still many years left, he shall pay proportionately for his redemption some of his sale price.
LEV|25|52|If there remain but a few years until the year of jubilee, he shall calculate and pay for his redemption in proportion to his years of service.
LEV|25|53|He shall treat him as a servant hired year by year. He shall not rule ruthlessly over him in your sight.
LEV|25|54|And if he is not redeemed by these means, then he and his children with him shall be released in the year of jubilee.
LEV|25|55|For it is to me that the people of Israel are servants. They are my servants whom I brought out of the land of Egypt: I am the LORD your God.
LEV|26|1|"You shall not make idols for yourselves or erect an image or pillar, and you shall not set up a figured stone in your land to bow down to it, for I am the LORD your God.
LEV|26|2|You shall keep my Sabbaths and reverence my sanctuary: I am the LORD.
LEV|26|3|"If you walk in my statutes and observe my commandments and do them,
LEV|26|4|then I will give you your rains in their season, and the land shall yield its increase, and the trees of the field shall yield their fruit.
LEV|26|5|Your threshing shall last to the time of the grape harvest, and the grape harvest shall last to the time for sowing. And you shall eat your bread to the full and dwell in your land securely.
LEV|26|6|I will give peace in the land, and you shall lie down, and none shall make you afraid. And I will remove harmful beasts from the land, and the sword shall not go through your land.
LEV|26|7|You shall chase your enemies, and they shall fall before you by the sword.
LEV|26|8|Five of you shall chase a hundred, and a hundred of you shall chase ten thousand, and your enemies shall fall before you by the sword.
LEV|26|9|I will turn to you and make you fruitful and multiply you and will confirm my covenant with you.
LEV|26|10|You shall eat old store long kept, and you shall clear out the old to make way for the new.
LEV|26|11|I will make my dwelling among you, and my soul shall not abhor you.
LEV|26|12|And I will walk among you and will be your God, and you shall be my people.
LEV|26|13|I am the LORD your God, who brought you out of the land of Egypt, that you should not be their slaves. And I have broken the bars of your yoke and made you walk erect.
LEV|26|14|"But if you will not listen to me and will not do all these commandments,
LEV|26|15|if you spurn my statutes, and if your soul abhors my rules, so that you will not do all my commandments, but break my covenant,
LEV|26|16|then I will do this to you: I will visit you with panic, with wasting disease and fever that consume the eyes and make the heart ache. And you shall sow your seed in vain, for your enemies shall eat it.
LEV|26|17|I will set my face against you, and you shall be struck down before your enemies. Those who hate you shall rule over you, and you shall flee when none pursues you.
LEV|26|18|And if in spite of this you will not listen to me, then I will discipline you again sevenfold for your sins,
LEV|26|19|and I will break the pride of your power, and I will make your heavens like iron and your earth like bronze.
LEV|26|20|And your strength shall be spent in vain, for your land shall not yield its increase, and the trees of the land shall not yield their fruit.
LEV|26|21|"Then if you walk contrary to me and will not listen to me, I will continue striking you, sevenfold for your sins.
LEV|26|22|And I will let loose the wild beasts against you, which shall bereave you of your children and destroy your livestock and make you few in number, so that your roads shall be deserted.
LEV|26|23|"And if by this discipline you are not turned to me but walk contrary to me,
LEV|26|24|then I also will walk contrary to you, and I myself will strike you sevenfold for your sins.
LEV|26|25|And I will bring a sword upon you, that shall execute vengeance for the covenant. And if you gather within your cities, I will send pestilence among you, and you shall be delivered into the hand of the enemy.
LEV|26|26|When I break your supply of bread, ten women shall bake your bread in a single oven and shall dole out your bread again by weight, and you shall eat and not be satisfied.
LEV|26|27|"But if in spite of this you will not listen to me, but walk contrary to me,
LEV|26|28|then I will walk contrary to you in fury, and I myself will discipline you sevenfold for your sins.
LEV|26|29|You shall eat the flesh of your sons, and you shall eat the flesh of your daughters.
LEV|26|30|And I will destroy your high places and cut down your incense altars and cast your dead bodies upon the dead bodies of your idols, and my soul will abhor you.
LEV|26|31|And I will lay your cities waste and will make your sanctuaries desolate, and I will not smell your pleasing aromas.
LEV|26|32|And I myself will devastate the land, so that your enemies who settle in it shall be appalled at it.
LEV|26|33|And I will scatter you among the nations, and I will unsheathe the sword after you, and your land shall be a desolation, and your cities shall be a waste.
LEV|26|34|"Then the land shall enjoy its Sabbaths as long as it lies desolate, while you are in your enemies' land; then the land shall rest, and enjoy its Sabbaths.
LEV|26|35|As long as it lies desolate it shall have rest, the rest that it did not have on your Sabbaths when you were dwelling in it.
LEV|26|36|And as for those of you who are left, I will send faintness into their hearts in the lands of their enemies. The sound of a driven leaf shall put them to flight, and they shall flee as one flees from the sword, and they shall fall when none pursues.
LEV|26|37|They shall stumble over one another, as if to escape a sword, though none pursues. And you shall have no power to stand before your enemies.
LEV|26|38|And you shall perish among the nations, and the land of your enemies shall eat you up.
LEV|26|39|And those of you who are left shall rot away in your enemies' lands because of their iniquity, and also because of the iniquities of their fathers they shall rot away like them.
LEV|26|40|"But if they confess their iniquity and the iniquity of their fathers in their treachery that they committed against me, and also in walking contrary to me,
LEV|26|41|so that I walked contrary to them and brought them into the land of their enemies- if then their uncircumcised heart is humbled and they make amends for their iniquity,
LEV|26|42|then I will remember my covenant with Jacob, and I will remember my covenant with Isaac and my covenant with Abraham, and I will remember the land.
LEV|26|43|But the land shall be abandoned by them and enjoy its Sabbaths while it lies desolate without them, and they shall make amends for their iniquity, because they spurned my rules and their soul abhorred my statutes.
LEV|26|44|Yet for all that, when they are in the land of their enemies, I will not spurn them, neither will I abhor them so as to destroy them utterly and break my covenant with them, for I am the LORD their God.
LEV|26|45|But I will for their sake remember the covenant with their forefathers, whom I brought out of the land of Egypt in the sight of the nations, that I might be their God: I am the LORD."
LEV|26|46|These are the statutes and rules and laws that the LORD made between him and the people of Israel through Moses on Mount Sinai.
LEV|27|1|The LORD spoke to Moses, saying,
LEV|27|2|"Speak to the people of Israel and say to them, If anyone makes a special vow to the LORD involving the valuation of persons,
LEV|27|3|then the valuation of a male from twenty years old up to sixty years old shall be fifty shekels of silver, according to the shekel of the sanctuary.
LEV|27|4|If the person is a female, the valuation shall be thirty shekels.
LEV|27|5|If the person is from five years old up to twenty years old, the valuation shall be for a male twenty shekels, and for a female ten shekels.
LEV|27|6|If the person is from a month old up to five years old, the valuation shall be for a male five shekels of silver, and for a female the valuation shall be three shekels of silver.
LEV|27|7|And if the person is sixty years old or over, then the valuation for a male shall be fifteen shekels, and for a female ten shekels.
LEV|27|8|And if someone is too poor to pay the valuation, then he shall be made to stand before the priest, and the priest shall value him; the priest shall value him according to what the vower can afford.
LEV|27|9|"If the vow is an animal that may be offered as an offering to the LORD, all of it that he gives to the LORD is holy.
LEV|27|10|He shall not exchange it or make a substitute for it, good for bad, or bad for good; and if he does in fact substitute one animal for another, then both it and the substitute shall be holy.
LEV|27|11|And if it is any unclean animal that may not be offered as an offering to the LORD, then he shall stand the animal before the priest,
LEV|27|12|and the priest shall value it as either good or bad; as the priest values it, so it shall be.
LEV|27|13|But if he wishes to redeem it, he shall add a fifth to the valuation.
LEV|27|14|"When a man dedicates his house as a holy gift to the LORD, the priest shall value it as either good or bad; as the priest values it, so it shall stand.
LEV|27|15|And if the donor wishes to redeem his house, he shall add a fifth to the valuation price, and it shall be his.
LEV|27|16|"If a man dedicates to the LORD part of the land that is his possession, then the valuation shall be in proportion to its seed. A homer of barley seed shall be valued at fifty shekels of silver.
LEV|27|17|If he dedicates his field from the year of jubilee, the valuation shall stand,
LEV|27|18|but if he dedicates his field after the jubilee, then the priest shall calculate the price according to the years that remain until the year of jubilee, and a deduction shall be made from the valuation.
LEV|27|19|And if he who dedicates the field wishes to redeem it, then he shall add a fifth to its valuation price, and it shall remain his.
LEV|27|20|But if he does not wish to redeem the field, or if he has sold the field to another man, it shall not be redeemed anymore.
LEV|27|21|But the field, when it is released in the jubilee, shall be a holy gift to the LORD, like a field that has been devoted. The priest shall be in possession of it.
LEV|27|22|If he dedicates to the LORD a field that he has bought, which is not a part of his possession,
LEV|27|23|then the priest shall calculate the amount of the valuation for it up to the year of jubilee, and the man shall give the valuation on that day as a holy gift to the LORD.
LEV|27|24|In the year of jubilee the field shall return to him from whom it was bought, to whom the land belongs as a possession.
LEV|27|25|Every valuation shall be according to the shekel of the sanctuary: twenty gerahs shall make a shekel.
LEV|27|26|"But a firstborn of animals, which as a firstborn belongs to the LORD, no man may dedicate; whether ox or sheep, it is the LORD's.
LEV|27|27|And if it is an unclean animal, then he shall buy it back at the valuation, and add a fifth to it; or, if it is not redeemed, it shall be sold at the valuation.
LEV|27|28|"But no devoted thing that a man devotes to the LORD, of anything that he has, whether man or beast, or of his inherited field, shall be sold or redeemed; every devoted thing is most holy to the LORD.
LEV|27|29|No one devoted, who is to be devoted for destruction from mankind, shall be ransomed; he shall surely be put to death.
LEV|27|30|"Every tithe of the land, whether of the seed of the land or of the fruit of the trees, is the LORD's; it is holy to the LORD.
LEV|27|31|If a man wishes to redeem some of his tithe, he shall add a fifth to it.
LEV|27|32|And every tithe of herds and flocks, every tenth animal of all that pass under the herdsman's staff, shall be holy to the LORD.
LEV|27|33|One shall not differentiate between good or bad, neither shall he make a substitute for it; and if he does substitute for it, then both it and the substitute shall be holy; it shall not be redeemed."
LEV|27|34|These are the commandments that the LORD commanded Moses for the people of Israel on Mount Sinai.
