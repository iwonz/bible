EZEK|1|1|在三十年四月初五，我在 迦巴魯河 邊被擄的人當中，那時天開了，我看見上帝的異象。
EZEK|1|2|正是 約雅斤 王被擄的第五年四月初五，
EZEK|1|3|在 迦勒底 人之地的 迦巴魯河 邊，耶和華的話特地臨到 布西 的兒子 以西結 祭司，耶和華的手按在他身上。
EZEK|1|4|我觀看，看哪，狂風從北方颳來，有一朵大雲閃爍著火，周圍有光輝，其中的火好像閃耀的金屬；
EZEK|1|5|又從其中顯出四個活物的形像。他們的形狀是這樣：有人的形像，
EZEK|1|6|各有四張臉，四個翅膀。
EZEK|1|7|他們的腿是直的，腳掌好像牛犢的蹄，燦爛如磨亮的銅。
EZEK|1|8|在四面的翅膀以下有人的手。這四個活物的臉和翅膀是這樣：
EZEK|1|9|翅膀彼此相接，行走時並不轉彎，各自往前直行。
EZEK|1|10|至於臉的形像：四個活物各有人的臉，右面有獅子的臉，左面有牛的臉，也有鷹的臉；
EZEK|1|11|這就是他們的臉 。他們的翅膀向上張開，各有兩個翅膀彼此相接，用另外兩個翅膀遮體。
EZEK|1|12|他們各自往前直行。靈往哪裏去，他們就往哪裏去，行走時並不轉彎。
EZEK|1|13|至於四活物的形像，就如燒著火炭的形狀，又如火把的形狀。有火在四活物中間來回移動，這火有光輝，從火中發出閃電。
EZEK|1|14|這些活物往來奔走，好像電光一閃。
EZEK|1|15|我觀看活物，看哪，有四張臉的活物旁邊各有一個輪子在地上。
EZEK|1|16|輪子的形狀結構 好像耀眼的水蒼玉。四輪都是一個樣式，形狀 結構好像輪中套輪。
EZEK|1|17|輪子行走的時候，向四方直行，行走時並不轉彎。
EZEK|1|18|至於輪圈，高而可畏；四個輪圈周圍佈滿眼睛。
EZEK|1|19|活物行走，輪子也在旁邊行走；活物離地上升，輪子也上升。
EZEK|1|20|靈往哪裏去，活物就往哪裏去；輪子在活物旁邊上升，因為活物的靈在輪中。
EZEK|1|21|活物行走，輪子也行走；活物站住，輪子也站住；活物離地上升，輪子也在旁邊上升，因為活物的靈在輪中。
EZEK|1|22|活物的頭上面有穹蒼的形像，像耀眼驚人的水晶，鋪張在活物的頭頂上。
EZEK|1|23|穹蒼之下，活物的翅膀伸直，彼此相對，每個活物用兩個翅膀遮住自己；每個活物用兩個翅膀遮住自己 ，就是自己的身體。
EZEK|1|24|活物行走的時候，我聽見翅膀的響聲，像大水的聲音，像全能者的聲音，又像軍隊鬧鬨的聲音。活物站住的時候，翅膀垂下。
EZEK|1|25|在他們頭上的穹蒼之上有聲音。他們站住的時候，翅膀垂下。
EZEK|1|26|在他們頭上的穹蒼之上有寶座的形像，彷彿藍寶石的樣子；寶座的形像上方有彷彿人的樣子的形像。
EZEK|1|27|我見他的腰以上有彷彿閃耀的金屬，周圍有彷彿火的形狀，又見他的腰以下有彷彿火的形狀，周圍也有光輝。
EZEK|1|28|下雨的日子，雲中彩虹的形狀怎樣，周圍光輝的形狀也是怎樣。 這就是耶和華榮耀形像的樣式，我一看見就臉伏於地。我又聽見一位說話者的聲音。
EZEK|2|1|他對我說：「人子啊，你站起來，我要和你說話。」
EZEK|2|2|他對我說話的時候，靈進入我裏面，使我站起來，我就聽見他對我說話。
EZEK|2|3|他對我說：「人子啊，我差你往悖逆我的國家， 以色列 人那裏去，他們是悖逆我的。他們和他們的祖先違背我，直到今日。
EZEK|2|4|這些人厚著臉皮，心裏剛硬。我差你到他們那裏去，你要對他們說：『主耶和華如此說。』
EZEK|2|5|他們是悖逆之家，他們或聽，或不聽，必知道在他們中間有了先知。
EZEK|2|6|你，人子啊，雖有荊棘和蒺藜在你那裏，你又住在蠍子中間，總不要怕他們，也不要怕他們的話；他們雖是悖逆之家，但你不要怕他們的話，也不要因他們的臉色驚惶。
EZEK|2|7|他們或聽，或不聽，你只管將我的話告訴他們；他們是極其悖逆的。
EZEK|2|8|「但是你，人子啊，要聽我對你說的話，不要像那悖逆之家一樣悖逆，要開口吃我所賜給你的。」
EZEK|2|9|我觀看，看哪，有一隻手向我伸來；看哪，手中有一書卷。
EZEK|2|10|他在我面前展開書卷，它內外都寫著字，上面所寫的有哀號、嘆息、悲痛的話。
EZEK|3|1|他對我說：「人子啊，要吃你所得到的，吃下這書卷；然後要去，對 以色列 家宣講。」
EZEK|3|2|於是我張開了口，他就使我吃這書卷。
EZEK|3|3|他對我說：「人子啊，要吃我所賜給你的這書卷，塞滿你的肚腹。」我就吃了，口中覺得其甜如蜜。
EZEK|3|4|他對我說：「人子啊，你要到 以色列 家那裏去，對他們傳講我的話。
EZEK|3|5|你奉差遣不是往那說話艱澀、言語難懂的民那裏，而是往 以色列 家去；
EZEK|3|6|你不是往那說話艱澀、言語難懂的許多民族那裏去，他們的話你不懂。然而，我若差你往他們那裏去，他們會聽從你。
EZEK|3|7|以色列 家卻不肯聽從你，因為他們不肯聽從我；原來 以色列 全家是額頭堅硬、心裏剛愎的人。
EZEK|3|8|看哪，我使你的臉堅硬，對抗他們的臉；使你的額頭堅硬，對抗他們的額頭。
EZEK|3|9|我使你的額頭像金剛石，比火石更堅硬。他們雖是悖逆之家，但你不要怕他們，也不要因他們的臉色而驚惶。」
EZEK|3|10|他又對我說：「人子啊，我對你說的一切話，你心裏要領會，耳朵要聽。
EZEK|3|11|要到被擄的人，到你本國百姓那裏去，他們或聽，或不聽，你要對他們宣講，告訴他們這是主耶和華說的。」
EZEK|3|12|那時，靈將我舉起，我就聽見在我身後有極大震動的聲音：「耶和華的榮耀，從他所在之處，是應當稱頌的！」
EZEK|3|13|有活物的翅膀相碰的聲音，也有活物旁邊輪子的聲音，是極大震動的聲音。
EZEK|3|14|於是靈將我舉起，帶著我走。我就去了，十分苦惱，我的靈火熱；耶和華的手重重地按在我身上。
EZEK|3|15|我就來到 提勒‧亞畢 那些住在 迦巴魯河 邊被擄的人那裏，到他們住的地方 ，在他們中間驚愕地坐了七日。
EZEK|3|16|過了七日，耶和華的話臨到我，說：
EZEK|3|17|「人子啊，我立你作 以色列 家的守望者，所以你要聽我口中的話，替我警戒他們。
EZEK|3|18|我何時指著惡人說：『他必要死』；你若不警戒他，也不勸告他，使他離開惡行，拯救他的性命，這惡人必死在罪孽之中；我卻要從你手裏討他的血債。
EZEK|3|19|倘若你警戒惡人，他仍不轉離罪惡，也不離開惡行，他必死在罪孽之中，你卻救了自己的命。
EZEK|3|20|但是義人若轉離他的義而作惡，我要把絆腳石放在他面前，他必死亡；因你沒有警戒他，他必死在罪中，他素來所行的義不被記念；我卻要從你手裏討他的血債。
EZEK|3|21|倘若你警戒義人，使他不犯罪，他就不犯罪；他因領受警戒就必存活，你也救了自己的命。」
EZEK|3|22|在那裏耶和華的手按在我身上。他對我說：「起來，到平原去，我要在那裏和你說話。」
EZEK|3|23|於是我起來，到平原去，看哪，耶和華的榮耀停在那裏，正如我在 迦巴魯河 邊所見到的一樣，我就臉伏於地。
EZEK|3|24|靈進入我裏面，使我站起來。耶和華對我說：「你進屋裏去，把門關上。
EZEK|3|25|你，人子，看哪，人要用繩索捆綁你，使你不能出去到他們中間。
EZEK|3|26|我必使你的舌頭貼住上膛，以致你啞口，不能作責備他們的人；他們原是悖逆之家。
EZEK|3|27|但我對你說話的時候，必使你開口，你就要對他們說：『主耶和華如此說。』聽的，讓他聽；不聽的，任他不聽，因為他們是悖逆之家。」
EZEK|4|1|「你，人子啊，拿一塊磚，擺在你面前，將一座城 耶路撒冷 畫在上面。
EZEK|4|2|你要圍攻這城，築堡壘，建土堆，安營攻擊，周圍設撞城槌攻城，
EZEK|4|3|又要拿一個鐵盤放在你和城的中間，作為鐵牆。你要把你的臉對著這城，使城被困。你要圍攻這城，這要成為 以色列 家的預兆。
EZEK|4|4|「你要向左側臥，承擔 以色列 家的罪孽；按你向左側臥的日數，擔當他們的罪孽。
EZEK|4|5|我已將他們作惡的年數定了日期，就是三百九十天，你要如此擔當 以色列 家的罪孽。
EZEK|4|6|這些日子結束之後，你還要向右側臥，擔當 猶大 家的罪孽。我為你定了四十天，一天頂一年。
EZEK|4|7|你要把你的臉對著被困的 耶路撒冷 ，露出膀臂，說預言攻擊這城。
EZEK|4|8|看哪，我用繩索捆綁你，使你不能從這邊翻到那邊，直等到你圍困的日子結束。
EZEK|4|9|「你要取小麥、大麥、豆子、紅豆、小米、粗麥，裝在一個器皿裏，為自己做餅；在你側臥的三百九十天吃這餅。
EZEK|4|10|你所吃食物的量是每天二十舍客勒，要按時吃。
EZEK|4|11|你喝水的量是每天六分之一欣，要按時喝。
EZEK|4|12|你要吃這餅像大麥餅一樣，在眾人眼前用人的糞烤它。」
EZEK|4|13|耶和華說：「 以色列 人在我趕他們到的列國中，也必這樣吃不潔淨的食物。」
EZEK|4|14|我說：「唉！主耶和華，看哪，我從來未曾被玷污，從幼年到如今沒有吃過自然死的，或被野獸撕裂的，那不潔淨的肉也未曾入我的口。」
EZEK|4|15|於是他對我說：「看，我給你牛糞代替人糞，你要在上面烤你的餅。」
EZEK|4|16|他又對我說：「人子，看哪，我必斷絕 耶路撒冷 糧食的供應 。他們要帶著憂慮限量吃餅；帶著驚惶限量喝水。
EZEK|4|17|他們因缺糧缺水，彼此驚惶，在自己的罪孽中消滅。」
EZEK|5|1|「你，人子啊，拿一把快刀當作剃刀，用這刀剃你的頭髮和鬍鬚，然後用天平將鬚髮分成幾份。
EZEK|5|2|圍困的日子滿了，你要把三分之一放在城中用火焚燒；三分之一放在城的四圍用刀砍碎；三分之一任風吹散，我要拔刀追趕它們。
EZEK|5|3|你要從其中取幾根鬚髮，用衣服的邊包起來，
EZEK|5|4|再從其中取一些扔在火裏，在火中焚燒；必有火從其中出來燒盡 以色列 全家。
EZEK|5|5|主耶和華如此說：這就是 耶路撒冷 。我曾將它安置在列國中，列邦都在它的四圍。
EZEK|5|6|耶路撒冷 行惡，違背我的典章，過於列國；干犯我的律例，過於四圍的列邦。它棄絕我的典章，也沒有遵行我的律例。
EZEK|5|7|所以主耶和華如此說：因為你們混亂，過於四圍的列國，不遵行我的律例，不順從我的典章，甚至也不順從四圍列國的規條 ，
EZEK|5|8|所以主耶和華如此說：看哪，我，我必與你為敵，必在列國眼前，在你中間施行審判；
EZEK|5|9|並且因你一切可憎的事，我要在你中間行未曾行過，將來也不會行的事。
EZEK|5|10|在你中間，父親要吃兒子，兒子要吃父親。我必向你施行審判，將你剩下的人分散四方 。
EZEK|5|11|主耶和華說：我指著我的永生起誓，因你用一切可憎之物、可厭的事玷污我的聖所，所以，我要把你剃光 ，我的眼必不顧惜你，也不可憐你。
EZEK|5|12|你的百姓三分之一必遭瘟疫而死，因饑荒在你們中間而消滅；三分之一必在你四圍倒在刀下；我必將三分之一分散四方，要拔刀追趕他們。
EZEK|5|13|「我要這樣發盡我的怒氣；我向他們發的憤怒停止以後，自己就得到平息。當我向他們發盡我的憤怒時，他們就知道我─耶和華所說的是出於妒忌。
EZEK|5|14|在四圍的列國中，我要使你成為荒涼，在所有過路人的眼前看為羞辱。
EZEK|5|15|這樣，我必以怒氣、憤怒和烈怒的責備，向你施行審判。那時，它 就在四圍的列國中成為羞辱、譏刺、警戒、驚駭；這是我─耶和華說的。
EZEK|5|16|我向滅亡的人射出饑荒的惡箭，將它們射出，毀滅你們；那時，我要加重你們的饑荒，斷絕你們糧食的供應。
EZEK|5|17|我要令饑荒和惡獸臨到你，使你喪失兒女。瘟疫和流血的事必在你那裏盛行，我也要使刀劍臨到你。這是我─耶和華說的。」
EZEK|6|1|耶和華的話臨到我，說：
EZEK|6|2|「人子啊，你要面向 以色列 的眾山說預言。
EZEK|6|3|你要說： 以色列 的眾山哪，要聽主耶和華的話。主耶和華對大山、小岡、水溝、山谷如此說：看哪，我要使刀劍臨到你們，也必毀壞你們的丘壇。
EZEK|6|4|你們的祭壇要荒廢，香壇必打碎。我要使你們當中被殺的人仆倒在你們的偶像面前，
EZEK|6|5|將 以色列 人的屍首放在他們的偶像面前，把你們的骸骨拋散在祭壇的四周圍。
EZEK|6|6|無論你們住在何處，城鎮要變為廢墟，丘壇也必毀壞，以至於你們的祭壇荒廢，被定罪 ，偶像打碎消除，香壇砍倒；你們所做的被塗去。
EZEK|6|7|被殺的人必仆倒在你們中間，你們就知道我是耶和華。
EZEK|6|8|「我必留下一些人，你們中有人得以在列國中脫離刀劍，分散在列邦。
EZEK|6|9|那些逃脫的人，必在被擄所到的各國中記得我，我心裏何等傷痛，因他們起淫心，離棄我，淫蕩的眼追隨偶像。他們因所做一切可憎的惡事，必厭惡自己。
EZEK|6|10|他們必知道我是耶和華；我說過要使這災禍臨到他們身上，並非空話。
EZEK|6|11|「主耶和華如此說：你當擊掌頓足，說：哀哉！ 以色列 家做了這一切可憎的惡事，必仆倒在刀劍、饑荒、瘟疫之下。
EZEK|6|12|在遠方的，必遭瘟疫而死；在近處的，必倒在刀劍之下；那存留被圍困的，必因饑荒而死；我要在他們身上發盡我的憤怒。
EZEK|6|13|被殺的要仆倒在祭壇四圍的偶像中，在各高岡、各山頂、各青翠的樹下，和各茂密的橡樹下，就是他們獻馨香的祭給一切偶像的地方。那時，他們就知道我是耶和華。
EZEK|6|14|我必伸手攻擊他們，使他們的地荒廢，從 第伯拉他 的曠野起 ，一切的住處都荒涼。他們就知道我是耶和華。」
EZEK|7|1|耶和華的話又臨到我，說：
EZEK|7|2|「你，人子啊，主耶和華對 以色列 地如此說：結局，結局臨到了地的四境！
EZEK|7|3|現在你的結局已經來臨；我要使我的怒氣臨到你，也要按你的行為審判你，照你所做一切可憎的事懲罰你。
EZEK|7|4|我的眼必不顧惜你，也不可憐你，卻要按你所做的報應你，照你們中間可憎的事懲罰你；你就知道我是耶和華。
EZEK|7|5|「主耶和華如此說：災難，惟一的災難 ，看哪，臨近了！
EZEK|7|6|結局到了，結局到了，它要醒起來攻擊你。看哪，它已來到！
EZEK|7|7|境內的居民哪，厄運臨到你；時候到了，日子近了，有鬧鬨，但不是山上歡呼的聲音。
EZEK|7|8|我快要將我的憤怒傾倒在你身上，向你發盡我的怒氣，按你的行為審判你，照你所做一切可憎的事懲罰你。
EZEK|7|9|我的眼必不顧惜你，也不可憐你，必按你所做的報應你，照你中間可憎的事懲罰你；你就知道擊打你的是我─耶和華。
EZEK|7|10|「看哪，那日子！看哪，已來到！厄運已經發生！杖已開花，驕傲已發芽。
EZEK|7|11|殘暴興起，成了罰惡的杖。他們將一無所有，他們的富足 、他們的財寶 都不復存在；他們中間也不再有尊榮。
EZEK|7|12|時候到了，日子近了，買主不可歡喜，賣主也不用愁煩，因為烈怒已經臨到他們眾人身上。
EZEK|7|13|賣主即使存活，也不能討回所賣的，因為這異象關乎他們眾人；誰都不能討回，也沒有人能在罪孽中使自己的生命剛強。」
EZEK|7|14|「他們吹了角，預備齊全，卻無一人出戰，因為我的烈怒臨到他們眾人身上。
EZEK|7|15|外有刀劍，內有瘟疫、饑荒。在田野的，必因刀劍而死；在城中的，必遭饑荒、瘟疫吞滅。
EZEK|7|16|其中倖存的要逃脫，各人因自己的罪孽在山上發出悲聲，如谷中的鴿子哀鳴；
EZEK|7|17|雙手發軟，膝蓋軟弱如水，
EZEK|7|18|腰束麻布，戰慄籠罩他們；各人臉上羞愧，頭上光禿。
EZEK|7|19|他們要把銀子拋棄在街上，看金子如污穢之物。正當耶和華發怒的日子，金銀不能拯救他們，不能滿足食慾，也不能使肚腹飽滿，反倒成了自己罪孽的絆腳石。
EZEK|7|20|他們用所誇耀華美的妝飾製造可憎可厭的偶像，所以我使他們看它如污穢之物。
EZEK|7|21|我必將它交給外邦人為掠物，交給地上的惡人為擄物；他們要褻瀆它。
EZEK|7|22|他們褻瀆我寶貴之所 ，強盜也進去褻瀆它。我必轉臉不顧 以色列 人 。
EZEK|7|23|「要製造鎖鏈；因為遍地都有流血的罪，滿城都是殘暴的事。
EZEK|7|24|所以，我要使列國中最兇惡的人前來佔據他們的房屋；我要止息殘暴人的驕傲，他們的聖所也要被褻瀆。
EZEK|7|25|毀滅來到；他們求平安，卻沒有平安。
EZEK|7|26|災害加上災害，風聲接連風聲；他們要向先知尋求異象，但祭司的教誨、長老的謀略都必斷絕。
EZEK|7|27|君王要悲哀，官長要披絕望為衣，這地百姓的手都發顫。我必照他們所做的待他們，按他們所應得的審判他們，他們就知道我是耶和華。」
EZEK|8|1|第六年六月初五，我坐在家中； 猶大 的眾長老坐在我面前。在那裏主耶和華的手降在我身上。
EZEK|8|2|我觀看，看哪，有形像彷彿火 的形狀，從他腰部以下形狀是火，從他腰部以上有光輝的形狀，好像閃耀的金屬。
EZEK|8|3|他伸出一隻手的樣式，抓住我的一綹頭髮，靈就將我舉到天地中間；在上帝的異象中，他帶我到 耶路撒冷 朝北的內院門口，在那裏有惹動妒忌的偶像的座位，它惹動了妒忌。
EZEK|8|4|看哪，在那裏有 以色列 上帝的榮耀，形狀與我在平原所見的一樣。
EZEK|8|5|上帝對我說：「人子啊，你舉目向北觀看。」我就舉目向北觀看，看哪，祭壇門北邊的門口有那惹動妒忌的偶像。
EZEK|8|6|他又對我說：「人子啊，你看見 以色列 家所做的嗎？他們在這裏做了極其可憎的事，使我遠離我的聖所。你還要看見另有極其可憎的事。」
EZEK|8|7|他領我到院子門口。我觀看，看哪，牆上有一個洞。
EZEK|8|8|他對我說：「人子啊，你要挖牆。」我就挖牆。看哪，有一扇門。
EZEK|8|9|他說：「你進去，看他們在這裏所做可憎的惡事。」
EZEK|8|10|於是我進去看。看哪，四面牆上刻著各樣爬行的動物、可憎的走獸和 以色列 家各樣的偶像。
EZEK|8|11|以色列 家的七十個長老站在這些像前， 沙番 的兒子 雅撒尼亞 也站在其中，各人手拿他的香爐，煙雲的香氣上騰。
EZEK|8|12|他對我說：「人子啊，你看見 以色列 家的長老，暗中在自己偶像的房間裏所做的嗎？因為他們說：『耶和華看不見我們；耶和華已經離棄這地。』」
EZEK|8|13|他又說：「你還要看見他們所做另外極其可憎的事。」
EZEK|8|14|他領我到耶和華殿朝北的門口。看哪，在那裏有婦女們坐著，為 搭模斯 哭泣。
EZEK|8|15|他對我說：「人子啊，你看見了嗎？你還要看見比這更可憎的事。」
EZEK|8|16|然後他領我到耶和華殿的內院。看哪，在耶和華殿門口、走廊和祭壇中間，約有二十五個人背向耶和華的殿，面向東方，向東拜太陽。
EZEK|8|17|他對我說：「人子啊，你看見了嗎？ 猶大 家在這裏行可憎的事還算為小嗎？他們遍地行殘暴，再三惹我發怒。看哪，他們手拿枝條舉向鼻前 ！
EZEK|8|18|因此，我也要以憤怒行事。我的眼必不顧惜，也不可憐他們；他們雖在我耳邊大聲呼求，我還是不聽。」
EZEK|9|1|他在我耳邊大聲喊叫，說：「上前來啊，懲罰這城的人，手中要各拿毀滅的兵器。」
EZEK|9|2|看哪，有六個人從朝北的 上門 而來，各人手裏拿著致命的兵器；他們當中有一人身穿細麻衣，腰間繫著文士用的墨盒。他們進來，站在銅的祭壇旁。
EZEK|9|3|在基路伯之上， 以色列 上帝的榮耀從那裏上升，到殿的入口處。上帝召那身穿細麻衣、腰間繫著墨盒的人前來。
EZEK|9|4|耶和華對他說：「你去走遍 耶路撒冷 全城，那些為城中所做可憎之事嘆息哀哭的人，你要在他們額上做記號。」
EZEK|9|5|我耳中聽見耶和華對其餘的人說：「要跟隨他走遍全城去擊殺。你們的眼不要顧惜，也不要可憐他們。
EZEK|9|6|要將年老的、年輕的、少女、孩童和婦女，從我的聖所開始全都殺盡，只是不可挨近凡有記號的人。」於是他們從殿前的長老殺起。
EZEK|9|7|他對他們說：「要使這殿污穢，使院中遍滿被殺的人。你們出去吧！」他們就出去，在城中擊殺。
EZEK|9|8|他們擊殺的時候，只剩我一人，我就臉伏在地上，呼喊說：「唉！主耶和華啊，你將憤怒傾倒在 耶路撒冷 ，豈要把 以色列 所剩餘的人都滅絕嗎？」
EZEK|9|9|他對我說：「 以色列 家和 猶大 家的罪孽極其重大。遍地都有流血的事，滿城有冤屈，因為他們說：『耶和華已經離棄這地，他看不見我們。』
EZEK|9|10|因此，我的眼必不顧惜，也不可憐他們，要照他們所做的報應在他們頭上。」
EZEK|9|11|看哪，那身穿細麻衣、腰間繫著墨盒的人回覆這事說：「我已經照你所吩咐的做了。」
EZEK|10|1|我觀看，看哪，在穹蒼之中，也就是基路伯的頭上，有藍寶石的形狀，彷彿寶座的形像顯在他們上面。
EZEK|10|2|耶和華對那身穿細麻衣的人說：「你進到基路伯下面旋轉的輪子中，從基路伯之間取出火炭裝滿兩手掌，撒在城上。」 我親眼看見他進去。
EZEK|10|3|那人進去的時候，基路伯站在殿的南邊，雲彩充滿了內院。
EZEK|10|4|耶和華的榮耀從基路伯那裏上升，到殿的入口處；殿內滿佈雲彩，院子也充滿了耶和華榮耀的光輝。
EZEK|10|5|基路伯翅膀的響聲傳到外院，好像全能上帝說話的聲音。
EZEK|10|6|耶和華吩咐那身穿細麻衣的人說：「要從基路伯之間旋轉的輪子中取火。」那人就進去站在一個輪子旁邊。
EZEK|10|7|基路伯中的一個基路伯伸手到基路伯中間的火那裏，取一些放在那身穿細麻衣人的手掌中，那人拿了就出去。
EZEK|10|8|在基路伯翅膀以下，顯出有人手的樣式。
EZEK|10|9|我又觀看，看哪，這些基路伯的旁邊有四個輪子。一個基路伯旁有一個輪子，另一個基路伯旁也有一個輪子；輪子的形狀好像水蒼玉石。
EZEK|10|10|至於四輪的形狀，都是一個樣式，好像輪中套輪。
EZEK|10|11|輪子行走的時候，向四方都能直行，行走時並不轉彎。頭轉向何方，它們也隨著向何方行走，行走時並不轉彎。
EZEK|10|12|基路伯的全身，連背帶手和翅膀，並輪子周圍都佈滿眼睛。他們四個的輪子都是如此。
EZEK|10|13|我耳中聽見這些輪子稱為「旋轉的輪」。
EZEK|10|14|基路伯各有四張臉：第一是基路伯的臉，第二是人的臉，第三是獅子的臉，第四是鷹的臉。
EZEK|10|15|基路伯升上去了；這就是我在 迦巴魯河 邊所看見的活物。
EZEK|10|16|基路伯行走，輪子也在旁邊行走。基路伯展開翅膀，離地上升，輪子也不轉離他們的旁邊。
EZEK|10|17|基路伯站住，輪子也站住；基路伯上升，輪子也跟著上升，因為活物的靈在輪中。
EZEK|10|18|耶和華的榮耀離開殿的入口處，停在基路伯之上。
EZEK|10|19|基路伯展開翅膀，在我眼前離地上升；他們離去的時候，輪子在旁邊，都停在耶和華殿的東門口。在他們上面有 以色列 上帝的榮耀。
EZEK|10|20|這是我在 迦巴魯河 邊所見的活物，他們在 以色列 上帝之下；因此我知道他們是基路伯。
EZEK|10|21|他們各有四張臉、四個翅膀，翅膀以下有人手的樣式。
EZEK|10|22|至於他們臉的模樣，以及身體的形像 ，正是我從前在 迦巴魯河 邊所看見的。他們各自往前直行。
EZEK|11|1|靈將我舉起，帶我到耶和華聖殿面向東方的東門。看哪，門口有二十五個人。我見其中有百姓的領袖 押朔 的兒子 雅撒尼亞 和 比拿雅 的兒子 毗拉提 。
EZEK|11|2|耶和華對我說：「人子啊，他們就是圖謀罪孽，在這城中設計惡謀的人。
EZEK|11|3|他們說：『蓋房屋的時候尚未臨近；這城是鍋，我們是肉。』
EZEK|11|4|人子啊，因此你當說預言，說預言攻擊他們。」
EZEK|11|5|耶和華的靈降在我身上，對我說：「你當說，耶和華如此說： 以色列 家啊，你們所說的，你們心裏所想的，我都知道。
EZEK|11|6|你們在這城裏大行屠殺，被殺的人遍滿街道。
EZEK|11|7|所以主耶和華如此說：你們在城中殺的人是肉，這城是鍋；你們卻要從其中被帶出去。
EZEK|11|8|你們怕刀劍，我卻要使刀劍臨到你們。這是主耶和華說的。
EZEK|11|9|我要把你們從這城中帶出去，交在外邦人的手裏，且要在你們中間施行審判。
EZEK|11|10|你們要仆倒在刀下；我必在 以色列 的邊界審判你們，你們就知道我是耶和華。
EZEK|11|11|這城必不作你們的鍋，你們也不作鍋中的肉。我要在 以色列 的邊界審判你們，
EZEK|11|12|你們就知道我是耶和華；因為你們不遵行我的律例，也不順從我的典章，卻隨從你們四圍列國的規條。」
EZEK|11|13|我正說預言的時候， 比拿雅 的兒子 毗拉提 死了。於是我臉伏在地，大聲呼叫說：「唉！主耶和華啊，你要把 以色列 剩餘的人都滅絕淨盡嗎？」
EZEK|11|14|耶和華的話臨到我，說：
EZEK|11|15|「人子啊， 耶路撒冷 的居民對你的兄弟、你的本家、你的親屬、 以色列 全家所有的人說：『你們遠離耶和華吧！這地是賜給我們為業的。』
EZEK|11|16|所以你當說：『主耶和華如此說：我雖將 以色列 全家遠遠流放到列國，使他們分散在列邦，我卻要在他們所到的列邦，暫時作他們的聖所。』
EZEK|11|17|你當說：『主耶和華如此說：我必從萬民中召集你們，從分散的列邦中聚集你們，又將 以色列 地賜給你們。』
EZEK|11|18|他們到了那裏，必從其中除掉一切可憎之物、可厭的事。
EZEK|11|19|我要使他們有合一的心，也要將新靈放在你們 裏面，又從他們的肉體中除掉石心，賜給他們肉心，
EZEK|11|20|使他們順從我的律例，謹守遵行我的典章。他們要作我的子民，我要作他們的上帝。
EZEK|11|21|至於那些心中隨從可憎之物、可厭的事的人，我必照他們所做的報應在他們頭上。這是主耶和華說的。」
EZEK|11|22|於是，基路伯展開翅膀，輪子都在他們旁邊；在他們上面有 以色列 上帝的榮耀。
EZEK|11|23|耶和華的榮耀從城中上升，停在城東的那座山上。
EZEK|11|24|靈將我舉起，在異象中上帝的靈將我帶回 迦勒底 地，到被擄的人那裏；之後我所見的異象就離我上升去了。
EZEK|11|25|我就把耶和華指示我的一切事都說給被擄的人聽。
EZEK|12|1|耶和華的話臨到我，說：
EZEK|12|2|「人子啊，你住在悖逆之家中；他們有眼可看卻看不見，有耳可聽卻聽不到，因為他們是悖逆之家。
EZEK|12|3|所以人子啊，你要收拾被擄時需用的物件，白天在他們眼前離去，在他們眼前離開你所住的地方，移到別處去；他們雖是悖逆之家，或者可以領悟。
EZEK|12|4|你要白天在他們眼前拿出你被擄時需用的物件。到了晚上，要在他們眼前離去，像被擄的人離去一樣。
EZEK|12|5|你要在他們眼前挖通牆壁，從其中將物件帶出去 。
EZEK|12|6|到天黑時，在他們眼前背在肩上帶走 ，並要蒙住臉看不見地，因為我要使你成為 以色列 家的預兆。」
EZEK|12|7|我就照著所吩咐的去做，白天拿出被擄時需用的物件。到了晚上，用手挖通牆壁；天黑的時候，在他們眼前背在肩上帶走。
EZEK|12|8|次日早晨，耶和華的話臨到我，說：
EZEK|12|9|「人子啊， 以色列 家，就是那悖逆之家，豈不是問你說：『你在做甚麼呢？』
EZEK|12|10|你要對他們說：『主耶和華如此說：這是關乎 耶路撒冷 君王和其中 以色列 全家的默示。』
EZEK|12|11|你要說：『我是你們的預兆：我怎樣做，他們所遭遇的也必這樣，他們必被擄去，作俘虜。』
EZEK|12|12|他們中間的君王也必在天黑時把物件背在肩上帶走。他們要挖通牆壁，從其中帶出去 。他必蒙住臉，眼看不見地。
EZEK|12|13|我要把我的網撒在他身上，他就被我的羅網纏住。我要帶他到 迦勒底 人之地的 巴比倫 ；他沒有看見那地，就死在那裏。
EZEK|12|14|我要把四圍幫助他的和他所有的軍隊分散到四方 ，也要拔刀追趕他們。
EZEK|12|15|我把他們驅逐到列國，分散在列邦的時候，他們就知道我是耶和華。
EZEK|12|16|我卻要留下他們當中幾個人得免刀劍、饑荒、瘟疫，使他們在所到的列國述說自己所做一切可憎的事；他們就知道我是耶和華。」
EZEK|12|17|耶和華的話臨到我，說：
EZEK|12|18|「人子啊，你吃飯時必戰抖，喝水時必驚惶憂慮。
EZEK|12|19|你要對這地的百姓說：主耶和華論 以色列 地的 耶路撒冷 居民如此說，他們吃飯時必憂慮，喝水時必驚惶，因其中居民所行殘暴的事，這地必然荒廢，一無所存。
EZEK|12|20|有人居住的城鎮必變為廢墟，地必荒涼；你們就知道我是耶和華。」
EZEK|12|21|耶和華的話臨到我，說：
EZEK|12|22|「人子啊，在 以色列 地你們怎麼有這俗語說：『日子延長，一切異象卻落了空』呢？
EZEK|12|23|你要告訴他們說：『主耶和華如此說：我必令這俗語止息， 以色列 中不再有人引用這俗語。』你卻要對他們說：『日子臨近，一切的異象都必應驗。』
EZEK|12|24|從此以後， 以色列 家不再有虛假的異象和奉承的占卜。
EZEK|12|25|我─耶和華說話，所說的必定實現，不再耽延。你們這悖逆之家啊，你們在世的日子，我所說的話必定實現。這是主耶和華說的。」
EZEK|12|26|耶和華的話臨到我，說：
EZEK|12|27|「人子，看哪， 以色列 家的人說：『他所見的異象是許多日子以後的事，所說的預言是指著遙遠的時候。』
EZEK|12|28|所以你要對他們說：『主耶和華如此說：我的話不再有一句耽延，我所說的話必定實現。』這是主耶和華說的。」
EZEK|13|1|耶和華的話臨到我，說：
EZEK|13|2|「人子啊，你要說預言，攻擊 以色列 中說預言的先知，對那些隨心說預言的人說：『你們當聽耶和華的話。』」
EZEK|13|3|主耶和華如此說：「禍哉！那些愚頑的先知，隨從自己的心意，卻一無所見
EZEK|13|4|以色列 啊，你的先知好像廢墟中的狐狸，
EZEK|13|5|沒有上去堵住缺口，也沒有為 以色列 家重修城牆，使它在耶和華的日子來臨時，可以在戰爭中站得住。
EZEK|13|6|他們看見的是虛假，是謊詐的占卜，說是耶和華說的；其實耶和華並沒有差遣他們，他們卻指望那話必站立得住。
EZEK|13|7|你們豈不是見了虛假的異象嗎？豈不是說了謊詐的占卜嗎？你們說，這是耶和華說的，其實我沒有說過。」
EZEK|13|8|所以主耶和華如此說：「因你們說的是虛假，見的是謊詐，所以，看哪，我要敵對你們。這是主耶和華說的。
EZEK|13|9|我的手必攻擊那見虛假異象、用謊詐占卜的先知，他們必不列在我百姓的會中，不錄在 以色列 家的名冊上，也不能進入 以色列 地；你們就知道我是主耶和華。
EZEK|13|10|他們誘惑我的百姓，說：『平安！』其實沒有平安，就像有人築牆壁，看哪，他們倒去粉刷它。
EZEK|13|11|所以你要對那些粉刷的人說：『牆要倒塌，暴雨漫過。你們大冰雹啊，要降下 ，狂風要吹裂這牆。』
EZEK|13|12|看哪，這牆倒塌，人豈不是要問你們說：『你們所粉刷的在哪裏呢？』」
EZEK|13|13|所以主耶和華如此說：「我要發怒，使狂風吹裂它，在怒中令暴雨漫過，又發怒降下大冰雹，毀壞它。
EZEK|13|14|我要這樣拆毀你們那粉飾的牆，把它夷為平地，以致根基露出；牆一倒塌，你們也要在其中滅亡。你們就知道我是耶和華。
EZEK|13|15|我要對牆和粉刷它的人發盡我的憤怒，我 要對你們說：『牆沒有了！粉刷它的人也沒有了！』
EZEK|13|16|這就是 以色列 的先知，他們指著 耶路撒冷 說預言，見到這城平安的異象，其實沒有平安。這是主耶和華說的。」
EZEK|13|17|「你，人子啊，要面向你百姓中隨心說預言的婦女們，說預言攻擊她們，
EZEK|13|18|說，主耶和華如此說：『這些婦女有禍了！她們為眾人的手腕縫驅邪帶，替身材高矮不同的人做頭巾，為要獵取人的性命。難道你們要獵取我百姓的性命，使自己存活嗎？
EZEK|13|19|你們為幾把大麥、幾塊餅，在我的百姓中褻瀆我，對那肯聽謊言的百姓說謊言，讓不該死的人死，讓不該活的人活。』」
EZEK|13|20|所以主耶和華如此說：「看哪，我要對付你們那用以獵取人，如獵飛鳥般的驅邪帶。我要把驅邪帶從你們的手腕扯去，釋放那些如飛鳥被你們獵取的人。
EZEK|13|21|我也必撕裂你們的頭巾，救我百姓脫離你們的手，使他們不再被獵取，落在你們手中；你們就知道我是耶和華。
EZEK|13|22|我未曾使義人傷心，你們卻以謊話使他傷心，且又堅固惡人的手，不使他回轉離開惡道得以存活。
EZEK|13|23|所以，你們必不再看見虛假的異象，也不再行占卜的事；我要救我的百姓脫離你們的手；你們就知道我是耶和華。」
EZEK|14|1|有幾個 以色列 的長老到我這裏來，坐在我面前。
EZEK|14|2|耶和華的話臨到我，說：
EZEK|14|3|「人子啊，這些人在心中設立偶像，把陷自己於罪的絆腳石放在面前，我真的能讓他們求問嗎？
EZEK|14|4|所以你要告訴他們，對他們說：『主耶和華如此說： 以色列 家的人，凡在心中設立偶像，把陷自己於罪的絆腳石放在面前，卻來到先知那裏的，我─耶和華在他所求的事上，必因他拜許多偶像向他施行報應 ，
EZEK|14|5|為要奪回 以色列 家的心，他們全都拜偶像，與我疏遠了。』
EZEK|14|6|「所以你要對 以色列 家說：『主耶和華如此說：回轉吧！回轉離開你們的偶像，轉臉離開一切可憎的事。』
EZEK|14|7|因為 以色列 家的人，或在 以色列 中寄居的外人，凡與我隔絕，在心中設立偶像，把陷自己於罪的絆腳石放在面前，卻來到先知那裏，要為自己的事求問我的，我─耶和華必親自報應他。
EZEK|14|8|我要向那人變臉，使他成為警戒和笑柄，並且我要把他從我民中剪除；你們就知道我是耶和華。
EZEK|14|9|先知若被騙說了一句預言，是我─耶和華騙了那先知，我要伸手攻擊他，把他從我百姓 以色列 中除滅。
EZEK|14|10|他們必擔當自己的罪孽。先知的罪孽和求問之人的罪孽都一樣，
EZEK|14|11|使 以色列 家不再走迷離開我，也不再因各樣的罪過玷污自己，卻要作我的子民，我也作他們的上帝。這是主耶和華說的。」
EZEK|14|12|耶和華的話臨到我，說：
EZEK|14|13|「人子啊，若有一國犯罪干犯我，我也伸手攻擊它，斷絕他們糧食的供應，使饑荒臨到那地，將人與牲畜從其中剪除；
EZEK|14|14|雖有 挪亞 、 但以理 、 約伯 這三人在那裏，他們只能因自己的義救自己的命。這是主耶和華說的。
EZEK|14|15|我若使惡獸經過那地，大肆蹂躪，使地荒涼，以致因這些獸，人都不得經過；
EZEK|14|16|雖有這三人在其中，主耶和華說：我指著我的永生起誓，他們不能救兒子女兒，只有他們自己可以得救，那地仍然荒涼。
EZEK|14|17|或者我使刀劍臨到那地，說：『讓刀劍穿越那地』，以致我把人與牲畜從其中剪除；
EZEK|14|18|雖有這三人在其中，主耶和華說：我指著我的永生起誓，他們不能救兒子女兒，只有他們自己可以得救。
EZEK|14|19|或者我叫瘟疫流行那地，把我的憤怒帶著血傾在其中，好使人與牲畜從其中剪除；
EZEK|14|20|雖有 挪亞 、 但以理 、 約伯 在那裏，主耶和華說：我指著我的永生起誓，他們不能救兒子女兒，只能因自己的義救自己的命。
EZEK|14|21|「主耶和華如此說：我若將這四樣大災，就是刀劍、饑荒、惡獸、瘟疫降在 耶路撒冷 ，將人與牲畜從其中剪除，豈不是更嚴重嗎？
EZEK|14|22|看哪，在那裏必有倖免於難的人帶著兒子女兒；看哪，他們來到你們這裏；你們看見他們的所作所為，就會因我降給 耶路撒冷 的災禍，因我降給它的一切，得到安慰。
EZEK|14|23|你們因看見他們的所作所為，得到安慰，就會知道我在 耶路撒冷 所做的並非毫無緣故。這是主耶和華說的。」
EZEK|15|1|耶和華的話臨到我，說：
EZEK|15|2|「人子啊，葡萄樹比一切其他的樹，就是樹林裏眾樹木的樹枝，有甚麼長處呢？
EZEK|15|3|可以從其中取木料來做工嗎？人可以拿來做釘子，掛東西在上面嗎？
EZEK|15|4|看哪，它已經拋在火中當柴燒，火既燒了兩頭，中間也燒焦了，它還有甚麼用處呢？
EZEK|15|5|看哪，它完整的時候尚且不能拿來做工，何況被火燒焦了，還能拿來做工嗎？
EZEK|15|6|所以，主耶和華如此說：我怎樣使林中樹裏的葡萄樹在火中當柴燒，我也必照樣對待 耶路撒冷 的居民。
EZEK|15|7|我必向他們變臉；他們雖從火中逃出來，火仍要燒滅他們。我向他們變臉的時候，你們就知道我是耶和華。
EZEK|15|8|我必使這地荒涼，因為他們做了背叛的事。這是主耶和華說的。」
EZEK|16|1|耶和華的話臨到我，說：
EZEK|16|2|「人子啊，你要使 耶路撒冷 知道它那些可憎的事。
EZEK|16|3|你要說，主耶和華對 耶路撒冷 如此說：你的根源，你的出身，是在 迦南 地；你的父親是 亞摩利 人，母親是 赫 人。
EZEK|16|4|論到你出世的景況，在你出生的日子沒有人為你斷臍帶，也沒有用水清洗，使你潔淨；沒有人撒鹽在你身上，也沒有人用布包你。
EZEK|16|5|沒有人顧惜你，為你做一件這樣的事來可憐你。你卻被扔在田野上面，因你出生的日子就被厭惡。
EZEK|16|6|「我從你旁邊經過，見你在血中打滾，就對你說：『你雖在血中，卻要活下去！』我又說：『你雖在血中，卻要活下去！』
EZEK|16|7|我使你成長如田間所生長的；你就漸長，美而又美 ，兩乳成形，頭髮秀長，但你仍然赤身露體。
EZEK|16|8|「我從你旁邊經過看見你，看哪，正是你渴慕愛情的時候，我就用我衣服的邊搭在你身上，遮蓋你的赤體；又向你起誓，與你立約，你就歸我。這是主耶和華說的。
EZEK|16|9|那時我用水洗你，洗淨你身上的血，又用油抹你。
EZEK|16|10|我使你身穿錦繡衣裳，腳穿海狗皮鞋，用細麻布裹著你，精緻衣料披在你身上。
EZEK|16|11|我用首飾打扮你：我把手鐲戴在你手上，項鏈在你頸上，
EZEK|16|12|我也把環子戴在你鼻上，耳環在你耳上，華冠在你頭上。
EZEK|16|13|這樣，你就有金銀的首飾，穿的是細麻衣和精緻衣料，以及錦繡衣裳；吃的是細麵、蜂蜜和油。你也極其美貌，配登王后之位。
EZEK|16|14|你美貌的名聲傳到列國，因我加給你榮華，使你完美。這是主耶和華說的。
EZEK|16|15|「只是你仗著自己美貌，又憑著你的名聲行淫。你向路人縱情淫亂，你的美貌就屬於他的了 。
EZEK|16|16|你拿你的衣服為自己做成彩色丘壇，在其上行淫。這樣的事本不該有，以後也不該發生。
EZEK|16|17|你拿我所賜給你的那些美麗的金銀寶物，為自己製造男性的偶像，與它們行淫；
EZEK|16|18|你拿你的錦繡衣裳為它們披上，把我的膏油和香料擺在它們面前；
EZEK|16|19|你把我賜給你的食物，就是我賜給你享用的細麵、油和蜂蜜，都擺在它們面前作為馨香的供物。事情就是這樣。這是主耶和華說的。
EZEK|16|20|你拿你為我所生的兒女獻給它們吞噬。你的淫亂豈是小事？
EZEK|16|21|你竟把我的兒女殺了，使他們經火獻給它們！
EZEK|16|22|你做這一切可憎和淫亂的事，並未追念你幼年的日子，那時你赤身露體，在血中打滾。」
EZEK|16|23|「你有禍了！你有禍了！這是主耶和華說的。你做這一切惡事之後，
EZEK|16|24|又為自己建造土墩，在各廣場上築起高臺。
EZEK|16|25|你在各個街頭建造高臺，使你的美貌變為可憎；又向所有過路的人招手 ，多行淫亂。
EZEK|16|26|你也和你那放縱情慾的鄰邦 埃及 人行淫，增添你的淫亂，惹我發怒。
EZEK|16|27|看哪，我伸手攻擊你，減少你的福分，卻將你交給恨惡你的 非利士 人 ，讓他們任意待你。他們為你的淫行也感到羞恥。
EZEK|16|28|你尚且不滿意，又與 亞述 人行淫，但與他們行淫之後，仍不滿足；
EZEK|16|29|於是你與那稱為貿易之地的 迦勒底 多行淫亂，即使這樣，你仍不滿足。
EZEK|16|30|「你的心何等脆弱！這是主耶和華說的。你做這一切事，都是不知羞恥的妓女所做的，
EZEK|16|31|在各個街頭建造土墩，在各廣場上築高臺；但你藐視行淫的賞金，又不像妓女。
EZEK|16|32|你這行淫的妻子啊，竟然接外人，替代丈夫。
EZEK|16|33|凡妓女都是得人贈禮，你反倒餽贈你所愛的人，倒貼他們，使他們從四圍來與你行淫。
EZEK|16|34|你的淫行與其他婦女相反，不是人要求與你行淫；是你給人賞金，不是人給你賞金；你是相反的。」
EZEK|16|35|「你這妓女啊，要聽耶和華的話。
EZEK|16|36|主耶和華如此說：因你放縱情慾，露出下體，與你所愛的行淫，因你敬拜一切可憎的偶像，就像 自己兒女的血獻給它們，
EZEK|16|37|所以，看哪，我要聚集所有與你交歡的情人，不論是你所愛的或你所恨的，聚集他們從四圍到你那裏來；我要在他們面前暴露你的下體，使他們看盡你的下體。
EZEK|16|38|我也要審判你，如審判淫婦和流人血的婦女一樣。我要在憤怒和妒忌中使流血的罪歸到你身上。
EZEK|16|39|我要把你交在他們手中；他們必拆毀你的土墩，毀壞你的高臺，剝去你的衣服，奪取你美麗的寶物，留下你赤身露體。
EZEK|16|40|他們必聚集眾人攻擊你，用石頭打死你，用刀劍刺透你，
EZEK|16|41|用火焚燒你的房屋，在許多婦女眼前審判你。我必使你不再行淫，你也不再給賞金。
EZEK|16|42|我止息了向你所發的憤怒，我的妒忌也離開了你；這樣，我就平靜，不再惱怒。
EZEK|16|43|因你不追念幼年的日子，反而在這一切的事上惹我發烈怒，所以，看哪，我必照你所做的報應在你頭上。在你一切可憎的事上，你不是還行了淫亂嗎？這是主耶和華說的。」
EZEK|16|44|「看哪，凡說俗語的必用這俗語攻擊你，說：『有其母必有其女。』
EZEK|16|45|你實在是你母親的女兒，厭棄丈夫和兒女；你也是你姊妹的姊妹，厭棄丈夫和兒女。你的母親是 赫 人，父親是 亞摩利 人。
EZEK|16|46|你的姊姊是 撒瑪利亞 ，她和她的女兒們住在你北邊；你的妹妹是 所多瑪 ，她和她的女兒們住在你南邊。
EZEK|16|47|你不只效法她們的行為，照她們可憎的事去做，不消多時 ，你所做的一切就比她們更惡。
EZEK|16|48|主耶和華說：我指著我的永生起誓，你的妹妹 所多瑪 與她的女兒們並未做你和你女兒們所做的事。
EZEK|16|49|看哪，你的妹妹 所多瑪 的罪孽是這樣：她和她的女兒們都驕傲，糧源充足，大享安逸，卻不扶持困苦和貧窮人的手。
EZEK|16|50|她們狂傲，在我面前做可憎的事，我看見了就把她們除掉。
EZEK|16|51|撒瑪利亞 所犯的罪不及你的一半，你所做可憎的事比她更多；比起你所做這一切可憎的事，你的姊妹倒顯為義。
EZEK|16|52|你既為你的姊妹辯護，就要擔當自己的羞辱。因你所犯的罪比她們更可憎，她們比你倒顯為義；你既使你的姊妹顯為義，就要抱愧，擔當自己的羞辱。」
EZEK|16|53|「我必使她們被擄的歸回，使 所多瑪 和她的女兒們、 撒瑪利亞 和她的女兒們，並與你一起被擄的都歸回；
EZEK|16|54|好使你擔當自己的羞辱，為所做的一切抱愧，讓她們得到安慰。
EZEK|16|55|你的妹妹 所多瑪 和她的女兒們必回復原狀； 撒瑪利亞 和她的女兒們必回復原狀；你和你的女兒們也必回復原狀。
EZEK|16|56|在你驕傲的日子，你的妹妹 所多瑪 豈不是你口中的笑柄嗎？
EZEK|16|57|在你的惡行顯露以前，那受了凌辱的 亞蘭 女兒們和 亞蘭 四圍 非利士 的女兒們，都在四圍藐視你。
EZEK|16|58|耶和華說：你的淫蕩和可憎之事，你自己要擔當。」
EZEK|16|59|「主耶和華如此說：你這輕看誓言而背約的，我必照你所做的報應你。
EZEK|16|60|然而我要追念在你幼年時我與你所立的約，也要與你立定永約。
EZEK|16|61|當你接納你的姊姊和妹妹時，你要追念你所行的，自覺慚愧；並且我要將她們賞給你做女兒，卻不是按著我與你所立的約。
EZEK|16|62|我要堅定與你所立的約，你就知道我是耶和華，
EZEK|16|63|使你在我赦免你一切惡行時，心中追念，自覺慚愧，又因羞辱就不再開口。這是主耶和華說的。」
EZEK|17|1|耶和華的話臨到我，說：
EZEK|17|2|「人子啊，你要向 以色列 家出謎語，設比喻，
EZEK|17|3|說，主耶和華如此說：有一隻大鷹，翅膀大，翎毛長，羽毛豐滿，色彩繽紛；牠飛到 黎巴嫩 ，啄去香柏樹梢，
EZEK|17|4|啄斷它頂端的嫩枝，叼到貿易之地，放在商業城中。
EZEK|17|5|牠又從這地取了一些種子，種在肥沃的田裏，栽於豐沛的水源旁，如種植柳樹。
EZEK|17|6|它漸漸生長，成為低矮蔓生的葡萄樹；樹枝伸向那鷹，根部在牠下面。這樣，它就長成了一棵葡萄樹，生出枝子，長出枝幹。
EZEK|17|7|「有一隻 大鷹，翅膀大，羽毛多。看哪，葡萄樹從栽種它的苗圃向這鷹伸出根來，長出枝子，期盼從牠得到澆灌。
EZEK|17|8|這棵樹栽於肥田豐沛的水源旁，原是為了生枝、結果，成為佳美的葡萄樹。
EZEK|17|9|你要說，主耶和華如此說：這棵葡萄樹豈能發旺呢？鷹豈不拔出它的根來，摘光它的果子，使它枯乾，連長出的嫩葉都枯萎了嗎？要把它連根拔除，並不需要費大力或動用許多人。
EZEK|17|10|看哪，葡萄樹雖然栽種了，豈能發旺呢？一經東風擊打，豈不全然枯乾了嗎？它必在生長的苗圃中枯乾了。」
EZEK|17|11|耶和華的話臨到我，說：
EZEK|17|12|「你要對那悖逆之家說：你們不知道這些事是甚麼意思嗎？你要這樣說，看哪， 巴比倫 王曾到 耶路撒冷 ，把其中的君王和官長帶到 巴比倫 去，
EZEK|17|13|又從 以色列 王室後裔中選取一人，與他立約，令他發誓，又擄走國中有勢力的人，
EZEK|17|14|使王國衰弱，不再強盛，只能靠守盟約方得生存。
EZEK|17|15|他卻背叛 巴比倫 王，差派使者前往 埃及 ，要求 埃及 人給他馬匹和許多人。他豈能亨通呢？這樣做的人豈能逃脫呢？他背了約豈能逃脫呢？
EZEK|17|16|主耶和華說：我指著我的永生起誓，他定要死在 巴比倫 ，就是 巴比倫 王所在之處；因為 巴比倫 王立他為王，他竟輕看向王所起的誓，背棄王與他所立的約。
EZEK|17|17|當敵人建土堆，築堡壘，要殲滅許多人時，法老雖有強大軍隊和大批人馬，在戰場上還是不能幫助他。
EZEK|17|18|他輕看誓言，背棄盟約，看哪，雖已投降 ，卻又做這一切的事，他必不能逃脫。
EZEK|17|19|所以主耶和華如此說：我指著我的永生起誓，他既輕看我的誓言，背棄我的約，我必使這罪歸到他頭上。
EZEK|17|20|我要把我的網撒在他身上，他就被我的羅網纏住。我要帶他到 巴比倫 ，在那裏因他背叛我的罪懲罰他。
EZEK|17|21|所有逃跑的 軍隊必倒在刀下；剩餘的也必分散四方 。你們就知道說這話的是我─耶和華。」
EZEK|17|22|主耶和華如此說：「我要從香柏樹高高的樹梢摘取並栽上，從頂端的嫩枝中折下一嫩枝，栽於極高的山上，
EZEK|17|23|栽在 以色列 高處的山上。它就生枝、結果，成為高大的香柏樹，各類飛禽中的鳥都來宿在其下，宿在枝子的蔭下 。
EZEK|17|24|田野的樹木因此就知道是我─耶和華使高樹矮小，使矮樹高大，使綠樹枯乾，使枯樹發旺。我─耶和華說了這話，就必成就。」
EZEK|18|1|耶和華的話又臨到我，說：
EZEK|18|2|「你們在 以色列 地何以有這俗語，『父親吃了酸葡萄，兒子牙齒就酸倒』呢？
EZEK|18|3|主耶和華說：我指著我的永生起誓，你們在 以色列 必不再引用這俗語。
EZEK|18|4|看哪，所有的生命都是屬我的；父親的生命怎樣屬我，兒子的生命也照樣屬我；然而犯罪的，他必定死。
EZEK|18|5|「人若是公義，行公平公義的事：
EZEK|18|6|未曾在山上吃祭物，未曾向 以色列 家的偶像舉目；未曾污辱鄰舍的妻，也未曾在婦人的經期間親近她；
EZEK|18|7|未曾虧負人，而是將欠債之人的抵押品還給他；未曾搶奪人的物件，卻把食物給飢餓的人吃，把衣服給赤身的人穿；
EZEK|18|8|未曾向人取利息，也未曾索取高利，反倒縮手不作惡，在人與人之間施行誠實的判斷；
EZEK|18|9|遵行我的律例，謹守我的典章，按誠實行事 ；這人是公義的，必要存活。這是主耶和華說的。
EZEK|18|10|「他若生了兒子，兒子作強盜，流人的血，作父親的 雖然未犯此過，兒子卻對弟兄 行了以上所說的惡，在山上吃祭物，污辱鄰舍的妻；
EZEK|18|11|
EZEK|18|12|虧負困苦和貧窮的人，搶奪別人的物件，不歸還抵押品，卻向偶像舉目，做可憎的事；
EZEK|18|13|向人取利息，索取高利，這人豈能存活呢？他不能存活。他因做這一切可憎的事，必要死亡，他的血要歸到自己身上。
EZEK|18|14|「看哪，他若生了兒子，兒子見父親所犯的一切罪，他見了，卻不照樣去做；
EZEK|18|15|他未曾在山上吃祭物，未曾向 以色列 家的偶像舉目，未曾污辱鄰舍的妻；
EZEK|18|16|也未曾虧負人，未曾取人的抵押品，未曾搶奪人的物件，卻把食物給飢餓的人吃，把衣服給赤身的人穿，
EZEK|18|17|縮手不害困苦人，未曾向人索取利息或高利；反倒順從我的典章，遵行我的律例；如此，他必不因父親的罪孽死亡，定要存活。
EZEK|18|18|至於他父親，因為施行欺壓，搶奪弟兄，在百姓中行不善，看哪，他必因自己的罪孽死亡。
EZEK|18|19|「你們還說：『兒子為甚麼不擔當父親的罪孽呢？』兒子若行公平公義的事，謹守遵行我一切的律例，他必要存活。
EZEK|18|20|惟有犯罪的，卻必死亡。兒子不擔當父親的罪孽，父親也不擔當兒子的罪孽。義人的善果要歸自己，惡人的惡報也要歸自己。
EZEK|18|21|「惡人若回轉離開所做的一切罪惡，謹守我的一切律例，行公平公義的事，他必要存活，不致死亡。
EZEK|18|22|他所犯的一切罪過都不被記念；他因所行的義，必要存活。
EZEK|18|23|惡人死亡，豈是我所喜悅的呢？我豈不是喜悅他回轉離開所行的道而存活嗎？這是主耶和華說的。
EZEK|18|24|至於義人，他若轉離義行而作惡，照著惡人所做一切可憎的事去做，豈能存活呢？他所行的一切義都不被記念；反而因所行的惡、所犯的罪死亡。
EZEK|18|25|「你們卻說：『主的道不公平！』 以色列 家啊，你們要聽，我的道不公平嗎？你們的道不是不公平嗎？
EZEK|18|26|義人若轉離義行而作惡，他就因這些惡而死亡。他要死在他所作的惡中。
EZEK|18|27|惡人若回轉離開所行的惡，行公平公義的事，他必救自己的命；
EZEK|18|28|因為他省察，回轉離開所犯的一切罪過，他必要存活，不致死亡。
EZEK|18|29|以色列 家還說：『主的道不公平！』 以色列 家啊，我的道不公平嗎？你們的道不是不公平嗎？
EZEK|18|30|所以， 以色列 家啊，我必按你們各人所做的審判你們。當回轉，回轉離開你們一切的罪過，免得罪孽成為你們的絆腳石。這是主耶和華說的。
EZEK|18|31|你們要把所犯的一切罪過盡行拋棄，為自己造一個新的心和新的靈。 以色列 家啊，你們為甚麼要死呢？
EZEK|18|32|我不喜歡有任何人死亡，所以你們當回轉，要存活！這是主耶和華說的。」
EZEK|19|1|你當為 以色列 的領袖們唱哀歌，
EZEK|19|2|說： 你的母親在獅子中 是怎樣的母獅呢？ 牠蹲伏在少壯獅子中， 養育小獅子。
EZEK|19|3|牠養大了其中一隻小獅子， 成了少壯獅子， 學會抓食， 牠就吃人。
EZEK|19|4|列國聽見了就把牠逮住在他們的坑裏， 用鉤子拉牠到 埃及 地去。
EZEK|19|5|母獅見自己等候， 期望落空， 就從小獅子中取一隻 ， 養為少壯獅子；
EZEK|19|6|牠在眾獅子中徜徉， 長大成為少壯獅子， 學會抓食， 牠就吃人。
EZEK|19|7|牠拆毀他們的宮殿 ， 使他們的城鎮變為廢墟； 因牠咆哮的聲音， 遍地和其中所充滿的都荒廢了。
EZEK|19|8|於是四圍列國 從各省前來攻擊牠， 把網撒在牠身上， 把牠逮住在他們的坑裏。
EZEK|19|9|他們又用鉤子鉤住牠，把牠放入籠中， 帶到 巴比倫 王那裏， 把牠押進城堡， 以色列 山上就不再聽見牠的聲音。
EZEK|19|10|你的母親如葡萄樹， 在葡萄園中 ， 栽於水邊，因為水多， 就多結果子，多生枝子；
EZEK|19|11|它長出堅固的枝幹， 可作統治者的權杖。 這枝幹高舉在茂密的樹枝中， 可見樹身高大，枝子繁多。
EZEK|19|12|但在烈怒中它被拔出，摔在地上； 東風吹乾其果子， 那堅固的枝幹因折斷而枯乾， 被火燒燬；
EZEK|19|13|如今這葡萄樹移植於曠野， 在乾旱無水之地，
EZEK|19|14|火從枝幹中發出， 燒滅它的枝條和它的果子 ， 以致不再有堅固的枝幹， 可作統治者的權杖。 這是哀傷之歌，成為一首哀歌。
EZEK|20|1|第七年五月初十，有 以色列 的幾個長老前來求問耶和華，坐在我面前。
EZEK|20|2|耶和華的話臨到我，說：
EZEK|20|3|「人子啊，你要告訴 以色列 的長老，對他們說，主耶和華如此說：你們來是為求問我嗎？主耶和華說：我指著我的永生起誓，我必不讓你們求問。
EZEK|20|4|人子啊，你要審問他們嗎？你要審問嗎？你當使他們知道他們祖先那些可憎的事；
EZEK|20|5|你要對他們說，主耶和華如此說：當日我揀選 以色列 ，對 雅各 家的後裔起誓，在 埃及 地向他們顯現，起誓說：我是耶和華─你們的上帝；
EZEK|20|6|那日我向他們起誓，要領他們出 埃及 地，到我為他們所找到的流奶與蜜之地，就是全地中最美好之地。
EZEK|20|7|我對他們說，你們各人要拋棄眼中所喜愛的可憎之物，不可用 埃及 的偶像玷污自己。我是耶和華─你們的上帝。
EZEK|20|8|他們卻悖逆我，不肯聽從我，不拋棄他們眼中所喜愛的可憎之物，離棄 埃及 的偶像。 「我就說，在 埃及 地，我要把我的憤怒傾倒在他們身上，向他們發盡我的怒氣。
EZEK|20|9|我這麼做是為了我名的緣故，免得我的名在他們所居住之列國眼中被褻瀆；我曾在這些列國眼前向他們顯現，領他們出了 埃及 地。
EZEK|20|10|我領他們出 埃及 地，帶他們到曠野。
EZEK|20|11|我將我的律例賜給他們，將我的典章指示他們；人若遵行就必因此存活。
EZEK|20|12|我將我的安息日賜給他們，在我與他們中間作記號，讓他們知道我─耶和華是使他們分別為聖的。
EZEK|20|13|以色列 家卻在曠野中悖逆我，不順從我的律例，厭棄我的典章；人若遵行就必因此存活。他們卻大大干犯我的安息日。 「因此我說，我要在曠野把我的憤怒傾倒在他們身上，滅絕他們。
EZEK|20|14|我這麼做是為了我名的緣故，免得我的名在列國眼中被褻瀆，因為在這些列國眼前我領了他們出來。
EZEK|20|15|並且我在曠野向他們起誓，必不領他們進入我所賜的流奶與蜜之地，就是全地中最美好之地；
EZEK|20|16|因為他們厭棄我的典章，不順從我的律例，干犯我的安息日，他們的心隨從自己的偶像。
EZEK|20|17|雖然如此，我的眼仍顧惜他們，不毀滅他們，不在曠野把他們滅絕淨盡。
EZEK|20|18|「我在曠野對他們的兒女說：『不要遵行你們祖先的律例，不要謹守他們的規條，也不要用他們的偶像玷污自己。
EZEK|20|19|我是耶和華─你們的上帝，你們要順從我的律例，謹守遵行我的典章，
EZEK|20|20|且以我的安息日為聖。這日必在我與你們中間作記號，使你們知道我是耶和華─你們的上帝。』
EZEK|20|21|只是他們的兒女悖逆我，不順從我的律例，也不謹守遵行我的典章；人若遵行就必因此存活。他們卻干犯我的安息日。 「因此我說，我要在曠野把我的憤怒傾倒在他們身上，向他們發盡我的怒氣。
EZEK|20|22|但我卻縮手而未如此行；我這麼做是為了我名的緣故，免得我的名在列國眼中被褻瀆，因為在這些列國眼前我領了他們出來。
EZEK|20|23|並且我在曠野向他們起誓，要把他們驅散到列國，分散在列邦；
EZEK|20|24|因為他們不遵行我的典章，厭棄我的律例，干犯我的安息日，眼目向著他們祖先的偶像。
EZEK|20|25|我也任他們遵行那無益的律例，隨從那不能使人存活的規條。
EZEK|20|26|他們使所有頭生的經火，我就任憑他們在這供物上玷污自己；我令他們驚恐，他們就知道我是耶和華。
EZEK|20|27|「人子啊，你要告訴 以色列 家，對他們說，主耶和華如此說：你們的祖先在背叛我的事上再次褻瀆了我；
EZEK|20|28|我領他們到我起誓應許賜給他們的地，他們看見各高岡、各茂密的樹，就在那裏獻祭，獻上惹我發怒的供物，也在那裏焚燒馨香的祭，獻澆酒祭。
EZEK|20|29|我就對他們說：你們去的那丘壇叫甚麼呢？它名叫 巴麻 ，直到今日。
EZEK|20|30|所以你要對 以色列 家說，主耶和華如此說：你們仍要照你們祖先所做的玷污自己嗎？還要照他們可憎的事行淫嗎？
EZEK|20|31|當你們獻上供物，使你們兒子經火的時候，你們仍用各樣的偶像玷污自己，直到今日。 以色列 家啊，我豈能讓你們求問呢？主耶和華說：我指著我的永生起誓，我必不讓你們求問。
EZEK|20|32|「你們說：『我們要像列國和列邦的宗族一樣，去事奉木頭與石頭。』你們所起的心意萬不能成就。」
EZEK|20|33|「主耶和華說：我指著我的永生起誓，我要作王，用大能的手和伸出的膀臂，並傾倒出來的憤怒治理你們。
EZEK|20|34|我必用大能的手和伸出的膀臂，並傾倒出來的憤怒，把你們從萬民中領出來，從被趕散到的列邦聚集你們。
EZEK|20|35|我必帶你們到萬民的曠野，在那裏當面審判你們。
EZEK|20|36|我怎樣在 埃及 地的曠野審判你們的祖先，也必照樣審判你們。這是主耶和華說的。
EZEK|20|37|我要使你們從杖下經過，按著約的拘束 帶領你們。
EZEK|20|38|我必從你們中間除盡叛逆和得罪我的人；我將他們從所寄居的地方領出來，他們卻不得進入 以色列 地，你們就知道我是耶和華。
EZEK|20|39|「你們， 以色列 家啊，主耶和華如此說：你們若不聽從我，從今以後就讓各人去事奉他的偶像吧，只是不可再以你們的供物和偶像褻瀆我的聖名。
EZEK|20|40|「在我的聖山，就是 以色列 高處的山， 以色列 全家，那地所有的人，都要在那裏事奉我。在那裏我悅納他們，並要你們獻供物和初熟的土產，以及一切的聖物。這是主耶和華說的。
EZEK|20|41|我把你們從萬民中領出來，從被趕散到的列邦聚集你們，那時我必悅納你們如同悅納馨香之祭，我要在列國眼前，在你們中間顯為聖。
EZEK|20|42|我領你們進入 以色列 地，就是我起誓應許賜給你們列祖之地，那時你們就知道我是耶和華。
EZEK|20|43|你們在那裏要追念那玷污自己的所作所為，又要因所行的一切惡事厭惡自己。
EZEK|20|44|以色列 家啊，我為我名的緣故，沒有照著你們的惡行和你們的敗壞對待你們；你們就知道我是耶和華。這是主耶和華說的。」
EZEK|20|45|耶和華的話臨到我，說：
EZEK|20|46|「人子啊，你要面向南方，向南方傳講 ，向 尼革夫 田野的樹林說預言。
EZEK|20|47|你要對 尼革夫 的樹林說，要聽耶和華的話。主耶和華如此說：看哪，我要在你那裏點火，燒滅你們中間所有的綠樹和枯樹，猛烈的火焰必不熄滅；從南到北，人的臉都被燒焦。
EZEK|20|48|凡血肉之軀都知道是我─耶和華點了火，這火必不熄滅。」
EZEK|20|49|於是我說：「唉！主耶和華啊，人都指著我說：他不是說比喻的人嗎？」
EZEK|21|1|耶和華的話臨到我，說：
EZEK|21|2|「人子啊，把你的臉正對著 耶路撒冷 ，對著聖所 傳講 ，向 以色列 地說預言。
EZEK|21|3|你要向 以色列 地說，耶和華如此說：看哪，我與你為敵，拔刀出鞘，把義人和惡人從你中間剪除。
EZEK|21|4|因為我要剪除你當中的義人和惡人，所以我的刀要出鞘，從南到北攻擊所有的血肉之軀；
EZEK|21|5|凡血肉之軀都知道我─耶和華已拔刀出鞘，刀必不再入鞘。
EZEK|21|6|你，人子啊，要嘆息，在他們眼前斷了腰，愁苦地嘆息。
EZEK|21|7|若有人對你說：『你為甚麼嘆息呢？』你就說：『因為有風聲傳來，人心惶惶，雙手發軟，精神衰敗，膝弱如水。看哪，它臨近了，一定會發生。』這是主耶和華說的。」
EZEK|21|8|耶和華的話臨到我，說：
EZEK|21|9|「人子啊，你要預言說，耶和華如此吩咐，你要說： 有刀，刀已磨快， 又擦亮了；
EZEK|21|10|磨快為要大大殺戮， 擦亮為要像閃電。 我們豈能快樂呢？ 它藐視我兒的權杖和一切的木頭 。
EZEK|21|11|它已經交給人擦亮，可以掌握使用；這刀已經磨快擦亮，好交在行殺戮的人手中。
EZEK|21|12|人子啊，你要呼喊哀號，因為這刀將臨到我的百姓，臨到 以色列 所有的領袖身上。他們和我的百姓都要交在刀下，所以你要捶胸 。
EZEK|21|13|因為這是一個考驗，若它藐視權杖，也不算一回事，又怎麼樣呢？這是主耶和華說的。」
EZEK|21|14|「人子啊，你要拍掌預言，使這刀三番兩次臨到；這是致人死傷的刀，就是包圍人，使人大受死傷的刀。
EZEK|21|15|我設立這恐嚇 的刀，攻擊他們一切的城門，為要使他們的心驚慌害怕，許多人因而跌倒。唉！它 造得像閃電，磨得尖利 ，要行殺戮。
EZEK|21|16|刀啊，要行動一致 ，向右邊，或指向左邊；面向哪方，就向哪方。
EZEK|21|17|我也要拍掌，使我的憤怒平息。這是我─耶和華說的。」
EZEK|21|18|耶和華的話臨到我，說：
EZEK|21|19|「人子啊，你要畫定兩條路線，使 巴比倫 王的刀過來，這兩條路必從同一地分出來；要在通往城裏的路口畫手作指標。
EZEK|21|20|你要劃定一條路，使刀來到 亞捫 人的 拉巴 ，來到 猶大 ，在堅固城 耶路撒冷 。
EZEK|21|21|因為 巴比倫 王站在岔路上，在兩條路口占卜。他搖籤 求問神像，察看肝臟；
EZEK|21|22|右手是 耶路撒冷 的占卜，以便安設撞城槌，張口喊殺 ，揚聲呼叫，建土堆，築堡壘，以撞城槌攻打城門。
EZEK|21|23|在那些曾鄭重起誓的 猶大 人眼中，這是虛假的占卜；但 巴比倫 王要使他們想起自己的罪孽，以便俘擄他們。」
EZEK|21|24|於是，主耶和華如此說：「因你們的過犯顯露，你們的罪孽被記得，以致你們的罪惡在你們一切的行為上都彰顯出來；你們既被記得，就被擄在掌中。
EZEK|21|25|你這褻瀆行惡的 以色列 王啊，你的日子，最後懲罰的時刻已來臨。
EZEK|21|26|主耶和華如此說：當除掉榮冕，摘下華冠，景況已不復從前；要使卑者升為高，使高者降為卑。
EZEK|21|27|我要將這國傾覆，傾覆，再傾覆；這國必不存在，直等到那應得的人來到，我就將國賜給他。」
EZEK|21|28|「人子啊，你要說預言；你要說，論到 亞捫 人和他們的凌辱，主耶和華吩咐我如此說：有刀，拔出來的刀，已經擦亮，為了行殺戮；它亮如閃電以行吞滅。
EZEK|21|29|他們為你見虛假的異象，行謊詐的占卜，使你倒在褻瀆之惡人的頸項上；他們的日子，最後懲罰的時刻已來臨。
EZEK|21|30|你收刀入鞘吧！我要在你受造之處、生長之地懲罰你。
EZEK|21|31|我要把我的憤怒傾倒在你身上，把我烈怒的火噴在你身上；又將你交在善於殺滅、畜牲一般的人手中。
EZEK|21|32|你要成為火中之柴，你的血必在地裏；你必不再被記得，因為這是我─耶和華說的。」
EZEK|22|1|耶和華的話臨到我，說：
EZEK|22|2|「你，人子啊，你要審問，審問這流人血的城嗎？要使它知道它一切可憎的事。
EZEK|22|3|你要說，主耶和華如此說：那在其中流人血的城啊，它的時刻已到，它製造偶像玷污了自己。
EZEK|22|4|你因流了人的血，算為有罪；因所製造的偶像，玷污自己；你使你的日子臨近，你的年數已來到 。所以我使你承受列國的凌辱和列邦的譏誚。
EZEK|22|5|你這惡名昭彰、混亂的城啊，離你或遠或近的國家都必譏誚你。
EZEK|22|6|「看哪， 以色列 的領袖在你那裏，為了流人的血各逞其能。
EZEK|22|7|你那裏有輕慢父母的，在你當中有欺壓寄居者的，你那裏也有虧負孤兒寡婦的。
EZEK|22|8|你藐視我的聖物，干犯我的安息日。
EZEK|22|9|你那裏有為流人血而毀謗人的，你那裏有在山上吃祭物的，在你當中也有行淫亂的，
EZEK|22|10|有露父親下體的 ，有玷辱經期中不潔淨之婦人的。
EZEK|22|11|這人與鄰舍的妻子行可憎的事，那人行淫污辱媳婦，在你那裏還有人污辱他的姊妹，父親的女兒。
EZEK|22|12|你那裏有收取報酬而流人血的。你取利息，又索取高利；欺壓鄰舍，奪取財物；你竟然忘了我。這是主耶和華說的。
EZEK|22|13|「看哪，我因你所得不義之財和你們中間所流的血，就擊打手掌。
EZEK|22|14|到了我對付你的日子，你的心豈能忍受呢？你的手還能有力嗎？我─耶和華說了這話，就必成就。
EZEK|22|15|我要把你驅散到列國，分散在列邦。我也必除掉你們中間的污穢。
EZEK|22|16|你在列國眼前因自己所做的被侮辱 ，你就知道我是耶和華。」
EZEK|22|17|耶和華的話臨到我，說：
EZEK|22|18|「人子啊，我看 以色列 家為渣滓。他們是爐中的銅、錫、鐵、鉛，是煉銀的渣滓 。
EZEK|22|19|所以主耶和華如此說：因你們全都成為渣滓，所以，看哪，我必將你們聚集在 耶路撒冷 中。
EZEK|22|20|人怎樣把銀、銅、鐵、鉛、錫聚在爐中，吹火使它鎔化；照樣，我也要在我的怒氣和憤怒中聚集你們，把你們安置在城中，使你們鎔化。
EZEK|22|21|我必聚集你們，把我烈怒的火吹在你們身上，你們就在其中鎔化。
EZEK|22|22|銀子怎樣在爐中鎔化，你們也必照樣在城中鎔化，因此就知道是我─耶和華把憤怒傾倒在你們身上。」
EZEK|22|23|耶和華的話臨到我，說：
EZEK|22|24|「人子啊，你要向這地說：你是未被潔淨 之地，在我盛怒的日子，沒有雨水在其上。
EZEK|22|25|其中的先知同謀背叛 ，如咆哮的獅子抓撕掠物。他們吞滅人命，搶奪財寶，使這地寡婦增多。
EZEK|22|26|其中的祭司曲解我的律法，褻瀆我的聖物，不分別聖與俗，也不使人分辨潔淨和不潔淨，又遮眼不顧我的安息日；在他們中間連我也被褻慢了。
EZEK|22|27|其中的領袖彷彿野狼抓撕掠物，流人的血，傷害人命，為得不義之財。
EZEK|22|28|其中的先知為他們粉刷，見虛假的異象，行謊詐的占卜，說：『主耶和華如此說』，其實耶和華並沒有說。
EZEK|22|29|這地的百姓慣行欺壓搶奪之事，虧負困苦和貧窮的人，欺壓寄居者，沒有公平。
EZEK|22|30|我在他們中間尋找一人重修城牆，在我面前為這地站在缺口上，使我不致滅絕它，卻連一個也找不著。
EZEK|22|31|所以我把憤怒傾倒在他們身上，用烈怒之火消滅他們，照他們所做的報應在他們頭上。這是主耶和華說的。」
EZEK|23|1|耶和華的話臨到我，說：
EZEK|23|2|「人子啊，有兩個女子，是一母所生，
EZEK|23|3|她們在 埃及 行淫，年少時就開始行淫；在那裏任人擁抱胸懷，撫弄她們少女的乳房。
EZEK|23|4|她們的名字，大的叫 阿荷拉 ，妹妹叫 阿荷利巴 。她們都歸於我，生了兒女。論到她們的名字， 阿荷拉 是 撒瑪利亞 ， 阿荷利巴 是 耶路撒冷 。
EZEK|23|5|「 阿荷拉 歸我之後卻仍行淫，戀慕所愛的人，就是 亞述 人，都是戰士 ，
EZEK|23|6|穿著藍衣，作省長、副省長，全都是俊美的年輕人，騎著馬的騎士。
EZEK|23|7|阿荷拉 與 亞述 人中所有的美男子放縱淫行，她因拜所戀慕之人的一切偶像，玷污了自己。
EZEK|23|8|她從 埃及 的時候，就沒有離開過淫亂；因為她年輕時，有人與她同寢，撫弄她少女的乳房，和她縱慾行淫。
EZEK|23|9|因此，我把她交在她所愛的人手中，就是她所戀慕的 亞述 人手中。
EZEK|23|10|他們暴露她的下體，擄掠她的兒女，用刀殺了她；他們向她施行審判，使她在婦女中留下臭名。
EZEK|23|11|「她妹妹 阿荷利巴 雖然看見了，卻還是縱慾，比姊姊更加腐敗，行淫亂比姊姊更甚。
EZEK|23|12|她戀慕 亞述 人，就是省長和副省長，披掛整齊的戰士，騎著馬的騎士，全都是俊美的年輕人。
EZEK|23|13|我看見她被污辱，姊妹二人同行一路。
EZEK|23|14|阿荷利巴 又加增淫行，她看見牆上刻有人像，就是鮮紅色的 迦勒底 人雕刻的像。
EZEK|23|15|它們腰間繫著帶子，頭上有飄揚的裹頭巾，都是將軍的樣子， 巴比倫 人的形像； 迦勒底 是他們的出生地。
EZEK|23|16|阿荷利巴 一看見就戀慕他們，派遣使者往 迦勒底 他們那裏去。
EZEK|23|17|巴比倫 人來到她那裏，上了她愛情的床，與她行淫污辱她。她被污辱，隨後她的心卻與他們生疏。
EZEK|23|18|這樣，她既暴露淫行，暴露下體；我的心就與她生疏，像先前與她的姊姊生疏一樣。
EZEK|23|19|她仍繼續增添淫行，追念她年輕時在 埃及 地行淫的日子，
EZEK|23|20|戀慕情人的身壯精足，如驢似馬。
EZEK|23|21|這樣，你就渴望年輕時的淫蕩；那時， 埃及 人因你年輕時的胸懷，撫弄你的乳房 。」
EZEK|23|22|阿荷利巴 啊，主耶和華如此說：「看哪，我要激起先前你喜愛，而後生疏的人前來攻擊你。我必使他們前來，在你四圍攻擊你；
EZEK|23|23|有 巴比倫 人、 迦勒底 眾人、 比割 人、 書亞 人、 哥亞 人，還有 亞述 眾人與他們一起，都是俊美的年輕人。他們是省長、副省長、將軍、有名聲的，全都騎著馬。
EZEK|23|24|他們用兵器、 戰車、輜重車，率領大軍前來攻擊你。他們要拿大小盾牌，戴著頭盔，在你四圍擺陣攻擊你。我要把審判交給他們，他們必按著自己的規條審判你。
EZEK|23|25|我要向你傾洩我的妒忌，使他們以憤怒對待你。他們必割去你的鼻子和耳朵，你剩餘的人必倒在刀下。他們必擄去你的兒女，你所剩餘的必被火焚燒。
EZEK|23|26|他們必剝去你的衣服，奪取你美麗的寶物。
EZEK|23|27|這樣，我必止息你的淫行和你從 埃及 地就開始犯的淫亂，使你不再仰望 亞述 ，也不再追念 埃及 。
EZEK|23|28|主耶和華如此說：看哪，我必把你交在你所恨惡的人手中，就是你心與他生疏的人手中。
EZEK|23|29|他們要以恨惡對待你，奪取你勞碌得來的一切，留下你赤身露體。你淫亂的下體，連你的淫行和淫蕩，都必顯露。
EZEK|23|30|人必向你行這些事；因為你隨從外邦人行淫，用他們的偶像玷污自己。
EZEK|23|31|你走了你姊姊的路，所以我必把她的杯交在你的手中。」
EZEK|23|32|主耶和華如此說： 「你必喝你姊姊的杯， 那杯又深又廣， 盛得很多， 使你遭受嗤笑譏刺。
EZEK|23|33|你必酩酊大醉， 滿有愁苦。 你姊姊 撒瑪利亞 的杯， 驚駭和淒涼的杯，
EZEK|23|34|你必喝它，並且喝乾。 甚至咀嚼杯片， 撕裂自己的胸脯； 因為我曾說過。 這是主耶和華說的。」
EZEK|23|35|主耶和華如此說：「因你忘記我，將我丟在背後，所以你要擔當你的淫行和淫蕩。」
EZEK|23|36|耶和華對我說：「人子啊，你要審問 阿荷拉 與 阿荷利巴 嗎？要指出她們所做可憎的事。
EZEK|23|37|她們行姦淫，手中有血。她們與偶像行姦淫，使她們為我所生的兒女經火，給它們當食物。
EZEK|23|38|此外，她們還向我這樣做：同一天又玷污我的聖所，干犯我的安息日。
EZEK|23|39|她們殺了兒女獻給偶像，當天又進入我的聖所，褻瀆了它。看哪，這就是她們在我殿中所做的。
EZEK|23|40|「況且你們兩姊妹派人從遠方召人來。使者到了他們那裏，看哪，他們就來了。為了他們，你們沐浴，畫眼影，佩戴首飾，
EZEK|23|41|坐在華美的床上，前面擺設桌子，把我的香料和膏油放在其上。
EZEK|23|42|在那裏有一群人歡樂的聲音；有許多的平民，從曠野來的醉漢 ，把鐲子戴在她們手上，把華冠戴在她們頭上。
EZEK|23|43|「我論到這久行姦淫而色衰的婦人說：現在人們還要與她行淫，她也要與人行淫。
EZEK|23|44|人去到 阿荷拉 和 阿荷利巴 二淫婦那裏 ，好像與妓女行淫。
EZEK|23|45|義人必按照審判淫婦和流人血之婦人的規條，審判她們；因為她們是淫婦，她們的手中有血。」
EZEK|23|46|主耶和華如此說：「我要讓軍隊上來攻擊她們，使她們驚駭，成為擄物。
EZEK|23|47|這軍隊必用石頭打死她們，用刀劍殺害她們，又殺戮她們的兒女，用火焚燒她們的房屋。
EZEK|23|48|我必使這地不再有淫行，所有的婦女都受警戒，不再效法你們的淫行 。
EZEK|23|49|人必因你們的淫行報應你們；你們要擔當拜偶像的罪，因此你們就知道我是主耶和華。」
EZEK|24|1|第九年十月初十，耶和華的話臨到我，說：
EZEK|24|2|「人子啊，你要記錄這一天的名稱，這特別的一天， 巴比倫 王圍困 耶路撒冷 ，就在這特別的一天。
EZEK|24|3|你要向這悖逆之家設比喻，對他們說，主耶和華如此說： 把鍋放在火上， 放好了，倒水在其中；
EZEK|24|4|要將肉塊，一切肥美的肉塊， 腿和肩都放在鍋裏， 要裝滿上等的骨頭；
EZEK|24|5|要取羊群中最好的， 把柴 堆在下面， 把它煮開， 骨頭煮在其中。
EZEK|24|6|「主耶和華如此說：禍哉！這流人血的城，就是長銹的鍋。它的銹未曾除掉，要將肉塊從其中一一取出，不必抽籤。
EZEK|24|7|這城所流的血還在城中，血倒在光滑的磐石上，沒有倒在地上，用土掩蓋；
EZEK|24|8|是我使這城所流的血倒在光滑的磐石上，不得掩蓋，為要惹動憤怒，施行報應。
EZEK|24|9|所以主耶和華如此說：禍哉！這流人血的城，我必親自加大柴堆。
EZEK|24|10|你要添上木柴，使火著旺，將肉煮爛，加上香料 ，烤焦骨頭；
EZEK|24|11|你要把空鍋放在炭火上，將鍋燒熱，把銅燒紅，鎔化其中的污穢，除淨其上的銹。
EZEK|24|12|然而這一切勞碌無效 ，它厚厚的銹，即使用火也除不掉。
EZEK|24|13|雖然我想潔淨你污穢的淫行，你卻不潔淨，你的污穢再也不能潔淨，直等我止息了向你發的憤怒。
EZEK|24|14|我─耶和華說了這話，時候到了，就必成就；必不退縮，不顧惜，也不憐憫。人必照你的所作所為審判你。這是主耶和華說的。」
EZEK|24|15|耶和華的話臨到我，說：
EZEK|24|16|「人子，看哪，我要以災病奪取你眼中所喜愛的，你卻不可悲哀哭泣，也不可流淚，
EZEK|24|17|只可嘆息，不可出聲，不可辦理喪事；裹上頭巾，腳上穿鞋，不可摀著鬍鬚，也不可吃一般人的食物 。」
EZEK|24|18|到了早晨我把這事告訴百姓，晚上我的妻子就死了。次日早晨我就遵命而行。
EZEK|24|19|百姓對我說：「你這樣做跟我們有甚麼關係，你不告訴我們嗎？」
EZEK|24|20|我對他們說：「耶和華的話臨到我，說：
EZEK|24|21|『你告訴 以色列 家，主耶和華如此說：我要使我的聖所被褻瀆，就是你們憑勢力所誇耀、眼裏所喜愛、心中所愛惜的；並且你們所遺留的兒女必倒在刀下。
EZEK|24|22|那時，你們要照我所做的去做。你們不可摀著鬍鬚，也不可吃一般人的食物。
EZEK|24|23|你們頭要裹上頭巾，腳要穿上鞋；不可悲哀哭泣。你們必因自己的罪孽衰殘，相對嘆息。
EZEK|24|24|以西結 必這樣成為你們的預兆；凡他所做的，你們也必照樣做。那事來到，你們就知道我是主耶和華。』」
EZEK|24|25|「你，人子啊，那日當我除掉他們所倚靠的保障、所歡喜的榮耀，並眼中所喜愛的，心裏所重看的兒女時，
EZEK|24|26|逃脫的人豈不來到你這裏，使你耳聞這事嗎？
EZEK|24|27|那日你要向逃脫的人開口說話，不再啞口無言。你必這樣成為他們的預兆，他們就知道我是耶和華。」
EZEK|25|1|耶和華的話臨到我，說：
EZEK|25|2|「人子啊，你要面向 亞捫 人說預言，攻擊他們。
EZEK|25|3|你要對 亞捫 人說，當聽主耶和華的話。主耶和華如此說：我的聖所遭褻瀆， 以色列 地變荒涼， 猶大 家被擄掠；那時，你因這些事說『啊哈』，
EZEK|25|4|所以，看哪，我要把你交給東方人為業；他們必在你中間安營居住，設立居所，吃你的果子，喝你的奶。
EZEK|25|5|我必使 拉巴 成為牧放駱駝之地，使 亞捫 成為羊群躺臥之處，你們就知道我是耶和華。
EZEK|25|6|主耶和華如此說：因你們拍手頓足，幸災樂禍，藐視 以色列 地，
EZEK|25|7|所以，看哪，我要伸手攻擊你，把你交給列國作為擄物。我必從萬民中剪除你，從列邦中消滅你。我必除滅你，你就知道我是耶和華。」
EZEK|25|8|「主耶和華如此說：因 摩押 和 西珥 人說『看哪， 猶大 家與列國無異』，
EZEK|25|9|所以，看哪，我要破開 摩押 邊界的城鎮，就是 摩押 人所誇耀的城鎮， 伯‧耶施末 、 巴力‧免 、 基列亭 ，
EZEK|25|10|令東方人前來攻擊 亞捫 人。我必將 亞捫 交給他們為業，使 亞捫 人在列國中不再被記念。
EZEK|25|11|我也必向 摩押 施行審判，他們就知道我是耶和華。」
EZEK|25|12|「主耶和華如此說：因為 以東 向 猶大 家報仇，因向他們報仇而大大顯為有罪，
EZEK|25|13|所以主耶和華如此說：我要伸手攻擊 以東 ，將人與牲畜剪除，使 以東 從 提幔 起，直到 底但 ，地變荒涼，人也都倒在刀下。
EZEK|25|14|我要藉我子民 以色列 的手報復 以東 ；他們必照我的怒氣，按我的憤怒對待 以東 ， 以東 人就知道施報的是我。這是主耶和華說的。」
EZEK|25|15|「主耶和華如此說：因 非利士 人報仇，就是心存輕蔑報仇；他們永懷仇恨，意圖毀滅，
EZEK|25|16|所以主耶和華如此說：看哪，我要伸手攻擊 非利士 人，剪除 基利提 人，滅絕沿海剩餘的居民。
EZEK|25|17|我要大大報復他們，發怒斥責他們。我報復他們的時候，他們就知道我是耶和華。」
EZEK|26|1|第十一年某月初一，耶和華的話臨到我，說：
EZEK|26|2|「人子啊，因 推羅 向 耶路撒冷 說：『啊哈！那眾民之門已經破壞，向我敞開；它既變為廢墟，我必豐盛。』
EZEK|26|3|所以，主耶和華如此說： 推羅 ，看哪，我與你為敵，使許多國家湧上攻擊你，如同海洋使波浪湧上一樣。
EZEK|26|4|他們要破壞 推羅 的城牆，拆毀它的城樓。我也要刮淨它的塵土，使它成為光滑的磐石。
EZEK|26|5|推羅 必成為海中的曬網場，因為我曾說過， 這是主耶和華說的。它必成為列國的擄物，
EZEK|26|6|推羅 鄉間鄰近的城鎮 必遭刀劍滅絕，他們就知道我是耶和華。」
EZEK|26|7|主耶和華如此說：「看哪，我必使諸王之王，就是 巴比倫 王 尼布甲尼撒 ，率領馬匹、戰車、騎兵、軍隊和許多人從北方來攻擊 推羅 。
EZEK|26|8|他必用刀劍殺滅你鄉間鄰近的城鎮，也必築堡壘，建土堆，舉盾牌攻擊你。
EZEK|26|9|他要安設撞城槌攻破你的城牆，以刀劍拆毀你的城樓。
EZEK|26|10|因他馬匹眾多，塵土必揚起遮蔽你。他進入你的城門，如同進入已有缺口之城。那時，你的城牆必因騎兵、車輪和戰車的響聲震動。
EZEK|26|11|他的馬蹄必踐踏你所有的街道；他必用刀劍殺戮你的居民。你堅固的柱子 必倒在地上。
EZEK|26|12|人必擄獲你的財寶，掠奪你的貨財；他們要破壞你的城牆，拆毀你華美的房屋，將你的石頭、木頭、塵土都拋在水中。
EZEK|26|13|我要使你唱歌的聲音止息；人不再聽見你彈琴的聲音。
EZEK|26|14|我必使你成為光滑的磐石，作曬網的場所。你不得再被建造，因為我─耶和華已這樣說了。這是主耶和華說的。」
EZEK|26|15|主耶和華對 推羅 如此說：「在你中間行殺戮，受傷的人唉哼時，海島豈不都因你傾倒的響聲震動嗎？
EZEK|26|16|那時沿海的君王都要從寶座下來，除去朝服，脫下錦衣，披上戰兢，坐在地上，不停發抖，為你而驚駭。
EZEK|26|17|他們必為你作哀歌，向你說： 『你這聞名之城， 航海之人居住， 海上最為堅固的， 你和居民使所有住在沿海的人 無不驚恐， 現在竟然毀滅了！
EZEK|26|18|如今在你傾覆的日子， 海島都要戰兢； 海中的群島見你歸於無有 就都驚惶。』」
EZEK|26|19|主耶和華如此說：「 推羅 啊 ，我要使你變為荒涼，如無人居住的城鎮；又使深水漫過你，大水淹沒你。
EZEK|26|20|那時，我要使你和下到地府的人同去，到古時候的人那裏；我要使你和下到地府的人一同住在地的深處，在久已荒廢的地方，使你那裏不再有人居住；我要在活人之地顯榮耀 。
EZEK|26|21|我必叫你令人驚恐，使你不再存留於世；人雖尋找你，卻永不尋見。這是主耶和華說的。」
EZEK|27|1|耶和華的話臨到我，說：
EZEK|27|2|「人子啊，要為 推羅 作哀歌。
EZEK|27|3|你要對位於海口，跟許多海島的百姓做生意的 推羅 說，主耶和華如此說： 推羅 啊，你曾說： 『我全然美麗。』
EZEK|27|4|你的疆界在海的中心， 造你的使你全然美麗。
EZEK|27|5|他們用 示尼珥 的松樹作你的甲板， 用 黎巴嫩 的香柏樹作桅杆，
EZEK|27|6|用 巴珊 的橡樹作你的槳， 用鑲嵌象牙的 基提 海島黃楊木 為艙板。
EZEK|27|7|你的帆是用 埃及 繡花細麻布做的， 可作你的大旗； 你的篷是用 以利沙島 的藍色和紫色布做的。
EZEK|27|8|西頓 和 亞發 的居民為你划槳； 推羅 啊，你們中間的智慧人為你掌舵。
EZEK|27|9|迦巴勒 的長者和智者 在你中間修補裂縫； 海上一切的船隻和水手 都在你那裏進行貨物交易。
EZEK|27|10|「 波斯 人、 路德 人、 弗 人在你的軍營中作戰士；他們在你們中間懸掛盾牌和頭盔，彰顯你的尊榮。
EZEK|27|11|亞發 人和你的軍隊都駐守在四圍的城牆上，你的城樓上也有勇士；他們懸掛盾牌，成全你的美麗。
EZEK|27|12|「 他施 因你多有財物，就作你的客商，他們帶著銀、鐵、錫、鉛前來換你的商品。
EZEK|27|13|雅完 、 土巴 、 米設 都與你交易，以人口和銅器換你的貨物。
EZEK|27|14|陀迦瑪 族用馬匹、戰馬和騾子換你的商品。
EZEK|27|15|底但 人與你交易，許多海島成為你的碼頭；他們拿象牙、黑檀木與你交換。
EZEK|27|16|亞蘭 因你貨品充裕，就作你的客商；他們用綠寶石、紫色布、刺繡、細麻布、珊瑚、紅寶石換你的商品。
EZEK|27|17|猶大 和 以色列 地都與你交易；他們用 米匿 的小麥、餅、蜜、油、乳香換你的貨物。
EZEK|27|18|大馬士革 也因你貨品充裕，多有各類財物，就帶來 黑本 酒和白羊毛與你交易。
EZEK|27|19|威但 和從 烏薩 來的 雅完 人 為了你的貨物，以加工的鐵、桂皮、香菖蒲換你的商品。
EZEK|27|20|底但 以騎馬用的座墊毯子與你交換。
EZEK|27|21|阿拉伯 和 基達 所有的領袖都作你的客商，用羔羊、公綿羊、公山羊與你交換。
EZEK|27|22|示巴 和 拉瑪 的商人也來與你交易，他們用各類上好的香料、各類的寶石和黃金換你的商品。
EZEK|27|23|哈蘭 、 干尼 、 伊甸 、 示巴 商人、 亞述 和 基抹 都與你交易。
EZEK|27|24|這些商人將美好的貨物包在藍色的繡花包袱內，又將華麗的衣服裝在香柏木的箱子裏，用繩索捆著，以此與你交易 。
EZEK|27|25|他施 的船隻為你運貨， 你在海中滿載貨物，極其沉重。
EZEK|27|26|划槳的把你划到水深之處， 東風在海中將你擊破。
EZEK|27|27|你的財寶、商品、貨物、 水手、掌舵的、 修補船縫的、進行貨物交易的， 並你那裏所有的戰士 和你中間所有的軍隊， 在你傾覆的日子都必沉在海底。
EZEK|27|28|因掌舵者的呼聲， 郊野就必震動。
EZEK|27|29|所有划槳的 都從他們的船下來； 水手和所有在海上掌舵的， 都要登岸。
EZEK|27|30|他們必為你放聲痛哭， 撒塵土於頭上， 在灰中打滾；
EZEK|27|31|又為你使頭光禿， 用麻布束腰， 號咷痛哭， 痛苦至極。
EZEK|27|32|他們哀號的時候， 為你作哀歌， 為你痛哭： 有何城如 推羅 ， 在海中沉寂呢？
EZEK|27|33|你由海上運出商品， 使許多民族充裕； 你以許多財寶貨物 令地上的君王豐富。
EZEK|27|34|在深水中被海浪打破的時候， 你的貨物和你中間所有的軍隊都下沉。
EZEK|27|35|海島所有的居民為你驚奇， 他們的君王都甚恐慌，面帶愁容。
EZEK|27|36|萬民中的商人向你發噓聲； 你令人驚恐， 不再存留於世，直到永遠。」
EZEK|28|1|耶和華的話臨到我，說：
EZEK|28|2|「人子啊，你要對 推羅 的君王說，主耶和華如此說： 你心裏高傲，說：『我是神明； 我在海中坐諸神之位。』 雖然你把你的心比作神明的心， 你卻不過是人，並不是神明！
EZEK|28|3|看哪，你比 但以理 更有智慧， 任何祕密都不能向你隱藏。
EZEK|28|4|你靠自己的智慧聰明得了財寶， 把金銀收入庫房；
EZEK|28|5|你靠自己的大智慧以貿易增添財寶， 又因你的財寶心裏高傲；
EZEK|28|6|所以主耶和華如此說： 因你把你的心比作神明的心，
EZEK|28|7|所以，看哪，我必使外國人， 就是列國中兇暴的人臨到你這裏； 他們要拔刀摧毀你用智慧得來的美物， 污損你的榮光。
EZEK|28|8|他們必使你墜入地府； 你要像被刺殺之人的死，死在海中。
EZEK|28|9|在殺你的人面前， 你還能說『我是神明』嗎？ 在殺害你的人手中， 你不過是人，並不是神明。
EZEK|28|10|你要死在陌生人手中， 像未受割禮之人的死， 因為我曾說過， 這是主耶和華說的。」
EZEK|28|11|耶和華的話臨到我，說：
EZEK|28|12|「人子啊，要為 推羅 王作哀歌，對他說，主耶和華如此說： 你曾是完美的典範， 智慧充足，全然美麗。
EZEK|28|13|你在 伊甸 ─上帝的園中， 佩戴各樣寶石， 就是紅寶石、紅璧璽、金剛石、 水蒼玉、紅瑪瑙、碧玉、 藍寶石、綠寶石、紅玉； 你的寶石有黃金的底座，手工精巧 ， 都是在你受造之日預備的。
EZEK|28|14|我指定你為受膏的基路伯， 看守保護； 你在上帝的聖山上； 往來在如火的寶石中。
EZEK|28|15|你從受造之日起行為正直， 直到後來查出你的不義。
EZEK|28|16|你因貿易發達， 暴力充斥其中，以致犯罪， 所以我污辱你，使你離開上帝的山。 守護者基路伯啊， 我已將你從如火的寶石中殲滅。
EZEK|28|17|你因美麗心中高傲， 因榮光而敗壞智慧， 我已將你拋棄在地， 把你擺在君王面前， 好叫他們目睹眼見。
EZEK|28|18|你因罪孽眾多，貿易不公， 褻瀆了你的聖所； 因此我使火從你中間發出， 燒滅了你， 使你在所有觀看的人眼前 變為地上的灰燼。
EZEK|28|19|萬民中凡認識你的 都必為你驚奇。 你令人驚恐， 不再存留於世，直到永遠。」
EZEK|28|20|耶和華的話臨到我，說：
EZEK|28|21|「人子啊，你要面向 西頓 ，向它說預言。
EZEK|28|22|你要說，主耶和華如此說： 『 西頓 ，看哪，我與你為敵， 我要在你中間得榮耀。』 我在它中間施行審判、顯為聖的時候， 人就知道我是耶和華。
EZEK|28|23|我必令瘟疫進入 西頓 ， 使血流在街上。 刀劍從四圍臨到它， 被殺的要仆倒在其中； 人就知道我是耶和華。」
EZEK|28|24|「四圍恨惡 以色列 家的人，對他們必不再如刺人的荊棘，傷人的蒺藜；他們就知道我是主耶和華。」
EZEK|28|25|主耶和華如此說：「我將分散在萬民中的 以色列 家召集回來，在列國眼前向他們顯為聖的時候，他們仍可在我所賜給我僕人 雅各 之地居住。
EZEK|28|26|他們要在這地上安然居住。我向四圍恨惡他們的眾人施行審判之後，他們要建造房屋，栽葡萄園，安然居住，他們就知道我是耶和華─他們的上帝。」
EZEK|29|1|第十年十月十二日，耶和華的話臨到我，說：
EZEK|29|2|「人子啊，你要面向 埃及 王法老，向他和 埃及 全地說預言。
EZEK|29|3|你要說，主耶和華如此說： 埃及 王法老， 你這臥在自己江河中的海怪， 看哪，我與你為敵。 你曾說：『我的 尼羅河 是我的， 是我為自己造的。』
EZEK|29|4|我必用鉤子鉤住你的腮頰， 令江河中的魚貼住你的鱗甲； 我要把你和所有貼著鱗甲的魚 從你的江河中拉上來。
EZEK|29|5|我要把你和江河中的魚全都拋棄在曠野； 你必仆倒在田間， 無人收殮，無人掩埋。 我已將你給了地上的走獸、空中的飛鳥作食物。
EZEK|29|6|「 埃及 所有的居民必定知道我是耶和華。因為你已成為 以色列 家蘆葦的杖；
EZEK|29|7|他們用手掌一握，你就斷裂，傷了他們的肩；他們靠著你，你卻折斷，閃了他們的腰 。
EZEK|29|8|所以主耶和華如此說：我必使刀劍臨到你，把人與牲畜從你中間剪除。
EZEK|29|9|埃及 地必荒蕪廢棄，他們就知道我是耶和華。 「因為法老說『 尼羅河 是我的，是我所造的』，
EZEK|29|10|所以，看哪，我必與你和你的江河為敵，使 埃及 地，從 密奪 到 色弗尼 ，直到 古實 邊界，全然廢棄荒蕪。
EZEK|29|11|人的腳不經過，獸的蹄也不經過，四十年之久無人居住。
EZEK|29|12|我要使 埃及 地成為荒蕪中最荒蕪的地，使它的城鎮變為荒廢中最荒廢的城鎮，共四十年之久。我必將 埃及 人分散到列國，四散在列邦。
EZEK|29|13|「主耶和華如此說：滿了四十年後，我必招聚分散在萬民中的 埃及 人。
EZEK|29|14|我要令 埃及 被擄的人歸回，使他們回到本地 巴特羅 。在那裏，他們必成為弱小的國家，
EZEK|29|15|成為列國中最低微的，不再自高於列邦之上。我必使他們變為小國，不再轄制列邦。
EZEK|29|16|埃及 必不再作 以色列 家的倚靠，卻使 以色列 家想起他們仰賴 埃及 的罪。他們就知道我是主耶和華。」
EZEK|29|17|第二十七年正月初一，耶和華的話臨到我，說：
EZEK|29|18|「人子啊， 巴比倫 王 尼布甲尼撒 令他的軍兵大力攻打 推羅 ，以致頭都光禿，肩都磨破；然而他和軍兵雖然為攻打 推羅 花這麼多力氣，卻沒有從那裏得到甚麼犒賞。
EZEK|29|19|所以主耶和華如此說：我要將 埃及 地賜給 巴比倫 王 尼布甲尼撒 ；他必擄掠 埃及 的財富，搶奪它的擄物，擄掠它的掠物，用以犒賞他的軍兵。
EZEK|29|20|我將 埃及 地賜給他，犒賞他，因他們為我效勞。這是主耶和華說的。
EZEK|29|21|「當那日，我必使 以色列 家壯大 ，又必使你─ 以西結 在他們中間開口；他們就知道我是耶和華。」
EZEK|30|1|耶和華的話臨到我，說：
EZEK|30|2|「人子啊，你要說預言；你要說，主耶和華如此說： 哀哉這日！你們應當哭號，
EZEK|30|3|因為日子近了， 耶和華的日子臨近了； 那是密雲之日， 是列國受罰 之期。
EZEK|30|4|必有刀劍臨到 埃及 ； 被殺的人仆倒在 埃及 時， 古實 人顫驚不已。 埃及 的財富遭擄掠， 根基被拆毀。
EZEK|30|5|古實 人、 弗 人、 路德 人、混居的各族和 古伯 人，以及盟國的人都要與 埃及 人一同倒在刀下。」
EZEK|30|6|耶和華如此說： 扶助 埃及 的必傾倒， 埃及 驕傲的權勢必降為卑， 從 密奪 到 色弗尼 ，人必倒在刀下。 這是主耶和華說的。
EZEK|30|7|埃及 成為荒涼中最荒涼的國， 它的城鎮變為荒廢中最荒廢的城鎮。
EZEK|30|8|我在 埃及 放火， 幫助 埃及 的，都遭滅絕； 那時，他們就知道我是耶和華。
EZEK|30|9|「到那日，必有使者從我面前乘船出去，使安逸無慮的 古實 人驚懼；當 埃及 遭難的日子，痛苦也必臨到他們。看哪，這事臨近了！
EZEK|30|10|主耶和華如此說： 我要藉 巴比倫 王 尼布甲尼撒 的手 除滅 埃及 的軍隊。
EZEK|30|11|他和隨從他的人， 就是列國中兇暴的人， 要前來毀滅這地， 拔刀攻擊 埃及 ， 使遍地佈滿被殺的人。
EZEK|30|12|我要使江河乾涸， 將這地賣在惡人手中； 我要藉外國人的手， 使這地和其中所充滿的變為荒蕪； 這是我─耶和華說的。
EZEK|30|13|「主耶和華如此說： 我要毀滅偶像， 從 挪弗 除掉神像； 不再有君王出自 埃及 地， 我要使 埃及 地的人懼怕。
EZEK|30|14|我必令 巴特羅 荒涼， 在 瑣安 放火， 向 挪 施行審判。
EZEK|30|15|我要將我的憤怒傾倒在 訓 ， 埃及 的堡壘上， 要剪除 挪 的眾民。
EZEK|30|16|我必在 埃及 放火， 訓 必大大痛苦， 挪 被攻破， 挪弗 終日遭敵侵襲。
EZEK|30|17|亞文 和 比‧伯實 的年輕人必倒在刀下， 這些城鎮將被擄掠。
EZEK|30|18|我在 答比匿 折斷 埃及 的軛 ， 使它驕傲的權勢止息。 那時，日光必退去； 至於這城，必有密雲遮蔽， 鄰近的城鎮 也遭擄掠。
EZEK|30|19|我要如此向 埃及 施行審判， 他們就知道我是耶和華。」
EZEK|30|20|第十一年正月初七，耶和華的話臨到我，說：
EZEK|30|21|「人子啊，我已折斷 埃及 王法老的一隻膀臂；看哪，無人為他敷藥，也無人為他包紮繃帶，使他有力持刀。
EZEK|30|22|因此，主耶和華如此說：看哪，我與 埃及 王法老為敵，要折斷他的膀臂，折斷強壯的和已受傷的，使刀從他手中掉落。
EZEK|30|23|我必將 埃及 人分散到列國，四散在列邦。
EZEK|30|24|我要使 巴比倫 王的膀臂有力，把我的刀交在他手中；卻要折斷法老的膀臂，使他在 巴比倫 王面前呻吟，如同被殺的人一樣。
EZEK|30|25|我要使 巴比倫 王的膀臂強壯，法老的膀臂卻要下垂；當我把我的刀交在 巴比倫 王手中時，他要舉刀攻擊 埃及 地，他們就知道我是耶和華。
EZEK|30|26|我必將 埃及 人分散到列國，四散在列邦；他們就知道我是耶和華。」
EZEK|31|1|第十一年三月初一，耶和華的話臨到我，說：
EZEK|31|2|「人子啊，你要對 埃及 王法老和他的軍隊說： 論到你的強盛，誰能與你相比呢？
EZEK|31|3|看哪， 亞述 是 黎巴嫩 的香柏樹， 枝條榮美，蔭密如林， 極其高大，樹頂高聳入雲。
EZEK|31|4|眾水使它生長， 深水使它長高； 所栽之地有江河環繞， 汊出的水道流至田野的樹木。
EZEK|31|5|所以它高大超過田野的樹木； 生長時因水源豐沛， 枝子繁多，枝條增長。
EZEK|31|6|空中所有的飛鳥在枝子上搭窩， 野地所有的走獸在枝條下生子， 所有的大國也在它的蔭下居住。
EZEK|31|7|它樹大枝長，極為榮美， 因它的根在眾水之旁。
EZEK|31|8|上帝園中的香柏樹不能遮蔽它； 松樹不及它的枝子， 楓樹不及它的枝條， 上帝園中的樹都沒有它榮美。
EZEK|31|9|我使它枝條繁多， 極為榮美； 在上帝的園中， 伊甸 所有的樹都嫉妒它。」
EZEK|31|10|所以主耶和華如此說：「因它 高大，樹頂高聳入雲，心高氣傲，
EZEK|31|11|我要把它交給 列國中強人的手裏，他們必定按它的罪惡懲治它。我已經驅逐它。
EZEK|31|12|外國人，就是列國中兇暴的人，已把它砍斷拋棄。它的枝條掉落山間和一切谷中，枝子折斷，落在地上一切河道。地上的萬民都離開它的遮蔭，拋棄了它。
EZEK|31|13|空中的飛鳥都棲身在掉落的樹幹上，野地的走獸也都躺臥在它的枝條中。
EZEK|31|14|為了要使水邊的樹木枝幹不再長高，樹頂也不再高聳入雲；那些得水滋潤的，不再屹立於其中。因為它們和下到地府的人一起，都被交與死亡，到了地底下。」
EZEK|31|15|主耶和華如此說：「它墜落陰間的那日，我為它遮蓋深淵，攔住江河，使眾水停流，以表哀悼。我使 黎巴嫩 為它悲哀，田野的樹木都因它枯萎。
EZEK|31|16|我把它扔到陰間，與下到地府的人一同墜落。那時，列國聽見墜落的響聲就震驚； 伊甸 一切的樹木，就是 黎巴嫩 中得水滋潤、最佳最美的樹，在地底下都得了安慰。
EZEK|31|17|這些樹也要與它同下陰間，到被刀所殺的人那裏；它們曾作它的膀臂 ，在列國中曾居住在它的蔭下。
EZEK|31|18|在這樣的榮耀與威勢中， 伊甸 樹木有誰能與你相比呢？然而你要與 伊甸 的樹木一同到地底下；在未受割禮的人中，與被刀所殺的人一同躺下。 「法老和他的軍隊正是如此。這是主耶和華說的。」
EZEK|32|1|第十二年十二月初一，耶和華的話臨到我，說：
EZEK|32|2|「人子啊，你要為 埃及 王法老作哀歌，說： 你在列國中，如同少壯獅子， 卻像海裏的海怪， 衝出江河， 以爪攪動諸水， 使江河渾濁。
EZEK|32|3|主耶和華如此說： 許多民族聚集時， 我要將我的網撒在你身上， 他們要把你拉上來。
EZEK|32|4|我要把你丟在地上， 拋在田野， 使空中的飛鳥落在你身上， 遍地的野獸因你得以飽足。
EZEK|32|5|我要將你的肉丟在山間， 用你巨大的屍首 填滿山谷。
EZEK|32|6|我要以你所流的血 浸透大地， 漫過山頂， 溢滿河道。
EZEK|32|7|我毀滅你時， 要遮蔽諸天， 使眾星昏暗； 我必以密雲遮掩太陽， 月亮也不放光。
EZEK|32|8|我要使天上發亮的光體 在你上面變為昏暗， 使你的地也變為黑暗。 這是主耶和華說的。
EZEK|32|9|「我使你在列國，在你所不認識的列邦中滅亡 。那時，我必使許多民族的心因你愁煩。
EZEK|32|10|當我在他們面前舉起我的刀，我要使許多民族因你驚恐，他們的君王也必因你極其恐慌。在你仆倒的日子，他們各人為自己的性命時時戰兢。
EZEK|32|11|主耶和華如此說： 巴比倫 王的刀必臨到你。
EZEK|32|12|我必藉勇士的刀使你的軍隊仆倒；這些勇士都是列國中兇暴的人。 他們必使 埃及 的驕傲歸於無有， 埃及 的軍隊必被滅絕。
EZEK|32|13|我要除滅眾水旁一切的走獸， 人的腳必不再攪渾這水， 獸的蹄也不攪渾這水。
EZEK|32|14|那時，我必使他們的水澄清， 使他們的江河像油緩流。 這是主耶和華說的。
EZEK|32|15|我使 埃及 地荒廢， 使這地空無一物， 又擊殺其中所有的居民； 那時，他們就知道我是耶和華。
EZEK|32|16|「這是一首為人所吟唱的哀歌；列國的女子要唱這哀歌，她們要為 埃及 和它的軍隊唱這哀歌。這是主耶和華說的。」
EZEK|32|17|第十二年某月 十五日，耶和華的話臨到我，說：
EZEK|32|18|「人子啊，你要為 埃及 的軍隊哀號，把他們和強盛之國 一同扔到地底下，與那些下到地府的人在一起。
EZEK|32|19|『你的美麗勝過誰呢？ 墜落吧，與未受割禮的人躺在一起！』
EZEK|32|20|他們要仆倒在被刀所殺的人當中。 埃及 被交給刀劍，人要把它和它的軍隊拉走。
EZEK|32|21|強壯的勇士要在陰間對 埃及 王和他的盟友說話；他們未受割禮，被刀劍所殺，已經墜落躺下。
EZEK|32|22|「 亞述 和它的全軍在那裏，四圍都是墳墓；他們全都是被殺倒在刀下的人。
EZEK|32|23|他們的墳墓在地府極深之處，它的眾軍環繞它的墳墓，他們全都是被殺倒在刀下的人，曾在活人之地使人驚恐。
EZEK|32|24|「 以攔 在那裏，它的全軍環繞它的墳墓；他們全都是被殺倒在刀下、未受割禮而到地底下的，曾在活人之地使人驚恐；他們與下到地府的人一同擔當羞辱。
EZEK|32|25|人為它和它的軍隊在被殺的人中設立床榻，四圍都是墳墓；他們都是未受割禮被刀所殺的，曾在活人之地使人驚恐；他們與下到地府的人一同擔當羞辱。 以攔 已列在被殺的人中。
EZEK|32|26|「 米設 、 土巴 和他們的全軍都在那裏，四圍都是墳墓；他們都是未受割禮被刀所殺的，曾在活人之地使人驚恐。
EZEK|32|27|他們不得與那未受割禮 仆倒的勇士躺在一起；這些勇士帶著兵器下到陰間，頭枕著刀劍，骨頭帶著本身的罪孽，曾在活人之地使人驚恐。
EZEK|32|28|法老啊，你必與未受割禮的人一起毀滅，與被刀所殺的人躺在一起。
EZEK|32|29|「 以東 在那裏，它的君王和所有官長雖然英勇，還是與被刀所殺的人同列；他們必與未受割禮的和下到地府的人躺在一起。
EZEK|32|30|「在那裏有北方的眾王子和所有的 西頓 人，全都與被殺的人一同下去。他們雖然英勇，使人驚恐，還是蒙羞。他們未受割禮，和被刀所殺的人躺在一起，與下到地府的人一同擔當羞辱。
EZEK|32|31|「法老看見他們，就為他的軍兵，就是被刀所殺屬法老的人和他的全軍感到安慰。這是主耶和華說的。
EZEK|32|32|我任憑法老在活人之地使人驚恐，法老和他的軍兵必躺在未受割禮和被刀所殺的人中。這是主耶和華說的。」
EZEK|33|1|耶和華的話臨到我，說：
EZEK|33|2|「人子啊，你要吩咐本國的百姓，對他們說：我使刀劍臨到哪一國，哪一國的百姓從他們中間選立一人，作為守望者。
EZEK|33|3|守望者見刀劍臨到那地，若吹角警戒百姓，
EZEK|33|4|有人聽見角聲卻不受警戒，刀劍來除滅了他，這人的血必歸到自己頭上。
EZEK|33|5|他聽見角聲，不受警戒，他的血必歸到自己身上；他若受警戒，就救了自己的命。
EZEK|33|6|倘若守望者見刀劍臨到，卻不吹角，以致百姓未受警戒，刀劍來殺了他們中間的一個人，這人雖然因自己的罪孽而死，我卻要從守望者的手裏討他的血債。
EZEK|33|7|「人子啊，我照樣立你作 以色列 家的守望者；你要聽我口中的話，替我警戒他們。
EZEK|33|8|我對惡人說：『惡人哪，你必要死！』你若不開口警戒惡人，使他離開所行的道，這惡人必因自己的罪孽而死，我卻要從你手裏討他的血債。
EZEK|33|9|但是你，你若警戒惡人，叫他離棄所行的道，他仍不轉離，他必因自己的罪孽而死，你卻救了自己的命。」
EZEK|33|10|「人子啊，你要對 以色列 家說：你們曾這樣說：『我們的過犯罪惡在自己身上，我們必因此消滅，怎能存活呢？』
EZEK|33|11|你要對他們說，主耶和華說：我指著我的永生起誓，我斷不喜悅惡人死亡，惟喜悅惡人轉離他所行的道而存活。 以色列 家啊，你們回轉，回轉離開惡道吧！何必死亡呢？
EZEK|33|12|人子啊，你要對本國的百姓說：義人的義，在他犯罪之日不能救他；至於惡人的惡，在他轉離惡行之日不會使他傾倒；義人在他犯罪之日不能因自己的義存活。
EZEK|33|13|我對義人說：『你必存活！』他若倚靠自己的義作惡，所行的義就不被記念；他必因所作的惡死亡。
EZEK|33|14|我對惡人說：『你必死亡！』他若轉離他的罪惡，行公平公義的事；
EZEK|33|15|惡人若歸還抵押品，歸回所搶奪的東西，遵行生命的律例，不再作惡；他必存活，不致死亡。
EZEK|33|16|他所犯的一切罪必不被記念；他行了公平公義的事，必要存活。
EZEK|33|17|「你本國的百姓說：『主的道不公平。』其實他們，他們的道才是不公平。
EZEK|33|18|義人轉離自己的義作惡，他必因此而死亡。
EZEK|33|19|惡人轉離他的惡，行公平公義的事，他必因此而存活。
EZEK|33|20|你們還說：『主的道不公平。』 以色列 家啊，我必按你們各人所行的審判你們。」
EZEK|33|21|我們被擄後第十二年的十月初五，有人從 耶路撒冷 逃到我這裏，說：「城已被攻破。」
EZEK|33|22|逃來的人到的前一天晚上，耶和華的手按在我身上，開我的口。第二天早晨，等那人來到我這裏，我的口就開了，不再說不出話來。
EZEK|33|23|耶和華的話臨到我，說：
EZEK|33|24|「人子啊，住在 以色列 荒廢之地的人說：『 亞伯拉罕 一人能得這地為業，我們人數眾多，這地更是給我們為業的。』
EZEK|33|25|所以你要對他們說，主耶和華如此說：你們吃帶血的食物，向偶像舉目，並且流人的血，你們還能得這地為業嗎？
EZEK|33|26|你們倚靠自己的刀劍行可憎的事，人人污辱鄰舍的妻，你們還能得這地為業嗎？
EZEK|33|27|你要對他們這樣說，主耶和華如此說：我指著我的永生起誓，在廢墟的，必倒在刀下；在田野的，必交給野獸吞吃；在堡壘和洞中的，必遭瘟疫而死。
EZEK|33|28|我必使這地荒廢荒涼，它驕傲的權勢也必止息； 以色列 的山都必荒廢，無人經過。
EZEK|33|29|我因他們所做一切可憎的事，使地荒廢荒涼；那時，他們就知道我是耶和華。」
EZEK|33|30|「你，人子啊，你本國的百姓在城牆旁邊、在房屋門口談論你。弟兄對弟兄彼此說：『來吧！聽聽有甚麼話從耶和華而出。』
EZEK|33|31|他們如同百姓前來，來到你這裏，坐在你面前彷彿是我的子民。他們聽了你的話，卻不實行；因為他們口裏說愛，心卻追隨財利。
EZEK|33|32|看哪，他們看你如同一個唱情歌的人 ，聲音優雅、善於奏樂；他們聽了你的話，卻不實行。
EZEK|33|33|看哪，這話就要應驗；應驗時，他們就知道在他們中間有了先知。」
EZEK|34|1|耶和華的話臨到我，說：
EZEK|34|2|「人子啊，你要向 以色列 的牧人說預言，對他們說，主耶和華如此說：禍哉！ 以色列 的牧人只知牧養自己。牧人豈不當牧養群羊嗎？
EZEK|34|3|你們吃肥油 、穿羊毛、宰殺肥羊，卻不牧養群羊。
EZEK|34|4|瘦弱的，你們不調養；有病的，你們不醫治；受傷的，你們未包紮；被逐的，你們不去領回；失喪的，你們不尋找；卻用暴力嚴嚴地轄制牠們 。
EZEK|34|5|牠們因無牧人就分散；既分散，就成為一切野獸的食物。
EZEK|34|6|我的羊流落眾山之間和各高岡上，分散在全地，無人去尋，無人去找。
EZEK|34|7|「所以，你們這些牧人要聽耶和華的話。
EZEK|34|8|主耶和華說：我指著我的永生起誓，我的羊因無牧人就成為掠物，也作了一切野獸的食物。我的牧人不尋找我的羊；這些牧人只知餵養自己，並不餵養我的羊。
EZEK|34|9|所以你們這些牧人要聽耶和華的話。
EZEK|34|10|主耶和華如此說：看哪，我必與牧人為敵，從他們手裏討回我的羊，使他們不再牧放群羊；牧人也不再餵養自己。我必救我的羊脫離他們的口，不再作他們的食物。」
EZEK|34|11|「主耶和華如此說：『看哪，我必親自尋找我的羊，將牠們尋見。
EZEK|34|12|牧人在羊群四散的日子怎樣尋找他的羊，我必照樣尋找我的羊。這些羊在密雲黑暗的日子散在各處，我要從那裏救回牠們。
EZEK|34|13|我要從萬民中領出牠們，從各國聚集牠們，引領牠們歸回故土。我要在 以色列 山上，在一切溪水旁邊，在境內所有可居住的地牧養牠們。
EZEK|34|14|我要在肥美的草場牧養牠們。牠們的圈必在 以色列 高處的山上，牠們必躺臥在佳美的圈內，在 以色列 山肥美的草場上吃草。
EZEK|34|15|我要親自牧養我的群羊，使牠們得以躺臥。這是主耶和華說的。
EZEK|34|16|失喪的，我必尋找；被逐的，我必領回；受傷的，我必包紮；有病的，我必醫治；只是肥的壯的，我要除滅 ；我必秉公牧養牠們。』
EZEK|34|17|「我的羊群哪，論到你們，主耶和華如此說：看哪，我要在羊與羊中間、公綿羊與公山羊中間施行審判。
EZEK|34|18|你們在肥美的草場上吃草還以為是小事嗎？竟用你們的腳踐踏剩下的草；你們喝了清水，竟用你們的腳攪渾剩下的水。
EZEK|34|19|至於我的羊，只能吃你們所踐踏的，喝你們所攪渾的。
EZEK|34|20|「所以，主耶和華對牠們如此說：看哪，我要親自在肥羊和瘦羊中間施行審判。
EZEK|34|21|因為你們用側邊用肩推擠一切瘦弱的羊，又用角牴撞，使牠們四散在外；
EZEK|34|22|所以，我要拯救我的群羊，牠們必不再作掠物；我也要在羊和羊中間施行審判。
EZEK|34|23|我必在他們之上立一牧人 ，就是我的僕人 大衛 ，牧養牠們；他必牧養他們，作他們的牧人。
EZEK|34|24|我─耶和華必作他們的上帝，我的僕人 大衛 要在他們中間作王。這是我─耶和華說的。
EZEK|34|25|「我要與他們立平安的約，使惡獸從境內斷絕；他們在曠野也能安然居住，在樹林也能躺臥。
EZEK|34|26|我要使他們和我山岡的四圍蒙福；我也必叫時雨落下，使福如甘霖降下。
EZEK|34|27|田野的樹木必結果子，地也必有出產；他們要在自己的土地安然居住。我折斷他們所負的軛，救他們脫離奴役他們之人的手；那時，他們就知道我是耶和華。
EZEK|34|28|他們必不再作外邦人的掠物，地上的野獸也不再吞吃他們；他們卻要安然居住，無人使他們驚嚇。
EZEK|34|29|我必為他們建立聞名的 栽種之地；他們在境內就不再為饑荒所滅，也不再受列國的羞辱。
EZEK|34|30|他們必知道我─耶和華他們的上帝與他們同在，並知道他們， 以色列 家，是我的子民。這是主耶和華說的。
EZEK|34|31|你們這些人，你們是我的羊，我草場上的羊；我是你們的上帝。這是主耶和華說的。」
EZEK|35|1|耶和華的話臨到我，說：
EZEK|35|2|「人子啊，你要面向 西珥山 ，向它說預言，
EZEK|35|3|對它說，主耶和華如此說： 西珥山 ，看哪，我與你為敵，必伸手攻擊你，使你荒涼荒廢。
EZEK|35|4|我必使你的城鎮變為廢墟，使你成為荒涼；你就知道我是耶和華。
EZEK|35|5|因為你永懷仇恨，在 以色列 人遭遇災難、罪孽到了盡頭時，把他們交給刀劍，
EZEK|35|6|所以主耶和華說：我指著我的永生起誓，我必使你遭遇血的報應，血必追趕你；你既不恨惡血，血必追趕你。
EZEK|35|7|我要使 西珥山 荒涼荒廢，把來往經過的人從它那裏剪除。
EZEK|35|8|我要使 西珥山 佈滿被殺的人。被刀殺的要倒在小山和山谷，並一切的溪水中。
EZEK|35|9|我必使你永遠荒涼，使你的城鎮無人居住，你們就知道我是耶和華。
EZEK|35|10|「因為你曾說『這二國、這二邦必歸我，我們必得為業』，其實耶和華仍在那裏；
EZEK|35|11|所以主耶和華說：我指著我的永生起誓，我必照你因仇恨向他們發的怒氣和嫉妒對待你；我審判你的時候，要在他們中間顯明自己。
EZEK|35|12|你必知道我─耶和華已聽見你一切凌辱的話，是針對 以色列 群山說的：『這些山荒涼了，它們是給我們作食物的。』
EZEK|35|13|你們用口向我說誇大的話，增多與我敵對的話，我都聽見了。
EZEK|35|14|主耶和華如此說：全地歡樂的時候，我必使你荒涼。
EZEK|35|15|你怎樣因 以色列 家的地業荒涼而喜樂，我也要照你所做的對待你。 西珥山 哪，你和 以東 全地都必荒涼；人就知道 我是耶和華。」
EZEK|36|1|「人子啊，你要對 以色列 群山說預言： 以色列 群山哪，要聽耶和華的話。
EZEK|36|2|主耶和華如此說，因仇敵說：『啊哈！這古老的丘壇都歸我們為業了！』
EZEK|36|3|所以你要預言，說：主耶和華如此說：因為敵人使你荒涼，四圍踐踏你，要叫你歸其餘的列國為業，使你們成為各族的話柄與百姓的笑談；
EZEK|36|4|因此， 以色列 群山哪，要聽主耶和華的話。對那遭四圍其餘列國佔據、譏刺的大山小岡、水溝山谷、荒廢之地、被棄之城，主耶和華如此說；
EZEK|36|5|所以，主耶和華如此說：我因妒火中燒，就責備其餘的列國和 以東 的眾人。他們快樂滿懷，心存恨惡，將我的地佔為己有，視為被拋棄的掠物。
EZEK|36|6|所以，你要指著 以色列 地說預言，對大山小岡、水溝山谷說，主耶和華如此說：看哪，我在妒忌和憤怒中宣佈：因你們曾受列國的羞辱，
EZEK|36|7|所以我起誓說，你們四圍的列國要擔當自己的羞辱。這是主耶和華說的。
EZEK|36|8|「 以色列 群山哪，要長出枝條，為我子民 以色列 結出果子，因為他們即將來到。
EZEK|36|9|看哪，我是幫助你們的，我要轉向你們，使你們得以耕作栽種。
EZEK|36|10|我要使 以色列 全家在你們那裏人數增多，城鎮有人居住，廢墟重新建造。
EZEK|36|11|我要使人丁和牲畜在你們那裏加增，他們必生養眾多。我要使你們那裏像以前一樣有人居住，並要賜福，比先前更多；你們就知道我是耶和華。
EZEK|36|12|我要使我的子民 以色列 在你們那裏行走，他們必得你為業；你就成為他們的產業，不再使他們喪失兒女。
EZEK|36|13|主耶和華如此說，因為人對你們說『你是吞吃人的，又使國民喪失兒女』，
EZEK|36|14|所以你必不再吞吃人，也不再使國民喪失兒女。這是主耶和華說的。
EZEK|36|15|我使你不再聽見列國的羞辱；你必不再受萬民的辱罵，也不再使國民絆跌。這是主耶和華說的。」
EZEK|36|16|耶和華的話臨到我，說：
EZEK|36|17|「人子啊， 以色列 家住本地的時候，所作所為使那地玷污。他們的行為在我面前，好像婦人在經期中那樣污穢。
EZEK|36|18|所以我因他們在那地流人的血，且以偶像使那地玷污，就把我的憤怒傾倒在他們身上。
EZEK|36|19|我將他們分散到列國，四散在列邦，按他們的所作所為懲罰他們。
EZEK|36|20|他們到了 所去的列國，使我的聖名被褻瀆；因為人談論他們說，這是耶和華的子民，卻從耶和華的地出來。
EZEK|36|21|但我顧惜我的聖名，就是 以色列 家在所到的列國中褻瀆的。
EZEK|36|22|「所以，你要對 以色列 家說，主耶和華如此說： 以色列 家啊，我做這事不是為你們，而是為了我的聖名，就是你們在所到的列國中褻瀆的。
EZEK|36|23|我要使我至大的名顯為聖；這名在列國中已遭褻瀆，是你們在他們中間褻瀆的。我在他們眼前，在你們身上顯為聖的時候，他們就知道我是耶和華。這是主耶和華說的。
EZEK|36|24|我必從列國帶領你們，從列邦聚集你們，領你們回到本地。
EZEK|36|25|我必灑清水在你們身上，你們就潔淨了。我要潔淨你們，使你們脫離一切的污穢，棄絕一切的偶像。
EZEK|36|26|我也要賜給你們一顆新心，將新靈放在你們裏面，又從你們的肉體中除掉石心，賜給你們肉心。
EZEK|36|27|我必將我的靈放在你們裏面，使你們順從我的律例，謹守遵行我的典章。
EZEK|36|28|你們必住在我所賜給你們祖先之地；你們要作我的子民，我要作你們的上帝。
EZEK|36|29|我要救你們脫離一切的污穢，也要令五穀豐登，使你們不再遭遇饑荒。
EZEK|36|30|我要使樹木多結果子，田地多出土產，好叫你們不再因饑荒被列國凌辱。
EZEK|36|31|那時，你們必追念自己的惡行和不好的作為，就因你們的罪孽和可憎的事厭惡自己。
EZEK|36|32|你們要知道，我這樣做不是為你們。 以色列 家啊，你們當為自己的行為抱愧蒙羞。這是主耶和華說的。
EZEK|36|33|「主耶和華如此說：我潔淨你們，使你們脫離一切罪孽的日子，必使城鎮有人居住，廢墟重新建造。
EZEK|36|34|這荒蕪的土地，曾被過路的人看為荒蕪，現今卻得以耕種。
EZEK|36|35|他們必說：『這荒蕪之地，現在成了像 伊甸園 一樣；這荒涼、荒廢、毀壞的城鎮，現今堅固，有人居住。』
EZEK|36|36|那時，在你們四圍其餘的列國必知道，我─耶和華修造那毀壞之處，開墾那荒蕪之地。我─耶和華說了這話，就必成就。
EZEK|36|37|「主耶和華如此說：我要回應 以色列 家的求問，成全他們，增添他們的人數，使他們多如羊群。
EZEK|36|38|在 耶路撒冷 守節時，作為祭物所獻的羊群有多少，照樣，荒涼的城鎮必為人群所充滿；他們就知道我是耶和華。」
EZEK|37|1|耶和華的手按在我身上。耶和華藉著他的靈帶我出去，把我放在平原中，平原遍滿骸骨。
EZEK|37|2|他使我從骸骨的四圍經過，看哪，平原上面的骸骨甚多，看哪，極其枯乾。
EZEK|37|3|他對我說：「人子啊，這些骸骨能活過來嗎？」我說：「主耶和華啊，你是知道的。」
EZEK|37|4|他又對我說：「你要向這些骸骨說預言，對它們說：枯乾的骸骨啊，要聽耶和華的話。
EZEK|37|5|主耶和華對這些骸骨如此說：『看哪，我必使氣息 進入你們裏面，你們就要活過來。
EZEK|37|6|我要給你們加上筋，長出肉，又給你們包上皮，使氣息進入你們裏面，你們就要活過來；你們就知道我是耶和華。』」
EZEK|37|7|於是，我遵命說預言。正說預言的時候，有響聲，看哪，有地震；骨與骨彼此接連。
EZEK|37|8|我觀看，看哪，骸骨上面有筋，長了肉，又包上皮，只是裏面還沒有氣息。
EZEK|37|9|耶和華對我說：「人子啊，你要說預言，向風 說預言。你要說，耶和華如此說：氣息啊，要從四方 而來，吹在這些被殺的人身上，使他們活過來。」
EZEK|37|10|於是我遵命說預言，氣息就進入骸骨，骸骨就活過來，並且用腳站起來，成為極大的軍隊。
EZEK|37|11|他對我說：「人子啊，這些骸骨就是 以色列 全家。他們說：『看哪，我們的骨頭枯乾了，我們的指望失去了，我們滅絕淨盡了！』
EZEK|37|12|所以你要說預言，對他們說，主耶和華如此說：我的子民，看哪，我要打開你們的墳墓，把你們帶出墳墓，領你們進入 以色列 地。
EZEK|37|13|我的子民哪，我打開你們的墳墓，把你們帶出墳墓時，你們就知道我是耶和華。
EZEK|37|14|我必將我的靈放在你們裏面，你們就要活過來。我把你們安置在本地，你們就知道我─耶和華說了這話，就必成就。這是耶和華說的。」
EZEK|37|15|耶和華的話臨到我，說：
EZEK|37|16|「人子啊，你要取一根木杖，在其上寫『為 猶大 和他的盟友 以色列 人』；又取一根 木杖，在其上寫『為 約瑟 ，就是 以法蓮 的杖，和他的盟友 以色列 全家』。
EZEK|37|17|你要將這兩根木杖彼此相接，連成一根，使它們在你手中合而為一。
EZEK|37|18|當你本國的子民對你說：『你這是甚麼意思，你不指示我們嗎？』
EZEK|37|19|你就對他們說，主耶和華如此說：看哪，我要將 約瑟 和他的盟友 以色列 支派的杖，就是在 以法蓮 手中的那根，與 猶大 的杖接連成為一根，在我手中合而為一。
EZEK|37|20|你要在他們眼前，把寫了字的那兩根杖拿在手中，
EZEK|37|21|對他們說，主耶和華如此說：看哪，我要從 以色列 人所到的列國帶領他們，從四圍聚集他們，領他們回到本地。
EZEK|37|22|我要使他們在這地，在 以色列 群山上成為一國，必有一王作他們全體的王。他們不再成為二國，絕不再分為二國。
EZEK|37|23|他們不再因偶像和可憎的物，並一切的罪過玷污自己。我卻要救他們離開一切犯罪所住的地方 ；我要潔淨他們，如此，他們要作我的子民，我要作他們的上帝。』
EZEK|37|24|「我的僕人 大衛 要作他們的王；他們全體必歸一個牧人。他們必順從我的典章，謹守遵行我的律例。
EZEK|37|25|他們要住在我賜給我僕人 雅各 的地上，就是你們列祖所住之地。他們和他們的子孫，並子孫的子孫，都永遠住在那裏。我的僕人 大衛 要作他們的王，直到永遠；
EZEK|37|26|並且我要與他們立平安的約，作為永約。我要安頓他們，使他們人數增多，又在他們中間設立我的聖所，直到永遠。
EZEK|37|27|我的居所必在他們中間；我要作他們的上帝，他們要作我的子民。
EZEK|37|28|我的聖所在 以色列 人中間直到永遠，列國就知道是我─耶和華使 以色列 分別為聖。」
EZEK|38|1|耶和華的話臨到我，說：
EZEK|38|2|「人子啊，你要面向 瑪各 地的 歌革 ，就是 米設 和 土巴 的大王，向他說預言。
EZEK|38|3|你要說，主耶和華如此說： 米設 和 土巴 的大王 歌革 ，看哪，我與你為敵。
EZEK|38|4|我要把你掉轉過來，用鉤子鉤住你的腮頰，把你和你的軍兵、馬匹、騎兵都帶走。他們全都披掛整齊，成為大軍，佩帶大小盾牌，各人拿著刀劍；
EZEK|38|5|他們當中有 波斯 人、 古實 人和 弗 人，都帶著盾牌和頭盔；
EZEK|38|6|還有 歌篾 人和他的軍隊，北方極遠的 陀迦瑪 族和他的軍隊，這許多民族都跟著你。
EZEK|38|7|「你和聚集到你那裏的軍隊都要預備，預備妥當，你要作他們的守衛。
EZEK|38|8|過了多日，你必被差派；到末後之年，你要來到那脫離刀劍、從列國召集回來的人所住之地，來到 以色列 常久荒涼的山上；他們都從列國中被領出，在那裏安然居住。
EZEK|38|9|你和你的全軍，並跟隨你的許多民族都要上來，如暴風刮來，如密雲遮蓋地面。
EZEK|38|10|「主耶和華如此說：那時，你的心必起意念，圖謀惡計，
EZEK|38|11|說：『我要上那無牆的鄉村之地，到那安靜的居民那裏，他們無牆，無門、無閂，安然居住。
EZEK|38|12|我去那裏要搶財為擄物，奪貨為掠物，反手攻擊那從前荒涼、現在有人居住之地，又攻擊那從列國招聚出來、得了牲畜財貨、住在地的高處的百姓。』
EZEK|38|13|示巴 人、 底但 人、 他施 的商人和他們的少壯獅子都對你說：『你來是要搶財為擄物嗎？你聚集軍隊是要奪貨為掠物，奪取金銀，擄去牲畜、財貨，搶奪許多財寶為擄物嗎？』
EZEK|38|14|「人子啊，你要因此說預言，對 歌革 說，主耶和華如此說：我的子民 以色列 安然居住時，你是知道的。
EZEK|38|15|你從你的地方，從北方極遠處率領許多民族前來，他們都騎著馬，是一隊強而多的軍兵。
EZEK|38|16|歌革 啊，你必上來攻擊我的子民 以色列 ，如密雲遮蓋地面。末後的日子，我必領你來攻擊我的地，我藉你在列國眼前顯為聖的時候，他們就要認識我。
EZEK|38|17|主耶和華如此說：我在古時藉我僕人 以色列 眾先知所說的，不就是你嗎？ 他們在那些日子，多年說預言，我必領你來攻擊 以色列 人。」
EZEK|38|18|「主耶和華說： 歌革 上來攻擊 以色列 地的時候，我的怒氣要從鼻孔裏發出。
EZEK|38|19|我在妒忌和如火的烈怒中說：那日在 以色列 地必有大震動，
EZEK|38|20|甚至海中的魚、天空的鳥、野地的獸，和地上爬的各種爬行動物，並地面上的眾人，因見我的面就都震動；山嶺崩裂，陡巖塌陷，一切的牆都必坍塌。
EZEK|38|21|我必令刀劍在我的眾山攻擊 歌革 ；人要用刀劍殺害弟兄。這是主耶和華說的。
EZEK|38|22|我要用瘟疫和血懲罰他。我也必降暴雨、大冰雹、火及硫磺在他和他的軍隊，並跟隨他的許多民族身上。
EZEK|38|23|我必顯為大，顯為聖，在許多國家眼前顯明自己；他們就知道我是耶和華。」
EZEK|39|1|「你，人子啊，要向 歌革 說預言。你要說，主耶和華如此說： 米設 和 土巴 的大王 歌革 ，看哪，我與你為敵。
EZEK|39|2|我要把你調轉過來，帶領你，從北方極遠的地方上來，帶你到 以色列 的群山上。
EZEK|39|3|我要打落你左手的弓，打掉你右手的箭。
EZEK|39|4|你和你的全軍，並跟隨你的列國的人，都必倒在 以色列 的群山上。我要將你給各類攫食的飛鳥和野地的走獸作食物。
EZEK|39|5|你必倒在田野，因為我曾說過，這是主耶和華說的。
EZEK|39|6|我要降火在 瑪各 和海島安然居住的人身上，他們就知道我是耶和華。
EZEK|39|7|「我要在我的子民 以色列 中彰顯我的聖名，不容我的聖名再被褻瀆，列國就知道我─耶和華是 以色列 中的聖者。
EZEK|39|8|看哪，時候到了，必然成就，這就是我曾說過的日子。這是主耶和華說的。
EZEK|39|9|「住 以色列 城鎮的人要出去生火，用軍器燃燒，就是大小盾牌、弓箭、棍棒、槍矛；用它們來燒火，直燒了七年。
EZEK|39|10|他們不必從田野撿柴，也不必從森林伐木，因為他們要用這些軍器燒火。他們要搶奪那搶奪他們的人，擄掠那擄掠他們的人。這是主耶和華說的。」
EZEK|39|11|「當那日，我要把 以色列 境內、海東邊的 旅人谷 給 歌革 在那裏作墳地 ，阻擋了旅行的人 。在那裏，人要埋葬 歌革 和他的軍兵，稱那地為 哈們‧歌革谷 。
EZEK|39|12|以色列 家的人要用七個月埋葬他們，好使那地潔淨。
EZEK|39|13|那地所有的百姓都來埋葬他們。當我得榮耀的日子，這事必叫百姓得名聲。這是主耶和華說的。
EZEK|39|14|他們要分派人專職巡查遍地，埋葬那遺留在地面上入侵者的屍首，好潔淨全地。過了七個月，他們還要再巡查。
EZEK|39|15|巡查的人要遍行全地，見有人的骸骨，就在旁邊立一標記，等埋葬的人來將骸骨葬在 哈們‧歌革谷 ，
EZEK|39|16|且有一城要取名為 哈摩那 。他們必這樣潔淨那地。
EZEK|39|17|「你，人子啊，主耶和華如此說：你要向各類的飛鳥和野地的走獸說：你們要聚集，來吧，從四方聚集來吃我為你們準備的祭物，就是在 以色列 的群山上豐盛的祭物，叫你們吃肉、喝血。
EZEK|39|18|你們要吃勇士的肉，喝地上領袖的血，如吃公綿羊、羔羊、公山羊、公牛；他們全都是 巴珊 的肥畜。
EZEK|39|19|你們吃我為你們準備的祭物，必吃油脂直到飽了，喝血直到醉了。
EZEK|39|20|你們要因我席上的馬匹、騎兵、勇士和所有的戰士而飽足。這是主耶和華說的。」
EZEK|39|21|「我要在列國中彰顯我的榮耀，萬國就必看見我怎樣把手加在他們身上，施行審判。
EZEK|39|22|從那日以後， 以色列 家就知道我是耶和華─他們的上帝，
EZEK|39|23|列國也必知道， 以色列 家被擄掠是因他們的罪孽。他們得罪我，我就轉臉不顧他們，將他們交在敵人手中，使他們全都倒在刀下。
EZEK|39|24|我照他們的污穢和罪過待他們，轉臉不顧他們。
EZEK|39|25|「所以主耶和華如此說：現在，我要使 雅各 被擄的人歸回，要憐憫 以色列 全家，又為我的聖名發熱心。
EZEK|39|26|我將他們從萬民中領回，從仇敵之地召來，在許多國家的眼前，在他們身上顯為聖，他們在本地安然居住，無人使他們驚嚇，那時，他們要擔當 自己的羞辱和干犯我的一切罪。
EZEK|39|27|
EZEK|39|28|我使他們被擄到列國，後又聚集他們回到本地，不再留一人在那裏，那時他們就知道我是耶和華─他們的上帝。
EZEK|39|29|我不再轉臉不顧他們，因我已將我的靈澆灌 以色列 家。這是主耶和華說的。」
EZEK|40|1|我們被擄的第二十五年， 耶路撒冷城 攻破後十四年，正在年初，某月初十，就在那一天，耶和華的手按在我身上，把我帶到那裏。
EZEK|40|2|在上帝的異象中，他帶我到 以色列 地，把我安置在一座極高的山上；在山的南邊有彷彿一座城的建築物。
EZEK|40|3|他帶我到那裏，看哪，有一人面貌 如銅，手拿麻繩和丈量的蘆葦竿，站在門口。
EZEK|40|4|那人對我說：「人子啊，凡我所指示你的，你都要用眼看，用耳聽，並要放在心上。我帶你到這裏來，為要指示你；凡你所見的，都要告訴 以色列 家。」
EZEK|40|5|看哪，殿外四圍有牆。那人手拿丈量的蘆葦竿，長六肘，每肘再加一掌。他量圍牆，寬一竿，高一竿。
EZEK|40|6|他到了朝東的門，就上臺階，量這門的門檻，寬一竿；這門檻寬一竿。
EZEK|40|7|又有守衛房，每間長一竿，寬一竿，守衛房之間相隔五肘。挨著通往殿之門走廊的門檻，一竿。
EZEK|40|8|他量通往殿之門的走廊，一竿。
EZEK|40|9|他量門的走廊，八肘；牆柱，二肘；門的走廊通往殿那裏。
EZEK|40|10|往東的門有守衛房：這旁三間，那旁三間，大小都一樣；這邊和那邊的牆柱，大小也一樣。
EZEK|40|11|他量門的入口，寬十肘，門長十三肘。
EZEK|40|12|守衛房前有矮牆，一肘，那邊的矮牆也是一肘；守衛房這邊六肘，那邊也是六肘。
EZEK|40|13|他量門，從守衛房這邊的房頂到那邊的房頂，寬二十五肘；入口與入口相對。
EZEK|40|14|他量牆柱，六十肘，院子的四周圍有挨著牆柱的門。
EZEK|40|15|從大門入口到裏面門的走廊，五十肘。
EZEK|40|16|守衛房和四圍挨著牆柱的門，都有嵌壁式的窗戶，廊子也有；裏面到處都有窗戶，牆柱上雕刻著棕樹。
EZEK|40|17|他帶我到外院，看哪，院子的四圍有房間，有石板地；石板地上有三十個房間。
EZEK|40|18|沿著門側邊的石板地，就是下面的石板地，與門的長度相同。
EZEK|40|19|他量寬度，從下門的前面到內院外的前面，東向北向一百肘。
EZEK|40|20|他量外院朝北的門的長和寬。
EZEK|40|21|門的守衛房，這旁三間，那旁三間；牆柱和廊子，與第一個門的大小一樣。長五十肘，寬二十五肘。
EZEK|40|22|其窗戶和廊子，並雕刻的棕樹，與朝東的門大小一樣。要登七個臺階才能上到這門，前面 有廊子。
EZEK|40|23|內院有門與這門相對，北面東面都是如此。他從這門量到那門，共一百肘。
EZEK|40|24|他帶我往南去，看哪，朝南有門，他量門的牆柱 和廊子，大小與先前一樣。
EZEK|40|25|門兩旁與廊子的周圍都有窗戶，和先前量的窗戶一樣。門長五十肘，寬二十五肘。
EZEK|40|26|要登七個臺階才能上到這門，前面 有廊子；牆柱上雕刻著棕樹，這邊一棵，那邊一棵。
EZEK|40|27|內院朝南也有門，從這門量到朝南的那門，共一百肘。
EZEK|40|28|他帶我從南門到內院，他量南門，大小與先前一樣。
EZEK|40|29|守衛房和牆柱、廊子，大小與先前一樣。門兩旁與廊子的周圍都有窗戶。門長五十肘，寬二十五肘。
EZEK|40|30|周圍有廊子，長二十五肘，寬五肘。
EZEK|40|31|廊子朝著外院，牆柱上雕刻著棕樹。要登八個臺階才能上到這門。
EZEK|40|32|他帶我到內院的東邊，他量那門，大小與先前一樣。
EZEK|40|33|守衛房和牆柱、廊子，大小與先前一樣。門兩旁與廊子的周圍都有窗戶。長五十肘，寬二十五肘。
EZEK|40|34|廊子朝著外院。牆柱兩邊都雕刻著棕樹。要登八個臺階才能上到這門。
EZEK|40|35|他帶我到北門，他量了，大小與先前一樣，
EZEK|40|36|就是量守衛房和牆柱、廊子。門的周圍都有窗戶；門長五十肘，寬二十五肘。
EZEK|40|37|牆柱 朝著外院。牆柱兩邊都雕刻著棕樹。要登八個臺階才能上到這門。
EZEK|40|38|有房間和它的入口在門的牆柱 旁，那裏是洗燔祭牲的地方。
EZEK|40|39|在門的走廊內，這邊有兩張桌子，那邊也有兩張桌子，其上可宰殺燔祭牲、贖罪祭牲和贖愆祭牲。
EZEK|40|40|上到北門的入口，朝向外面的這邊有兩張桌子，門的走廊那邊也有兩張桌子。
EZEK|40|41|門這邊有四張桌子，那邊也有四張桌子，共八張，在其上宰殺祭牲。
EZEK|40|42|為燔祭牲的四張桌子是用石頭鑿成的，長一肘半，寬一肘半，高一肘。宰殺燔祭牲和其他祭牲所用的器皿可放在其上。
EZEK|40|43|有鉤子，寬一掌，掛在廊內的四周圍。桌子上可放祭牲的肉。
EZEK|40|44|從外面進到內門，內院裏有房間，為歌唱的人而設 ；一間在北門旁，朝南，又有一間在南 門旁，朝北。
EZEK|40|45|他對我說：「這朝南的房間是為了聖殿供職的祭司，
EZEK|40|46|那朝北的房間是為了祭壇前供職的祭司；這些祭司是 利未 人中 撒督 的子孫，近前來事奉耶和華的。」
EZEK|40|47|他又量內院，長一百肘，寬一百肘，是正方的。祭壇就在殿前。
EZEK|40|48|於是他帶我到殿前的走廊，量走廊的牆柱。這面寬五肘，那面寬五肘。 門的兩旁，這邊三肘，那邊三肘。
EZEK|40|49|走廊長二十肘，寬十一肘 。要登臺階 才能上到走廊。靠近牆柱又有柱子，這邊一根，那邊一根。
EZEK|41|1|他帶我到殿那裏，他量牆柱：這面寬六肘，那面寬六肘，寬窄與會幕相同 。
EZEK|41|2|門口寬十肘。門的兩旁，這邊五肘，那邊五肘。他又量了殿，長四十肘，寬二十肘。
EZEK|41|3|他到內殿量門的牆柱，二肘，門口六肘，門的兩旁各寬七肘。
EZEK|41|4|他量內殿，長二十肘，寬二十肘。他對我說：「這是至聖所。」
EZEK|41|5|他又量殿的牆，六肘；圍著殿有廂房，各寬四肘。
EZEK|41|6|廂房有三層，層疊而上，每層排列三十間。殿的牆四周有凸出的牆支撐廂房，廂房就不必以殿的牆為支柱。
EZEK|41|7|這圍繞著殿的廂房越高越寬；廂房圍著殿懸疊而上，所以越上面越寬，從下一層，到中一層，到上一層。
EZEK|41|8|我又見有高臺圍繞著殿，作為廂房的根基，高足足有一竿，就是六大肘。
EZEK|41|9|廂房的外牆寬五肘。殿的廂房和那邊的房間中間還有空地，寬二十肘，圍繞著殿。
EZEK|41|10|
EZEK|41|11|廂房的門口向著空地：一門向北，一門向南。周圍的空地寬五肘。
EZEK|41|12|在西邊空地之後有房子，寬七十肘，長九十肘，牆四圍厚五肘。
EZEK|41|13|這樣，他量了殿，長一百肘，又量空地和那房子並牆，共長一百肘。
EZEK|41|14|殿的前面和東邊的空地，寬一百肘。
EZEK|41|15|他量了空地後面的那房子，並兩旁的樓廊，共長一百肘。 內殿、院的走廊、
EZEK|41|16|門檻 、嵌壁式的窗戶，並對著門檻的三層樓廊，周圍都鑲上木板；地板到窗戶，窗戶都關著，
EZEK|41|17|直到門以上，就是到內殿和外殿內外四圍牆壁，都這樣測量。
EZEK|41|18|牆上雕刻基路伯和棕樹，基路伯和基路伯之間有一棵棕樹，每基路伯有兩張臉；
EZEK|41|19|人的臉向著這邊的棕樹，獅子的臉向著那邊的棕樹，殿內四周圍都是如此。
EZEK|41|20|從地板到門的上面，都有基路伯和棕樹。殿的牆就是這樣。
EZEK|41|21|殿的門柱是方的。至聖所的前面有個東西形狀像
EZEK|41|22|木頭做的壇，高三肘，長二肘 。壇角和底座 ，並四面，都是木頭做的。他對我說：「這是耶和華面前的供桌。」
EZEK|41|23|殿和聖所各有一個雙層門。
EZEK|41|24|每個門有兩扇，每扇又有兩個摺疊頁；這一扇有兩頁，另一扇也有兩頁。
EZEK|41|25|殿的門扇上雕刻著基路伯和棕樹，與刻在牆上的一樣。在外面門的走廊前有木頭做的飛簷。
EZEK|41|26|門的走廊這邊和那邊都有嵌壁式的窗戶和棕樹；殿的廂房和飛簷也是這樣。
EZEK|42|1|他帶我出來往北，到外院，又帶我進入一個房間，一面對著空地，一面對著北邊的房子。
EZEK|42|2|前面長一百肘，寬五十肘，有門向北；
EZEK|42|3|對著內院那二十肘 ，又對著外院的石板地，在第三層樓有樓廊對著樓廊。
EZEK|42|4|那些房間前有一條走道，寬十肘，往裏面有寬一肘的通道 。房門都向北。
EZEK|42|5|房間因為樓廊佔掉一些地方，所以房子的上層比中下兩層窄。
EZEK|42|6|房間分三層，卻不像外院的屋子用柱子支撐，而是從地面往上，所以一層比一層更窄。
EZEK|42|7|外面有一道牆，長五十肘，在房間前面，與朝外院的房間平行。
EZEK|42|8|靠著外院的房間長五十肘，看哪，朝聖殿的長一百肘。
EZEK|42|9|這些房間下面的東邊有一個入口，從外院可由此進入；
EZEK|42|10|其寬如院牆。朝東 也有房間，一面對著空地，一面對著房子。
EZEK|42|11|這些房間前的通道與北邊房間的通道一樣；長、寬、出口、樣式和入口都相同。
EZEK|42|12|在東邊通道的開端，正對著那道牆有門可以進入，與向南邊房間的門一樣。
EZEK|42|13|他對我說：「面對空地南邊的房間和北邊的房間，都是聖的房間；親近耶和華的祭司當在那裏吃至聖的東西，也當在那裏存放至聖的東西，就是素祭、贖罪祭和贖愆祭，因此處為聖。
EZEK|42|14|祭司進聖所，出來的時候，不可直接到外院，要在那裏放下他們供職的衣服，因為這是聖衣；要穿上別的衣服才可以到百姓所在之處。」
EZEK|42|15|他量完了內殿的大小，就帶我出朝東的門，去量院的四周圍。
EZEK|42|16|他用丈量的蘆葦竿量東面，五百竿 ；又轉去
EZEK|42|17|用丈量的蘆葦竿量北面，五百竿；又轉去
EZEK|42|18|用丈量的蘆葦竿量南面，五百竿。
EZEK|42|19|他又轉到西面，用丈量的蘆葦竿去量，五百竿。
EZEK|42|20|他量四面，長五百，寬五百，四周圍有牆，為要分別聖與俗。
EZEK|43|1|以後，他帶我到一座門，就是朝東的門。
EZEK|43|2|看哪， 以色列 上帝的榮光從東而來，他的聲音如同眾水的響聲，地因他的榮耀發光。
EZEK|43|3|我所見的異象如同從前我 來滅城的時候所見的異象，又如我在 迦巴魯河 邊所見的異象，我就臉伏於地。
EZEK|43|4|耶和華的榮光從朝東的門照入殿中。
EZEK|43|5|靈將我舉起，帶入內院，看哪，耶和華的榮光充滿了殿。
EZEK|43|6|我聽見有一位從殿中向我說話，有一人站在我旁邊。
EZEK|43|7|他對我說：「人子啊，這是我寶座之地，是我腳掌所踏之地。我要住在這裏，住在 以色列 人中間直到永遠。 以色列 家和他們的君王不可再以淫行，或在高處以君王的屍首 玷污我的聖名。
EZEK|43|8|因他們使自己的門檻挨近我的門檻，使自己的門框挨近我的門框，又使他們與我之間僅隔一牆，並且行可憎的事，玷污我的聖名，所以我發怒滅絕他們。
EZEK|43|9|現在，他們當從我面前遠離淫行和君王的屍首，我就要住在他們中間，直到永遠。
EZEK|43|10|「你，人子啊，要將這殿指示 以色列 家，讓他們量殿的大小 ，使他們因自己的罪孽羞愧。
EZEK|43|11|他們若因自己所做的一切感到羞愧，你就要將殿的規模、樣式、出口、入口，以及有關整體規模的條例、禮儀、律法指示他們 ，在他們眼前寫下，使他們遵照殿整體的規模和條例去做。
EZEK|43|12|這是殿的律法：山頂上四周圍的全地界都稱為至聖；看哪，這就是殿的律法 。」
EZEK|43|13|這些是祭壇的大小，以肘來量，這肘是一肘一掌。底座高一肘，邊寬一肘，四周圍有邊，高一虎口；這是祭壇的座 。
EZEK|43|14|從底座到下層的臺座，二肘，邊寬一肘。從小臺座到大臺座，四肘，邊寬一肘。
EZEK|43|15|壇上的爐臺，高四肘，從爐臺向上突起四個角。
EZEK|43|16|這爐臺長十二肘，寬十二肘，四面見方。
EZEK|43|17|臺座長十四肘，寬十四肘，四面見方。四周圍有邊，高半肘，底座四圍的邊寬一肘。有臺階朝東。
EZEK|43|18|他對我說：「人子啊，主耶和華如此說：這些是建造祭壇，為要在其上獻燔祭，把血灑在上面的條例：
EZEK|43|19|你要將一頭公牛犢作為贖罪祭，交給那近前來事奉我的 利未 家的祭司 撒督 的後裔；這是主耶和華說的。
EZEK|43|20|你要取那公牛犢的一些血，抹在壇的四角和臺座的四角，並周圍的邊上。你要這樣潔淨壇，為壇贖罪。
EZEK|43|21|你又要將那作贖罪祭的公牛燒在聖所外面，殿的預定之處。
EZEK|43|22|次日，要將無殘疾的公山羊獻為贖罪祭；要潔淨壇，像用公牛潔淨一樣。
EZEK|43|23|你潔淨了壇，就要將一頭無殘疾的公牛犢和羊群中一隻無殘疾的公綿羊
EZEK|43|24|奉到耶和華面前。祭司要撒鹽在其上，獻給耶和華為燔祭。
EZEK|43|25|七日內，你要每日獻一隻公山羊為贖罪祭，也要獻一頭公牛犢和羊群中的一隻公綿羊，都要沒有殘疾的。
EZEK|43|26|七日內祭司要為壇贖罪，使它潔淨，把它分別為聖。
EZEK|43|27|滿了七日，自八日以後，祭司要在壇上獻你們的燔祭和平安祭；我必悅納你們。這是主耶和華說的。」
EZEK|44|1|他又帶我回到聖所朝東的外門，那門關閉了。
EZEK|44|2|耶和華對我說：「這門必須關閉，不可敞開，誰也不可由其中進入；因為耶和華─ 以色列 的上帝已經由其中進入，所以必須關閉。
EZEK|44|3|至於君王，他必按君王的位分坐在其內，在耶和華面前吃餅。他必由這門的走廊而入，也必由此而出。」
EZEK|44|4|他又帶我由北門來到殿前。我觀看，看哪，耶和華的榮光充滿耶和華的殿，我就臉伏於地。
EZEK|44|5|耶和華對我說：「人子啊，我對你所說耶和華殿中一切的條例和律法，你要留心，用眼看，用耳聽，要留心殿的入口和聖所一切的出口。
EZEK|44|6|你要對那悖逆的 以色列 家說，主耶和華如此說： 以色列 家啊，你們行這一切可憎的事，夠了吧！
EZEK|44|7|你們把我的食物，就是脂肪和血獻上的時候，竟把心和肉體未受割禮的外邦人領進我的聖所，玷污我的殿；你們行這一切可憎的事，違背了我的約。
EZEK|44|8|你們未盡看守我聖物的職責，竟派別人在我的聖所替你們盡看守之責。
EZEK|44|9|「主耶和華如此說：所有心和肉體未受割禮的外邦人，就是住在 以色列 中間的任何外邦人，都不可進入我的聖所。」
EZEK|44|10|「 以色列 人走迷的時候， 利未 人遠離我，隨從他們的偶像走迷離開我，他們必擔當自己的罪孽。
EZEK|44|11|他們必在我的聖所當僕役，照管殿門，在殿裏伺候；他們要為百姓宰殺燔祭牲和其他祭牲，站在百姓面前伺候他們。
EZEK|44|12|因為這些 利未 人曾在偶像前伺候他們，成了 以色列 家罪孽的絆腳石，所以我向他們起誓：他們必擔當自己的罪孽。這是主耶和華說的。
EZEK|44|13|他們不可親近我，作事奉我的祭司，也不可挨近我任何一件聖物，就是至聖的物；他們卻要擔當自己的羞辱和所行可憎之事的報應。
EZEK|44|14|我要指派他們在殿裏看守，辦理殿中一切事務，做一切當做的工。」
EZEK|44|15|「 以色列 人走迷離開我的時候， 利未 家的祭司 撒督 的子孫仍然盡看守我聖所的職責；因此他們必親近我，事奉我，並且侍立在我面前，把脂肪與血獻給我。這是主耶和華說的。
EZEK|44|16|只有他們可以進我的聖所，來到我的桌前事奉我，守我吩咐的職責。
EZEK|44|17|他們進內院的門要穿細麻衣，在內院門和殿內供職時不可穿羊毛衣服。
EZEK|44|18|他們要頭戴細麻布的頭巾，腰穿細麻布的褲子；不可穿容易出汗的衣服。
EZEK|44|19|他們出到外院，到外院 百姓那裏，要脫下供職所穿的衣服，放在聖的房間內，換上別的衣服，免得因他們的衣服使百姓成為聖。
EZEK|44|20|他們不可剃頭，也不可留長髮，頭髮一定要修剪。
EZEK|44|21|祭司進內院時不可喝酒。
EZEK|44|22|他們不可娶寡婦或被休的婦人為妻，只可娶 以色列 後裔中的處女，或祭司的寡婦。
EZEK|44|23|他們要教導我的子民分辨聖與俗，使他們知道潔淨和不潔淨的分別。
EZEK|44|24|有爭訟的事，他們應當審判，按我的典章審判。他們要在我的節期守我的律法和條例，也當以我的安息日為聖日。
EZEK|44|25|祭司不可挨近死屍使自己不潔淨，只可為父親、母親、兒子、女兒、兄弟和未出嫁的姊妹使自己不潔淨。
EZEK|44|26|他潔淨之後，他們必須再為他計算七天。
EZEK|44|27|當他進內院，入聖所，在聖所中事奉的日子，要為自己獻上贖罪祭。這是主耶和華說的。
EZEK|44|28|「祭司必有產業，我就是他們的產業。不可在 以色列 中給他們基業，我就是他們的基業。
EZEK|44|29|素祭、贖罪祭和贖愆祭他們都可以吃， 以色列 中一切永獻的祭物都歸他們。
EZEK|44|30|各樣上好的初熟之物和所獻的供物，都要歸祭司。你們也要將最先的麵團給祭司；這樣，福氣就必臨到你們的家。
EZEK|44|31|無論是鳥是獸，凡自然死去的，或是被撕裂的，祭司都不可吃。」
EZEK|45|1|你們抽籤分地為業，要獻上一份作為獻給耶和華的聖地，長二萬五千肘 ，寬二萬 肘。整個地區都作為聖地。
EZEK|45|2|再從其中劃出一塊作為聖所，長五百肘，寬五百肘，四面見方；四圍再加五十肘的空地。
EZEK|45|3|從這整個範圍要劃出長二萬五千肘，寬一萬肘的地，其中要有聖所，是至聖的。
EZEK|45|4|這是地上的一塊聖地，要歸給在聖所供職、親近事奉耶和華的祭司，作為他們房屋用地與聖所的聖地。
EZEK|45|5|其餘長二萬五千肘，寬一萬肘，要歸給在殿中供職的 利未 人，作為他們二十間房屋 的地業。
EZEK|45|6|在那塊獻上的聖地旁邊，你們要劃分造城的地業，寬五千肘，長二萬五千肘，歸 以色列 全家。
EZEK|45|7|劃歸君王的地要在獻上的聖地和城用地的兩旁，面對著聖地，又面對城的用地，西至西邊的疆界，東至東邊的疆界，從西到東，長度與每支派所分得的一樣。
EZEK|45|8|這地要在 以色列 中歸君王為業。我所立的君王必不再欺壓我的子民，卻要按支派把地分給 以色列 家。
EZEK|45|9|主耶和華如此說：「 以色列 的王啊，你們夠了吧！要除掉殘暴和搶奪的事，行公平和公義，不可再勒索我的百姓。這是主耶和華說的。
EZEK|45|10|「你們要用公道的天平、公道的伊法、公道的罷特。
EZEK|45|11|伊法要與罷特等量；一罷特為賀梅珥的十分之一，一伊法也是賀梅珥的十分之一，都以賀梅珥為計算單位。
EZEK|45|12|一舍客勒是二十季拉；二十舍客勒，二十五舍客勒，十五舍客勒，合起來為你們的一彌那。
EZEK|45|13|「你們當獻的供物是這樣：一賀梅珥麥子要獻六分之一伊法，一賀梅珥大麥也要獻六分之一伊法。
EZEK|45|14|獻油的條例是這樣，按油的罷特：每一歌珥油，即十罷特或一賀梅珥，要獻十分之一罷特，原來十罷特等於一賀梅珥。
EZEK|45|15|從 以色列 水源豐沛的草場上，每二百隻羊中要獻一隻羔羊。這都可作素祭、燔祭、平安祭，來為民贖罪。這是主耶和華說的。
EZEK|45|16|這地所有的百姓都要帶這些供物到 以色列 王那裏。
EZEK|45|17|王的本分是在節期、初一、安息日，就是 以色列 家一切的盛會，奉上燔祭、素祭、澆酒祭。他要獻上贖罪祭、素祭、燔祭和平安祭，為 以色列 家贖罪。」
EZEK|45|18|主耶和華如此說：「正月初一，你要取無殘疾的公牛犢，潔淨聖所。
EZEK|45|19|祭司要取一些贖罪祭牲的血，抹在殿的門柱上和祭壇臺座的四角上，並內院的門框上。
EZEK|45|20|本月初七，你也要為誤犯罪的和因無知而犯罪的這樣做；你們要為聖殿贖罪。
EZEK|45|21|「正月十四日，你們要守逾越節，七天的節期都要吃無酵餅。
EZEK|45|22|當日，王要為自己和全國百姓預備一頭公牛作贖罪祭。
EZEK|45|23|節期的七天內，每天他要預備無殘疾的七頭公牛、七隻公綿羊，給耶和華為燔祭；每天又要預備一隻公山羊為贖罪祭。
EZEK|45|24|他也要預備素祭，為一頭公牛同獻一伊法細麵，為一隻公綿羊同獻一伊法細麵，每一伊法加一欣油。
EZEK|45|25|七月十五日守節的時候，七天他都要像這樣預備贖罪祭、燔祭、素祭和油。」
EZEK|46|1|主耶和華如此說：「內院朝東的門，在六個工作的日子必須關閉；惟有安息日和初一要敞開。
EZEK|46|2|王從外面要由門的走廊進入，站在門框旁邊；祭司要為他預備燔祭和平安祭，王要在門的門檻那裏敬拜，然後退出。這門直到晚上不可關閉。
EZEK|46|3|安息日和初一，這地的百姓要在這門口，在耶和華面前敬拜。
EZEK|46|4|安息日，王要用六隻無殘疾的羔羊、一隻無殘疾的公綿羊，獻給耶和華為燔祭；
EZEK|46|5|同獻的素祭，要為公綿羊獻一伊法細麵，為羔羊則按照他的力量獻，一伊法要加一欣油。
EZEK|46|6|初一，他要獻一頭無殘疾的公牛犢、六隻羔羊、一隻公綿羊，全都要用無殘疾的。
EZEK|46|7|他也要預備素祭，為公牛獻一伊法細麵，為公綿羊獻一伊法細麵，為羔羊則按照他的力量獻，一伊法要加一欣油。
EZEK|46|8|王進入的時候要由這門的走廊而入，也要從原路出去。
EZEK|46|9|「在各節期，這地的百姓朝見耶和華的時候，從北門進入敬拜的，要由南門而出；從南門進入的，要由北門而出。不可從進入的門出去，要往前直行，從對面的門出去。
EZEK|46|10|他們進入時，王也跟他們一同進入；他們出去，他也要出去。
EZEK|46|11|「在節期和盛會的日子同獻的素祭，要為一頭公牛獻一伊法細麵，為一隻公綿羊獻一伊法細麵，為羔羊則按照各人的力量獻，一伊法要加一欣油。
EZEK|46|12|王奉獻甘心祭，就是向耶和華甘心獻的燔祭或平安祭時，當有人為他開朝東的門。他就獻上燔祭和平安祭，與安息日所獻的一樣，然後退出。他出去之後，當有人將門關閉。」
EZEK|46|13|「每日，你要取一隻無殘疾一歲的羔羊獻給耶和華為燔祭；要每天早晨獻上。
EZEK|46|14|每天早晨你也要預備同獻的素祭，六分之一伊法細麵，並三分之一欣油，調和細麵。這素祭要經常獻給耶和華，作為永遠的定例。
EZEK|46|15|每天早晨要這樣獻上羔羊、素祭和油，為經常獻的燔祭。」
EZEK|46|16|主耶和華如此說：「王若將禮物賜給他的任何一個兒子，這就成為兒子的產業，可留給子孫，是他們所承受的地業。
EZEK|46|17|倘若王將他產業的一份賜給他的一個臣僕，這就成為他臣僕的產業，直到自由之年，然後地要歸還王；王的產業終究要歸自己的兒子。
EZEK|46|18|王不可奪取百姓的產業，以致趕逐他們離開自己的地業；他應該從自己的地業中將產業賜給子孫，免得我的子民離開自己的地業，四散各處。」
EZEK|46|19|他帶領我從大門旁邊的入口，進到朝北為祭司所預備聖的房間，看哪，西邊盡頭有一塊土地。
EZEK|46|20|他對我說：「這是祭司煮贖愆祭牲、贖罪祭牲，烤素祭的地方，免得帶出外院，使百姓成為聖。」
EZEK|46|21|他又帶我出到外院，使我經過院子的四個角落，看哪，院子的每個角落都有一個小院子。
EZEK|46|22|院子四個角落有小院子，周圍有牆，每個小院子長四十肘 ，寬三十肘；四個角落的小院子大小都一樣，
EZEK|46|23|小院子周圍各有一排石牆，每排石牆下面有爐灶。
EZEK|46|24|他對我說：「這些是煮肉用的屋子，殿內的僕役要在這裏煮百姓的祭物。」
EZEK|47|1|他帶我回到殿門，看哪，有水從殿的門檻下面往東流出，因為這殿是朝東的。水從殿的側面，就是右邊，從祭壇的南邊往下流。
EZEK|47|2|他帶我出北門，又領我從外邊轉到朝東的外門，看哪，水從右邊流出。
EZEK|47|3|他手拿繩子往東出去，量了一千肘，使我涉水而過，水到腳踝。
EZEK|47|4|他又量了一千，使我涉水而過，水就到膝；再量了一千，使我過去，水就到腰；
EZEK|47|5|又量了一千，水已成河，無法過去；因為水勢高漲成河，只能游泳，無法走過。
EZEK|47|6|他對我說：「人子啊，你看見了嗎？」 他帶我回到河邊。
EZEK|47|7|我回到河邊時，看哪，河這邊與那邊的岸上有極多的樹木。
EZEK|47|8|他對我說：「這水往東方流，下到 亞拉巴 ，直到海。所流出來的水，一入海 就使水變淡 。
EZEK|47|9|這兩條河 所到之處，凡滋生的動物都必存活；這水流到那裏，使那裏的水變淡，因此裏面有極多的魚。這河水所到之處，百物都必存活。
EZEK|47|10|必有漁夫站在河邊，從 隱‧基底 直到 隱‧以革蓮 ，全都成了曬 網的場所。那裏的魚各從其類，好像大海的魚甚多。
EZEK|47|11|但是沼澤與池塘的水無法變淡，只能作產鹽之用。
EZEK|47|12|河這邊與那邊的岸上必生長各類樹木，可作食物；葉子不枯乾，果子不斷絕。每月必結新果子，因為這水是從聖所流出來的。樹上的果子必作食物，葉子可以治病。」
EZEK|47|13|主耶和華如此說：「這是你們按 以色列 十二支派分地為業的地界， 約瑟 要得兩份。
EZEK|47|14|你們承受這地為業，要彼此均分；我曾起誓應許將這地賜給你們的列祖，這地必歸你們為業。
EZEK|47|15|「這地的疆界如下：北界從 大海 往 希特倫 ，直到 西達達 口；
EZEK|47|16|又往 哈馬 、 比羅他 、 西伯蓮 ( 西伯蓮 在 大馬士革 的邊界與 哈馬 的邊界中間)，到 浩蘭 邊界的 哈撒‧哈提干 。
EZEK|47|17|這樣，疆界是從 大海 往 大馬士革 地界上的 哈薩‧以難 ，北邊以 哈馬 為界。這是北界。
EZEK|47|18|「東界在 浩蘭 和 大馬士革 中間， 基列 和 以色列 地的中間，以 約旦河 為界。你們要量疆界直到東海 。這是東界。
EZEK|47|19|「南界是從 他瑪 到 加低斯 的 米利巴 水，經 埃及 溪谷 ，直到 大海 。這是南界。
EZEK|47|20|「西界就是 大海 ，從南界直到 哈馬口 對面。這是西界。
EZEK|47|21|「你們要為自己按 以色列 的支派分這地。
EZEK|47|22|要抽籤分這地為業，歸自己和那在你們中間寄居，生兒育女的外人。你們要看他們如本地出生的 以色列 人，他們要在 以色列 支派中與你們同得地業。
EZEK|47|23|外人寄居在哪個支派，你們就在哪裏將地業分給他們。這是主耶和華說的。」
EZEK|48|1|眾支派的名字如下：從北邊盡頭，由 希特倫 往 哈馬 口，到 大馬士革 地界上的 哈薩‧以難 。北邊靠著 哈馬 地，從東到西是 但 的一份。
EZEK|48|2|靠著 但 的地界，從東到西，是 亞設 的一份。
EZEK|48|3|靠著 亞設 的地界，從東到西，是 拿弗他利 的一份。
EZEK|48|4|靠著 拿弗他利 的地界，從東到西，是 瑪拿西 的一份。
EZEK|48|5|靠著 瑪拿西 的地界，從東到西，是 以法蓮 的一份。
EZEK|48|6|靠著 以法蓮 的地界，從東到西，是 呂便 的一份。
EZEK|48|7|靠著 呂便 的地界，從東到西，是 猶大 的一份。
EZEK|48|8|靠著 猶大 的地界，從東到西，必有你們所當獻的聖地，寬二萬五千肘 ；長短與各族從東到西所分的地相同，聖所當在其中。
EZEK|48|9|你們獻給耶和華的聖地要長二萬五千肘，寬一萬肘。
EZEK|48|10|這聖地要歸祭司，北長二萬五千肘，西寬一萬肘，東寬一萬肘，南長二萬五千肘。耶和華的聖所當在其中。
EZEK|48|11|這地要歸 撒督 的子孫中成為聖的祭司，他們謹守我所吩咐的；當 以色列 人走迷的時候，他們不像那些 利未 人走迷了。
EZEK|48|12|在聖地中要特別保留一份歸他們，為至聖，緊鄰著 利未 人的地界。
EZEK|48|13|利未 人所得的地長二萬五千肘，寬一萬肘，與祭司的地界相等，都長二萬五千肘，寬一萬肘。
EZEK|48|14|這地不可賣，不可換；這上好的部分不可轉讓給別人，因為它歸耶和華為聖。
EZEK|48|15|剩下的地長二萬五千肘、寬五千肘，要作公用，為造城、蓋房、空地之用；城要在中間。
EZEK|48|16|以下是城的大小：北面四千五百肘，南面四千五百肘，東面四千五百肘，西面四千五百肘。
EZEK|48|17|城要有空地，向北二百五十肘，向南二百五十肘，向東二百五十肘，向西二百五十肘。
EZEK|48|18|靠著聖地並排剩餘的，東長一萬肘，西長一萬肘；它與聖地並排，其中所出產的要作城內工人的食物。
EZEK|48|19|以色列 支派中所有在城內做工的，都要耕種這地。
EZEK|48|20|你們要將整塊四方的聖地，長二萬五千肘，寬二萬五千肘，連同城的用地都獻作聖地。
EZEK|48|21|聖地和城的用地兩邊剩餘的要歸給王。地的東邊，南北二萬五千肘，東至東界；西邊，南北二萬五千肘，西至西界；靠著各支派所分的地，都要歸給王。聖地和殿的聖所要在其中。
EZEK|48|22|利未 人的地與城的用地都在王的地中間， 猶大 邊界和 便雅憫 邊界之間，要歸給王。
EZEK|48|23|論到其餘的支派，從東到西，是 便雅憫 的一份。
EZEK|48|24|靠著 便雅憫 的地界，從東到西，是 西緬 的一份。
EZEK|48|25|靠著 西緬 的地界，從東到西，是 以薩迦 的一份。
EZEK|48|26|靠著 以薩迦 的地界，從東到西，是 西布倫 的一份。
EZEK|48|27|靠著 西布倫 的地界，從東到西，是 迦得 的一份。
EZEK|48|28|靠著 迦得 南邊的地界，界限從 他瑪 到 加低斯 的 米利巴 水，經 埃及 溪谷 ，直到 大海 。
EZEK|48|29|這就是你們要抽籤分給 以色列 支派為業之地，是他們各支派所得的份。這是主耶和華說的。
EZEK|48|30|以下是城的出口：北面四千五百肘，
EZEK|48|31|城的各門要按 以色列 的支派命名。北面有三個門，一為 呂便 門，一為 猶大 門，一為 利未 門。
EZEK|48|32|東面四千五百肘，有三個門，一為 約瑟 門，一為 便雅憫 門，一為 但 門。
EZEK|48|33|南面四千五百肘，有三個門，一為 西緬 門，一為 以薩迦 門，一為 西布倫 門。
EZEK|48|34|西面四千五百肘，有三個門，一為 迦得 門，一為 亞設 門，一為 拿弗他利 門。
EZEK|48|35|城的周圍共一萬八千肘。從此以後，這城的名字必稱為「耶和華的所在」。
