NUM|1|1|And the LORD spake unto Moses in the wilderness of Sinai, in the tabernacle of the congregation, on the first day of the second month, in the second year after they were come out of the land of Egypt, saying,
NUM|1|2|Take ye the sum of all the congregation of the children of Israel, after their families, by the house of their fathers, with the number of their names, every male by their polls;
NUM|1|3|From twenty years old and upward, all that are able to go forth to war in Israel: thou and Aaron shall number them by their armies.
NUM|1|4|And with you there shall be a man of every tribe; every one head of the house of his fathers.
NUM|1|5|And these are the names of the men that shall stand with you: of the tribe of Reuben; Elizur the son of Shedeur.
NUM|1|6|Of Simeon; Shelumiel the son of Zurishaddai.
NUM|1|7|Of Judah; Nahshon the son of Amminadab.
NUM|1|8|Of Issachar; Nethaneel the son of Zuar.
NUM|1|9|Of Zebulun; Eliab the son of Helon.
NUM|1|10|Of the children of Joseph: of Ephraim; Elishama the son of Ammihud: of Manasseh; Gamaliel the son of Pedahzur.
NUM|1|11|Of Benjamin; Abidan the son of Gideoni.
NUM|1|12|Of Dan; Ahiezer the son of Ammishaddai.
NUM|1|13|Of Asher; Pagiel the son of Ocran.
NUM|1|14|Of Gad; Eliasaph the son of Deuel.
NUM|1|15|Of Naphtali; Ahira the son of Enan.
NUM|1|16|These were the renowned of the congregation, princes of the tribes of their fathers, heads of thousands in Israel.
NUM|1|17|And Moses and Aaron took these men which are expressed by their names:
NUM|1|18|And they assembled all the congregation together on the first day of the second month, and they declared their pedigrees after their families, by the house of their fathers, according to the number of the names, from twenty years old and upward, by their polls.
NUM|1|19|As the LORD commanded Moses, so he numbered them in the wilderness of Sinai.
NUM|1|20|And the children of Reuben, Israel's eldest son, by their generations, after their families, by the house of their fathers, according to the number of the names, by their polls, every male from twenty years old and upward, all that were able to go forth to war;
NUM|1|21|Those that were numbered of them, even of the tribe of Reuben, were forty and six thousand and five hundred.
NUM|1|22|Of the children of Simeon, by their generations, after their families, by the house of their fathers, those that were numbered of them, according to the number of the names, by their polls, every male from twenty years old and upward, all that were able to go forth to war;
NUM|1|23|Those that were numbered of them, even of the tribe of Simeon, were fifty and nine thousand and three hundred.
NUM|1|24|Of the children of Gad, by their generations, after their families, by the house of their fathers, according to the number of the names, from twenty years old and upward, all that were able to go forth to war;
NUM|1|25|Those that were numbered of them, even of the tribe of Gad, were forty and five thousand six hundred and fifty.
NUM|1|26|Of the children of Judah, by their generations, after their families, by the house of their fathers, according to the number of the names, from twenty years old and upward, all that were able to go forth to war;
NUM|1|27|Those that were numbered of them, even of the tribe of Judah, were threescore and fourteen thousand and six hundred.
NUM|1|28|Of the children of Issachar, by their generations, after their families, by the house of their fathers, according to the number of the names, from twenty years old and upward, all that were able to go forth to war;
NUM|1|29|Those that were numbered of them, even of the tribe of Issachar, were fifty and four thousand and four hundred.
NUM|1|30|Of the children of Zebulun, by their generations, after their families, by the house of their fathers, according to the number of the names, from twenty years old and upward, all that were able to go forth to war;
NUM|1|31|Those that were numbered of them, even of the tribe of Zebulun, were fifty and seven thousand and four hundred.
NUM|1|32|Of the children of Joseph, namely, of the children of Ephraim, by their generations, after their families, by the house of their fathers, according to the number of the names, from twenty years old and upward, all that were able to go forth to war;
NUM|1|33|Those that were numbered of them, even of the tribe of Ephraim, were forty thousand and five hundred.
NUM|1|34|Of the children of Manasseh, by their generations, after their families, by the house of their fathers, according to the number of the names, from twenty years old and upward, all that were able to go forth to war;
NUM|1|35|Those that were numbered of them, even of the tribe of Manasseh, were thirty and two thousand and two hundred.
NUM|1|36|Of the children of Benjamin, by their generations, after their families, by the house of their fathers, according to the number of the names, from twenty years old and upward, all that were able to go forth to war;
NUM|1|37|Those that were numbered of them, even of the tribe of Benjamin, were thirty and five thousand and four hundred.
NUM|1|38|Of the children of Dan, by their generations, after their families, by the house of their fathers, according to the number of the names, from twenty years old and upward, all that were able to go forth to war;
NUM|1|39|Those that were numbered of them, even of the tribe of Dan, were threescore and two thousand and seven hundred.
NUM|1|40|Of the children of Asher, by their generations, after their families, by the house of their fathers, according to the number of the names, from twenty years old and upward, all that were able to go forth to war;
NUM|1|41|Those that were numbered of them, even of the tribe of Asher, were forty and one thousand and five hundred.
NUM|1|42|Of the children of Naphtali, throughout their generations, after their families, by the house of their fathers, according to the number of the names, from twenty years old and upward, all that were able to go forth to war;
NUM|1|43|Those that were numbered of them, even of the tribe of Naphtali, were fifty and three thousand and four hundred.
NUM|1|44|These are those that were numbered, which Moses and Aaron numbered, and the princes of Israel, being twelve men: each one was for the house of his fathers.
NUM|1|45|So were all those that were numbered of the children of Israel, by the house of their fathers, from twenty years old and upward, all that were able to go forth to war in Israel;
NUM|1|46|Even all they that were numbered were six hundred thousand and three thousand and five hundred and fifty.
NUM|1|47|But the Levites after the tribe of their fathers were not numbered among them.
NUM|1|48|For the LORD had spoken unto Moses, saying,
NUM|1|49|Only thou shalt not number the tribe of Levi, neither take the sum of them among the children of Israel:
NUM|1|50|But thou shalt appoint the Levites over the tabernacle of testimony, and over all the vessels thereof, and over all things that belong to it: they shall bear the tabernacle, and all the vessels thereof; and they shall minister unto it, and shall encamp round about the tabernacle.
NUM|1|51|And when the tabernacle setteth forward, the Levites shall take it down: and when the tabernacle is to be pitched, the Levites shall set it up: and the stranger that cometh nigh shall be put to death.
NUM|1|52|And the children of Israel shall pitch their tents, every man by his own camp, and every man by his own standard, throughout their hosts.
NUM|1|53|But the Levites shall pitch round about the tabernacle of testimony, that there be no wrath upon the congregation of the children of Israel: and the Levites shall keep the charge of the tabernacle of testimony.
NUM|1|54|And the children of Israel did according to all that the LORD commanded Moses, so did they.
NUM|2|1|And the LORD spake unto Moses and unto Aaron, saying,
NUM|2|2|Every man of the children of Israel shall pitch by his own standard, with the ensign of their father's house: far off about the tabernacle of the congregation shall they pitch.
NUM|2|3|And on the east side toward the rising of the sun shall they of the standard of the camp of Judah pitch throughout their armies: and Nahshon the son of Amminadab shall be captain of the children of Judah.
NUM|2|4|And his host, and those that were numbered of them, were threescore and fourteen thousand and six hundred.
NUM|2|5|And those that do pitch next unto him shall be the tribe of Issachar: and Nethaneel the son of Zuar shall be captain of the children of Issachar.
NUM|2|6|And his host, and those that were numbered thereof, were fifty and four thousand and four hundred.
NUM|2|7|Then the tribe of Zebulun: and Eliab the son of Helon shall be captain of the children of Zebulun.
NUM|2|8|And his host, and those that were numbered thereof, were fifty and seven thousand and four hundred.
NUM|2|9|All that were numbered in the camp of Judah were an hundred thousand and fourscore thousand and six thousand and four hundred, throughout their armies. These shall first set forth.
NUM|2|10|On the south side shall be the standard of the camp of Reuben according to their armies: and the captain of the children of Reuben shall be Elizur the son of Shedeur.
NUM|2|11|And his host, and those that were numbered thereof, were forty and six thousand and five hundred.
NUM|2|12|And those which pitch by him shall be the tribe of Simeon: and the captain of the children of Simeon shall be Shelumiel the son of Zurishaddai.
NUM|2|13|And his host, and those that were numbered of them, were fifty and nine thousand and three hundred.
NUM|2|14|Then the tribe of Gad: and the captain of the sons of Gad shall be Eliasaph the son of Reuel.
NUM|2|15|And his host, and those that were numbered of them, were forty and five thousand and six hundred and fifty.
NUM|2|16|All that were numbered in the camp of Reuben were an hundred thousand and fifty and one thousand and four hundred and fifty, throughout their armies. And they shall set forth in the second rank.
NUM|2|17|Then the tabernacle of the congregation shall set forward with the camp of the Levites in the midst of the camp: as they encamp, so shall they set forward, every man in his place by their standards.
NUM|2|18|On the west side shall be the standard of the camp of Ephraim according to their armies: and the captain of the sons of Ephraim shall be Elishama the son of Ammihud.
NUM|2|19|And his host, and those that were numbered of them, were forty thousand and five hundred.
NUM|2|20|And by him shall be the tribe of Manasseh: and the captain of the children of Manasseh shall be Gamaliel the son of Pedahzur.
NUM|2|21|And his host, and those that were numbered of them, were thirty and two thousand and two hundred.
NUM|2|22|Then the tribe of Benjamin: and the captain of the sons of Benjamin shall be Abidan the son of Gideoni.
NUM|2|23|And his host, and those that were numbered of them, were thirty and five thousand and four hundred.
NUM|2|24|All that were numbered of the camp of Ephraim were an hundred thousand and eight thousand and an hundred, throughout their armies. And they shall go forward in the third rank.
NUM|2|25|The standard of the camp of Dan shall be on the north side by their armies: and the captain of the children of Dan shall be Ahiezer the son of Ammishaddai.
NUM|2|26|And his host, and those that were numbered of them, were threescore and two thousand and seven hundred.
NUM|2|27|And those that encamp by him shall be the tribe of Asher: and the captain of the children of Asher shall be Pagiel the son of Ocran.
NUM|2|28|And his host, and those that were numbered of them, were forty and one thousand and five hundred.
NUM|2|29|Then the tribe of Naphtali: and the captain of the children of Naphtali shall be Ahira the son of Enan.
NUM|2|30|And his host, and those that were numbered of them, were fifty and three thousand and four hundred.
NUM|2|31|All they that were numbered in the camp of Dan were an hundred thousand and fifty and seven thousand and six hundred. They shall go hindmost with their standards.
NUM|2|32|These are those which were numbered of the children of Israel by the house of their fathers: all those that were numbered of the camps throughout their hosts were six hundred thousand and three thousand and five hundred and fifty.
NUM|2|33|But the Levites were not numbered among the children of Israel; as the LORD commanded Moses.
NUM|2|34|And the children of Israel did according to all that the LORD commanded Moses: so they pitched by their standards, and so they set forward, every one after their families, according to the house of their fathers.
NUM|3|1|These also are the generations of Aaron and Moses in the day that the LORD spake with Moses in mount Sinai.
NUM|3|2|And these are the names of the sons of Aaron; Nadab the firstborn, and Abihu, Eleazar, and Ithamar.
NUM|3|3|These are the names of the sons of Aaron, the priests which were anointed, whom he consecrated to minister in the priest's office.
NUM|3|4|And Nadab and Abihu died before the LORD, when they offered strange fire before the LORD, in the wilderness of Sinai, and they had no children: and Eleazar and Ithamar ministered in the priest's office in the sight of Aaron their father.
NUM|3|5|And the LORD spake unto Moses, saying,
NUM|3|6|Bring the tribe of Levi near, and present them before Aaron the priest, that they may minister unto him.
NUM|3|7|And they shall keep his charge, and the charge of the whole congregation before the tabernacle of the congregation, to do the service of the tabernacle.
NUM|3|8|And they shall keep all the instruments of the tabernacle of the congregation, and the charge of the children of Israel, to do the service of the tabernacle.
NUM|3|9|And thou shalt give the Levites unto Aaron and to his sons: they are wholly given unto him out of the children of Israel.
NUM|3|10|And thou shalt appoint Aaron and his sons, and they shall wait on their priest's office: and the stranger that cometh nigh shall be put to death.
NUM|3|11|And the LORD spake unto Moses, saying,
NUM|3|12|And I, behold, I have taken the Levites from among the children of Israel instead of all the firstborn that openeth the matrix among the children of Israel: therefore the Levites shall be mine;
NUM|3|13|Because all the firstborn are mine; for on the day that I smote all the firstborn in the land of Egypt I hallowed unto me all the firstborn in Israel, both man and beast: mine shall they be: I am the LORD.
NUM|3|14|And the LORD spake unto Moses in the wilderness of Sinai, saying,
NUM|3|15|Number the children of Levi after the house of their fathers, by their families: every male from a month old and upward shalt thou number them.
NUM|3|16|And Moses numbered them according to the word of the LORD, as he was commanded.
NUM|3|17|And these were the sons of Levi by their names; Gershon, and Kohath, and Merari.
NUM|3|18|And these are the names of the sons of Gershon by their families; Libni, and Shimei.
NUM|3|19|And the sons of Kohath by their families; Amram, and Izehar, Hebron, and Uzziel.
NUM|3|20|And the sons of Merari by their families; Mahli, and Mushi. These are the families of the Levites according to the house of their fathers.
NUM|3|21|Of Gershon was the family of the Libnites, and the family of the Shimites: these are the families of the Gershonites.
NUM|3|22|Those that were numbered of them, according to the number of all the males, from a month old and upward, even those that were numbered of them were seven thousand and five hundred.
NUM|3|23|The families of the Gershonites shall pitch behind the tabernacle westward.
NUM|3|24|And the chief of the house of the father of the Gershonites shall be Eliasaph the son of Lael.
NUM|3|25|And the charge of the sons of Gershon in the tabernacle of the congregation shall be the tabernacle, and the tent, the covering thereof, and the hanging for the door of the tabernacle of the congregation,
NUM|3|26|And the hangings of the court, and the curtain for the door of the court, which is by the tabernacle, and by the altar round about, and the cords of it for all the service thereof.
NUM|3|27|And of Kohath was the family of the Amramites, and the family of the Izeharites, and the family of the Hebronites, and the family of the Uzzielites: these are the families of the Kohathites.
NUM|3|28|In the number of all the males, from a month old and upward, were eight thousand and six hundred, keeping the charge of the sanctuary.
NUM|3|29|The families of the sons of Kohath shall pitch on the side of the tabernacle southward.
NUM|3|30|And the chief of the house of the father of the families of the Kohathites shall be Elizaphan the son of Uzziel.
NUM|3|31|And their charge shall be the ark, and the table, and the candlestick, and the altars, and the vessels of the sanctuary wherewith they minister, and the hanging, and all the service thereof.
NUM|3|32|And Eleazar the son of Aaron the priest shall be chief over the chief of the Levites, and have the oversight of them that keep the charge of the sanctuary.
NUM|3|33|Of Merari was the family of the Mahlites, and the family of the Mushites: these are the families of Merari.
NUM|3|34|And those that were numbered of them, according to the number of all the males, from a month old and upward, were six thousand and two hundred.
NUM|3|35|And the chief of the house of the father of the families of Merari was Zuriel the son of Abihail: these shall pitch on the side of the tabernacle northward.
NUM|3|36|And under the custody and charge of the sons of Merari shall be the boards of the tabernacle, and the bars thereof, and the pillars thereof, and the sockets thereof, and all the vessels thereof, and all that serveth thereto,
NUM|3|37|And the pillars of the court round about, and their sockets, and their pins, and their cords.
NUM|3|38|But those that encamp before the tabernacle toward the east, even before the tabernacle of the congregation eastward, shall be Moses, and Aaron and his sons, keeping the charge of the sanctuary for the charge of the children of Israel; and the stranger that cometh nigh shall be put to death.
NUM|3|39|All that were numbered of the Levites, which Moses and Aaron numbered at the commandment of the LORD, throughout their families, all the males from a month old and upward, were twenty and two thousand.
NUM|3|40|And the LORD said unto Moses, Number all the firstborn of the males of the children of Israel from a month old and upward, and take the number of their names.
NUM|3|41|And thou shalt take the Levites for me (I am the LORD) instead of all the firstborn among the children of Israel; and the cattle of the Levites instead of all the firstlings among the cattle of the children of Israel.
NUM|3|42|And Moses numbered, as the LORD commanded him, all the firstborn among the children of Israel.
NUM|3|43|And all the firstborn males by the number of names, from a month old and upward, of those that were numbered of them, were twenty and two thousand two hundred and threescore and thirteen.
NUM|3|44|And the LORD spake unto Moses, saying,
NUM|3|45|Take the Levites instead of all the firstborn among the children of Israel, and the cattle of the Levites instead of their cattle; and the Levites shall be mine: I am the LORD.
NUM|3|46|And for those that are to be redeemed of the two hundred and threescore and thirteen of the firstborn of the children of Israel, which are more than the Levites;
NUM|3|47|Thou shalt even take five shekels apiece by the poll, after the shekel of the sanctuary shalt thou take them: (the shekel is twenty gerahs:)
NUM|3|48|And thou shalt give the money, wherewith the odd number of them is to be redeemed, unto Aaron and to his sons.
NUM|3|49|And Moses took the redemption money of them that were over and above them that were redeemed by the Levites:
NUM|3|50|Of the firstborn of the children of Israel took he the money; a thousand three hundred and threescore and five shekels, after the shekel of the sanctuary:
NUM|3|51|And Moses gave the money of them that were redeemed unto Aaron and to his sons, according to the word of the LORD, as the LORD commanded Moses.
NUM|4|1|And the LORD spake unto Moses and unto Aaron, saying,
NUM|4|2|Take the sum of the sons of Kohath from among the sons of Levi, after their families, by the house of their fathers,
NUM|4|3|From thirty years old and upward even until fifty years old, all that enter into the host, to do the work in the tabernacle of the congregation.
NUM|4|4|This shall be the service of the sons of Kohath in the tabernacle of the congregation, about the most holy things:
NUM|4|5|And when the camp setteth forward, Aaron shall come, and his sons, and they shall take down the covering vail, and cover the ark of testimony with it:
NUM|4|6|And shall put thereon the covering of badgers' skins, and shall spread over it a cloth wholly of blue, and shall put in the staves thereof.
NUM|4|7|And upon the table of showbread they shall spread a cloth of blue, and put thereon the dishes, and the spoons, and the bowls, and covers to cover withal: and the continual bread shall be thereon:
NUM|4|8|And they shall spread upon them a cloth of scarlet, and cover the same with a covering of badgers' skins, and shall put in the staves thereof.
NUM|4|9|And they shall take a cloth of blue, and cover the candlestick of the light, and his lamps, and his tongs, and his snuffdishes, and all the oil vessels thereof, wherewith they minister unto it:
NUM|4|10|And they shall put it and all the vessels thereof within a covering of badgers' skins, and shall put it upon a bar.
NUM|4|11|And upon the golden altar they shall spread a cloth of blue, and cover it with a covering of badgers' skins, and shall put to the staves thereof:
NUM|4|12|And they shall take all the instruments of ministry, wherewith they minister in the sanctuary, and put them in a cloth of blue, and cover them with a covering of badgers' skins, and shall put them on a bar:
NUM|4|13|And they shall take away the ashes from the altar, and spread a purple cloth thereon:
NUM|4|14|And they shall put upon it all the vessels thereof, wherewith they minister about it, even the censers, the fleshhooks, and the shovels, and the basins, all the vessels of the altar; and they shall spread upon it a covering of badgers' skins, and put to the staves of it.
NUM|4|15|And when Aaron and his sons have made an end of covering the sanctuary, and all the vessels of the sanctuary, as the camp is to set forward; after that, the sons of Kohath shall come to bear it: but they shall not touch any holy thing, lest they die. These things are the burden of the sons of Kohath in the tabernacle of the congregation.
NUM|4|16|And to the office of Eleazar the son of Aaron the priest pertaineth the oil for the light, and the sweet incense, and the daily meat offering, and the anointing oil, and the oversight of all the tabernacle, and of all that therein is, in the sanctuary, and in the vessels thereof.
NUM|4|17|And the LORD spake unto Moses and unto Aaron saying,
NUM|4|18|Cut ye not off the tribe of the families of the Kohathites from among the Levites:
NUM|4|19|But thus do unto them, that they may live, and not die, when they approach unto the most holy things: Aaron and his sons shall go in, and appoint them every one to his service and to his burden:
NUM|4|20|But they shall not go in to see when the holy things are covered, lest they die.
NUM|4|21|And the LORD spake unto Moses, saying,
NUM|4|22|Take also the sum of the sons of Gershon, throughout the houses of their fathers, by their families;
NUM|4|23|From thirty years old and upward until fifty years old shalt thou number them; all that enter in to perform the service, to do the work in the tabernacle of the congregation.
NUM|4|24|This is the service of the families of the Gershonites, to serve, and for burdens:
NUM|4|25|And they shall bear the curtains of the tabernacle, and the tabernacle of the congregation, his covering, and the covering of the badgers' skins that is above upon it, and the hanging for the door of the tabernacle of the congregation,
NUM|4|26|And the hangings of the court, and the hanging for the door of the gate of the court, which is by the tabernacle and by the altar round about, and their cords, and all the instruments of their service, and all that is made for them: so shall they serve.
NUM|4|27|At the appointment of Aaron and his sons shall be all the service of the sons of the Gershonites, in all their burdens, and in all their service: and ye shall appoint unto them in charge all their burdens.
NUM|4|28|This is the service of the families of the sons of Gershon in the tabernacle of the congregation: and their charge shall be under the hand of Ithamar the son of Aaron the priest.
NUM|4|29|As for the sons of Merari, thou shalt number them after their families, by the house of their fathers;
NUM|4|30|From thirty years old and upward even unto fifty years old shalt thou number them, every one that entereth into the service, to do the work of the tabernacle of the congregation.
NUM|4|31|And this is the charge of their burden, according to all their service in the tabernacle of the congregation; the boards of the tabernacle, and the bars thereof, and the pillars thereof, and sockets thereof,
NUM|4|32|And the pillars of the court round about, and their sockets, and their pins, and their cords, with all their instruments, and with all their service: and by name ye shall reckon the instruments of the charge of their burden.
NUM|4|33|This is the service of the families of the sons of Merari, according to all their service, in the tabernacle of the congregation, under the hand of Ithamar the son of Aaron the priest.
NUM|4|34|And Moses and Aaron and the chief of the congregation numbered the sons of the Kohathites after their families, and after the house of their fathers,
NUM|4|35|From thirty years old and upward even unto fifty years old, every one that entereth into the service, for the work in the tabernacle of the congregation:
NUM|4|36|And those that were numbered of them by their families were two thousand seven hundred and fifty.
NUM|4|37|These were they that were numbered of the families of the Kohathites, all that might do service in the tabernacle of the congregation, which Moses and Aaron did number according to the commandment of the LORD by the hand of Moses.
NUM|4|38|And those that were numbered of the sons of Gershon, throughout their families, and by the house of their fathers,
NUM|4|39|From thirty years old and upward even unto fifty years old, every one that entereth into the service, for the work in the tabernacle of the congregation,
NUM|4|40|Even those that were numbered of them, throughout their families, by the house of their fathers, were two thousand and six hundred and thirty.
NUM|4|41|These are they that were numbered of the families of the sons of Gershon, of all that might do service in the tabernacle of the congregation, whom Moses and Aaron did number according to the commandment of the LORD.
NUM|4|42|And those that were numbered of the families of the sons of Merari, throughout their families, by the house of their fathers,
NUM|4|43|From thirty years old and upward even unto fifty years old, every one that entereth into the service, for the work in the tabernacle of the congregation,
NUM|4|44|Even those that were numbered of them after their families, were three thousand and two hundred.
NUM|4|45|These be those that were numbered of the families of the sons of Merari, whom Moses and Aaron numbered according to the word of the LORD by the hand of Moses.
NUM|4|46|All those that were numbered of the Levites, whom Moses and Aaron and the chief of Israel numbered, after their families, and after the house of their fathers,
NUM|4|47|From thirty years old and upward even unto fifty years old, every one that came to do the service of the ministry, and the service of the burden in the tabernacle of the congregation.
NUM|4|48|Even those that were numbered of them, were eight thousand and five hundred and fourscore,
NUM|4|49|According to the commandment of the LORD they were numbered by the hand of Moses, every one according to his service, and according to his burden: thus were they numbered of him, as the LORD commanded Moses.
NUM|5|1|And the LORD spake unto Moses, saying,
NUM|5|2|Command the children of Israel, that they put out of the camp every leper, and every one that hath an issue, and whosoever is defiled by the dead:
NUM|5|3|Both male and female shall ye put out, without the camp shall ye put them; that they defile not their camps, in the midst whereof I dwell.
NUM|5|4|And the children of Israel did so, and put them out without the camp: as the LORD spake unto Moses, so did the children of Israel.
NUM|5|5|And the LORD spake unto Moses, saying,
NUM|5|6|Speak unto the children of Israel, When a man or woman shall commit any sin that men commit, to do a trespass against the LORD, and that person be guilty;
NUM|5|7|Then they shall confess their sin which they have done: and he shall recompense his trespass with the principal thereof, and add unto it the fifth part thereof, and give it unto him against whom he hath trespassed.
NUM|5|8|But if the man have no kinsman to recompense the trespass unto, let the trespass be recompensed unto the LORD, even to the priest; beside the ram of the atonement, whereby an atonement shall be made for him.
NUM|5|9|And every offering of all the holy things of the children of Israel, which they bring unto the priest, shall be his.
NUM|5|10|And every man's hallowed things shall be his: whatsoever any man giveth the priest, it shall be his.
NUM|5|11|And the LORD spake unto Moses, saying,
NUM|5|12|Speak unto the children of Israel, and say unto them, If any man's wife go aside, and commit a trespass against him,
NUM|5|13|And a man lie with her carnally, and it be hid from the eyes of her husband, and be kept close, and she be defiled, and there be no witness against her, neither she be taken with the manner;
NUM|5|14|And the spirit of jealousy come upon him, and he be jealous of his wife, and she be defiled: or if the spirit of jealousy come upon him, and he be jealous of his wife, and she be not defiled:
NUM|5|15|Then shall the man bring his wife unto the priest, and he shall bring her offering for her, the tenth part of an ephah of barley meal; he shall pour no oil upon it, nor put frankincense thereon; for it is an offering of jealousy, an offering of memorial, bringing iniquity to remembrance.
NUM|5|16|And the priest shall bring her near, and set her before the LORD:
NUM|5|17|And the priest shall take holy water in an earthen vessel; and of the dust that is in the floor of the tabernacle the priest shall take, and put it into the water:
NUM|5|18|And the priest shall set the woman before the LORD, and uncover the woman's head, and put the offering of memorial in her hands, which is the jealousy offering: and the priest shall have in his hand the bitter water that causeth the curse:
NUM|5|19|And the priest shall charge her by an oath, and say unto the woman, If no man have lain with thee, and if thou hast not gone aside to uncleanness with another instead of thy husband, be thou free from this bitter water that causeth the curse:
NUM|5|20|But if thou hast gone aside to another instead of thy husband, and if thou be defiled, and some man have lain with thee beside thine husband:
NUM|5|21|Then the priest shall charge the woman with an oath of cursing, and the priest shall say unto the woman, The LORD make thee a curse and an oath among thy people, when the LORD doth make thy thigh to rot, and thy belly to swell;
NUM|5|22|And this water that causeth the curse shall go into thy bowels, to make thy belly to swell, and thy thigh to rot: And the woman shall say, Amen, amen.
NUM|5|23|And the priest shall write these curses in a book, and he shall blot them out with the bitter water:
NUM|5|24|And he shall cause the woman to drink the bitter water that causeth the curse: and the water that causeth the curse shall enter into her, and become bitter.
NUM|5|25|Then the priest shall take the jealousy offering out of the woman's hand, and shall wave the offering before the LORD, and offer it upon the altar:
NUM|5|26|And the priest shall take an handful of the offering, even the memorial thereof, and burn it upon the altar, and afterward shall cause the woman to drink the water.
NUM|5|27|And when he hath made her to drink the water, then it shall come to pass, that, if she be defiled, and have done trespass against her husband, that the water that causeth the curse shall enter into her, and become bitter, and her belly shall swell, and her thigh shall rot: and the woman shall be a curse among her people.
NUM|5|28|And if the woman be not defiled, but be clean; then she shall be free, and shall conceive seed.
NUM|5|29|This is the law of jealousies, when a wife goeth aside to another instead of her husband, and is defiled;
NUM|5|30|Or when the spirit of jealousy cometh upon him, and he be jealous over his wife, and shall set the woman before the LORD, and the priest shall execute upon her all this law.
NUM|5|31|Then shall the man be guiltless from iniquity, and this woman shall bear her iniquity.
NUM|6|1|And the LORD spake unto Moses, saying,
NUM|6|2|Speak unto the children of Israel, and say unto them, When either man or woman shall separate themselves to vow a vow of a Nazarite, to separate themselves unto the LORD:
NUM|6|3|He shall separate himself from wine and strong drink, and shall drink no vinegar of wine, or vinegar of strong drink, neither shall he drink any liquor of grapes, nor eat moist grapes, or dried.
NUM|6|4|All the days of his separation shall he eat nothing that is made of the vine tree, from the kernels even to the husk.
NUM|6|5|All the days of the vow of his separation there shall no razor come upon his head: until the days be fulfilled, in the which he separateth himself unto the LORD, he shall be holy, and shall let the locks of the hair of his head grow.
NUM|6|6|All the days that he separateth himself unto the LORD he shall come at no dead body.
NUM|6|7|He shall not make himself unclean for his father, or for his mother, for his brother, or for his sister, when they die: because the consecration of his God is upon his head.
NUM|6|8|All the days of his separation he is holy unto the LORD.
NUM|6|9|And if any man die very suddenly by him, and he hath defiled the head of his consecration; then he shall shave his head in the day of his cleansing, on the seventh day shall he shave it.
NUM|6|10|And on the eighth day he shall bring two turtles, or two young pigeons, to the priest, to the door of the tabernacle of the congregation:
NUM|6|11|And the priest shall offer the one for a sin offering, and the other for a burnt offering, and make an atonement for him, for that he sinned by the dead, and shall hallow his head that same day.
NUM|6|12|And he shall consecrate unto the LORD the days of his separation, and shall bring a lamb of the first year for a trespass offering: but the days that were before shall be lost, because his separation was defiled.
NUM|6|13|And this is the law of the Nazarite, when the days of his separation are fulfilled: he shall be brought unto the door of the tabernacle of the congregation:
NUM|6|14|And he shall offer his offering unto the LORD, one he lamb of the first year without blemish for a burnt offering, and one ewe lamb of the first year without blemish for a sin offering, and one ram without blemish for peace offerings,
NUM|6|15|And a basket of unleavened bread, cakes of fine flour mingled with oil, and wafers of unleavened bread anointed with oil, and their meat offering, and their drink offerings.
NUM|6|16|And the priest shall bring them before the LORD, and shall offer his sin offering, and his burnt offering:
NUM|6|17|And he shall offer the ram for a sacrifice of peace offerings unto the LORD, with the basket of unleavened bread: the priest shall offer also his meat offering, and his drink offering.
NUM|6|18|And the Nazarite shall shave the head of his separation at the door of the tabernacle of the congregation, and shall take the hair of the head of his separation, and put it in the fire which is under the sacrifice of the peace offerings.
NUM|6|19|And the priest shall take the sodden shoulder of the ram, and one unleavened cake out of the basket, and one unleavened wafer, and shall put them upon the hands of the Nazarite, after the hair of his separation is shaven:
NUM|6|20|And the priest shall wave them for a wave offering before the LORD: this is holy for the priest, with the wave breast and heave shoulder: and after that the Nazarite may drink wine.
NUM|6|21|This is the law of the Nazarite who hath vowed, and of his offering unto the LORD for his separation, beside that that his hand shall get: according to the vow which he vowed, so he must do after the law of his separation.
NUM|6|22|And the LORD spake unto Moses, saying,
NUM|6|23|Speak unto Aaron and unto his sons, saying, On this wise ye shall bless the children of Israel, saying unto them,
NUM|6|24|The LORD bless thee, and keep thee:
NUM|6|25|The LORD make his face shine upon thee, and be gracious unto thee:
NUM|6|26|The LORD lift up his countenance upon thee, and give thee peace.
NUM|6|27|And they shall put my name upon the children of Israel, and I will bless them.
NUM|7|1|And it came to pass on the day that Moses had fully set up the tabernacle, and had anointed it, and sanctified it, and all the instruments thereof, both the altar and all the vessels thereof, and had anointed them, and sanctified them;
NUM|7|2|That the princes of Israel, heads of the house of their fathers, who were the princes of the tribes, and were over them that were numbered, offered:
NUM|7|3|And they brought their offering before the LORD, six covered wagons, and twelve oxen; a wagon for two of the princes, and for each one an ox: and they brought them before the tabernacle.
NUM|7|4|And the LORD spake unto Moses, saying,
NUM|7|5|Take it of them, that they may be to do the service of the tabernacle of the congregation; and thou shalt give them unto the Levites, to every man according to his service.
NUM|7|6|And Moses took the wagons and the oxen, and gave them unto the Levites.
NUM|7|7|Two wagons and four oxen he gave unto the sons of Gershon, according to their service:
NUM|7|8|And four wagons and eight oxen he gave unto the sons of Merari, according unto their service, under the hand of Ithamar the son of Aaron the priest.
NUM|7|9|But unto the sons of Kohath he gave none: because the service of the sanctuary belonging unto them was that they should bear upon their shoulders.
NUM|7|10|And the princes offered for dedicating of the altar in the day that it was anointed, even the princes offered their offering before the altar.
NUM|7|11|And the LORD said unto Moses, They shall offer their offering, each prince on his day, for the dedicating of the altar.
NUM|7|12|And he that offered his offering the first day was Nahshon the son of Amminadab, of the tribe of Judah:
NUM|7|13|And his offering was one silver charger, the weight thereof was an hundred and thirty shekels, one silver bowl of seventy shekels, after the shekel of the sanctuary; both of them were full of fine flour mingled with oil for a meat offering:
NUM|7|14|One spoon of ten shekels of gold, full of incense:
NUM|7|15|One young bullock, one ram, one lamb of the first year, for a burnt offering:
NUM|7|16|One kid of the goats for a sin offering:
NUM|7|17|And for a sacrifice of peace offerings, two oxen, five rams, five he goats, five lambs of the first year: this was the offering of Nahshon the son of Amminadab.
NUM|7|18|On the second day Nethaneel the son of Zuar, prince of Issachar, did offer:
NUM|7|19|He offered for his offering one silver charger, the weight whereof was an hundred and thirty shekels, one silver bowl of seventy shekels, after the shekel of the sanctuary; both of them full of fine flour mingled with oil for a meat offering:
NUM|7|20|One spoon of gold of ten shekels, full of incense:
NUM|7|21|One young bullock, one ram, one lamb of the first year, for a burnt offering:
NUM|7|22|One kid of the goats for a sin offering:
NUM|7|23|And for a sacrifice of peace offerings, two oxen, five rams, five he goats, five lambs of the first year: this was the offering of Nethaneel the son of Zuar.
NUM|7|24|On the third day Eliab the son of Helon, prince of the children of Zebulun, did offer:
NUM|7|25|His offering was one silver charger, the weight whereof was an hundred and thirty shekels, one silver bowl of seventy shekels, after the shekel of the sanctuary; both of them full of fine flour mingled with oil for a meat offering:
NUM|7|26|One golden spoon of ten shekels, full of incense:
NUM|7|27|One young bullock, one ram, one lamb of the first year, for a burnt offering:
NUM|7|28|One kid of the goats for a sin offering:
NUM|7|29|And for a sacrifice of peace offerings, two oxen, five rams, five he goats, five lambs of the first year: this was the offering of Eliab the son of Helon.
NUM|7|30|On the fourth day Elizur the son of Shedeur, prince of the children of Reuben, did offer:
NUM|7|31|His offering was one silver charger of the weight of an hundred and thirty shekels, one silver bowl of seventy shekels, after the shekel of the sanctuary; both of them full of fine flour mingled with oil for a meat offering:
NUM|7|32|One golden spoon of ten shekels, full of incense:
NUM|7|33|One young bullock, one ram, one lamb of the first year, for a burnt offering:
NUM|7|34|One kid of the goats for a sin offering:
NUM|7|35|And for a sacrifice of peace offerings, two oxen, five rams, five he goats, five lambs of the first year: this was the offering of Elizur the son of Shedeur.
NUM|7|36|On the fifth day Shelumiel the son of Zurishaddai, prince of the children of Simeon, did offer:
NUM|7|37|His offering was one silver charger, the weight whereof was an hundred and thirty shekels, one silver bowl of seventy shekels, after the shekel of the sanctuary; both of them full of fine flour mingled with oil for a meat offering:
NUM|7|38|One golden spoon of ten shekels, full of incense:
NUM|7|39|One young bullock, one ram, one lamb of the first year, for a burnt offering:
NUM|7|40|One kid of the goats for a sin offering:
NUM|7|41|And for a sacrifice of peace offerings, two oxen, five rams, five he goats, five lambs of the first year: this was the offering of Shelumiel the son of Zurishaddai.
NUM|7|42|On the sixth day Eliasaph the son of Deuel, prince of the children of Gad, offered:
NUM|7|43|His offering was one silver charger of the weight of an hundred and thirty shekels, a silver bowl of seventy shekels, after the shekel of the sanctuary; both of them full of fine flour mingled with oil for a meat offering:
NUM|7|44|One golden spoon of ten shekels, full of incense:
NUM|7|45|One young bullock, one ram, one lamb of the first year, for a burnt offering:
NUM|7|46|One kid of the goats for a sin offering:
NUM|7|47|And for a sacrifice of peace offerings, two oxen, five rams, five he goats, five lambs of the first year: this was the offering of Eliasaph the son of Deuel.
NUM|7|48|On the seventh day Elishama the son of Ammihud, prince of the children of Ephraim, offered:
NUM|7|49|His offering was one silver charger, the weight whereof was an hundred and thirty shekels, one silver bowl of seventy shekels, after the shekel of the sanctuary; both of them full of fine flour mingled with oil for a meat offering:
NUM|7|50|One golden spoon of ten shekels, full of incense:
NUM|7|51|One young bullock, one ram, one lamb of the first year, for a burnt offering:
NUM|7|52|One kid of the goats for a sin offering:
NUM|7|53|And for a sacrifice of peace offerings, two oxen, five rams, five he goats, five lambs of the first year: this was the offering of Elishama the son of Ammihud.
NUM|7|54|On the eighth day offered Gamaliel the son of Pedahzur, prince of the children of Manasseh:
NUM|7|55|His offering was one silver charger of the weight of an hundred and thirty shekels, one silver bowl of seventy shekels, after the shekel of the sanctuary; both of them full of fine flour mingled with oil for a meat offering:
NUM|7|56|One golden spoon of ten shekels, full of incense:
NUM|7|57|One young bullock, one ram, one lamb of the first year, for a burnt offering:
NUM|7|58|One kid of the goats for a sin offering:
NUM|7|59|And for a sacrifice of peace offerings, two oxen, five rams, five he goats, five lambs of the first year: this was the offering of Gamaliel the son of Pedahzur.
NUM|7|60|On the ninth day Abidan the son of Gideoni, prince of the children of Benjamin, offered:
NUM|7|61|His offering was one silver charger, the weight whereof was an hundred and thirty shekels, one silver bowl of seventy shekels, after the shekel of the sanctuary; both of them full of fine flour mingled with oil for a meat offering:
NUM|7|62|One golden spoon of ten shekels, full of incense:
NUM|7|63|One young bullock, one ram, one lamb of the first year, for a burnt offering:
NUM|7|64|One kid of the goats for a sin offering:
NUM|7|65|And for a sacrifice of peace offerings, two oxen, five rams, five he goats, five lambs of the first year: this was the offering of Abidan the son of Gideoni.
NUM|7|66|On the tenth day Ahiezer the son of Ammishaddai, prince of the children of Dan, offered:
NUM|7|67|His offering was one silver charger, the weight whereof was an hundred and thirty shekels, one silver bowl of seventy shekels, after the shekel of the sanctuary; both of them full of fine flour mingled with oil for a meat offering:
NUM|7|68|One golden spoon of ten shekels, full of incense:
NUM|7|69|One young bullock, one ram, one lamb of the first year, for a burnt offering:
NUM|7|70|One kid of the goats for a sin offering:
NUM|7|71|And for a sacrifice of peace offerings, two oxen, five rams, five he goats, five lambs of the first year: this was the offering of Ahiezer the son of Ammishaddai.
NUM|7|72|On the eleventh day Pagiel the son of Ocran, prince of the children of Asher, offered:
NUM|7|73|His offering was one silver charger, the weight whereof was an hundred and thirty shekels, one silver bowl of seventy shekels, after the shekel of the sanctuary; both of them full of fine flour mingled with oil for a meat offering:
NUM|7|74|One golden spoon of ten shekels, full of incense:
NUM|7|75|One young bullock, one ram, one lamb of the first year, for a burnt offering:
NUM|7|76|One kid of the goats for a sin offering:
NUM|7|77|And for a sacrifice of peace offerings, two oxen, five rams, five he goats, five lambs of the first year: this was the offering of Pagiel the son of Ocran.
NUM|7|78|On the twelfth day Ahira the son of Enan, prince of the children of Naphtali, offered:
NUM|7|79|His offering was one silver charger, the weight whereof was an hundred and thirty shekels, one silver bowl of seventy shekels, after the shekel of the sanctuary; both of them full of fine flour mingled with oil for a meat offering:
NUM|7|80|One golden spoon of ten shekels, full of incense:
NUM|7|81|One young bullock, one ram, one lamb of the first year, for a burnt offering:
NUM|7|82|One kid of the goats for a sin offering:
NUM|7|83|And for a sacrifice of peace offerings, two oxen, five rams, five he goats, five lambs of the first year: this was the offering of Ahira the son of Enan.
NUM|7|84|This was the dedication of the altar, in the day when it was anointed, by the princes of Israel: twelve chargers of silver, twelve silver bowls, twelve spoons of gold:
NUM|7|85|Each charger of silver weighing an hundred and thirty shekels, each bowl seventy: all the silver vessels weighed two thousand and four hundred shekels, after the shekel of the sanctuary:
NUM|7|86|The golden spoons were twelve, full of incense, weighing ten shekels apiece, after the shekel of the sanctuary: all the gold of the spoons was an hundred and twenty shekels.
NUM|7|87|All the oxen for the burnt offering were twelve bullocks, the rams twelve, the lambs of the first year twelve, with their meat offering: and the kids of the goats for sin offering twelve.
NUM|7|88|And all the oxen for the sacrifice of the peace offerings were twenty and four bullocks, the rams sixty, the he goats sixty, the lambs of the first year sixty. This was the dedication of the altar, after that it was anointed.
NUM|7|89|And when Moses was gone into the tabernacle of the congregation to speak with him, then he heard the voice of one speaking unto him from off the mercy seat that was upon the ark of testimony, from between the two cherubim: and he spake unto him.
NUM|8|1|And the LORD spake unto Moses, saying,
NUM|8|2|Speak unto Aaron and say unto him, When thou lightest the lamps, the seven lamps shall give light over against the candlestick.
NUM|8|3|And Aaron did so; he lighted the lamps thereof over against the candlestick, as the LORD commanded Moses.
NUM|8|4|And this work of the candlestick was of beaten gold, unto the shaft thereof, unto the flowers thereof, was beaten work: according unto the pattern which the LORD had showed Moses, so he made the candlestick.
NUM|8|5|And the LORD spake unto Moses, saying,
NUM|8|6|Take the Levites from among the children of Israel, and cleanse them.
NUM|8|7|And thus shalt thou do unto them, to cleanse them: Sprinkle water of purifying upon them, and let them shave all their flesh, and let them wash their clothes, and so make themselves clean.
NUM|8|8|Then let them take a young bullock with his meat offering, even fine flour mingled with oil, and another young bullock shalt thou take for a sin offering.
NUM|8|9|And thou shalt bring the Levites before the tabernacle of the congregation: and thou shalt gather the whole assembly of the children of Israel together:
NUM|8|10|And thou shalt bring the Levites before the LORD: and the children of Israel shall put their hands upon the Levites:
NUM|8|11|And Aaron shall offer the Levites before the LORD for an offering of the children of Israel, that they may execute the service of the LORD.
NUM|8|12|And the Levites shall lay their hands upon the heads of the bullocks: and thou shalt offer the one for a sin offering, and the other for a burnt offering, unto the LORD, to make an atonement for the Levites.
NUM|8|13|And thou shalt set the Levites before Aaron, and before his sons, and offer them for an offering unto the LORD.
NUM|8|14|Thus shalt thou separate the Levites from among the children of Israel: and the Levites shall be mine.
NUM|8|15|And after that shall the Levites go in to do the service of the tabernacle of the congregation: and thou shalt cleanse them, and offer them for an offering.
NUM|8|16|For they are wholly given unto me from among the children of Israel; instead of such as open every womb, even instead of the firstborn of all the children of Israel, have I taken them unto me.
NUM|8|17|For all the firstborn of the children of Israel are mine, both man and beast: on the day that I smote every firstborn in the land of Egypt I sanctified them for myself.
NUM|8|18|And I have taken the Levites for all the firstborn of the children of Israel.
NUM|8|19|And I have given the Levites as a gift to Aaron and to his sons from among the children of Israel, to do the service of the children of Israel in the tabernacle of the congregation, and to make an atonement for the children of Israel: that there be no plague among the children of Israel, when the children of Israel come nigh unto the sanctuary.
NUM|8|20|And Moses, and Aaron, and all the congregation of the children of Israel, did to the Levites according unto all that the LORD commanded Moses concerning the Levites, so did the children of Israel unto them.
NUM|8|21|And the Levites were purified, and they washed their clothes; and Aaron offered them as an offering before the LORD; and Aaron made an atonement for them to cleanse them.
NUM|8|22|And after that went the Levites in to do their service in the tabernacle of the congregation before Aaron, and before his sons: as the LORD had commanded Moses concerning the Levites, so did they unto them.
NUM|8|23|And the LORD spake unto Moses, saying,
NUM|8|24|This is it that belongeth unto the Levites: from twenty and five years old and upward they shall go in to wait upon the service of the tabernacle of the congregation:
NUM|8|25|And from the age of fifty years they shall cease waiting upon the service thereof, and shall serve no more:
NUM|8|26|But shall minister with their brethren in the tabernacle of the congregation, to keep the charge, and shall do no service. Thus shalt thou do unto the Levites touching their charge.
NUM|9|1|And the LORD spake unto Moses in the wilderness of Sinai, in the first month of the second year after they were come out of the land of Egypt, saying,
NUM|9|2|Let the children of Israel also keep the passover at his appointed season.
NUM|9|3|In the fourteenth day of this month, at even, ye shall keep it in his appointed season: according to all the rites of it, and according to all the ceremonies thereof, shall ye keep it.
NUM|9|4|And Moses spake unto the children of Israel, that they should keep the passover.
NUM|9|5|And they kept the passover on the fourteenth day of the first month at even in the wilderness of Sinai: according to all that the LORD commanded Moses, so did the children of Israel.
NUM|9|6|And there were certain men, who were defiled by the dead body of a man, that they could not keep the passover on that day: and they came before Moses and before Aaron on that day:
NUM|9|7|And those men said unto him, We are defiled by the dead body of a man: wherefore are we kept back, that we may not offer an offering of the LORD in his appointed season among the children of Israel?
NUM|9|8|And Moses said unto them, Stand still, and I will hear what the LORD will command concerning you.
NUM|9|9|And the LORD spake unto Moses, saying,
NUM|9|10|Speak unto the children of Israel, saying, If any man of you or of your posterity shall be unclean by reason of a dead body, or be in a journey afar off, yet he shall keep the passover unto the LORD.
NUM|9|11|The fourteenth day of the second month at even they shall keep it, and eat it with unleavened bread and bitter herbs.
NUM|9|12|They shall leave none of it unto the morning, nor break any bone of it: according to all the ordinances of the passover they shall keep it.
NUM|9|13|But the man that is clean, and is not in a journey, and forbeareth to keep the passover, even the same soul shall be cut off from among his people: because he brought not the offering of the LORD in his appointed season, that man shall bear his sin.
NUM|9|14|And if a stranger shall sojourn among you, and will keep the passover unto the LORD; according to the ordinance of the passover, and according to the manner thereof, so shall he do: ye shall have one ordinance, both for the stranger, and for him that was born in the land.
NUM|9|15|And on the day that the tabernacle was reared up the cloud covered the tabernacle, namely, the tent of the testimony: and at even there was upon the tabernacle as it were the appearance of fire, until the morning.
NUM|9|16|So it was alway: the cloud covered it by day, and the appearance of fire by night.
NUM|9|17|And when the cloud was taken up from the tabernacle, then after that the children of Israel journeyed: and in the place where the cloud abode, there the children of Israel pitched their tents.
NUM|9|18|At the commandment of the LORD the children of Israel journeyed, and at the commandment of the LORD they pitched: as long as the cloud abode upon the tabernacle they rested in their tents.
NUM|9|19|And when the cloud tarried long upon the tabernacle many days, then the children of Israel kept the charge of the LORD, and journeyed not.
NUM|9|20|And so it was, when the cloud was a few days upon the tabernacle; according to the commandment of the LORD they abode in their tents, and according to the commandment of the LORD they journeyed.
NUM|9|21|And so it was, when the cloud abode from even unto the morning, and that the cloud was taken up in the morning, then they journeyed: whether it was by day or by night that the cloud was taken up, they journeyed.
NUM|9|22|Or whether it were two days, or a month, or a year, that the cloud tarried upon the tabernacle, remaining thereon, the children of Israel abode in their tents, and journeyed not: but when it was taken up, they journeyed.
NUM|9|23|At the commandment of the LORD they rested in the tents, and at the commandment of the LORD they journeyed: they kept the charge of the LORD, at the commandment of the LORD by the hand of Moses.
NUM|10|1|And the LORD spake unto Moses, saying,
NUM|10|2|Make thee two trumpets of silver; of a whole piece shalt thou make them: that thou mayest use them for the calling of the assembly, and for the journeying of the camps.
NUM|10|3|And when they shall blow with them, all the assembly shall assemble themselves to thee at the door of the tabernacle of the congregation.
NUM|10|4|And if they blow but with one trumpet, then the princes, which are heads of the thousands of Israel, shall gather themselves unto thee.
NUM|10|5|When ye blow an alarm, then the camps that lie on the east parts shall go forward.
NUM|10|6|When ye blow an alarm the second time, then the camps that lie on the south side shall take their journey: they shall blow an alarm for their journeys.
NUM|10|7|But when the congregation is to be gathered together, ye shall blow, but ye shall not sound an alarm.
NUM|10|8|And the sons of Aaron, the priests, shall blow with the trumpets; and they shall be to you for an ordinance for ever throughout your generations.
NUM|10|9|And if ye go to war in your land against the enemy that oppresseth you, then ye shall blow an alarm with the trumpets; and ye shall be remembered before the LORD your God, and ye shall be saved from your enemies.
NUM|10|10|Also in the day of your gladness, and in your solemn days, and in the beginnings of your months, ye shall blow with the trumpets over your burnt offerings, and over the sacrifices of your peace offerings; that they may be to you for a memorial before your God: I am the LORD your God.
NUM|10|11|And it came to pass on the twentieth day of the second month, in the second year, that the cloud was taken up from off the tabernacle of the testimony.
NUM|10|12|And the children of Israel took their journeys out of the wilderness of Sinai; and the cloud rested in the wilderness of Paran.
NUM|10|13|And they first took their journey according to the commandment of the LORD by the hand of Moses.
NUM|10|14|In the first place went the standard of the camp of the children of Judah according to their armies: and over his host was Nahshon the son of Amminadab.
NUM|10|15|And over the host of the tribe of the children of Issachar was Nethaneel the son of Zuar.
NUM|10|16|And over the host of the tribe of the children of Zebulun was Eliab the son of Helon.
NUM|10|17|And the tabernacle was taken down; and the sons of Gershon and the sons of Merari set forward, bearing the tabernacle.
NUM|10|18|And the standard of the camp of Reuben set forward according to their armies: and over his host was Elizur the son of Shedeur.
NUM|10|19|And over the host of the tribe of the children of Simeon was Shelumiel the son of Zurishaddai.
NUM|10|20|And over the host of the tribe of the children of Gad was Eliasaph the son of Deuel.
NUM|10|21|And the Kohathites set forward, bearing the sanctuary: and the other did set up the tabernacle against they came.
NUM|10|22|And the standard of the camp of the children of Ephraim set forward according to their armies: and over his host was Elishama the son of Ammihud.
NUM|10|23|And over the host of the tribe of the children of Manasseh was Gamaliel the son of Pedahzur.
NUM|10|24|And over the host of the tribe of the children of Benjamin was Abidan the son of Gideoni.
NUM|10|25|And the standard of the camp of the children of Dan set forward, which was the rearward of all the camps throughout their hosts: and over his host was Ahiezer the son of Ammishaddai.
NUM|10|26|And over the host of the tribe of the children of Asher was Pagiel the son of Ocran.
NUM|10|27|And over the host of the tribe of the children of Naphtali was Ahira the son of Enan.
NUM|10|28|Thus were the journeyings of the children of Israel according to their armies, when they set forward.
NUM|10|29|And Moses said unto Hobab, the son of Raguel the Midianite, Moses' father in law, We are journeying unto the place of which the LORD said, I will give it you: come thou with us, and we will do thee good: for the LORD hath spoken good concerning Israel.
NUM|10|30|And he said unto him, I will not go; but I will depart to mine own land, and to my kindred.
NUM|10|31|And he said, Leave us not, I pray thee; forasmuch as thou knowest how we are to encamp in the wilderness, and thou mayest be to us instead of eyes.
NUM|10|32|And it shall be, if thou go with us, yea, it shall be, that what goodness the LORD shall do unto us, the same will we do unto thee.
NUM|10|33|And they departed from the mount of the LORD three days' journey: and the ark of the covenant of the LORD went before them in the three days' journey, to search out a resting place for them.
NUM|10|34|And the cloud of the LORD was upon them by day, when they went out of the camp.
NUM|10|35|And it came to pass, when the ark set forward, that Moses said, Rise up, LORD, and let thine enemies be scattered; and let them that hate thee flee before thee.
NUM|10|36|And when it rested, he said, Return, O LORD, unto the many thousands of Israel.
NUM|11|1|And when the people complained, it displeased the LORD: and the LORD heard it; and his anger was kindled; and the fire of the LORD burnt among them, and consumed them that were in the uttermost parts of the camp.
NUM|11|2|And the people cried unto Moses; and when Moses prayed unto the LORD, the fire was quenched.
NUM|11|3|And he called the name of the place Taberah: because the fire of the LORD burnt among them.
NUM|11|4|And the mixed multitude that was among them fell a lusting: and the children of Israel also wept again, and said, Who shall give us flesh to eat?
NUM|11|5|We remember the fish, which we did eat in Egypt freely; the cucumbers, and the melons, and the leeks, and the onions, and the garlic:
NUM|11|6|But now our soul is dried away: there is nothing at all, beside this manna, before our eyes.
NUM|11|7|And the manna was as coriander seed, and the color thereof as the color of bdellium.
NUM|11|8|And the people went about, and gathered it, and ground it in mills, or beat it in a mortar, and baked it in pans, and made cakes of it: and the taste of it was as the taste of fresh oil.
NUM|11|9|And when the dew fell upon the camp in the night, the manna fell upon it.
NUM|11|10|Then Moses heard the people weep throughout their families, every man in the door of his tent: and the anger of the LORD was kindled greatly; Moses also was displeased.
NUM|11|11|And Moses said unto the LORD, Wherefore hast thou afflicted thy servant? and wherefore have I not found favor in thy sight, that thou layest the burden of all this people upon me?
NUM|11|12|Have I conceived all this people? have I begotten them, that thou shouldest say unto me, Carry them in thy bosom, as a nursing father beareth the sucking child, unto the land which thou swarest unto their fathers?
NUM|11|13|Whence should I have flesh to give unto all this people? for they weep unto me, saying, Give us flesh, that we may eat.
NUM|11|14|I am not able to bear all this people alone, because it is too heavy for me.
NUM|11|15|And if thou deal thus with me, kill me, I pray thee, out of hand, if I have found favor in thy sight; and let me not see my wretchedness.
NUM|11|16|And the LORD said unto Moses, Gather unto me seventy men of the elders of Israel, whom thou knowest to be the elders of the people, and officers over them; and bring them unto the tabernacle of the congregation, that they may stand there with thee.
NUM|11|17|And I will come down and talk with thee there: and I will take of the spirit which is upon thee, and will put it upon them; and they shall bear the burden of the people with thee, that thou bear it not thyself alone.
NUM|11|18|And say thou unto the people, Sanctify yourselves against to morrow, and ye shall eat flesh: for ye have wept in the ears of the LORD, saying, Who shall give us flesh to eat? for it was well with us in Egypt: therefore the LORD will give you flesh, and ye shall eat.
NUM|11|19|Ye shall not eat one day, nor two days, nor five days, neither ten days, nor twenty days;
NUM|11|20|But even a whole month, until it come out at your nostrils, and it be loathsome unto you: because that ye have despised the LORD which is among you, and have wept before him, saying, Why came we forth out of Egypt?
NUM|11|21|And Moses said, The people, among whom I am, are six hundred thousand footmen; and thou hast said, I will give them flesh, that they may eat a whole month.
NUM|11|22|Shall the flocks and the herds be slain for them, to suffice them? or shall all the fish of the sea be gathered together for them, to suffice them?
NUM|11|23|And the LORD said unto Moses, Is the LORD's hand waxed short? thou shalt see now whether my word shall come to pass unto thee or not.
NUM|11|24|And Moses went out, and told the people the words of the LORD, and gathered the seventy men of the elders of the people, and set them round about the tabernacle.
NUM|11|25|And the LORD came down in a cloud, and spake unto him, and took of the spirit that was upon him, and gave it unto the seventy elders: and it came to pass, that, when the spirit rested upon them, they prophesied, and did not cease.
NUM|11|26|But there remained two of the men in the camp, the name of the one was Eldad, and the name of the other Medad: and the spirit rested upon them; and they were of them that were written, but went not out unto the tabernacle: and they prophesied in the camp.
NUM|11|27|And there ran a young man, and told Moses, and said, Eldad and Medad do prophesy in the camp.
NUM|11|28|And Joshua the son of Nun, the servant of Moses, one of his young men, answered and said, My lord Moses, forbid them.
NUM|11|29|And Moses said unto him, Enviest thou for my sake? would God that all the LORD's people were prophets, and that the LORD would put his spirit upon them!
NUM|11|30|And Moses gat him into the camp, he and the elders of Israel.
NUM|11|31|And there went forth a wind from the LORD, and brought quails from the sea, and let them fall by the camp, as it were a day's journey on this side, and as it were a day's journey on the other side, round about the camp, and as it were two cubits high upon the face of the earth.
NUM|11|32|And the people stood up all that day, and all that night, and all the next day, and they gathered the quails: he that gathered least gathered ten homers: and they spread them all abroad for themselves round about the camp.
NUM|11|33|And while the flesh was yet between their teeth, ere it was chewed, the wrath of the LORD was kindled against the people, and the LORD smote the people with a very great plague.
NUM|11|34|And he called the name of that place Kibrothhattaavah: because there they buried the people that lusted.
NUM|11|35|And the people journeyed from Kibrothhattaavah unto Hazeroth; and abode at Hazeroth.
NUM|12|1|And Miriam and Aaron spake against Moses because of the Ethiopian woman whom he had married: for he had married an Ethiopian woman.
NUM|12|2|And they said, Hath the LORD indeed spoken only by Moses? hath he not spoken also by us? And the LORD heard it.
NUM|12|3|(Now the man Moses was very meek, above all the men which were upon the face of the earth.)
NUM|12|4|And the LORD spake suddenly unto Moses, and unto Aaron, and unto Miriam, Come out ye three unto the tabernacle of the congregation. And they three came out.
NUM|12|5|And the LORD came down in the pillar of the cloud, and stood in the door of the tabernacle, and called Aaron and Miriam: and they both came forth.
NUM|12|6|And he said, Hear now my words: If there be a prophet among you, I the LORD will make myself known unto him in a vision, and will speak unto him in a dream.
NUM|12|7|My servant Moses is not so, who is faithful in all mine house.
NUM|12|8|With him will I speak mouth to mouth, even apparently, and not in dark speeches; and the similitude of the LORD shall he behold: wherefore then were ye not afraid to speak against my servant Moses?
NUM|12|9|And the anger of the LORD was kindled against them; and he departed.
NUM|12|10|And the cloud departed from off the tabernacle; and, behold, Miriam became leprous, white as snow: and Aaron looked upon Miriam, and, behold, she was leprous.
NUM|12|11|And Aaron said unto Moses, Alas, my lord, I beseech thee, lay not the sin upon us, wherein we have done foolishly, and wherein we have sinned.
NUM|12|12|Let her not be as one dead, of whom the flesh is half consumed when he cometh out of his mother's womb.
NUM|12|13|And Moses cried unto the LORD, saying, Heal her now, O God, I beseech thee.
NUM|12|14|And the LORD said unto Moses, If her father had but spit in her face, should she not be ashamed seven days? let her be shut out from the camp seven days, and after that let her be received in again.
NUM|12|15|And Miriam was shut out from the camp seven days: and the people journeyed not till Miriam was brought in again.
NUM|12|16|And afterward the people removed from Hazeroth, and pitched in the wilderness of Paran.
NUM|13|1|And the LORD spake unto Moses, saying,
NUM|13|2|Send thou men, that they may search the land of Canaan, which I give unto the children of Israel: of every tribe of their fathers shall ye send a man, every one a ruler among them.
NUM|13|3|And Moses by the commandment of the LORD sent them from the wilderness of Paran: all those men were heads of the children of Israel.
NUM|13|4|And these were their names: of the tribe of Reuben, Shammua the son of Zaccur.
NUM|13|5|Of the tribe of Simeon, Shaphat the son of Hori.
NUM|13|6|Of the tribe of Judah, Caleb the son of Jephunneh.
NUM|13|7|Of the tribe of Issachar, Igal the son of Joseph.
NUM|13|8|Of the tribe of Ephraim, Oshea the son of Nun.
NUM|13|9|Of the tribe of Benjamin, Palti the son of Raphu.
NUM|13|10|Of the tribe of Zebulun, Gaddiel the son of Sodi.
NUM|13|11|Of the tribe of Joseph, namely, of the tribe of Manasseh, Gaddi the son of Susi.
NUM|13|12|Of the tribe of Dan, Ammiel the son of Gemalli.
NUM|13|13|Of the tribe of Asher, Sethur the son of Michael.
NUM|13|14|Of the tribe of Naphtali, Nahbi the son of Vophsi.
NUM|13|15|Of the tribe of Gad, Geuel the son of Machi.
NUM|13|16|These are the names of the men which Moses sent to spy out the land. And Moses called Oshea the son of Nun Jehoshua.
NUM|13|17|And Moses sent them to spy out the land of Canaan, and said unto them, Get you up this way southward, and go up into the mountain:
NUM|13|18|And see the land, what it is, and the people that dwelleth therein, whether they be strong or weak, few or many;
NUM|13|19|And what the land is that they dwell in, whether it be good or bad; and what cities they be that they dwell in, whether in tents, or in strong holds;
NUM|13|20|And what the land is, whether it be fat or lean, whether there be wood therein, or not. And be ye of good courage, and bring of the fruit of the land. Now the time was the time of the first ripe grapes.
NUM|13|21|So they went up, and searched the land from the wilderness of Zin unto Rehob, as men come to Hamath.
NUM|13|22|And they ascended by the south, and came unto Hebron; where Ahiman, Sheshai, and Talmai, the children of Anak, were. (Now Hebron was built seven years before Zoan in Egypt.)
NUM|13|23|And they came unto the brook of Eshcol, and cut down from thence a branch with one cluster of grapes, and they bare it between two upon a staff; and they brought of the pomegranates, and of the figs.
NUM|13|24|The place was called the brook Eshcol, because of the cluster of grapes which the children of Israel cut down from thence.
NUM|13|25|And they returned from searching of the land after forty days.
NUM|13|26|And they went and came to Moses, and to Aaron, and to all the congregation of the children of Israel, unto the wilderness of Paran, to Kadesh; and brought back word unto them, and unto all the congregation, and showed them the fruit of the land.
NUM|13|27|And they told him, and said, We came unto the land whither thou sentest us, and surely it floweth with milk and honey; and this is the fruit of it.
NUM|13|28|Nevertheless the people be strong that dwell in the land, and the cities are walled, and very great: and moreover we saw the children of Anak there.
NUM|13|29|The Amalekites dwell in the land of the south: and the Hittites, and the Jebusites, and the Amorites, dwell in the mountains: and the Canaanites dwell by the sea, and by the coast of Jordan.
NUM|13|30|And Caleb stilled the people before Moses, and said, Let us go up at once, and possess it; for we are well able to overcome it.
NUM|13|31|But the men that went up with him said, We be not able to go up against the people; for they are stronger than we.
NUM|13|32|And they brought up an evil report of the land which they had searched unto the children of Israel, saying, The land, through which we have gone to search it, is a land that eateth up the inhabitants thereof; and all the people that we saw in it are men of a great stature.
NUM|13|33|And there we saw the giants, the sons of Anak, which come of the giants: and we were in our own sight as grasshoppers, and so we were in their sight.
NUM|14|1|And all the congregation lifted up their voice, and cried; and the people wept that night.
NUM|14|2|And all the children of Israel murmured against Moses and against Aaron: and the whole congregation said unto them, Would God that we had died in the land of Egypt! or would God we had died in this wilderness!
NUM|14|3|And wherefore hath the LORD brought us unto this land, to fall by the sword, that our wives and our children should be a prey? were it not better for us to return into Egypt?
NUM|14|4|And they said one to another, Let us make a captain, and let us return into Egypt.
NUM|14|5|Then Moses and Aaron fell on their faces before all the assembly of the congregation of the children of Israel.
NUM|14|6|And Joshua the son of Nun, and Caleb the son of Jephunneh, which were of them that searched the land, rent their clothes:
NUM|14|7|And they spake unto all the company of the children of Israel, saying, The land, which we passed through to search it, is an exceeding good land.
NUM|14|8|If the LORD delight in us, then he will bring us into this land, and give it us; a land which floweth with milk and honey.
NUM|14|9|Only rebel not ye against the LORD, neither fear ye the people of the land; for they are bread for us: their defense is departed from them, and the LORD is with us: fear them not.
NUM|14|10|But all the congregation bade stone them with stones. And the glory of the LORD appeared in the tabernacle of the congregation before all the children of Israel.
NUM|14|11|And the LORD said unto Moses, How long will this people provoke me? and how long will it be ere they believe me, for all the signs which I have showed among them?
NUM|14|12|I will smite them with the pestilence, and disinherit them, and will make of thee a greater nation and mightier than they.
NUM|14|13|And Moses said unto the LORD, Then the Egyptians shall hear it, (for thou broughtest up this people in thy might from among them;)
NUM|14|14|And they will tell it to the inhabitants of this land: for they have heard that thou LORD art among this people, that thou LORD art seen face to face, and that thy cloud standeth over them, and that thou goest before them, by day time in a pillar of a cloud, and in a pillar of fire by night.
NUM|14|15|Now if thou shalt kill all this people as one man, then the nations which have heard the fame of thee will speak, saying,
NUM|14|16|Because the LORD was not able to bring this people into the land which he sware unto them, therefore he hath slain them in the wilderness.
NUM|14|17|And now, I beseech thee, let the power of my Lord be great, according as thou hast spoken, saying,
NUM|14|18|The LORD is long-suffering, and of great mercy, forgiving iniquity and transgression, and by no means clearing the guilty, visiting the iniquity of the fathers upon the children unto the third and fourth generation.
NUM|14|19|Pardon, I beseech thee, the iniquity of this people according unto the greatness of thy mercy, and as thou hast forgiven this people, from Egypt even until now.
NUM|14|20|And the LORD said, I have pardoned according to thy word:
NUM|14|21|But as truly as I live, all the earth shall be filled with the glory of the LORD.
NUM|14|22|Because all those men which have seen my glory, and my miracles, which I did in Egypt and in the wilderness, and have tempted me now these ten times, and have not hearkened to my voice;
NUM|14|23|Surely they shall not see the land which I sware unto their fathers, neither shall any of them that provoked me see it:
NUM|14|24|But my servant Caleb, because he had another spirit with him, and hath followed me fully, him will I bring into the land whereinto he went; and his seed shall possess it.
NUM|14|25|(Now the Amalekites and the Canaanites dwelt in the valley.) Tomorrow turn you, and get you into the wilderness by the way of the Red sea.
NUM|14|26|And the LORD spake unto Moses and unto Aaron, saying,
NUM|14|27|How long shall I bear with this evil congregation, which murmur against me? I have heard the murmurings of the children of Israel, which they murmur against me.
NUM|14|28|Say unto them, As truly as I live, saith the LORD, as ye have spoken in mine ears, so will I do to you:
NUM|14|29|Your carcasses shall fall in this wilderness; and all that were numbered of you, according to your whole number, from twenty years old and upward which have murmured against me.
NUM|14|30|Doubtless ye shall not come into the land, concerning which I sware to make you dwell therein, save Caleb the son of Jephunneh, and Joshua the son of Nun.
NUM|14|31|But your little ones, which ye said should be a prey, them will I bring in, and they shall know the land which ye have despised.
NUM|14|32|But as for you, your carcasses, they shall fall in this wilderness.
NUM|14|33|And your children shall wander in the wilderness forty years, and bear your whoredoms, until your carcasses be wasted in the wilderness.
NUM|14|34|After the number of the days in which ye searched the land, even forty days, each day for a year, shall ye bear your iniquities, even forty years, and ye shall know my breach of promise.
NUM|14|35|I the LORD have said, I will surely do it unto all this evil congregation, that are gathered together against me: in this wilderness they shall be consumed, and there they shall die.
NUM|14|36|And the men, which Moses sent to search the land, who returned, and made all the congregation to murmur against him, by bringing up a slander upon the land,
NUM|14|37|Even those men that did bring up the evil report upon the land, died by the plague before the LORD.
NUM|14|38|But Joshua the son of Nun, and Caleb the son of Jephunneh, which were of the men that went to search the land, lived still.
NUM|14|39|And Moses told these sayings unto all the children of Israel: and the people mourned greatly.
NUM|14|40|And they rose up early in the morning, and gat them up into the top of the mountain, saying, Lo, we be here, and will go up unto the place which the LORD hath promised: for we have sinned.
NUM|14|41|And Moses said, Wherefore now do ye transgress the commandment of the LORD? but it shall not prosper.
NUM|14|42|Go not up, for the LORD is not among you; that ye be not smitten before your enemies.
NUM|14|43|For the Amalekites and the Canaanites are there before you, and ye shall fall by the sword: because ye are turned away from the LORD, therefore the LORD will not be with you.
NUM|14|44|But they presumed to go up unto the hill top: nevertheless the ark of the covenant of the LORD, and Moses, departed not out of the camp.
NUM|14|45|Then the Amalekites came down, and the Canaanites which dwelt in that hill, and smote them, and discomfited them, even unto Hormah.
NUM|15|1|And the LORD spake unto Moses, saying,
NUM|15|2|Speak unto the children of Israel, and say unto them, When ye be come into the land of your habitations, which I give unto you,
NUM|15|3|And will make an offering by fire unto the LORD, a burnt offering, or a sacrifice in performing a vow, or in a freewill offering, or in your solemn feasts, to make a sweet savor unto the LORD, of the herd or of the flock:
NUM|15|4|Then shall he that offereth his offering unto the LORD bring a meat offering of a tenth deal of flour mingled with the fourth part of an hin of oil.
NUM|15|5|And the fourth part of an hin of wine for a drink offering shalt thou prepare with the burnt offering or sacrifice, for one lamb.
NUM|15|6|Or for a ram, thou shalt prepare for a meat offering two tenth deals of flour mingled with the third part of an hin of oil.
NUM|15|7|And for a drink offering thou shalt offer the third part of an hin of wine, for a sweet savor unto the LORD.
NUM|15|8|And when thou preparest a bullock for a burnt offering, or for a sacrifice in performing a vow, or peace offerings unto the LORD:
NUM|15|9|Then shall he bring with a bullock a meat offering of three tenth deals of flour mingled with half an hin of oil.
NUM|15|10|And thou shalt bring for a drink offering half an hin of wine, for an offering made by fire, of a sweet savor unto the LORD.
NUM|15|11|Thus shall it be done for one bullock, or for one ram, or for a lamb, or a kid.
NUM|15|12|According to the number that ye shall prepare, so shall ye do to every one according to their number.
NUM|15|13|All that are born of the country shall do these things after this manner, in offering an offering made by fire, of a sweet savor unto the LORD.
NUM|15|14|And if a stranger sojourn with you, or whosoever be among you in your generations, and will offer an offering made by fire, of a sweet savor unto the LORD; as ye do, so he shall do.
NUM|15|15|One ordinance shall be both for you of the congregation, and also for the stranger that sojourneth with you, an ordinance for ever in your generations: as ye are, so shall the stranger be before the LORD.
NUM|15|16|One law and one manner shall be for you, and for the stranger that sojourneth with you.
NUM|15|17|And the LORD spake unto Moses, saying,
NUM|15|18|Speak unto the children of Israel, and say unto them, When ye come into the land whither I bring you,
NUM|15|19|Then it shall be, that, when ye eat of the bread of the land, ye shall offer up an heave offering unto the LORD.
NUM|15|20|Ye shall offer up a cake of the first of your dough for an heave offering: as ye do the heave offering of the threshingfloor, so shall ye heave it.
NUM|15|21|Of the first of your dough ye shall give unto the LORD an heave offering in your generations.
NUM|15|22|And if ye have erred, and not observed all these commandments, which the LORD hath spoken unto Moses,
NUM|15|23|Even all that the LORD hath commanded you by the hand of Moses, from the day that the LORD commanded Moses, and henceforward among your generations;
NUM|15|24|Then it shall be, if ought be committed by ignorance without the knowledge of the congregation, that all the congregation shall offer one young bullock for a burnt offering, for a sweet savor unto the LORD, with his meat offering, and his drink offering, according to the manner, and one kid of the goats for a sin offering.
NUM|15|25|And the priest shall make an atonement for all the congregation of the children of Israel, and it shall be forgiven them; for it is ignorance: and they shall bring their offering, a sacrifice made by fire unto the LORD, and their sin offering before the LORD, for their ignorance:
NUM|15|26|And it shall be forgiven all the congregation of the children of Israel, and the stranger that sojourneth among them; seeing all the people were in ignorance.
NUM|15|27|And if any soul sin through ignorance, then he shall bring a she goat of the first year for a sin offering.
NUM|15|28|And the priest shall make an atonement for the soul that sinneth ignorantly, when he sinneth by ignorance before the LORD, to make an atonement for him; and it shall be forgiven him.
NUM|15|29|Ye shall have one law for him that sinneth through ignorance, both for him that is born among the children of Israel, and for the stranger that sojourneth among them.
NUM|15|30|But the soul that doeth ought presumptuously, whether he be born in the land, or a stranger, the same reproacheth the LORD; and that soul shall be cut off from among his people.
NUM|15|31|Because he hath despised the word of the LORD, and hath broken his commandment, that soul shall utterly be cut off; his iniquity shall be upon him.
NUM|15|32|And while the children of Israel were in the wilderness, they found a man that gathered sticks upon the sabbath day.
NUM|15|33|And they that found him gathering sticks brought him unto Moses and Aaron, and unto all the congregation.
NUM|15|34|And they put him in ward, because it was not declared what should be done to him.
NUM|15|35|And the LORD said unto Moses, The man shall be surely put to death: all the congregation shall stone him with stones without the camp.
NUM|15|36|And all the congregation brought him without the camp, and stoned him with stones, and he died; as the LORD commanded Moses.
NUM|15|37|And the LORD spake unto Moses, saying,
NUM|15|38|Speak unto the children of Israel, and bid them that they make them fringes in the borders of their garments throughout their generations, and that they put upon the fringe of the borders a ribband of blue:
NUM|15|39|And it shall be unto you for a fringe, that ye may look upon it, and remember all the commandments of the LORD, and do them; and that ye seek not after your own heart and your own eyes, after which ye use to go a whoring:
NUM|15|40|That ye may remember, and do all my commandments, and be holy unto your God.
NUM|15|41|I am the LORD your God, which brought you out of the land of Egypt, to be your God: I am the LORD your God.
NUM|16|1|Now Korah, the son of Izhar, the son of Kohath, the son of Levi, and Dathan and Abiram, the sons of Eliab, and On, the son of Peleth, sons of Reuben, took men:
NUM|16|2|And they rose up before Moses, with certain of the children of Israel, two hundred and fifty princes of the assembly, famous in the congregation, men of renown:
NUM|16|3|And they gathered themselves together against Moses and against Aaron, and said unto them, Ye take too much upon you, seeing all the congregation are holy, every one of them, and the LORD is among them: wherefore then lift ye up yourselves above the congregation of the LORD?
NUM|16|4|And when Moses heard it, he fell upon his face:
NUM|16|5|And he spake unto Korah and unto all his company, saying, Even to morrow the LORD will show who are his, and who is holy; and will cause him to come near unto him: even him whom he hath chosen will he cause to come near unto him.
NUM|16|6|This do; Take you censers, Korah, and all his company;
NUM|16|7|And put fire therein, and put incense in them before the LORD to morrow: and it shall be that the man whom the LORD doth choose, he shall be holy: ye take too much upon you, ye sons of Levi.
NUM|16|8|And Moses said unto Korah, Hear, I pray you, ye sons of Levi:
NUM|16|9|Seemeth it but a small thing unto you, that the God of Israel hath separated you from the congregation of Israel, to bring you near to himself to do the service of the tabernacle of the LORD, and to stand before the congregation to minister unto them?
NUM|16|10|And he hath brought thee near to him, and all thy brethren the sons of Levi with thee: and seek ye the priesthood also?
NUM|16|11|For which cause both thou and all thy company are gathered together against the LORD: and what is Aaron, that ye murmur against him?
NUM|16|12|And Moses sent to call Dathan and Abiram, the sons of Eliab: which said, We will not come up:
NUM|16|13|Is it a small thing that thou hast brought us up out of a land that floweth with milk and honey, to kill us in the wilderness, except thou make thyself altogether a prince over us?
NUM|16|14|Moreover thou hast not brought us into a land that floweth with milk and honey, or given us inheritance of fields and vineyards: wilt thou put out the eyes of these men? we will not come up.
NUM|16|15|And Moses was very wroth, and said unto the LORD, Respect not thou their offering: I have not taken one ass from them, neither have I hurt one of them.
NUM|16|16|And Moses said unto Korah, Be thou and all thy company before the LORD, thou, and they, and Aaron, to morrow:
NUM|16|17|And take every man his censer, and put incense in them, and bring ye before the LORD every man his censer, two hundred and fifty censers; thou also, and Aaron, each of you his censer.
NUM|16|18|And they took every man his censer, and put fire in them, and laid incense thereon, and stood in the door of the tabernacle of the congregation with Moses and Aaron.
NUM|16|19|And Korah gathered all the congregation against them unto the door of the tabernacle of the congregation: and the glory of the LORD appeared unto all the congregation.
NUM|16|20|And the LORD spake unto Moses and unto Aaron, saying,
NUM|16|21|Separate yourselves from among this congregation, that I may consume them in a moment.
NUM|16|22|And they fell upon their faces, and said, O God, the God of the spirits of all flesh, shall one man sin, and wilt thou be wroth with all the congregation?
NUM|16|23|And the LORD spake unto Moses, saying,
NUM|16|24|Speak unto the congregation, saying, Get you up from about the tabernacle of Korah, Dathan, and Abiram.
NUM|16|25|And Moses rose up and went unto Dathan and Abiram; and the elders of Israel followed him.
NUM|16|26|And he spake unto the congregation, saying, Depart, I pray you, from the tents of these wicked men, and touch nothing of theirs, lest ye be consumed in all their sins.
NUM|16|27|So they gat up from the tabernacle of Korah, Dathan, and Abiram, on every side: and Dathan and Abiram came out, and stood in the door of their tents, and their wives, and their sons, and their little children.
NUM|16|28|And Moses said, Hereby ye shall know that the LORD hath sent me to do all these works; for I have not done them of mine own mind.
NUM|16|29|If these men die the common death of all men, or if they be visited after the visitation of all men; then the LORD hath not sent me.
NUM|16|30|But if the LORD make a new thing, and the earth open her mouth, and swallow them up, with all that appertain unto them, and they go down quick into the pit; then ye shall understand that these men have provoked the LORD.
NUM|16|31|And it came to pass, as he had made an end of speaking all these words, that the ground clave asunder that was under them:
NUM|16|32|And the earth opened her mouth, and swallowed them up, and their houses, and all the men that appertained unto Korah, and all their goods.
NUM|16|33|They, and all that appertained to them, went down alive into the pit, and the earth closed upon them: and they perished from among the congregation.
NUM|16|34|And all Israel that were round about them fled at the cry of them: for they said, Lest the earth swallow us up also.
NUM|16|35|And there came out a fire from the LORD, and consumed the two hundred and fifty men that offered incense.
NUM|16|36|And the LORD spake unto Moses, saying,
NUM|16|37|Speak unto Eleazar the son of Aaron the priest, that he take up the censers out of the burning, and scatter thou the fire yonder; for they are hallowed.
NUM|16|38|The censers of these sinners against their own souls, let them make them broad plates for a covering of the altar: for they offered them before the LORD, therefore they are hallowed: and they shall be a sign unto the children of Israel.
NUM|16|39|And Eleazar the priest took the brazen censers, wherewith they that were burnt had offered; and they were made broad plates for a covering of the altar:
NUM|16|40|To be a memorial unto the children of Israel, that no stranger, which is not of the seed of Aaron, come near to offer incense before the LORD; that he be not as Korah, and as his company: as the LORD said to him by the hand of Moses.
NUM|16|41|But on the morrow all the congregation of the children of Israel murmured against Moses and against Aaron, saying, Ye have killed the people of the LORD.
NUM|16|42|And it came to pass, when the congregation was gathered against Moses and against Aaron, that they looked toward the tabernacle of the congregation: and, behold, the cloud covered it, and the glory of the LORD appeared.
NUM|16|43|And Moses and Aaron came before the tabernacle of the congregation.
NUM|16|44|And the LORD spake unto Moses, saying,
NUM|16|45|Get you up from among this congregation, that I may consume them as in a moment. And they fell upon their faces.
NUM|16|46|And Moses said unto Aaron, Take a censer, and put fire therein from off the altar, and put on incense, and go quickly unto the congregation, and make an atonement for them: for there is wrath gone out from the LORD; the plague is begun.
NUM|16|47|And Aaron took as Moses commanded, and ran into the midst of the congregation; and, behold, the plague was begun among the people: and he put on incense, and made an atonement for the people.
NUM|16|48|And he stood between the dead and the living; and the plague was stayed.
NUM|16|49|Now they that died in the plague were fourteen thousand and seven hundred, beside them that died about the matter of Korah.
NUM|16|50|And Aaron returned unto Moses unto the door of the tabernacle of the congregation: and the plague was stayed.
NUM|17|1|And the LORD spake unto Moses, saying,
NUM|17|2|Speak unto the children of Israel, and take of every one of them a rod according to the house of their fathers, of all their princes according to the house of their fathers twelve rods: write thou every man's name upon his rod.
NUM|17|3|And thou shalt write Aaron's name upon the rod of Levi: for one rod shall be for the head of the house of their fathers.
NUM|17|4|And thou shalt lay them up in the tabernacle of the congregation before the testimony, where I will meet with you.
NUM|17|5|And it shall come to pass, that the man's rod, whom I shall choose, shall blossom: and I will make to cease from me the murmurings of the children of Israel, whereby they murmur against you.
NUM|17|6|And Moses spake unto the children of Israel, and every one of their princes gave him a rod apiece, for each prince one, according to their fathers' houses, even twelve rods: and the rod of Aaron was among their rods.
NUM|17|7|And Moses laid up the rods before the LORD in the tabernacle of witness.
NUM|17|8|And it came to pass, that on the morrow Moses went into the tabernacle of witness; and, behold, the rod of Aaron for the house of Levi was budded, and brought forth buds, and bloomed blossoms, and yielded almonds.
NUM|17|9|And Moses brought out all the rods from before the LORD unto all the children of Israel: and they looked, and took every man his rod.
NUM|17|10|And the LORD said unto Moses, Bring Aaron's rod again before the testimony, to be kept for a token against the rebels; and thou shalt quite take away their murmurings from me, that they die not.
NUM|17|11|And Moses did so: as the LORD commanded him, so did he.
NUM|17|12|And the children of Israel spake unto Moses, saying, Behold, we die, we perish, we all perish.
NUM|17|13|Whosoever cometh any thing near unto the tabernacle of the LORD shall die: shall we be consumed with dying?
NUM|18|1|And the LORD said unto Aaron, Thou and thy sons and thy father's house with thee shall bear the iniquity of the sanctuary: and thou and thy sons with thee shall bear the iniquity of your priesthood.
NUM|18|2|And thy brethren also of the tribe of Levi, the tribe of thy father, bring thou with thee, that they may be joined unto thee, and minister unto thee: but thou and thy sons with thee shall minister before the tabernacle of witness.
NUM|18|3|And they shall keep thy charge, and the charge of all the tabernacle: only they shall not come nigh the vessels of the sanctuary and the altar, that neither they, nor ye also, die.
NUM|18|4|And they shall be joined unto thee, and keep the charge of the tabernacle of the congregation, for all the service of the tabernacle: and a stranger shall not come nigh unto you.
NUM|18|5|And ye shall keep the charge of the sanctuary, and the charge of the altar: that there be no wrath any more upon the children of Israel.
NUM|18|6|And I, behold, I have taken your brethren the Levites from among the children of Israel: to you they are given as a gift for the LORD, to do the service of the tabernacle of the congregation.
NUM|18|7|Therefore thou and thy sons with thee shall keep your priest's office for everything of the altar, and within the vail; and ye shall serve: I have given your priest's office unto you as a service of gift: and the stranger that cometh nigh shall be put to death.
NUM|18|8|And the LORD spake unto Aaron, Behold, I also have given thee the charge of mine heave offerings of all the hallowed things of the children of Israel; unto thee have I given them by reason of the anointing, and to thy sons, by an ordinance for ever.
NUM|18|9|This shall be thine of the most holy things, reserved from the fire: every oblation of theirs, every meat offering of theirs, and every sin offering of theirs, and every trespass offering of theirs which they shall render unto me, shall be most holy for thee and for thy sons.
NUM|18|10|In the most holy place shalt thou eat it; every male shall eat it: it shall be holy unto thee.
NUM|18|11|And this is thine; the heave offering of their gift, with all the wave offerings of the children of Israel: I have given them unto thee, and to thy sons and to thy daughters with thee, by a statute for ever: every one that is clean in thy house shall eat of it.
NUM|18|12|All the best of the oil, and all the best of the wine, and of the wheat, the firstfruits of them which they shall offer unto the LORD, them have I given thee.
NUM|18|13|And whatsoever is first ripe in the land, which they shall bring unto the LORD, shall be thine; every one that is clean in thine house shall eat of it.
NUM|18|14|Every thing devoted in Israel shall be thine.
NUM|18|15|Every thing that openeth the matrix in all flesh, which they bring unto the LORD, whether it be of men or beasts, shall be thine: nevertheless the firstborn of man shalt thou surely redeem, and the firstling of unclean beasts shalt thou redeem.
NUM|18|16|And those that are to be redeemed from a month old shalt thou redeem, according to thine estimation, for the money of five shekels, after the shekel of the sanctuary, which is twenty gerahs.
NUM|18|17|But the firstling of a cow, or the firstling of a sheep, or the firstling of a goat, thou shalt not redeem; they are holy: thou shalt sprinkle their blood upon the altar, and shalt burn their fat for an offering made by fire, for a sweet savor unto the LORD.
NUM|18|18|And the flesh of them shall be thine, as the wave breast and as the right shoulder are thine.
NUM|18|19|All the heave offerings of the holy things, which the children of Israel offer unto the LORD, have I given thee, and thy sons and thy daughters with thee, by a statute for ever: it is a covenant of salt for ever before the LORD unto thee and to thy seed with thee.
NUM|18|20|And the LORD spake unto Aaron, Thou shalt have no inheritance in their land, neither shalt thou have any part among them: I am thy part and thine inheritance among the children of Israel.
NUM|18|21|And, behold, I have given the children of Levi all the tenth in Israel for an inheritance, for their service which they serve, even the service of the tabernacle of the congregation.
NUM|18|22|Neither must the children of Israel henceforth come nigh the tabernacle of the congregation, lest they bear sin, and die.
NUM|18|23|But the Levites shall do the service of the tabernacle of the congregation, and they shall bear their iniquity: it shall be a statute for ever throughout your generations, that among the children of Israel they have no inheritance.
NUM|18|24|But the tithes of the children of Israel, which they offer as an heave offering unto the LORD, I have given to the Levites to inherit: therefore I have said unto them, Among the children of Israel they shall have no inheritance.
NUM|18|25|And the LORD spake unto Moses, saying,
NUM|18|26|Thus speak unto the Levites, and say unto them, When ye take of the children of Israel the tithes which I have given you from them for your inheritance, then ye shall offer up an heave offering of it for the LORD, even a tenth part of the tithe.
NUM|18|27|And this your heave offering shall be reckoned unto you, as though it were the corn of the threshingfloor, and as the fulness of the winepress.
NUM|18|28|Thus ye also shall offer an heave offering unto the LORD of all your tithes, which ye receive of the children of Israel; and ye shall give thereof the LORD's heave offering to Aaron the priest.
NUM|18|29|Out of all your gifts ye shall offer every heave offering of the LORD, of all the best thereof, even the hallowed part thereof out of it.
NUM|18|30|Therefore thou shalt say unto them, When ye have heaved the best thereof from it, then it shall be counted unto the Levites as the increase of the threshingfloor, and as the increase of the winepress.
NUM|18|31|And ye shall eat it in every place, ye and your households: for it is your reward for your service in the tabernacle of the congregation.
NUM|18|32|And ye shall bear no sin by reason of it, when ye have heaved from it the best of it: neither shall ye pollute the holy things of the children of Israel, lest ye die.
NUM|19|1|And the LORD spake unto Moses and unto Aaron, saying,
NUM|19|2|This is the ordinance of the law which the LORD hath commanded, saying, Speak unto the children of Israel, that they bring thee a red heifer without spot, wherein is no blemish, and upon which never came yoke:
NUM|19|3|And ye shall give her unto Eleazar the priest, that he may bring her forth without the camp, and one shall slay her before his face:
NUM|19|4|And Eleazar the priest shall take of her blood with his finger, and sprinkle of her blood directly before the tabernacle of the congregation seven times:
NUM|19|5|And one shall burn the heifer in his sight; her skin, and her flesh, and her blood, with her dung, shall he burn:
NUM|19|6|And the priest shall take cedar wood, and hyssop, and scarlet, and cast it into the midst of the burning of the heifer.
NUM|19|7|Then the priest shall wash his clothes, and he shall bathe his flesh in water, and afterward he shall come into the camp, and the priest shall be unclean until the even.
NUM|19|8|And he that burneth her shall wash his clothes in water, and bathe his flesh in water, and shall be unclean until the even.
NUM|19|9|And a man that is clean shall gather up the ashes of the heifer, and lay them up without the camp in a clean place, and it shall be kept for the congregation of the children of Israel for a water of separation: it is a purification for sin.
NUM|19|10|And he that gathereth the ashes of the heifer shall wash his clothes, and be unclean until the even: and it shall be unto the children of Israel, and unto the stranger that sojourneth among them, for a statute for ever.
NUM|19|11|He that toucheth the dead body of any man shall be unclean seven days.
NUM|19|12|He shall purify himself with it on the third day, and on the seventh day he shall be clean: but if he purify not himself the third day, then the seventh day he shall not be clean.
NUM|19|13|Whosoever toucheth the dead body of any man that is dead, and purifieth not himself, defileth the tabernacle of the LORD; and that soul shall be cut off from Israel: because the water of separation was not sprinkled upon him, he shall be unclean; his uncleanness is yet upon him.
NUM|19|14|This is the law, when a man dieth in a tent: all that come into the tent, and all that is in the tent, shall be unclean seven days.
NUM|19|15|And every open vessel, which hath no covering bound upon it, is unclean.
NUM|19|16|And whosoever toucheth one that is slain with a sword in the open fields, or a dead body, or a bone of a man, or a grave, shall be unclean seven days.
NUM|19|17|And for an unclean person they shall take of the ashes of the burnt heifer of purification for sin, and running water shall be put thereto in a vessel:
NUM|19|18|And a clean person shall take hyssop, and dip it in the water, and sprinkle it upon the tent, and upon all the vessels, and upon the persons that were there, and upon him that touched a bone, or one slain, or one dead, or a grave:
NUM|19|19|And the clean person shall sprinkle upon the unclean on the third day, and on the seventh day: and on the seventh day he shall purify himself, and wash his clothes, and bathe himself in water, and shall be clean at even.
NUM|19|20|But the man that shall be unclean, and shall not purify himself, that soul shall be cut off from among the congregation, because he hath defiled the sanctuary of the LORD: the water of separation hath not been sprinkled upon him; he is unclean.
NUM|19|21|And it shall be a perpetual statute unto them, that he that sprinkleth the water of separation shall wash his clothes; and he that toucheth the water of separation shall be unclean until even.
NUM|19|22|And whatsoever the unclean person toucheth shall be unclean; and the soul that toucheth it shall be unclean until even.
NUM|20|1|Then came the children of Israel, even the whole congregation, into the desert of Zin in the first month: and the people abode in Kadesh; and Miriam died there, and was buried there.
NUM|20|2|And there was no water for the congregation: and they gathered themselves together against Moses and against Aaron.
NUM|20|3|And the people chode with Moses, and spake, saying, Would God that we had died when our brethren died before the LORD!
NUM|20|4|And why have ye brought up the congregation of the LORD into this wilderness, that we and our cattle should die there?
NUM|20|5|And wherefore have ye made us to come up out of Egypt, to bring us in unto this evil place? it is no place of seed, or of figs, or of vines, or of pomegranates; neither is there any water to drink.
NUM|20|6|And Moses and Aaron went from the presence of the assembly unto the door of the tabernacle of the congregation, and they fell upon their faces: and the glory of the LORD appeared unto them.
NUM|20|7|And the LORD spake unto Moses, saying,
NUM|20|8|Take the rod, and gather thou the assembly together, thou, and Aaron thy brother, and speak ye unto the rock before their eyes; and it shall give forth his water, and thou shalt bring forth to them water out of the rock: so thou shalt give the congregation and their beasts drink.
NUM|20|9|And Moses took the rod from before the LORD, as he commanded him.
NUM|20|10|And Moses and Aaron gathered the congregation together before the rock, and he said unto them, Hear now, ye rebels; must we fetch you water out of this rock?
NUM|20|11|And Moses lifted up his hand, and with his rod he smote the rock twice: and the water came out abundantly, and the congregation drank, and their beasts also.
NUM|20|12|And the LORD spake unto Moses and Aaron, Because ye believed me not, to sanctify me in the eyes of the children of Israel, therefore ye shall not bring this congregation into the land which I have given them.
NUM|20|13|This is the water of Meribah; because the children of Israel strove with the LORD, and he was sanctified in them.
NUM|20|14|And Moses sent messengers from Kadesh unto the king of Edom, Thus saith thy brother Israel, Thou knowest all the travail that hath befallen us:
NUM|20|15|How our fathers went down into Egypt, and we have dwelt in Egypt a long time; and the Egyptians vexed us, and our fathers:
NUM|20|16|And when we cried unto the LORD, he heard our voice, and sent an angel, and hath brought us forth out of Egypt: and, behold, we are in Kadesh, a city in the uttermost of thy border:
NUM|20|17|Let us pass, I pray thee, through thy country: we will not pass through the fields, or through the vineyards, neither will we drink of the water of the wells: we will go by the king's high way, we will not turn to the right hand nor to the left, until we have passed thy borders.
NUM|20|18|And Edom said unto him, Thou shalt not pass by me, lest I come out against thee with the sword.
NUM|20|19|And the children of Israel said unto him, We will go by the high way: and if I and my cattle drink of thy water, then I will pay for it: I will only, without doing anything else, go through on my feet.
NUM|20|20|And he said, Thou shalt not go through. And Edom came out against him with much people, and with a strong hand.
NUM|20|21|Thus Edom refused to give Israel passage through his border: wherefore Israel turned away from him.
NUM|20|22|And the children of Israel, even the whole congregation, journeyed from Kadesh, and came unto mount Hor.
NUM|20|23|And the LORD spake unto Moses and Aaron in mount Hor, by the coast of the land of Edom, saying,
NUM|20|24|Aaron shall be gathered unto his people: for he shall not enter into the land which I have given unto the children of Israel, because ye rebelled against my word at the water of Meribah.
NUM|20|25|Take Aaron and Eleazar his son, and bring them up unto mount Hor:
NUM|20|26|And strip Aaron of his garments, and put them upon Eleazar his son: and Aaron shall be gathered unto his people, and shall die there.
NUM|20|27|And Moses did as the LORD commanded: and they went up into mount Hor in the sight of all the congregation.
NUM|20|28|And Moses stripped Aaron of his garments, and put them upon Eleazar his son; and Aaron died there in the top of the mount: and Moses and Eleazar came down from the mount.
NUM|20|29|And when all the congregation saw that Aaron was dead, they mourned for Aaron thirty days, even all the house of Israel.
NUM|21|1|And when king Arad the Canaanite, which dwelt in the south, heard tell that Israel came by the way of the spies; then he fought against Israel, and took some of them prisoners.
NUM|21|2|And Israel vowed a vow unto the LORD, and said, If thou wilt indeed deliver this people into my hand, then I will utterly destroy their cities.
NUM|21|3|And the LORD hearkened to the voice of Israel, and delivered up the Canaanites; and they utterly destroyed them and their cities: and he called the name of the place Hormah.
NUM|21|4|And they journeyed from mount Hor by the way of the Red sea, to compass the land of Edom: and the soul of the people was much discouraged because of the way.
NUM|21|5|And the people spake against God, and against Moses, Wherefore have ye brought us up out of Egypt to die in the wilderness? for there is no bread, neither is there any water; and our soul loatheth this light bread.
NUM|21|6|And the LORD sent fiery serpents among the people, and they bit the people; and much people of Israel died.
NUM|21|7|Therefore the people came to Moses, and said, We have sinned, for we have spoken against the LORD, and against thee; pray unto the LORD, that he take away the serpents from us. And Moses prayed for the people.
NUM|21|8|And the LORD said unto Moses, Make thee a fiery serpent, and set it upon a pole: and it shall come to pass, that every one that is bitten, when he looketh upon it, shall live.
NUM|21|9|And Moses made a serpent of brass, and put it upon a pole, and it came to pass, that if a serpent had bitten any man, when he beheld the serpent of brass, he lived.
NUM|21|10|And the children of Israel set forward, and pitched in Oboth.
NUM|21|11|And they journeyed from Oboth, and pitched at Ijeabarim, in the wilderness which is before Moab, toward the sunrising.
NUM|21|12|From thence they removed, and pitched in the valley of Zared.
NUM|21|13|From thence they removed, and pitched on the other side of Arnon, which is in the wilderness that cometh out of the coasts of the Amorites: for Arnon is the border of Moab, between Moab and the Amorites.
NUM|21|14|Wherefore it is said in the book of the wars of the LORD, What he did in the Red sea, and in the brooks of Arnon,
NUM|21|15|And at the stream of the brooks that goeth down to the dwelling of Ar, and lieth upon the border of Moab.
NUM|21|16|And from thence they went to Beer: that is the well whereof the LORD spake unto Moses, Gather the people together, and I will give them water.
NUM|21|17|Then Israel sang this song, Spring up, O well; sing ye unto it:
NUM|21|18|The princes digged the well, the nobles of the people digged it, by the direction of the lawgiver, with their staves. And from the wilderness they went to Mattanah:
NUM|21|19|And from Mattanah to Nahaliel: and from Nahaliel to Bamoth:
NUM|21|20|And from Bamoth in the valley, that is in the country of Moab, to the top of Pisgah, which looketh toward Jeshimon.
NUM|21|21|And Israel sent messengers unto Sihon king of the Amorites, saying,
NUM|21|22|Let me pass through thy land: we will not turn into the fields, or into the vineyards; we will not drink of the waters of the well: but we will go along by the king's high way, until we be past thy borders.
NUM|21|23|And Sihon would not suffer Israel to pass through his border: but Sihon gathered all his people together, and went out against Israel into the wilderness: and he came to Jahaz, and fought against Israel.
NUM|21|24|And Israel smote him with the edge of the sword, and possessed his land from Arnon unto Jabbok, even unto the children of Ammon: for the border of the children of Ammon was strong.
NUM|21|25|And Israel took all these cities: and Israel dwelt in all the cities of the Amorites, in Heshbon, and in all the villages thereof.
NUM|21|26|For Heshbon was the city of Sihon the king of the Amorites, who had fought against the former king of Moab, and taken all his land out of his hand, even unto Arnon.
NUM|21|27|Wherefore they that speak in proverbs say, Come into Heshbon, let the city of Sihon be built and prepared:
NUM|21|28|For there is a fire gone out of Heshbon, a flame from the city of Sihon: it hath consumed Ar of Moab, and the lords of the high places of Arnon.
NUM|21|29|Woe to thee, Moab! thou art undone, O people of Chemosh: he hath given his sons that escaped, and his daughters, into captivity unto Sihon king of the Amorites.
NUM|21|30|We have shot at them; Heshbon is perished even unto Dibon, and we have laid them waste even unto Nophah, which reacheth unto Medeba.
NUM|21|31|Thus Israel dwelt in the land of the Amorites.
NUM|21|32|And Moses sent to spy out Jaazer, and they took the villages thereof, and drove out the Amorites that were there.
NUM|21|33|And they turned and went up by the way of Bashan: and Og the king of Bashan went out against them, he, and all his people, to the battle at Edrei.
NUM|21|34|And the LORD said unto Moses, Fear him not: for I have delivered him into thy hand, and all his people, and his land; and thou shalt do to him as thou didst unto Sihon king of the Amorites, which dwelt at Heshbon.
NUM|21|35|So they smote him, and his sons, and all his people, until there was none left him alive: and they possessed his land.
NUM|22|1|And the children of Israel set forward, and pitched in the plains of Moab on this side Jordan by Jericho.
NUM|22|2|And Balak the son of Zippor saw all that Israel had done to the Amorites.
NUM|22|3|And Moab was sore afraid of the people, because they were many: and Moab was distressed because of the children of Israel.
NUM|22|4|And Moab said unto the elders of Midian, Now shall this company lick up all that are round about us, as the ox licketh up the grass of the field. And Balak the son of Zippor was king of the Moabites at that time.
NUM|22|5|He sent messengers therefore unto Balaam the son of Beor to Pethor, which is by the river of the land of the children of his people, to call him, saying, Behold, there is a people come out from Egypt: behold, they cover the face of the earth, and they abide over against me:
NUM|22|6|Come now therefore, I pray thee, curse me this people; for they are too mighty for me: peradventure I shall prevail, that we may smite them, and that I may drive them out of the land: for I wot that he whom thou blessest is blessed, and he whom thou cursest is cursed.
NUM|22|7|And the elders of Moab and the elders of Midian departed with the rewards of divination in their hand; and they came unto Balaam, and spake unto him the words of Balak.
NUM|22|8|And he said unto them, Lodge here this night, and I will bring you word again, as the LORD shall speak unto me: and the princes of Moab abode with Balaam.
NUM|22|9|And God came unto Balaam, and said, What men are these with thee?
NUM|22|10|And Balaam said unto God, Balak the son of Zippor, king of Moab, hath sent unto me, saying,
NUM|22|11|Behold, there is a people come out of Egypt, which covereth the face of the earth: come now, curse me them; peradventure I shall be able to overcome them, and drive them out.
NUM|22|12|And God said unto Balaam, Thou shalt not go with them; thou shalt not curse the people: for they are blessed.
NUM|22|13|And Balaam rose up in the morning, and said unto the princes of Balak, Get you into your land: for the LORD refuseth to give me leave to go with you.
NUM|22|14|And the princes of Moab rose up, and they went unto Balak, and said, Balaam refuseth to come with us.
NUM|22|15|And Balak sent yet again princes, more, and more honorable than they.
NUM|22|16|And they came to Balaam, and said to him, Thus saith Balak the son of Zippor, Let nothing, I pray thee, hinder thee from coming unto me:
NUM|22|17|For I will promote thee unto very great honor, and I will do whatsoever thou sayest unto me: come therefore, I pray thee, curse me this people.
NUM|22|18|And Balaam answered and said unto the servants of Balak, If Balak would give me his house full of silver and gold, I cannot go beyond the word of the LORD my God, to do less or more.
NUM|22|19|Now therefore, I pray you, tarry ye also here this night, that I may know what the LORD will say unto me more.
NUM|22|20|And God came unto Balaam at night, and said unto him, If the men come to call thee, rise up, and go with them; but yet the word which I shall say unto thee, that shalt thou do.
NUM|22|21|And Balaam rose up in the morning, and saddled his ass, and went with the princes of Moab.
NUM|22|22|And God's anger was kindled because he went: and the angel of the LORD stood in the way for an adversary against him. Now he was riding upon his ass, and his two servants were with him.
NUM|22|23|And the ass saw the angel of the LORD standing in the way, and his sword drawn in his hand: and the ass turned aside out of the way, and went into the field: and Balaam smote the ass, to turn her into the way.
NUM|22|24|But the angel of the LORD stood in a path of the vineyards, a wall being on this side, and a wall on that side.
NUM|22|25|And when the ass saw the angel of the LORD, she thrust herself unto the wall, and crushed Balaam's foot against the wall: and he smote her again.
NUM|22|26|And the angel of the LORD went further, and stood in a narrow place, where was no way to turn either to the right hand or to the left.
NUM|22|27|And when the ass saw the angel of the LORD, she fell down under Balaam: and Balaam's anger was kindled, and he smote the ass with a staff.
NUM|22|28|And the LORD opened the mouth of the ass, and she said unto Balaam, What have I done unto thee, that thou hast smitten me these three times?
NUM|22|29|And Balaam said unto the ass, Because thou hast mocked me: I would there were a sword in mine hand, for now would I kill thee.
NUM|22|30|And the ass said unto Balaam, Am not I thine ass, upon which thou hast ridden ever since I was thine unto this day? was I ever wont to do so unto thee? And he said, Nay.
NUM|22|31|Then the LORD opened the eyes of Balaam, and he saw the angel of the LORD standing in the way, and his sword drawn in his hand: and he bowed down his head, and fell flat on his face.
NUM|22|32|And the angel of the LORD said unto him, Wherefore hast thou smitten thine ass these three times? behold, I went out to withstand thee, because thy way is perverse before me:
NUM|22|33|And the ass saw me, and turned from me these three times: unless she had turned from me, surely now also I had slain thee, and saved her alive.
NUM|22|34|And Balaam said unto the angel of the LORD, I have sinned; for I knew not that thou stoodest in the way against me: now therefore, if it displease thee, I will get me back again.
NUM|22|35|And the angel of the LORD said unto Balaam, Go with the men: but only the word that I shall speak unto thee, that thou shalt speak. So Balaam went with the princes of Balak.
NUM|22|36|And when Balak heard that Balaam was come, he went out to meet him unto a city of Moab, which is in the border of Arnon, which is in the utmost coast.
NUM|22|37|And Balak said unto Balaam, Did I not earnestly send unto thee to call thee? wherefore camest thou not unto me? am I not able indeed to promote thee to honor?
NUM|22|38|And Balaam said unto Balak, Lo, I am come unto thee: have I now any power at all to say any thing? the word that God putteth in my mouth, that shall I speak.
NUM|22|39|And Balaam went with Balak, and they came unto Kirjathhuzoth.
NUM|22|40|And Balak offered oxen and sheep, and sent to Balaam, and to the princes that were with him.
NUM|22|41|And it came to pass on the morrow, that Balak took Balaam, and brought him up into the high places of Baal, that thence he might see the utmost part of the people.
NUM|23|1|And Balaam said unto Balak, Build me here seven altars, and prepare me here seven oxen and seven rams.
NUM|23|2|And Balak did as Balaam had spoken; and Balak and Balaam offered on every altar a bullock and a ram.
NUM|23|3|And Balaam said unto Balak, Stand by thy burnt offering, and I will go: peradventure the LORD will come to meet me: and whatsoever he showeth me I will tell thee. And he went to an high place.
NUM|23|4|And God met Balaam: and he said unto him, I have prepared seven altars, and I have offered upon every altar a bullock and a ram.
NUM|23|5|And the LORD put a word in Balaam's mouth, and said, Return unto Balak, and thus thou shalt speak.
NUM|23|6|And he returned unto him, and, lo, he stood by his burnt sacrifice, he, and all the princes of Moab.
NUM|23|7|And he took up his parable, and said, Balak the king of Moab hath brought me from Aram, out of the mountains of the east, saying, Come, curse me Jacob, and come, defy Israel.
NUM|23|8|How shall I curse, whom God hath not cursed? or how shall I defy, whom the LORD hath not defied?
NUM|23|9|For from the top of the rocks I see him, and from the hills I behold him: lo, the people shall dwell alone, and shall not be reckoned among the nations.
NUM|23|10|Who can count the dust of Jacob, and the number of the fourth part of Israel? Let me die the death of the righteous, and let my last end be like his!
NUM|23|11|And Balak said unto Balaam, What hast thou done unto me? I took thee to curse mine enemies, and, behold, thou hast blessed them altogether.
NUM|23|12|And he answered and said, Must I not take heed to speak that which the LORD hath put in my mouth?
NUM|23|13|And Balak said unto him, Come, I pray thee, with me unto another place, from whence thou mayest see them: thou shalt see but the utmost part of them, and shalt not see them all: and curse me them from thence.
NUM|23|14|And he brought him into the field of Zophim, to the top of Pisgah, and built seven altars, and offered a bullock and a ram on every altar.
NUM|23|15|And he said unto Balak, Stand here by thy burnt offering, while I meet the LORD yonder.
NUM|23|16|And the LORD met Balaam, and put a word in his mouth, and said, Go again unto Balak, and say thus.
NUM|23|17|And when he came to him, behold, he stood by his burnt offering, and the princes of Moab with him. And Balak said unto him, What hath the LORD spoken?
NUM|23|18|And he took up his parable, and said, Rise up, Balak, and hear; hearken unto me, thou son of Zippor:
NUM|23|19|God is not a man, that he should lie; neither the son of man, that he should repent: hath he said, and shall he not do it? or hath he spoken, and shall he not make it good?
NUM|23|20|Behold, I have received commandment to bless: and he hath blessed; and I cannot reverse it.
NUM|23|21|He hath not beheld iniquity in Jacob, neither hath he seen perverseness in Israel: the LORD his God is with him, and the shout of a king is among them.
NUM|23|22|God brought them out of Egypt; he hath as it were the strength of an unicorn.
NUM|23|23|Surely there is no enchantment against Jacob, neither is there any divination against Israel: according to this time it shall be said of Jacob and of Israel, What hath God wrought!
NUM|23|24|Behold, the people shall rise up as a great lion, and lift up himself as a young lion: he shall not lie down until he eat of the prey, and drink the blood of the slain.
NUM|23|25|And Balak said unto Balaam, Neither curse them at all, nor bless them at all.
NUM|23|26|But Balaam answered and said unto Balak, Told not I thee, saying, All that the LORD speaketh, that I must do?
NUM|23|27|And Balak said unto Balaam, Come, I pray thee, I will bring thee unto another place; peradventure it will please God that thou mayest curse me them from thence.
NUM|23|28|And Balak brought Balaam unto the top of Peor, that looketh toward Jeshimon.
NUM|23|29|And Balaam said unto Balak, Build me here seven altars, and prepare me here seven bullocks and seven rams.
NUM|23|30|And Balak did as Balaam had said, and offered a bullock and a ram on every altar.
NUM|24|1|And when Balaam saw that it pleased the LORD to bless Israel, he went not, as at other times, to seek for enchantments, but he set his face toward the wilderness.
NUM|24|2|And Balaam lifted up his eyes, and he saw Israel abiding in his tents according to their tribes; and the spirit of God came upon him.
NUM|24|3|And he took up his parable, and said, Balaam the son of Beor hath said, and the man whose eyes are open hath said:
NUM|24|4|He hath said, which heard the words of God, which saw the vision of the Almighty, falling into a trance, but having his eyes open:
NUM|24|5|How goodly are thy tents, O Jacob, and thy tabernacles, O Israel!
NUM|24|6|As the valleys are they spread forth, as gardens by the river's side, as the trees of lign aloes which the LORD hath planted, and as cedar trees beside the waters.
NUM|24|7|He shall pour the water out of his buckets, and his seed shall be in many waters, and his king shall be higher than Agag, and his kingdom shall be exalted.
NUM|24|8|God brought him forth out of Egypt; he hath as it were the strength of an unicorn: he shall eat up the nations his enemies, and shall break their bones, and pierce them through with his arrows.
NUM|24|9|He couched, he lay down as a lion, and as a great lion: who shall stir him up? Blessed is he that blesseth thee, and cursed is he that curseth thee.
NUM|24|10|And Balak's anger was kindled against Balaam, and he smote his hands together: and Balak said unto Balaam, I called thee to curse mine enemies, and, behold, thou hast altogether blessed them these three times.
NUM|24|11|Therefore now flee thou to thy place: I thought to promote thee unto great honor; but, lo, the LORD hath kept thee back from honor.
NUM|24|12|And Balaam said unto Balak, Spake I not also to thy messengers which thou sentest unto me, saying,
NUM|24|13|If Balak would give me his house full of silver and gold, I cannot go beyond the commandment of the LORD, to do either good or bad of mine own mind; but what the LORD saith, that will I speak?
NUM|24|14|And now, behold, I go unto my people: come therefore, and I will advertise thee what this people shall do to thy people in the latter days.
NUM|24|15|And he took up his parable, and said, Balaam the son of Beor hath said, and the man whose eyes are open hath said:
NUM|24|16|He hath said, which heard the words of God, and knew the knowledge of the most High, which saw the vision of the Almighty, falling into a trance, but having his eyes open:
NUM|24|17|I shall see him, but not now: I shall behold him, but not nigh: there shall come a Star out of Jacob, and a Sceptre shall rise out of Israel, and shall smite the corners of Moab, and destroy all the children of Sheth.
NUM|24|18|And Edom shall be a possession, Seir also shall be a possession for his enemies; and Israel shall do valiantly.
NUM|24|19|Out of Jacob shall come he that shall have dominion, and shall destroy him that remaineth of the city.
NUM|24|20|And when he looked on Amalek, he took up his parable, and said, Amalek was the first of the nations; but his latter end shall be that he perish for ever.
NUM|24|21|And he looked on the Kenites, and took up his parable, and said, Strong is thy dwelling place, and thou puttest thy nest in a rock.
NUM|24|22|Nevertheless the Kenite shall be wasted, until Asshur shall carry thee away captive.
NUM|24|23|And he took up his parable, and said, Alas, who shall live when God doeth this!
NUM|24|24|And ships shall come from the coast of Chittim, and shall afflict Asshur, and shall afflict Eber, and he also shall perish for ever.
NUM|24|25|And Balaam rose up, and went and returned to his place: and Balak also went his way.
NUM|25|1|And Israel abode in Shittim, and the people began to commit whoredom with the daughters of Moab.
NUM|25|2|And they called the people unto the sacrifices of their gods: and the people did eat, and bowed down to their gods.
NUM|25|3|And Israel joined himself unto Baalpeor: and the anger of the LORD was kindled against Israel.
NUM|25|4|And the LORD said unto Moses, Take all the heads of the people, and hang them up before the LORD against the sun, that the fierce anger of the LORD may be turned away from Israel.
NUM|25|5|And Moses said unto the judges of Israel, Slay ye every one his men that were joined unto Baalpeor.
NUM|25|6|And, behold, one of the children of Israel came and brought unto his brethren a Midianitish woman in the sight of Moses, and in the sight of all the congregation of the children of Israel, who were weeping before the door of the tabernacle of the congregation.
NUM|25|7|And when Phinehas, the son of Eleazar, the son of Aaron the priest, saw it, he rose up from among the congregation, and took a javelin in his hand;
NUM|25|8|And he went after the man of Israel into the tent, and thrust both of them through, the man of Israel, and the woman through her belly. So the plague was stayed from the children of Israel.
NUM|25|9|And those that died in the plague were twenty and four thousand.
NUM|25|10|And the LORD spake unto Moses, saying,
NUM|25|11|Phinehas, the son of Eleazar, the son of Aaron the priest, hath turned my wrath away from the children of Israel, while he was zealous for my sake among them, that I consumed not the children of Israel in my jealousy.
NUM|25|12|Wherefore say, Behold, I give unto him my covenant of peace:
NUM|25|13|And he shall have it, and his seed after him, even the covenant of an everlasting priesthood; because he was zealous for his God, and made an atonement for the children of Israel.
NUM|25|14|Now the name of the Israelite that was slain, even that was slain with the Midianitish woman, was Zimri, the son of Salu, a prince of a chief house among the Simeonites.
NUM|25|15|And the name of the Midianitish woman that was slain was Cozbi, the daughter of Zur; he was head over a people, and of a chief house in Midian.
NUM|25|16|And the LORD spake unto Moses, saying,
NUM|25|17|Vex the Midianites, and smite them:
NUM|25|18|For they vex you with their wiles, wherewith they have beguiled you in the matter of Peor, and in the matter of Cozbi, the daughter of a prince of Midian, their sister, which was slain in the day of the plague for Peor's sake.
NUM|26|1|And it came to pass after the plague, that the LORD spake unto Moses and unto Eleazar the son of Aaron the priest, saying,
NUM|26|2|Take the sum of all the congregation of the children of Israel, from twenty years old and upward, throughout their fathers' house, all that are able to go to war in Israel.
NUM|26|3|And Moses and Eleazar the priest spake with them in the plains of Moab by Jordan near Jericho, saying,
NUM|26|4|Take the sum of the people, from twenty years old and upward; as the LORD commanded Moses and the children of Israel, which went forth out of the land of Egypt.
NUM|26|5|Reuben, the eldest son of Israel: the children of Reuben; Hanoch, of whom cometh the family of the Hanochites: of Pallu, the family of the Palluites:
NUM|26|6|Of Hezron, the family of the Hezronites: of Carmi, the family of the Carmites.
NUM|26|7|These are the families of the Reubenites: and they that were numbered of them were forty and three thousand and seven hundred and thirty.
NUM|26|8|And the sons of Pallu; Eliab.
NUM|26|9|And the sons of Eliab; Nemuel, and Dathan, and Abiram. This is that Dathan and Abiram, which were famous in the congregation, who strove against Moses and against Aaron in the company of Korah, when they strove against the LORD:
NUM|26|10|And the earth opened her mouth, and swallowed them up together with Korah, when that company died, what time the fire devoured two hundred and fifty men: and they became a sign.
NUM|26|11|Notwithstanding the children of Korah died not.
NUM|26|12|The sons of Simeon after their families: of Nemuel, the family of the Nemuelites: of Jamin, the family of the Jaminites: of Jachin, the family of the Jachinites:
NUM|26|13|Of Zerah, the family of the Zarhites: of Shaul, the family of the Shaulites.
NUM|26|14|These are the families of the Simeonites, twenty and two thousand and two hundred.
NUM|26|15|The children of Gad after their families: of Zephon, the family of the Zephonites: of Haggi, the family of the Haggites: of Shuni, the family of the Shunites:
NUM|26|16|Of Ozni, the family of the Oznites: of Eri, the family of the Erites:
NUM|26|17|Of Arod, the family of the Arodites: of Areli, the family of the Arelites.
NUM|26|18|These are the families of the children of Gad according to those that were numbered of them, forty thousand and five hundred.
NUM|26|19|The sons of Judah were Er and Onan: and Er and Onan died in the land of Canaan.
NUM|26|20|And the sons of Judah after their families were; of Shelah, the family of the Shelanites: of Pharez, the family of the Pharzites: of Zerah, the family of the Zarhites.
NUM|26|21|And the sons of Pharez were; of Hezron, the family of the Hezronites: of Hamul, the family of the Hamulites.
NUM|26|22|These are the families of Judah according to those that were numbered of them, threescore and sixteen thousand and five hundred.
NUM|26|23|Of the sons of Issachar after their families: of Tola, the family of the Tolaites: of Pua, the family of the Punites:
NUM|26|24|Of Jashub, the family of the Jashubites: of Shimron, the family of the Shimronites.
NUM|26|25|These are the families of Issachar according to those that were numbered of them, threescore and four thousand and three hundred.
NUM|26|26|Of the sons of Zebulun after their families: of Sered, the family of the Sardites: of Elon, the family of the Elonites: of Jahleel, the family of the Jahleelites.
NUM|26|27|These are the families of the Zebulunites according to those that were numbered of them, threescore thousand and five hundred.
NUM|26|28|The sons of Joseph after their families were Manasseh and Ephraim.
NUM|26|29|Of the sons of Manasseh: of Machir, the family of the Machirites: and Machir begat Gilead: of Gilead come the family of the Gileadites.
NUM|26|30|These are the sons of Gilead: of Jeezer, the family of the Jeezerites: of Helek, the family of the Helekites:
NUM|26|31|And of Asriel, the family of the Asrielites: and of Shechem, the family of the Shechemites:
NUM|26|32|And of Shemida, the family of the Shemidaites: and of Hepher, the family of the Hepherites.
NUM|26|33|And Zelophehad the son of Hepher had no sons, but daughters: and the names of the daughters of Zelophehad were Mahlah, and Noah, Hoglah, Milcah, and Tirzah.
NUM|26|34|These are the families of Manasseh, and those that were numbered of them, fifty and two thousand and seven hundred.
NUM|26|35|These are the sons of Ephraim after their families: of Shuthelah, the family of the Shuthalhites: of Becher, the family of the Bachrites: of Tahan, the family of the Tahanites.
NUM|26|36|And these are the sons of Shuthelah: of Eran, the family of the Eranites.
NUM|26|37|These are the families of the sons of Ephraim according to those that were numbered of them, thirty and two thousand and five hundred. These are the sons of Joseph after their families.
NUM|26|38|The sons of Benjamin after their families: of Bela, the family of the Belaites: of Ashbel, the family of the Ashbelites: of Ahiram, the family of the Ahiramites:
NUM|26|39|Of Shupham, the family of the Shuphamites: of Hupham, the family of the Huphamites.
NUM|26|40|And the sons of Bela were Ard and Naaman: of Ard, the family of the Ardites: and of Naaman, the family of the Naamites.
NUM|26|41|These are the sons of Benjamin after their families: and they that were numbered of them were forty and five thousand and six hundred.
NUM|26|42|These are the sons of Dan after their families: of Shuham, the family of the Shuhamites. These are the families of Dan after their families.
NUM|26|43|All the families of the Shuhamites, according to those that were numbered of them, were threescore and four thousand and four hundred.
NUM|26|44|Of the children of Asher after their families: of Jimna, the family of the Jimnites: of Jesui, the family of the Jesuites: of Beriah, the family of the Beriites.
NUM|26|45|Of the sons of Beriah: of Heber, the family of the Heberites: of Malchiel, the family of the Malchielites.
NUM|26|46|And the name of the daughter of Asher was Sarah.
NUM|26|47|These are the families of the sons of Asher according to those that were numbered of them; who were fifty and three thousand and four hundred.
NUM|26|48|Of the sons of Naphtali after their families: of Jahzeel, the family of the Jahzeelites: of Guni, the family of the Gunites:
NUM|26|49|Of Jezer, the family of the Jezerites: of Shillem, the family of the Shillemites.
NUM|26|50|These are the families of Naphtali according to their families: and they that were numbered of them were forty and five thousand and four hundred.
NUM|26|51|These were the numbered of the children of Israel, six hundred thousand and a thousand seven hundred and thirty.
NUM|26|52|And the LORD spake unto Moses, saying,
NUM|26|53|Unto these the land shall be divided for an inheritance according to the number of names.
NUM|26|54|To many thou shalt give the more inheritance, and to few thou shalt give the less inheritance: to every one shall his inheritance be given according to those that were numbered of him.
NUM|26|55|Notwithstanding the land shall be divided by lot: according to the names of the tribes of their fathers they shall inherit.
NUM|26|56|According to the lot shall the possession thereof be divided between many and few.
NUM|26|57|And these are they that were numbered of the Levites after their families: of Gershon, the family of the Gershonites: of Kohath, the family of the Kohathites: of Merari, the family of the Merarites.
NUM|26|58|These are the families of the Levites: the family of the Libnites, the family of the Hebronites, the family of the Mahlites, the family of the Mushites, the family of the Korathites. And Kohath begat Amram.
NUM|26|59|And the name of Amram's wife was Jochebed, the daughter of Levi, whom her mother bare to Levi in Egypt: and she bare unto Amram Aaron and Moses, and Miriam their sister.
NUM|26|60|And unto Aaron was born Nadab, and Abihu, Eleazar, and Ithamar.
NUM|26|61|And Nadab and Abihu died, when they offered strange fire before the LORD.
NUM|26|62|And those that were numbered of them were twenty and three thousand, all males from a month old and upward: for they were not numbered among the children of Israel, because there was no inheritance given them among the children of Israel.
NUM|26|63|These are they that were numbered by Moses and Eleazar the priest, who numbered the children of Israel in the plains of Moab by Jordan near Jericho.
NUM|26|64|But among these there was not a man of them whom Moses and Aaron the priest numbered, when they numbered the children of Israel in the wilderness of Sinai.
NUM|26|65|For the LORD had said of them, They shall surely die in the wilderness. And there was not left a man of them, save Caleb the son of Jephunneh, and Joshua the son of Nun.
NUM|27|1|Then came the daughters of Zelophehad, the son of Hepher, the son of Gilead, the son of Machir, the son of Manasseh, of the families of Manasseh the son of Joseph: and these are the names of his daughters; Mahlah, Noah, and Hoglah, and Milcah, and Tirzah.
NUM|27|2|And they stood before Moses, and before Eleazar the priest, and before the princes and all the congregation, by the door of the tabernacle of the congregation, saying,
NUM|27|3|Our father died in the wilderness, and he was not in the company of them that gathered themselves together against the LORD in the company of Korah; but died in his own sin, and had no sons.
NUM|27|4|Why should the name of our father be done away from among his family, because he hath no son? Give unto us therefore a possession among the brethren of our father.
NUM|27|5|And Moses brought their cause before the LORD.
NUM|27|6|And the LORD spake unto Moses, saying,
NUM|27|7|The daughters of Zelophehad speak right: thou shalt surely give them a possession of an inheritance among their father's brethren; and thou shalt cause the inheritance of their father to pass unto them.
NUM|27|8|And thou shalt speak unto the children of Israel, saying, If a man die, and have no son, then ye shall cause his inheritance to pass unto his daughter.
NUM|27|9|And if he have no daughter, then ye shall give his inheritance unto his brethren.
NUM|27|10|And if he have no brethren, then ye shall give his inheritance unto his father's brethren.
NUM|27|11|And if his father have no brethren, then ye shall give his inheritance unto his kinsman that is next to him of his family, and he shall possess it: and it shall be unto the children of Israel a statute of judgment, as the LORD commanded Moses.
NUM|27|12|And the LORD said unto Moses, Get thee up into this mount Abarim, and see the land which I have given unto the children of Israel.
NUM|27|13|And when thou hast seen it, thou also shalt be gathered unto thy people, as Aaron thy brother was gathered.
NUM|27|14|For ye rebelled against my commandment in the desert of Zin, in the strife of the congregation, to sanctify me at the water before their eyes: that is the water of Meribah in Kadesh in the wilderness of Zin.
NUM|27|15|And Moses spake unto the LORD, saying,
NUM|27|16|Let the LORD, the God of the spirits of all flesh, set a man over the congregation,
NUM|27|17|Which may go out before them, and which may go in before them, and which may lead them out, and which may bring them in; that the congregation of the LORD be not as sheep which have no shepherd.
NUM|27|18|And the LORD said unto Moses, Take thee Joshua the son of Nun, a man in whom is the spirit, and lay thine hand upon him;
NUM|27|19|And set him before Eleazar the priest, and before all the congregation; and give him a charge in their sight.
NUM|27|20|And thou shalt put some of thine honor upon him, that all the congregation of the children of Israel may be obedient.
NUM|27|21|And he shall stand before Eleazar the priest, who shall ask counsel for him after the judgment of Urim before the LORD: at his word shall they go out, and at his word they shall come in, both he, and all the children of Israel with him, even all the congregation.
NUM|27|22|And Moses did as the LORD commanded him: and he took Joshua, and set him before Eleazar the priest, and before all the congregation:
NUM|27|23|And he laid his hands upon him, and gave him a charge, as the LORD commanded by the hand of Moses.
NUM|28|1|And the LORD spake unto Moses, saying,
NUM|28|2|Command the children of Israel, and say unto them, My offering, and my bread for my sacrifices made by fire, for a sweet savor unto me, shall ye observe to offer unto me in their due season.
NUM|28|3|And thou shalt say unto them, This is the offering made by fire which ye shall offer unto the LORD; two lambs of the first year without spot day by day, for a continual burnt offering.
NUM|28|4|The one lamb shalt thou offer in the morning, and the other lamb shalt thou offer at even;
NUM|28|5|And a tenth part of an ephah of flour for a meat offering, mingled with the fourth part of an hin of beaten oil.
NUM|28|6|It is a continual burnt offering, which was ordained in mount Sinai for a sweet savor, a sacrifice made by fire unto the LORD.
NUM|28|7|And the drink offering thereof shall be the fourth part of an hin for the one lamb: in the holy place shalt thou cause the strong wine to be poured unto the LORD for a drink offering.
NUM|28|8|And the other lamb shalt thou offer at even: as the meat offering of the morning, and as the drink offering thereof, thou shalt offer it, a sacrifice made by fire, of a sweet savor unto the LORD.
NUM|28|9|And on the sabbath day two lambs of the first year without spot, and two tenth deals of flour for a meat offering, mingled with oil, and the drink offering thereof:
NUM|28|10|This is the burnt offering of every sabbath, beside the continual burnt offering, and his drink offering.
NUM|28|11|And in the beginnings of your months ye shall offer a burnt offering unto the LORD; two young bullocks, and one ram, seven lambs of the first year without spot;
NUM|28|12|And three tenth deals of flour for a meat offering, mingled with oil, for one bullock; and two tenth deals of flour for a meat offering, mingled with oil, for one ram;
NUM|28|13|And a several tenth deal of flour mingled with oil for a meat offering unto one lamb; for a burnt offering of a sweet savor, a sacrifice made by fire unto the LORD.
NUM|28|14|And their drink offerings shall be half an hin of wine unto a bullock, and the third part of an hin unto a ram, and a fourth part of an hin unto a lamb: this is the burnt offering of every month throughout the months of the year.
NUM|28|15|And one kid of the goats for a sin offering unto the LORD shall be offered, beside the continual burnt offering, and his drink offering.
NUM|28|16|And in the fourteenth day of the first month is the passover of the LORD.
NUM|28|17|And in the fifteenth day of this month is the feast: seven days shall unleavened bread be eaten.
NUM|28|18|In the first day shall be an holy convocation; ye shall do no manner of servile work therein:
NUM|28|19|But ye shall offer a sacrifice made by fire for a burnt offering unto the LORD; two young bullocks, and one ram, and seven lambs of the first year: they shall be unto you without blemish:
NUM|28|20|And their meat offering shall be of flour mingled with oil: three tenth deals shall ye offer for a bullock, and two tenth deals for a ram;
NUM|28|21|A several tenth deal shalt thou offer for every lamb, throughout the seven lambs:
NUM|28|22|And one goat for a sin offering, to make an atonement for you.
NUM|28|23|Ye shall offer these beside the burnt offering in the morning, which is for a continual burnt offering.
NUM|28|24|After this manner ye shall offer daily, throughout the seven days, the meat of the sacrifice made by fire, of a sweet savor unto the LORD: it shall be offered beside the continual burnt offering, and his drink offering.
NUM|28|25|And on the seventh day ye shall have an holy convocation; ye shall do no servile work.
NUM|28|26|Also in the day of the firstfruits, when ye bring a new meat offering unto the LORD, after your weeks be out, ye shall have an holy convocation; ye shall do no servile work:
NUM|28|27|But ye shall offer the burnt offering for a sweet savor unto the LORD; two young bullocks, one ram, seven lambs of the first year;
NUM|28|28|And their meat offering of flour mingled with oil, three tenth deals unto one bullock, two tenth deals unto one ram,
NUM|28|29|A several tenth deal unto one lamb, throughout the seven lambs;
NUM|28|30|And one kid of the goats, to make an atonement for you.
NUM|28|31|Ye shall offer them beside the continual burnt offering, and his meat offering, (they shall be unto you without blemish) and their drink offerings.
NUM|29|1|And in the seventh month, on the first day of the month, ye shall have an holy convocation; ye shall do no servile work: it is a day of blowing the trumpets unto you.
NUM|29|2|And ye shall offer a burnt offering for a sweet savor unto the LORD; one young bullock, one ram, and seven lambs of the first year without blemish:
NUM|29|3|And their meat offering shall be of flour mingled with oil, three tenth deals for a bullock, and two tenth deals for a ram,
NUM|29|4|And one tenth deal for one lamb, throughout the seven lambs:
NUM|29|5|And one kid of the goats for a sin offering, to make an atonement for you:
NUM|29|6|Beside the burnt offering of the month, and his meat offering, and the daily burnt offering, and his meat offering, and their drink offerings, according unto their manner, for a sweet savor, a sacrifice made by fire unto the LORD.
NUM|29|7|And ye shall have on the tenth day of this seventh month an holy convocation; and ye shall afflict your souls: ye shall not do any work therein:
NUM|29|8|But ye shall offer a burnt offering unto the LORD for a sweet savor; one young bullock, one ram, and seven lambs of the first year; they shall be unto you without blemish:
NUM|29|9|And their meat offering shall be of flour mingled with oil, three tenth deals to a bullock, and two tenth deals to one ram,
NUM|29|10|A several tenth deal for one lamb, throughout the seven lambs:
NUM|29|11|One kid of the goats for a sin offering; beside the sin offering of atonement, and the continual burnt offering, and the meat offering of it, and their drink offerings.
NUM|29|12|And on the fifteenth day of the seventh month ye shall have an holy convocation; ye shall do no servile work, and ye shall keep a feast unto the LORD seven days:
NUM|29|13|And ye shall offer a burnt offering, a sacrifice made by fire, of a sweet savor unto the LORD; thirteen young bullocks, two rams, and fourteen lambs of the first year; they shall be without blemish:
NUM|29|14|And their meat offering shall be of flour mingled with oil, three tenth deals unto every bullock of the thirteen bullocks, two tenth deals to each ram of the two rams,
NUM|29|15|And a several tenth deal to each lamb of the fourteen lambs:
NUM|29|16|And one kid of the goats for a sin offering; beside the continual burnt offering, his meat offering, and his drink offering.
NUM|29|17|And on the second day ye shall offer twelve young bullocks, two rams, fourteen lambs of the first year without spot:
NUM|29|18|And their meat offering and their drink offerings for the bullocks, for the rams, and for the lambs, shall be according to their number, after the manner:
NUM|29|19|And one kid of the goats for a sin offering; beside the continual burnt offering, and the meat offering thereof, and their drink offerings.
NUM|29|20|And on the third day eleven bullocks, two rams, fourteen lambs of the first year without blemish;
NUM|29|21|And their meat offering and their drink offerings for the bullocks, for the rams, and for the lambs, shall be according to their number, after the manner:
NUM|29|22|And one goat for a sin offering; beside the continual burnt offering, and his meat offering, and his drink offering.
NUM|29|23|And on the fourth day ten bullocks, two rams, and fourteen lambs of the first year without blemish:
NUM|29|24|Their meat offering and their drink offerings for the bullocks, for the rams, and for the lambs, shall be according to their number, after the manner:
NUM|29|25|And one kid of the goats for a sin offering; beside the continual burnt offering, his meat offering, and his drink offering.
NUM|29|26|And on the fifth day nine bullocks, two rams, and fourteen lambs of the first year without spot:
NUM|29|27|And their meat offering and their drink offerings for the bullocks, for the rams, and for the lambs, shall be according to their number, after the manner:
NUM|29|28|And one goat for a sin offering; beside the continual burnt offering, and his meat offering, and his drink offering.
NUM|29|29|And on the sixth day eight bullocks, two rams, and fourteen lambs of the first year without blemish:
NUM|29|30|And their meat offering and their drink offerings for the bullocks, for the rams, and for the lambs, shall be according to their number, after the manner:
NUM|29|31|And one goat for a sin offering; beside the continual burnt offering, his meat offering, and his drink offering.
NUM|29|32|And on the seventh day seven bullocks, two rams, and fourteen lambs of the first year without blemish:
NUM|29|33|And their meat offering and their drink offerings for the bullocks, for the rams, and for the lambs, shall be according to their number, after the manner:
NUM|29|34|And one goat for a sin offering; beside the continual burnt offering, his meat offering, and his drink offering.
NUM|29|35|On the eighth day ye shall have a solemn assembly: ye shall do no servile work therein:
NUM|29|36|But ye shall offer a burnt offering, a sacrifice made by fire, of a sweet savor unto the LORD: one bullock, one ram, seven lambs of the first year without blemish:
NUM|29|37|Their meat offering and their drink offerings for the bullock, for the ram, and for the lambs, shall be according to their number, after the manner:
NUM|29|38|And one goat for a sin offering; beside the continual burnt offering, and his meat offering, and his drink offering.
NUM|29|39|These things ye shall do unto the LORD in your set feasts, beside your vows, and your freewill offerings, for your burnt offerings, and for your meat offerings, and for your drink offerings, and for your peace offerings.
NUM|29|40|And Moses told the children of Israel according to all that the LORD commanded Moses.
NUM|30|1|And Moses spake unto the heads of the tribes concerning the children of Israel, saying, This is the thing which the LORD hath commanded.
NUM|30|2|If a man vow a vow unto the LORD, or swear an oath to bind his soul with a bond; he shall not break his word, he shall do according to all that proceedeth out of his mouth.
NUM|30|3|If a woman also vow a vow unto the LORD, and bind herself by a bond, being in her father's house in her youth;
NUM|30|4|And her father hear her vow, and her bond wherewith she hath bound her soul, and her father shall hold his peace at her; then all her vows shall stand, and every bond wherewith she hath bound her soul shall stand.
NUM|30|5|But if her father disallow her in the day that he heareth; not any of her vows, or of her bonds wherewith she hath bound her soul, shall stand: and the LORD shall forgive her, because her father disallowed her.
NUM|30|6|And if she had at all an husband, when she vowed, or uttered ought out of her lips, wherewith she bound her soul;
NUM|30|7|And her husband heard it, and held his peace at her in the day that he heard it: then her vows shall stand, and her bonds wherewith she bound her soul shall stand.
NUM|30|8|But if her husband disallowed her on the day that he heard it; then he shall make her vow which she vowed, and that which she uttered with her lips, wherewith she bound her soul, of none effect: and the LORD shall forgive her.
NUM|30|9|But every vow of a widow, and of her that is divorced, wherewith they have bound their souls, shall stand against her.
NUM|30|10|And if she vowed in her husband's house, or bound her soul by a bond with an oath;
NUM|30|11|And her husband heard it, and held his peace at her, and disallowed her not: then all her vows shall stand, and every bond wherewith she bound her soul shall stand.
NUM|30|12|But if her husband hath utterly made them void on the day he heard them; then whatsoever proceeded out of her lips concerning her vows, or concerning the bond of her soul, shall not stand: her husband hath made them void; and the LORD shall forgive her.
NUM|30|13|Every vow, and every binding oath to afflict the soul, her husband may establish it, or her husband may make it void.
NUM|30|14|But if her husband altogether hold his peace at her from day to day; then he establisheth all her vows, or all her bonds, which are upon her: he confirmeth them, because he held his peace at her in the day that he heard them.
NUM|30|15|But if he shall any ways make them void after that he hath heard them; then he shall bear her iniquity.
NUM|30|16|These are the statutes, which the LORD commanded Moses, between a man and his wife, between the father and his daughter, being yet in her youth in her father's house.
NUM|31|1|And the LORD spake unto Moses, saying,
NUM|31|2|Avenge the children of Israel of the Midianites: afterward shalt thou be gathered unto thy people.
NUM|31|3|And Moses spake unto the people, saying, Arm some of yourselves unto the war, and let them go against the Midianites, and avenge the LORD of Midian.
NUM|31|4|Of every tribe a thousand, throughout all the tribes of Israel, shall ye send to the war.
NUM|31|5|So there were delivered out of the thousands of Israel, a thousand of every tribe, twelve thousand armed for war.
NUM|31|6|And Moses sent them to the war, a thousand of every tribe, them and Phinehas the son of Eleazar the priest, to the war, with the holy instruments, and the trumpets to blow in his hand.
NUM|31|7|And they warred against the Midianites, as the LORD commanded Moses; and they slew all the males.
NUM|31|8|And they slew the kings of Midian, beside the rest of them that were slain; namely, Evi, and Rekem, and Zur, and Hur, and Reba, five kings of Midian: Balaam also the son of Beor they slew with the sword.
NUM|31|9|And the children of Israel took all the women of Midian captives, and their little ones, and took the spoil of all their cattle, and all their flocks, and all their goods.
NUM|31|10|And they burnt all their cities wherein they dwelt, and all their goodly castles, with fire.
NUM|31|11|And they took all the spoil, and all the prey, both of men and of beasts.
NUM|31|12|And they brought the captives, and the prey, and the spoil, unto Moses, and Eleazar the priest, and unto the congregation of the children of Israel, unto the camp at the plains of Moab, which are by Jordan near Jericho.
NUM|31|13|And Moses, and Eleazar the priest, and all the princes of the congregation, went forth to meet them without the camp.
NUM|31|14|And Moses was wroth with the officers of the host, with the captains over thousands, and captains over hundreds, which came from the battle.
NUM|31|15|And Moses said unto them, Have ye saved all the women alive?
NUM|31|16|Behold, these caused the children of Israel, through the counsel of Balaam, to commit trespass against the LORD in the matter of Peor, and there was a plague among the congregation of the LORD.
NUM|31|17|Now therefore kill every male among the little ones, and kill every woman that hath known man by lying with him.
NUM|31|18|But all the women children, that have not known a man by lying with him, keep alive for yourselves.
NUM|31|19|And do ye abide without the camp seven days: whosoever hath killed any person, and whosoever hath touched any slain, purify both yourselves and your captives on the third day, and on the seventh day.
NUM|31|20|And purify all your raiment, and all that is made of skins, and all work of goats' hair, and all things made of wood.
NUM|31|21|And Eleazar the priest said unto the men of war which went to the battle, This is the ordinance of the law which the LORD commanded Moses;
NUM|31|22|Only the gold, and the silver, the brass, the iron, the tin, and the lead,
NUM|31|23|Every thing that may abide the fire, ye shall make it go through the fire, and it shall be clean: nevertheless it shall be purified with the water of separation: and all that abideth not the fire ye shall make go through the water.
NUM|31|24|And ye shall wash your clothes on the seventh day, and ye shall be clean, and afterward ye shall come into the camp.
NUM|31|25|And the LORD spake unto Moses, saying,
NUM|31|26|Take the sum of the prey that was taken, both of man and of beast, thou, and Eleazar the priest, and the chief fathers of the congregation:
NUM|31|27|And divide the prey into two parts; between them that took the war upon them, who went out to battle, and between all the congregation:
NUM|31|28|And levy a tribute unto the LORD of the men of war which went out to battle: one soul of five hundred, both of the persons, and of the beeves, and of the asses, and of the sheep:
NUM|31|29|Take it of their half, and give it unto Eleazar the priest, for an heave offering of the LORD.
NUM|31|30|And of the children of Israel's half, thou shalt take one portion of fifty, of the persons, of the beeves, of the asses, and of the flocks, of all manner of beasts, and give them unto the Levites, which keep the charge of the tabernacle of the LORD.
NUM|31|31|And Moses and Eleazar the priest did as the LORD commanded Moses.
NUM|31|32|And the booty, being the rest of the prey which the men of war had caught, was six hundred thousand and seventy thousand and five thousand sheep,
NUM|31|33|And threescore and twelve thousand beeves,
NUM|31|34|And threescore and one thousand asses,
NUM|31|35|And thirty and two thousand persons in all, of women that had not known man by lying with him.
NUM|31|36|And the half, which was the portion of them that went out to war, was in number three hundred thousand and seven and thirty thousand and five hundred sheep:
NUM|31|37|And the LORD's tribute of the sheep was six hundred and threescore and fifteen.
NUM|31|38|And the beeves were thirty and six thousand; of which the LORD's tribute was threescore and twelve.
NUM|31|39|And the asses were thirty thousand and five hundred; of which the LORD's tribute was threescore and one.
NUM|31|40|And the persons were sixteen thousand; of which the LORD's tribute was thirty and two persons.
NUM|31|41|And Moses gave the tribute, which was the LORD's heave offering, unto Eleazar the priest, as the LORD commanded Moses.
NUM|31|42|And of the children of Israel's half, which Moses divided from the men that warred,
NUM|31|43|(Now the half that pertained unto the congregation was three hundred thousand and thirty thousand and seven thousand and five hundred sheep,
NUM|31|44|And thirty and six thousand beeves,
NUM|31|45|And thirty thousand asses and five hundred,
NUM|31|46|And sixteen thousand persons;)
NUM|31|47|Even of the children of Israel's half, Moses took one portion of fifty, both of man and of beast, and gave them unto the Levites, which kept the charge of the tabernacle of the LORD; as the LORD commanded Moses.
NUM|31|48|And the officers which were over thousands of the host, the captains of thousands, and captains of hundreds, came near unto Moses:
NUM|31|49|And they said unto Moses, Thy servants have taken the sum of the men of war which are under our charge, and there lacketh not one man of us.
NUM|31|50|We have therefore brought an oblation for the LORD, what every man hath gotten, of jewels of gold, chains, and bracelets, rings, earrings, and tablets, to make an atonement for our souls before the LORD.
NUM|31|51|And Moses and Eleazar the priest took the gold of them, even all wrought jewels.
NUM|31|52|And all the gold of the offering that they offered up to the LORD, of the captains of thousands, and of the captains of hundreds, was sixteen thousand seven hundred and fifty shekels.
NUM|31|53|(For the men of war had taken spoil, every man for himself.)
NUM|31|54|And Moses and Eleazar the priest took the gold of the captains of thousands and of hundreds, and brought it into the tabernacle of the congregation, for a memorial for the children of Israel before the LORD.
NUM|32|1|Now the children of Reuben and the children of Gad had a very great multitude of cattle: and when they saw the land of Jazer, and the land of Gilead, that, behold, the place was a place for cattle;
NUM|32|2|The children of Gad and the children of Reuben came and spake unto Moses, and to Eleazar the priest, and unto the princes of the congregation, saying,
NUM|32|3|Ataroth, and Dibon, and Jazer, and Nimrah, and Heshbon, and Elealeh, and Shebam, and Nebo, and Beon,
NUM|32|4|Even the country which the LORD smote before the congregation of Israel, is a land for cattle, and thy servants have cattle:
NUM|32|5|Wherefore, said they, if we have found grace in thy sight, let this land be given unto thy servants for a possession, and bring us not over Jordan.
NUM|32|6|And Moses said unto the children of Gad and to the children of Reuben, Shall your brethren go to war, and shall ye sit here?
NUM|32|7|And wherefore discourage ye the heart of the children of Israel from going over into the land which the LORD hath given them?
NUM|32|8|Thus did your fathers, when I sent them from Kadeshbarnea to see the land.
NUM|32|9|For when they went up unto the valley of Eshcol, and saw the land, they discouraged the heart of the children of Israel, that they should not go into the land which the LORD had given them.
NUM|32|10|And the LORD's anger was kindled the same time, and he sware, saying,
NUM|32|11|Surely none of the men that came up out of Egypt, from twenty years old and upward, shall see the land which I sware unto Abraham, unto Isaac, and unto Jacob; because they have not wholly followed me:
NUM|32|12|Save Caleb the son of Jephunneh the Kenezite, and Joshua the son of Nun: for they have wholly followed the LORD.
NUM|32|13|And the LORD's anger was kindled against Israel, and he made them wander in the wilderness forty years, until all the generation, that had done evil in the sight of the LORD, was consumed.
NUM|32|14|And, behold, ye are risen up in your fathers' stead, an increase of sinful men, to augment yet the fierce anger of the LORD toward Israel.
NUM|32|15|For if ye turn away from after him, he will yet again leave them in the wilderness; and ye shall destroy all this people.
NUM|32|16|And they came near unto him, and said, We will build sheepfolds here for our cattle, and cities for our little ones:
NUM|32|17|But we ourselves will go ready armed before the children of Israel, until we have brought them unto their place: and our little ones shall dwell in the fenced cities because of the inhabitants of the land.
NUM|32|18|We will not return unto our houses, until the children of Israel have inherited every man his inheritance.
NUM|32|19|For we will not inherit with them on yonder side Jordan, or forward; because our inheritance is fallen to us on this side Jordan eastward.
NUM|32|20|And Moses said unto them, If ye will do this thing, if ye will go armed before the LORD to war,
NUM|32|21|And will go all of you armed over Jordan before the LORD, until he hath driven out his enemies from before him,
NUM|32|22|And the land be subdued before the LORD: then afterward ye shall return, and be guiltless before the LORD, and before Israel; and this land shall be your possession before the LORD.
NUM|32|23|But if ye will not do so, behold, ye have sinned against the LORD: and be sure your sin will find you out.
NUM|32|24|Build you cities for your little ones, and folds for your sheep; and do that which hath proceeded out of your mouth.
NUM|32|25|And the children of Gad and the children of Reuben spake unto Moses, saying, Thy servants will do as my lord commandeth.
NUM|32|26|Our little ones, our wives, our flocks, and all our cattle, shall be there in the cities of Gilead:
NUM|32|27|But thy servants will pass over, every man armed for war, before the Lord to battle, as my lord saith.
NUM|32|28|So concerning them Moses commanded Eleazar the priest, and Joshua the son of Nun, and the chief fathers of the tribes of the children of Israel:
NUM|32|29|And Moses said unto them, If the children of Gad and the children of Reuben will pass with you over Jordan, every man armed to battle, before the LORD, and the land shall be subdued before you; then ye shall give them the land of Gilead for a possession:
NUM|32|30|But if they will not pass over with you armed, they shall have possessions among you in the land of Canaan.
NUM|32|31|And the children of Gad and the children of Reuben answered, saying, As the LORD hath said unto thy servants, so will we do.
NUM|32|32|We will pass over armed before the LORD into the land of Canaan, that the possession of our inheritance on this side Jordan may be ours.
NUM|32|33|And Moses gave unto them, even to the children of Gad, and to the children of Reuben, and unto half the tribe of Manasseh the son of Joseph, the kingdom of Sihon king of the Amorites, and the kingdom of Og king of Bashan, the land, with the cities thereof in the coasts, even the cities of the country round about.
NUM|32|34|And the children of Gad built Dibon, and Ataroth, and Aroer,
NUM|32|35|And Atroth, Shophan, and Jaazer, and Jogbehah,
NUM|32|36|And Bethnimrah, and Bethharan, fenced cities: and folds for sheep.
NUM|32|37|And the children of Reuben built Heshbon, and Elealeh, and Kirjathaim,
NUM|32|38|And Nebo, and Baalmeon, (their names being changed,) and Shibmah: and gave other names unto the cities which they builded.
NUM|32|39|And the children of Machir the son of Manasseh went to Gilead, and took it, and dispossessed the Amorite which was in it.
NUM|32|40|And Moses gave Gilead unto Machir the son of Manasseh; and he dwelt therein.
NUM|32|41|And Jair the son of Manasseh went and took the small towns thereof, and called them Havothjair.
NUM|32|42|And Nobah went and took Kenath, and the villages thereof, and called it Nobah, after his own name.
NUM|33|1|These are the journeys of the children of Israel, which went forth out of the land of Egypt with their armies under the hand of Moses and Aaron.
NUM|33|2|And Moses wrote their goings out according to their journeys by the commandment of the LORD: and these are their journeys according to their goings out.
NUM|33|3|And they departed from Rameses in the first month, on the fifteenth day of the first month; on the morrow after the passover the children of Israel went out with an high hand in the sight of all the Egyptians.
NUM|33|4|For the Egyptians buried all their firstborn, which the LORD had smitten among them: upon their gods also the LORD executed judgments.
NUM|33|5|And the children of Israel removed from Rameses, and pitched in Succoth.
NUM|33|6|And they departed from Succoth, and pitched in Etham, which is in the edge of the wilderness.
NUM|33|7|And they removed from Etham, and turned again unto Pihahiroth, which is before Baalzephon: and they pitched before Migdol.
NUM|33|8|And they departed from before Pihahiroth, and passed through the midst of the sea into the wilderness, and went three days' journey in the wilderness of Etham, and pitched in Marah.
NUM|33|9|And they removed from Marah, and came unto Elim: and in Elim were twelve fountains of water, and threescore and ten palm trees; and they pitched there.
NUM|33|10|And they removed from Elim, and encamped by the Red sea.
NUM|33|11|And they removed from the Red sea, and encamped in the wilderness of Sin.
NUM|33|12|And they took their journey out of the wilderness of Sin, and encamped in Dophkah.
NUM|33|13|And they departed from Dophkah, and encamped in Alush.
NUM|33|14|And they removed from Alush, and encamped at Rephidim, where was no water for the people to drink.
NUM|33|15|And they departed from Rephidim, and pitched in the wilderness of Sinai.
NUM|33|16|And they removed from the desert of Sinai, and pitched at Kibrothhattaavah.
NUM|33|17|And they departed from Kibrothhattaavah, and encamped at Hazeroth.
NUM|33|18|And they departed from Hazeroth, and pitched in Rithmah.
NUM|33|19|And they departed from Rithmah, and pitched at Rimmonparez.
NUM|33|20|And they departed from Rimmonparez, and pitched in Libnah.
NUM|33|21|And they removed from Libnah, and pitched at Rissah.
NUM|33|22|And they journeyed from Rissah, and pitched in Kehelathah.
NUM|33|23|And they went from Kehelathah, and pitched in mount Shapher.
NUM|33|24|And they removed from mount Shapher, and encamped in Haradah.
NUM|33|25|And they removed from Haradah, and pitched in Makheloth.
NUM|33|26|And they removed from Makheloth, and encamped at Tahath.
NUM|33|27|And they departed from Tahath, and pitched at Tarah.
NUM|33|28|And they removed from Tarah, and pitched in Mithcah.
NUM|33|29|And they went from Mithcah, and pitched in Hashmonah.
NUM|33|30|And they departed from Hashmonah, and encamped at Moseroth.
NUM|33|31|And they departed from Moseroth, and pitched in Benejaakan.
NUM|33|32|And they removed from Benejaakan, and encamped at Horhagidgad.
NUM|33|33|And they went from Horhagidgad, and pitched in Jotbathah.
NUM|33|34|And they removed from Jotbathah, and encamped at Ebronah.
NUM|33|35|And they departed from Ebronah, and encamped at Eziongaber.
NUM|33|36|And they removed from Eziongaber, and pitched in the wilderness of Zin, which is Kadesh.
NUM|33|37|And they removed from Kadesh, and pitched in mount Hor, in the edge of the land of Edom.
NUM|33|38|And Aaron the priest went up into mount Hor at the commandment of the LORD, and died there, in the fortieth year after the children of Israel were come out of the land of Egypt, in the first day of the fifth month.
NUM|33|39|And Aaron was an hundred and twenty and three years old when he died in mount Hor.
NUM|33|40|And king Arad the Canaanite, which dwelt in the south in the land of Canaan, heard of the coming of the children of Israel.
NUM|33|41|And they departed from mount Hor, and pitched in Zalmonah.
NUM|33|42|And they departed from Zalmonah, and pitched in Punon.
NUM|33|43|And they departed from Punon, and pitched in Oboth.
NUM|33|44|And they departed from Oboth, and pitched in Ijeabarim, in the border of Moab.
NUM|33|45|And they departed from Iim, and pitched in Dibongad.
NUM|33|46|And they removed from Dibongad, and encamped in Almondiblathaim.
NUM|33|47|And they removed from Almondiblathaim, and pitched in the mountains of Abarim, before Nebo.
NUM|33|48|And they departed from the mountains of Abarim, and pitched in the plains of Moab by Jordan near Jericho.
NUM|33|49|And they pitched by Jordan, from Bethjesimoth even unto Abelshittim in the plains of Moab.
NUM|33|50|And the LORD spake unto Moses in the plains of Moab by Jordan near Jericho, saying,
NUM|33|51|Speak unto the children of Israel, and say unto them, When ye are passed over Jordan into the land of Canaan;
NUM|33|52|Then ye shall drive out all the inhabitants of the land from before you, and destroy all their pictures, and destroy all their molten images, and quite pluck down all their high places:
NUM|33|53|And ye shall dispossess the inhabitants of the land, and dwell therein: for I have given you the land to possess it.
NUM|33|54|And ye shall divide the land by lot for an inheritance among your families: and to the more ye shall give the more inheritance, and to the fewer ye shall give the less inheritance: every man's inheritance shall be in the place where his lot falleth; according to the tribes of your fathers ye shall inherit.
NUM|33|55|But if ye will not drive out the inhabitants of the land from before you; then it shall come to pass, that those which ye let remain of them shall be pricks in your eyes, and thorns in your sides, and shall vex you in the land wherein ye dwell.
NUM|33|56|Moreover it shall come to pass, that I shall do unto you, as I thought to do unto them.
NUM|34|1|And the LORD spake unto Moses, saying,
NUM|34|2|Command the children of Israel, and say unto them, When ye come into the land of Canaan; (this is the land that shall fall unto you for an inheritance, even the land of Canaan with the coasts thereof:)
NUM|34|3|Then your south quarter shall be from the wilderness of Zin along by the coast of Edom, and your south border shall be the outmost coast of the salt sea eastward:
NUM|34|4|And your border shall turn from the south to the ascent of Akrabbim, and pass on to Zin: and the going forth thereof shall be from the south to Kadeshbarnea, and shall go on to Hazaraddar, and pass on to Azmon:
NUM|34|5|And the border shall fetch a compass from Azmon unto the river of Egypt, and the goings out of it shall be at the sea.
NUM|34|6|And as for the western border, ye shall even have the great sea for a border: this shall be your west border.
NUM|34|7|And this shall be your north border: from the great sea ye shall point out for you mount Hor:
NUM|34|8|From mount Hor ye shall point out your border unto the entrance of Hamath; and the goings forth of the border shall be to Zedad:
NUM|34|9|And the border shall go on to Ziphron, and the goings out of it shall be at Hazarenan: this shall be your north border.
NUM|34|10|And ye shall point out your east border from Hazarenan to Shepham:
NUM|34|11|And the coast shall go down from Shepham to Riblah, on the east side of Ain; and the border shall descend, and shall reach unto the side of the sea of Chinnereth eastward:
NUM|34|12|And the border shall go down to Jordan, and the goings out of it shall be at the salt sea: this shall be your land with the coasts thereof round about.
NUM|34|13|And Moses commanded the children of Israel, saying, This is the land which ye shall inherit by lot, which the LORD commanded to give unto the nine tribes, and to the half tribe:
NUM|34|14|For the tribe of the children of Reuben according to the house of their fathers, and the tribe of the children of Gad according to the house of their fathers, have received their inheritance; and half the tribe of Manasseh have received their inheritance:
NUM|34|15|The two tribes and the half tribe have received their inheritance on this side Jordan near Jericho eastward, toward the sunrising.
NUM|34|16|And the LORD spake unto Moses, saying,
NUM|34|17|These are the names of the men which shall divide the land unto you: Eleazar the priest, and Joshua the son of Nun.
NUM|34|18|And ye shall take one prince of every tribe, to divide the land by inheritance.
NUM|34|19|And the names of the men are these: Of the tribe of Judah, Caleb the son of Jephunneh.
NUM|34|20|And of the tribe of the children of Simeon, Shemuel the son of Ammihud.
NUM|34|21|Of the tribe of Benjamin, Elidad the son of Chislon.
NUM|34|22|And the prince of the tribe of the children of Dan, Bukki the son of Jogli.
NUM|34|23|The prince of the children of Joseph, for the tribe of the children of Manasseh, Hanniel the son of Ephod.
NUM|34|24|And the prince of the tribe of the children of Ephraim, Kemuel the son of Shiphtan.
NUM|34|25|And the prince of the tribe of the children of Zebulun, Elizaphan the son of Parnach.
NUM|34|26|And the prince of the tribe of the children of Issachar, Paltiel the son of Azzan.
NUM|34|27|And the prince of the tribe of the children of Asher, Ahihud the son of Shelomi.
NUM|34|28|And the prince of the tribe of the children of Naphtali, Pedahel the son of Ammihud.
NUM|34|29|These are they whom the LORD commanded to divide the inheritance unto the children of Israel in the land of Canaan.
NUM|35|1|And the LORD spake unto Moses in the plains of Moab by Jordan near Jericho, saying,
NUM|35|2|Command the children of Israel, that they give unto the Levites of the inheritance of their possession cities to dwell in; and ye shall give also unto the Levites suburbs for the cities round about them.
NUM|35|3|And the cities shall they have to dwell in; and the suburbs of them shall be for their cattle, and for their goods, and for all their beasts.
NUM|35|4|And the suburbs of the cities, which ye shall give unto the Levites, shall reach from the wall of the city and outward a thousand cubits round about.
NUM|35|5|And ye shall measure from without the city on the east side two thousand cubits, and on the south side two thousand cubits, and on the west side two thousand cubits, and on the north side two thousand cubits; and the city shall be in the midst: this shall be to them the suburbs of the cities.
NUM|35|6|And among the cities which ye shall give unto the Levites there shall be six cities for refuge, which ye shall appoint for the manslayer, that he may flee thither: and to them ye shall add forty and two cities.
NUM|35|7|So all the cities which ye shall give to the Levites shall be forty and eight cities: them shall ye give with their suburbs.
NUM|35|8|And the cities which ye shall give shall be of the possession of the children of Israel: from them that have many ye shall give many; but from them that have few ye shall give few: every one shall give of his cities unto the Levites according to his inheritance which he inheriteth.
NUM|35|9|And the LORD spake unto Moses, saying,
NUM|35|10|Speak unto the children of Israel, and say unto them, When ye be come over Jordan into the land of Canaan;
NUM|35|11|Then ye shall appoint you cities to be cities of refuge for you; that the slayer may flee thither, which killeth any person at unawares.
NUM|35|12|And they shall be unto you cities for refuge from the avenger; that the manslayer die not, until he stand before the congregation in judgment.
NUM|35|13|And of these cities which ye shall give six cities shall ye have for refuge.
NUM|35|14|Ye shall give three cities on this side Jordan, and three cities shall ye give in the land of Canaan, which shall be cities of refuge.
NUM|35|15|These six cities shall be a refuge, both for the children of Israel, and for the stranger, and for the sojourner among them: that every one that killeth any person unawares may flee thither.
NUM|35|16|And if he smite him with an instrument of iron, so that he die, he is a murderer: the murderer shall surely be put to death.
NUM|35|17|And if he smite him with throwing a stone, wherewith he may die, and he die, he is a murderer: the murderer shall surely be put to death.
NUM|35|18|Or if he smite him with an hand weapon of wood, wherewith he may die, and he die, he is a murderer: the murderer shall surely be put to death.
NUM|35|19|The revenger of blood himself shall slay the murderer: when he meeteth him, he shall slay him.
NUM|35|20|But if he thrust him of hatred, or hurl at him by laying of wait, that he die;
NUM|35|21|Or in enmity smite him with his hand, that he die: he that smote him shall surely be put to death; for he is a murderer: the revenger of blood shall slay the murderer, when he meeteth him.
NUM|35|22|But if he thrust him suddenly without enmity, or have cast upon him any thing without laying of wait,
NUM|35|23|Or with any stone, wherewith a man may die, seeing him not, and cast it upon him, that he die, and was not his enemy, neither sought his harm:
NUM|35|24|Then the congregation shall judge between the slayer and the revenger of blood according to these judgments:
NUM|35|25|And the congregation shall deliver the slayer out of the hand of the revenger of blood, and the congregation shall restore him to the city of his refuge, whither he was fled: and he shall abide in it unto the death of the high priest, which was anointed with the holy oil.
NUM|35|26|But if the slayer shall at any time come without the border of the city of his refuge, whither he was fled;
NUM|35|27|And the revenger of blood find him without the borders of the city of his refuge, and the revenger of blood kill the slayer; he shall not be guilty of blood:
NUM|35|28|Because he should have remained in the city of his refuge until the death of the high priest: but after the death of the high priest the slayer shall return into the land of his possession.
NUM|35|29|So these things shall be for a statute of judgment unto you throughout your generations in all your dwellings.
NUM|35|30|Whoso killeth any person, the murderer shall be put to death by the mouth of witnesses: but one witness shall not testify against any person to cause him to die.
NUM|35|31|Moreover ye shall take no satisfaction for the life of a murderer, which is guilty of death: but he shall be surely put to death.
NUM|35|32|And ye shall take no satisfaction for him that is fled to the city of his refuge, that he should come again to dwell in the land, until the death of the priest.
NUM|35|33|So ye shall not pollute the land wherein ye are: for blood it defileth the land: and the land cannot be cleansed of the blood that is shed therein, but by the blood of him that shed it.
NUM|35|34|Defile not therefore the land which ye shall inhabit, wherein I dwell: for I the LORD dwell among the children of Israel.
NUM|36|1|And the chief fathers of the families of the children of Gilead, the son of Machir, the son of Manasseh, of the families of the sons of Joseph, came near, and spake before Moses, and before the princes, the chief fathers of the children of Israel:
NUM|36|2|And they said, The LORD commanded my lord to give the land for an inheritance by lot to the children of Israel: and my lord was commanded by the LORD to give the inheritance of Zelophehad our brother unto his daughters.
NUM|36|3|And if they be married to any of the sons of the other tribes of the children of Israel, then shall their inheritance be taken from the inheritance of our fathers, and shall be put to the inheritance of the tribe whereunto they are received: so shall it be taken from the lot of our inheritance.
NUM|36|4|And when the jubilee of the children of Israel shall be, then shall their inheritance be put unto the inheritance of the tribe whereunto they are received: so shall their inheritance be taken away from the inheritance of the tribe of our fathers.
NUM|36|5|And Moses commanded the children of Israel according to the word of the LORD, saying, The tribe of the sons of Joseph hath said well.
NUM|36|6|This is the thing which the LORD doth command concerning the daughters of Zelophehad, saying, Let them marry to whom they think best; only to the family of the tribe of their father shall they marry.
NUM|36|7|So shall not the inheritance of the children of Israel remove from tribe to tribe: for every one of the children of Israel shall keep himself to the inheritance of the tribe of his fathers.
NUM|36|8|And every daughter, that possesseth an inheritance in any tribe of the children of Israel, shall be wife unto one of the family of the tribe of her father, that the children of Israel may enjoy every man the inheritance of his fathers.
NUM|36|9|Neither shall the inheritance remove from one tribe to another tribe; but every one of the tribes of the children of Israel shall keep himself to his own inheritance.
NUM|36|10|Even as the LORD commanded Moses, so did the daughters of Zelophehad:
NUM|36|11|For Mahlah, Tirzah, and Hoglah, and Milcah, and Noah, the daughters of Zelophehad, were married unto their father's brothers' sons:
NUM|36|12|And they were married into the families of the sons of Manasseh the son of Joseph, and their inheritance remained in the tribe of the family of their father.
NUM|36|13|These are the commandments and the judgments, which the LORD commanded by the hand of Moses unto the children of Israel in the plains of Moab by Jordan near Jericho.
