ESTH|1|1|This is what happened during the time of Xerxes, the Xerxes who ruled over 127 provinces stretching from India to Cush:
ESTH|1|2|At that time King Xerxes reigned from his royal throne in the citadel of Susa,
ESTH|1|3|and in the third year of his reign he gave a banquet for all his nobles and officials. The military leaders of Persia and Media, the princes, and the nobles of the provinces were present.
ESTH|1|4|For a full 180 days he displayed the vast wealth of his kingdom and the splendor and glory of his majesty.
ESTH|1|5|When these days were over, the king gave a banquet, lasting seven days, in the enclosed garden of the king's palace, for all the people from the least to the greatest, who were in the citadel of Susa.
ESTH|1|6|The garden had hangings of white and blue linen, fastened with cords of white linen and purple material to silver rings on marble pillars. There were couches of gold and silver on a mosaic pavement of porphyry, marble, mother-of-pearl and other costly stones.
ESTH|1|7|Wine was served in goblets of gold, each one different from the other, and the royal wine was abundant, in keeping with the king's liberality.
ESTH|1|8|By the king's command each guest was allowed to drink in his own way, for the king instructed all the wine stewards to serve each man what he wished.
ESTH|1|9|Queen Vashti also gave a banquet for the women in the royal palace of King Xerxes.
ESTH|1|10|On the seventh day, when King Xerxes was in high spirits from wine, he commanded the seven eunuchs who served him-Mehuman, Biztha, Harbona, Bigtha, Abagtha, Zethar and Carcas-
ESTH|1|11|to bring before him Queen Vashti, wearing her royal crown, in order to display her beauty to the people and nobles, for she was lovely to look at.
ESTH|1|12|But when the attendants delivered the king's command, Queen Vashti refused to come. Then the king became furious and burned with anger.
ESTH|1|13|Since it was customary for the king to consult experts in matters of law and justice, he spoke with the wise men who understood the times
ESTH|1|14|and were closest to the king-Carshena, Shethar, Admatha, Tarshish, Meres, Marsena and Memucan, the seven nobles of Persia and Media who had special access to the king and were highest in the kingdom.
ESTH|1|15|"According to law, what must be done to Queen Vashti?" he asked. "She has not obeyed the command of King Xerxes that the eunuchs have taken to her."
ESTH|1|16|Then Memucan replied in the presence of the king and the nobles, "Queen Vashti has done wrong, not only against the king but also against all the nobles and the peoples of all the provinces of King Xerxes.
ESTH|1|17|For the queen's conduct will become known to all the women, and so they will despise their husbands and say, 'King Xerxes commanded Queen Vashti to be brought before him, but she would not come.'
ESTH|1|18|This very day the Persian and Median women of the nobility who have heard about the queen's conduct will respond to all the king's nobles in the same way. There will be no end of disrespect and discord.
ESTH|1|19|"Therefore, if it pleases the king, let him issue a royal decree and let it be written in the laws of Persia and Media, which cannot be repealed, that Vashti is never again to enter the presence of King Xerxes. Also let the king give her royal position to someone else who is better than she.
ESTH|1|20|Then when the king's edict is proclaimed throughout all his vast realm, all the women will respect their husbands, from the least to the greatest."
ESTH|1|21|The king and his nobles were pleased with this advice, so the king did as Memucan proposed.
ESTH|1|22|He sent dispatches to all parts of the kingdom, to each province in its own script and to each people in its own language, proclaiming in each people's tongue that every man should be ruler over his own household.
ESTH|2|1|Later when the anger of King Xerxes had subsided, he remembered Vashti and what she had done and what he had decreed about her.
ESTH|2|2|Then the king's personal attendants proposed, "Let a search be made for beautiful young virgins for the king.
ESTH|2|3|Let the king appoint commissioners in every province of his realm to bring all these beautiful girls into the harem at the citadel of Susa. Let them be placed under the care of Hegai, the king's eunuch, who is in charge of the women; and let beauty treatments be given to them.
ESTH|2|4|Then let the girl who pleases the king be queen instead of Vashti." This advice appealed to the king, and he followed it.
ESTH|2|5|Now there was in the citadel of Susa a Jew of the tribe of Benjamin, named Mordecai son of Jair, the son of Shimei, the son of Kish,
ESTH|2|6|who had been carried into exile from Jerusalem by Nebuchadnezzar king of Babylon, among those taken captive with Jehoiachin king of Judah.
ESTH|2|7|Mordecai had a cousin named Hadassah, whom he had brought up because she had neither father nor mother. This girl, who was also known as Esther, was lovely in form and features, and Mordecai had taken her as his own daughter when her father and mother died.
ESTH|2|8|When the king's order and edict had been proclaimed, many girls were brought to the citadel of Susa and put under the care of Hegai. Esther also was taken to the king's palace and entrusted to Hegai, who had charge of the harem.
ESTH|2|9|The girl pleased him and won his favor. Immediately he provided her with her beauty treatments and special food. He assigned to her seven maids selected from the king's palace and moved her and her maids into the best place in the harem.
ESTH|2|10|Esther had not revealed her nationality and family background, because Mordecai had forbidden her to do so.
ESTH|2|11|Every day he walked back and forth near the courtyard of the harem to find out how Esther was and what was happening to her.
ESTH|2|12|Before a girl's turn came to go in to King Xerxes, she had to complete twelve months of beauty treatments prescribed for the women, six months with oil of myrrh and six with perfumes and cosmetics.
ESTH|2|13|And this is how she would go to the king: Anything she wanted was given her to take with her from the harem to the king's palace.
ESTH|2|14|In the evening she would go there and in the morning return to another part of the harem to the care of Shaashgaz, the king's eunuch who was in charge of the concubines. She would not return to the king unless he was pleased with her and summoned her by name.
ESTH|2|15|When the turn came for Esther (the girl Mordecai had adopted, the daughter of his uncle Abihail) to go to the king, she asked for nothing other than what Hegai, the king's eunuch who was in charge of the harem, suggested. And Esther won the favor of everyone who saw her.
ESTH|2|16|She was taken to King Xerxes in the royal residence in the tenth month, the month of Tebeth, in the seventh year of his reign.
ESTH|2|17|Now the king was attracted to Esther more than to any of the other women, and she won his favor and approval more than any of the other virgins. So he set a royal crown on her head and made her queen instead of Vashti.
ESTH|2|18|And the king gave a great banquet, Esther's banquet, for all his nobles and officials. He proclaimed a holiday throughout the provinces and distributed gifts with royal liberality.
ESTH|2|19|When the virgins were assembled a second time, Mordecai was sitting at the king's gate.
ESTH|2|20|But Esther had kept secret her family background and nationality just as Mordecai had told her to do, for she continued to follow Mordecai's instructions as she had done when he was bringing her up.
ESTH|2|21|During the time Mordecai was sitting at the king's gate, Bigthana and Teresh, two of the king's officers who guarded the doorway, became angry and conspired to assassinate King Xerxes.
ESTH|2|22|But Mordecai found out about the plot and told Queen Esther, who in turn reported it to the king, giving credit to Mordecai.
ESTH|2|23|And when the report was investigated and found to be true, the two officials were hanged on a gallows. All this was recorded in the book of the annals in the presence of the king.
ESTH|3|1|After these events, King Xerxes honored Haman son of Hammedatha, the Agagite, elevating him and giving him a seat of honor higher than that of all the other nobles.
ESTH|3|2|All the royal officials at the king's gate knelt down and paid honor to Haman, for the king had commanded this concerning him. But Mordecai would not kneel down or pay him honor.
ESTH|3|3|Then the royal officials at the king's gate asked Mordecai, "Why do you disobey the king's command?"
ESTH|3|4|Day after day they spoke to him but he refused to comply. Therefore they told Haman about it to see whether Mordecai's behavior would be tolerated, for he had told them he was a Jew.
ESTH|3|5|When Haman saw that Mordecai would not kneel down or pay him honor, he was enraged.
ESTH|3|6|Yet having learned who Mordecai's people were, he scorned the idea of killing only Mordecai. Instead Haman looked for a way to destroy all Mordecai's people, the Jews, throughout the whole kingdom of Xerxes.
ESTH|3|7|In the twelfth year of King Xerxes, in the first month, the month of Nisan, they cast the pur (that is, the lot) in the presence of Haman to select a day and month. And the lot fell on the twelfth month, the month of Adar.
ESTH|3|8|Then Haman said to King Xerxes, "There is a certain people dispersed and scattered among the peoples in all the provinces of your kingdom whose customs are different from those of all other people and who do not obey the king's laws; it is not in the king's best interest to tolerate them.
ESTH|3|9|If it pleases the king, let a decree be issued to destroy them, and I will put ten thousand talents of silver into the royal treasury for the men who carry out this business."
ESTH|3|10|So the king took his signet ring from his finger and gave it to Haman son of Hammedatha, the Agagite, the enemy of the Jews.
ESTH|3|11|"Keep the money," the king said to Haman, "and do with the people as you please."
ESTH|3|12|Then on the thirteenth day of the first month the royal secretaries were summoned. They wrote out in the script of each province and in the language of each people all Haman's orders to the king's satraps, the governors of the various provinces and the nobles of the various peoples. These were written in the name of King Xerxes himself and sealed with his own ring.
ESTH|3|13|Dispatches were sent by couriers to all the king's provinces with the order to destroy, kill and annihilate all the Jews-young and old, women and little children-on a single day, the thirteenth day of the twelfth month, the month of Adar, and to plunder their goods.
ESTH|3|14|A copy of the text of the edict was to be issued as law in every province and made known to the people of every nationality so they would be ready for that day.
ESTH|3|15|Spurred on by the king's command, the couriers went out, and the edict was issued in the citadel of Susa. The king and Haman sat down to drink, but the city of Susa was bewildered.
ESTH|4|1|When Mordecai learned of all that had been done, he tore his clothes, put on sackcloth and ashes, and went out into the city, wailing loudly and bitterly.
ESTH|4|2|But he went only as far as the king's gate, because no one clothed in sackcloth was allowed to enter it.
ESTH|4|3|In every province to which the edict and order of the king came, there was great mourning among the Jews, with fasting, weeping and wailing. Many lay in sackcloth and ashes.
ESTH|4|4|When Esther's maids and eunuchs came and told her about Mordecai, she was in great distress. She sent clothes for him to put on instead of his sackcloth, but he would not accept them.
ESTH|4|5|Then Esther summoned Hathach, one of the king's eunuchs assigned to attend her, and ordered him to find out what was troubling Mordecai and why.
ESTH|4|6|So Hathach went out to Mordecai in the open square of the city in front of the king's gate.
ESTH|4|7|Mordecai told him everything that had happened to him, including the exact amount of money Haman had promised to pay into the royal treasury for the destruction of the Jews.
ESTH|4|8|He also gave him a copy of the text of the edict for their annihilation, which had been published in Susa, to show to Esther and explain it to her, and he told him to urge her to go into the king's presence to beg for mercy and plead with him for her people.
ESTH|4|9|Hathach went back and reported to Esther what Mordecai had said.
ESTH|4|10|Then she instructed him to say to Mordecai,
ESTH|4|11|"All the king's officials and the people of the royal provinces know that for any man or woman who approaches the king in the inner court without being summoned the king has but one law: that he be put to death. The only exception to this is for the king to extend the gold scepter to him and spare his life. But thirty days have passed since I was called to go to the king."
ESTH|4|12|When Esther's words were reported to Mordecai,
ESTH|4|13|he sent back this answer: "Do not think that because you are in the king's house you alone of all the Jews will escape.
ESTH|4|14|For if you remain silent at this time, relief and deliverance for the Jews will arise from another place, but you and your father's family will perish. And who knows but that you have come to royal position for such a time as this?"
ESTH|4|15|Then Esther sent this reply to Mordecai:
ESTH|4|16|"Go, gather together all the Jews who are in Susa, and fast for me. Do not eat or drink for three days, night or day. I and my maids will fast as you do. When this is done, I will go to the king, even though it is against the law. And if I perish, I perish."
ESTH|4|17|So Mordecai went away and carried out all of Esther's instructions.
ESTH|5|1|On the third day Esther put on her royal robes and stood in the inner court of the palace, in front of the king's hall. The king was sitting on his royal throne in the hall, facing the entrance.
ESTH|5|2|When he saw Queen Esther standing in the court, he was pleased with her and held out to her the gold scepter that was in his hand. So Esther approached and touched the tip of the scepter.
ESTH|5|3|Then the king asked, "What is it, Queen Esther? What is your request? Even up to half the kingdom, it will be given you."
ESTH|5|4|"If it pleases the king," replied Esther, "let the king, together with Haman, come today to a banquet I have prepared for him."
ESTH|5|5|"Bring Haman at once," the king said, "so that we may do what Esther asks." So the king and Haman went to the banquet Esther had prepared.
ESTH|5|6|As they were drinking wine, the king again asked Esther, "Now what is your petition? It will be given you. And what is your request? Even up to half the kingdom, it will be granted."
ESTH|5|7|Esther replied, "My petition and my request is this:
ESTH|5|8|If the king regards me with favor and if it pleases the king to grant my petition and fulfill my request, let the king and Haman come tomorrow to the banquet I will prepare for them. Then I will answer the king's question."
ESTH|5|9|Haman went out that day happy and in high spirits. But when he saw Mordecai at the king's gate and observed that he neither rose nor showed fear in his presence, he was filled with rage against Mordecai.
ESTH|5|10|Nevertheless, Haman restrained himself and went home. Calling together his friends and Zeresh, his wife,
ESTH|5|11|Haman boasted to them about his vast wealth, his many sons, and all the ways the king had honored him and how he had elevated him above the other nobles and officials.
ESTH|5|12|"And that's not all," Haman added. "I'm the only person Queen Esther invited to accompany the king to the banquet she gave. And she has invited me along with the king tomorrow.
ESTH|5|13|But all this gives me no satisfaction as long as I see that Jew Mordecai sitting at the king's gate."
ESTH|5|14|His wife Zeresh and all his friends said to him, "Have a gallows built, seventy-five feet high, and ask the king in the morning to have Mordecai hanged on it. Then go with the king to the dinner and be happy." This suggestion delighted Haman, and he had the gallows built.
ESTH|6|1|That night the king could not sleep; so he ordered the book of the chronicles, the record of his reign, to be brought in and read to him.
ESTH|6|2|It was found recorded there that Mordecai had exposed Bigthana and Teresh, two of the king's officers who guarded the doorway, who had conspired to assassinate King Xerxes.
ESTH|6|3|"What honor and recognition has Mordecai received for this?" the king asked. "Nothing has been done for him," his attendants answered.
ESTH|6|4|The king said, "Who is in the court?" Now Haman had just entered the outer court of the palace to speak to the king about hanging Mordecai on the gallows he had erected for him.
ESTH|6|5|His attendants answered, "Haman is standing in the court.Bring him in," the king ordered.
ESTH|6|6|When Haman entered, the king asked him, "What should be done for the man the king delights to honor?" Now Haman thought to himself, "Who is there that the king would rather honor than me?"
ESTH|6|7|So he answered the king, "For the man the king delights to honor,
ESTH|6|8|have them bring a royal robe the king has worn and a horse the king has ridden, one with a royal crest placed on its head.
ESTH|6|9|Then let the robe and horse be entrusted to one of the king's most noble princes. Let them robe the man the king delights to honor, and lead him on the horse through the city streets, proclaiming before him, 'This is what is done for the man the king delights to honor!'"
ESTH|6|10|"Go at once," the king commanded Haman. "Get the robe and the horse and do just as you have suggested for Mordecai the Jew, who sits at the king's gate. Do not neglect anything you have recommended."
ESTH|6|11|So Haman got the robe and the horse. He robed Mordecai, and led him on horseback through the city streets, proclaiming before him, "This is what is done for the man the king delights to honor!"
ESTH|6|12|Afterward Mordecai returned to the king's gate. But Haman rushed home, with his head covered in grief,
ESTH|6|13|and told Zeresh his wife and all his friends everything that had happened to him. His advisers and his wife Zeresh said to him, "Since Mordecai, before whom your downfall has started, is of Jewish origin, you cannot stand against him-you will surely come to ruin!"
ESTH|6|14|While they were still talking with him, the king's eunuchs arrived and hurried Haman away to the banquet Esther had prepared.
ESTH|7|1|So the king and Haman went to dine with Queen Esther,
ESTH|7|2|and as they were drinking wine on that second day, the king again asked, "Queen Esther, what is your petition? It will be given you. What is your request? Even up to half the kingdom, it will be granted."
ESTH|7|3|Then Queen Esther answered, "If I have found favor with you, O king, and if it pleases your majesty, grant me my life-this is my petition. And spare my people-this is my request.
ESTH|7|4|For I and my people have been sold for destruction and slaughter and annihilation. If we had merely been sold as male and female slaves, I would have kept quiet, because no such distress would justify disturbing the king. "
ESTH|7|5|King Xerxes asked Queen Esther, "Who is he? Where is the man who has dared to do such a thing?"
ESTH|7|6|Esther said, "The adversary and enemy is this vile Haman." Then Haman was terrified before the king and queen.
ESTH|7|7|The king got up in a rage, left his wine and went out into the palace garden. But Haman, realizing that the king had already decided his fate, stayed behind to beg Queen Esther for his life.
ESTH|7|8|Just as the king returned from the palace garden to the banquet hall, Haman was falling on the couch where Esther was reclining. The king exclaimed, "Will he even molest the queen while she is with me in the house?" As soon as the word left the king's mouth, they covered Haman's face.
ESTH|7|9|Then Harbona, one of the eunuchs attending the king, said, "A gallows seventy-five feet high stands by Haman's house. He had it made for Mordecai, who spoke up to help the king." The king said, "Hang him on it!"
ESTH|7|10|So they hanged Haman on the gallows he had prepared for Mordecai. Then the king's fury subsided.
ESTH|8|1|That same day King Xerxes gave Queen Esther the estate of Haman, the enemy of the Jews. And Mordecai came into the presence of the king, for Esther had told how he was related to her.
ESTH|8|2|The king took off his signet ring, which he had reclaimed from Haman, and presented it to Mordecai. And Esther appointed him over Haman's estate.
ESTH|8|3|Esther again pleaded with the king, falling at his feet and weeping. She begged him to put an end to the evil plan of Haman the Agagite, which he had devised against the Jews.
ESTH|8|4|Then the king extended the gold scepter to Esther and she arose and stood before him.
ESTH|8|5|"If it pleases the king," she said, "and if he regards me with favor and thinks it the right thing to do, and if he is pleased with me, let an order be written overruling the dispatches that Haman son of Hammedatha, the Agagite, devised and wrote to destroy the Jews in all the king's provinces.
ESTH|8|6|For how can I bear to see disaster fall on my people? How can I bear to see the destruction of my family?"
ESTH|8|7|King Xerxes replied to Queen Esther and to Mordecai the Jew, "Because Haman attacked the Jews, I have given his estate to Esther, and they have hanged him on the gallows.
ESTH|8|8|Now write another decree in the king's name in behalf of the Jews as seems best to you, and seal it with the king's signet ring-for no document written in the king's name and sealed with his ring can be revoked."
ESTH|8|9|At once the royal secretaries were summoned-on the twenty-third day of the third month, the month of Sivan. They wrote out all Mordecai's orders to the Jews, and to the satraps, governors and nobles of the 127 provinces stretching from India to Cush. These orders were written in the script of each province and the language of each people and also to the Jews in their own script and language.
ESTH|8|10|Mordecai wrote in the name of King Xerxes, sealed the dispatches with the king's signet ring, and sent them by mounted couriers, who rode fast horses especially bred for the king.
ESTH|8|11|The king's edict granted the Jews in every city the right to assemble and protect themselves; to destroy, kill and annihilate any armed force of any nationality or province that might attack them and their women and children; and to plunder the property of their enemies.
ESTH|8|12|The day appointed for the Jews to do this in all the provinces of King Xerxes was the thirteenth day of the twelfth month, the month of Adar.
ESTH|8|13|A copy of the text of the edict was to be issued as law in every province and made known to the people of every nationality so that the Jews would be ready on that day to avenge themselves on their enemies.
ESTH|8|14|The couriers, riding the royal horses, raced out, spurred on by the king's command. And the edict was also issued in the citadel of Susa.
ESTH|8|15|Mordecai left the king's presence wearing royal garments of blue and white, a large crown of gold and a purple robe of fine linen. And the city of Susa held a joyous celebration.
ESTH|8|16|For the Jews it was a time of happiness and joy, gladness and honor.
ESTH|8|17|In every province and in every city, wherever the edict of the king went, there was joy and gladness among the Jews, with feasting and celebrating. And many people of other nationalities became Jews because fear of the Jews had seized them.
ESTH|9|1|On the thirteenth day of the twelfth month, the month of Adar, the edict commanded by the king was to be carried out. On this day the enemies of the Jews had hoped to overpower them, but now the tables were turned and the Jews got the upper hand over those who hated them.
ESTH|9|2|The Jews assembled in their cities in all the provinces of King Xerxes to attack those seeking their destruction. No one could stand against them, because the people of all the other nationalities were afraid of them.
ESTH|9|3|And all the nobles of the provinces, the satraps, the governors and the king's administrators helped the Jews, because fear of Mordecai had seized them.
ESTH|9|4|Mordecai was prominent in the palace; his reputation spread throughout the provinces, and he became more and more powerful.
ESTH|9|5|The Jews struck down all their enemies with the sword, killing and destroying them, and they did what they pleased to those who hated them.
ESTH|9|6|In the citadel of Susa, the Jews killed and destroyed five hundred men.
ESTH|9|7|They also killed Parshandatha, Dalphon, Aspatha,
ESTH|9|8|Poratha, Adalia, Aridatha,
ESTH|9|9|Parmashta, Arisai, Aridai and Vaizatha,
ESTH|9|10|the ten sons of Haman son of Hammedatha, the enemy of the Jews. But they did not lay their hands on the plunder.
ESTH|9|11|The number of those slain in the citadel of Susa was reported to the king that same day.
ESTH|9|12|The king said to Queen Esther, "The Jews have killed and destroyed five hundred men and the ten sons of Haman in the citadel of Susa. What have they done in the rest of the king's provinces? Now what is your petition? It will be given you. What is your request? It will also be granted."
ESTH|9|13|"If it pleases the king," Esther answered, "give the Jews in Susa permission to carry out this day's edict tomorrow also, and let Haman's ten sons be hanged on gallows."
ESTH|9|14|So the king commanded that this be done. An edict was issued in Susa, and they hanged the ten sons of Haman.
ESTH|9|15|The Jews in Susa came together on the fourteenth day of the month of Adar, and they put to death in Susa three hundred men, but they did not lay their hands on the plunder.
ESTH|9|16|Meanwhile, the remainder of the Jews who were in the king's provinces also assembled to protect themselves and get relief from their enemies. They killed seventy-five thousand of them but did not lay their hands on the plunder.
ESTH|9|17|This happened on the thirteenth day of the month of Adar, and on the fourteenth they rested and made it a day of feasting and joy.
ESTH|9|18|The Jews in Susa, however, had assembled on the thirteenth and fourteenth, and then on the fifteenth they rested and made it a day of feasting and joy.
ESTH|9|19|That is why rural Jews-those living in villages-observe the fourteenth of the month of Adar as a day of joy and feasting, a day for giving presents to each other.
ESTH|9|20|Mordecai recorded these events, and he sent letters to all the Jews throughout the provinces of King Xerxes, near and far,
ESTH|9|21|to have them celebrate annually the fourteenth and fifteenth days of the month of Adar
ESTH|9|22|as the time when the Jews got relief from their enemies, and as the month when their sorrow was turned into joy and their mourning into a day of celebration. He wrote them to observe the days as days of feasting and joy and giving presents of food to one another and gifts to the poor.
ESTH|9|23|So the Jews agreed to continue the celebration they had begun, doing what Mordecai had written to them.
ESTH|9|24|For Haman son of Hammedatha, the Agagite, the enemy of all the Jews, had plotted against the Jews to destroy them and had cast the pur (that is, the lot) for their ruin and destruction.
ESTH|9|25|But when the plot came to the king's attention, he issued written orders that the evil scheme Haman had devised against the Jews should come back onto his own head, and that he and his sons should be hanged on the gallows.
ESTH|9|26|(Therefore these days were called Purim, from the word pur.) Because of everything written in this letter and because of what they had seen and what had happened to them,
ESTH|9|27|the Jews took it upon themselves to establish the custom that they and their descendants and all who join them should without fail observe these two days every year, in the way prescribed and at the time appointed.
ESTH|9|28|These days should be remembered and observed in every generation by every family, and in every province and in every city. And these days of Purim should never cease to be celebrated by the Jews, nor should the memory of them die out among their descendants.
ESTH|9|29|So Queen Esther, daughter of Abihail, along with Mordecai the Jew, wrote with full authority to confirm this second letter concerning Purim.
ESTH|9|30|And Mordecai sent letters to all the Jews in the 127 provinces of the kingdom of Xerxes-words of goodwill and assurance-
ESTH|9|31|to establish these days of Purim at their designated times, as Mordecai the Jew and Queen Esther had decreed for them, and as they had established for themselves and their descendants in regard to their times of fasting and lamentation.
ESTH|9|32|Esther's decree confirmed these regulations about Purim, and it was written down in the records.
ESTH|10|1|King Xerxes imposed tribute throughout the empire, to its distant shores.
ESTH|10|2|And all his acts of power and might, together with a full account of the greatness of Mordecai to which the king had raised him, are they not written in the book of the annals of the kings of Media and Persia?
ESTH|10|3|Mordecai the Jew was second in rank to King Xerxes, preeminent among the Jews, and held in high esteem by his many fellow Jews, because he worked for the good of his people and spoke up for the welfare of all the Jews.
