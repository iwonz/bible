JAS|1|1|James, a servant of God and of the Lord Jesus Christ, To the twelve tribes scattered among the nations: Greetings.
JAS|1|2|Consider it pure joy, my brothers, whenever you face trials of many kinds,
JAS|1|3|because you know that the testing of your faith develops perseverance.
JAS|1|4|Perseverance must finish its work so that you may be mature and complete, not lacking anything.
JAS|1|5|If any of you lacks wisdom, he should ask God, who gives generously to all without finding fault, and it will be given to him.
JAS|1|6|But when he asks, he must believe and not doubt, because he who doubts is like a wave of the sea, blown and tossed by the wind.
JAS|1|7|That man should not think he will receive anything from the Lord;
JAS|1|8|he is a double-minded man, unstable in all he does.
JAS|1|9|The brother in humble circumstances ought to take pride in his high position.
JAS|1|10|But the one who is rich should take pride in his low position, because he will pass away like a wild flower.
JAS|1|11|For the sun rises with scorching heat and withers the plant; its blossom falls and its beauty is destroyed. In the same way, the rich man will fade away even while he goes about his business.
JAS|1|12|Blessed is the man who perseveres under trial, because when he has stood the test, he will receive the crown of life that God has promised to those who love him.
JAS|1|13|When tempted, no one should say, "God is tempting me." For God cannot be tempted by evil, nor does he tempt anyone;
JAS|1|14|but each one is tempted when, by his own evil desire, he is dragged away and enticed.
JAS|1|15|Then, after desire has conceived, it gives birth to sin; and sin, when it is full-grown, gives birth to death.
JAS|1|16|Don't be deceived, my dear brothers.
JAS|1|17|Every good and perfect gift is from above, coming down from the Father of the heavenly lights, who does not change like shifting shadows.
JAS|1|18|He chose to give us birth through the word of truth, that we might be a kind of firstfruits of all he created.
JAS|1|19|My dear brothers, take note of this: Everyone should be quick to listen, slow to speak and slow to become angry,
JAS|1|20|for man's anger does not bring about the righteous life that God desires.
JAS|1|21|Therefore, get rid of all moral filth and the evil that is so prevalent and humbly accept the word planted in you, which can save you.
JAS|1|22|Do not merely listen to the word, and so deceive yourselves. Do what it says.
JAS|1|23|Anyone who listens to the word but does not do what it says is like a man who looks at his face in a mirror
JAS|1|24|and, after looking at himself, goes away and immediately forgets what he looks like.
JAS|1|25|But the man who looks intently into the perfect law that gives freedom, and continues to do this, not forgetting what he has heard, but doing it--he will be blessed in what he does.
JAS|1|26|If anyone considers himself religious and yet does not keep a tight rein on his tongue, he deceives himself and his religion is worthless.
JAS|1|27|Religion that God our Father accepts as pure and faultless is this: to look after orphans and widows in their distress and to keep oneself from being polluted by the world.
JAS|2|1|My brothers, as believers in our glorious Lord Jesus Christ, don't show favoritism.
JAS|2|2|Suppose a man comes into your meeting wearing a gold ring and fine clothes, and a poor man in shabby clothes also comes in.
JAS|2|3|If you show special attention to the man wearing fine clothes and say, "Here's a good seat for you," but say to the poor man, "You stand there" or "Sit on the floor by my feet,"
JAS|2|4|have you not discriminated among yourselves and become judges with evil thoughts?
JAS|2|5|Listen, my dear brothers: Has not God chosen those who are poor in the eyes of the world to be rich in faith and to inherit the kingdom he promised those who love him?
JAS|2|6|But you have insulted the poor. Is it not the rich who are exploiting you? Are they not the ones who are dragging you into court?
JAS|2|7|Are they not the ones who are slandering the noble name of him to whom you belong?
JAS|2|8|If you really keep the royal law found in Scripture, "Love your neighbor as yourself," you are doing right.
JAS|2|9|But if you show favoritism, you sin and are convicted by the law as lawbreakers.
JAS|2|10|For whoever keeps the whole law and yet stumbles at just one point is guilty of breaking all of it.
JAS|2|11|For he who said, "Do not commit adultery," also said, "Do not murder." If you do not commit adultery but do commit murder, you have become a lawbreaker.
JAS|2|12|Speak and act as those who are going to be judged by the law that gives freedom,
JAS|2|13|because judgment without mercy will be shown to anyone who has not been merciful. Mercy triumphs over judgment!
JAS|2|14|What good is it, my brothers, if a man claims to have faith but has no deeds? Can such faith save him?
JAS|2|15|Suppose a brother or sister is without clothes and daily food.
JAS|2|16|If one of you says to him, "Go, I wish you well; keep warm and well fed," but does nothing about his physical needs, what good is it?
JAS|2|17|In the same way, faith by itself, if it is not accompanied by action, is dead.
JAS|2|18|But someone will say, "You have faith; I have deeds." Show me your faith without deeds, and I will show you my faith by what I do.
JAS|2|19|You believe that there is one God. Good! Even the demons believe that--and shudder.
JAS|2|20|You foolish man, do you want evidence that faith without deeds is useless?
JAS|2|21|Was not our ancestor Abraham considered righteous for what he did when he offered his son Isaac on the altar?
JAS|2|22|You see that his faith and his actions were working together, and his faith was made complete by what he did.
JAS|2|23|And the scripture was fulfilled that says, "Abraham believed God, and it was credited to him as righteousness," and he was called God's friend.
JAS|2|24|You see that a person is justified by what he does and not by faith alone.
JAS|2|25|In the same way, was not even Rahab the prostitute considered righteous for what she did when she gave lodging to the spies and sent them off in a different direction?
JAS|2|26|As the body without the spirit is dead, so faith without deeds is dead.
JAS|3|1|Not many of you should presume to be teachers, my brothers, because you know that we who teach will be judged more strictly.
JAS|3|2|We all stumble in many ways. If anyone is never at fault in what he says, he is a perfect man, able to keep his whole body in check.
JAS|3|3|When we put bits into the mouths of horses to make them obey us, we can turn the whole animal.
JAS|3|4|Or take ships as an example. Although they are so large and are driven by strong winds, they are steered by a very small rudder wherever the pilot wants to go.
JAS|3|5|Likewise the tongue is a small part of the body, but it makes great boasts. Consider what a great forest is set on fire by a small spark.
JAS|3|6|The tongue also is a fire, a world of evil among the parts of the body. It corrupts the whole person, sets the whole course of his life on fire, and is itself set on fire by hell.
JAS|3|7|All kinds of animals, birds, reptiles and creatures of the sea are being tamed and have been tamed by man,
JAS|3|8|but no man can tame the tongue. It is a restless evil, full of deadly poison.
JAS|3|9|With the tongue we praise our Lord and Father, and with it we curse men, who have been made in God's likeness.
JAS|3|10|Out of the same mouth come praise and cursing. My brothers, this should not be.
JAS|3|11|Can both fresh water and salt water flow from the same spring?
JAS|3|12|My brothers, can a fig tree bear olives, or a grapevine bear figs? Neither can a salt spring produce fresh water.
JAS|3|13|Who is wise and understanding among you? Let him show it by his good life, by deeds done in the humility that comes from wisdom.
JAS|3|14|But if you harbor bitter envy and selfish ambition in your hearts, do not boast about it or deny the truth.
JAS|3|15|Such "wisdom" does not come down from heaven but is earthly, unspiritual, of the devil.
JAS|3|16|For where you have envy and selfish ambition, there you find disorder and every evil practice.
JAS|3|17|But the wisdom that comes from heaven is first of all pure; then peace-loving, considerate, submissive, full of mercy and good fruit, impartial and sincere.
JAS|3|18|Peacemakers who sow in peace raise a harvest of righteousness.
JAS|4|1|What causes fights and quarrels among you? Don't they come from your desires that battle within you?
JAS|4|2|You want something but don't get it. You kill and covet, but you cannot have what you want. You quarrel and fight. You do not have, because you do not ask God.
JAS|4|3|When you ask, you do not receive, because you ask with wrong motives, that you may spend what you get on your pleasures.
JAS|4|4|You adulterous people, don't you know that friendship with the world is hatred toward God? Anyone who chooses to be a friend of the world becomes an enemy of God.
JAS|4|5|Or do you think Scripture says without reason that the spirit he caused to live in us envies intensely?
JAS|4|6|But he gives us more grace. That is why Scripture says: "God opposes the proud but gives grace to the humble."
JAS|4|7|Submit yourselves, then, to God. Resist the devil, and he will flee from you.
JAS|4|8|Come near to God and he will come near to you. Wash your hands, you sinners, and purify your hearts, you double-minded.
JAS|4|9|Grieve, mourn and wail. Change your laughter to mourning and your joy to gloom.
JAS|4|10|Humble yourselves before the Lord, and he will lift you up.
JAS|4|11|Brothers, do not slander one another. Anyone who speaks against his brother or judges him speaks against the law and judges it. When you judge the law, you are not keeping it, but sitting in judgment on it.
JAS|4|12|There is only one Lawgiver and Judge, the one who is able to save and destroy. But you--who are you to judge your neighbor?
JAS|4|13|Now listen, you who say, "Today or tomorrow we will go to this or that city, spend a year there, carry on business and make money."
JAS|4|14|Why, you do not even know what will happen tomorrow. What is your life? You are a mist that appears for a little while and then vanishes.
JAS|4|15|Instead, you ought to say, "If it is the Lord's will, we will live and do this or that."
JAS|4|16|As it is, you boast and brag. All such boasting is evil.
JAS|4|17|Anyone, then, who knows the good he ought to do and doesn't do it, sins.
JAS|5|1|Now listen, you rich people, weep and wail because of the misery that is coming upon you.
JAS|5|2|Your wealth has rotted, and moths have eaten your clothes.
JAS|5|3|Your gold and silver are corroded. Their corrosion will testify against you and eat your flesh like fire. You have hoarded wealth in the last days.
JAS|5|4|Look! The wages you failed to pay the workmen who mowed your fields are crying out against you. The cries of the harvesters have reached the ears of the Lord Almighty.
JAS|5|5|You have lived on earth in luxury and self-indulgence. You have fattened yourselves in the day of slaughter.
JAS|5|6|You have condemned and murdered innocent men, who were not opposing you.
JAS|5|7|Be patient, then, brothers, until the Lord's coming. See how the farmer waits for the land to yield its valuable crop and how patient he is for the autumn and spring rains.
JAS|5|8|You too, be patient and stand firm, because the Lord's coming is near.
JAS|5|9|Don't grumble against each other, brothers, or you will be judged. The Judge is standing at the door!
JAS|5|10|Brothers, as an example of patience in the face of suffering, take the prophets who spoke in the name of the Lord.
JAS|5|11|As you know, we consider blessed those who have persevered. You have heard of Job's perseverance and have seen what the Lord finally brought about. The Lord is full of compassion and mercy.
JAS|5|12|Above all, my brothers, do not swear--not by heaven or by earth or by anything else. Let your "Yes" be yes, and your "No," no, or you will be condemned.
JAS|5|13|Is any one of you in trouble? He should pray. Is anyone happy? Let him sing songs of praise.
JAS|5|14|Is any one of you sick? He should call the elders of the church to pray over him and anoint him with oil in the name of the Lord.
JAS|5|15|And the prayer offered in faith will make the sick person well; the Lord will raise him up. If he has sinned, he will be forgiven.
JAS|5|16|Therefore confess your sins to each other and pray for each other so that you may be healed. The prayer of a righteous man is powerful and effective.
JAS|5|17|Elijah was a man just like us. He prayed earnestly that it would not rain, and it did not rain on the land for three and a half years.
JAS|5|18|Again he prayed, and the heavens gave rain, and the earth produced its crops.
JAS|5|19|My brothers, if one of you should wander from the truth and someone should bring him back,
JAS|5|20|remember this: Whoever turns a sinner from the error of his way will save him from death and cover over a multitude of sins.
