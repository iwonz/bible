LAM|1|1|唉！先前人口稠密的城市， 現在為何獨坐！ 先前在列國中為大的， 現在竟如寡婦！ 先前在各省中為王后的， 現在竟成為服苦役的人！
LAM|1|2|她 夜間痛哭，淚流滿頰， 在所有親愛的人中，找不到一個安慰她的。 她的朋友都以詭詐待她， 成為她的仇敵。
LAM|1|3|猶大 被擄， 遭遇苦難，多服勞役。 她住在列國中，得不著安息； 追逼她的在狹窄之地追上她。
LAM|1|4|錫安 的道路因無人前來過節就哀傷， 她的城門荒涼， 祭司嘆息， 少女悲傷； 她自己充滿痛苦。
LAM|1|5|她的敵人作主， 她的仇敵亨通； 耶和華因她過犯多而使她受苦， 她的孩童在敵人面前去作俘虜。
LAM|1|6|錫安 的威榮全都失去。 她的領袖如找不著草場的鹿， 在追趕的人面前無力行走。
LAM|1|7|耶路撒冷 在困苦窘迫之時， 就追想古時一切的榮華。 她的百姓落在敵人手中，無人幫助； 敵人看見，就因她的毀滅嗤笑。
LAM|1|8|耶路撒冷 犯了大罪， 因此成為不潔淨； 素來尊敬她的，見她裸露就都藐視她， 她自己也嘆息退後。
LAM|1|9|她的污穢是在下襬上； 她未曾思想自己的結局， 她的敗落令人驚詫， 無人安慰她。 「耶和華啊，求你看顧我的苦難， 因為仇敵強大。」
LAM|1|10|敵人伸手奪取她的一切貴重物品； 她眼見列國侵入她的聖所， 你曾吩咐他們不可進入你的集會。
LAM|1|11|她的百姓都嘆息，尋求食物； 他們用貴重物品換取糧食，要救性命。 「耶和華啊，求你觀看， 留意我多麼卑微。」
LAM|1|12|所有過路的人哪，願這事不要發生在你們身上 。 你們要留意觀看， 有像這樣臨到我的痛苦沒有？ 耶和華在他發烈怒的日子使我受苦。
LAM|1|13|他從高處降火進入我的骨頭， 剋制了我； 他張開網，絆我的腳， 使我退後， 又令我終日淒涼發昏。
LAM|1|14|他用手綁我罪過的軛， 捲繞著加在我頸項上； 他使我力量衰敗。 主將我交在我不能抵擋的人手中。
LAM|1|15|主棄絕我們當中所有的勇士， 聚集會眾攻擊我， 要壓碎我的年輕人。 主踹下少女 猶大 ， 在醡酒池中。
LAM|1|16|我因這些事哭泣， 眼淚汪汪； 因為那安慰我、使我重新得力的， 離我甚遠。 我的兒女孤苦， 因為仇敵得勝了。
LAM|1|17|錫安 伸出雙手，卻無人安慰。 論到 雅各 ，耶和華已經出令， 使四圍的人作他的仇敵； 耶路撒冷 在他們中間成為不潔淨。
LAM|1|18|耶和華是公義的！ 我違背了他的命令。 萬民哪，請聽， 來看我的痛苦； 我的少女和壯丁都被擄去。
LAM|1|19|我招呼我所親愛的， 他們卻欺騙了我。 我的祭司和長老尋找食物，要救性命的時候， 就在城中斷了氣。
LAM|1|20|耶和華啊，求你觀看， 因為我在急難中； 我的心腸煩亂， 我心在我裏面翻轉， 因我大大背逆。 在外，刀劍使人喪亡； 在家，猶如死亡。
LAM|1|21|有人聽見我嘆息 ， 卻無人安慰我！ 我所有的仇敵聽見我的患難就喜樂， 因這是你所做的。 你使你所宣告的日子來臨， 願他們像我一樣。
LAM|1|22|願他們的惡行都呈現在你面前； 你怎樣因我一切的罪過待我， 求你也照樣待他們； 因我嘆息甚多，心中發昏。
LAM|2|1|唉！主竟發怒，使黑雲遮蔽 錫安 ！ 他將 以色列 的華美從天扔在地上， 在他發怒的日子並不顧念自己的腳凳。
LAM|2|2|主吞滅 雅各 一切的住處，並不顧惜。 他發怒傾覆 猶大 的堡壘， 將它們夷為平地， 凌辱這國與她的領袖。
LAM|2|3|他發烈怒，砍斷 以色列 一切的角， 在仇敵面前收回右手。 他將 雅各 燒燬，如火焰四圍吞滅。
LAM|2|4|他張弓好像仇敵， 他站立舉起右手， 如同敵人殺戮我們眼目所喜愛的。 他在 錫安 的帳棚 傾倒憤怒，如火一般。
LAM|2|5|主如仇敵吞滅 以色列 ， 吞滅它一切的宮殿， 毀壞境內的堡壘； 在 猶大 加添悲傷和哭號。
LAM|2|6|他摧毀自己的帳幕如摧毀園子， 毀壞自己的會幕。 耶和華使節慶和安息日在 錫安 盡被遺忘， 又在極其憤怒中厭棄君王與祭司。
LAM|2|7|耶和華撇棄自己的祭壇， 憎惡自己的聖所， 把宮殿的牆交給仇敵。 他們在耶和華的殿中喧嚷， 如在節慶之日一樣。
LAM|2|8|耶和華定意拆毀 錫安 的城牆； 他拉了準繩， 不將手收回，定要毀滅。 他使城郭和城牆都悲哀， 一同衰敗。
LAM|2|9|錫安 的門陷入地裏， 主毀壞，折斷她的門閂。 她的君王和官長都置身列國中，沒有律法； 她的先知也不再從耶和華領受異象。
LAM|2|10|錫安 的長老坐在地上，默默無聲； 他們揚起塵土落在頭上，腰束麻布； 耶路撒冷 的少女垂頭至地。
LAM|2|11|我的眼睛流淚，以致失明； 我的心腸煩亂，肝膽落地， 都因我的百姓 遭毀滅， 又因孩童和吃奶的在城內的廣場上昏厥。
LAM|2|12|他們如受傷的人在城內廣場上昏厥， 在母親的懷裏將要喪命時， 就對母親說：「餅和酒在哪裏呢？」
LAM|2|13|耶路撒冷 啊，我可用甚麼向你證明 呢？ 我可用甚麼與你相比呢？ 少女 錫安 哪，我拿甚麼和你比較，好安慰你呢？ 因你的裂傷大如海； 誰能醫治你呢？
LAM|2|14|你的先知為你看見虛假和粉飾的異象， 並未揭露你的罪孽， 使你被擄的歸回； 卻傳給你虛假與誤導人的默示。
LAM|2|15|凡過路的都向你拍掌。 他們向 耶路撒冷 嗤笑，搖頭： 「這就是人稱為全美的、 稱為全地所喜悅的城嗎？」
LAM|2|16|你所有的仇敵 張口來攻擊你； 他們嗤笑，切齒，說： 「我們把她吞滅了， 這是我們所盼望的日子！ 我們終於等到了，親眼看見了！」
LAM|2|17|耶和華成就了他所定的， 應驗了他古時所命定的。 他傾覆，並不顧惜， 他使仇敵向你誇耀， 使你敵人的角高舉。
LAM|2|18|他們的心哀求主。 錫安 的城牆啊， 願你日夜淚流如河，不讓自己休息， 你眼中的瞳人也不歇息。
LAM|2|19|夜間每逢時辰開始，要起來呼喊， 在主面前傾心吐意如水。 你的孩童在街頭上挨餓昏厥， 你要為他們的性命向主舉手。
LAM|2|20|耶和華啊，求你觀看， 留意你向誰這樣行。 婦人豈可吃自己所生、所撫育的嬰孩嗎？ 祭司和先知豈可在主的聖所中被殺嗎？
LAM|2|21|年輕人和老年人躺臥在街上， 我的少女和壯丁都倒在刀下。 你在發怒的日子殺了他們， 你殺戮，並不顧惜。
LAM|2|22|你從四圍招聚使我驚嚇的人， 像在節慶的日子一樣。 耶和華發怒的日子， 無人逃脫，無人生還。 我所撫育養大的， 仇敵都殺盡了。
LAM|3|1|因耶和華憤怒的杖， 我是遭遇困苦的人。
LAM|3|2|他驅趕我走入黑暗， 沒有光明。
LAM|3|3|他反手攻擊我， 終日不停。
LAM|3|4|他使我皮肉枯乾， 折斷我的骨頭。
LAM|3|5|他築壘攻擊我， 以苦楚和艱難圍困我；
LAM|3|6|使我住在幽暗之處， 像死了許久的人一樣。
LAM|3|7|他圍住我，使我無法脫身； 他使我的銅鏈沉重。
LAM|3|8|儘管我哀號求救， 他仍攔阻我的禱告。
LAM|3|9|他用鑿過的石頭擋住我的道路， 使我的路徑彎曲。
LAM|3|10|他向我如埋伏的熊， 如在隱密處的獅子。
LAM|3|11|他使我轉離正路， 把我撕碎 ，使我淒涼。
LAM|3|12|他拉弓，命我站立， 作為箭靶；
LAM|3|13|把箭袋中的箭 射入我的肺腑。
LAM|3|14|我成了全體百姓的笑柄， 成了他們終日的歌曲。
LAM|3|15|他使我受盡苦楚， 飽食茵蔯；
LAM|3|16|用沙石磨斷我的牙， 以灰塵覆蓋我。
LAM|3|17|你使我遠離平安， 我忘了何為福樂。
LAM|3|18|於是我說：「我的力量衰敗， 在耶和華那裏我毫無指望！」
LAM|3|19|求你記得我的困苦和流離， 它如茵蔯和苦膽一般；
LAM|3|20|我心想念這些， 就在我裏面憂悶 。
LAM|3|21|但我的心回轉過來， 因此就有指望；
LAM|3|22|因耶和華的慈愛，我們不致滅絕 ， 因他的憐憫永不斷絕，
LAM|3|23|每早晨，這些都是新的； 你的信實極其廣大！
LAM|3|24|我心裏說：「耶和華是我的福分， 因此，我要仰望他。」
LAM|3|25|凡等候耶和華，心裏尋求他的， 耶和華必施恩給他。
LAM|3|26|人仰望耶和華， 安靜等候他的救恩， 這是好的。
LAM|3|27|人在年輕時負軛， 這是好的。
LAM|3|28|他當安靜獨坐， 因為這是耶和華加在他身上的。
LAM|3|29|讓他臉伏於地 吧！ 或者還會有指望。
LAM|3|30|讓人打他耳光， 使他飽受凌辱吧！
LAM|3|31|主必不永遠撇棄，
LAM|3|32|他雖使人憂愁， 還要照他豐盛的慈愛施憐憫；
LAM|3|33|他並不存心要人受苦， 令世人憂愁。
LAM|3|34|把世上所有的囚犯 踹在腳下，
LAM|3|35|在至高者面前 扭曲人的公正，
LAM|3|36|在人的訴訟上 顛倒是非， 這都是主看不中的。
LAM|3|37|若非主發命令， 誰能說了就成呢？
LAM|3|38|是禍，是福， 不都出於至高者的口嗎？
LAM|3|39|人都有自己的罪， 活人有甚麼好發怨言的呢？
LAM|3|40|讓我們省察，檢討自己的行為， 歸向耶和華吧！
LAM|3|41|讓我們獻上我們的心， 向天上的上帝舉手！
LAM|3|42|我們犯罪悖逆， 你並未赦免。
LAM|3|43|你渾身是怒氣，追趕我們； 你施行殺戮，並不顧惜。
LAM|3|44|你以密雲圍著自己， 禱告不能穿透。
LAM|3|45|你使我們在萬民中 成為污物和垃圾。
LAM|3|46|我們所有的仇敵 張口來攻擊我們；
LAM|3|47|驚嚇和陷阱臨到我們， 殘害和毀滅也臨到我們。
LAM|3|48|因我百姓 遭毀滅， 我的眼睛淚流成河。
LAM|3|49|我的眼睛流淚不停， 流淚不止，
LAM|3|50|直等到耶和華垂顧， 從天上觀看。
LAM|3|51|為我城中的百姓 ， 我眼所見的使我心痛。
LAM|3|52|無故與我為敵的追逼我， 像追捕雀鳥一樣。
LAM|3|53|他們要在坑中了結我的性命， 丟石頭在我身上。
LAM|3|54|眾水淹沒我的頭， 我說：「我沒命了！」
LAM|3|55|耶和華啊， 在極深的地府裏，我求告你的名。
LAM|3|56|我的聲音你聽見了， 求你不要掩耳不聽 我的呼聲，我的求救。
LAM|3|57|我求告你的時候， 你臨近我，說：「不要懼怕！」
LAM|3|58|主啊，你為我伸冤， 你救贖了我的命。
LAM|3|59|耶和華啊，你已看見我的委屈， 求你為我主持正義。
LAM|3|60|他們要報復，謀害我， 你都看見了。
LAM|3|61|耶和華啊，你聽見他們的辱罵， 他們害我的一切計謀，
LAM|3|62|那些起來攻擊我的人嘴唇所說的話 和他們終日攻擊我的計謀。
LAM|3|63|求你留意！ 他們無論坐下或起來， 我都是他們的笑柄。
LAM|3|64|耶和華啊，求你照他們手所做的 向他們施行報應。
LAM|3|65|求你使他們心裏剛硬， 使你的詛咒臨到他們。
LAM|3|66|求你發怒追趕他們， 從耶和華的地上 除滅他們。
LAM|4|1|唉！黃金竟然無光！ 純金竟然變色！ 聖所的石頭散落在街上。
LAM|4|2|錫安 寶貝的孩子雖然好比精金， 現在竟當作陶匠手所做的瓦瓶！
LAM|4|3|野狗尚且哺乳其子， 我百姓 的婦人反倒殘忍， 如曠野的鴕鳥一般；
LAM|4|4|吃奶孩子的舌頭因乾渴貼住上膛， 孩童求餅，卻無人擘給他們。
LAM|4|5|素來吃美好食物的， 如今遭遺棄在街上； 素來穿著朱紅衣裳長大的， 如今卻擁抱糞堆。
LAM|4|6|我百姓的罪孽比 所多瑪 的罪還大； 所多瑪 雖無人伸手攻擊， 轉眼之間就被傾覆。
LAM|4|7|錫安 的拿細耳人 比雪純淨， 比奶更白； 他們的身體比寶石更紅， 身軀之美如藍寶石一般。
LAM|4|8|但如今他們的面貌比煤炭更黑， 在街上無人認識； 他們的皮膚緊貼骨頭， 枯乾形同槁木。
LAM|4|9|被刀劍刺殺的 勝過因飢餓而死 的； 飢餓者由於缺乏田裏的出產 就消瘦而亡 。
LAM|4|10|當我百姓遭毀滅的時候， 慈心的婦人親手烹煮自己的兒女為食物。
LAM|4|11|耶和華發盡他的憤怒， 傾倒他的烈怒， 用火焚燒 錫安 ， 燒燬 錫安 的根基。
LAM|4|12|地上的君王和世上的居民都不信 敵人和仇敵竟能進入 耶路撒冷 的城門。
LAM|4|13|這都因她先知的罪惡和祭司的罪孽， 他們在城中流了義人的血。
LAM|4|14|他們如盲人在街上徘徊， 又被血玷污， 以致人不敢摸他們的衣服。
LAM|4|15|人向他們喊著： 「你這不潔淨的，走開！ 走開！走開！不要摸我！」 他們逃走流浪的時候， 列國中有人說： 「他們不可再寄居此地。」
LAM|4|16|耶和華親自趕散他們， 不再眷顧他們； 不看重祭司，也不厚待長老。
LAM|4|17|我們的眼目徒然仰望幫助，以致失明， 我們從瞭望臺所守望的，竟是一個不能救人的國！
LAM|4|18|仇敵追逐我們的腳蹤， 使我們不敢在自己的街上行走。 我們的結局臨近， 日子已滿， 我們的結局已經來到。
LAM|4|19|追趕我們的比空中的鷹更快； 他們在山上追逼我們， 在曠野埋伏，等候我們。
LAM|4|20|耶和華的受膏者是我們鼻中的氣， 被抓到他們的坑裏， 論到他，我們曾說： 「我們必在他蔭下， 在列國中存活。」
LAM|4|21|住 烏斯 地的 以東 啊，儘管歡喜快樂， 苦杯必傳到你那裏； 你要喝醉，裸露自己。
LAM|4|22|錫安 哪，你罪孽的懲罰已經結束， 耶和華必不再使你被擄去。 以東 啊，耶和華必懲罰你的罪孽， 揭露你的罪惡。
LAM|5|1|耶和華啊，求你顧念我們所遭遇的， 留意看我們所受的凌辱。
LAM|5|2|我們的產業歸陌生人， 我們的房屋歸外邦人。
LAM|5|3|我們是無父的孤兒， 我們的母親如同寡婦。
LAM|5|4|我們出銀錢才得水喝， 我們的柴也是用錢買來的。
LAM|5|5|我們被追趕，迫及頸項， 疲乏卻不得歇息。
LAM|5|6|我們束手投降 埃及 和 亞述 ， 為要得糧吃飽。
LAM|5|7|我們的祖先犯罪，而今他們不在了， 我們卻擔當他們的罪孽。
LAM|5|8|奴僕轄制我們， 無人救我們脫離他們的手。
LAM|5|9|因曠野有刀劍， 我們冒生命的危險才能得糧食。
LAM|5|10|因饑荒的乾熱， 我們的皮膚熱如火爐。
LAM|5|11|他們在 錫安 玷污婦人， 在 猶大 城鎮污辱少女。
LAM|5|12|他們吊起領袖的手， 使長老臉上無光。
LAM|5|13|年輕人扛磨石， 孩童背木柴而跌倒。
LAM|5|14|城門口不再有老年人， 年輕人也不再奏樂。
LAM|5|15|我們心中的快樂止息， 跳舞轉為悲哀。
LAM|5|16|冠冕從我們的頭上掉落； 我們有禍了，因為犯了罪。
LAM|5|17|因這些事我們心裏發昏， 眼睛昏花。
LAM|5|18|錫安山 荒涼， 狐狸行在其上。
LAM|5|19|耶和華啊，你治理直到永遠， 你的寶座萬代長存。
LAM|5|20|你為何全然忘記我們？ 為何長久離棄我們？
LAM|5|21|耶和華啊，求你使我們回轉歸向你， 我們就得以回轉。 求你更新我們的年日，像古時一樣，
LAM|5|22|難道你全然棄絕了我們， 向我們大發烈怒？
