JUDE|1|1|耶穌基督的僕人、 雅各 的兄弟 猶大 ，寫信給那些被召、在父上帝裏蒙愛、為耶穌基督保守的人。
JUDE|1|2|願憐憫、平安 、慈愛多多加給你們！
JUDE|1|3|親愛的，我一直很迫切地想要寫信給你們，論到我們同享的救恩，但我覺得有必要現在就寫信勸你們，要為從前一次交付給聖徒的真道竭力奮鬥。
JUDE|1|4|因為有些人偷偷地進來，就是早就被判定受懲罰的不虔誠的人，他們把我們上帝的恩典變為放縱情慾的機會，並且不認獨一的主宰—我們的主耶穌基督。
JUDE|1|5|這一切的事，你們雖然知道，我卻仍要提醒你們：從前主 只一次就 救了他的百姓出 埃及 地，後來卻把那些不信的滅絕了。
JUDE|1|6|至於那些不守本位、離開自己住處的天使，主用鎖鏈把他們永遠拘留在黑暗裏，等候大日子的審判。
JUDE|1|7|同樣， 所多瑪 、 蛾摩拉 和周圍城鎮的人也跟著他們一樣犯淫亂，隨從逆性的情慾，以致遭受永不熄滅之火的懲罰，作為眾人的鑒戒。
JUDE|1|8|照樣，這些做夢的人也污穢身體，輕慢掌權者，毀謗眾尊榮者。
JUDE|1|9|天使長 米迦勒 為 摩西 的屍首與魔鬼爭辯的時候，尚且不敢用毀謗的話譴責他，只說：「主責備你吧！」
JUDE|1|10|但這些人毀謗他們所不知道的。他們與那些沒有理性的牲畜一樣，只做本性所知道的事，敗壞了自己。
JUDE|1|11|他們有禍了！因為他們走 該隱 的道路，又為財利往 巴蘭 的錯謬裏直奔，並在 可拉 的背叛中滅亡了。
JUDE|1|12|這樣的人是你們愛筵上的污點 ；他們無所懼怕地同你們宴樂，彷彿牧人只顧餵飽自己。他們是無雨的浮雲，被風飄蕩；是秋天沒有果子的樹，死而又死，連根被拔出來；
JUDE|1|13|是海裏的狂浪，湧出自己可恥的沫子來；是流蕩的星，有漆黑的幽暗永遠為他們保留著。
JUDE|1|14|亞當 的七世孫 以諾 曾預言這些人說：「看哪，主帶著他的千萬聖者來臨，
JUDE|1|15|要審判眾人，證實一切不敬虔的人所妄行一切不敬虔的事，又證實不敬虔的罪人所說頂撞他的剛愎的話。」
JUDE|1|16|這些人喜出怨言，責怪他人，隨從自己的情慾而行，口說誇大的話，為自己的利益諂媚人。
JUDE|1|17|親愛的，至於你們，要記得我們主耶穌基督的使徒從前所說的話。
JUDE|1|18|他們曾對你們說過，末世必有好嘲弄的人隨從自己不敬虔的私慾而行。
JUDE|1|19|這就是那些好結黨分派、屬乎血氣、沒有聖靈的人。
JUDE|1|20|親愛的，至於你們，要在至聖的真道上造就自己，藉著聖靈禱告，
JUDE|1|21|保守自己常在上帝的愛中，仰望我們主耶穌基督的憐憫，進入永生。
JUDE|1|22|有些人心中猶疑 ，你們要憐憫 他們；
JUDE|1|23|有些人你們要從火中搶出來，搭救他們 ；有些人你們要存懼怕的心憐憫他們，連那被情慾污染的衣服也要厭惡。
JUDE|1|24|願那能保守你們不失腳，使你們無瑕無疵、歡歡喜喜站在他榮耀之前的、
JUDE|1|25|我們的救主獨一的上帝，藉著我們的主耶穌基督，得享榮耀、威嚴、能力、權柄，從萬古以前，到現今，直到永永遠遠。阿們！
