2KGS|1|1|А по смерті Ахава збунтувався Моав на Ізраїля.
2KGS|1|2|А Ахазія випав через ґрати в своїй горниці, що в Самарії, та й захворів. І послав він послів, і сказав до них: Ідіть, запитайте Ваал-Зевува, екронського бога, чи видужаю я з своєї цієї хвороби?
2KGS|1|3|А Ангол Господній говорив до тішб'янина Іллі: Устань, вийди назустріч послів самарійського царя та й скажи їм: Чи через те, що нема в Ізраїлі Бога, ви йдете питатися Ваал-Зевува, екронського бога?
2KGS|1|4|Тому так сказав Господь: Із того ліжка, що на нього ти ліг, не встанеш із нього, бо напевно помреш!... І пішов Ілля.
2KGS|1|5|І вернулися посли до царя, а він сказав до них: Що це ви вернулися?
2KGS|1|6|А вони відказали йому: Назустріч нам вийшов один чоловік, і сказав нам: Ідіть, верніться до царя, що послав вас, і скажіть йому: Так сказав Господь: Чи через те, що нема в Ізраїлі Бога, ти посилаєш вивідати Ваал-Зевува, екронського бога? Тому те ложе, що на нього ти ліг, не встанеш із нього, бо напевно помреш...
2KGS|1|7|А він їм сказав: Якого вигляду той чоловік, що вийшов назустріч вас, і говорив вам оці слова?
2KGS|1|8|Вони ж відказали: Це чоловік волохатий, а шкуряний пояс оперезаний на стегнах його. А він сказав: Це тішб'янин Ілля!
2KGS|1|9|І послав він до нього п'ятдесятника та його п'ятдесятку. І вийшов він до нього, аж ось він сидить на верхів'ї гори. І сказав він до нього: Чоловіче Божий, цар сказав: Зійди ж ізвідти!
2KGS|1|10|А Ілля відповів і говорив до того п'ятдесятника: А якщо я Божий чоловік, нехай зійде з неба огонь, і нехай пожере тебе та п'ятдесятку твою! І зійшов із неба огонь, і пожер його та його п'ятдесятку...
2KGS|1|11|І цар знову послав до нього іншого п'ятдесятника та його п'ятдесятку. І він відповів і сказав до нього: Чоловіче Божий, отак сказав цар: Зійди ж скоро!
2KGS|1|12|І відповів Ілля та й сказав до нього: Якщо я Божий чоловік, нехай зійде з неба огонь, і нехай пожере тебе та твою п'ятдесятку! І зійшов із неба Божий огонь, і пожер його та його п'ятдесятку...
2KGS|1|13|І знову послав він третього п'ятдесятника та його п'ятдесятку. І вийшов, і прийшов третій п'ятдесятник, та й упав на коліна свої перед Іллею, і благав його та до нього говорив: Чоловіче Божий, нехай же буде дорога душа моя та душа твоїх рабів, тих п'ятидесяти, в очах твоїх!
2KGS|1|14|Ось зійшов був огонь із неба, та й пожер тих двох перших п'ятдесятників та їхні п'ятдесятки; а тепер нехай буде дорога душа моя в очах твоїх!
2KGS|1|15|А Ангол Господній сказав до Іллі: Зійди з ним, не бійся його! І він устав, і зійшов з ним до царя,
2KGS|1|16|Та й сказав до нього: Так сказав Господь: Тому, що ти посилав послів, щоб вивідати від Ваал-Зевува, екронського бога, ніби в Ізраїлі нема Бога, щоб вивідати слова Його, тому те ложе, що на нього ти ліг, не встанеш із нього, бо напевно помреш!
2KGS|1|17|І той помер, за словом Господа, що говорив до Іллі, а замість нього зацарював Єгорам, другого року Єгорама, сина Йосафата, Юдиного царя, бо не було в нього сина.
2KGS|1|18|А решта діл Ахазії, що він зробив був, ото вони написані в Книзі Хроніки Ізраїлевих царів.
2KGS|2|1|І сталося, коли Господь мав узяти Іллю в вихрі на небо, то йшов Ілля та Єлисей із Ґілґалу.
2KGS|2|2|І сказав Ілля до Єлисея: Сиди тут, бо Господь послав мене аж до Бет-Елу. Та Єлисей відказав: Як живий Господь і жива душа твоя, я не залишу тебе! І зійшли вони до Бет-Елу.
2KGS|2|3|І повиходили бет-ельські пророчі сини до Єлисея та й сказали до нього: Чи ти знаєш, що сьогодні Господь бере пана твого від тебе? А він відказав: Я також знаю, мовчіть!
2KGS|2|4|І сказав йому Ілля: Єлисею, сиди тут, бо Господь послав мене до Єрихону. Та той відказав: Як живий Господь і жива душа твоя, я не залишу тебе! І прийшли вони до Єрихону.
2KGS|2|5|І підійшли єрихонські пророчі сини до Єлисея та й сказали до нього: Чи ти знаєш, що сьогодні Господь бере пана твого від тебе? А він відказав: Я також знаю, мовчіть!
2KGS|2|6|І сказав йому Ілля: Сиди тут, бо Господь послав мене до Йордану! Та той відказав: Як живий Господь і жива душа твоя, я не залишу тебе! І пішли вони обоє.
2KGS|2|7|І п'ятдесят чоловіка пророчих синів також пішли, і стали навпроти здалека, а вони обидва стали над Йорданом.
2KGS|2|8|І взяв Ілля плаща свого, і згорнув, і вдарив по воді, і вона розділилась пополовині туди та сюди...
2KGS|2|9|І сталося, як вони перейшли, то Ілля сказав до Єлисея: Проси, що маю зробити тобі, поки я буду взятий від тебе! І сказав Єлисей: Нехай же буде на мені подвійний твій дух!
2KGS|2|10|А той відказав: Тяжкого зажадав ти! Якщо ти побачиш мене, що буду взятий від тебе, буде тобі так, а якщо ні не буде.
2KGS|2|11|І сталося, як вони все йшли та говорили, аж ось появився огняний віз та огняні коні, і розлучили їх одного від одного. І вознісся Ілля в вихрі на небо...
2KGS|2|12|А Єлисей це бачив, і він закричав: Батьку мій, батьку мій, возе Ізраїлів та верхівці його! Та вже не побачив його... І схопився він сильно за одежу свою та й роздер її на дві частині.
2KGS|2|13|І підняв він Іллевого плаща, що спав із нього, і вернувся, і став на березі Йордану.
2KGS|2|14|І взяв він Іллевого плаща, що спав із нього, і вдарив по воді та сказав: Де Господь, Бог Іллі? І також він ударив по воді, і вона розділилася пополовині туди та сюди!...
2KGS|2|15|І побачили його знавпроти єрихонські пророчі сини, та й сказали: На Єлисеї спочив дух Іллів! І пішли вони назустріч йому, і попадали перед ним до землі,
2KGS|2|16|та й сказали до нього: Ось із твоїми рабами є п'ятдесят чоловіка хоробрих, нехай вони підуть та пошукають твого пана, а ну ж забрав його Дух Господній, і кинув його на одну з гір або в одну з долин! А той відказав: Не посилайте!
2KGS|2|17|Та вони сильно благали його, аж докучили йому, то він сказав: Посилайте! І послали вони п'ятдесят чоловіка, і шукали три дні, та не знайшли його.
2KGS|2|18|І вони вернулися до нього (а він мешкав в Єрихоні). І сказав він до них: Чи ж не казав я вам: Не йдіть?
2KGS|2|19|І сказали люди того міста Єлисеєві: Ось положення цього міста хороше, як пан бачить, та вода нехороша, а земля неплідна.
2KGS|2|20|А він сказав: Подайте мені нового дзбанка, і покладіть туди соли. І вони подали йому.
2KGS|2|21|І він вийшов до джерела води, і кинув туди соли й сказав: Так сказав Господь: Уздоровив Я цю воду, не буде вже звідти смерти, ані непліддя!
2KGS|2|22|І була вилікувана та вода, і так є аж до цього дня, за словом Єлисея, яке він говорив.
2KGS|2|23|І відійшов він звідти до Бет-Елу. А коли він ішов дорогою, то малі хлопці виходили з того міста й насміхалися з нього, і казали йому: Ходи, лисий! Ходи, лисий!
2KGS|2|24|І він обернувся назад і побачив їх, та й прокляв їх Іменем Господнім. І вийшли дві ведмедиці з лісу, і розірвали з них сорок і двоє дітей...
2KGS|2|25|А він пішов звідти до гори Кармел, а звідти вернувся до Самарії.
2KGS|3|1|А Єгорам, Ахавів син, зацарював над Ізраїлем у Самарії, у вісімнадцятому році Йосафата, Юдиного царя, і царював дванадцять років.
2KGS|3|2|І чинив він лихо в Господніх очах, тільки не так, як батько його та мати його, він викинув Ваалового боввана, що зробив був батько його.
2KGS|3|3|Проте гріхів Єровоама, Неватового сина, що вводив у гріх Ізраїля, він тримався, і не відставав від них.
2KGS|3|4|А Меша, цар моавський, розводив дрібну худобу, і давав Ізраїлевому цареві сто тисяч ягнят та сто тисяч рунних баранів.
2KGS|3|5|І сталося, як помер Ахав, то збунтувався моавський цар проти Ізраїлевого царя.
2KGS|3|6|І вийшов того дня цар Єгорам із Самарії, і перелічив усього Ізраїля.
2KGS|3|7|І пішов він, і послав до Йосафата, царя Юдиного, говорячи: Збунтувався проти мене цар моавський. Чи підеш зо мною на війну до Моаву? А той відказав: Вийду. Я як ти, мій народ як твій народ, мої коні як твої коні!
2KGS|3|8|І сказав: Котрою дорогою підемо? А той відказав: Дорогою едомської пустині.
2KGS|3|9|І пішов цар Ізраїлів, і цар Юдин, і цар едомський, і йшли обхідною дорогою сім день. І не було води таборові та худобі, що була при них.
2KGS|3|10|І сказав Ізраїлів цар: Ах, Господь викликав трьох оцих царів, щоб віддати їх у руку Моава.
2KGS|3|11|І сказав Йосафат: Чи нема тут Господнього пророка, щоб через нього вивідати слово Господа? І відповів один із слуг Ізраїлевого царя й сказав: Тут є Єлисей, Шафатів син, що служив Іллі.
2KGS|3|12|І сказав Йосафат: Слово Господнє з ним! І зійшли до нього цар Ізраїлів, і Йосафат, і цар едомський.
2KGS|3|13|І сказав Єлисей до Ізраїлевого царя: Що тобі до мене? Іди до пророків батька свого та до пророків своєї матері! А Ізраїлів цар відказав йому: Ні, бо Господь покликав трьох цих царів, щоб віддати їх у руку Моава.
2KGS|3|14|І сказав Єлисей: Як живий Господь Саваот, що я стою перед лицем Його, коли б я не зважав на Йосафата, Юдиного царя, не споглянув би на тебе, і не побачив би я тебе.
2KGS|3|15|А тепер приведіть мені гусляра. І сталося, коли грав гусляр, то на Єлисеї була Господня рука,
2KGS|3|16|і він сказав: Так сказав Господь: Накопайте на цій долині яму за ямою!
2KGS|3|17|Бо так сказав Господь: Не побачите вітру, і не побачите дощу, а потік цей буде наповнений водою. І будете пити ви, та череди ваші, та ваша худоба.
2KGS|3|18|Та буде цього мало в Господніх очах, і Він видасть і Моава в вашу руку.
2KGS|3|19|І ви поб'єте всяке укріплене місто та всяке місто вибране, і всяке добре дерево повалите, і всі водні джерела загатите, і всяку добру полеву ділянку завалите камінням.
2KGS|3|20|І сталося ранком, коли приноситься хлібна жертва, аж ось полилася вода з едомської дороги. І наповнилася земля водою.
2KGS|3|21|А ввесь Моав почув, що ті царі вийшли воювати з ними. І вони скликали всіх, хто носить пояса й старше, і поставали на границі.
2KGS|3|22|І повставали вони рано вранці, і сонце засвітило над водою. І побачили моавляни навпроти воду, червону, як кров.
2KGS|3|23|І казали вони: Це кров, рубаючися, порубалися царі мечами, і позабивали один одного. А тепер на здобич, Моаве!
2KGS|3|24|І прийшли вони до Ізраїлевого табору. І встав Ізраїль та й побив моавлян, і ті повтікали перед ними. І вони ввійшли до них, і били моавлян,
2KGS|3|25|а міста руйнували, і на всяку добру польову ділянку усі кидали свого каменя й закидали її, і всяке джерело води загачували, і валили всяке добре дерево, й аж тільки в Кір-Харешеті позоставили каміння його. І оточили тарани, та й били його.
2KGS|3|26|І побачив моавський цар, що бій перемагає його, і взяв він сім сотень чоловіка, що орудують мечем, щоб продертися до едомського царя, та не зміг.
2KGS|3|27|І він узяв свого перворідного сина, що мав царювати замість нього, і приніс його цілопаленням на мурі... І повстав великий гнів на Ізраїля, і вони відступили від нього, і вернулися до свого краю.
2KGS|4|1|А одна з жінок пророчих синів кликала до Єлисея, говорячи: Помер раб твій, мій чоловік! А ти знаєш, що раб твій боявся Господа. А позичальник прийшов ось, щоб забрати собі двоє дітей моїх за рабів...
2KGS|4|2|І сказав до неї Єлисей: Що я зроблю тобі? Розкажи мені, що є в тебе в домі. А та відказала: Нічого нема в домі твоєї невільниці, є тільки горня оливи.
2KGS|4|3|А він сказав: Іди, позич собі настороні посуд від усіх сусідок твоїх, посуд порожній. Не бери мало!
2KGS|4|4|І ввійдеш, і замкнеш двері за собою та за синами своїми, і поналиваєш у всі ті посудини, а повні повідставляй.
2KGS|4|5|І пішла вона від нього, і замкнула двері за собою та за синами своїми. Вони подавали їй посуд, а вона наливала.
2KGS|4|6|І сталося, коли понаповнювано посуд, то сказала вона до сина свого: Подай мені ще посуду! А він відказав їй: Нема вже посуду. І спинилася олива.
2KGS|4|7|І вона прийшла, і донесла Божому чоловікові. І він сказав: Іди, продай ту оливу, та й заплати своєму позичальникові. А ти та сини твої будете жити на позостале.
2KGS|4|8|І сталося певного дня, і прийшов Єлисей до Шунаму, а там була багата жінка, і вона сильно просила його до себе поїсти хліба. І бувало, скільки разів приходив він, заходив туди їсти хліб.
2KGS|4|9|І сказала вона до чоловіка свого: Ось я познала, що Божий чоловік, який завжди приходить до нас, він святий.
2KGS|4|10|Зробім же малу муровану горницю, і поставимо йому там ліжко, і стола, і стільця, і свічника. І коли він приходитиме до нас, то заходитиме туди.
2KGS|4|11|Одного разу прийшов він туди, і зайшов до горниці та й ліг там.
2KGS|4|12|І сказав він до свого слуги Ґехазі: Поклич оцю шунамітянку! І той покликав її, і вона стала перед ним.
2KGS|4|13|І сказав він до нього: Скажи їй: Ось ти старанно піклувалася про всі наші потреби. Що зробити тобі за це? Чи є що, щоб сказати про тебе цареві або начальникові війська? А вона відказала: Ні, я сиджу серед народу свого!
2KGS|4|14|І сказав він: Що ж зробити їй? А Ґехазі відказав: Та вона не має сина, а чоловік її старий.
2KGS|4|15|А він сказав: Поклич її. І він покликав її, і вона стала при вході.
2KGS|4|16|І він сказав: На цей означений час, коли саме цей час вернеться, ти обійматимеш сина! А вона відказала: Ні, пане, чоловіче Божий, не говори неправди своїй невільниці!
2KGS|4|17|Та зачала та жінка, і породила сина на той означений час, того саме часу, про який говорив до неї Єлисей.
2KGS|4|18|І росло те дитя. А одного разу вийшло воно до свого батька до женців.
2KGS|4|19|І сказало воно до свого батька: Голова моя, голова моя!... А той сказав слузі: Занеси його до його матері!
2KGS|4|20|І той поніс його, і приніс його до його матері. І сиділо воно на її колінах аж до полудня, та й померло...
2KGS|4|21|І ввійшла вона, і поклала його на ліжко Божого чоловіка, і замкнула за ним двері та й вийшла.
2KGS|4|22|І покликала вона свого чоловіка та й сказала: Пришли мені одного із слуг та одну з ослиць, і я поїду до Божого чоловіка й вернуся.
2KGS|4|23|А він сказав: Чому ти їдеш до нього? Сьогодні не новомісяччя й не субота. А вона відказала: Добре!
2KGS|4|24|І осідлала вона ослицю, і сказала до свого слуги: Поганяй та йди. Не затримуй мені в їзді, аж поки не скажу тобі.
2KGS|4|25|І поїхала вона, і приїхала до Божого чоловіка, до гори Кармел. І сталося, як Божий чоловік побачив її здалека, то сказав до слуги свого Ґехазі: Ось та шунамітянка!
2KGS|4|26|Побіжи ж назустріч їй та й скажи їй: Чи все гаразд тобі, чи гаразд чоловікові твоєму, чи гаразд дитині? А та відказала: Усе гаразд!
2KGS|4|27|І прийшла вона до Божого чоловіка на гору, і сильно схопила за ноги його. А Ґехазі підійшов, щоб відіпхнути її, та Божий чоловік сказав: Позостав її, бо затурбована душа її, а Господь затаїв це передо мною й не сказав мені.
2KGS|4|28|А вона сказала: Чи я жадала сина від пана? Чи я не говорила: Не впроваджуй мене в обману?
2KGS|4|29|І він сказав до Ґехазі: Опережи стегна свої, і візьми мою палицю в руку свою та й іди. Коли спіткаєш кого, не повітаєш його, а коли хто повітає тебе, не відповіси йому. І покладеш мою палицю на хлопцеве обличчя.
2KGS|4|30|А мати того хлопця сказала: Як живий Господь і жива душа твоя, я не полишу тебе! І він устав і пішов за нею.
2KGS|4|31|А Ґехазі пішов перед ними, і поклав ту палицю на хлопцеве обличчя, та не було ані голосу, ані чуття. І вернувся він навпроти нього, і доніс йому, говорячи: Не збудився той хлопець!
2KGS|4|32|І ввійшов Єлисей у дім, аж ось той хлопець лежить мертвий на ліжку його!...
2KGS|4|33|І ввійшов він, і замкнув двері за ними обома, та й молився до Господа.
2KGS|4|34|І ввійшов він, і ліг на того хлопця, і поклав уста свої на уста його, а очі свої на очі його, і долоні свої на долоні його. І схилився над ним, і стало тепле тіло тієї дитини!...
2KGS|4|35|І він знову ходив по дому раз сюди, а раз туди. І ввійшов він, і знову схилився над ним, і чхнув той хлопець аж до семи раз. І розплющив той хлопець очі свої.
2KGS|4|36|І покликав він Ґехазі та й сказав: Поклич ту шунамітянку! І той покликав її. І прийшла вона до нього, і він сказав: Забери свого сина!
2KGS|4|37|І ввійшла вона, і впала до його ніг, і вклонилася до землі. І взяла вона сина свого та й вийшла...
2KGS|4|38|І вернувся Єлисей до Ґілґалу. А в Краю був голод, і пророчі сини сиділи перед ним. І сказав він до свого хлопця: Пристав великого горшка, і звари їжу для пророчих синів.
2KGS|4|39|І вийшов один на поле, щоб назбирати ярини, і знайшов там витку рослину, і назбирав із неї повну свою одежу диких огірків. І він прийшов, і накришив до горшка їжі, бо вони не знали того.
2KGS|4|40|І поналивали вони людям їжі. І сталося, як вони їли ту їжу, то закричали й сказали: Смерть у горшку, чоловіче Божий! І не могли вони їсти...
2KGS|4|41|А він сказав: Дайте муки! І він всипав її до горшка і сказав: Наливай народові, і нехай їдять! І вже не було нічого злого в горшку.
2KGS|4|42|І прийшов один чоловік із Баал-Шалішу, і приніс Божому чоловікові хліб первоплоду, двадцять ячмінних хлібців та зерна в колосках у своїй торбі. І сказав Єлисей: Дай народові, і нехай вони їдять!
2KGS|4|43|А слуга його сказав: Що оце покладу я перед сотнею чоловіка? Та він відказав: Дай народові, і нехай їдять, бо так сказав Господь: Їжте й позоставте!
2KGS|4|44|І він поклав перед ними, і вони їли й позоставили, за словом Господнім.
2KGS|5|1|А Нааман, начальник війська сирійського царя, був муж великий перед своїм паном, вельмиповажаний, бо через нього Господь дав перемогу Сирії. І був це муж дуже хоробрий, але прокажений.
2KGS|5|2|А сирійці вийшли були ордами, і взяли до неволі з Ізраїлевого краю малу дівчину, і вона услуговувала жінці Наамана.
2KGS|5|3|І сказала вона до своєї пані: Ох, коли б пан мій побував у того пророка, що в Самарії, то він вилікував би його від прокази його!
2KGS|5|4|А Нааман прийшов, і доніс своєму панові, говорячи: Отак і отак говорила та дівчина, що з Ізраїлевого краю.
2KGS|5|5|І сказав сирійський цар: Тож піди, а я пошлю свого листа до Ізраїлевого царя. І той пішов, і взяв із собою десять талантів срібла та шість тисяч шеклів золота, і десять змін одежі.
2KGS|5|6|І він приніс до Ізраїлевого царя такого листа: Ось тепер, як прийде оцей лист до тебе, то знай: ото послав я до тебе свого раба Наамана, а ти вилікуєш його від прокази його.
2KGS|5|7|І сталося, як Ізраїлів цар перечитав цього листа, то роздер свої шати й сказав: Чи я Бог, щоб убивати чи лишати при житті, що той посилає до мене, щоб я вилікував чоловіка від прокази його? Тож знайте й дивіться це він шукає проти мене зачіпки.
2KGS|5|8|І сталося, як почув Єлисей, Божий чоловік, що Ізраїлів цар роздер шати свої, то послав до царя, говорячи: Нащо роздер ти шати свої? Нехай той прийде до мене, і пізнає, що є пророк ув Ізраїлі!
2KGS|5|9|І прибув Нааман зо своїми кіньми та з колесницею своєю, і став при вході Єлисеєвого дому.
2KGS|5|10|І послав Єлисей до нього посла, говорячи: Іди, і вимиєшся сім раз у Йордані, і вигоїться тіло твоє тобі, й очистишся.
2KGS|5|11|І розгнівався Нааман, і пішов і сказав: Ось я подумав був: він вийде до мене, і стане, і закличе Ім'я Господа, Бога свого, і покладе свою руку на те місце, і вилікує прокаженого...
2KGS|5|12|Чи ж не ліпші Авана та Парпар, дамаські річки, від усіх Ізраїлевих вод? Чи не міг я вимитися в них, і стати чистим? І повернувся він, і пішов у гніві.
2KGS|5|13|І підійшли його раби, і говорили до нього, і сказали: Батьку мій, коли б велику річ говорив тобі той пророк, чи ж ти не зробив би? А що ж, коли він сказав тобі тільки: Умийся і будеш чистий!
2KGS|5|14|І зійшов він, і занурився в Йордані сім раз, за словом Божого чоловіка. І сталося тіло його, як тіло малого хлопця, і став він чистий!
2KGS|5|15|І вернувся до Божого чоловіка він та ввесь табір його. І прийшов він, і став перед ним та й сказав: Оце пізнав я, що на всій землі нема Бога, а тільки в Ізраїлі! А тепер візьми дарунка від свого раба.
2KGS|5|16|Та Єлисей відказав: Як живий Господь, що стою перед лицем Його, я не візьму! А той сильно просив його взяти, та він відмовився.
2KGS|5|17|І сказав Нааман: А як ні, то нехай буде дано твоєму рабові землі, скільки понесуть два мули, бо твій раб не буде вже приносити цілопалення та жертву іншим богам, а тільки Господеві!
2KGS|5|18|Тільки оцю річ нехай простить Господь твоєму рабові: коли мій пан прийде до Ріммонового дому, щоб там поклонятися, і опиратиметься на мою руку, то й я схилюся в Ріммоновім домі. Коли я кланятимуся в Ріммоновім домі, то нехай простить Господь твоєму рабові цю річ!
2KGS|5|19|А той відказав: Іди з миром! І відійшов від нього на невелику відстань.
2KGS|5|20|І сказав Ґехазі, слуга Єлисея, чоловіка Божого: Ось мій пан стримав цього сиріянина Наамана, щоб нічого не взяти з руки його, що він приніс. Як живий Господь, побіжу за ним і візьму щось від нього!...
2KGS|5|21|І погнався Ґехазі за Нааманом. І побачив Нааман бігуна за собою, і зіскочив із воза навпроти нього й сказав: Чи все гаразд?
2KGS|5|22|А той відказав: Гаразд! Пан мій послав мене, говорячи: Ось тепер прийшла до мене з Єфремових гір двоє юнаків, пророчі сини. Дай їм талант срібла та дві зміні одежі!
2KGS|5|23|А Нааман відказав: Будь ласкав, візьми два таланти! І він упрошував його. І зав'язав він два таланти срібла в дві торбі, та дві зміні одежі, і дав своїм слугам, а вони понесли перед ним.
2KGS|5|24|І прийшов він до згір'я, і взяв з їхньої руки, і вмістив у домі, а тих людей відпустив, і вони пішли.
2KGS|5|25|А він прийшов та й став перед паном своїм. І сказав до нього Єлисей: Звідки ти, Ґехазі? А той відказав: Нікуди не ходив твій раб, ані туди, ані сюди...
2KGS|5|26|І сказав Єлисей до нього: Чи моє серце не ходило з тобою, коли обернувся той муж зо свого воза назустріч тобі? Чи час брати срібло та брати одежі, і оливки, і виноградника, і худобу дрібну та худобу велику, і рабів, і невільниць?
2KGS|5|27|Тож Нааманова проказа нехай приліпиться до тебе та до насіння твого навіки! І той вийшов від нього прокажений, побілівши, як сніг!...
2KGS|6|1|І сказали пророчі сини до Єлисея: Ось те місце, де ми сидимо перед тобою, затісне для нас.
2KGS|6|2|Ходім аж до Йордану, і візьмімо звідти кожен по одній деревині, і зробимо собі місце, щоб сидіти там. А він сказав: Ідіть.
2KGS|6|3|І сказав один: Будь же ласкавий, і ходи зо своїми рабами! А він сказав: Я піду.
2KGS|6|4|І пішов він із ними, і вони прийшли до Йордану, і рубали дерево.
2KGS|6|5|І сталося, коли один валив деревину, то впала сокира до води. А той скрикнув і сказав: Ох, пане мій, таж вона позичена!
2KGS|6|6|І сказав Божий чоловік: Куди вона впала? А той показав йому те місце. І він відрубав кусок дерева й кинув туди, і випливла сокира!...
2KGS|6|7|І він сказав: Витягни собі! А той простяг свою руку і взяв...
2KGS|6|8|Сирійський цар воював з Ізраїлем. І радився він зо слугами своїми, говорячи: На такому то й такому то місці буде моє таборування.
2KGS|6|9|А Божий чоловік послав до Ізраїлевого царя, говорячи: Стережися переходити оце місце, бо там сходяться сиріяни!
2KGS|6|10|І послав Ізраїлів цар до того місця, про яке говорив йому Божий чоловік та остерігав його; і він стерігся там не раз і не два.
2KGS|6|11|І сильно занепокоїлося серце сирійського царя про ту річ, і він покликав своїх слуг та й сказав до них: Чи не розповісте мені, хто з наших зраджує перед Ізраїльським царем?
2KGS|6|12|І сказав один з його слуг: Ні, пане мій царю, це не наш, а це Єлисей, той пророк, що в Ізраїлі, доносить Ізраїлевому цареві ті слова, що ти говориш у спальні своїй!...
2KGS|6|13|А він відказав: Ідіть, і подивіться, де він, і я пошлю й візьму його! І донесено йому, кажучи: Ось він у Дотані!
2KGS|6|14|І послав він туди коні, і колесниці та військо. І прийшли вони вночі й оточили те місто.
2KGS|6|15|А слуга Божого чоловіка встав рано і вийшов, аж ось військо оточує місто, і коні, і колесниці! І сказав його слуга до нього: Ох, пане мій, що будемо робити?
2KGS|6|16|А той відказав: Не бійся, бо ті, що з нами, численніші від тих, що з ними.
2KGS|6|17|І молився Єлисей і говорив: Господи, розкрий йому очі, і нехай він побачить! І відкрив Господь очі того слуги, і він побачив, аж ось гора повна коней та огняних колесниць навколо Єлисея!...
2KGS|6|18|І зійшли сирійці до нього, а Єлисей помолився до Господа й сказав: Удар цей люд сліпотою! І Він ударив їх сліпотою за Єлисеєвим словом...
2KGS|6|19|І сказав до них Єлисей: Це не та дорога й не те місто. Ідіть за мною, й я проведу вас до того чоловіка, якого ви шукаєте. І він завів їх у Самарію.
2KGS|6|20|І сталося, як прийшли вони до Самарії, то Єлисей сказав: Господи, відкрий оці очі, і нехай вони побачать! І Господь відкрив їхні очі, і вони побачили, аж ось вони в середині Самарії!...
2KGS|6|21|І сказав Ізраїлів цар до Єлисея, коли побачив їх: Чи побити їх, чи побити, мій батьку?
2KGS|6|22|А той відказав: Не вбивай! Чи ти повбиваєш тих, кого ти взяв до неволі своїм мечем та своїм списом? Поклади хліб та воду перед ними, і нехай вони їдять та п'ють, і нехай ідуть до свого пана.
2KGS|6|23|І справив цар для них велику гостину, і вони їли й пили; і він відпустив їх, і вони пішли до свого пана. І сирійські орди вже більш не входили до Ізраїлевого Краю.
2KGS|6|24|І сталося по тому, і зібрав Бен-Гадад, сирійський цар, увесь свій табір, і він зійшов і обліг Самарію.
2KGS|6|25|І був великий голод у Самарії. І ось ті облягали їх, а осляча голова коштувала вісімдесят шеклів срібла, а чвертка каву голубиного помету п'ять шеклів срібла.
2KGS|6|26|І сталося, проходив Ізраїлів цар по мурі, а одна жінка крикнула до нього, говорячи: Поможи, пане царю!
2KGS|6|27|А він відказав: Як тобі не поможе Господь, звідки я поможу тобі? Чи з току, або з чавила?
2KGS|6|28|І сказав до неї цар: Що тобі? А та відказала: Оця жінка сказала мені: Дай свого сина, і ми з'їмо його сьогодні, а мого сина з'їмо взавтра.
2KGS|6|29|І зварили ми мого сина та й з'їли його... І сказала я до неї другого дня: Дай сина свого, і ми з'їмо його, та вона сховала свого сина.
2KGS|6|30|І сталося, як цар почув слова цієї жінки, то роздер шати свої, і він ходив по мурі. І народ побачив, аж ось веретище на тілі його зо споду!
2KGS|6|31|І він сказав: Отак нехай зробить мені Бог, і так нехай додасть, якщо позостанеться голова Єлисея, Шафатового сина, на ньому сьогодні!
2KGS|6|32|А Єлисей сидів у своєму домі, а з ним сиділи старші. І послав цар чоловіка від себе. Поки прийшов посол до нього, то він сказав до старших: Чи ви бачите, що цей син убивника послав зняти мою голову? Глядіть, як прийде цей посол, то замкніть двері, і притиснете його в дверях. Ось і шарудіння ніг пана його за ним.
2KGS|6|33|Ще він говорив із ними, аж ось приходить до нього посланець. І він сказав: Отаке зло від Господа! Чого ще чекати від Господа?
2KGS|7|1|І сказав Єлисей: Послухайте слово Господнє: Так сказав Господь: Цього часу взавтра буде сея пшеничної муки за шекля, і дві сеї ячменю за шекля в брамі Самарії.
2KGS|7|2|І відповів Божому чоловікові вельможа царя, що він на його руку спирався, і сказав: Якби Господь поробив отвори в небі, чи сталася б ця річ? А той відказав: Ось ти побачиш своїми очима, та їсти звідти не будеш.
2KGS|7|3|І були при вході до брами чотири прокажені чоловіки. І сказали вони один до одного: Чого ми сидимо тут, аж поки не помремо?
2KGS|7|4|Якщо ми скажемо: Увійдімо до міста, а в місті голод, то помремо там; а якщо сидітимемо тут, то теж помремо. Отож, ходіть, і перейдімо до сирійського табору, якщо там позоставлять нас при житті, будемо жити, а якщо заб'ють нас, то помремо...
2KGS|7|5|І встали вони надвечір, щоб іти до сирійського табору. І прибули вони до краю сирійського табору, аж ось нема там нікого!
2KGS|7|6|Бо Господь учинив, що сирійський табір почув стукотняву колесниць і їржання коней, та галас великого війська. І сказали вони один до одного: Ось Ізраїлів цар найняв на нас хіттейських царів та царів єгипетських, щоб пішли на нас!
2KGS|7|7|І встали вони, і повтікали надвечір, і полишили свої намети, й осли свої, і табір, як він був, та й повтікали, спасаючи життя своє!
2KGS|7|8|І прийшли ті прокажені аж до краю табору, і ввійшли до одного намету, і їли й пили, і повиносили звідти срібло й золото та вбрання, і пішли й заховали. І вони знову ввійшли до іншого намету, і повиносили звідти, і пішли та й сховали.
2KGS|7|9|І сказали вони один до одного: Неслушно ми робимо. Цей день він день доброї звістки, а ми мовчимо. Як ми будемо чекати аж до ранішнього світла, то впаде на нас провина. А тепер ходімо, і ввійдімо й донесімо царевому дому!
2KGS|7|10|І прийшли вони, і покликали міських воротарів, та й донесли їм, говорячи: Увійшли ми до сирійського табору, а там нема ані людини, ані людського голосу, а тільки поприв'язувані коні та поприв'язувані осли, та намети, як вони були!
2KGS|7|11|І воротарі покликали, і донесли про це до самого царського дому.
2KGS|7|12|І встав цар уночі й сказав своїм слугам: Розкажу я вам, що нам зробили сирійці. Вони знають, що ми голодні, і повиходили з табору, щоб сховатися на полі, говорячи: Коли ті повиходять із міста, то ми схопимо їх живих, та й увійдемо до міста!
2KGS|7|13|І відповів один із його слуг і сказав: Нехай візьмуть п'ятеро позосталих коней, що лишилися в ньому, у місті. Ось вони, (із усього війська Ізраїлевого тільки й лишилися, із усього війська Ізраїля, що згинуло), і пошлемо, і побачимо.
2KGS|7|14|І взяли вони дві колесниці з кіньми, і цар послав їх услід за сирійським табором, говорячи: Ідіть і подивіться.
2KGS|7|15|І пішли вони за ними аж до Йордану, аж ось уся дорога повна вбрання та речей, що покидали сирійці, як поспішали! І вернулися ці посли, і донесли цареві.
2KGS|7|16|І вийшов народ, і розграбували сирійський табір. І коштувала сея пшеничної муки по шеклю, і дві сеї ячменю по шеклю за словом Господнім!
2KGS|7|17|І цар призначив того вельможу, що на його руку він опирався, доглядати над брамою. Та затоптав його народ у брамі, і він помер, як казав був Божий чоловік, який говорив, коли приходив до нього цар.
2KGS|7|18|І сталося, коли Божий чоловік говорив до царя, кажучи: Дві сеї ячменю по шеклю, і сея пшеничної муки по шеклю буде того часу взавтра в брамі Самарії,
2KGS|7|19|то цей вельможа відповів Божому чоловікові й сказав: Якби Господь поробив отвори в небі, чи сталася б ця річ? А той відказав: Ось ти побачиш своїми очима, та їсти звідти не будеш.
2KGS|7|20|І сталося йому так, і затоптав його народ у брамі, і він помер...
2KGS|8|1|А Єлисей говорив до жінки, що її сина він воскресив, кажучи: Устань та й іди ти та дім твій, і мешкай дебудь, бо Господь прикликав голод, і він прийшов до краю на сім літ.
2KGS|8|2|І встала та жінка, і зробила за словом Божого чоловіка. І пішла вона та її дім, і замешкала в филистимському краї сім літ.
2KGS|8|3|І сталося наприкінці семи років, вернулася та жінка з филистимського краю, і пішла до царя благати за свій дім та за своє поле.
2KGS|8|4|А цар говорив до Ґехазі, слуги Божого чоловіка, кажучи: Розкажи мені про все те велике, що зробив Єлисей.
2KGS|8|5|І сталося, як він оповідав цареві, що той воскресив померлого, аж ось та жінка, що він воскресив сина її, благає царя за свій дім та за своє поле.
2KGS|8|6|І сказав Ґехазі: Пане мій царю, оце та жінка, і це той син її, що воскресив Єлисей!
2KGS|8|7|І прийшов Єлисей до Дамаску, а Бен-Гадад, сирійський цар, хворий. І донесено йому, кажучи: Божий чоловік прийшов аж сюди!
2KGS|8|8|І сказав цар до Газаїла: Візьми в свою руку подарунка, та й іди зустріти чоловіка Божого. І запитайся Господа через нього, кажучи: Чи видужаю я від оцієї хвороби?
2KGS|8|9|І пішов Газаїл спіткати його, і взяв подарунка в руку свою, та зо всього добра Дамаску тягару на сорок верблюдів. І прийшов, і став перед ним та й сказав: Син твій Бен-Гадад, цар сирійський, послав мене до тебе, питаючи: Чи видужаю я з оцієї хвороби?
2KGS|8|10|І сказав до нього Єлисей: Іди, скажи йому: Жити житимеш, та Господь показав мені, що напевно помре він.
2KGS|8|11|І наставив він обличчя своє на нього, і довго вдивлявся, аж той збентежився. І заплакав Божий чоловік.
2KGS|8|12|А Газаїл сказав: Чого плаче мій пан? А той відказав: Бо знаю, що ти зробиш лихо Ізраїлевим синам: їхні твердині пустиш з огнем, і їхніх вояків позабиваєш мечем, і дітей їхніх порозбиваєш, а їхне вагітне посічеш...
2KGS|8|13|А Газаїл сказав: Та що таке твій раб, цей пес, що зробить таку велику річ? І сказав Єлисей: Господь показав мені тебе царем над Сирією!
2KGS|8|14|І пішов він від Єлисея, і прийшов до свого пана. А той сказав йому: Що говорив тобі Єлисей? І він сказав: Говорив мені: жити житимеш!
2KGS|8|15|І сталося другого дня, і взяв він покривало, і намочив у воді, і поклав на його обличчя, і той помер. І зацарював Газаїл замість нього.
2KGS|8|16|А п'ятого року Йорама, Ахавого сина, Ізраїлевого царя, за Йосафата, Юдиного царя, зацарював Єгорам, син Йосафатів, цар Юдин.
2KGS|8|17|Він був віку тридцяти й двох літ, коли зацарював, а царював вісім літ в Єрусалимі.
2KGS|8|18|І ходив він дорогою Ізраїлевих царів, як робив Ахавів дім, бо Ахавова дочка була йому за жінку. І робив він зло в Господніх очах.
2KGS|8|19|Та не хотів Господь погубити Юду ради раба Свого Давида, як обіцяв був йому дати світильника йому та синам його по всі дні.
2KGS|8|20|За його днів збунтувався був Едом, вийшли з-під Юдиної руки, і настановили над собою царя.
2KGS|8|21|І пішов Йорам до Цаіру, а з ним усі колесниці. І сталося, коли він уночі встав і побив Едома, що оточив був його, і керівників колесниць, то народ повтікав до наметів своїх.
2KGS|8|22|І збунтувався Едом, і вийшов з-під Юдиної руки, і так є аж до цього дня. Тоді того часу збунтувалася й Лівна.
2KGS|8|23|А решта діл Йорама, та все, що він зробив, ось вони написані в Книзі Хроніки Юдиних царів.
2KGS|8|24|І спочив Йорам із батьками своїми, і був похований із батьками своїми в Давидовому Місті, а замість нього зацарював син його Ахазія.
2KGS|8|25|У дванадцятому році Йорама, Ахавого сина, Ізраїлевого царя, зацарював Ахазія, син Єгорама, Юдиного царя.
2KGS|8|26|Ахазія був віку двадцяти і двох літ, коли він зацарював, і царював він один рік в Єрусалимі. А ім'я його матері Аталія, дочка Омрі, Ізраїлевого царя.
2KGS|8|27|І ходив він дорогою Ахавого дому, і робив зло в Господніх очах, як і Ахавів дім, бо він був зять Ахавого дому.
2KGS|8|28|І пішов він з Йорамом, Ахавовим сином, на війну з Газаїлом, сирійським царем, до ґілеадського Рамоту, та побили сиріяни Йорама.
2KGS|8|29|І вернувся цар Йорам лікуватися в Їзреелі від тих ран, що вчинили йому сиріяни в Рамі, як він воював з Газаїлом, сирійським царем. А Ахазія, Єгорамів син, цар Юдин, зійшов побачити Йорама, Ахавового сина, в Їзреелі, бо той був слабий.
2KGS|9|1|А пророк Єлисей покликав одного з пророчих синів і сказав йому: Підпережи свої стегна, і візьми це горня оливи в свою руку, і йди до ґілеадського Рамоту.
2KGS|9|2|І прийдеш туди, і побач там Єгу, сина Йосафата, Німшієвого сина. І ти ввійдеш, і візьмеш його з-між братів його, і введеш його до внутрішньої кімнати.
2KGS|9|3|І візьмеш горня цієї оливи, і виллєш на його голову та й скажеш: Так сказав Господь: Помазую тебе на царя над Ізраїлем! А по тому відчиниш двері й утечеш, і не будеш чекати.
2KGS|9|4|І пішов той слуга, слуга пророка, до ґілеадського Рамоту.
2KGS|9|5|І прийшов він, аж ось сидять керівники війська. І він сказав: Слово мені до тебе, о керівнику! А Єгу відказав: До кого з усіх нас? І той сказав: До тебе, о керівнику!
2KGS|9|6|І він устав, і вийшов до дому, а той вилив оливу на його голову. І сказав він йому: Так сказав Господь, Бог Ізраїля: Помазую тебе на царя над народом Господнім, над Ізраїлем!...
2KGS|9|7|І ти поб'єш дім Ахава, пана свого, і помстиш за кров Моїх рабів пророків, і за кров усіх Господніх рабів від руки Єзавелі.
2KGS|9|8|І згине ввесь Ахавів дім, і вигублю Ахавові навіть те, що мочиться на стіну, і невільного та вільного в Ізраїлі!
2KGS|9|9|І зроблю Ахавів дім, як дім Єровоама, Неватового сина, і як дім Баші, сина Ахійїного.
2KGS|9|10|А Єзавелю з'їдять пси в Їзреелевій ділянці, і не буде, хто б її поховав. І відчинив він двері та й утік...
2KGS|9|11|А Єгу вийшов до слуг свого пана, і вони сказали йому: Чи все гаразд? Чого приходив той несамовитий до тебе? А він відказав: Ви знаєте того чоловіка та його мову.
2KGS|9|12|А вони відказали: Неправда! Розкажи ж нам! І той сказав: Отак і так сказав він до мене, говорячи: Так сказав Господь: Помазую тебе на царя над Ізраїлем!
2KGS|9|13|А ті поспішно взяли кожен шати свої, і постелили під ним на верху сходів. І засурмили вони в сурму, і сказали: Зацарював Єгу!
2KGS|9|14|І змовився Єгу, син Йосафата, Німшієвого сина, проти Йорама. А Йорам стеріг ґілеадського Рамота, він та ввесь Ізраїль перед Газаїлом, сирійським царем.
2KGS|9|15|І вернувся цар Єгорам лікуватися в Їзреелі від ран, що вчинили йому сиріяни, як він воював з Газаїлом, сирійським царем. І сказав Єгу: Якщо згода ваша на те, нехай не вийде жоден утікач із міста, щоб піти донести в Їзреелі.
2KGS|9|16|І сів верхи Єгу, і поїхав до Їзреелу, бо Йорам лежав там. А Ахазія, цар Юдин, зійшов побачити Йорама.
2KGS|9|17|А на башті в Їзреелі стояв вартовий. І побачив він натовп Єгуїв, як він ішов, і сказав: Я бачу натовп! А Єгорам відказав: Візьми верхівця, і пошли назустріч їм, і нехай він скаже: Чи все гаразд?
2KGS|9|18|І відправився верхівець назустріч йому, і сказав: Так сказав цар: Чи все гаразд? А Єгу відказав: Що тобі до того? Повертай за мною! І доніс вартовий, говорячи: Прийшов той посол аж до них, та не вернувся.
2KGS|9|19|І послав він другого верхівця, і він прийшов до них та й сказав: Так сказав цар: Чи все гаразд? А Єгу відказав: Що тобі до гаразду? Повертай за мною!
2KGS|9|20|І доніс вартовий, говорячи: Прийшов він аж до них, та не вернувся. А кінна їзда, як їзда Єгу, Німшієвого сина, бо їде несамовито.
2KGS|9|21|І сказав Єгорам: Запрягай! І запріг його колесницю. І відправився Єгорам, Ізраїлів цар, та Ахазія, Юдин цар, кожен своєю колесницею, щоб зустріти Єгу, і спіткали його в ділянці їзреелянина Навота.
2KGS|9|22|І сталося, як Єгорам побачив Єгу, то сказав: Чи все гаразд, Єгу? А той відказав: Який гаразд при перелюбі твоєї матері Єзавелі та її багатьох чарів?
2KGS|9|23|І обернув Єгорам руки свої та й утік. І сказав він Ахазії: Зрада, Ахазіє!
2KGS|9|24|А Єгу взяв лука в руку свою, і вдарив Єгорама між його раменами, і пробила стріла його серце, і він похилився на колесниці своїй...
2KGS|9|25|І сказав Єгу до Бідкара, вельможі свого: Візьми, кинь його на ділянці поля їзреелянина Навота. Бо пам'ятай, я й ти їхали вдвох за Ахавом, батьком його, а Господь прорік на нього оце пророцтво:
2KGS|9|26|Поправді кажу, що бачив Я вчора кров Навота та кров синів його, говорить Господь, і відплачу тобі на цій же ділянці, говорить Господь. А тепер кинь його на цій ділянці за словом Господнім.
2KGS|9|27|А Ахазія, Юдин цар, побачив це, і втікав дорогою на Бет-Гаґґан, а Єгу погнався за ним і сказав: Убийте й його на колесниці! І поранили його в Маале-Ґурі, що при Ївлеамі, а він утік до Меґіддо та й помер там.
2KGS|9|28|А раби його відвезли його верхи до Єрусалиму, та й поховали його в його гробі з батьками його в Давидовому Місті.
2KGS|9|29|А в одинадцятому році Йорама, Ахавового сина, над Юдою зацарював Ахазія.
2KGS|9|30|І прийшов Єгу до Їзрееля, а Єзавель почула про це, і нафарбувала очі свої, і прикрасила голову свою, та й виглянула через вікно.
2KGS|9|31|А Єгу входить до брами. І сказала вона: Чи все гаразд, Зімрі, убивце пана свого?
2KGS|9|32|І підняв він обличчя своє до вікна та й сказав: Хто зо мною, хто? І виглянули до нього два-три євнухи.
2KGS|9|33|А він сказав: Скиньте її! І викинули її, і бризнула кров її на стіну та на коні. І він топтав її...
2KGS|9|34|І він увійшов, і їв та пив, та й сказав: Підіть до тієї проклятої, і поховайте її, бо все ж таки вона царева дочка!
2KGS|9|35|І пішли поховати її, та не знайшли з неї нічого, а тільки черепа, та ноги, та долоні рук...
2KGS|9|36|І вони вернулися, і донесли йому про це. А він відказав: Це слово Господа, що казав був через раба Свого тішб'янина Іллю, говорячи: В Їзреелевій ділянці пси з'їдять Єзавелине тіло!
2KGS|9|37|І буде Єзавелин труп, як погній на поверхні поля в Їзреелевій ділянці, так що не скажуть: Це Єзавель...
2KGS|10|1|А Ахав мав сімдесят синів у Самарії. І понаписував Єгу листи, і порозсилав до Самарії, до провідників Їзреелу, до старших і до виховників Ахавових синів, говорячи:
2KGS|10|2|Як тільки прийде лист цей до вас, а з вами сини вашого пана, і з вами колесниці, і коні, і твердині, і зброя,
2KGS|10|3|то виберіть найліпшого та найвідповіднішого з синів вашого пана, і посадіть його на трон вашого батька, та й воюйте за дім вашого пана!
2KGS|10|4|А вони дуже-дуже налякалися й сказали: Ось два царі не встояли перед ним, якже встоїмо ми?
2KGS|10|5|І послали ті, що були над домом та над тим містом, і старші, і виховники до Єгу, говорячи: Ми раби твої, і зробимо все, що ти нам скажеш. Та ми не настановимо царем нікого, що добре в очах твоїх, те роби!
2KGS|10|6|А він написав до них другого листа, пишучи: Якщо ви мої, і слухняні моєму голосові, візьміть голови мужів, синів вашого пана, і прийдіть до мене цього часу взавтра до Їзреелу (а царських синів було сімдесят чоловіка, при міських вельможах, що виховали їх).
2KGS|10|7|І сталося, як прийшов той лист до них, то побрали вони царських синів, та й позабивали сімдесят чоловіка. І поскладали вони їхні голови в кошики, та й послали до нього в Їзреел...
2KGS|10|8|І прибув посол, і доніс йому, кажучи: Принесли голови царських синів! А він сказав: Покладіть їх на дві купі при вході до брами до ранку.
2KGS|10|9|І сталося вранці, і він вийшов і став, і сказав до всього народу: Ви невинні. Я вчинив змову на свого пана й убив його. А хто повбивав усіх цих?
2KGS|10|10|Знайте ж тепер, що з Господнього слова не проминеться нічого, що Господь говорив на Ахавів дім, і Господь зробив те, що говорив був через раба Свого Іллю.
2KGS|10|11|І Єгу повбивав усіх позосталих з Ахавого дому в Їзреелі, і всіх вельмож його, і знайомих його, і священиків його, так, що не позоставив йому і врятованого!
2KGS|10|12|І встав він і відійшов, і пішов до Самарії. А коли він був на дорозі при Бет-Екед-Гароімі,
2KGS|10|13|то спіткав братів Ахазії, Юдиного царя, і сказав: Хто ви? А ті відказали: Ми Ахазієві брати, а йдемо запитати про гаразд царевих синів та синів цариці!
2KGS|10|14|А він сказав: Схопіть їх живих! І схопили їх живих, і позабивали їх до ями Бет-Екеду, сорок і два чоловіка, і він не позоставив ані одного з них!
2KGS|10|15|І пішов він ізвідти, і спіткав Єгонадава, Рехавового сина, що йшов навпроти нього, і привітав його та й сказав до нього: Чи твоє серце щире до мене, як моє серце до тебе? А Єгонадав відказав: Так! Дай же свою руку! І той дав руку свою, і підняв його до себе до колесниці,
2KGS|10|16|і сказав: Іди ж зо мною, і приглянься до моєї запопадливости для Господа! І посадили його в колесницю його.
2KGS|10|17|І прибув він до Самарії, і повбивав усіх позосталих в Ахава в Самарії, і вибив аж до кінця його, за словом Господа, що говорив до був Іллі.
2KGS|10|18|І зібрав Єгу ввесь народ і сказав до них: Ахав мало служив Ваалові, Єгу служитиме йому більше!
2KGS|10|19|А тепер покличте до мене всіх пророків Ваала, усіх, хто служить йому, та всіх священиків. Нехай нікого не бракуватиме, бо в мене велика жертва для Ваала. Кожен, хто буде відсутній, не буде живий! А Єгу зробив це підступом, щоб вигубити тих, хто служить Ваалові.
2KGS|10|20|І сказав Єгу: Оголосіть святочні збори для Ваала! І вони оголосили.
2KGS|10|21|І послав Єгу по всьому Ізраїлю. І посходилися всі, хто служить Ваалові, і не позостався ніхто, хто не прийшов би. І прибули вони до Ваалового дому, і переповнився Ваалів дім від входу до входу.
2KGS|10|22|І сказав він тому, хто над царською шатнею: Винеси одежу для всіх тих, хто служить Ваалові. І той виніс їм ту одежу.
2KGS|10|23|І ввійшов Єгу та Єгонадав, Рехавів син, до Ваалового дому, і сказав до Ваалових служителів: Пошукайте й подивіться, щоб не був тут із вами ніхто з Господніх слуг, а тільки самі ті, хто служить Ваалові.
2KGS|10|24|І ввійшли вони, щоб принести жертви та цілопалення. А Єгу поставив собі назовні вісімдесят чоловіка й сказав: Кожен, у кого втече хто з тих людей, що я ввів на ваші руки, життя його буде за життя того!
2KGS|10|25|І сталося, як скінчив він приряджувати цілопалення, то Єгу сказав до бігунів та до старшин: Увійдіть, повбивайте їх, нехай ніхто не вийде!... І повбивали їх вістрям меча, і поскидали їх ті бігуни та старшини. Потому пішли до міста Ваалового дому.
2KGS|10|26|І повиносили вони бовванів Ваалового дому, і попалили те.
2KGS|10|27|І розбили вони Ваалового боввана, і розбили Ваалів дім, та й зробили з нього нечисте місце, і так є аж до сьогодні.
2KGS|10|28|І вигубив Єгу Ваала з Ізраїля.
2KGS|10|29|Тільки не відступив він від гріхів Єровоама, Неватового сина, що вводив у гріх Ізраїля, від золотих тельців, що в Бет-Елі та що в Дані.
2KGS|10|30|І сказав Господь до Єгу: Тому, що ти добре зробив угодне в очах Моїх, зробив Ахавовому домові все, що було на серці Моєму, сидітимуть сини твої на Ізраїлевому троні аж до четвертого покоління.
2KGS|10|31|Та Єгу не пильнував ходити за Законом Господа, Бога Ізраїля, усім своїм серцем, не відступив від гріхів Єровоама, що вводив у гріх Ізраїля.
2KGS|10|32|За тих днів розпочав Господь відрубувати від Ізраїля частини, і побив їх Газаїл в усій Ізраїлевій країні,
2KGS|10|33|від Йордану на схід сонця, увесь край Ґілеаду, Ґадів, Рувимів та Манасіїн, від Ароеру, що над потоком Арнон, і Ґілеад та Башан.
2KGS|10|34|А решта діл Єгу, і все, що він зробив, і вся лицарськість його, ось вони написані в Книзі Хроніки Ізраїлевих царів.
2KGS|10|35|І спочив Єгу зо своїми батьками, і поховали його в Самарії, а замість нього зацарював син його Єгоахаз.
2KGS|10|36|А дні, що царював Єгу над Ізраїлем у Самарії, були двадцять і вісім літ.
2KGS|11|1|А коли Аталія, мати Ахазії, побачила, що помер її син, то встала та й вигубила все цареве насіння.
2KGS|11|2|А Єгошева, дочка царя Йорама, сестра Ахазії, взяла Йоаша, сина Ахазії, та й викрала його з-поміж вбиваних царських синів, його та няньку його, і сховала в спальній кімнаті. І сховали його від Аталії, і він не був забитий.
2KGS|11|3|І ховався він із нею в Господньому домі шість років, а Аталія царювала над краєм.
2KGS|11|4|А сьомого року послав Єгояда, і взяв сотників із карійців та бігунів, і привів їх до себе до Господнього дому, і склав із ними умову, і заприсягнув їх у Господньому домі, і показав їм царського сина.
2KGS|11|5|І він наказав їм, говорячи: Оце та річ, яку зробите. Третина з вас, що приходите в суботу, будете виконувати сторожу царського дому.
2KGS|11|6|А третина буде в брамі Сур, а третина у брамі за бігунами, і будете виконувати сторожу дому на зміну.
2KGS|11|7|А дві частині з вас, усі, що відходять у суботу, будуть виконувати сторожу Господнього дому при цареві.
2KGS|11|8|І оточите царя навколо, кожен із своєю зброєю в руці своїй; а хто ввійшов би до рядів, нехай буде забитий. І будете ви з царем при виході його та при вході його.
2KGS|11|9|І зробили сотники все, що наказав священик Єгояда. І взяли кожен людей своїх, що приходять у суботу та виходять у суботу, і прийшли до священика Єгояди.
2KGS|11|10|І дав священик сотникам списи та щити, що належали цареві Давидові, що були в Господньому домі.
2KGS|11|11|І поставали бігуни, кожен зо зброєю своєю в руці своїй, від правого боку дому аж до лівого боку дому, при жертівнику та при домі, навколо біля царя.
2KGS|11|12|А він вивів царевого сина, і поклав на нього корону та нараменники. І зробили вони його царем, і помазали його, і вдарили в долоні та й крикнули: Нехай живе цар!
2KGS|11|13|І почула Аталія голос бігунів та народу, і прийшла до народу до Господнього дому.
2KGS|11|14|І побачила вона, аж ось цар стоїть за звичаєм на помості, а при царі зверхники та сурми, а ввесь народ краю тішиться та сурмить у сурми. І роздерла Аталія шати свої та й крикнула: Зрада, зрада!
2KGS|11|15|А священик Єгояда наказав сотникам, поставленим над військом, і сказав до них: Випровадьте її поза ряди, а хто піде за нею, того забийте мечем! Бо священик сказав: Нехай вона не буде забита в Господньому домі!
2KGS|11|16|І зробили їй прохід, і вона прийшла Кінським входом до царського дому, і там була забита.
2KGS|11|17|І склав Єгояда заповіта між Господом та між царем і між народом, щоб був народом Господнім, і між царем та між народом.
2KGS|11|18|І ввійшов увесь народ Краю до Ваалового дому, та й порозбивали його та жертівники його, і бовванів його зовсім поламали, а Маттана, Ваалового священика, убили перед жертівниками. А при Господньому домі священик поставив варти.
2KGS|11|19|І взяв він сотників і карійців, і бігунів та ввесь народ краю, і вивели царя з Господнього дому. І ввійшли вони через браму бігунів до царського дому, і той сів на царському троні.
2KGS|11|20|І тішився ввесь народ краю, а місто заспокоїлось. А Аталію вбили мечем у царському домі.
2KGS|11|21|(12-1) Єгоаш був віку семи років, коли зацарював.
2KGS|12|1|(12-2) Сьомого року Єгу зацарював Єгоаш, і сорок років царював він в Єрусалимі. А ім'я його матері Ців'я, з Беер-Шеви.
2KGS|12|2|(12-3) І робив Єгоаш угодне в Господніх очах по всі дні, коли вказував йому священик Єгояда.
2KGS|12|3|(12-4) Тільки пагірки не були понищені, народ ще приносив жертви та кадив на пагірках.
2KGS|12|4|(12-5) І сказав Єгоаш до священика: Усе посвячене срібло, що буде внесене до Господнього дому, срібло перелічених людей, срібло за душі за вартістю їх, усе срібло, скільки людині спаде на серце принести до Господнього дому,
2KGS|12|5|(12-6) візьмуть собі священики, кожен від знайомого свого, і вони зроблять направу Господнього дому в усьому, що буде знайдене там на направу.
2KGS|12|6|(12-7) І сталося двадцятого й третього року царя Єгоаша, священики не направили ушкодження храму.
2KGS|12|7|(12-8) І покликав цар Єгоаш священика Єгояду й священиків, та й сказав їм: Чому ви не направляєте ушкодження храму? А тепер не беріть срібла від ваших знайомих, а на направу ушкодження храму віддасте його.
2KGS|12|8|(12-9) І погодилися священики не брати срібла від народу, і не направляти ушкодження храму.
2KGS|12|9|(12-10) І взяв священик Єгояда одну скриньку, і продовбав дірку на віку її, і поставив її при жертівнику праворуч, як входити до Господнього дому. І давали туди священики, що стерегли порога, усе срібло, що приносилося до Господнього дому.
2KGS|12|10|(12-11) І бувало, як вони бачили, що намножилося те срібло в скрині, то приходив царський писар та великий священик, і вони в'язали в мішки та рахували срібло, знайдене в Господньому домі.
2KGS|12|11|(12-12) І давали те перелічене срібло на руки робітникам праці, поставленим до Господнього дому, а вони давали його теслям та будівничим, що робили в Господньому домі.
2KGS|12|12|(12-13) І мулярам, і каменярам, і на закуп дерева та тесаного каменя, та на направу ушкодження Господнього дому, та на все, що йшло на храм для направи.
2KGS|12|13|(12-14) Тільки не робилися для Господнього дому срібні чаші, ножиці, кропильниці, сурми, усяка річ золота та річ срібна з того срібла, що приносилося до Господнього дому,
2KGS|12|14|(12-15) бо його давали робітникам праці та направляли ним дім Господній.
2KGS|12|15|(12-16) І не облічували тих людей, яким давали те срібло до їхніх рук, щоб вони давали робітникам праці, бо ті робили чесно.
2KGS|12|16|(12-17) Срібло ж жертви за провину та жертов за гріх не вносилося до Господнього дому, воно було для священиків.
2KGS|12|17|(12-18) Вийшов тоді Газаїл, сирійський цар, та й воював з Ґатом, і здобув його. І намірився Газаїл іти на Єрусалим.
2KGS|12|18|(12-19) І взяв Єгоаш, Юдин цар, усі святі речі, що присвятили були Йосафат, і Єгорам, і Ахазія, батьки його, царі Юдині, та святі речі свої, і все золото, що знайшлося в скарбницях Господнього дому та дому царського, та й послав Газаїлові, цареві сирійському, і той відійшов від Єрусалиму...
2KGS|12|19|(12-20) А решта діл Йоаша, і все, що він зробив, он вони написані в Книзі Хроніки Юдиних царів.
2KGS|12|20|(12-21) І встали його слуги, і вчинили змову, та й забили Йоаша в Бет-Мілло, де йдеться до Сілли.
2KGS|12|21|(12-22) Йозахар, Шім'атів син, та Єгозавад, Шомерів син, його слуги, забили його, і він помер. І поховали його з батьками його в Давидовім Місті, а замість нього зацарював син його Амація.
2KGS|13|1|Двадцятого й третього року Йоаша, сина Ахазії, Юдиного царя, зацарював над Ізраїлем у Самарії Єгоахаз, син Єгу, на сімнадцять літ.
2KGS|13|2|І робив він зло в Господніх очах, і ходив у гріхах Єровоама, Неватового сина, що вводив у гріх Ізраїля, і не відхилявся від того.
2KGS|13|3|І запалився гнів Господа на Ізраїля, і Він дав їх у руку Газаїла, царя сирійського, та в руку Бен-Гадада, Газаїлового сина, на всі ті дні.
2KGS|13|4|Та вблагав Єгоахаз лице Господнє, і Господь його вислухав, бо бачив Він горе Ізраїля, бо тиснув їх сирійський цар.
2KGS|13|5|І дав Господь Ізраїлеві спасителя, і вони вийшли з-під руки Сирії. І сиділи Ізраїлеві сини в своїх наметах, як давніш.
2KGS|13|6|Тільки не відійшли вони з гріхів дому Єровоама, що вводив у гріх Ізраїля, і сам у тому ходив, і Астарта стояла в Самарії.
2KGS|13|7|А Сирія не позоставила Єгоахазові народу, як тільки п'ятдесят верхівців та десять возів, та десять тисяч піхоти, бо їх вигубив сирійський цар, і зробив їх порохом на топтання.
2KGS|13|8|А решта діл Єгоахаза, і все, що він робив, та його лицарськість, он вони написані в Книзі Ізраїлевих царів.
2KGS|13|9|І спочив Єгоахаз з батьками своїми, і поховали його в Самарії, а замість нього зацарював син його Йоаш.
2KGS|13|10|Тридцятого й сьомого року Йоаша, Юдиного царя, зацарював над Ізраїлем у Самарії Йоаш, Єгоахазів син, на шістнадцять літ.
2KGS|13|11|І робив він зле в Господніх очах, і не відходив від усіх гріхів Єровоама, Неватового сина, що вводив у гріх Ізраїля, і в тому ходив.
2KGS|13|12|А решта діл Йоаша, і все, що він робив, і лицарськість його, як він воював з Амацією, Юдиним царем, он вони написані в Книзі Хроніки Ізраїлевих царів.
2KGS|13|13|І спочив Йоаш з батьками своїми, а Єровоам сів на троні його. І був похований Йоаш у Самарії, з Ізраїлевими царями.
2KGS|13|14|А Єлисей заслаб на недугу, що з неї й помер. І зійшов до нього Йоаш, Ізраїлів цар, і плакав над ним і говорив: Батьку мій, батьку мій, колеснице Ізраїлева та верхівці його!
2KGS|13|15|І сказав йому Єлисей: Візьми лука та стріли. І приніс той до нього лука та стріли.
2KGS|13|16|А він сказав Ізраїлевому цареві: Поклади свою руку на лука! І той поклав свою руку. А Єлисей поклав свої руки на руки цареві.
2KGS|13|17|І він сказав: Відчини вікно на схід! І той відчинив. І сказав Єлисей: Стріляй! І той вистрілив, а він сказав: Стріла спасіння Господнього, і стріла спасіння проти Сирії. І поб'єш ти Сирію в Афеку аж до кінця!
2KGS|13|18|І він сказав: Візьми стріли! І той узяв, а він сказав до Ізраїлевого царя: Удар по землі! І він ударив три рази та й став.
2KGS|13|19|І розгнівався на нього Божий чоловік і сказав: Щоб ти був ударив п'ять або шість раз, тоді побив би Сирію аж до кінця! А тепер тільки три рази поб'єш ти Сирію.
2KGS|13|20|І спочив Єлисей, і поховали його. А моавські орди прийшли до Краю наступного року.
2KGS|13|21|І сталося, як ховали одного чоловіка, то погребальники побачили ті орди, та й кинули того чоловіка до Єлисеєвого гробу. А коли впав і доторкнувся той чоловік до Єлисеєвих костей, то воскрес, і встав на ноги свої...
2KGS|13|22|А Газаїл, сирійський цар, тиснув Ізраїля всі дні Єгоахаза.
2KGS|13|23|Та Господь був милостивий до них, і змилувався над ними, і звернувся до них ради заповіта Свого з Авраамом, Ісаком та Яковом, і не хотів вигубити їх, і не відкинув їх від Свого лиця аж дотепер.
2KGS|13|24|І спочив Газаїл, сирійський цар, а замість нього зацарював син його Бен-Гадад.
2KGS|13|25|І Йоаш, Єгоахазів син, узяв назад ті міста з руки Бен-Гадада, Газаїлового сина, що взяв був із руки Єгоахаза, свого батька, у війні. Три рази побив його Йоаш, і вернув Ізраїлеві міста.
2KGS|14|1|Другого року Йоаша, Йоахазового сина, Ізраїлевого царя, зацарював Амація, Йоашів син, цар Юдин.
2KGS|14|2|Він був віку двадцяти й п'яти літ, коли зацарював, і царював в Єрусалимі двадцять і дев'ять років. А ім'я його матері Єгоаддан, з Єрусалиму.
2KGS|14|3|І робив він угодне в Господніх очах, тільки не так, як його батько Давид, він робив усе, що робив його батько Йоаш.
2KGS|14|4|Тільки пагірки не були знищені, народ приносив жертву та кадив на пагірках.
2KGS|14|5|І сталося, як зміцнилося царство в руці його, то він повбивав своїх слуг, що забили його батька царя.
2KGS|14|6|А синів убійників він не позабивав, як написано в Книзі Мойсеєвого Закону, що наказав був Господь, говорячи: Не будуть забиті батьки за синів, а сини не будуть забиті за батьків, а тільки кожен за гріх свій буде забитий.
2KGS|14|7|Він побив Едома в Соляній долині, десять тисяч, і взяв у війні Селу, і назвав ім'я їй: Йоктеїл, і так вона зветься аж до цього дня.
2KGS|14|8|Тоді Амація послав послів до Йоаша, сина Єгоахаза, сина Єгу, Ізраїлевого царя, говорячи: Іди ж, поміряємось!
2KGS|14|9|І послав Йоаш, Ізраїлів цар, до Амації, Юдиного царя, говорячи: Терен, що на Ливані, послав до кедрини, що на Ливані, кажучи: Дай же дочку свою моєму синові за жінку! Та перейшла польова звірина, що на Ливані, і витоптала той терен.
2KGS|14|10|Побити побив ти Едома, і піднесло тебе твоє серце. Пишайся собі та сиди в своїм домі! І пощо будеш ти дрочитися зо злом, бо впадеш ти та Юда з тобою?
2KGS|14|11|Та не послухався Амація. І вийшов Йоаш, Ізраїлів цар, і помірялися він та Амація, цар Юдин, у Юдиному Бет-Шемеші.
2KGS|14|12|І був розбитий Юда Ізраїлем, і повтікали кожен до намету свого.
2KGS|14|13|А Йоаш, цар Ізраїлів, схопив Амацію, Юдиного царя, сина Йоаша, сина Ахазії, у Бет-Шемеші, і прибув до Єрусалиму, і зруйнував єрусалимський мур від Єфремової брами аж до брами наріжної, чотири сотні ліктів.
2KGS|14|14|І забрав він усе золото й срібло, та ввесь посуд, що знаходився в Господньому домі та в скарбницях дому царевого, та запоручників, і вернувся в Самарію.
2KGS|14|15|А решта діл Йоаша, що зробив він, та лицарськість його, і як воював з Амацією, Юдиним царем, ось вони написані в Книзі Хроніки Ізраїлевих царів.
2KGS|14|16|І спочив Йоаш зо своїми батьками, і був похований у Самарії з Ізраїлевими царями, а замість нього зацарював син його Єровоам.
2KGS|14|17|І жив Амація, Йоашів син, цар Юдин, по смерті Йоаша, Єгоахазового сина, Ізраїлевого царя, п'ятнадцять літ.
2KGS|14|18|А решта діл Амації, ось вони написані в Книзі Хроніки Юдиних царів.
2KGS|14|19|І вчинили на нього змову в Єрусалимі, та він утік до Лахішу. І послали за ним до Лахішу, і вбили його там.
2KGS|14|20|І повезли його на конях, і він був похований з батьками своїми в Давидовому Місті.
2KGS|14|21|І взяв ввесь Юдин народ Азарію, а він був віку шістнадцяти літ, і настановили його царем замість батька його Амації.
2KGS|14|22|Він збудував Елат, і вернув його Юді, як цар спочив зо своїми батьками.
2KGS|14|23|П'ятнадцятого року Амації, сина Йоаша, Юдиного царя, зацарював Єровоам, син Йоаша, Ізраїлевого царя, у Самарії, на сорок і один рік.
2KGS|14|24|І робив він зло в Господніх очах, не відступався від усіх гріхів Єровоама, Неватового сина, що вводив у гріх Ізраїля.
2KGS|14|25|Він вернув Ізраїлеву границю відти, де йдеться до Гамату, аж до степового моря, за словом Господа, Бога Ізраїля, що говорив через раба Свого Йону, сина пророка Амміттая, що з Ґат-Гахеферу,
2KGS|14|26|бо Господь побачив Ізраїлеву біду, дуже гірку, і не було вже невільного та вільного, і не було помічника Ізраїлеві.
2KGS|14|27|Та не говорив Господь знищити Ізраїлеве ім'я з-під неба, і споміг їх рукою Єровоама, Йоашового сина.
2KGS|14|28|А решта діл Єровоама та лицарськість його, як воював, і як вернув Юді Дамаск та Хамат в Ізраїлі, ось вони написані в Книзі Хроніки Ізраїлевих царів.
2KGS|14|29|І спочив Єровоам із батьками своїми та з Ізраїлевими царями, а замість нього зацарював син його Захарій.
2KGS|15|1|Двадцятого й сьомого року Єровоама, Ізраїлевого царя, зацарював Азарія, син Амації, Юдиного царя.
2KGS|15|2|Він був віку шістнадцяти літ, коли зацарював, і царював в Єрусалимі п'ятдесят і два роки. А ім'я його матері Єхолія, з Єрусалиму.
2KGS|15|3|І робив він угодне в Господніх очах, усе так, як робив його батько Амація.
2KGS|15|4|Тільки пагірки не були знищені, народ ще приносив жертву та кадив на пагірках.
2KGS|15|5|І вдарив Господь царя, і він був прокажений аж до дня своєї смерти, і сидів ув осібному домі. А над домом був Йотам, царів син, він судив народ Краю.
2KGS|15|6|А решта діл Азарії та все, що він робив, ось вони написані в Книзі Хроніки Юдиних царів.
2KGS|15|7|І спочив Азарія з своїми батьками, і його поховали з його батьками в Давидовому Місті, а замість нього зацарював син його Йотам.
2KGS|15|8|Тридцятого й восьмого року Азарії, Юдиного царя, зацарював над Ізраїлем у Самарії Захарій, син Єровоама, на шість місяців.
2KGS|15|9|І робив він зле в Господніх очах, як робили батьки його, не відступився від гріхів Єровоама, Наватового сина, що вводив у гріх Ізраїля.
2KGS|15|10|І вчинив змову на нього Шаллум, Явешів син, і бив його перед народом і вбив його, і зацарював замість нього.
2KGS|15|11|А решта діл Захарія, ось вони написані в Книзі Хроніки Ізраїлевих царів.
2KGS|15|12|Оце Господнє слово, що Він промовляв до Єгу, говорячи: Сини чотирьох поколінь будуть сидіти тобі на Ізраїлевому троні. І сталося так.
2KGS|15|13|Шаллум, Явешів син, зацарював тридцятого й дев'ятого року Уззійї, Юдиного царя, і царював місяць часу в Самарії.
2KGS|15|14|І пішов Менахем, Ґадіїв син, з Тірци, і прибув у Самарію, та й побив Шаллума, Явешового сина, в Самарії, і вбив його, і зацарював замість нього.
2KGS|15|15|А решта днів Шаллума та змова його, яку він учинив був, ото вони написані в Книзі Хроніки Ізраїлевих царів.
2KGS|15|16|Тоді побив Менахем місто Тіфсах та все, що в ньому, і границі його від Тірци, бо не відчинило воно брами. І він вибив його, а все вагітне повитинав.
2KGS|15|17|Тридцятого й дев'ятого року Азарії, Юдиного царя, зацарював над Ізраїлем у Самарії Менахем, Ґадіїв син, на десять літ.
2KGS|15|18|І робив він зле в Господніх очах, не вступився від гріхів Єровоама, Неватового сина, що вводив у гріх Ізраїля. За його днів
2KGS|15|19|прийшов Пул, асирійський цар, на край. І дав Менахем Пулові тисячу талантів срібла, щоб його руки були з ним, щоб зміцнити царство в його руці.
2KGS|15|20|А Менахем розклав це срібло на Ізраїля, на всіх вояків, щоб дати асирійському цареві, по п'ятдесят шеклів срібла від кожного чоловіка. І вернувся асирійський цар, і не стояв там у Краю.
2KGS|15|21|А решта діл Менахема та все, що він робив, ото вони написані в Книзі Хроніки Ізраїлевих царів.
2KGS|15|22|І спочив Менахем з батьками своїми, а замість нього зацарював син його Пекахія.
2KGS|15|23|П'ятдесятого року Азарії, Юдиного царя, зацарював над Ізраїлем у Самарії Пекахія, син Менахемів, на два роки.
2KGS|15|24|І робив він зло в Господніх очах, не відступався від гріхів Єровоама, Неватового сина, що вводив у гріх Ізраїля.
2KGS|15|25|І вчинив на нього змову Пеках, син Ремалії, старшина його, і забив його в палаті царського дому, з Арґовом та з Ар'єм, а з ним було п'ятдесят чоловіка з ґілеадян. І він убив його, і зацарював замість нього.
2KGS|15|26|А решта діл Пекахії та все, що він робив, ото вони написані в Книзі Хроніки Ізраїлевих царів.
2KGS|15|27|П'ятдесятого й другого року Азарії, Юдиного царя, зацарював у Самарії над Ізраїлем Пеках, син Ремалії, на двадцять років.
2KGS|15|28|І робив він зло в Господніх очах, ні відступався від гріхів Єровоама, Неватового сина, що вводив у гріх Ізраїля.
2KGS|15|29|За днів Пекаха, Ізраїлевого царя, прийшов Тіґлат-Піл'есер, цар асирійський, взяв Іййона, і Авел-Бет-Мааху, і Йоноаха, і Кедеша, і Хацора, і Ґілеада, і Ґаліла, увесь край Нефталимів, та й вигнав їх до Асирії.
2KGS|15|30|А Осія, син Елин, склав змову на Пекаха, сина Ремалії, і вдарив його та й убив його, і зацарював замість нього двадцятого року Йотама, Уззійїного сина.
2KGS|15|31|А решта діл Пекаха та все, що він зробив, ото вони написані в Книзі Хроніки Ізраїлевих царів.
2KGS|15|32|Другого року Пекаха, сина Ремалії, Ізраїлевого царя, зацарював Йотам, син Уззійї, Юдиного царя.
2KGS|15|33|Він був віку двадцяти й п'яти років, коли зацарював, і шістнадцять літ царював в Єрусалимі. А ім'я його матері Єруша, Садокова дочка.
2KGS|15|34|І робив він угодне в Господніх очах, усе, що робив був його батько Уззійя, робив він.
2KGS|15|35|Тільки пагірки не були знищені, народ іще приносив жертви та кадив на пагірках. Він збудував горішню браму Господнього дому.
2KGS|15|36|А решта діл Йотама та все, що він зробив, ото вони написані в Книзі Хроніки Юдиних царів.
2KGS|15|37|За тих днів зачав Господь посилати на Юду Реціна, сирійського царя, та Пекаха, сина Ремалії.
2KGS|15|38|І спочив Йотам із своїми батьками, і був похований з батьками своїми в Місті Давида, свого батька, а замість нього зацарював син його Ахаз.
2KGS|16|1|Сімнадцятого року Пекаха, сина Ремалії, зацарював Ахаз, син Йотама, Юдиного царя.
2KGS|16|2|Ахаз був віку двадцяти літ, коли він зацарював, і царював в Єрусалимі шістнадцять років, і не робив угодного в очах Господа, Бога свого, як батько його Давид.
2KGS|16|3|І ходив він дорогою Ізраїлевих царів, і навіть сина свого провів через огонь для Молоха, за гидотою тих народів, що Господь вигнав їх перед Ізраїлевими синами.
2KGS|16|4|І приносив він жертву та кадив на пагірках, і на згір'ях, та під усяким зеленим деревом.
2KGS|16|5|Тоді прийшов Рецін, сирійський цар, та Пеках, син Ремалії, Ізраїлів цар, на війну до Єрусалиму. І облягли вони Ахаза, та не змогли звоювати.
2KGS|16|6|Того часу Рецін, сирійський цар, вернув Едомові Елата, і вигнав юдеїв з Елоту. І едомляни прибули до Елату, й осілися там, і живуть тут аж до цього дня.
2KGS|16|7|І послав Ахаз послів до Тіґлат-Пелесера, асирійського царя, говорячи: Я твій раб та син твій, вийди й спаси мене з руки сирійського царя та з руки царя Ізраїлевого, що повстають на мене.
2KGS|16|8|І взяв Ахаз срібло та золото, знайдене в Господньому домі та в скарбницях дому царевого, і послав дарунка до асирійського царя.
2KGS|16|9|І послухав його асирійський цар. І пішов асирійський цар на Дамаск і взяв його, а його мешканців вигнав до Кіру, а Реціна вбив.
2KGS|16|10|І пішов цар Ахаз назустріч Тіґлат-Піл'есера, асирійського царя, до Дамаску, і побачив дамаського жертівника. І послав цар Ахаз до священика Урії подобу жертівника та взір його всієї його будови.
2KGS|16|11|І збудував священик Урія жертівника, як усе, що послав був цар Ахаз із Дамаску, так зробив священик Урія до приходу царя Ахаза з Дамаску.
2KGS|16|12|І прибув цар із Дамаску, і побачив цар того жертівника, і приступив цар до жертівника, і приніс на ньому жертву.
2KGS|16|13|І спалив він своє цілопалення та свою жертву хлібну, і вилив свою ливну жертву, і покропив кров'ю своїх мирних жертов того жертівника.
2KGS|16|14|А мідяного жертівника, що перед Господнім лицем, він переставив із переднього боку храму, з-поміж жертівника та з-поміж Господнього дому, і поставив його на бік жертівника на північ.
2KGS|16|15|І наказав цар Ахаз священикові Урії, говорячи: На великому жертівнику пали ранішнє цілопалення та вечірню хлібну жертву, і цілопалення цареве та хлібну його жертву, і цілопалення всього народу Краю та хлібну їхню жертву, і їхні ливні жертви. І всю кров цілопалення та всю кров жертви покропиш на нього. А щодо мідяного жертівника, то я розважу.
2KGS|16|16|І зробив священик Урія все так, як наказав був цар Ахаз.
2KGS|16|17|А цар Ахаз повідрубував рами підстав, і відсунув із них умивальницю, і зняв море з мідяних волів, що під ним, і поставив його на камінну підлогу.
2KGS|16|18|І закритий суботній перехід, що збудували при храмі, і зовнішній царський вхід він обернув до Господнього дому задля асирійського царя.
2KGS|16|19|А решта діл Ахаза, що він зробив, ото вони написані в Книзі Хроніки Юдиних царів.
2KGS|16|20|І спочив Ахаз із батьками своїми, і був похований з батьками своїми в Давидовому Місті, а замість нього зацарював син його Хізкійя.
2KGS|17|1|Дванадцятого року Ахаза, Юдиного царя, зацарював над Ізраїлем у Самарії Осія, син Елин, на дев'ять років.
2KGS|17|2|І робив він зле в Господніх очах, тільки не так, як ті Ізраїлеві царі, що були перед ним.
2KGS|17|3|На нього вийшов Салманасар, цар асирійський, і Осія став йому за раба, і давав йому данину.
2KGS|17|4|Та асирійський цар знайшов в Осії змову, що він посилав послів до Со, єгипетського царя, та не приносив асирійському цареві данини, як рік-у-рік те робив був. І замкнув його асирійський цар, і зв'язав його в в'язничому домі.
2KGS|17|5|І вийшов асирійський цар на ввесь Край, і прийшов до Самарії, й облягав її три роки.
2KGS|17|6|Дев'ятого року Осії асирійський цар здобув Самарію, та й вигнав Ізраїля до Асирії, і осадив їх у Халаху, і в Хаворі над річкою Ґозан, і в містах Мідії.
2KGS|17|7|І сталося, коли Ізраїлеві сини грішили проти Господа, Бога свого, що випровадив їх з єгипетського краю з руки фараона, єгипетського царя, і боялися інших богів,
2KGS|17|8|і ходили уставами тих народів, що Господь повиганяв їх перед Ізраїлевими синами, та Ізраїлевих царів, які вони встановили,
2KGS|17|9|а Ізраїлеві сини вимишляли на Господа, Бога свого, слова, що не були слушні, і будували собі пагірки по всіх своїх містах, від вартової башти аж до твердинного міста,
2KGS|17|10|і ставили собі стовпи для богів та Астарти на кожному високому взгір'ї та під усяким зеленим деревом,
2KGS|17|11|і кадили там на всіх пагірках, як ті люди, що Господь повиганяв перед ними, і робили злі речі, щоб гнівити Господа,
2KGS|17|12|і служили бовванам, про яких Господь говорив їм: Не будете робити цієї речі,
2KGS|17|13|то Господь засвідчив в Ізраїлі та в Юді через усіх Своїх пророків та всіх прозорливців, говорячи: Верніться з ваших злих доріг, і додержуйте Моїх заповідей, уставів Моїх, згідно зо всім Законом, якого Я наказав був вашим батькам, і якого послав до вас через Моїх рабів пророків.
2KGS|17|14|Та не слухали вони, і робили твердою свою шию, як шия їхніх батьків, що не вірили в Господа, Бога свого.
2KGS|17|15|І нехтували вони постанови Його, і заповіта Його, що склав з їхніми батьками, і свідоцтва Його, що засвідчив на них, і пішли за гидотою й марнотами, та за народами, що були навколо них, про яких Господь наказав був їм не робити, як вони.
2KGS|17|16|І полишили вони всі заповіді Господа, Бога свого, і зробили собі литого боввана, двох телят, і зробили Астарту, і вклонялися всьому небесному військові та служили Ваалові.
2KGS|17|17|І вони переводили через огонь своїх синів та дочок своїх, і чарували чарами, і ворожили, і віддавалися робити зло в Господніх очах, щоб гнівити Його.
2KGS|17|18|І сильно розгнівався Господь на Ізраїля, і відкинув їх від Свого лиця, не позостало нікого, тільки саме Юдине плем'я.
2KGS|17|19|Та й Юда не додержував заповідей Господа, Бога свого, і ходили вони Ізраїлевими постановами, які вони встановили.
2KGS|17|20|І відвернувся Господь від усього Ізраїлевого насіння, і впокоряв їх, і давав їх у руку грабіжників, аж поки не кинув їх від лиця Свого,
2KGS|17|21|бо Ізраїль розірвав з Давидовим домом, і вони зробили царем Єровоама, Неватового сина, а Єровоам відвернув Ізраїля від Господа, і вводив їх у великий гріх.
2KGS|17|22|І ходили Ізраїлеві сини в усіх Єровоамових гріхах, які він робив, не відступалися з того,
2KGS|17|23|аж поки Господь не відкинув Ізраїля від лиця Свого, як говорив був через усіх Своїх рабів пророків. І пішов Ізраїль на вигнання з своєї землі до Асирії, і він там аж до цього дня.
2KGS|17|24|І спровадив асирійський цар людей з Вавилону, і з Кути, і з Авви, і з Гамоту, і з Сефарваїму, й оселив по містах Самарії замість Ізраїлевих синів. І посіли вони Самарію, й осілися по містах її.
2KGS|17|25|І сталося, на початку пробування їх там не боялися вони Господа, і Господь послав на них левів, і вони нищили їх.
2KGS|17|26|І сказали вони до асирійського царя, говорячи: Ті люди, яких ти вигнав та оселив по містах Самарії, не знають прав Бога цього Краю, і Він послав на них оцих левів, і ось вони нищать їх, бо вони не знають права Бога цього Краю.
2KGS|17|27|І наказав асирійський цар, говорячи: Відведіть туди одного зо священиків, яких вигнали звідти, і підуть, і осядуть там, і він навчатиме їх права Бога цього краю.
2KGS|17|28|І прибув один із священиків, яких вигнали з Самарії, й осівся в Бет-Елі, і він навчав їх, як мають боятися Господа.
2KGS|17|29|Та крім того кожен народ робив свого бога, і ставили їх у пагірковому місці, що робили попередні самаряни, кожен народ по своїх містах, де вони сиділи.
2KGS|17|30|А вавилоняни зробили Сукот-Бенота, а кутяни зробили Нереґала, а гаматяни зробили Ашіму,
2KGS|17|31|а авв'яни зробили Нівхаза та Тартака, а мешканці Сефарваїму палили синів своїх ув огні Адраммелехові й Анаммелехові, сефарваїмським богам.
2KGS|17|32|І при тому вони боялися Господа, і настановили собі з-серед себе священиків пагірків, і вони приносили їм жертви в пагірковому місці.
2KGS|17|33|Вони боялися Господа, і богам своїм служили за правом тих народів, звідки повиганяли їх.
2KGS|17|34|Аж до цього дня вони роблять за колишнім правом, вони не бояться Господа, і не роблять за уставами своїми та за правом своїм, ані за Законом, ані за заповіддю, як наказав був Господь синам Якова, якому дав ім'я Ізраїля.
2KGS|17|35|І склав Господь із ними заповіта, і наказав їм, говорячи: Не будете боятися інших богів, і не будете вклонятися їм, і не будете служити їм, і не будете приносити жертов їм,
2KGS|17|36|а тільки Господа, що вивів вас із єгипетського краю великою силою та витягненим раменом, Його будете боятися, і Йому будете вклонятися, і Йому будете приносити жертви.
2KGS|17|37|І устави, і права, і Закона, і заповідь, які написав вам, будете додержувати, щоб виконувати по всі дні, а богів інших не будете боятися.
2KGS|17|38|А заповіта, що Я склав із вами, не забудете, і не будете боятися інших богів,
2KGS|17|39|а тільки Господа, Бога вашого, будете боятися, і Він вирятує вас із руки всіх ваших ворогів.
2KGS|17|40|Та не послухали вони, бо все робили за своїм попереднім звичаєм.
2KGS|17|41|І ті народи все боялися Господа, але служили бовванам своїм. Так само сини їхні та сини їхніх синів, як робили батьки їхні, так роблять вони аж до цього дня.
2KGS|18|1|І сталося третього року Осії, сина Елиного, Ізраїлевого царя, зацарював Єзекія, син Ахазів, цар Юдин.
2KGS|18|2|Він був віку двадцяти й п'яти літ, коли зацарював, і царював в Єрусалимі двадцять і дев'ять літ. А ім'я його матері Аві, дочка Захарія.
2KGS|18|3|І робив він угодне в Господніх очах, усе так, як робив був його батько Давид.
2KGS|18|4|Він понищив пагірки, і поламав стовпи для богів, і стяв Астарту, і розбив мідяного змія, якого зробив був Мойсей, бо аж до цих днів Ізраїлеві сини все кадили йому й кликали його: Нехуштан.
2KGS|18|5|Він надіявся на Господа, Бога Ізраїля, і такого, як він, не було між усіма царями Юдиними, ані між тими, що були перед ним.
2KGS|18|6|І міцно тримався він Господа, не відступався від Нього, і додержував заповіді Його, що наказав був Господь Мойсеєві.
2KGS|18|7|І був Господь із ним, у всьому, куди він ходив, він мав поводження. І збунтувався він на асирійського царя, і не служив йому.
2KGS|18|8|Він побив филистимлян аж до Аззи та границі її від вартової башти аж до твердинного міста.
2KGS|18|9|І сталося четвертого року царя Єзекії, це сьомий рік Осії, Елиного сина, Ізраїлевого царя, пішов Салманасар, цар асирійський, на Самарію, та й обліг її.
2KGS|18|10|І здобув він її по трьох роках: шостого року Єзекії, це дев'ятий рік Осії, Ізраїлевого царя, була здобута Самарія.
2KGS|18|11|І вигнав асирійський цар Ізраїля до Асирії, і попровадив їх у Халах, і в Хавор, над річку Ґазан, та до мідійських міст.
2KGS|18|12|Це за те, що не слухалися вони голосу Господа, Бога свого, і переступали заповіта Його; усього, що наказав був Мойсей, раб Господній, вони ані не слухали, ані не робили.
2KGS|18|13|А чотирнадцятого року царя Єзекії прийшов Санхерів, цар асирійський, на всі укріплені Юдині міста, та й захопив їх.
2KGS|18|14|І послав Єзекія, цар Юдин, до царя асирійського, до Лахішу, говорячи: Згрішив я! Відійди від мене, а що накладеш на мене, понесу. І наклав асирійський цар на Єзекію, Юдиного царя, три сотні талантів срібла та тридцять талантів золота.
2KGS|18|15|І віддав Єзекія все срібло, знайдене в Господньому домі та в царевих скарбницях.
2KGS|18|16|Того часу Єзекія відрубав золото з дверей Господнього дому та зо стовпів, що покрив був Єзекія, Юдин цар, золотом, і дав його асирійському цареві.
2KGS|18|17|А асирійський цар послав із Лахішу до царя Єзекії головного командувача, і великого євнуха та великого чашника з великим військом до Єрусалиму. І пішли вони, і прийшли та й стали над водотягом горішнього ставу, що на битій дорозі до поля Валюшників.
2KGS|18|18|І кликнули вони до царя, і до них вийшов Еліяким, син Хілкійї, начальник палати, і писар Шевна, та Йоах, син Асафів, канцлер.
2KGS|18|19|І сказав до них великий чашник: Скажіть Єзекії: Отак сказав великий цар, цар асирійський: Що це за надія, на яку ти надієшся?
2KGS|18|20|Чи думаєш ти, що слово уст, то вже рада та сила до війни? На кого тепер надієшся, що збунтувався проти мене?
2KGS|18|21|Тепер оце ти надієшся собі опертися на оту поламану очеретину, на Єгипет, що коли хто опирається на неї, то вона входить у долоню йому й продірявлює її. Отакий фараон, цар єгипетський, для всіх, хто надіється на нього.
2KGS|18|22|А коли ви скажете мені: Ми надіємось на Господа, Бога нашого, то чи ж Він не Той, що Єзекія понищив пагірки Його та жертівники Його, і сказав Юді та Єрусалимові: перед оцим тільки жертівником будете вклонятися в Єрусалимі?
2KGS|18|23|А тепер піди в заклад із моїм паном, асирійським царем, і я дам тобі дві тисячі коней, якщо ти зможеш собі дати на них верхівців.
2KGS|18|24|І як же ти проженеш хоч одного намісника з найменших слуг мого пана? А ти собі надієшся на Єгипет ради колесниць та верхівців!
2KGS|18|25|Тепер же, чи без Господа прийшов я на це місце, щоб знищити його? Господь сказав був мені: Піди на той край та знищ його!
2KGS|18|26|І сказав Еліяким, син Хілкійї, і Шевна та Йоах до великого чашника: Говори до своїх рабів по-арамейському, бо ми розуміємо, і не говори з нами по-юдейському в слух тих людей, що на мурі.
2KGS|18|27|І сказав до них великий чашник: Чи пан мій послав мене говорити ці слова до твого пана та до тебе? Хіба не до цих людей, що сидять на мурі, щоб із вами їсти свій кал та пити свою сечу?
2KGS|18|28|І став великий чашник, і кликнув гучним голосом по-юдейському, і говорив і сказав: Послухайте слово великого царя, царя асирійського:
2KGS|18|29|Так сказав цар: Нехай не дурить вас Єзекія, бо він не зможе врятувати вас від руки його!
2KGS|18|30|І нехай не запевняє вас Єзекія Господом, говорячи: Рятуючи, врятує вас Господь, і не буде дано цього міста в руку царя асирійського.
2KGS|18|31|Не слухайте Єзекії, бо так сказав цар асирійський: Примиріться зо мною, та й вийдіть до мене, та й їжте кожен свій виноград та кожен фіґу свою, і пийте кожен воду зо своєї копанки,
2KGS|18|32|аж поки я не прийду й не візьму вас до краю такого ж, як ваш Край, до краю збіжжя та виноградного соку, до краю хліба та виноградників, до краю оливки, оливного соку та меду, щоб ви жили й не вмирали! І не слухайте Єзекії, коли він намовляє вас, говорячи: Господь порятує нас!
2KGS|18|33|Чи справді врятували боги тих народів, кожен свій край від руки асирійського царя?
2KGS|18|34|Де боги Гамату та Арпаду? Де боги Сефарваїму, Гени та Івви? Чи врятували вони Самарію від моєї руки?
2KGS|18|35|Котрий з-поміж усіх богів цих країв урятував свій край від моєї руки, то невже ж Господь урятує Єрусалим від моєї руки?
2KGS|18|36|І мовчав той народ, і не відповів йому ані слова, бо це був наказ царя, що сказав: Не відповідайте йому!
2KGS|18|37|І прийшов Еліяким, син Хілкійї, начальник палати, і писар Шевна, і Йоах, Асафів син, канцлер, із роздертими шатами, до Єзекії, і донесли йому слова великого чашника.
2KGS|19|1|І сталося, як почув це цар Єзекія, то роздер свої шати та накрився веретою, і ввійшов до Господнього дому.
2KGS|19|2|І послав він Еліякима, начальника палати, і писаря Шевну, та старших із священиків, покритих веретами, до пророка Ісаї, Амосового сина.
2KGS|19|3|І сказали вони до нього: Так сказав Єзекія: Цей день це день горя й картання та наруги! Бо підійшли діти аж до виходу утроби, та немає сили породити!
2KGS|19|4|Може почує Господь, Бог твій, всі слова великого чашника, що його послав асирійський цар, пан його, на образу Живого Бога, і Господь, Бог твій, покарає за слова, які чув, а ти принесеш молитву за рештку, що ще знаходиться.
2KGS|19|5|І прийшли раби царя Єзекії до Ісаї.
2KGS|19|6|І сказав їм Ісая: Так скажете вашому панові: Так сказав Господь: Не бійся тих слів, що почув ти, якими ображали Мене слуги асирійського царя!
2KGS|19|7|Ось Я дам в нього духа, і він почує звістку, і вернеться до свого краю. І Я вражу його мечем у його краї.
2KGS|19|8|І вернувся великий чашник, і знайшов асирійського царя, що воював проти Лівни, бо почув, що той рушив із Лахішу.
2KGS|19|9|А коли він почув про Тіргаку, царя етіопського, таке: Ось він вийшов воювати з тобою! то вернувся, і послав послів до Єзекії, говорячи:
2KGS|19|10|Так скажете до Єзекії, Юдиного царя, говорячи: Нехай не зводить тебе Бог твій, що ти надієшся на Нього, кажучи: Не буде даний Єрусалим у руку асирійського царя.
2KGS|19|11|Ось ти чув, що зробили асирійські царі всім краям, щоб учинити їх закляттям, а ти будеш урятований?
2KGS|19|12|Чи врятували їх боги тих народів, яких понищили батьки мої: Гозана, і Харана, і Рецефа, і синів Едена, що в Телассарі?
2KGS|19|13|Де він, цар Гамату, і цар Арпаду, і цар міста Сефарваїму, Гени та Івви?
2KGS|19|14|І взяв Єзекія ті листи з руки послів, і прочитав їх, і ввійшов у Господній дім. І Єзекія розгорнув одного листа перед Господнім лицем.
2KGS|19|15|І Єзекія молився перед Господнім лицем і сказав: Господи, Боже Ізраїлів, що сидиш на херувимах! Ти Той єдиний Бог для всіх царств землі, Ти створив небеса та землю!
2KGS|19|16|Нахили, Господи, ухо Своє та й почуй! Відкрий, Господи, очі Свої та й побач, і почуй слова Санхеріва, що прислав ображати Живого Бога!
2KGS|19|17|Справді, Господи, асирійські царі попустошили ті народи та їхній край.
2KGS|19|18|І кинули вони їхніх богів на огонь, бо не боги вони, а тільки чин людських рук, дерево та камінь, і понищили їх.
2KGS|19|19|А тепер, Господи, Боже наш, спаси нас від руки його, і нехай знають усі царства землі, що Ти Господь, Бог єдиний!
2KGS|19|20|І послав Ісая, Амосів син, до Єзекії, говорячи: Так сказав Господь, Бог Ізраїлів: Я почув те, про що ти молився до Мене, про Санхеріва, царя асирійського.
2KGS|19|21|Ось те слово, яке Господь говорив про нього: Гордує тобою, сміється із тебе дівиця, сіонська дочка, вслід тобі головою хитає дочка Єрусалиму!
2KGS|19|22|Кого лаяв ти та ображав, і на кого повищив ти голос та вгору підніс свої очі? На Святого Ізраїлевого!
2KGS|19|23|Через послів своїх Господа ти ображав та казав: Із безліччю своїх колесниць я вийшов на гори високі, на боки Ливану, і позрубую кедри високі його, добірні його кипариси, і вийду аж на вершок його на нічліг, у гущину його саду.
2KGS|19|24|Я копаю та п'ю чужу воду, і стопою своєї ноги повисушую я всі єгипетські ріки!
2KGS|19|25|Хіба ти не чув, що віддавна зробив Я оце, що за днів стародавніх Я це був створив? Тепер же спровадив Я це, що ти нищиш міста поукріплювані, на купу румовищ обертаєш їх...
2KGS|19|26|А мешканці їхні безсилі, настрашені та побентежені. Вони стали, як зілля оте польове, мов трава зеленіюча, як трава на дахах, як попалене збіжжя, яке не доспіло...
2KGS|19|27|І сидіння твоє, і твій вихід та вхід твій Я знаю, і твоє проти Мене обурення.
2KGS|19|28|За твоє проти Мене обурення, що гординя твоя надійшла до ушей Моїх, то на ніздрі твої Я сережку привішу, а вудило Моє в твої уста, і тебе поверну Я тією дорогою, якою прийшов ти!
2KGS|19|29|А оце тобі знак: їжте цього року збіжжя самосійне, а другого року саморосле, а третього року сійте та жніть, і садіть виноградники, та й їжте їх плід.
2KGS|19|30|А врятоване Юдиного дому, що лишилося, пустить коріння додолу, і свого плода дасть угору.
2KGS|19|31|Бо з Єрусалиму вийде позостале, а рештки від гори Сіону. Ревність Господа Саваота зробить це!
2KGS|19|32|Тому так сказав Господь про асирійського царя: Він не ввійде до міста оцього, і туди він не кине стріли, і щитом її не попередить, і вала на нього не висипле!
2KGS|19|33|Якою дорогою прийде, то нею повернеться, у місто ж оце він не ввійде, говорить Господь!
2KGS|19|34|І це місто Я обороню на спасіння його ради Себе та ради Давида, Мойого раба!
2KGS|19|35|І сталося тієї ночі, і вийшов Ангол Господній, і забив в асирійському таборі сто й вісімдесят і п'ять тисяч. І повставали вони рано вранці, аж ось усі мертві трупи!...
2KGS|19|36|А Санхерів, асирійський цар, рушив та й пішов, і вернувся й осівся в Ніневії.
2KGS|19|37|І сталося, коли він молився в домі Нісроха, свого бога, то Адраммелех та Шар'ецер убили його мечем, а самі втекли до краю Арарат. А замість нього зацарював син його Есар-Хаддон.
2KGS|20|1|Тими днями смертельно захворів був Єзекія. І прийшов до нього Ісая, Амосів син, пророк, і сказав до нього: Так сказав Господь: Заряди своїм домом, бо ти вмреш, а не видужаєш.
2KGS|20|2|А той відвернув обличчя своє до стіни, і помолився до Господа, говорячи:
2KGS|20|3|О, Господи, згадай же, що я ходив перед лицем Твоїм правдою та цілим серцем, і робив я добре в очах Твоїх. І заплакав Єзекія ревним плачем...
2KGS|20|4|І сталося, Ісая не вийшов ще з середини міста, а до нього було Господнє слово, говорячи:
2KGS|20|5|Вернися, і скажеш до Єзекії, володаря Мого народу: Так сказав Господь, Бог батька твого Давида: Почув Я молитву твою, побачив Я сльозу твою! Ось Я вилікую тебе, третього дня зійдеш ти до Господнього дому!
2KGS|20|6|І до днів твоїх Я додам п'ятнадцять літ, і з руки асирійського царя врятую тебе та це місто, й обороню це місто ради Себе та ради раба Свого Давида.
2KGS|20|7|А Ісая сказав: Візьміть грудку фіґ. І взяли й поклали на того гнояка, і він видужав...
2KGS|20|8|І сказав Єзекія до Ісаї: Який знак, що Господь мене вилікує, і що я третього дня зійду до Господнього дому?
2KGS|20|9|І сказав Ісая: Ось тобі знак той від Господа, що Господь зробить ту річ, про яку говорив: Чого хочеш, щоб пішла тінь уперед на десять ступенів, чи щоб вернулася на десять ступенів?
2KGS|20|10|І сказав Єзекія: Легко тіні похилитися вперед на десять ступенів; ні, а нехай тінь вернеться назад на десять ступенів!
2KGS|20|11|І кликнув пророк Ісая до Господа, і Він завернув тінь на ступенях, де вона спускалася на ступені Ахазові, на десять ступенів...
2KGS|20|12|Того часу послав Беродах-Бал'адан, син Бал'аданів, вавилонський цар, листа та дарунка до Єзекії, бо прочув був, що Єзекія захворів.
2KGS|20|13|І вислухав їх Єзекія, і показав їм усю скарбницю свою, і срібло, і золото, і пахощі, і добру оливу, і всю зброївню свою, і все, що знаходилося в його скарбницях. Не було речі, якої не показав би їм Єзекія в домі своїм та в усім володінні своїм.
2KGS|20|14|І прийшов пророк Ісая до царя Єзекії та й сказав до нього: Що говорили ці люди? І звідки вони прийшли до тебе? А Єзекія сказав: Вони прийшли з далекого краю, з Вавилону.
2KGS|20|15|І той сказав: Що вони бачили в домі твоїм? І Єзекія сказав: Усе, що в домі моїм, вони бачили, не було речі, якої не показав би я їм у скарбницях своїх.
2KGS|20|16|І сказав Ісая до Єзекії: Послухай Господнього слова:
2KGS|20|17|Ось приходять дні, і все, що в домі твоєму, і що були зібрали батьки твої аж до цього дня, буде винесене до Вавилону. Нічого не позостанеться, говорить Господь!
2KGS|20|18|А з синів твоїх, що вийдуть із тебе, яких ти породиш, декого заберуть, і вони будуть євнухами в палатах вавилонського царя!
2KGS|20|19|І сказав Єзекія до Ісаї: Добре Господнє слово, яке ти сказав! І подумав собі: Так, мир та безпека буде за моїх днів!
2KGS|20|20|А решта діл Єзекії та вся лицарськість його, і як він зробив става та водотяга, і впровадив воду до міста, ото вони написані в Книзі Хроніки Юдиних царів.
2KGS|20|21|І спочив Єзекія зо своїми батьками, а замість нього зацарював син його Манасія.
2KGS|21|1|Манасія був віку дванадцяти літ, коли він зацарював, і царював в Єрусалимі п'ятдесят і п'ять літ. А ім'я його матері Хевці-Ваг.
2KGS|21|2|І робив він зло в Господніх очах, за гидотою тих народів, яких Господь повиганяв з-перед обличчя Ізраїлевих синів.
2KGS|21|3|І він знову побудував пагірки, що їх винищив був його батько Єзекія, і понаставляв жертівників Ваалові, і зробив Астарту, як зробив був Ахав, Ізраїлів цар, і вклонявся всім небесним світилам та служив їм.
2KGS|21|4|І побудував він жертівники в Господньому домі, про якого сказав був Господь: В Єрусалимі покладу Я Ім'я Своє!
2KGS|21|5|І побудував він жертівники для всіх небесних світил на обох подвір'ях Господнього дому.
2KGS|21|6|І він перепровадив свого сина через огонь, і гадав, і ворожив, і настановив викликувачів духів померлих та духів віщих, і багато робив зла в очах Господа, щоб гнівити Його.
2KGS|21|7|І поставив він боввана Астарти, якого зробив, у домі, про якого Господь сказав був до Давида та до сина його Соломона: У цьому домі та в Єрусалимі, що його Я вибрав зо всіх Ізраїлевих племен, покладу Я Ім'я Своє навіки!
2KGS|21|8|І більше не мандруватиме Ізраїлева нога з тієї землі, яку Я дав їхнім батькам, якщо тільки вони будуть пильнувати робити все так, як наказав Я їм, та ввесь Закон, що наказав їм Мій раб Мойсей.
2KGS|21|9|Та не послухалися вони. І Манасія звів їх до того, щоб робити гірше від тих народів, яких Господь вигубив з-перед обличчя Ізраїлевих синів.
2KGS|21|10|І говорив Господь через Своїх рабів пророків, кажучи:
2KGS|21|11|За те, що Манасія, цар Юдин, зробив ці гидоти, учинив гірше від усього, що робили були амореяни, що були перед ним, і ввів у гріх також Юду божками своїми,
2KGS|21|12|тому так сказав Господь, Бог Ізраїлів: Ось Я наводжу таке зло на Єрусалим та на Юду, що в кожного, хто почує про це, задзвенить в обох вухах!...
2KGS|21|13|І протягну Я на Єрусалим мірку Самарії, та вагу Ахавого дому, і витру Єрусалим, як витирають миску: витер і перевернув її догори дном!
2KGS|21|14|І Я покину останок наділу Мого, і дам їх у руку їхнім ворогам, і вони будуть на грабіж та на здобич для всіх їхніх ворогів,
2KGS|21|15|тому, що вони робили зло в Моїх очах, і все гнівили Мене від дня, коли вийшли їхні батьки з Єгипту, й аж до дня цього...
2KGS|21|16|А також Манасія пролив дуже багато невинної крови, аж наповнив нею Єрусалим від входу до входу, окрім свого гріха, що ввів у гріх Юду, щоб чинити зле в Господніх очах.
2KGS|21|17|А решта діл Манасії, та все, що він зробив, і гріх його, яким він грішив, ото вони написані в Книзі Хроніки Юдиних царів.
2KGS|21|18|І спочив Манасія з батьками своїми, і був похований в садку свого дому, в Уззиному садку, а замість нього зацарював син його Амон.
2KGS|21|19|Амон був віку двадцяти й двох років, коли він зацарював, і царював він в Єрусалимі два роки. А ім'я його матері Мешуллемет, дочка Харуца з Йотви.
2KGS|21|20|І робив він зло в Господніх очах, як робив його батько Манасія.
2KGS|21|21|І ходив він усією тією дорогою, якою ходив його батько, і служив тим бовванам, яким служив батько його, і вклонявся їм.
2KGS|21|22|І покинув він Господа, Бога батьків своїх, і не ходив Господньою дорогою.
2KGS|21|23|І вчинили змову слуги Амона на нього, і вбили царя в його домі.
2KGS|21|24|Та народ Краю перебив усіх змовників на царя Амона. І народ настановив царем Краю замість нього сина його Йосію.
2KGS|21|25|А решта діл Амона, усе, що робив він, ото вони написані в Книзі Хроніки Юдиних царів.
2KGS|21|26|І поховали його в його гробі в Уззиному садку, а замість нього зацарював син його Йосія.
2KGS|22|1|Йосія був віку восьми літ, коли він зацарював, і царював в Єрусалимі тридцять і один рік. А ім'я його матері Єдида, дочка Адаї з Боцкату.
2KGS|22|2|І робив він угодне в Господніх очах, і ходив усією дорогою свого батька Давида, і не вступався ані праворуч, ані ліворуч.
2KGS|22|3|І сталося вісімнадцятого року царя Йосії, послав цар Шафана, сина Ацалії, Мешулламового сина, писаря, до Господнього дому, говорячи:
2KGS|22|4|Піди до Хілкійї, первосвященика, і нехай перелічить те срібло, що знесене до Господнього дому, що зібрали від народу сторожі порога.
2KGS|22|5|І нехай дадуть його на руку виконавцям роботи, поставленим у Господньому домі, а ті нехай дадуть його тим, хто працює в Господньому домі, щоб направляти ушкодження храму,
2KGS|22|6|теслярам, і будівничим, і мулярам, щоб купувати дерево та тесане каміння на направу храму.
2KGS|22|7|Тільки нехай не облічуються з ними про те срібло, що дане на їхню руку, бо чесно вони роблять.
2KGS|22|8|І сказав Хілкійя, первосвященик, до писаря Шафана: Я знайшов у Господньому домі Книгу Закону! І дав Хілкійя ту Книгу Шафанові, і той перечитав її.
2KGS|22|9|І ввійшов писар Шафан до царя, і приніс цареві вістку, і сказав: Раби твої висипали те срібло, що знайдене в домі, і дали його на руку виконавцям роботи, поставленим у Господньому домі.
2KGS|22|10|І доніс писар Шафан цареві, говорячи: Священик Хілкійя дав мені книгу. І Шафан перечитав її перед царем.
2KGS|22|11|І сталося, як цар почув слова Книги Закону, то роздер свої шати...
2KGS|22|12|І наказав цар священикові Хілкійї, і Ахікамові, Шафановому синові, і Ахборові, Міхаїному синові, і писареві Шафанові, і Асаї, царевому слузі, говорячи:
2KGS|22|13|Ідіть, зверніться до Господа про мене й про народ, та про всього Юду, про слова цієї знайденої книги. Великий бо гнів Господній, що запалився на нас за те, що батьки наші не слухалися слів цієї книги, щоб робити все, що написано про нас.
2KGS|22|14|І пішов священик Хілкійя, і Ахікам, і Ахбор, і Шафан, і Асая до пророчиці Хулди, жінки Шаллума, сина Тікви, сина Хархасового, сторожа шат, вона сиділа в Єрусалимі, на Новому Місті, і говорили до неї.
2KGS|22|15|А вона сказала до них: Так говорить Господь, Бог Ізраїлів: Скажіть чоловікові, що послав вас до мене:
2KGS|22|16|Так говорить Господь: Ось Я наведу лихо на оце місце та на мешканців його, усі слова тієї книги, що читав Юдин цар,
2KGS|22|17|за те, що вони покинули Мене, і кадили іншим богам, щоб гнівити Мене всім ділом своїх рук. І розпалився Мій гнів на це місце, і він не погасне!
2KGS|22|18|А Юдиному цареві, що послав вас звернутися до Господа, скажете йому так: Так говорить Господь, Бог Ізраїлів, ті слова, які ти чув:
2KGS|22|19|За те, що зм'якло твоє серце, і ти впокорився перед Господнім лицем, коли почув, що Я говорив про це місце та про мешканців його, що вони стануть спустошенням та прокляттям, і що ти роздер шати свої та плакав перед Моїм лицем, то Я також почув, говорить Господь.
2KGS|22|20|Тому то Я прилучу тебе до батьків твоїх, і ти будеш прилучений до гробів своїх у мирі, і очі твої не побачать усього того лиха, що Я наводжу на оце місце. І вони принесли цю вістку цареві.
2KGS|23|1|А цар послав, і зібрали до нього всіх старших Юди та Єрусалиму.
2KGS|23|2|І ввійшов до Господнього дому цар та кожен муж Юди, а з ним усі мешканці Єрусалиму, і священики, і пророки, і ввесь народ від малого й аж до великого, і він прочитав до їхніх ушей усі слова Книги Заповіту, знайденої в Господньому домі.
2KGS|23|3|І став цар на підвищенні, і склав заповіта перед Господнім лицем, щоб ходити за Господом та додержувати заповіді Його, і свідчення Його, і постанови Його всім серцем та всією душею, щоб виконати слова того заповіту, що написані в тій книзі. І ввесь народ пристав до заповіту.
2KGS|23|4|І наказав цар Хілкійї, великому священикові, й іншим священикам та сторожам порога, щоб повиносили з Господнього храму всі речі, зроблені для Ваала та для Астарти, та для всіх небесних світил. І він попалив їх поза Єрусалимом на кедронських полях, а їхній порох відніс до Бет-Елу.
2KGS|23|5|І він поскидав жерців, що їх понаставляли були Юдині царі, і що вони кадили на пагірках по Юдиних містах та в околицях Єрусалиму, і кадили для Ваала, і для сонця, і для місяця, і для планет, і для всіх небесних світил.
2KGS|23|6|І він виніс Астарту з Господнього дому поза Єрусалим до кедронської долини, та й спалив її в кедронській долині, і стер на порох, а її порох кинув на гроби звичайних людей.
2KGS|23|7|І він порозбивав доми культу блудодійників, що були при Господньому домі, де жінки ткали завісу для Астарти.
2KGS|23|8|І він випровадив усіх священиків з Юдиних міст, і опоганив пагірки, де священики кадили, від Ґеви аж до Беер-Шеви, і порозбивав пагірки брам, що були при вході брами Ісуса, зверхника міста, що ліворуч тому, хто входив до брами міста.
2KGS|23|9|Але священики пагірків не входили до Господнього жертівника в Єрусалимі, а тільки їли прісне серед своїх братів.
2KGS|23|10|І він опоганив місце ставлення на огні, що в долині Гінномового сина, щоб ніхто не переводив через огонь сина свого та дочку свою для Молоха.
2KGS|23|11|І він повідставляв коні, яких давали Юдині царі для сонця, від входу до Господнього дому, при кімнаті євнуха Нетан-Мелеха, що був у Парварімі, а колесниці сонця попалив ув огні.
2KGS|23|12|А жертівники, що були на даху Ахазової горниці, що поробили Юдині царі, та жертівники, що поробив Манасія на двох подвір'ях Господнього дому, цар порозбивав. І він звідти побіг, і кинув їхній порох до кедронського потоку.
2KGS|23|13|А пагірки, що навпроти Єрусалиму, праворуч гори Згуби, які побудував був Соломон, Ізраїлів цар, для Астарти, гидоти сидонської, і для Кемота, гидоти моавської, і для Мілкома, гидоти Аммонових синів, цар поопоганював.
2KGS|23|14|І він порозбивав стовпи для богів, і постинав посвячені дерева, а їхнє місце наповнив людськими кістками.
2KGS|23|15|А також жертівника, що в Бет-Елі, пагірка, що зробив був Єровоам, син Неватів, що ввів у гріх Ізраїля, також жертівника цього та цього пагірка він розбив, і спалив того пагірка та стер на порох, і Астарту спалив.
2KGS|23|16|І обернувся Йосія, та й побачив гроби, що були там на горі. І послав він, і позабирав кості з гробів, і попалив на жертівнику, і опоганив його, за словом Господнім, яке кликав був Божий чоловік, що прорікав оці речі.
2KGS|23|17|І сказав цар: Що це за надгробок, що я бачу? А люди того міста сказали йому: Це надгробок Божого чоловіка, що прийшов з Юдеї й прорік оці речі, які зробив ти на жертівнику в Бет-Елі.
2KGS|23|18|А він сказав: Дайте йому спокій, нехай ніхто не рухає костей його. І зберегли його кості, кості того пророка, що прийшов був із Самарії.
2KGS|23|19|А також усі доми пагірків, що по самарійських містах, що поробили були Ізраїлеві царі, щоб гнівити Господа, Йосія понищив, і зробив з ними те саме, що зробив у Бет-Елі.
2KGS|23|20|І порізав він усіх священиків пагірків, що були там, на жертівниках, і попалив на них людські кості, та й вернувся до Єрусалиму.
2KGS|23|21|І наказав цар усьому народові, говорячи: Справте Пасху для Господа, вашого Бога, як написано в оцій Книзі Заповіту.
2KGS|23|22|Бо не справлялася ця Пасха від днів суддів, що судили Ізраїля, по всі дні царів Ізраїлевих та царів Юдиних.
2KGS|23|23|І тільки вісімнадцятого року царя Йосії справлялася Пасха для Господа в Єрусалимі.
2KGS|23|24|А також викликачів духів померлих, і духів віщих, і домових божків, і бовванів, і всякі гидоти, що появилися в Юдинім краї та в Єрусалимі, повинищував Йосія, щоб поставити слова Закону, написані в книзі, що знайшов священик Хілкійя в Господньому домі.
2KGS|23|25|А такого царя, як він, не було перед ним, що навернувся б до Господа всім своїм серцем, і всією душею своєю, і всією силою своєю, за всім Мойсеєвим Законом, і по ньому не повставав такий, як він.
2KGS|23|26|Тільки не спинився Господь від ревности Свого великого гніву, яким запалився Його гнів на Юду за всі огірчення, якими гнівив Його Манасія.
2KGS|23|27|І сказав Господь: Також Юду відкину Я від лиця Свого, як відкинув Я Ізраїля, і відкину це місто, яке вибрав, Єрусалим, та цей храм, про який Я сказав: Ім'я Моє буде там!
2KGS|23|28|А решта діл Йосії та все, що він робив, ото вони написані в Книзі Хроніки Юдиних царів.
2KGS|23|29|За його днів пішов фараон Нехо, єгипетський цар, на асирійського царя, на річку Єфрат. І вийшов цар Йосія навпроти нього, та той убив його в Меґіддо, коли він побачив його...
2KGS|23|30|І його раби повезли його мертвого з Меґіддо, і привезли його до Єрусалиму, і поховали його в гробівці його. А народ Краю взяв Єгоахаза, сина Йосії, і помазали його, та й настановили його царем замість його батька.
2KGS|23|31|Єгоахаз був віку двадцяти й трьох літ, коли він зацарював, і царював в Єрусалимі три місяці. А ім'я його матері Хамуталь, дочка Єремії, з Лівни.
2KGS|23|32|І робив він зло в Господніх очах, усе так, як робили його батьки.
2KGS|23|33|І фараон Нехо зв'язав його в Рівлі, в гаматському краї, щоб він не царював в Єрусалимі, і наклав кару на цей край, сто талантів срібла та талант золота.
2KGS|23|34|А царем настановив фараон Нехо Ел'якима, сина Йосії, замість батька його Йосії, і змінив ім'я його на Єгояким. А Єгоахаза він узяв, і той прибув до Єгипту та й помер там.
2KGS|23|35|І Єгояким давав фараонові срібла та золота; тільки розклав це на Край, щоб давати те срібло на фараонів наказ, він стягав те срібло та золото з народу Краю за оцінкою землі кожного, щоб віддати фараонові Нехо.
2KGS|23|36|Єгояким був віку двадцяти й п'яти літ, коли він зацарював, і одинадцять років царював в Єрусалимі. А ім'я його матері Зевуда, дочка Педаї, з Руми.
2KGS|23|37|І робив він зло в Господніх очах, усе так, як робили батьки його.
2KGS|24|1|За його днів прийшов Навуходоносор, цар вавилонський, а Єгояким був йому три роки невільником, та потому збунтувався на нього.
2KGS|24|2|А Господь послав на нього орди халдеїв, і орди сирійські, і орди моавські, та орди синів Аммона. І він послав їх на Юду, щоб вигубити їх за словом Господа, що Він говорив через рабів Своїх пророків.
2KGS|24|3|Тільки на наказ Господа сталося це на Юду, щоб відкинути його від лиця Його за гріхи Манасії, за все, що він робив,
2KGS|24|4|а також за неповинну кров, яку він пролив, і наповнив Єрусалим неповинною кров'ю; і не хотів Господь простити.
2KGS|24|5|А решта Єгоякимових діл, та все, що він робив, ото вони описані в Книзі Хроніки Юдиних царів.
2KGS|24|6|І спочив Єгояким зо своїми батьками, а замість нього зацарював син його Єгояхін.
2KGS|24|7|І більше вже не виходив єгипетський цар зо свого краю, бо вавилонський цар забрав усе від Єгипетського потоку аж до річки Ефрату, усе, що належало єгипетському цареві.
2KGS|24|8|Єгояхін був віку вісімнадцяти літ, коли він зацарював, і царював в Єрусалимі три місяці. А ім'я його матері Нехушта, дочка Елнатана, з Єрусалиму.
2KGS|24|9|І робив він зло в Господніх очах, усе так, як робив його батько.
2KGS|24|10|Того часу прийшли до Єрусалиму раби Навуходоносора, царя вавилонського, і місто попало в облогу.
2KGS|24|11|І прийшов Навуходоносор, вавилонський цар, на місто, а його раби облягали його.
2KGS|24|12|І вийшов Єгояхін, цар Юдин, до вавилонського царя, він та мати його, і слуги його, і князі його, і євнухи його, і вавилонський цар узяв його восьмого року свого царювання.
2KGS|24|13|І позабирав він звідти всі скарби Господнього дому та скарби дому царевого, і повідрубував всі золоті речі, які поробив був Соломон, цар Ізраїлів, у Господньому храмі, як говорив Господь.
2KGS|24|14|І повиводив він увесь Єрусалим, і всіх князів, і всіх лицарів військових, десять тисяч пішло до неволі, і всіх теслів та ковалів. Не позоставив нікого, окрім нужденного народу Краю...
2KGS|24|15|І він вивів до Вавилону Єгояхіна та цареву матір, і царських жінок, і його євнухів, і видатних у Краї, усіх випровадив у неволю з Єрусалиму до Вавилону.
2KGS|24|16|І всіх військових, сім тисяч, і теслів та ковалів тисячу, усіх лицарів, що займалися війною, вивів їх вавилонський цар у неволю до Вавилону.
2KGS|24|17|А царем настановив вавилонський цар Маттанію, дядька Єгояхіна, замість нього, і перемінив ім'я його на Седекію.
2KGS|24|18|Седекія був віку двадцяти й одного року, коли він зацарював, і він царював в Єрусалимі одинадцять років. А ім'я його матері Хамуталь, дочка Єремії з Лівни.
2KGS|24|19|І робив він зло в Господніх очах, усе так, як робив був Єгояким.
2KGS|24|20|Бо за Господній гнів сталося це на Єрусалим та на Юду, і Він відкинув їх від Свого лиця. І Седекія збунтувався проти вавилонського царя.
2KGS|25|1|І сталося дев'ятого року його царювання, десятого місяця, десятого дня місяця, прийшов Навуходоносор, цар вавилонський, він та все військо його, на Єрусалим, і розтаборився проти нього, і побудували проти нього вала навколо.
2KGS|25|2|І було місто в облозі аж до одинадцятого року царя Седекії.
2KGS|25|3|Дев'ятого дня місяця настав сильний голод у місті, і не було хліба для народу Краю.
2KGS|25|4|І пробитий був пролім у мурі міста, і всі вояки повтікали вночі дорогою брами між двома мурами, що при царському садку, бо халдеї були при місті навколо. А цар утік дорогою в степ.
2KGS|25|5|А халдейське військо погналося за царем, та й догнали його в єрихонських степах, а все його військо розпорошилося від нього.
2KGS|25|6|І схопили царя, і відвели його до вавилонського царя до Рівли, і там його той засудив.
2KGS|25|7|А синів Седекії зарізали на його очах, а очі Седекії він вибрав, і скував його двома мідяними кайданами, та й відвів його до Вавилону...
2KGS|25|8|А п'ятого місяця, сьомого дня місяця, це дев'ятнадцятий рік царя Навуходоносора, вавилонського царя, прийшов до Єрусалиму Невузар'адан, начальник царської сторожі, слуга вавилонського царя.
2KGS|25|9|І він спалив дім Господній та дім царевий, і всі доми в Єрусалимі, і кожен великий дім спалив огнем.
2KGS|25|10|І мури навколо Єрусалиму порозбивало все халдейське військо, що було з начальником царської сторожі.
2KGS|25|11|А решту народу, що позостався в місті, і тих, що перебігли до вавилонського царя, і решту простого люду повиганяв Невузар'адан, начальник царської сторожі.
2KGS|25|12|А з бідноти Краю начальник царської сторожі позоставив декого за винярів та за рільників.
2KGS|25|13|А мідяні стовпи, що в Господньому домі, і підстави, і мідяне море, що в Господньому домі, халдеї поламали, і віднесли їхню мідь до Вавилону.
2KGS|25|14|І горнята, і лопатки, і ножі, і ложки, і ввесь мідяний посуд, що вживається при службі, позабирали.
2KGS|25|15|І кадильниці, і чаші, усе, що було золоте забрав золото, а що було срібне срібло взяв начальник царської сторожі.
2KGS|25|16|Два стовпи, одне море та ті підстави, що Соломон поробив був для Господнього дому, не було й ваги для всіх цих речей!
2KGS|25|17|Вісімнадцять ліктів високість одного стовпа й одна мідяна маковиця, а високість маковиці три лікті, та мережка, і гранатові яблука на маковиці навколо, усе мідь. І для другого стовпа з мережкою так само.
2KGS|25|18|І начальник царської сторожі взяв Сераю, первосвященика, і Цефанію, другого священика, та трьох сторожів порога.
2KGS|25|19|А з міста взяв він одного євнуха, що був начальником над військовими, та п'ять чоловіка з тих, що бачать цареве обличчя, що були знайдені в місті, і писаря, зверхника військових відділів, що записував народ Краю до військових відділів, і шістдесят чоловіка з народу Краю, що знаходилися в місті.
2KGS|25|20|І позабирав їх Невузар'адан, начальник царської сторожі, і відвів їх до вавилонсього царя, до Рівли.
2KGS|25|21|І вдарив їх вавилонський цар, і повбивав їх у Рівлі, у гаматовому краї. І пішов Юда на вигнання з своєї землі.
2KGS|25|22|А народ, що позостався в Юдиному краї, якого позоставив Навуходоносор, вавилонський цар, то настановив над ним Ґедалію, сина Ахікама, Шафанового сина.
2KGS|25|23|І почули всі військові зверхники, вони та люди, що вавилонський цар настановив Ґедалію, то поприходили до Ґедалії до Міцпи і Ізмаїл, син Нетаніїн, і Йоханан, син Кареахів, і Серая, син нетофатянина Танхумета, і Яазанія, син маахатянина, вони та їхні люди.
2KGS|25|24|І присягнув Ґедалія їм та їхнім людям, і сказав їм: Не бійтеся бути підданими халдейцям, осядьте в Краї та служіть вавилонському цареві, і буде вам добре!
2KGS|25|25|І сталося сьомого місяця, прийшов Ізмаїл, син Нетанії, Елішамового сина, з царського насіння, та десять мужів із ним, і вдарили вони Ґедалію, і він помер, і юдеїв, і халдеїв, що були з ними в Міцпі.
2KGS|25|26|І знявся ввесь народ, від малого й аж до великого, та зверхники військ, і пішов до Єгипту, бо боявся халдеїв.
2KGS|25|27|І сталося тридцятого й сьомого року неволі Єгояхіна, Юдиного царя, дванадцятого місяця, двадцять сьомого дня місяця, Евіл-Меродах, цар вавилонський, у році свого зацарювання, змилувався над Єгояхіном, Юдиним царем, і вивів його з дому ув'язнення.
2KGS|25|28|І він говорив із ним ласкаво, і поставив трона його понад трона царів, що були з ним у Вавилоні.
2KGS|25|29|І змінив в'язничну одежу його, і він завжди їв хліб перед ним по всі дні свого життя.
2KGS|25|30|А їжа його, їжа стала, видавалася йому від царя, щоденне щоденно, по всі дні його життя.
