GEN|1|1|In principio creavit Deus caelum et terram.
GEN|1|2|Terra autem erat inanis et vacua, et tenebrae super faciem abyssi, et spiritus Dei ferebatur super aquas.
GEN|1|3|Dixitque Deus: " Fiat lux ". Et facta est lux.
GEN|1|4|Et vidit Deus lucem quod esset bona et divisit Deus lucem ac tenebras.
GEN|1|5|Appellavitque Deus lucem Diem et tenebras Noctem. Factumque est vespere et mane, dies unus.
GEN|1|6|Dixit quoque Deus: " Fiat firmamentum in medio aquarum et dividat aquas ab aquis ".
GEN|1|7|Et fecit Deus firmamentum divisitque aquas, quae erant sub firmamento, ab his, quae erant super firmamentum. Et factum est ita.
GEN|1|8|Vocavitque Deus firmamentum Caelum. Et factum est vespere et mane, dies secundus.
GEN|1|9|Dixit vero Deus: " Congregentur aquae, quae sub caelo sunt, in locum unum, et appareat arida ". Factumque est ita.
GEN|1|10|Et vocavit Deus aridam Terram congregationesque aquarum appellavit Maria. Et vidit Deus quod esset bonum.
GEN|1|11|Et ait Deus: " Germinet terra herbam virentem et herbam facientem semen et lignum pomiferum faciens fructum iuxta genus suum, cuius semen in semetipso sit super terram ". Et factum est ita.
GEN|1|12|Et protulit terra herbam virentem et herbam afferentem semen iuxta genus suum lignumque faciens fructum, qui habet in semetipso sementem secundum speciem suam. Et vidit Deus quod esset bonum.
GEN|1|13|Et factum est vespere et mane, dies tertius.
GEN|1|14|Dixit autem Deus: " Fiant luminaria in firmamento caeli, ut dividant diem ac noctem et sint in signa et tempora et dies et annos,
GEN|1|15|ut luceant in firmamento caeli et illuminent terram. Et factum est ita.
GEN|1|16|Fecitque Deus duo magna luminaria: luminare maius, ut praeesset diei, et luminare minus, ut praeesset nocti, et stellas.
GEN|1|17|Et posuit eas Deus in firmamento caeli, ut lucerent super terram
GEN|1|18|et praeessent diei ac nocti et dividerent lucem ac tenebras. Et vidit Deus quod esset bonum.
GEN|1|19|Et factum est vespere et mane, dies quartus.
GEN|1|20|Dixit etiam Deus: " Pullulent aquae reptile animae viventis, et volatile volet super terram sub firmamento caeli ".
GEN|1|21|Creavitque Deus cete grandia et omnem animam viventem atque motabilem, quam pullulant aquae secundum species suas, et omne volatile secundum genus suum. Et vidit Deus quod esset bonum;
GEN|1|22|benedixitque eis Deus dicens: " Crescite et multiplicamini et replete aquas maris, avesque multiplicentur super terram ".
GEN|1|23|Et factum est vespere et mane, dies quintus.
GEN|1|24|Dixit quoque Deus: " Producat terra animam viventem in genere suo, iumenta et reptilia et bestias terrae secundum species suas ". Factumque est ita.
GEN|1|25|Et fecit Deus bestias terrae iuxta species suas et iumenta secundum species suas et omne reptile terrae in genere suo. Et vidit Deus quod esset bonum.
GEN|1|26|Et ait Deus: " Faciamus hominem ad imaginem et similitudinem nostram; et praesint piscibus maris et volatilibus caeli et bestiis universaeque terrae omnique reptili, quod movetur in terra ".
GEN|1|27|Et creavit Deus hominem ad imaginem suam;ad imaginem Dei creavit illum;masculum et feminam creavit eos.
GEN|1|28|Benedixitque illis Deus et ait illis Deus: " Crescite et multiplicamini et replete terram et subicite eam et dominamini piscibus maris et volatilibus caeli et universis animantibus, quae moventur super terram ".
GEN|1|29|Dixitque Deus: " Ecce dedi vobis omnem herbam afferentem semen super terram et universa ligna, quae habent in semetipsis fructum ligni portantem sementem, ut sint vobis in escam
GEN|1|30|et cunctis animantibus terrae omnique volucri caeli et universis, quae moventur in terra et in quibus est anima vivens, omnem herbam virentem ad vescendum ". Et factum est ita.
GEN|1|31|Viditque Deus cuncta, quae fecit, et ecce erant valde bona. Et factum est vespere et mane, dies sextus.
GEN|2|1|Igitur perfecti sunt caeli et terra et omnis exercitus eorum.
GEN|2|2|Complevitque Deus die septimo opus suum, quod fecerat, et requievit die septimo ab universo opere, quod patrarat.
GEN|2|3|Et benedixit Deus diei septimo et sanctificavit illum, quia in ipso requieverat ab omni opere suo, quod creavit Deus, ut faceret.
GEN|2|4|Istae sunt generationes caeli et terrae, quando creata sunt.In die quo fecit Dominus Deus terram et caelum ­
GEN|2|5|omne virgultum agri, antequam oriretur in terra, omnisque herba regionis, priusquam germinaret; non enim pluerat Dominus Deus super terram, et homo non erat, qui operaretur humum,
GEN|2|6|sed fons ascendebat e terra irrigans universam superficiem terrae ­
GEN|2|7|tunc formavit Dominus Deus hominem pulverem de humo et inspiravit in nares eius spiraculum vitae, et factus est homo in animam viventem.
GEN|2|8|Et plantavit Dominus Deus paradisum in Eden ad orientem, in quo posuit hominem, quem formaverat.
GEN|2|9|Produxitque Dominus Deus de humo omne lignum pulchrum visu et ad vescendum suave, lignum etiam vitae in medio paradisi lignumque scientiae boni et mali.
GEN|2|10|Et fluvius egrediebatur ex Eden ad irrigandum paradisum, qui inde dividitur in quattuor capita.
GEN|2|11|Nomen uni Phison: ipse est, qui circuit omnem terram Hevila, ubi est aurum;
GEN|2|12|et aurum terrae illius optimum est; ibi invenitur bdellium et lapis onychinus.
GEN|2|13|Et nomen fluvio secundo Geon: ipse est, qui circuit omnem terram Aethiopiae.
GEN|2|14|Nomen vero fluminis tertii Tigris: ipse vadit ad orientem Assyriae. Fluvius autem quartus ipse est Euphrates.
GEN|2|15|Tulit ergo Dominus Deus hominem et posuit eum in paradiso Eden, ut operaretur et custodiret illum;
GEN|2|16|praecepitque Dominus Deus homini dicens: " Ex omni ligno paradisi comede;
GEN|2|17|de ligno autem scientiae boni et mali ne comedas; in quocumque enim die comederis ex eo, morte morieris ".
GEN|2|18|Dixit quoque Dominus Deus: " Non est bonum esse hominem solum; faciam ei adiutorium simile sui ".
GEN|2|19|Formatis igitur Dominus Deus de humo cunctis animantibus agri et universis volatilibus caeli, adduxit ea ad Adam, ut videret quid vocaret ea; omne enim, quod vocavit Adam animae viventis, ipsum est nomen eius.
GEN|2|20|Appellavitque Adam nominibus suis cuncta pecora et universa volatilia caeli et omnes bestias agri; Adae vero non inveniebatur adiutor similis eius.
GEN|2|21|Immisit ergo Dominus Deus soporem in Adam. Cumque obdormisset, tulit unam de costis eius et replevit carnem pro ea;
GEN|2|22|et aedificavit Dominus Deus costam, quam tulerat de Adam, in mulierem et adduxit eam ad Adam.
GEN|2|23|Dixitque Adam: Haec nunc os ex ossibus meiset caro de carne mea!Haec vocabitur Virago,quoniam de viro sumpta est haec ".
GEN|2|24|Quam ob rem relinquet vir patrem suum et matrem et adhaerebit uxori suae; et erunt in carnem unam.
GEN|2|25|Erant autem uterque nudi, Adam scilicet et uxor eius, et non erubescebant.
GEN|3|1|Et serpens erat callidior cunctis animantibus agri, quae fecerat Dominus Deus. Qui dixit ad mulierem: " Verene praecepit vobis Deus, ut non comederetis de omni ligno paradisi? ".
GEN|3|2|Cui respondit mulier: " De fructu lignorum, quae sunt in paradiso, vescimur;
GEN|3|3|de fructu vero ligni, quod est in medio paradisi, praecepit nobis Deus, ne comederemus et ne tangeremus illud, ne moriamur ".
GEN|3|4|Dixit autem serpens ad mulierem: " Nequaquam morte moriemini!
GEN|3|5|Scit enim Deus quod in quocumque die comederitis ex eo, aperientur oculi vestri, et eritis sicut Deus scientes bonum et malum ".
GEN|3|6|Vidit igitur mulier quod bonum esset lignum ad vescendum et pulchrum oculis et desiderabile esset lignum ad intellegendum; et tulit de fructu illius et comedit deditque etiam viro suo secum, qui comedit.
GEN|3|7|Et aperti sunt oculi amborum. Cumque cognovissent esse se nudos, consuerunt folia ficus et fecerunt sibi perizomata.
GEN|3|8|Et cum audissent vocem Domini Dei deambulantis in paradiso ad auram post meridiem, abscondit se Adam et uxor eius a facie Domini Dei in medio ligni paradisi.
GEN|3|9|Vocavitque Dominus Deus Adam et dixit ei: " Ubi es? ".
GEN|3|10|Qui ait: " Vocem tuam audivi in paradiso et timui eo quod nudus essem et abscondi me ".
GEN|3|11|Cui dixit: " Quis enim indicavit tibi quod nudus esses, nisi quod ex ligno, de quo tibi praeceperam, ne comederes, comedisti? ".
GEN|3|12|Dixitque Adam: " Mulier, quam dedisti sociam mihi, ipsa dedit mihi de ligno, et comedi ".
GEN|3|13|Et dixit Dominus Deus ad mulierem: " Quid hoc fecisti? ". Quae respondit: " Serpens decepit me, et comedi ".
GEN|3|14|Et ait Dominus Deus ad serpentem: Quia fecisti hoc, maledictus esinter omnia pecoraet omnes bestias agri!Super pectus tuum gradieriset pulverem comedes cunctisdiebus vitae tuae.
GEN|3|15|Inimicitias ponam inter te et mulieremet semen tuum et semen illius;ipsum conteret caput tuum,et tu conteres calcaneum eius ".
GEN|3|16|Mulieri dixit: Multiplicabo aerumnas tuaset conceptus tuos:in dolore paries filios,et ad virum tuum erit appetitus tuus,ipse autem dominabitur tui ".
GEN|3|17|Adae vero dixit: " Quia audisti vocem uxoris tuae et comedisti de ligno, ex quo praeceperam tibi, ne comederes,maledicta humus propter te!In laboribus comedes ex eacunctis diebus vitae tuae.
GEN|3|18|Spinas et tribulos germinabit tibi,et comedes herbas terrae;
GEN|3|19|in sudore vultus tui vesceris pane,donec revertaris ad humum,de qua sumptus es,quia pulvis es et in pulverem reverteris ".
GEN|3|20|Et vocavit Adam nomen uxoris suae Eva, eo quod mater esset cunctorum viventium.
GEN|3|21|Fecit quoque Dominus Deus Adae et uxori eius tunicas pelliceas et induit eos.
GEN|3|22|Et ait Dominus Deus: " Ecce homo factus est quasi unus ex nobis, ut sciat bonum et malum; nunc ergo, ne mittat manum suam et sumat etiam de ligno vitae et comedat et vivat in aeternum! ".
GEN|3|23|Emisit eum Dominus Deus de paradiso Eden, ut operaretur humum, de qua sumptus est.
GEN|3|24|Eiecitque hominem et collocavit ad orientem paradisi Eden cherubim et flammeum gladium atque versatilem ad custodiendam viam ligni vitae.
GEN|4|1|Adam vero cognovit Evam uxo rem suam, quae concepit et peperit Cain dicens: " Acquisivi virum per Dominum ".
GEN|4|2|Rursusque peperit fratrem eius Abel. Et fuit Abel pastor ovium et Cain agricola.
GEN|4|3|Factum est autem post aliquot dies ut offerret Cain de fructibus agri munus Domino.
GEN|4|4|Abel quoque obtulit de primogenitis gregis sui et de adipibus eorum. Et respexit Dominus ad Abel et ad munus eius,
GEN|4|5|ad Cain vero et ad munus illius non respexit. Iratusque est Cain vehementer, et concidit vultus eius.
GEN|4|6|Dixitque Dominus ad eum: " Quare iratus es, et cur concidit facies tua?
GEN|4|7|Nonne si bene egeris, vultum attolles? Sin autem male, in foribus peccatum insidiabitur, et ad te erit appetitus eius, tu autem dominaberis illius ".
GEN|4|8|Dixitque Cain ad Abel fratrem suum: " Egrediamur foras ". Cumque essent in agro, consurrexit Cain adversus Abel fratrem suum et interfecit eum.
GEN|4|9|Et ait Dominus ad Cain: " Ubi est Abel frater tuus? ". Qui respondit: " Nescio. Num custos fratris mei sum ego? ".
GEN|4|10|Dixitque ad eum: " Quid fecisti? Vox sanguinis fratris tui clamat ad me de agro.
GEN|4|11|Nunc igitur maledictus eris procul ab agro, qui aperuit os suum et suscepit sanguinem fratris tui de manu tua!
GEN|4|12|Cum operatus fueris eum, amplius non dabit tibi fructus suos; vagus et profugus eris super terram ".
GEN|4|13|Dixitque Cain ad Dominum: " Maior est poena mea quam ut portem eam.
GEN|4|14|Ecce eicis me hodie a facie agri, et a facie tua abscondar et ero vagus et profugus in terra; omnis igitur, qui invenerit me, occidet me ".
GEN|4|15|Dixitque ei Dominus: " Nequaquam ita fiet, sed omnis qui occiderit Cain, septuplum punietur! ". Posuitque Dominus Cain signum, ut non eum interficeret omnis qui invenisset eum.
GEN|4|16|Egressusque Cain a facie Domini habitavit in terra Nod ad orientalem plagam Eden.
GEN|4|17|Cognovit autem Cain uxorem suam, quae concepit et peperit Henoch. Et aedificavit civitatem vocavitque nomen eius ex nomine filii sui Henoch.
GEN|4|18|Porro Henoch genuit Irad, et Irad genuit Maviael, et Maviael genuit Mathusael, et Mathusael genuit Lamech.
GEN|4|19|Qui accepit uxores duas: nomen uni Ada et nomen alteri Sella.
GEN|4|20|Genuitque Ada Iabel, qui fuit pater habitantium in tentoriis atque pastorum.
GEN|4|21|Et nomen fratris eius Iubal; ipse fuit pater omnium canentium cithara et organo.
GEN|4|22|Sella quoque genuit Tubalcain, qui fuit malleator et faber in cuncta opera aeris et ferri. Soror vero Tubalcain Noema.
GEN|4|23|Dixitque Lamech uxoribus suis: Ada et Sella, audite vocem meam; uxores Lamech, auscultate sermonem meum:occidi virum pro vulnere meoet adulescentulum pro livore meo;
GEN|4|24|septuplum ultio dabitur de Cain, de Lamech vero septuagies septies ".
GEN|4|25|Cognovit quoque Adam uxorem suam, et peperit filium vocavitque nomen eius Seth dicens: " Posuit mihi Deus semen aliud pro Abel, quem occidit Cain ".
GEN|4|26|Sed et Seth natus est filius, quem vocavit Enos. Tunc coeperunt invocare nomen Domini.
GEN|5|1|Hic est liber generationis Adam. In die qua creavit Deus homi nem, ad similitudinem Dei fecit illum.
GEN|5|2|Masculum et feminam creavit eos et benedixit illis; et vocavit nomen eorum Adam in die, quo creati sunt.
GEN|5|3|Vixit autem Adam centum triginta annis et genuit ad similitudinem et imaginem suam vocavitque nomen eius Seth.
GEN|5|4|Et facti sunt dies Adam, postquam genuit Seth, octingenti anni, genuitque filios et filias.
GEN|5|5|Et factum est omne tempus, quod vixit Adam, anni nongenti triginta, et mortuus est.
GEN|5|6|Vixit quoque Seth centum quinque annos et genuit Enos.
GEN|5|7|Vixitque Seth, postquam genuit Enos, octingentis septem annis genuitque filios et filias.
GEN|5|8|Et facti sunt omnes dies Seth nongentorum duodecim annorum, et mortuus est.
GEN|5|9|Vixit vero Enos nonaginta annis et genuit Cainan.
GEN|5|10|Et vixit Enos, postquam genuit Cainan, octingentis quindecim annis et genuit filios et filias.
GEN|5|11|Factique sunt omnes dies Enos nongentorum quinque annorum, et mortuus est.
GEN|5|12|Vixit quoque Cainan septuaginta annis et genuit Malaleel.
GEN|5|13|Et vixit Cainan, postquam genuit Malaleel, octingentos quadraginta annos genuitque filios et filias.
GEN|5|14|Et facti sunt omnes dies Cainan nongenti decem anni, et mortuus est.
GEN|5|15|Vixit autem Malaleel sexaginta quinque annos et genuit Iared.
GEN|5|16|Et vixit Malaleel, postquam genuit Iared, octingentis triginta annis et genuit filios et filias.
GEN|5|17|Et facti sunt omnes dies Malaleel octingenti nonaginta quinque anni, et mortuus est.
GEN|5|18|Vixitque Iared centum sexaginta duobus annis et genuit Henoch.
GEN|5|19|Et vixit Iared, postquam genuit Henoch, octingentos annos et genuit filios et filias.
GEN|5|20|Et facti sunt omnes dies Iared nongenti sexaginta duo anni, et mortuus est.
GEN|5|21|Porro Henoch vixit sexaginta quinque annis et genuit Mathusalam.
GEN|5|22|Et ambulavit Henoch cum Deo, postquam genuit Mathusalam, trecentis annis et genuit filios et filias.
GEN|5|23|Et facti sunt omnes dies Henoch trecenti sexaginta quinque anni,
GEN|5|24|ambulavitque cum Deo et non apparuit, quia tulit eum Deus.
GEN|5|25|Vixit quoque Mathusala centum octoginta septem annos et genuit Lamech.
GEN|5|26|Et vixit Mathusala, postquam genuit Lamech, septingentos octoginta duos annos et genuit filios et filias.
GEN|5|27|Et facti sunt omnes dies Mathusalae nongenti sexaginta novem anni, et mortuus est.
GEN|5|28|Vixit autem Lamech centum octoginta duobus annis et genuit filium
GEN|5|29|vocavitque nomen eius Noe dicens: " Iste consolabitur nos ab operibus nostris et labore manuum nostrarum in agro, cui maledixit Dominus ".
GEN|5|30|Vixitque Lamech, postquam genuit Noe, quingentos nonaginta quinque annos et genuit filios et filias.
GEN|5|31|Et facti sunt omnes dies Lamech septingenti septuaginta septem anni, et mortuus est.
GEN|5|32|Noe vero, cum quingentorum esset annorum, genuit Sem, Cham et Iapheth.
GEN|6|1|Cumque coepissent homines multiplicari super terram et fi lias procreassent,
GEN|6|2|videntes filii Dei filias hominum quod essent pulchrae, acceperunt sibi uxores ex omnibus, quas elegerant.
GEN|6|3|Dixitque Deus: " Non permanebit spiritus meus in homine in aeternum, quia caro est; eruntque dies illius centum viginti annorum ".
GEN|6|4|Gigantes erant super terram in diebus illis et etiam postquam ingressi sunt filii Dei ad filias hominum, illaeque eis genuerunt: isti sunt potentes a saeculo viri famosi.
GEN|6|5|Videns autem Dominus quod multa malitia hominum esset in terra, et cuncta cogitatio cordis eorum non intenta esset nisi ad malum omni tempore,
GEN|6|6|paenituit Dominum quod hominem fecisset in terra. Et tactus dolore cordis intrinsecus:
GEN|6|7|" Delebo, inquit, hominem, quem creavi, a facie terrae, ab homine usque ad pecus, usque ad reptile et usque ad volucres caeli; paenitet enim me fecisse eos ".
GEN|6|8|Noe vero invenit gratiam coram Domino.
GEN|6|9|Hae sunt generationes Noe: Noe vir iustus atque perfectus fuit in generatione sua; cum Deo ambulavit.
GEN|6|10|Et genuit tres filios: Sem, Cham et Iapheth.
GEN|6|11|Corrupta est autem terra coram Deo et repleta est iniquitate.
GEN|6|12|Cumque vidisset Deus terram esse corruptam ­ omnis quippe caro corruperat viam suam super terram ­
GEN|6|13|dixit ad Noe: " Finis universae carnis venit coram me; repleta est enim terra iniquitate a facie eorum, et ecce ego disperdam eos de terra.
GEN|6|14|Fac tibi arcam de lignis cupressinis; mansiunculas in arca facies et bitumine linies eam intrinsecus et extrinsecus.
GEN|6|15|Et sic facies eam: trecentorum cubitorum erit longitudo arcae, quinquaginta cubitorum latitudo et triginta cubitorum altitudo illius.
GEN|6|16|Fenestram in arca facies et cubito consummabis summitatem eius. Ostium autem arcae pones ex latere; tabulatum inferius, medium et superius facies in ea.
GEN|6|17|Ecce ego adducam diluvii aquas super terram, ut interficiam omnem carnem, in qua spiritus vitae est subter caelum: universa, quae in terra sunt, consumentur.
GEN|6|18|Ponamque foedus meum tecum; et ingredieris arcam tu et filii tui, uxor tua et uxores filiorum tuorum tecum.
GEN|6|19|Et ex cunctis animantibus universae carnis bina induces in arcam, ut vivant tecum, masculini sexus et feminini.
GEN|6|20|De volucribus iuxta genus suum et de iumentis in genere suo et ex omni reptili terrae secundum genus suum: bina de omnibus ingredientur ad te, ut possint vivere.
GEN|6|21|Tu autem tolle tecum ex omnibus escis, quae mandi possunt, et comportabis apud te; et erunt tam tibi quam illis in cibum ".
GEN|6|22|Fecit ergo Noe omnia, quae praeceperat illi Deus; sic fecit.
GEN|7|1|Dixitque Dominus ad Noe: " Ingredere tu et omnis domus tua arcam; te enim vidi iustum coram me in generatione hac.
GEN|7|2|Ex omnibus pecoribus mundis tolle septena septena, masculum et feminam; de pecoribus vero non mundis duo duo, masculum et feminam.
GEN|7|3|Sed et de volatilibus caeli septena septena, masculum et feminam, ut salvetur semen super faciem universae terrae.
GEN|7|4|Adhuc enim et post dies septem ego pluam super terram quadraginta diebus et quadraginta noctibus et delebo omnem substantiam, quam feci, de superficie terrae ".
GEN|7|5|Fecit ergo Noe omnia, quae mandaverat ei Dominus.
GEN|7|6|Eratque Noe sescentorum annorum, quando diluvii aquae inundaverunt super terram.
GEN|7|7|Et ingressus est Noe et filii eius, uxor eius et uxores filiorum eius cum eo in arcam propter aquas diluvii.
GEN|7|8|De pecoribus mundis et immundis et de volucribus et ex omni, quod movetur super terram,
GEN|7|9|duo et duo ingressa sunt ad Noe in arcam, masculus et femina, sicut praeceperat Deus Noe.
GEN|7|10|Cumque transissent septem dies, aquae diluvii inundaverunt super terram.
GEN|7|11|Anno sescentesimo vitae Noe, mense secundo, septimo decimo die mensis rupti sunt omnes fontes abyssi magnae, et cataractae caeli apertae sunt;
GEN|7|12|et facta est pluvia super terram quadraginta diebus et quadraginta noctibus.
GEN|7|13|In articulo diei illius ingressus est Noe et Sem et Cham et Iapheth filii eius, uxor illius et tres uxores filiorum eius cum eis in arcam.
GEN|7|14|Ipsi et omne animal secundum genus suum, universaque iumenta in genere suo, et omne reptile, quod movetur super terram in genere suo, cunctumque volatile secundum genus suum, universae aves omnesque volucres
GEN|7|15|ingressae sunt ad Noe in arcam, bina et bina ex omni carne, in qua erat spiritus vitae.
GEN|7|16|Et quae ingressa sunt, masculus et femina ex omni carne introierunt, sicut praeceperat ei Deus; et inclusit eum Dominus de foris.
GEN|7|17|Factumque est diluvium quadraginta diebus super terram, et multiplicatae sunt aquae et elevaverunt arcam in sublime a terra.
GEN|7|18|Vehementer enim inundaverunt et omnia repleverunt in superficie terrae; porro arca ferebatur super aquas.
GEN|7|19|Et aquae praevaluerunt nimis super terram, opertique sunt omnes montes excelsi sub universo caelo.
GEN|7|20|Quindecim cubitis altior fuit aqua super montes, quos operuerat.
GEN|7|21|Consumptaque est omnis caro, quae movebatur super terram, volucrum, pecorum, bestiarum omniumque reptilium, quae reptant super terram, et universi homines:
GEN|7|22|cuncta, in quibus spiraculum vitae in terra, mortua sunt.
GEN|7|23|Et delevit omnem substantiam, quae erat super terram, ab homine usque ad pecus, usque ad reptile et usque ad volucres caeli; et deleta sunt de terra. Remansit autem solus Noe et qui cum eo erant in arca.
GEN|7|24|Obtinueruntque aquae terram centum quinquaginta diebus.
GEN|8|1|Recordatus autem Deus Noe cunctorumque animantium et omnium iumentorum, quae erant cum eo in arca, adduxit spiritum super terram, et imminutae sunt aquae.
GEN|8|2|Et clausi sunt fontes abyssi et cataractae caeli, et prohibitae sunt pluviae de caelo.
GEN|8|3|Reversaeque sunt aquae de terra euntes et redeuntes et coeperunt minui post centum quinquaginta dies.
GEN|8|4|Requievitque arca mense septimo, decima septima die mensis super montes Ararat.
GEN|8|5|At vero aquae ibant et decrescebant usque ad decimum mensem; decimo enim mense, prima die mensis, apparuerunt cacumina montium.
GEN|8|6|Cumque transissent quadraginta dies, aperiens Noe fenestram arcae, quam fecerat, dimisit corvum;
GEN|8|7|qui egrediebatur exiens et rediens, donec siccarentur aquae super terram.
GEN|8|8|Emisit quoque columbam a se, ut videret si iam cessassent aquae super faciem terrae.
GEN|8|9|Quae, cum non invenisset, ubi requiesceret pes eius, reversa est ad eum in arcam; aquae enim erant super universam terram. Extenditque manum et apprehensam intulit in arcam.
GEN|8|10|Exspectatis autem ultra septem diebus aliis, rursum dimisit columbam ex arca.
GEN|8|11|At illa venit ad eum ad vesperam portans ramum olivae virentibus foliis in ore suo. Intellexit ergo Noe quod cessassent aquae super terram.
GEN|8|12|Exspectavitque nihilominus septem alios dies; et emisit columbam, quae non est reversa ultra ad eum.
GEN|8|13|Igitur sescentesimo primo anno, primo mense, prima die mensis, siccatae sunt aquae super terram; et aperiens Noe tectum arcae, et ecce aspexit viditque quod exsiccata erat superficies terrae.
GEN|8|14|Mense secundo, septima et vicesima die mensis, arefacta est terra.
GEN|8|15|Locutus est autem Deus ad Noe dicens:
GEN|8|16|" Egredere de arca tu et uxor tua, filii tui et uxores filiorum tuorum tecum.
GEN|8|17|Cuncta animantia, quae sunt apud te ex omni carne, tam in volatilibus quam in pecoribus et in universis reptilibus, quae reptant super terram, educ tecum, ut pullulent super terram et crescant et multiplicentur super eam ".
GEN|8|18|Egressus est ergo Noe et filii eius, uxor illius et uxores filiorum eius cum eo.
GEN|8|19|Sed et omnia animantia, iumenta, volatilia et reptilia, quae reptant super terram, secundum genus suum egressa sunt de arca.
GEN|8|20|Aedificavit autem Noe altare Domino; et tollens de cunctis pecoribus mundis et volucribus mundis obtulit holocausta super altare.
GEN|8|21|Odoratusque est Dominus odorem suavitatis et locutus est Dominus ad cor suum: " Nequaquam ultra maledicam terrae propter homines, quia cogitatio humani cordis in malum prona est ab adulescentia sua. Non igitur ultra percutiam omnem animam viventem, sicut feci.
GEN|8|22|Cunctis diebus terrae, sementis et messis, frigus et aestus, aestas et hiems, dies et nox non requiescent ".
GEN|9|1|Benedixitque Deus Noe et filiis eius et dixit ad eos: " Crescite et multiplicamini et implete terram.
GEN|9|2|Et terror vester ac tremor sit super cuncta animalia terrae et super omnes volucres caeli cum universis, quae moventur super terram; omnes pisces maris manui vestrae traditi sunt.
GEN|9|3|Omne, quod movetur et vivit, erit vobis in cibum; quasi holera virentia tradidi vobis omnia,
GEN|9|4|excepto quod carnem cum anima, quae est in sanguine, non comedetis.
GEN|9|5|Sanguinem enim animarum vestrarum requiram de manu cunctarum bestiarum; et de manu hominis, de manu viri fratris eius requiram animam hominis.
GEN|9|6|Quicumque effuderit humanum sanguinem,per hominem fundetur sanguis illius;ad imaginem quippe Deifactus est homo.
GEN|9|7|Vos autem crescite et multiplicamini et pullulate super terram et dominamini ei ".
GEN|9|8|Haec quoque dixit Deus ad Noe et ad filios eius cum eo:
GEN|9|9|" Ecce ego statuam pactum meum vobiscum et cum semine vestro post vos
GEN|9|10|et ad omnem animam viventem, quae est vobiscum tam in volucribus quam in iumentis et in omnibus bestiis terrae, quae sunt vobiscum, cunctis, quae egressa sunt de arca, universis bestiis terrae.
GEN|9|11|Statuam pactum meum vobiscum; et nequaquam ultra interficietur omnis caro aquis diluvii, neque erit deinceps diluvium dissipans terram ".
GEN|9|12|Dixitque Deus: " Hoc signum foederis, quod do inter me et vos et ad omnem animam viventem, quae est vobiscum, in generationes sempiternas:
GEN|9|13|arcum meum ponam in nubibus, et erit signum foederis inter me et inter terram.
GEN|9|14|Cumque obduxero nubibus caelum, apparebit arcus meus in nubibus,
GEN|9|15|et recordabor foederis mei vobiscum et cum omni anima vivente, quae carnem vegetat; et non erunt ultra aquae diluvii ad delendum universam carnem.
GEN|9|16|Eritque arcus in nubibus, et videbo illum et recordabor foederis sempiterni, quod pactum est inter Deum et omnem animam viventem universae carnis, quae est super terram ".
GEN|9|17|Dixitque Deus ad Noe: " Hoc erit signum foederis, quod constitui inter me et omnem carnem super terram ".
GEN|9|18|Erant ergo filii Noe, qui egressi sunt de arca, Sem, Cham et Iapheth. Porro Cham ipse est pater Chanaan.
GEN|9|19|Tres isti filii sunt Noe, et ab his disseminatum est omne hominum genus super universam terram.
GEN|9|20|Coepitque Noe agricola plantare vineam;
GEN|9|21|bibensque vinum inebriatus est et nudatus in tabernaculo suo.
GEN|9|22|Quod cum vidisset Cham pater Chanaan, verenda scilicet patris sui esse nudata, nuntiavit duobus fratribus suis foras.
GEN|9|23|At vero Sem et Iapheth pallium imposuerunt umeris suis et incedentes retrorsum operuerunt verecunda patris sui, faciesque eorum aversae erant, et patris virilia non viderunt.
GEN|9|24|Evigilans autem Noe ex vino, cum didicisset, quae fecerat ei filius suus minor,
GEN|9|25|ait:Maledictus Chanaan!Servus servorum erit fratribus suis ".
GEN|9|26|Dixitque:Benedictus Dominus Deus Sem!Sitque Chanaan servus eius.
GEN|9|27|Dilatet Deus Iapheth,et habitet in tabernaculis Sem,sitque Chanaan servus eius ".
GEN|9|28|Vixit autem Noe post diluvium trecentis quinquaginta annis.
GEN|9|29|Et impleti sunt omnes dies eius nongentorum quinquaginta annorum, et mortuus est.
GEN|10|1|Hae sunt generationes filio rum Noe, Sem, Cham et Ia pheth; natique sunt eis filii post diluvium.
GEN|10|2|Filii Iapheth: Gomer et Magog et Madai et Iavan et Thubal et Mosoch et Thiras.
GEN|10|3|Porro filii Gomer: Aschenez et Riphath et Thogorma.
GEN|10|4|Filii autem Iavan: Elisa et Tharsis, Cetthim et Rodanim.
GEN|10|5|Ab his divisae sunt insulae gentium in regionibus suis, unusquisque secundum linguam suam et familias suas in nationibus suis.
GEN|10|6|Filii autem Cham: Chus et Mesraim et Phut et Chanaan.
GEN|10|7|Filii Chus: Saba et Hevila et Sabatha et Regma et Sabathacha. Filii Regma: Saba et Dedan.
GEN|10|8|Porro Chus genuit Nemrod: ipse coepit esse potens in terra
GEN|10|9|et erat robustus venator coram Domino. Ob hoc exivit proverbium: " Quasi Nemrod robustus venator coram Domino ".
GEN|10|10|Fuit autem principium regni eius Babylon et Arach et Achad et Chalanne in terra Sennaar.
GEN|10|11|De terra illa egressus est in Assyriam et aedificavit Nineven et Rohobothir et Chale,
GEN|10|12|Resen quoque inter Nineven et Chale; haec est civitas magna.
GEN|10|13|At vero Mesraim genuit Ludim et Anamim et Laabim, Nephthuim
GEN|10|14|et Phetrusim et Chasluim et Caphtorim, de quibus egressi sunt Philisthim.
GEN|10|15|Chanaan autem genuit Sidonem primogenitum suum, Hetthaeum
GEN|10|16|et Iebusaeum et Amorraeum, Gergesaeum,
GEN|10|17|Hevaeum et Aracaeum, Sinaeum
GEN|10|18|et Aradium, Samaraeum et Emathaeum; et post haec disseminati sunt populi Chananaeorum.
GEN|10|19|Factique sunt termini Chanaan venientibus a Sidone Geraram usque Gazam, donec ingrediaris Sodomam et Gomorram et Adamam et Seboim usque Lesa.
GEN|10|20|Hi sunt filii Cham in cognationibus et linguis terrisque et gentibus suis.
GEN|10|21|De Sem quoque nati sunt, patre omnium filiorum Heber, fratre Iapheth maiore.
GEN|10|22|Filii Sem: Elam et Assur et Arphaxad et Lud et Aram.
GEN|10|23|Filii Aram: Us et Hul et Gether et Mes.
GEN|10|24|At vero Arphaxad genuit Sala, de quo ortus est Heber.
GEN|10|25|Natique sunt Heber filii duo: nomen uni Phaleg, eo quod in diebus eius divisa sit terra, et nomen fratris eius Iectan.
GEN|10|26|Qui Iectan genuit Elmodad et Saleph et Asarmoth, Iare
GEN|10|27|et Adoram et Uzal et Decla
GEN|10|28|et Ebal et Abimael, Saba
GEN|10|29|et Ophir et Hevila et Iobab. Omnes isti filii Iectan;
GEN|10|30|et facta est habitatio eorum de Messa pergentibus usque Sephar montem orientalem.
GEN|10|31|Isti filii Sem secundum cognationes et linguas et regiones in gentibus suis.
GEN|10|32|Hae familiae filiorum Noe iuxta generationes et nationes suas. Ab his divisae sunt gentes in terra post diluvium.
GEN|11|1|Erat autem universa terra labii unius et sermonum eo rundem.
GEN|11|2|Cumque proficiscerentur de oriente, invenerunt campum in terra Sennaar et habitaverunt in eo.
GEN|11|3|Dixitque alter ad proximum suum: " Venite, faciamus lateres et coquamus eos igni ". Habueruntque lateres pro saxis et bitumen pro caemento.
GEN|11|4|Et dixerunt: " Venite, faciamus nobis civitatem et turrim, cuius culmen pertingat ad caelum, et faciamus nobis nomen, ne dividamur super faciem universae terrae ".
GEN|11|5|Descendit autem Dominus, ut videret civitatem et turrim, quam aedificaverunt filii hominum,
GEN|11|6|et dixit Dominus: " Ecce unus est populus et unum labium omnibus; et hoc est initium operationis eorum, nec eis erit deinceps difficile, quidquid cogitaverint facere.
GEN|11|7|Venite igitur, descendamus et confundamus ibi linguam eorum, ut non intellegat unusquisque vocem proximi sui ".
GEN|11|8|Atque ita divisit eos Dominus ex illo loco super faciem universae terrae, et cessaverunt aedificare civitatem.
GEN|11|9|Et idcirco vocatum est nomen eius Babel, quia ibi confusum est labium universae terrae, et inde dispersit eos Dominus super faciem universae terrae.
GEN|11|10|Hae sunt generationes Sem. Sem centum erat annorum, quando genuit Arphaxad biennio post diluvium;
GEN|11|11|vixitque Sem, postquam genuit Arphaxad, quingentos annos et genuit filios et filias.
GEN|11|12|Porro Arphaxad vixit triginta quinque annos et genuit Sala.
GEN|11|13|Vixitque Arphaxad, postquam genuit Sala, quadringentis tribus annis et genuit filios et filias.
GEN|11|14|Sala quoque vixit triginta annis et genuit Heber.
GEN|11|15|Vixitque Sala, postquam genuit Heber, quadringentis tribus annis et genuit filios et filias.
GEN|11|16|Vixit autem Heber triginta quattuor annis et genuit Phaleg.
GEN|11|17|Et vixit Heber, postquam genuit Phaleg, quadringentis triginta annis et genuit filios et filias.
GEN|11|18|Vixit quoque Phaleg triginta annis et genuit Reu.
GEN|11|19|Vixitque Phaleg, postquam genuit Reu, ducentis novem annis et genuit filios et filias.
GEN|11|20|Vixit autem Reu triginta duobus annis et genuit Seruch.
GEN|11|21|Vixitque Reu, postquam genuit Seruch, ducentis septem annis et genuit filios et filias.
GEN|11|22|Vixit vero Seruch triginta annis et genuit Nachor.
GEN|11|23|Vixitque Seruch, postquam genuit Nachor, ducentos annos et genuit filios et filias.
GEN|11|24|Vixit autem Nachor viginti novem annis et genuit Thare.
GEN|11|25|Vixitque Nachor, postquam genuit Thare, centum decem et novem annos et genuit filios et filias.
GEN|11|26|Vixitque Thare septuaginta annis et genuit Abram, Nachor et Aran.
GEN|11|27|Hae sunt autem generationes Thare. Thare genuit Abram, Nachor et Aran. Porro Aran genuit Lot;
GEN|11|28|mortuusque est Aran ante Thare patrem suum in terra nativitatis suae in Ur Chaldaeorum.
GEN|11|29|Duxerunt autem Abram et Nachor uxores: nomen uxoris Abram Sarai, et nomen uxoris Nachor Melcha, filia Aran patris Melchae et patris Ieschae.
GEN|11|30|Erat autem Sarai sterilis nec habebat liberos.
GEN|11|31|Tulitque Thare Abram filium suum et Lot filium Aran filium filii sui et Sarai nurum suam, uxorem Abram filii sui, et eduxit eos de Ur Chaldaeorum, ut irent in terram Chanaan. Veneruntque usque Charran et habitaverunt ibi.
GEN|11|32|Et facti sunt dies Thare ducentorum quinque annorum, et mortuus est in Charran.
GEN|12|1|Dixit autem Dominus ad Abram: Egredere de terra tua et de cognatione tuaet de domo patris tuiin terram, quam monstrabo tibi.
GEN|12|2|Faciamque te in gentem magnamet benedicam tibiet magnificabo nomen tuum,erisque in benedictionem.
GEN|12|3|Benedicam benedicentibus tibiet maledicentibus tibi maledicam,atque in te benedicenturuniversae cognationes terrae! ".
GEN|12|4|Egressus est itaque Abram, sicut praeceperat ei Dominus, et ivit cum eo Lot. Septuaginta quinque annorum erat Abram, cum egrederetur de Charran.
GEN|12|5|Tulitque Sarai uxorem suam et Lot filium fratris sui universamque substantiam, quam acquisiverant, et animas, quas fecerant in Charran, et egressi sunt, ut irent in terram Chanaan; et venerunt in terram Chanaan.
GEN|12|6|Pertransivit Abram terram usque ad locum Sichem, usque ad Quercum Moreh. Chananaeus autem tunc erat in terra.
GEN|12|7|Apparuit autem Dominus Abram et dixit ei: " Semini tuo dabo terram hanc. Qui aedificavit ibi altare Domino, qui apparuerat ei.
GEN|12|8|Et inde transgrediens ad montem, qui erat contra orientem Bethel, tetendit ibi tabernaculum suum ab occidente habens Bethel et ab oriente Hai; aedificavit quoque ibi altare Domino et invocavit nomen Domini.
GEN|12|9|Perrexitque Abram de mansione in mansionem usque ad Nageb.
GEN|12|10|Facta est autem fames in terra; descenditque Abram in Aegyptum, ut peregrinaretur ibi; praevaluerat enim fames in terra.
GEN|12|11|Cumque prope esset, ut ingrederetur Aegyptum, dixit Sarai uxori suae: " Novi quod pulchra sis mulier
GEN|12|12|et quod, cum viderint te Aegyptii, dicturi sunt: "Uxor ipsius est"; et interficient me et te reservabunt.
GEN|12|13|Dic ergo, obsecro te, quod soror mea sis, ut bene sit mihi propter te, et vivat anima mea ob gratiam tui ".
GEN|12|14|Cum itaque ingressus esset Abram Aegyptum, viderunt Aegyptii mulierem quod esset pulchra nimis,
GEN|12|15|et viderunt eam principes pharaonis et laudaverunt eam apud illum; et sublata est mulier in domum pharaonis.
GEN|12|16|Abram vero bene usus est propter illam; fueruntque ei oves et boves et asini et servi et famulae et asinae et cameli.
GEN|12|17|Flagellavit autem Dominus pharaonem plagis maximis et domum eius propter Sarai uxorem Abram.
GEN|12|18|Vocavitque pharao Abram et dixit ei: " Quidnam est hoc quod fecisti mihi? Quare non indicasti mihi quod uxor tua esset?
GEN|12|19|Quam ob causam dixisti esse sororem tuam, ut tollerem eam mihi in uxorem? Nunc igitur, ecce coniux tua: accipe eam et vade! ".
GEN|12|20|Praecepitque pharao super Abram viris; et deduxerunt eum et uxorem illius et omnia, quae habebat.
GEN|13|1|Ascendit ergo Abram de Ae gypto ipse et uxor eius et om nia, quae habebat, et Lot cum eo ad Nageb.
GEN|13|2|Abram autem erat dives valde in pecoribus, argento et auro.
GEN|13|3|Et profectus est de mansione in mansionem a Nageb in Bethel usque ad locum, ubi prius fixerat tabernaculum inter Bethel et Hai,
GEN|13|4|in loco altaris, quod fecerat prius, et invocavit ibi nomen Domini.
GEN|13|5|Sed et Lot, qui ibat cum Abram, fuerunt greges ovium et armenta et tabernacula;
GEN|13|6|nec poterat eos capere terra, ut habitarent simul: erat quippe substantia eorum multa, et nequibant habitare communiter.
GEN|13|7|Unde et facta est rixa inter pastores gregum Abram et pastores gregum Lot. Eo autem tempore Chananaeus et Pherezaeus habitabant in illa terra.
GEN|13|8|Dixit ergo Abram ad Lot: " Ne, quaeso, sit iurgium inter me et te et inter pastores meos et pastores tuos: fratres enim sumus.
GEN|13|9|Nonne universa terra coram te est? Recede a me, obsecro: si ad sinistram ieris, ego dexteram tenebo; si tu dexteram elegeris, ego ad sinistram pergam ".
GEN|13|10|Elevatis itaque Lot oculis, vidit omnem circa regionem Iordanis, quae universa irrigabatur, antequam subverteret Dominus Sodomam et Gomorram, sicut paradisus Domini et sicut Aegyptus usque in Segor.
GEN|13|11|Elegitque sibi Lot omnem regionem circa Iordanem et recessit ad orientem; divisique sunt alterutrum a fratre suo.
GEN|13|12|Abram habitavit in terra Chanaan; Lot vero moratus est in oppidis, quae erant circa Iordanem, et tabernacula movit usque ad Sodomam.
GEN|13|13|Homines autem Sodomitae pessimi erant et peccatores coram Domino nimis.
GEN|13|14|Dixitque Dominus ad Abram, postquam divisus est Lot ab eo: " Leva oculos tuos et vide a loco, in quo nunc es, ad aquilonem et ad meridiem, ad orientem et ad occidentem:
GEN|13|15|omnem terram, quam conspicis, tibi dabo et semini tuo usque in sempiternum;
GEN|13|16|faciamque semen tuum sicut pulverem terrae: si quis potest hominum numerare pulverem terrae, semen quoque tuum numerare poterit.
GEN|13|17|Surge et perambula terram in longitudine et in latitudine sua, quia tibi daturus sum eam ".
GEN|13|18|Movens igitur tabernaculum suum, Abram venit et habitavit iuxta Quercus Mambre, quae sunt in Hebron, aedificavitque ibi altare Domino.
GEN|14|1|Factum est autem in illo tempore, ut Amraphel rex Sennaar et Arioch rex Ellasar et Chodorlahomor rex Elam et Thadal rex gentium
GEN|14|2|inirent bellum contra Bara regem Sodomae et contra Bersa regem Gomorrae et contra Sennaab regem Adamae et contra Semeber regem Seboim contraque regem Belae; ipsa est Segor.
GEN|14|3|Omnes hi convenerunt in vallem Siddim, quae nunc est mare Salis.
GEN|14|4|Duodecim annis servierant Chodorlahomor et tertio decimo anno recesserunt ab eo.
GEN|14|5|Igitur anno quarto decimo venit Chodorlahomor et reges, qui erant cum eo, percusseruntque Raphaim in Astharothcarnaim et Zuzim in Ham et Emim in Savecariathaim
GEN|14|6|et Chorraeos in montibus Seir usque ad Elpharan, quae est in deserto.
GEN|14|7|Reversique sunt et venerunt ad fontem Mesphat; ipsa est Cades. Et percusserunt omnem regionem Amalecitarum et etiam Amorraeum, qui habitabat in Asasonthamar.
GEN|14|8|Et egressi sunt rex Sodomae et rex Gomorrae rexque Adamae et rex Seboim necnon et rex Belae, quae est Segor; et direxerunt contra eos aciem in valle Siddim,
GEN|14|9|scilicet adversus Chodorlahomor regem Elam et Thadal regem gentium et Amraphel regem Sennaar et Arioch regem Ellasar: quattuor reges adversus quinque.
GEN|14|10|Vallis autem Siddim habebat puteos multos bituminis. Itaque rex Sodomae et Gomorrae terga verterunt cecideruntque illuc; et, qui remanserant, fugerunt ad montem.
GEN|14|11|Tulerunt autem omnem substantiam Sodomae et Gomorrae et universa, quae ad cibum pertinent, et abierunt;
GEN|14|12|ceperunt et Lot et substantiam eius, filium fratris Abram, qui habitabat in Sodoma.
GEN|14|13|Et ecce unus, qui evaserat, nuntiavit Abram Hebraeo, qui habitabat iuxta Quercus Mambre Amorraei fratris Eschol et fratris Aner; hi enim pepigerant foedus cum Abram.
GEN|14|14|Quod cum audisset Abram, captum videlicet Lot fratrem suum, numeravit expeditos vernaculos suos trecentos decem et octo et persecutus est usque Dan;
GEN|14|15|et, divisis sociis, irruit super eos nocte percussitque eos et persecutus est eos usque Hoba, quae est ad laevam Damasci;
GEN|14|16|reduxitque omnem substantiam, necnon et Lot fratrem suum cum substantia illius, mulieres quoque et populum.
GEN|14|17|Egressus est autem rex Sodomae in occursum eius, postquam reversus est a caede Chodorlahomor et regum, qui cum eo erant, in vallem Save, quae est vallis Regis.
GEN|14|18|At vero Melchisedech rex Salem proferens panem et vinum ­ erat enim sacerdos Dei altissimi ­
GEN|14|19|benedixit ei et ait: Benedictus Abram a Deo excelso, qui creavit caelum et terram
GEN|14|20|et benedictus Deus excelsus,qui tradidit hostes tuos in manus tuas ".Et dedit ei decimas ex omnibus.
GEN|14|21|Dixit autem rex Sodomae ad Abram: " Da mihi animas; substantiam tolle tibi ".
GEN|14|22|Qui respondit ei: " Levo manum meam ad Dominum, Deum excelsum, creatorem caeli et terrae,
GEN|14|23|a filo subteminis usque ad corrigiam caligae non accipiam ex omnibus, quae tua sunt, ne dicas: "Ego ditavi Abram";
GEN|14|24|exceptis his, quae comederunt iuvenes, et partibus virorum, qui venerunt mecum, Aner, Eschol et Mambre: isti accipient partes suas ".
GEN|15|1|His itaque transactis, factus est sermo Domini ad Abram per visionem dicens: "Noli timere, Abram! Ego protector tuus sum, et merces tua magna erit nimis ".
GEN|15|2|Dixitque Abram: " Domine Deus, quid dabis mihi? Ego vadam absque liberis, et heres domus meae erit Damascenus Eliezer ".
GEN|15|3|Addiditque Abram: " En mihi non dedisti semen, et ecce vernaculus meus heres meus erit ".
GEN|15|4|Sed ecce sermo Domini factus est ad eum: "Non erit hic heres tuus, sed qui egredietur de visceribus tuis, ipsum habebis heredem ".
GEN|15|5|Eduxitque eum foras et ait illi: " Suspice caelum et numera stellas, si potes ". Et dixit ei: " Sic erit semen tuum ".
GEN|15|6|Credidit Domino, et reputatum est ei ad iustitiam.
GEN|15|7|Dixitque ad eum: " Ego Dominus, qui eduxi te de Ur Chaldaeorum, ut darem tibi terram istam, et possideres eam ".
GEN|15|8|Et ille ait: " Domine Deus, unde scire possum quod possessurus sim eam?.
GEN|15|9|Respondens Dominus: " Sume, inquit, mihi vitulam triennem et capram trimam et arietem annorum trium, turturem quoque et columbam ".
GEN|15|10|Qui tollens universa haec divisit ea per medium et utrasque partes contra se altrinsecus posuit; aves autem non divisit.
GEN|15|11|Descenderuntque volucres super cadavera, et abigebat eas Abram.
GEN|15|12|Cumque sol occumberet, sopor irruit super Abram, et ecce horror magnus et tenebrosus invasit eum.
GEN|15|13|Dictumque est ad eum: " Scito praenoscens quod peregrinum futurum sit semen tuum in terra non sua, et subicient eos servituti et affligent quadringentis annis.
GEN|15|14|Verumtamen et gentem, cui servituri sunt, ego iudicabo, et post haec egredientur cum magna substantia.
GEN|15|15|Tu autem ibis ad patres tuos in pace, sepultus in senectute bona.
GEN|15|16|Generatione autem quarta revertentur huc; necdum enim completae sunt iniquitates Amorraeorum usque ad praesens tempus ".
GEN|15|17|Cum ergo occubuisset sol, facta est caligo tenebrosa, et apparuit clibanus fumans et lampas ignis transiens inter divisiones illas.
GEN|15|18|In illo die pepigit Dominus cum Abram foedus dicens: " Semini tuo dabo terram hanc a fluvio Aegypti usque ad magnum fluvium Euphraten,
GEN|15|19|Cinaeos et Cenezaeos, Cedmonaeos
GEN|15|20|et Hetthaeos et Pherezaeos, Raphaim quoque
GEN|15|21|et Amorraeos et Chananaeos et Gergesaeos et Iebusaeos ".
GEN|16|1|Sarai autem uxor Abram non genuerat ei liberos; sed habens ancillam Aegyptiam nomine Agar,
GEN|16|2|dixit marito suo: " Ecce conclusit me Dominus, ne parerem; ingredere ad ancillam meam, si forte saltem ex illa suscipiam filios ". Cumque ille acquiesceret deprecanti,
GEN|16|3|tulit Agar Aegyptiam ancillam suam post annos decem quam habitare coeperant in terra Chanaan, et dedit eam viro suo uxorem.
GEN|16|4|Qui ingressus est ad eam. At illa concepisse se videns despexit dominam suam.
GEN|16|5|Dixitque Sarai ad Abram: " Inique agis contra me; ego dedi ancillam meam in sinum tuum, quae videns quod conceperit, despectui me habet. Iudicet Dominus inter me et te ".
GEN|16|6|Cui respondens Abram: " Ecce, ait, ancilla tua in manu tua est; utere ea, ut libet ". Affligente igitur eam Sarai, aufugit ab ea.
GEN|16|7|Cumque invenisset illam angelus Domini iuxta fontem aquae in deserto, ad fontem in via Sur,
GEN|16|8|dixit: " Agar, ancilla Sarai, unde venis et quo vadis? ". Quae respondit: " A facie Sarai dominae meae ego fugio ".
GEN|16|9|Dixitque ei angelus Domini: " Revertere ad dominam tuam et humiliare sub manibus ipsius ".
GEN|16|10|Et dixit ei angelus Domini: " Multiplicans multiplicabo semen tuum, et non numerabitur prae multitudine ".
GEN|16|11|Et dixit ei angelus Domini: Ecce, concepisti et paries filiumvocabisque nomen eius Ismael,eo quod audierit Dominus afflictionem tuam.
GEN|16|12|Hic erit homo onagro similis;manus eius contra omnes,et manus omnium contra eum;et e regione universorum fratrum suorum figet tabernacula ".
GEN|16|13|Vocavit autem nomen Domini, qui loquebatur ad eam: " Tu Deus, qui vidisti me ". Dixit enim: " Profecto hic vidi posteriora videntis me ".
GEN|16|14|Propterea appellatur puteus ille Lahairoi (id est Viventis et Videntis me); ipse est inter Cades et Barad.
GEN|16|15|Peperitque Agar Abrae filium; qui vocavit nomen filii sui, quem pepererat Agar, Ismael.
GEN|16|16|Octoginta et sex annorum erat Abram, quando peperit ei Agar Ismaelem.
GEN|17|1|Postquam Abram nonaginta et novem annorum factus est, apparuit ei Dominus dixitque ad eum: " Ego Deus omnipotens, ambula coram me et esto perfectus.
GEN|17|2|Ponamque foedus meum inter me et te et multiplicabo te vehementer nimis.
GEN|17|3|Cecidit Abram pronus in faciem.
GEN|17|4|Dixitque ei Deus: " Ecce pactum meum tecum. Erisque pater multarum gentium,
GEN|17|5|nec ultra vocabitur nomen tuum Abram, sed Abraham erit nomen tuum, quia patrem multarum gentium constitui te.
GEN|17|6|Faciamque te crescere vehementissime et ponam te in gentes; regesque ex te egredientur.
GEN|17|7|Et statuam pactum meum inter me et te et inter semen tuum post te in generationibus suis foedere sempiterno, ut sim Deus tuus et seminis tui post te.
GEN|17|8|Daboque tibi et semini tuo post te terram peregrinationis tuae, omnem terram Chanaan in possessionem aeternam; eroque Deus eorum ".
GEN|17|9|Dixit iterum Deus ad Abraham: " Tu autem pactum meum custodies, et semen tuum post te in generationibus suis.
GEN|17|10|Hoc est pactum meum, quod observabitis, inter me et vos et semen tuum post te. Circumcidetur ex vobis omne masculinum,
GEN|17|11|et circumcidetis carnem praeputii vestri, ut sit in signum foederis inter me et vos.
GEN|17|12|Infans octo dierum circumcidetur in vobis: omne masculinum in generationibus vestris, tam vernaculus quam empticius ex omnibus alienigenis, quicumque non fuerit de stirpe vestra.
GEN|17|13|Circumcidetur vernaculus et empticius, eritque pactum meum in carne vestra in foedus aeternum.
GEN|17|14|Masculus, cuius praeputii caro circumcisa non fuerit, delebitur anima illa de populo suo; pactum meum irritum fecit.
GEN|17|15|Dixit quoque Deus ad Abraham: " Sarai uxorem tuam non vocabis nomen eius Sarai, sed Sara erit nomen eius.
GEN|17|16|Et benedicam ei; et ex illa quoque dabo tibi filium. Benedicturus sum eam, eritque in nationes; reges populorum orientur ex ea ".
GEN|17|17|Cecidit Abraham in faciem suam et risit dicens in corde suo: " Putasne centenario nascetur filius? Et Sara nonagenaria pariet? ".
GEN|17|18|Dixitque ad Deum: " Utinam Ismael vivat coram te ".
GEN|17|19|Et ait Deus: " Sara uxor tua pariet tibi filium, vocabisque nomen eius Isaac; et constituam pactum meum illi in foedus sempiternum et semini eius post eum.
GEN|17|20|Super Ismael quoque exaudivi te: ecce benedicam ei et crescere faciam et multiplicabo eum vehementissime; duodecim duces generabit, et faciam illum in gentem magnam.
GEN|17|21|Pactum vero meum statuam ad Isaac, quem pariet tibi Sara tempore isto in anno altero ".
GEN|17|22|Cumque cessasset loqui cum eo, ascendit Deus ab Abraham.
GEN|17|23|Tulit ergo Abraham Ismael filium suum et omnes vernaculos domus suae universosque, quos emerat: cunctos mares ex omnibus viris domus suae; et circumcidit carnem praeputii eorum statim in ipsa die, sicut praeceperat ei Deus.
GEN|17|24|Abraham nonaginta novem erat annorum, quando circumcisus est in carne praeputii sui;
GEN|17|25|et Ismael filius eius tredecim annos impleverat tempore circumcisionis suae.
GEN|17|26|Eadem die circumcisus est Abraham et Ismael filius eius;
GEN|17|27|et omnes viri domus illius, tam vernaculi quam empticii ex alienigenis, circumcisi sunt cum eo.
GEN|18|1|Apparuit autem ei Dominus iuxta Quercus Mambre se denti in ostio tabernaculi sui in ipso fervore diei.
GEN|18|2|Cumque elevasset oculos, apparuerunt ei tres viri stantes prope eum. Quos cum vidisset, cucurrit in occursum eorum de ostio tabernaculi et adoravit in terram
GEN|18|3|et dixit: " Domine mi, si inveni gratiam in oculis tuis, ne transeas servum tuum;
GEN|18|4|afferatur pauxillum aquae, et lavate pedes vestros et requiescite sub arbore.
GEN|18|5|Ponamque buccellam panis, et confortate cor vestrum, postea transibitis; idcirco enim declinastis ad servum vestrum ". Qui dixerunt: " Fac ut locutus es ".
GEN|18|6|Festinavit Abraham in tabernaculum ad Saram dixitque: " Accelera, tria sata similae commisce et fac subcinericios panes ".
GEN|18|7|Ipse vero ad armentum cucurrit et tulit inde vitulum tenerrimum et optimum deditque puero; qui festinavit et coxit illum.
GEN|18|8|Tulit quoque butyrum et lac et vitulum, quem coxerat, et posuit coram eis. Ipse vero stabat iuxta eos sub arbore; et comederunt.
GEN|18|9|Dixeruntque ad eum: " Ubi est Sara uxor tua? ". Ille respondit: " Ecce in tabernaculo est ".
GEN|18|10|Cui dixit: " Revertens veniam ad te tempore isto, et habebit filium Sara uxor tua ". Quo audito, Sara risit ad ostium tabernaculi, quod erat post eum.
GEN|18|11|Erant autem ambo senes provectaeque aetatis, et desierant Sarae fieri muliebria.
GEN|18|12|Quae risit occulte dicens: " Postquam consenui, et dominus meus vetulus est, voluptas mihi erit? ".
GEN|18|13|Dixit autem Dominus ad Abraham: " Quare risit Sara dicens: "Num vere paritura sum anus?"".
GEN|18|14|Numquid Domino est quidquam difficile? Revertar ad te hoc eodem tempore, et habebit Sara filium ".
GEN|18|15|Negavit Sara dicens: " Non risi ", timore perterrita. Ille autem dixit: Non; sed risisti ".
GEN|18|16|Cum ergo surrexissent inde viri, direxerunt oculos contra Sodomam; et Abraham simul gradiebatur deducens eos.
GEN|18|17|Dixitque Dominus: " Num celare potero Abraham, quae gesturus sum,
GEN|18|18|cum futurus sit in gentem magnam ac robustissimam, et benedicendae sint in illo omnes nationes terrae?
GEN|18|19|Nam elegi eum, ut praecipiat filiis suis et domui suae post se, ut custodiant viam Domini et faciant iustitiam et iudicium, ut adducat Dominus super Abraham omnia, quae locutus est ad eum ".
GEN|18|20|Dixit itaque Dominus: " Clamor contra Sodomam et Gomorram multiplicatus est, et peccatum eorum aggravatum est nimis.
GEN|18|21|Descendam et videbo utrum clamorem, qui venit ad me, opere compleverint an non; sciam ".
GEN|18|22|Converteruntque se inde viri et abierunt Sodomam; Abraham vero adhuc stabat coram Domino.
GEN|18|23|Et appropinquans ait: " Numquid vere perdes iustum cum impio?
GEN|18|24|Si forte fuerint quinquaginta iusti in civitate, vere perdes et non parces loco illi propter quinquaginta iustos, si fuerint in eo?
GEN|18|25|Absit a te, ut rem hanc facias et occidas iustum cum impio, fiatque iustus sicut impius; absit a te. Nonne iudex universae terrae faciet iudicium? ".
GEN|18|26|Dixitque Dominus: " Si invenero Sodomae quinquaginta iustos in medio civitatis, dimittam omni loco propter eos ".
GEN|18|27|Respondensque Abraham ait: " Ecce coepi loqui ad Dominum meum, cum sim pulvis et cinis.
GEN|18|28|Quid, si forte minus quinquaginta iustis quinque fuerint? Delebis propter quinque universam urbem? ". Et ait: " Non delebo, si invenero ibi quadraginta quinque ".
GEN|18|29|Rursumque locutus est ad eum: " Si forte inventi fuerint ibi quadraginta? ". Ait: " Non percutiam propter quadraginta ".
GEN|18|30|" Ne, quaeso, inquit, indignetur Dominus meus, si loquar. Si forte ibi inventi fuerint triginta? ". Respondit: " Non faciam, si invenero ibi triginta ".
GEN|18|31|" Ecce, ait, coepi loqui ad Dominum meum. Si forte inventi fuerint ibi viginti? ". Dixit: " Non interficiam propter viginti ".
GEN|18|32|" Obsecro, inquit, ne irascatur Dominus meus, si loquar adhuc semel. Si forte inventi fuerint ibi decem? ". Dixit: " Non delebo propter decem ".
GEN|18|33|Abiit Dominus, postquam cessavit loqui ad Abraham; et ille reversus est in locum suum.
GEN|19|1|Veneruntque duo angeli Sodomam vespere, sedente Lot in foribus civitatis. Qui cum vidisset eos, surrexit et ivit obviam eis adoravitque pronus in terram
GEN|19|2|et dixit: " Obsecro, domini mei, declinate in domum pueri vestri et pernoctate; lavate pedes vestros et mane proficiscemini in viam vestram ". Qui dixerunt: " Minime, sed in platea pernoctabimus ".
GEN|19|3|Compulit illos oppido, et diverterunt ad eum. Ingressisque domum illius fecit convivium et coxit azyma, et comederunt.
GEN|19|4|Prius autem quam irent cubitum, viri civitatis, viri Sodomae, vallaverunt domum a iuvene usque ad senem, omnis populus simul.
GEN|19|5|Vocaveruntque Lot et dixerunt ei: " Ubi sunt viri, qui introierunt ad te nocte? Educ illos ad nos, ut cognoscamus eos ".
GEN|19|6|Egressus ad eos Lot post tergum occludens ostium ait:
GEN|19|7|" Nolite, quaeso, fratres mei, nolite malum hoc facere.
GEN|19|8|Ecce, habeo duas filias, quae necdum cognoverunt virum; educam eas ad vos, et facite eis sicut placuerit vobis, dummodo viris istis nihil faciatis; ideo enim ingressi sunt sub umbra tecti mei ".
GEN|19|9|At illi dixerunt: " Recede illuc ". Et rursus: " Unus ingressus est, inquiunt, ut advena et vult iudicare? Te ergo ipsum magis quam hos affligemus ". Vimque faciebant Lot vehementissime, iamque prope erat, ut effringerent fores.
GEN|19|10|Et ecce miserunt manum viri et introduxerunt ad se Lot clauseruntque ostium;
GEN|19|11|et eos, qui foris erant, percusserunt caecitate a minimo usque ad maximum, ita ut ostium invenire non possent.
GEN|19|12|Dixerunt autem viri ad Lot: " Habes hic quempiam tuorum? Generum et filios et filias et omnes, qui tui sunt in urbe, educ de loco hoc:
GEN|19|13|delebimus enim locum istum, eo quod increverit clamor contra eos coram Domino, qui misit nos, ut perdamus eam ".
GEN|19|14|Egressus itaque Lot locutus est ad generos suos, qui accepturi erant filias eius, et dixit: " Surgite, egredimini de loco isto, quia delebit Dominus civitatem ". Et visus est eis quasi ludens loqui.
GEN|19|15|Cumque esset mane, cogebant eum angeli dicentes: " Surge, tolle uxorem tuam et duas filias, quas habes hic, ne pereas in scelere civitatis ".
GEN|19|16|Tardante illo, apprehenderunt viri manum eius et manum uxoris ac duarum filiarum eius, eo quod parceret Dominus illi.
GEN|19|17|Et eduxerunt eum posueruntque extra civitatem. Ibi locutus est: " Salvare, agitur de vita tua; noli respicere post tergum, nec stes in omni circa regione; sed in monte salvum te fac, ne pereas ".
GEN|19|18|Dixitque Lot ad eos: " Non, quaeso, Domine.
GEN|19|19|Ecce invenit servus tuus gratiam coram te, et magnificasti misericordiam tuam, quam fecisti mecum, ut salvares animam meam; nec possum in monte salvari, ne forte apprehendat me malum et moriar.
GEN|19|20|Ecce, civitas haec iuxta, ad quam possum fugere, parva, et salvabor in ea ­ numquid non modica est? ­ et vivet anima mea ".
GEN|19|21|Dixitque ad eum: " Ecce, etiam in hoc suscepi preces tuas, ut non subvertam urbem, pro qua locutus es.
GEN|19|22|Festina et salvare ibi, quia non potero facere quidquam, donec ingrediaris illuc ". Idcirco vocatum est nomen urbis illius Segor.
GEN|19|23|Sol egressus est super terram, et Lot ingressus est Segor.
GEN|19|24|Igitur Dominus pluit super Sodomam et Gomorram sulphur et ignem a Domino de caelo
GEN|19|25|et subvertit civitates has et omnem circa regionem, universos habitatores urbium et cuncta terrae virentia.
GEN|19|26|Respiciensque uxor eius post se versa est in statuam salis.
GEN|19|27|Abraham autem consurgens mane venit ad locum, ubi steterat prius cum Domino,
GEN|19|28|intuitus est Sodomam et Gomorram et universam terram regionis illius; viditque ascendentem favillam de terra quasi fornacis fumum.
GEN|19|29|Cum enim subverteret Deus civitates regionis illius, recordatus Abrahae liberavit Lot de subversione urbium, in quibus habitaverat.
GEN|19|30|Ascenditque Lot de Segor et mansit in monte, duae quoque filiae eius cum eo; timuerat enim manere in Segor. Et mansit in spelunca ipse et duae filiae eius.
GEN|19|31|Dixitque maior ad minorem: " Pater noster senex est, et nullus virorum remansit in terra, qui possit ingredi ad nos iuxta morem universae terrae.
GEN|19|32|Veni, inebriemus patrem nostrum vino dormiamusque cum eo, ut servare possimus ex patre nostro semen ".
GEN|19|33|Dederunt itaque patri suo bibere vinum nocte illa, et ingressa est maior dormivitque cum patre; at ille non sensit, nec quando accubuit filia nec quando surrexit.
GEN|19|34|Altera quoque die dixit maior ad minorem: " Ecce, dormivi heri cum patre meo; demus ei bibere vinum etiam hac nocte, et ingressa dormies cum eo, ut salvemus semen de patre nostro ".
GEN|19|35|Dederunt et illa nocte patri suo bibere vinum, ingressaque minor filia dormivit cum eo; et ne tunc quidem sensit, quando illa concubuerit vel quando surrexerit.
GEN|19|36|Conceperunt ergo duae filiae Lot de patre suo.
GEN|19|37|Peperitque maior filium et vocavit nomen eius Moab; ipse est pater Moabitarum usque in praesentem diem.
GEN|19|38|Minor quoque peperit filium et vocavit nomen eius Benammi (id est Filius populi mei); ipse est pater Ammonitarum usque hodie.
GEN|20|1|Profectus inde Abraham in terram Nageb, habitavit in ter Cades et Sur et peregrinatus est in Geraris.
GEN|20|2|Dixitque de Sara uxore sua: " Soror mea est ". Misit ergo Abimelech rex Gerarae et tulit eam.
GEN|20|3|Venit autem Deus ad Abimelech per somnium nocte et ait illi: " En morieris propter mulierem, quam tulisti; habet enim virum ".
GEN|20|4|Abimelech vero non tetigerat eam. Et ait: " Domine, num gentem etiam iustam interficies?
GEN|20|5|Nonne ipse dixit mihi: "Soror mea est", et ipsa quoque ait: "Frater meus est"? In simplicitate cordis mei et munditia manuum mearum feci hoc ".
GEN|20|6|Dixitque ad eum Deus per somnium: " Et ego scio quod simplici corde feceris; et ideo custodivi te, ne peccares in me, et non dimisi, ut tangeres eam.
GEN|20|7|Nunc igitur redde viro suo uxorem, quia propheta est; et orabit pro te, et vives. Si autem nolueris reddere, scito quod morte morieris tu et omnia, quae tua sunt ".
GEN|20|8|Statimque de nocte consurgens Abimelech vocavit omnes servos suos et locutus est universa verba haec in auribus eorum; timueruntque viri valde.
GEN|20|9|Vocavit autem Abimelech etiam Abraham et dixit ei: " Quid fecisti nobis? Quid peccavi in te, quia induxisti super me et super regnum meum peccatum grande? Quae non debuisti facere, fecisti mihi ".
GEN|20|10|Rursusque ait: " Quid vidisti, ut hoc faceres? ".
GEN|20|11|Respondit Abraham: " Cogitavi mecum: Certe non est timor Dei in loco isto, et interficient me propter uxorem meam.
GEN|20|12|Alias autem et vere soror mea est, filia patris mei et non filia matris meae, et duxi eam in uxorem.
GEN|20|13|Cum autem vagari me faceret Deus de domo patris mei, dixi ad eam: Hanc misericordiam facies mecum: in omni loco, ad quem ingrediemur, dices quod frater tuus sim ".
GEN|20|14|Tulit igitur Abimelech oves et boves et servos et ancillas et dedit Abraham; reddiditque illi Saram uxorem suam
GEN|20|15|et ait: " Ecce terra mea coram te; ubicumque tibi placuerit, habita ".
GEN|20|16|Sarae autem dixit: " Ecce mille argenteos dedi fratri tuo; ecce hoc erit tibi in velamen oculorum ad omnes, qui tecum sunt, et apud omnes iustificaberis ".
GEN|20|17|Orante autem Abraham, sanavit Deus Abimelech et uxorem ancillasque eius et pepererunt;
GEN|20|18|concluserat enim Dominus omnem vulvam domus Abimelech propter Saram uxorem Abraham.
GEN|21|1|Visitavit autem Dominus Saram, sicut promiserat, et implevit Sarae, quae locutus est;
GEN|21|2|concepitque et peperit Abrahae filium in senectute eius tempore, quo praedixerat ei Deus.
GEN|21|3|Vocavitque Abraham nomen filii sui, quem genuit ei Sara, Isaac
GEN|21|4|et circumcidit eum octavo die, sicut praeceperat ei Deus.
GEN|21|5|Cum Abraham centum esset annorum, natus est ei Isaac filius eius.
GEN|21|6|Dixitque Sara: Risum fecit mihi Deus;quicumque audierit, corridebit mihi?.
GEN|21|7|Rursumque ait: Quis auditurum crederet Abrahamquod Sara lactaret filios,quia peperit ei filiumiam seni? ".
GEN|21|8|Crevit igitur puer et ablactatus est. Fecitque Abraham grande convivium in die ablactationis eius.
GEN|21|9|Cumque vidisset Sara filium Agar Aegyptiae iocantem cum Isaac filio suo, dixit ad Abraham:
GEN|21|10|" Eice ancillam hanc et filium eius; non enim erit heres filius ancillae cum filio meo Isaac ".
GEN|21|11|Dure accepit hoc Abraham propter filium suum.
GEN|21|12|Cui dixit Deus: " Non tibi videatur asperum super puero et super ancilla tua; omnia, quae dixerit tibi Sara, audi vocem eius, quia in Isaac vocabitur tibi semen.
GEN|21|13|Sed et filium ancillae faciam in gentem magnam, quia semen tuum est ".
GEN|21|14|Surrexit itaque Abraham mane et tollens panem et utrem aquae imposuit scapulae eius tradiditque puerum et dimisit eam. Quae cum abisset, errabat in deserto Bersabee.
GEN|21|15|Cumque consumpta esset aqua in utre, abiecit puerum subter unum arbustum
GEN|21|16|et abiit; seditque e regione procul, quantum potest arcus iacere. Dixit enim: " Non videbo morientem puerum ". Et sedens contra levavit vocem suam et flevit.
GEN|21|17|Exaudivit autem Deus vocem pueri; vocavitque angelus Dei Agar de caelo dicens: " Quid tibi, Agar? Noli timere; exaudivit enim Deus vocem pueri de loco, in quo est.
GEN|21|18|Surge, tolle puerum et tene illum manu tua, quia in gentem magnam faciam eum ".
GEN|21|19|Aperuitque Deus oculos eius; quae videns puteum aquae abiit et implevit utrem deditque puero bibere.
GEN|21|20|Et fuit Deus cum eo; qui crevit et moratus est in solitudine factusque est iuvenis sagittarius.
GEN|21|21|Habitavitque in deserto Pharan; et accepit illi mater sua uxorem de terra Aegypti.
GEN|21|22|Eodem tempore dixit Abimelech et Phicol princeps exercitus eius ad Abraham: " Deus tecum est in universis, quae agis.
GEN|21|23|Iura ergo per Deum, ne noceas mihi et posteris meis stirpique meae; sed iuxta fidem, quam feci tibi, facies mihi et terrae, in qua versatus es advena ".
GEN|21|24|Dixitque Abraham: " Ego iurabo ".
GEN|21|25|Et increpavit Abraham Abimelech propter puteum aquae, quem vi abstulerant servi eius.
GEN|21|26|Responditque Abimelech: " Nescivi quis fecerit hanc rem; sed et tu non indicasti mihi, et ego non audivi praeter hodie ".
GEN|21|27|Tulit itaque Abraham oves et boves et dedit Abimelech; percusseruntque ambo foedus.
GEN|21|28|Et statuit Abraham septem agnas gregis seorsum.
GEN|21|29|Cui dixit Abimelech: " Quid sibi volunt septem agnae istae, quas stare fecisti seorsum? ".
GEN|21|30|At ille: " Septem, inquit, agnas accipies de manu mea, ut sint in testimonium mihi, quoniam ego fodi puteum istum ".
GEN|21|31|Idcirco vocatus est locus ille Bersabee, quia ibi uterque iuraverunt.
GEN|21|32|Et inierunt foedus in Bersabee.
GEN|21|33|Surrexit autem Abimelech et Phicol princeps militiae eius reversique sunt in terram Philisthim. Abraham vero plantavit nemus in Bersabee et invocavit ibi nomen Domini, Dei aeterni. 34 Et fuit colonus in terra Philisthim diebus multis.
GEN|22|1|Quae postquam gesta sunt, tentavit Deus Abraham et di xit ad eum: " Abraham ". Ille respondit: " Adsum ".
GEN|22|2|Ait: " Tolle filium tuum unigenitum, quem diligis, Isaac et vade in terram Moria; atque offer eum ibi in holocaustum super unum montium, quem monstravero tibi ".
GEN|22|3|Igitur Abraham de nocte consurgens stravit asinum suum ducens secum duos iuvenes suos et Isaac filium suum. Cumque concidisset ligna in holocaustum, surrexit et abiit ad locum, quem praeceperat ei Deus.
GEN|22|4|Die autem tertio, elevatis oculis, vidit locum procul
GEN|22|5|dixitque ad pueros suos: " Exspectate hic cum asino. Ego et puer illuc usque properantes, postquam adoraverimus, revertemur ad vos ".
GEN|22|6|Tulit quoque ligna holocausti et imposuit super Isaac filium suum; ipse vero portabat in manibus ignem et cultrum. Cumque duo pergerent simul,
GEN|22|7|dixit Isaac Abrahae patri suo: " Pater mi ". Ille respondit: " Quid vis, fili? ". " Ecce, inquit, ignis et ligna; ubi est victima holocausti? ".
GEN|22|8|Dixit Abraham: " Deus providebit sibi victimam holocausti, fili mi ".Pergebant ambo pariter;
GEN|22|9|et venerunt ad locum, quem ostenderat ei Deus, in quo aedificavit Abraham altare et desuper ligna composuit. Cumque colligasset Isaac filium suum, posuit eum in altari super struem lignorum
GEN|22|10|extenditque Abraham manum et arripuit cultrum, ut immolaret filium suum.
GEN|22|11|Et ecce angelus Domini de caelo clamavit: " Abraham, Abraham ". Qui respondit: " Adsum ".
GEN|22|12|Dixitque: " Non extendas manum tuam super puerum neque facias illi quidquam. Nunc cognovi quod times Deum et non pepercisti filio tuo unigenito propter me ".
GEN|22|13|Levavit Abraham oculos suos viditque arietem unum inter vepres haerentem cornibus; quem assumens obtulit holocaustum pro filio.
GEN|22|14|Appellavitque nomen loci illius: " Dominus videt ". Unde usque hodie dicitur: " In monte Dominus videtur ".
GEN|22|15|Vocavit autem angelus Domini Abraham secundo de caelo et dixit:
GEN|22|16|" Per memetipsum iuravi, dicit Dominus: quia fecisti hanc rem et non pepercisti filio tuo unigenito,
GEN|22|17|benedicam tibi et multiplicabo semen tuum sicut stellas caeli et velut arenam, quae est in litore maris. Possidebit semen tuum portas inimicorum suorum,
GEN|22|18|et benedicentur in semine tuo omnes gentes terrae, quia oboedisti voci meae ".
GEN|22|19|Reversus est Abraham ad pueros suos, et surrexerunt abieruntque Bersabee simul, et habitavit Abraham in Bersabee.
GEN|22|20|His ita gestis, nuntiatum est Abrahae quod Melcha quoque genuisset filios Nachor fratri suo:
GEN|22|21|Us primogenitum et Buz fratrem eius et Camuel patrem Aram
GEN|22|22|et Cased et Azau, Pheldas quoque et Iedlaph
GEN|22|23|ac Bathuel, de quo nata est Rebecca. Octo istos genuit Melcha Nachor fratri Abrahae. 24 Concubina vero illius, nomine Reuma, peperit Tabee et Gaham et Tahas et Maacha.
GEN|23|1|Vixit autem Sara centum viginti septem annis
GEN|23|2|et mortua est in Cariatharbe, quae est Hebron, in terra Chanaan; venitque Abraham, ut plangeret et fleret eam.
GEN|23|3|Cumque surrexisset ab officio funeris, locutus est ad filios Heth dicens:
GEN|23|4|" Advena sum et inquilinus apud vos; date mihi possessionem sepulcri vobiscum, ut sepeliam mortuum meum ".
GEN|23|5|Responderunt filii Heth dicentes:
GEN|23|6|" Audi nos, domine, princeps Dei es apud nos: in nobilissimo sepulcrorum nostrorum sepeli mortuum tuum; nullusque te prohibebit, quin in sepulcro eius sepelias mortuum tuum ".
GEN|23|7|Surrexit Abraham et adoravit populum terrae, filios videlicet Heth,
GEN|23|8|dixitque ad eos: " Si placet animae vestrae, ut sepeliam mortuum meum, audite me et intercedite pro me apud Ephron filium Seor,
GEN|23|9|ut det mihi speluncam Machpela, quam habet in extrema parte agri sui. Pecunia digna tradat eam mihi coram vobis in possessionem sepulcri ".
GEN|23|10|Sedebat autem Ephron in medio filiorum Heth. Responditque Ephron Hetthaeus ad Abraham, filiis Heth audientibus cunctis, qui ingrediebantur portam civitatis illius, dicens:
GEN|23|11|" Nequaquam ita fiat, domine mi, ausculta me. Agrum do tibi et speluncam, quae in eo est, praesentibus filiis populi mei; sepeli mortuum tuum ".
GEN|23|12|Adoravit Abraham coram populo terrae
GEN|23|13|et locutus est ad Ephron, audiente populo terrae: " Quaeso, ut audias me. Dabo pecuniam pro agro; suscipe eam, et sic sepeliam mortuum meum in eo ".
GEN|23|14|Respondit Ephron ad Abraham dicens ei:
GEN|23|15|" Domine mi, audi me. Terra quadringentorum siclorum argenti inter me et te quid est hoc? Sepeli mortuum tuum ".
GEN|23|16|Auscultavit Abraham Ephron et appendit pecuniam, quam Ephron postulaverat, audientibus filiis Heth, quadringentos siclos argenti, sicut mos erat apud negotiatores.
GEN|23|17|Confirmatusque est ager Ephronis, qui erat in Machpela respiciens Mambre, tam ipse quam spelunca in eo et omnes arbores eius in cunctis terminis eius per circuitum,
GEN|23|18|Abrahae in possessionem, videntibus filiis Heth cunctis, qui intrabant portam civitatis illius.
GEN|23|19|Deinde sepelivit Abraham Saram uxorem suam in spelunca agri Machpela, qui respiciebat Mambre ­ haec est Hebron ­ in terra Chanaan.
GEN|23|20|Et confirmatus est ager et antrum, quod erat in eo, Abrahae in possessionem sepulcri a filiis Heth.
GEN|24|1|Erat autem Abraham senex dierumque multorum; et Do minus in cunctis benedixerat ei.
GEN|24|2|Dixitque Abraham ad servum seniorem domus suae, qui praeerat omnibus, quae habebat: " Pone manum tuam subter femur meum,
GEN|24|3|ut adiurem te per Dominum, Deum caeli et Deum terrae, ut non accipias uxorem filio meo de filiabus Chananaeorum, inter quos habito;
GEN|24|4|sed ad terram et cognationem meam proficiscaris et inde accipias uxorem filio meo Isaac ".
GEN|24|5|Respondit servus: " Si noluerit mulier venire mecum in terram hanc, num reducere debeo filium tuum ad terram, a quo tu egressus es? ".
GEN|24|6|Dixit Abraham: " Cave, ne quando reducas illuc filium meum.
GEN|24|7|Dominus, Deus caeli, qui tulit me de domo patris mei et de terra nativitatis meae, qui locutus est mihi et iuravit mihi dicens: "Semini tuo dabo terram hanc", ipse mittet angelum suum coram te, et accipies inde uxorem filio meo.
GEN|24|8|Sin autem noluerit mulier sequi te, non teneberis iuramento; filium tantum meum ne reducas illuc ".
GEN|24|9|Posuit ergo servus manum sub femore Abraham domini sui et iuravit illi super hac re.
GEN|24|10|Tulitque servus decem camelos de grege domini sui et abiit ex omnibus bonis eius portans secum; profectusque perrexit in Aram Naharaim ad urbem Nachor.
GEN|24|11|Cumque camelos fecisset accumbere extra oppidum iuxta puteum aquae vespere, tempore quo solent mulieres egredi ad hauriendam aquam, dixit:
GEN|24|12|" Domine,Deus domini mei Abraham, occurre obsecro mihi hodie et fac misericordiam cum domino meo Abraham.
GEN|24|13|Ecce ego sto prope fontem aquae, et filiae habitatorum huius civitatis egredientur ad hauriendam aquam.
GEN|24|14|Igitur puella, cui ego dixero: "Inclina hydriam tuam, ut bibam", et illa responderit: "Bibe, quin et camelis tuis dabo potum", ipsa est, quam praeparasti servo tuo Isaac, et per hoc intellegam quod feceris misericordiam cum domino meo ".
GEN|24|15|Necdum intra se verba compleverat, et ecce Rebecca egrediebatur filia Bathuel filii Melchae uxoris Nachor fratris Abraham habens hydriam in scapula:
GEN|24|16|puella decora nimis, virgo et incognita viro. Descendit ad fontem et implevit hydriam ac revertebatur.
GEN|24|17|Occurritque ei servus et ait: " Pauxillum mihi ad sorbendum praebe aquae de hydria tua ".
GEN|24|18|Quae respondit: " Bibe, domine mi ". Celeriterque deposuit hydriam super ulnam suam et dedit ei potum.
GEN|24|19|Cumque ille bibisset, adiecit: " Quin et camelis tuis hauriam aquam, donec cuncti bibant ".
GEN|24|20|Effundensque hydriam in canalibus recurrit ad puteum, ut hauriret aquam; et haustam omnibus camelis dedit.
GEN|24|21|Ille autem contemplabatur eam tacitus, scire volens utrum prosperum fecisset iter suum Dominus an non.
GEN|24|22|Postquam ergo biberunt cameli, protulit vir anulum aureum pondo dimidii sicli pro naribus et duas armillas pro manibus eius pondo siclorum decem;
GEN|24|23|dixitque: " Cuius es filia? lndica mihi. Est in domo patris tui locus nobis ad pernoctandum? ".
GEN|24|24|Quae respondit: " Filia Bathuelis sum filii Melchae, quem peperit Nachor ".
GEN|24|25|Et addidit dicens: " Palearum quoque et pabuli plurimum est apud nos et locus ad pernoctandum ".
GEN|24|26|Inclinavit se homo et adoravit Dominum
GEN|24|27|dicens: " Benedictus Dominus, Deus domini mei Abraham, qui non abstulit misericordiam et veritatem suam a domino meo et recto itinere me perduxit in domum fratris domini mei ".
GEN|24|28|Cucurrit itaque puella et nuntiavit in domum matris suae omnia, quae evenerant.
GEN|24|29|Habebat autem Rebecca fratrem nomine Laban, qui festinus egressus est ad hominem, ubi erat fons.
GEN|24|30|Cumque vidisset anulum in naribus et armillas in manibus sororis suae et audisset cuncta verba referentis: " Haec locutus est mihi homo ", venit ad virum, qui stabat iuxta camelos et prope fontem aquae;
GEN|24|31|dixitque ad eum: " Ingredere, benedicte Domini, cur foris stas? Praeparavi domum et locum camelis ".
GEN|24|32|Et introduxit eum in hospitium ac destravit camelos; deditque paleas et pabulum camelis et aquam ad lavandos pedes eius et virorum, qui venerant cum eo.
GEN|24|33|Et apposuit in conspectu eius panem. Qui ait: " Non comedam, donec loquar sermones meos ". Respondit: " Loquere ".
GEN|24|34|At ille: " Servus, inquit, Abraham sum;
GEN|24|35|et Dominus benedixit domino meo valde, magnificatusque est; et dedit ei oves et boves, argentum et aurum, servos et ancillas, camelos et asinos.
GEN|24|36|Et peperit Sara uxor domini mei filium domino meo in senectute sua; deditque illi omnia, quae habuerat.
GEN|24|37|Et adiuravit me dominus meus dicens: "Non accipies uxorem filio meo de filiabus Chananaeorum, in quorum terra habito;
GEN|24|38|sed ad domum patris mei perges et de cognatione mea accipies uxorem filio meo".
GEN|24|39|Ego vero respondi domino meo: Quid, si noluerit venire mecum mulier?
GEN|24|40|"Dominus, ait, in cuius conspectu ambulo, mittet angelum suum tecum et diriget viam tuam; accipiesque uxorem filio meo de cognatione mea et de domo patris mei.
GEN|24|41|Innocens eris a maledictione mea, cum veneris ad propinquos meos, et non dederint tibi; tunc innocens eris a maledictione mea".
GEN|24|42|Veni ergo hodie ad fontem et dixi: Domine, Deus domini mei Abraham, si direxisti viam meam, in qua nunc ambulo,
GEN|24|43|ecce sto iuxta fontem aquae; et virgo, quae egredietur ad hauriendam aquam, audierit a me: "Da mihi pauxillum aquae ad bibendum ex hydria tua";
GEN|24|44|et dixerit mihi: "Et tu bibe, et camelis tuis hauriam", ipsa est mulier, quam praeparavit Dominus filio domini mei.
GEN|24|45|Dum haec tacitus mecum volverem, apparuit Rebecca veniens cum hydria, quam portabat in scapula; descenditque ad fontem et hausit aquam. Et aio ad eam: Da mihi paululum bibere.
GEN|24|46|Quae festina deposuit hydriam de umero et dixit mihi: "Et tu bibe, et camelis tuis potum tribuam". Bibi, et adaquavit camelos.
GEN|24|47|Interrogavique eam et dixi: Cuius es filia? Quae respondit: "Filia Bathuelis sum filii Nachor, quem peperit illi Melcha".Suspendi itaque anulum in naribus eius et armillas posui in manibus eius.
GEN|24|48|Pronusque adoravi Dominum benedicens Domino, Deo domini mei Abraham, qui perduxit me recto itinere, ut sumerem filiam fratris domini mei filio eius.
GEN|24|49|Quam ob rem, si facitis misericordiam et veritatem cum domino meo, indicate mihi; sin autem aliud placet, et hoc dicite mihi, ut vadam ad dexteram sive ad sinistram ".
GEN|24|50|Responderunt Laban et Bathuel: " A Domino egressus est sermo; non possumus extra placitum eius quidquam aliud loqui tecum.
GEN|24|51|En Rebecca coram te est; tolle eam et proficiscere, et sit uxor filii domini tui, sicut locutus est Dominus ".
GEN|24|52|Quod cum audisset puer Abraham, procidens adoravit in terram Dominum.
GEN|24|53|Prolatisque vasis argenteis et aureis ac vestibus, dedit ea Rebeccae; res pretiosas dedit fratri eius et matri.
GEN|24|54|Tunc comederunt et biberunt ipse et viri, qui erant cum eo, et pernoctaverunt ibi.Surgens autem mane locutus est puer: " Dimittite me, ut vadam ad dominum meum ".
GEN|24|55|Responderuntque frater eius et mater: " Maneat puella saltem decem dies apud nos et postea proficiscetur ".
GEN|24|56|" Nolite, ait, me retinere, quia Dominus direxit viam meam; dimittite me, ut pergam ad dominum meum ".
GEN|24|57|Dixerunt: " Vocemus puellam et quaeramus ipsius voluntatem ".
GEN|24|58|Cumque vocata venisset, sciscitati sunt: " Vis ire cum homine isto? ". Quae ait: " Vadam ".
GEN|24|59|Dimiserunt ergo Rebeccam sororem eorum et nutricem illius servumque Abraham et comites eius,
GEN|24|60|imprecantes prospera sorori suae atque dicentes: Soror nostra es,crescas in mille milia,et possideat semen tuumportas inimicorum suorum! ".
GEN|24|61|Igitur surrexit Rebecca et puellae illius et, ascensis camelis, secutae sunt virum; sumpsitque servus Rebeccam et abiit.
GEN|24|62|Isaac autem venerat a regione putei Lahairoi et habitabat in terra Nageb.
GEN|24|63|Et egressus est Isaac ad lamentandum in agro, inclinata iam die. Cumque levasset oculos, vidit camelos venientes.
GEN|24|64|Rebecca quoque levavit oculos et vidit Isaac; descenditque de camelo
GEN|24|65|et ait ad puerum: " Quis est ille homo, qui venit per agrum in occursum nobis? ". Dixitque ei: " Ipse est dominus meus ". At illa tollens cito velum operuit se.
GEN|24|66|Servus autem cuncta, quae gesserat, narravit Isaac;
GEN|24|67|qui introduxit eam in tabernaculum Sarae matris suae et accepit Rebeccam uxorem; et dilexit eam et consolatus est a morte matris suae.
GEN|25|1|Abraham vero aliam duxit uxorem nomine Ceturam,
GEN|25|2|quae peperit ei Zamran et Iecsan et Madan et Madian et Iesboc et Sue.
GEN|25|3|Iecsan quoque genuit Saba et Dedan. Filii Dedan fuerunt Assurim et Latusim et Loommim.
GEN|25|4|At vero ex Madian ortus est Epha et Opher et Henoch et Abida et Eldaa. Omnes hi filii Ceturae.
GEN|25|5|Deditque Abraham cuncta, quae possederat, Isaac;
GEN|25|6|filiis autem concubinarum suarum largitus est munera et separavit eos ab Isaac filio suo, dum adhuc ipse viveret, ad plagam orientalem.
GEN|25|7|Fuerunt autem dies vitae Abrahae centum septuaginta quinque anni.
GEN|25|8|Et deficiens mortuus est Abraham in senectute bona provectaeque aetatis et plenus dierum congregatusque est ad populum suum.
GEN|25|9|Et sepelierunt eum Isaac et Ismael filii sui in spelunca Machpela, quae sita est in agro Ephron filii Seor Hetthaei e regione Mambre,
GEN|25|10|quem emerat a filiis Heth. Ibi sepultus est ipse et Sara uxor eius.
GEN|25|11|Et post obitum illius benedixit Deus Isaac filio eius, qui habitabat iuxta puteum Lahairoi.
GEN|25|12|Hae sunt generationes Ismael filii Abrahae, quem peperit ei Agar Aegyptia famula Sarae.
GEN|25|13|Et haec nomina filiorum Ismael in vocabulis et generationibus suis: primogenitus Ismaelis Nabaioth, dein Cedar et Adbeel et Mabsam,
GEN|25|14|Masma quoque et Duma et Massa,
GEN|25|15|Hadad et Thema, Iethur et Naphis et Cedma.
GEN|25|16|Isti sunt filii Ismaelis, et haec nomina eorum per vicos et mansiones eorum: duodecim principes tribuum suarum.
GEN|25|17|Et facti sunt anni vitae Ismaelis centum triginta septem; deficiens mortuus est et appositus ad populum suum.
GEN|25|18|Habitaverunt autem ab Hevila usque Sur, quae respicit Aegyptum introeuntibus Assyriam. In faciem cunctorum fratrum suorum obiit.
GEN|25|19|Hae sunt generationes Isaac filii Abraham: Abraham genuit Isaac;
GEN|25|20|qui, cum quadraginta esset annorum, duxit uxorem Rebeccam filiam Bathuelis Aramaei de Paddanaram, sororem Laban Aramaei.
GEN|25|21|Deprecatusque est Isaac Dominum pro uxore sua, eo quod esset sterilis. Qui exaudivit eum et dedit conceptum Rebeccae.
GEN|25|22|Sed collidebantur in utero eius parvuli. Quae ait: " Si sic est, cur mihi? ". Perrexitque, ut consuleret Dominum.
GEN|25|23|Qui respondens ait: Duae gentes sunt in utero tuo,et duo populi ex ventre tuo dividentur;populusque populum superabit,et maior serviet minori ".
GEN|25|24|Iam tempus pariendi venerat, et ecce gemini in utero eius.
GEN|25|25|Qui primus egressus est rufus erat et totus quasi pallium pilosum; vocatumque est nomen eius Esau. Postea frater eius egrediens plantam Esau tenebat manu, et idcirco appellatum est nomen eius Iacob.
GEN|25|26|Sexagenarius erat Isaac, quando nati sunt parvuli.
GEN|25|27|Quibus adultis, factus est Esau vir gnarus venandi et homo agrestis; Iacob autem vir compositus et habitans in tabernaculis.
GEN|25|28|Isaac amabat Esau, eo quod de venationibus illius libenter vesceretur; et Rebecca diligebat Iacob.
GEN|25|29|Coxit autem Iacob pulmentum; ad quem, cum venisset Esau de agro lassus,
GEN|25|30|ait: " Da mihi de coctione hac rufa, quia oppido lassus sum ". Quam ob causam vocatum est nomen eius Edom (id est Rufus).
GEN|25|31|Cui dixit Iacob: " Vende mihi prius primogenita tua ".
GEN|25|32|Ille respondit: " En morior; quid mihi proderunt primogenita? ".
GEN|25|33|Ait Iacob: " Iura ergo mihi ". Iuravit et vendidit primogenita.
GEN|25|34|Et sic, accepto pane et lentis edulio, comedit et bibit; surrexit et abiit parvipendens quod primogenita vendidisset.
GEN|26|1|Orta autem fame super terram post eam sterilitatem, quae acciderat in diebus Abraham, abiit Isaac ad Abimelech regem Philisthim in Gerara.
GEN|26|2|Apparuitque ei Dominus et ait: " Ne descendas in Aegyptum, sed habita in terra, quam dixero tibi,
GEN|26|3|et peregrinare in ea; eroque tecum et benedicam tibi. Tibi enim et semini tuo dabo universas regiones has complens iuramentum, quod spopondi Abraham patri tuo,
GEN|26|4|et multiplicabo semen tuum sicut stellas caeli daboque posteris tuis universas regiones has; et benedicentur in semine tuo omnes gentes terrae,
GEN|26|5|eo quod oboedierit Abraham voci meae et custodierit praecepta et mandata mea et iustificationes legesque servaverit ".
GEN|26|6|Mansit itaque Isaac in Geraris.
GEN|26|7|Qui, cum interrogaretur a viris loci illius super uxore sua, respondit: Soror mea est ". Timuerat enim confiteri quod sibi esset sociata coniugio, reputans ne forte interficerent eum propter illius pulchritudinem.
GEN|26|8|Cumque pertransissent dies plurimi et ibidem moraretur, prospiciens Abimelech rex Philisthim per fenestram vidit eum iocantem cum Rebecca uxore sua.
GEN|26|9|Et, accersito eo, ait: " Perspicuum est quod uxor tua sit; cur mentitus es eam sororem tuam esse? ". Respondit: " Timui, ne morerer propter eam ".
GEN|26|10|Dixitque Abimelech: " Quare hoc fecisti nobis? Potuit coire quispiam de populo cum uxore tua, et induxeras super nos grande peccatum ". Praecepitque omni populo dicens:
GEN|26|11|" Qui tetigerit hominem hunc et uxorem eius, morte morietur ".
GEN|26|12|Sevit autem Isaac in terra illa et invenit in ipso anno centuplum; benedixitque ei Dominus.
GEN|26|13|Et locupletatus est homo et ibat proficiens atque succrescens, donec magnus vehementer effectus est;
GEN|26|14|habuitque possessionem ovium et armentorum et familiae plurimum.Ob haec invidentes ei Philisthim
GEN|26|15|omnes puteos, quos foderant servi patris illius in diebus Abraham, obstruxerunt implentes humo,
GEN|26|16|in tantum ut ipse Abimelech diceret ad Isaac: " Recede a nobis, quoniam potentior nostri factus es valde ".
GEN|26|17|Et ille discedens tentoria fixit ad torrentem Gerarae habitavitque ibi.
GEN|26|18|Rursum fodit puteos, quos foderant in diebus patris sui Abraham et quos, illo mortuo, obstruxerant Philisthim. Appellavitque eos eisdem nominibus, quibus ante pater vocaverat.
GEN|26|19|Foderunt servi Isaac in torrente et reppererunt ibi puteum aquae vivae.
GEN|26|20|Sed et ibi iurgium fuit pastorum Gerarae adversus pastores Isaac dicentium: " Nostra est aqua! ". Quam ob rem nomen putei vocavit Esec (id est Iurgium), quia iurgati sunt cum eo.
GEN|26|21|Foderunt autem et alium puteum, et pro illo quoque rixati sunt; appellavitque eum Sitna (id est Inimicitias).
GEN|26|22|Profectus inde fodit alium puteum, pro quo non contenderunt; itaque vocavit nomen eius Rehoboth (id est Latitudinem) dicens: " Nunc dilatavit nos Dominus, et crescemus in terra ".
GEN|26|23|Ascendit autem ex illo loco in Bersabee,
GEN|26|24|ubi apparuit ei Dominus in ipsa nocte dicens: Ego sum Deus Abraham patris tui.Noli timere, quia tecum sum;benedicam tibiet multiplicabo semen tuumpropter servum meum Abraham ".
GEN|26|25|Itaque aedificavit ibi altare et, invocato nomine Domini, extendit tabernaculum, et servi Isaac foderunt ibi puteum.
GEN|26|26|Abimelech autem venit ad eum de Geraris et Ochozath amicus illius et Phicol dux militum,
GEN|26|27|et locutus est eis Isaac: " Quid venistis ad me hominem, quem odistis et expulistis a vobis? ".
GEN|26|28|Qui responderunt: " Vidimus tecum esse Dominum et idcirco diximus: Sit iuramentum inter nos et te, et ineamus tecum foedus,
GEN|26|29|ut non facias nobis quidquam mali, sicut et nos non attigimus te et nihil fecimus tibi nisi bonum et cum pace dimisimus te. Tu es enim benedictus Domini ".
GEN|26|30|Fecit ergo eis convivium, et comederunt et biberunt.
GEN|26|31|Surgentesque mane iuraverunt sibi mutuo. Dimisitque eos Isaac, et profecti sunt ab eo cum pace.
GEN|26|32|Ecce autem venerunt in ipso die servi Isaac annuntiantes ei de puteo, quem foderant, atque dicentes: " Invenimus aquam ".
GEN|26|33|Unde appellavit eum Sabee (quod significat Abundantiam); et nomen urbi impositum est Bersabee usque in praesentem diem.
GEN|26|34|Esau vero quadragenarius duxit uxores Iudith filiam Beeri Hetthaei et Basemath filiam Elon Hetthaei.
GEN|26|35|Quae ambae offenderant animum Isaac et Rebeccae.
GEN|27|1|Senuit autem Isaac, et caligaverunt oculi eius, et videre non poterat. Vocavitque Esau filium suum maiorem et dixit ei: " Fili mi ". Qui respondit: " Adsum ".
GEN|27|2|Cui pater: " Vides, inquit, quod senuerim et ignorem diem mortis meae;
GEN|27|3|sume arma tua, pharetram et arcum, et egredere in agrum. Cumque venatu aliquid apprehenderis,
GEN|27|4|fac mihi inde pulmentum, sicut velle me nosti, et affer, ut comedam; et benedicat tibi anima mea, antequam moriar ".
GEN|27|5|Rebecca autem audierat Isaac loquentem cum Esau filio suo. Esau ergo abiit in agrum, ut venationem caperet et offerret eam.
GEN|27|6|Rebecca autem dixit filio suo Iacob: " Ecce, audivi patrem tuum loquentem cum Esau fratre tuo et dicentem ei:
GEN|27|7|"Affer mihi venationem tuam et fac cibos, ut comedam et benedicam tibi coram Domino, antequam moriar".
GEN|27|8|Nunc ergo, fili mi, audi vocem meam in eo, quod praecipio tibi.
GEN|27|9|Pergens ad gregem affer mihi duos haedos optimos, ut faciam ex eis escas patri tuo, quibus libenter vescitur.
GEN|27|10|Quas cum intuleris patri tuo, et comederit, benedicat tibi, priusquam moriatur ".
GEN|27|11|Cui ille respondit: " Nosti quod Esau frater meus homo pilosus sit, et ego lenis.
GEN|27|12|Si attrectaverit me pater meus et senserit, timeo, ne putet me sibi voluisse illudere; et inducam super me maledictionem pro benedictione".
GEN|27|13|Ad quem mater: " In me sit, ait, ista maledictio, fili mi; tantum audi vocem meam et perge afferque, quae dixi ".
GEN|27|14|Abiit et attulit deditque matri. Paravit illa cibos, sicut noverat velle patrem illius.
GEN|27|15|Et vestibus Esau valde bonis, quas apud se habebat domi, induit eum
GEN|27|16|pelliculasque haedorum circumdedit manibus et colli nuda protexit;
GEN|27|17|dedit pulmentum optimum et panes, quos coxerat, in manus filii sui Iacob.
GEN|27|18|Qui ingressus ad patrem suum dixit: " Pater mi ". At ille respondit: " Audio. Quis es tu, fili mi? ".
GEN|27|19|Dixitque Iacob ad patrem suum: " Ego sum Esau primogenitus tuus. Feci sicut praecepisti mihi; surge, sede et comede de venatione mea, ut benedicat mihi anima tua ".
GEN|27|20|Rursum Isaac ad filium suum: " Quomodo, inquit, tam cito invenire potuisti, fili mi? ". Qui respondit: " Voluntas Domini Dei tui fuit, ut occurreret mihi ".
GEN|27|21|Dixitque Isaac ad Iacob: " Accede huc, ut tangam te, fili mi, et probem, utrum tu sis filius meus Esau an non ".
GEN|27|22|Accessit ille ad patrem, et, palpato eo, dixit Isaac: " Vox quidem, vox Iacob est, sed manus, manus sunt Esau ".
GEN|27|23|Et non cognovit eum, quia pilosae manus similitudinem maioris expresserant. Benedixit ergo illi.
GEN|27|24|Ait: " Tu es filius meus Esau? ". Respondit: " Ego sum ".
GEN|27|25|At ille: " Affer, inquit, mihi, et comedam de venatione tua, fili mi, ut benedicat tibi anima mea ". Quos cum oblatos comedisset, obtulit ei etiam vinum. Quo hausto,
GEN|27|26|dixit ad eum Isaac pater eius: " Accede ad me et da mihi osculum, fili mi ".
GEN|27|27|Accessit et osculatus est eum. Statimque, ut sensit vestimentorum illius fragrantiam, benedicens illi ait: Ecce odor filii meisicut odor agri pleni,cui benedixit Dominus.
GEN|27|28|Det tibi Deus de rore caeliet de pinguedine terraeet abundantiam frumenti et vini.
GEN|27|29|Et serviant tibi populi,et adorent te nationes;esto dominus fratrum tuorum,et incurventur ante te filii matris tuae.Qui maledixerit tibi, sit maledictus;et, qui benedixerit tibi, sit benedictus! ".
GEN|27|30|Vix Isaac benedictionem Iacob finierat, et Iacob egressus erat a patre suo Isaac, venit Esau frater eius
GEN|27|31|coctosque de venatione cibos intulit patri dicens: " Surge, pater mi, et comede de venatione filii tui, ut benedicat mihi anima tua ".
GEN|27|32|Dixitque illi Isaac pater eius: " Quis enim es tu? ". Qui respondit: " Ego sum filius tuus primogenitus Esau ".
GEN|27|33|Expavit Isaac stupore vehementi ultra modum et ait: " Quis igitur ille est, qui dudum captam venationem attulit mihi, et comedi ex omnibus, priusquam tu venires? Benedixique ei, et erit benedictus! ".
GEN|27|34|Auditis Esau sermonibus patris, irrugiit clamore magno et amaro ultra modum et ait patri suo: " Benedic etiam mihi, pater mi! ".
GEN|27|35|Qui ait: " Venit germanus tuus fraudulenter et accepit benedictionem tuam ".
GEN|27|36|At ille subiunxit: " Iuste vocatum est nomen eius Iacob; supplantavit enim me en altera vice: primogenita mea ante tulit et nunc secundo surripuit benedictionem meam ".Rursumque ait: " Numquid non reservasti mihi benedictionem? ".
GEN|27|37|Respondit Isaac: " Ecce, dominum tuum illum constitui et omnes fratres eius servituti illius subiugavi; frumento et vino stabilivi eum. Et tibi post haec, fili mi, ultra quid faciam? ".
GEN|27|38|Dixitque Esau ad patrem suum: " Num unam tantum benedictionem habes, pater mi? Mihi quoque obsecro, ut benedicas! ". Cumque eiulatu magno fleret,
GEN|27|39|motus Isaac dixit ad eum: Ecce, procul a pinguedine terrae erit habitatio tuaet procul a rore caeli desuper.
GEN|27|40|De gladio tuo viveset fratri tuo servies.Tempusque veniet, cum excutiaset solvas iugum eius de cervicibus tuis ".
GEN|27|41|Oderat ergo Esau Iacob pro benedictione, qua benedixerat ei pater, dixitque in corde suo: " Appropinquabunt dies luctus patris mei, et occidam Iacob fratrem meum ".
GEN|27|42|Nuntiata sunt Rebeccae verba Esau filii eius maioris, quae mittens et vocans Iacob filium suum minorem dixit ad eum: " Ecce, Esau frater tuus minatur, ut occidat te.
GEN|27|43|Nunc ergo, fili mi, audi vocem meam et consurgens fuge ad Laban fratrem meum in Charran;
GEN|27|44|habitabisque cum eo dies paucos, donec requiescat furor fratris tui,
GEN|27|45|et cesset indignatio eius, obliviscaturque eorum, quae fecisti in eum. Postea mittam et adducam te inde huc. Cur utroque orbabor filio in uno die? ".
GEN|27|46|Dixit quoque Rebecca ad Isaac: " Taedet me vitae meae propter filias Heth; si acceperit Iacob uxorem de filiabus Heth sicut istis de filiabus terrae, nolo vivere ".
GEN|28|1|Vocavit itaque Isaac Iacob et benedixit eum praecepit que ei dicens: " Noli accipere coniugem de filiabus Chanaan;
GEN|28|2|surge, vade in Paddanaram ad domum Bathuel patris matris tuae et accipe tibi inde uxorem de filiabus Laban avunculi tui.
GEN|28|3|Deus autem omnipotens benedicat tibi et crescere te faciat atque multiplicet, ut sis in multitudinem populorum;
GEN|28|4|et det tibi benedictiones Abraham tibi et semini tuo tecum, ut possideas terram peregrinationis tuae, quam pollicitus est Deus avo tuo ".
GEN|28|5|Cumque dimisisset eum Isaac, profectus est in Paddanaram ad Laban filium Bathuel Aramaei fratrem Rebeccae matris Iacob et Esau.
GEN|28|6|Videns autem Esau quod benedixisset pater suus Iacob et misisset eum in Paddanaram, ut inde uxorem duceret, et quod post benedictionem praecepisset ei dicens: " Non accipies uxorem de filiabus Chanaan ",
GEN|28|7|quodque oboediens Iacob parentibus suis isset in Paddanaram;
GEN|28|8|probans quoque quod non libenter aspiceret filias Chanaan pater suus,
GEN|28|9|ivit ad Ismaelem et duxit uxorem, absque iis, quas habebat, Mahalath filiam Ismael filii Abraham sororem Nabaioth.
GEN|28|10|Igitur egressus Iacob de Bersabee pergebat Charran.
GEN|28|11|Cumque venisset ad quendam locum et vellet in eo requiescere post solis occubitum, tulit de lapidibus, qui iacebant, et supponens capiti suo dormivit in eodem loco.
GEN|28|12|Viditque in somnio scalam stantem super terram et cacumen illius tangens caelum, angelos quoque Dei ascendentes et descendentes per eam
GEN|28|13|et Dominum innixum scalae dicentem sibi: " Ego sum Dominus, Deus Abraham patris tui et Deus Isaac. Terram, in qua dormis, tibi dabo et semini tuo.
GEN|28|14|Eritque semen tuum quasi pulvis terrae; dilataberis ad occidentem et orientem et septentrionem et meridiem; et benedicentur in te et in semine tuo cunctae tribus terrae.
GEN|28|15|Et ecce, ego tecum sum et custodiam te, quocumque perrexeris, et reducam te in terram hanc; nec dimittam te, nisi complevero quae dixi tibi.
GEN|28|16|Cumque evigilasset Iacob de somno, ait: " Vere Dominus est in loco isto, et ego nesciebam ".
GEN|28|17|Pavensque: " Quam terribilis est, inquit, locus iste! Non est hic aliud nisi domus Dei et porta caeli ".
GEN|28|18|Surgens ergo Iacob mane tulit lapidem, quem supposuerat capiti suo, et erexit in titulum fundens oleum desuper.
GEN|28|19|Appellavitque nomen loci illius Bethel; prius autem urbs vocabatur Luza.
GEN|28|20|Vovit Iacob etiam votum dicens: " Si fuerit Deus mecum et custodierit me in via hac, per quam ambulo, et dederit mihi panem ad vescendum et vestimentum ad induendum,
GEN|28|21|reversusque fuero prospere ad domum patris mei, erit mihi Dominus in Deum,
GEN|28|22|et lapis iste, quem erexi in titulum, erit domus Dei; cunctorumque, quae dederis mihi, decimas offeram tibi ".
GEN|29|1|Profectus ergo Iacob venit in terram orientalium.
GEN|29|2|Et vidit puteum in agro, tres quoque greges ovium accubantes iuxta eum; nam ex illo adaquabantur pecora, et os eius grandi lapide claudebatur.
GEN|29|3|Morisque erat, ut, cunctis ovibus congregatis, devolverent lapidem et, refectis gregibus, rursum super os putei ponerent.
GEN|29|4|Dixitque ad pastores: " Fratres, unde estis? ". Qui responderunt: " De Charran ".
GEN|29|5|Quos interrogans: " Numquid, ait, nostis Laban filium Nachor? ". Dixerunt: " Novimus ".
GEN|29|6|" Sanusne est? ", inquit. " Valet, inquiunt, et ecce Rachel filia eius venit cum grege ".
GEN|29|7|Dixitque: " Adhuc multum diei superest, nec est tempus, ut congregentur greges; date potum ovibus et sic ad pastum eas reducite ".
GEN|29|8|Qui responderunt: " Non possumus, donec omnia pecora congregentur et amoveamus lapidem de ore putei, ut adaquemus greges ".
GEN|29|9|Adhuc loquebatur cum eis, et ecce Rachel veniebat cum ovibus patris sui; nam gregem ipsa pascebat.
GEN|29|10|Cum vidisset Iacob Rachel filiam Laban avunculi sui ovesque Laban avunculi sui, accedens amovit lapidem de ore putei
GEN|29|11|et adaquavit gregem Laban avunculi sui. Tunc Iacob osculatus est Rachel et elevata voce flevit;
GEN|29|12|et indicavit ei quod frater esset patris eius et filius Rebeccae. At illa festinans nuntiavit patri suo.
GEN|29|13|Qui cum audisset venisse Iacob filium sororis suae, cucurrit obviam ei; complexusque eum et in oscula ruens duxit in domum suam. Auditis autem omnibus, quae evenerant,
GEN|29|14|respondit: " Vere os meum es et caro mea! ".Et, postquam Iacob habitavit apud eum per dies mensis unius,
GEN|29|15|dixit ei Laban: " Num, quia frater meus es, gratis servies mihi? Dic quid mercedis accipias ".
GEN|29|16|Habebat vero filias duas: nomen maioris Lia, minor vero appellabatur Rachel;
GEN|29|17|sed Lia lippis erat oculis, Rachel decora et venusto aspectu.
GEN|29|18|Quam diligens Iacob ait: " Serviam tibi pro Rachel filia tua minore septem annis ".
GEN|29|19|Respondit Laban: " Melius est, ut tibi eam dem quam alteri viro; mane apud me ".
GEN|29|20|Servivit igitur Iacob pro Rachel septem annis, et videbantur illi pauci dies prae amoris magnitudine.
GEN|29|21|Dixitque ad Laban: " Da mihi uxorem meam, quia iam tempus expletum est, ut ingrediar ad eam ".
GEN|29|22|Qui, vocatis omnibus viris loci ad convivium, fecit nuptias.
GEN|29|23|Et vespere sumpsit Liam filiam suam et introduxit ad eum, et venit ad eam.
GEN|29|24|Et dedit Laban ancillam filiae Zelpham nomine.Facto mane, vidit, et ecce erat Lia.
GEN|29|25|Et dixit ad socerum suum: " Quid hoc fecisti mihi? Nonne pro Rachel servivi tibi? Quare imposuisti mihi? ".
GEN|29|26|Respondit Laban: " Non est in loco nostro consuetudinis, ut minorem ante maiorem tradamus ad nuptias.
GEN|29|27|Imple hebdomadam hanc, et alteram quoque dabo tibi pro opere, quo serviturus es mihi septem annis aliis ".
GEN|29|28|Acquievit placito et, hebdomada transacta, dedit ei Laban filiam suam Rachel uxorem,
GEN|29|29|cui servam Bilham tradidit.
GEN|29|30|Et ingressus etiam ad Rachel amavit eam plus quam Liam serviens apud eum septem annis aliis.
GEN|29|31|Videns autem Dominus quod despiceret Liam, aperuit vulvam eius, Rachel sterili permanente.
GEN|29|32|Et concepit Lia et genuit filium vocavitque nomen eius Ruben dicens: " Vidit Dominus humilitatem meam; nunc amabit me vir meus ".
GEN|29|33|Rursumque concepit et peperit filium et ait: " Quoniam audivit me Dominus haberi contemptui, dedit etiam istum mihi "; vocavitque nomen illius Simeon.
GEN|29|34|Concepit tertio et genuit alium filium dixitque: " Nunc quoque copulabitur mihi maritus meus, eo quod pepererim ei tres filios "; et idcirco appellavit nomen eius Levi.
GEN|29|35|Quarto concepit et peperit filium et ait: " Modo confitebor Domino "; et ob hoc vocavit eum Iudam. Cessavitque parere.
GEN|30|1|Cernens autem Rachel quod infecunda esset, invidit sorori et ait marito suo: " Da mihi liberos, alioquin moriar ".
GEN|30|2|Cui iratus respondit Iacob: " Num pro Deo ego sum, qui privavit te fructu ventris? ".
GEN|30|3|At illa: " Ecce, inquit, famula mea Bilha; ingredere ad illam, ut pariat super genua mea, et habeam ex illa et ego filios ".
GEN|30|4|Deditque illi Bilham famulam suam in coniugium. Quae,
GEN|30|5|ingresso ad se Iacob, concepit et peperit filium.
GEN|30|6|Dixitque Rachel: " Iudicavit mihi Deus et exaudivit vocem quoque meam dans mihi filium "; et idcirco appellavit nomen illius Dan.
GEN|30|7|Rursumque Bilha famula Rachel concepit et peperit Iacob alterum filium, et
GEN|30|8|ait Rachel: " Certamina Dei certavi cum sorore mea et invalui "; vocavitque eum Nephthali.
GEN|30|9|Sentiens Lia quod parere desisset, sumpsit Zelpham ancillam suam et tradidit eam Iacob in uxorem.
GEN|30|10|Quae peperit Iacob filium.
GEN|30|11|Dixitque Lia: " Feliciter! "; et idcirco vocavit nomen eius Gad.
GEN|30|12|Peperit quoque Zelpha ancilla Liae Iacob alterum filium.
GEN|30|13|Dixitque Lia: " Pro beatitudine mea! Beatam quippe me dicent mulieres; propterea appellavit eum Aser.
GEN|30|14|Egressus autem Ruben tempore messis triticeae, repperit in agro mandragoras, quas Liae matri suae detulit. Dixitque Rachel: " Da mihi partem de mandragoris filii tui ".
GEN|30|15|Illa respondit: " Parumne tibi videtur, quod praeripueris maritum mihi, ut etiam mandragoras filii mei auferas? ". Ait Rachel: " Dormiat ergo tecum hac nocte pro mandragoris filii tui ".
GEN|30|16|Redeuntique ad vesperam Iacob de agro egressa est in occursum eius Lia et: " Ad me, inquit, intrabis, quia mercede conduxi te pro mandragoris filii mei ". Dormivitque cum ea nocte illa.
GEN|30|17|Et exaudivit Deus Liam, concepitque et peperit Iacob filium quintum
GEN|30|18|et ait: " Dedit Deus mercedem mihi, quia dedi ancillam meam viro meo "; appellavitque nomen illius Issachar.
GEN|30|19|Rursum Lia concepit et peperit Iacob sextum filium
GEN|30|20|et ait: " Donavit me Deus dono bono; hac vice honorabit me maritus meus, eo quod genuerim ei sex filios "; et idcirco appellavit nomen eius Zabulon.
GEN|30|21|Post quem peperit filiam nomine Dinam.
GEN|30|22|Recordatus quoque Deus Rachelis exaudivit eam Deus et aperuit vulvam illius.
GEN|30|23|Quae concepit et peperit filium dicens: " Abstulit Deus opprobrium meum;
GEN|30|24|et vocavit nomen illius Ioseph dicens: " Addat mihi Dominus filium alterum! ".
GEN|30|25|Nato autem Ioseph, dixit Iacob ad Laban: " Dimitte me, ut revertar in patriam et ad terram meam.
GEN|30|26|Da mihi uxores et liberos meos, pro quibus servivi tibi, ut abeam; tu nosti servitutem, qua servivi tibi ".
GEN|30|27|Ait illi Laban: " Inveniam gratiam in conspectu tuo; augurio didici, quia benedixerit mihi Deus propter te.
GEN|30|28|Constitue mercedem tuam, quam dem tibi ".
GEN|30|29|At ille respondit: " Tu nosti quomodo servierim tibi et quanti in manibus meis facti sint greges tui.
GEN|30|30|Modicum habuisti, antequam venirem ad te, et nunc multiplicatum est vehementer, benedixitque tibi Dominus ad introitum meum. Nunc autem quando providebo etiam domui meae? ".
GEN|30|31|Dixitque Laban: " Quid tibi dabo? ". At ille ait: " Nihil mihi dabis; si feceris, quod postulo, iterum pascam et custodiam pecora tua.
GEN|30|32|Gyrabo omnes greges tuos hodie; separa cuncta pecora varia et maculosa et, quodcumque furvum in ovibus et maculosum variumque in capris fuerit, erit merces mea.
GEN|30|33|Respondebitque mihi cras iustitia mea; quando veneris, ut inspicias mercedem meam, omnia, quae non fuerint varia et maculosa in capris et furva in ovibus, furti me arguent ".
GEN|30|34|Dixit Laban: " Gratum habeo, quod petis! ".
GEN|30|35|Et separavit in die illo hircos striatos atque maculosos et omnes capras varias et maculosas, omne, in quo album erat, et omne furvum in ovibus, et tradidit in manu filiorum suorum.
GEN|30|36|Et posuit spatium itineris trium dierum inter se et Iacob, qui pascebat reliquos greges Laban.
GEN|30|37|Tollens ergo Iacob virgas virides populeas et amygdalinas et ex platanis, ex parte ita decorticavit eas, ut in his, quae spoliata fuerant, candor appareret.
GEN|30|38|Posuitque virgas, quas ex parte decorticaverat, in canalibus, ubi effundebatur aqua, ut, cum venissent greges ad bibendum, ante oculos haberent virgas et in aspectu earum conciperent.
GEN|30|39|Factumque est ut in ipso calore coitus greges intuerentur virgas et parerent striata et varia et maculosa.
GEN|30|40|Agnos autem segregavit Iacob et posuit gregem ex adverso striatorum et omnium furvorum in grege Laban et constituit sibi greges seorsum neque statuit eos cum grege Laban.
GEN|30|41|Quotiescumque igitur calefiebant pecora robusta, ponebat Iacob virgas in canalibus aquarum ante oculos pecorum, ut in earum contemplatione conciperent.
GEN|30|42|Quando vero pecora debilia erant, non ponebat eas. Factaque sunt debilia Laban et robusta Iacob;
GEN|30|43|ditatusque est homo ultra modum et habuit greges multos, ancillas et servos, camelos et asinos.
GEN|31|1|Postquam autem audivit verba filiorum Laban dicen tium: " Tulit Iacob omnia, quae fuerunt patris nostri, et de patris nostri facultate acquisivit has divitias ",
GEN|31|2|animadvertit quoque faciem Laban quod non esset erga se sicut heri et nudiustertius.
GEN|31|3|Et dixit Dominus ad Iacob: " Revertere in terram patrum tuorum et ad cognationem tuam, eroque tecum ".
GEN|31|4|Misit Iacob et vocavit Rachel et Liam in agrum, ubi pascebat greges,
GEN|31|5|dixitque eis: " Video faciem patris vestri quod non sit erga me sicut heri et nudiustertius; Deus autem patris mei fuit mecum,
GEN|31|6|et ipsae nostis quod totis viribus meis servierim patri vestro.
GEN|31|7|Sed pater vester circumvenit me et mutavit mercedem meam decem vicibus; et tamen non dimisit eum Deus, ut noceret mihi.
GEN|31|8|Si quando dixit: "Variae erunt mercedes tuae", pariebant omnes oves varios fetus. Quando vero e contrario ait: "Striata quaeque accipies pro mercede", omnes greges striata pepererunt.
GEN|31|9|Tulitque Deus substantiam patris vestri et dedit mihi.
GEN|31|10|Postquam enim conceptus gregis tempus advenerat, levavi oculos meos et vidi in somnis ascendentes mares super feminas, striatos et varios et respersos.
GEN|31|11|Dixitque angelus Dei ad me in somnis: "Iacob". Et ego respondi: Adsum.
GEN|31|12|Qui ait: "Leva oculos tuos et vide universos masculos ascendentes super feminas, striatos et varios atque respersos. Vidi enim omnia, quae fecit tibi Laban.
GEN|31|13|Ego sum Deus Bethel, ubi unxisti lapidem et votum vovisti mihi. Nunc ergo surge et egredere de terra hac revertens in terram nativitatis tuae".
GEN|31|14|Responderunt ei Rachel et Lia: " Numquid habemus adhuc partem et hereditatem in domo patris nostri?
GEN|31|15|Nonne quasi alienas reputavit nos et vendidit nos comeditque pretium nostrum?
GEN|31|16|Sed omnes opes, quas tulit Deus patri nostro, nobis abstulit ac filiis nostris; unde omnia, quae praecepit tibi Deus, fac ".
GEN|31|17|Surrexit itaque Iacob et imposuit liberos suos ac coniuges suas super camelos.
GEN|31|18|Tulitque omnes greges suos et omnem substantiam suam, quidquid in Paddanaram acquisierat, ut iret ad Isaac patrem suum in terram Chanaan.
GEN|31|19|Eo tempore Laban ierat ad tondendas oves, et Rachel furata est theraphim patris sui.
GEN|31|20|Iacob autem decepit cor Laban, non indicans ei quod fugeret.
GEN|31|21|Cumque fugisset cum omnibus, quae possidebat, et, amne transmisso, pergeret contra montem Galaad,
GEN|31|22|nuntiatum est Laban die tertio quod fugisset Iacob.
GEN|31|23|Qui, assumptis fratribus suis, persecutus est eum diebus septem et comprehendit eum in monte Galaad.
GEN|31|24|Venit autem Deus ad Laban Aramaeum per somnium noctis dixitque ei: Cave, ne quidquam loquaris contra Iacob!".
GEN|31|25|Iamque Iacob extenderat in monte tabernaculum, cum Laban, consecutus eum cum fratribus suis, in eodem monte Galaad fixit tentorium.
GEN|31|26|Et dixit ad Iacob: " Quare ita egisti et decepisti cor meum, abigens filias meas quasi captivas gladio?
GEN|31|27|Cur clam fugisti et decepisti me, non indicans mihi, ut prosequerer te cum gaudio et canticis et tympanis et citharis?
GEN|31|28|Non es passus, ut oscularer filios meos ac filias; stulte operatus es. Et nunc
GEN|31|29|valet quidem manus mea reddere tibi malum, sed Deus patris vestri heri dixit mihi: "Cave, ne loquaris contra Iacob quidquam!".
GEN|31|30|Esto, profectus es, quia desiderio tibi erat domus patris tui; cur furatus es deos meos? ".
GEN|31|31|Respondit Iacob: " Quia timui. Dixi enim, ne forte violenter auferres filias tuas a me.
GEN|31|32|Apud quemcumque inveneris deos tuos, non vivat! Coram fratribus nostris scrutare, quidquid tuorum apud me inveneris, et aufer ". Ignorabat enim Iacob quod Rachel furata esset theraphim.
GEN|31|33|Ingressus itaque Laban tabernacula Iacob et Liae et utriusque famulae, non invenit. Egressus de tentorio Liae, intravit tentorium Rachelis.
GEN|31|34|Illa autem absconderat theraphim in stramento cameli et sedit desuper. Scrutantique omne tentorium et nihil invenienti
GEN|31|35|ait: " Ne irascatur dominus meus, quod coram te assurgere nequeo, quia iuxta consuetudinem feminarum nunc accidit mihi ". Quaesivit ergo et non invenit theraphim.
GEN|31|36|Tumensque Iacob cum iurgio ait: " Quam ob culpam meam et ob quod peccatum meum sic persecutus es me,
GEN|31|37|quia scrutatus es omnem supellectilem meam? Quid invenisti de cuncta substantia domus tuae? Pone hic coram fratribus meis et fratribus tuis, et iudicent inter me et te.
GEN|31|38|Ecce, viginti annis fui tecum. Oves tuae et caprae non abortiverunt, arietes gregis tui non comedi;
GEN|31|39|nec dilaceratum a bestia ostendi tibi: ego damnum omne reddebam; quidquid die noctuque furto perierat, a me exigebas.
GEN|31|40|Die aestu consumebar et nocte gelu, fugiebatque somnus ab oculis meis.
GEN|31|41|Sic per viginti annos in domo tua servivi tibi: quattuordecim pro filiabus et sex pro gregibus tuis; immutasti quoque mercedem meam decem vicibus.
GEN|31|42|Nisi Deus patris mei, Deus Abraham et Timor Isaac, affuisset mihi, certemodo nudum me dimisisses; afflictionem meam et laborem manuum mearum respexit Deus et iudicavit heri ".
GEN|31|43|Respondit ei Laban: " Filiae filiae meae et filii filii mei et greges greges mei et omnia, quae cernis, mea sunt; et filiabus meis quid possum facere illis hodie et filiis earum, quos genuerunt?
GEN|31|44|Veni ergo, et ineamus foedus ego et tu, ut sit in testimonium inter me et te ".
GEN|31|45|Tulit itaque Iacob lapidem et erexit illum in titulum;
GEN|31|46|dixitque fratribus suis: " Afferte lapides ". Qui congregantes fecerunt tumulum comederuntque ibi super eum.
GEN|31|47|Quem vocavit Laban Iegarsahadutha (id est Tumulus testimonii), et Iacob Galed (uterque iuxta proprietatem linguae suae).
GEN|31|48|Dixitque Laban: " Tumulus iste testis erit inter me et te hodie "; et idcirco appellatum est nomen eius Galed (id est Tumulus testis)
GEN|31|49|et etiam Maspha (id est Specula), quia dixit: " Speculetur Dominus inter me et te, quando absconditi erimus ab invicem.
GEN|31|50|Si afflixeris filias meas et si introduxeris uxores alias super eas, cum nemo nobiscum sit, vide, Deus est testis inter me et te ".
GEN|31|51|Dixitque Laban ad Iacob: " En tumulus hic et lapis, quem erexi inter me et te.
GEN|31|52|Testis erit tumulus iste et lapis quod ego non transibo tumulum hunc pergens ad te, neque tu transibis tumulum hunc et lapidem hunc ad malum.
GEN|31|53|Deus Abraham et Deus Nachor iudicent inter nos ".Iuravit Iacob per Timorem patris sui Isaac;
GEN|31|54|immolatisque victimis in monte, vocavit fratres suos, ut ederent panem. Qui cum comedissent, pernoctaverunt in monte.
GEN|32|1|Laban vero de nocte consur gens osculatus est filios et fi lias suas et benedixit illis reversusque est in locum suum.
GEN|32|2|Iacob quoque abiit itinere, quo coeperat, fueruntque ei obviam angeli Dei.
GEN|32|3|Quos cum vidisset, ait: " Castra Dei sunt haec "; et appellavit nomen loci illius Mahanaim (id est Castra).
GEN|32|4|Misit autem nuntios ante se ad Esau fratrem suum in terram Seir, in regionem Edom.
GEN|32|5|Praecepitque eis dicens: " Sic loquimini domino meo Esau: Haec dicit servus tuus Iacob: Apud Laban peregrinatus sum et fui usque in praesentem diem.
GEN|32|6|Habeo boves et asinos, oves et servos atque ancillas; mittoque nunc legationem ad dominum meum, ut inveniam gratiam in conspectu tuo ".
GEN|32|7|Reversique sunt nuntii ad Iacob dicentes: " Venimus ad Esau fratrem tuum, et ecce properat in occursum tibi cum quadringentis viris ".
GEN|32|8|Timuit Iacob valde et perterritus divisit populum, qui secum erat, greges quoque et oves et boves et camelos in duas turmas
GEN|32|9|dicens: " Si venerit Esau ad unam turmam et percusserit eam, alia turma, quae reliqua est, salvabitur ".
GEN|32|10|Dixitque Iacob: " Deus patris mei Abraham et Deus patris mei Isaac, Domine, qui dixisti mihi: "Revertere in terram tuam et in locum nativitatis tuae, et benefaciam tibi",
GEN|32|11|minor sum cunctis miserationibus et cuncta veritate, quam explesti servo tuo. In baculo meo transivi Iordanem istum et nunc cum duabus turmis regredior.
GEN|32|12|Erue me de manu fratris mei, de manu Esau, quia valde eum timeo; ne forte veniens percutiat matrem cum filiis.
GEN|32|13|Tu locutus es quod bene mihi faceres et dilatares semen meum sicut arenam maris, quae prae multitudine numerari non potest ".
GEN|32|14|Mansit ibi nocte illa et sumpsit de his, quae habebat, munera Esau fratri suo:
GEN|32|15|capras ducentas, hircos viginti, oves ducentas et arietes viginti,
GEN|32|16|camelos fetas cum pullis suis triginta, vaccas quadraginta et tauros decem, asinas viginti et pullos earum decem.
GEN|32|17|Et misit per manus servorum suorum singulos seorsum greges dixitque pueris suis: " Antecedite me, et sit spatium inter gregem et gregem ".
GEN|32|18|Et praecepit priori dicens: " Si obvium habueris Esau fratrem meum, et interrogaverit te: "Cuius es?" et "Quo vadis?" et "Cuius sunt ista, quae sequeris?",
GEN|32|19|respondebis: Servi tui Iacob; munera misit domino meo Esau. Ipse quoque post nos venit ".
GEN|32|20|Similiter mandata dedit secundo ac tertio et cunctis, qui sequebantur greges, dicens: " Iisdem verbis loquimini ad Esau, cum inveneritis eum,
GEN|32|21|et addetis: Ipse quoque servus tuus Iacob iter nostrum insequitur. Dixit enim: Placabo illum muneribus, quae praecedunt, et postea videbo faciem eius: forsitan propitiabitur mihi ".
GEN|32|22|Praecesserunt itaque munera ante eum, ipse vero mansit nocte illa in castris.
GEN|32|23|Cumque nocte surrexisset, tulit duas uxores suas et totidem famulas cum undecim filiis et transivit vadum Iaboc;
GEN|32|24|sumptis ergo traductisque illis et omnibus, quae ad se pertinebant, per torrentem,
GEN|32|25|mansit solus.Et ecce vir luctabatur cum eo usque mane.
GEN|32|26|Qui cum videret quod eum superare non posset, tetigit acetabulum femoris eius, et statim luxatum est acetabulum femoris Iacob, cum luctaretur cum illo.
GEN|32|27|Dixitque: " Dimitte me, iam enim ascendit aurora ". Respondit: " Non dimittam te, nisi benedixeris mihi ".
GEN|32|28|Ait ad eum: " Quod nomen est tibi? ". Respondit: " Iacob ".
GEN|32|29|At ille: " Nequaquam, inquit, Iacob amplius appellabitur nomen tuum, sed Israel: quoniam certasti cum Deo et cum hominibus et praevaluisti! ".
GEN|32|30|Interrogavit eum Iacob: " Dic mihi, quo appellaris nomine? ". Respondit: " Cur quaeris nomen meum? ". Et benedixit ei in eodem loco.
GEN|32|31|Vocavitque Iacob nomen loci illius Phanuel dicens: " Vidi Deum facie ad faciem, et salva facta est anima mea ".
GEN|32|32|Ortusque est ei sol, cum transgrederetur Phanuel; ipse vero claudicabat propter femur.
GEN|32|33|Quam ob causam non comedunt filii Israel nervum, qui est in femore, usque in praesentem diem, eo quod tetigerit nervum femoris Iacob.
GEN|33|1|Elevans autem Iacob oculos suos vidit venientem Esau et cum eo quadringentos viros; divisitque filios Liae et Rachel ambarumque famularum.
GEN|33|2|Et posuit utramque ancillam et liberos earum in principio, Liam vero et filios eius in secundo loco, Rachel autem et Ioseph novissimos.
GEN|33|3|Et ipse praegrediens adoravit pronus in terram septies, donec appropinquaret ad fratrem suum.
GEN|33|4|Currens itaque Esau obviam fratri suo amplexatus est eum; stringensque collum eius osculatus est eum, et fleverunt.
GEN|33|5|Levatisque oculis, vidit mulieres et liberos earum et ait: " Qui sunt isti tibi? ". Respondit: " Liberi sunt, quos donavit mihi Deus servo tuo.
GEN|33|6|Et appropinquantes ancillae et filii earum incurvati sunt.
GEN|33|7|Accessit quoque Lia cum liberis suis et, cum similiter adorassent, extremi Ioseph et Rachel adoraverunt.
GEN|33|8|" Quaenam sunt, inquit, istae turmae, quas obvias habui? ". Respondit: " Ut invenirem gratiam coram domino meo ".
GEN|33|9|At ille: " Habeo, ait, plurima, frater mi; sint tua tibi ".
GEN|33|10|Dixit Iacob: " Noli ita, obsecro; sed, si inveni gratiam in oculis tuis, accipe munusculum de manibus meis; sic enim vidi faciem tuam quasi viderim vultum Dei, et mihi propitius fuisti.
GEN|33|11|Suscipe, quaeso, benedictionem, quae allata est tibi; quia Deus misertus est mihi, et habeo omnia ".Et, cum compelleret illum, suscepit
GEN|33|12|et ait: " Gradiamur simul, eroque socius itineris tui ".
GEN|33|13|Dixit Iacob: " Nosti, domine mi, quod parvulos habeam teneros et oves et boves fetas mecum; quas si plus in ambulando fecero laborare vel una die, morientur cuncti greges.
GEN|33|14|Praecedat dominus meus ante servum suum; et ego sequar paulatim secundum gressum pecorum ante me et secundum gressum parvulorum, donec veniam ad dominum meum in Seir ".
GEN|33|15|Respondit Esau: " Oro te, ut de populo, qui mecum est, saltem socii remaneant viae tuae". " Non est, inquit, necesse; hoc uno indigeo, ut inveniam gratiam in conspectu domini mei ".
GEN|33|16|Reversus est itaque illo die Esau itinere suo in Seir.
GEN|33|17|Et Iacob venit in Succoth, ubi, aedificata sibi domo et fixis tentoriis pro gregibus suis, appellavit nomen loci illius Succoth (id est Tabernacula).
GEN|33|18|Transivitque Iacob incolumis ad urbem Sichem, quae est in terra Chanaan, cum veniret de Paddanaram; et habitavit iuxta oppidum.
GEN|33|19|Emitque partem agri, in qua fixerat tabernaculum suum, a filiis Hemmor patris Sichem centum argenteis.
GEN|33|20|Et erexit ibi altare et vocavit illud: " Deus est Deus Israel ".
GEN|34|1|Egressa est autem Dina filia, quam Lia pepererat Iacob, ut videret filias regionis illius.
GEN|34|2|Quam cum vidisset Sichem filius Hemmor Hevaei principis terrae illius, adamavit eam et rapuit; et dormivit cum illa, vi opprimens illam.
GEN|34|3|Et conglutinata est anima eius cum ea, et amavit puellam et locutus est ad cor eius.
GEN|34|4|Dixitque ad Hemmor patrem suum: " Accipe mihi puellam hanc coniugem ".
GEN|34|5|Cum audisset Iacob quod violasset Dinam filiam suam, absentibus filiis et in pastu pecorum occupatis, siluit, donec redirent.
GEN|34|6|Egresso autem Hemmor patre Sichem, ut loqueretur ad Iacob,
GEN|34|7|ecce filii Iacob veniebant de agro, auditoque, quod acciderat, contristati et irati sunt valde, eo quod foedam rem esset operatus in Israel et, violata filia Iacob, rem illicitam perpetrasset.
GEN|34|8|Locutus est itaque Hemmor ad eos: " Sichem filii mei adhaesit anima filiae vestrae; date eam illi uxorem,
GEN|34|9|et iungamus vicissim conubia: filias vestras tradite nobis et filias nostras accipite vobis.
GEN|34|10|Et habitate nobiscum; terra in potestate vestra est: manete, perambulate et possidete eam ".
GEN|34|11|Sed et Sichem ad patrem et ad fratres eius ait: " Inveniam gratiam coram vobis et, quaecumque statueritis, dabo.
GEN|34|12|Augete mihi valde dotem et munera; libens tribuam, quod petieritis. Tantum date mihi puellam hanc uxorem ".
GEN|34|13|Responderunt filii Iacob Sichem et Hemmor patri eius in dolo ob stuprum sororis:
GEN|34|14|" Non possumus facere, quod petitis, dare sororem nostram homini incircumciso, opprobrium enim esset nobis.
GEN|34|15|In hoc tantum valebimus acquiescere vobis: si esse volueritis similes nostri, circumcidatur in vobis omne masculini sexus;
GEN|34|16|tunc dabimus et accipiemus mutuo filias nostras ac vestras et habitabimus vobiscum erimusque unus populus.
GEN|34|17|Si autem circumcidi nolueritis, tollemus filiam nostram et recedemus ".
GEN|34|18|Placuit oblatio eorum Hemmor et Sichem filio eius,
GEN|34|19|nec distulit adulescens quin statim, quod petebatur, expleret; amabat enim filiam Iacob valde, et ipse erat inclitus in omni domo patris sui.
GEN|34|20|Ingressique portam urbis, Hemmor et Sichem filius eius locuti sunt ad viros civitatis suae:
GEN|34|21|" Viri isti pacifici sunt erga nos; maneant in terra et perambulent eam, quae spatiosa et lata est eis; filias eorum accipiemus uxores et nostras illis dabimus.
GEN|34|22|Tantum in hoc valebunt viri acquiescere nobis, ut maneant nobiscum et efficiamur unus populus, si circumcidamus masculos nostros ritum gentis imitantes;
GEN|34|23|et pecora et substantia et armenta eorum nostra erunt. Tantum in hoc acquiescamus, et habitabunt nobiscum ".
GEN|34|24|Assensique sunt omnes, circumcisis cunctis maribus, qui egrediebantur e porta civitatis suae.
GEN|34|25|Et ecce, die tertio, quando gravissimus vulnerum dolor est, arreptis duo filii Iacob Simeon et Levi fratres Dinae gladiis, ingressi sunt urbem securi; interfectisque omnibus masculis,
GEN|34|26|Hemmor et Sichem pariter necaverunt, tollentes Dinam de domo Sichem sororem suam.
GEN|34|27|Filii Iacob irruerunt super occisos, et depopulati sunt urbem in ultionem stupri.
GEN|34|28|Oves eorum et armenta et asinos cunctaque, quae in civitate et in agris erant, tulerunt.
GEN|34|29|Omnes opes eorum, parvulos quoque et uxores duxerunt captivas et diripuerunt omnia, quae in domibus erant.
GEN|34|30|Iacob autem dixit ad Simeon et Levi: " Turbastis me et odiosum fecistis me Chananaeis et Pherezaeis habitatoribus terrae huius. Nos pauci sumus; illi congregati percutient me, et delebor ego et domus mea ".
GEN|34|31|Responderunt: " Numquid ut scorto abuti debuere sorore nostra? ".
GEN|35|1|Locutus est Deus ad Iacob: " Surge et ascende Bethel et habita ibi; facque altare Deo, qui apparuit tibi, quando fugiebas Esau fratrem tuum ".
GEN|35|2|Iacob vero, convocata omni domo sua, ait: " Abigite deos alienos, qui in medio vestri sunt, et mundamini ac mutate vestimenta vestra.
GEN|35|3|Surgamus et ascendamus in Bethel, ut faciamus ibi altare Deo, qui exaudivit me in die tribulationis meae et socius fuit itineris mei ".
GEN|35|4|Dederunt ergo ei omnes deos alienos, quos habebant, et inaures, quae erant in auribus eorum; at ille infodit ea subter Quercum, quae est prope urbem Sichem.
GEN|35|5|Cumque profecti essent, terror Dei invasit omnes per circuitum civitates, et non sunt ausi persequi filios Iacob.
GEN|35|6|Venit igitur Iacob Luzam, quae est in terra Chanaan, id est Bethel, ipse et omnis populus cum eo.
GEN|35|7|Aedificavitque ibi altare et appellavit nomen loci illius Deus Bethel; ibi enim apparuit ei Deus, cum fugeret fratrem suum.
GEN|35|8|Eodem tempore mortua est Debora nutrix Rebeccae et sepulta est ad radices Bethel subter quercum; vocatumque est nomen loci illius Quercus fletus.
GEN|35|9|Apparuit iterum Deus Iacob, postquam reversus est de Paddanaram, benedixitque ei
GEN|35|10|dicens: " Non vocaberis ultra Iacob, sed Israel erit nomen tuum ", et appellavit eum Israel.
GEN|35|11|Dixitque ei: " Ego Deus omnipotens. Cresce et multiplicare; gens et congregatio nationum erunt ex te, reges de lumbis tuis egredientur.
GEN|35|12|Terramque, quam dedi Abraham et Isaac, dabo tibi; et semini tuo post te dabo terram hanc ".
GEN|35|13|Et ascendit ab eo Deus.
GEN|35|14|Ille vero erexit titulum lapideum in loco, quo locutus ei fuerat Deus, libans super eum libamina et effundens oleum
GEN|35|15|vocansque nomen loci illius Bethel.
GEN|35|16|Egressi sunt de Bethel. Et adhuc spatium quoddam erat usque ad Ephratham, cum parturiret Rachel;
GEN|35|17|ob difficultatem partus periclitari coepit, dixitque ei obstetrix: " Noli timere, quia et hac vice habes filium ".
GEN|35|18|Egrediente autem anima et imminente iam morte, vocavit nomen filii sui Benoni (id est Filius doloris mei); pater vero appellavit eum Beniamin (id est Filius dextrae).
GEN|35|19|Mortua est ergo Rachel et sepulta est in via, quae ducit Ephratham; haec est Bethlehem.
GEN|35|20|Erexitque Iacob titulum super sepulcrum eius; hic est titulus monumenti Rachel usque in praesentem diem.
GEN|35|21|Egressus inde Israel, fixit tabernaculum trans Magdaleder (id est Turris gregis).
GEN|35|22|Cumque habitaret in illa regione, abiit Ruben et dormivit cum Bilha concubina patris sui; quod illum minime latuit.Erant autem filii Iacob duodecim.
GEN|35|23|Filii Liae: primogenitus Ruben et Simeon et Levi et Iudas et Issachar et Zabulon.
GEN|35|24|Filii Rachel: Ioseph et Beniamin.
GEN|35|25|Filii Bilhae ancillae Rachelis: Dan et Nephthali.
GEN|35|26|Filii Zelphae ancillae Liae: Gad et Aser. Hi sunt filii Iacob, qui nati sunt ei in Paddanaram.
GEN|35|27|Venit Iacob ad Isaac patrem suum in Mambre Cariatharbe, id est Hebron, ubi peregrinatus est Abraham et Isaac.
GEN|35|28|Et completi sunt dies Isaac centum octoginta annorum;
GEN|35|29|consumptusque aetate mortuus est et appositus est populo suo senex et plenus dierum. Et sepelierunt eum Esau et Iacob filii sui.
GEN|36|1|Hae sunt autem generationes Esau. Ipse est Edom.
GEN|36|2|Esau accepit uxores de filiabus Chanaan: Ada filiam Elon Hetthaei et Oolibama filiam Ana filii Sebeon Horraei;
GEN|36|3|Basemath quoque filiam Ismael sororem Nabaioth.
GEN|36|4|Peperit autem Ada Eliphaz, Basemath genuit Rahuel,
GEN|36|5|Oolibama genuit Iehus et Ialam et Core.Hi filii Esau, qui nati sunt ei in terra Chanaan.
GEN|36|6|Tulit autem Esau uxores suas et filios et filias et omnes animas domus suae et pecora armenta et cuncta, quae acquisierat in terra Chanaan, et abiit in terram Seir; recessitque a fratre suo Iacob.
GEN|36|7|Divites enim erant valde et simul habitare non poterant; nec sustinebat eos terra peregrinationis eorum prae multitudine gregum.
GEN|36|8|Habitavitque Esau in monte Seir. Ipse est Edom.
GEN|36|9|Hae autem sunt generationes Esau patris Edom in monte Seir,
GEN|36|10|et haec nomina filiorum eius: Eliphaz filius Ada uxoris Esau, Rahuel quoque filius Basemath uxoris eius.
GEN|36|11|Fueruntque Eliphaz filii: Theman, Omar, Sepho et Gatham et Cenez.
GEN|36|12|Erat autem Thamna concubina Eliphaz filii Esau, quae peperit ei Amalec. Hi sunt filii Ada uxoris Esau.
GEN|36|13|Filii autem Rahuel: Nahath et Zara, Samma et Meza; hi filii Basemath uxoris Esau.
GEN|36|14|Isti erant filii Oolibama filiae Ana filii Sebeon uxoris Esau, quos genuit ei: Iehus et Ialam et Core.
GEN|36|15|Hi duces filiorum Esau. Filii Eliphaz primogeniti Esau: dux Theman, dux Omar, dux Sepho, dux Cenez,
GEN|36|16|dux Core, dux Gatham, dux Amalec. Hi duces Eliphaz in terra Edom; hi filii Ada.
GEN|36|17|Hi filii Rahuel filii Esau: dux Nahath, dux Zara, dux Samma, dux Meza. Hi duces Rahuel in terra Edom; isti filii Basemath uxoris Esau.
GEN|36|18|Hi filii Oolibama uxoris Esau: dux Iehus, dux Ialam, dux Core. Hi duces Oolibama filiae Ana uxoris Esau.
GEN|36|19|Isti sunt filii Esau et hi duces eorum. Ipse est Edom.
GEN|36|20|Isti sunt filii Seir Horraei habitatores terrae: Lotan et Sobal et Sebeon et Ana
GEN|36|21|et Dison et Eser et Disan; hi duces Horraei filii Seir in terra Edom.
GEN|36|22|Facti sunt autem filii Lotan: Hori et Hemam; erat autem soror Lotan Thamna.
GEN|36|23|Et isti filii Sobal: Alvan et Manahath et Ebal, Sepho et Onam.
GEN|36|24|Et hi filii Sebeon: Aia et Ana. Iste est Ana, qui invenit aquas calidas in solitudine, cum pasceret asinos Sebeon patris sui.
GEN|36|25|Habuitque filium Dison et filiam Oolibama.
GEN|36|26|Et isti filii Dison: Hemdan et Eseban et Iethran et Charran.
GEN|36|27|Hi filii Eser: Bilhan et Zavan et Iacan.
GEN|36|28|Habuit autem filios Disan: Us et Aran.
GEN|36|29|Isti duces Horraeorum: dux Lotan, dux Sobal, dux Sebeon, dux Ana,
GEN|36|30|dux Dison, dux Eser, dux Disan; isti duces Horraeorum secundum tribus eorum in terra Seir.
GEN|36|31|Reges autem, qui regnaverunt in terra Edom, antequam haberent regem filii Israel, fuerunt hi.
GEN|36|32|Regnavit in Edom Bela filius Beor, nomenque urbis eius Denaba.
GEN|36|33|Mortuus est autem Bela, et regnavit pro eo Iobab filius Zarae de Bosra.
GEN|36|34|Cumque mortuus esset Iobab, regnavit pro eo Husam de terra Themanorum.
GEN|36|35|Hoc quoque mortuo, regnavit pro eo Adad filius Badad, qui percussit Madian in regione Moab; et nomen urbis eius Avith.
GEN|36|36|Cumque mortuus esset Adad, regnavit pro eo Semla de Masreca.
GEN|36|37|Hoc quoque mortuo, regnavit pro eo Saul de Rohoboth iuxta fluvium.
GEN|36|38|Cumque et hic obiisset, successit in regnum Baalhanan filius Achobor.
GEN|36|39|Isto quoque mortuo, regnavit pro eo Adad, nomenque urbis eius Phau; et appellabatur uxor eius Meetabel filia Matred filiae Mezaab.
GEN|36|40|Haec ergo nomina ducum Esau in cognationibus et locis et vocabulis suis: dux Thamna, dux Alva, dux Ietheth,
GEN|36|41|dux Oolibama, dux Ela, dux Phinon,
GEN|36|42|dux Cenez, dux Theman, dux Mabsar,
GEN|36|43|dux Magdiel, dux Iram.Hi duces Edom habitantes in terra imperii sui. Ipse est Esau pater Idumaeorum.
GEN|37|1|Habitavit autem Iacob in terra Chanaan, in qua pere grinatus est pater suus.
GEN|37|2|Hae sunt generationes Iacob.Ioseph, cum decem et scptem esset annorum, pascebat gregem cum fratribus suis adhuc puer; et erat cum filiis Bilhae et Zelphae uxorum patris sui; detulitque patri malam eorum famam.
GEN|37|3|Israel autem diligebat Ioseph super omnes filios suos, eo quod in senectute genuisset eum; fecitque ei tunicam talarem.
GEN|37|4|Videntes autem fratres eius quod a patre plus cunctis filiis amaretur, oderant eum nec poterant ei quidquam pacifice loqui.
GEN|37|5|Accidit quoque ut visum somnium referret fratribus suis; quae causa maioris odii seminarium fuit.
GEN|37|6|Dixitque ad eos: " Audite somnium meum, quod vidi.
GEN|37|7|Putabam ligare nos manipulos in agro, et quasi consurgere manipulum meum et stare, vestrosque manipulos circumstantes adorare manipulum meum ".
GEN|37|8|Responderunt fratres eius: " Numquid rex noster eris? Aut subiciemur dicioni tuae? ". Haec ergo causa somniorum atque sermonum, invidiae et odii fomitem ministravit.
GEN|37|9|Aliud quoque vidit somnium, quod narrans fratribus ait: " Vidi per somnium quasi solem et lunam et stellas undecim adorare me ".
GEN|37|10|Quod cum patri suo et fratribus retulisset, increpavit eum pater suus et dixit: " Quid sibi vult hoc somnium, quod vidisti? Num ego et mater tua et fratres tui adorabimus te proni in terram? ".
GEN|37|11|Invidebant igitur ei fratres sui; pater vero rem tacitus considerabat.
GEN|37|12|Cumque fratres illius in pascendis gregibus patris morarentur in Sichem,
GEN|37|13|dixit Israel ad Ioseph: " Fratres tui pascunt oves in Sichimis; veni, mittam te ad eos ". Quo respondente:
GEN|37|14|" Praesto sum ", ait ei: " Vade et vide, si cuncta prospera sint erga fratres tuos et pecora, et renuntia mihi quid agatur ". Missus de valle Hebron venit in Sichem;
GEN|37|15|invenitque eum vir errantem in agro et interrogavit quid quaereret.
GEN|37|16|At ille respondit: " Fratres meos quaero; indica mihi, ubi pascant greges ".
GEN|37|17|Dixitque ei vir: " Recesserunt de loco isto; audivi autem eos dicentes: Eamus in Dothain" ". Perrexit ergo Ioseph post fratres suos et invenit eos in Dothain.
GEN|37|18|Qui cum vidissent eum procul, antequam accederet ad eos, cogitaverunt illum occidere.
GEN|37|19|Et mutuo loquebantur: " Ecce somniator venit;
GEN|37|20|venite, occidamus eum et mittamus in unam cisternarum dicemusque: Fera pessima devoravit eum. Et tunc apparebit quid illi prosint somnia sua ".
GEN|37|21|Audiens autem hoc Ruben nitebatur liberare eum de manibus eorum et dixit:
GEN|37|22|" Non interficiamus animam eius ". Et dixit ad eos: " Non effundatis sanguinem; sed proicite eum in cisternam hanc, quae est in solitudine, manusque vestras servate innoxias ". Hoc autem dicebat volens eripere eum de manibus eorum et reddere patri suo.
GEN|37|23|Confestim igitur, ut pervenit ad fratres suos, nudaverunt eum tunica talari
GEN|37|24|miseruntque eum in cisternam, quae non habebat aquam.
GEN|37|25|Et sederunt, ut comederent panem. Attollentes autem oculos viderunt Ismaelitas viatorcs venire de Galaad et camelos eorum portantes tragacanthum et masticem et ladanum in Aegyptum.
GEN|37|26|Dixit ergo Iudas fratribus suis: " Quid nobis prodest, si occiderimus fratrem nostrum et celaverimus sanguinem ipsius?
GEN|37|27|Melius est ut vendatur Ismaelitis, et manus nostrae non polluantur; frater enim et caro nostra est ". Acquieverunt fratres sermonibus illius.
GEN|37|28|Et praetereuntibus Madianitis negotiatoribus, extrahentes Ioseph de cisterna, vendiderunt eum Ismaelitis viginti argenteis. Qui duxerunt eum in Aegyptum.
GEN|37|29|Reversusque Ruben ad cisternam non invenit puerum
GEN|37|30|et, scissis vestibus, pergens ad fratres suos ait: " Puer non comparet, et ego quo ibo? ".
GEN|37|31|Tulerunt autem tunicam eius et in sanguinem haedi, quem occiderant, tinxerunt
GEN|37|32|mittentes, qui ferrent ad patrem et dicerent: "Hanc invenimus; vide, utrum tunica talaris filii tui sit an non? ".
GEN|37|33|Quam cum agnovisset pater, ait: " Tunica filii mei est; fera pessima comedit eum, bestia devoravit Ioseph ".
GEN|37|34|Scissisque vestibus, indutus est cilicio lugens filium suum multo tempore.
GEN|37|35|Congregatis autem cunctis liberis eius, ut lenirent dolorem patris, noluit consolationem accipere et ait: " Descendam ad filium meum lugens in infernum ". Et flevit super eo pater eius.
GEN|37|36|Madianitae autem vendiderunt Ioseph in Aegypto Putiphari eunucho pharaonis, magistro satellitum.
GEN|38|1|Eo tempore descendens Iudas a fratribus suis divertit ad virum Odollamitem nomine Hiram.
GEN|38|2|Viditque ibi filiam hominis Chananaei vocabulo Sue et, accepta uxore, ingressus est ad eam.
GEN|38|3|Quae concepit et peperit filium vocavitque nomen eius Her.
GEN|38|4|Rursumque concepto fetu, natum filium nominavit Onan.
GEN|38|5|Tertium quoque peperit, quem appellavit Sela. Ipsa autem erat in Chasib, quando peperit illum.
GEN|38|6|Dedit autem Iudas uxorem primogenito suo Her nomine Thamar.
GEN|38|7|Fuit quoque Her primogenitus Iudae nequam in conspectu Domini, et ab eo occisus est.
GEN|38|8|Dixit ergo Iudas ad Onan: " Ingredere ad uxorem fratris tui et sociare illi, ut suscites semen fratri tuo ".
GEN|38|9|Ille, sciens non sibi nasci hunc filium, introiens ad uxorem fratris sui semen fundebat in terram, ne proles fratris nomine nasceretur.
GEN|38|10|Et idcirco occidit et eum Dominus, quod rem detestabilem fecerat.
GEN|38|11|Quam ob rem dixit Iudas Thamar nurui suae: " Esto vidua in domo patris tui, donec crescat Sela filius meus ". Timebat, enim, ne et ipse moreretur sicut fratres eius. Quae abiit et habitavit in domo patris sui.
GEN|38|12|Evolutis autem multis diebus, mortua est filia Sue uxor Iudae. Qui, post luctum consolatione suscepta, ascendebat ad tonsores ovium suarum ipse et Hiras amicus suus Odollamites in Thamnam.
GEN|38|13|Nuntiatumque est Thamar quod socer illius ascenderet in Thamnam ad tondendas oves.
GEN|38|14|Quae, depositis viduitatis vestibus, cooperuit se velo et, mutato habitu, sedit in porta Enaim in via, quae ducit Thamnam; eo quod crevisset Sela, et non eum accepisset maritum.
GEN|38|15|Quam cum vidisset Iudas, suspicatus est esse meretricem; operuerat enim vultum suum.
GEN|38|16|Declinansque ad eam in via ait: " Veni, coeam tecum "; nesciebat enim quod nurus sua esset. Qua respondente: " Quid mihi dabis, ut fruaris concubitu meo? ",
GEN|38|17|dixit: " Mittam tibi haedum de gregibus ". Rursum illa dicente: " Si dederis mihi arrabonem, donec mittas illum ",
GEN|38|18|ait Iudas: " Quid vis tibi pro arrabone dari? ". Respondit: " Sigillum tuum et funiculum et baculum, quem manu tenes ". Et dedit ei. In coitu cum eo mulier concepit
GEN|38|19|et surgens abiit; depositoque velo, induta est viduitatis vestibus.
GEN|38|20|Misit autem Iudas haedum per amicum suum Odollamitem, ut reciperet pignus, quod dederat mulieri. Qui cum non invenisset eam,
GEN|38|21|interrogavit homines loci illius: " Ubi est meretrix, quae sedebat in Enaim in via? ". Respondentibus cunctis: " Non fuit in loco isto meretrix,
GEN|38|22|reversus est ad Iudam et dixit ei: " Non inveni eam; sed et homines loci illius dixerunt mihi numquam ibi sedisse scortum ".
GEN|38|23|Ait Iudas: " Habeat sibi; ne simus in ludibrium. Ego misi haedum, quem promiseram, et tu non invenisti eam ".
GEN|38|24|Ecce autem post tres menses nuntiaverunt Iudae dicentes: " Fornicata est Thamar nurus tua et gravida est ex fornicatione ". Dixitque Iudas: " Producite eam, ut comburatur ".
GEN|38|25|Quae cum educeretur ad poenam, misit ad socerum suum dicens: " De viro, cuius haec sunt, concepi; cognosce cuius sit sigillum et funiculus et baculus ".
GEN|38|26|Qui, agnitis pignoribus, ait: " Iustior me est, quia non tradidi eam Sela filio meo ". Attamen ultra non cognovit illam.
GEN|38|27|Instante autem partu, apparuerunt gemini in utero; atque in ipsa effusione infantium unus protulit manum, in qua obstetrix ligavit coccinum dicens:
GEN|38|28|" Iste egressus est prior ".
GEN|38|29|Illo vero retrahente manum, egressus est frater eius; dixitque mulier: Qualem rupisti tibi rupturam? ". Et ob hanc causam vocatum est nomen eius Phares (id est Ruptura).
GEN|38|30|Postea egressus est frater eius, in cuius manu erat coccinum; qui appellatus est Zara (id est Ortus solis).
GEN|39|1|Igitur Ioseph ductus est in Aegyptum; emitque eum Pu tiphar eunuchus pharaonis, princeps satellitum, vir Aegyptius, de manu Ismaelitarum, a quibus perductus erat.
GEN|39|2|Fuitque Dominus cum eo, et erat vir in cunctis prospere agens habitabatque in domo domini sui.
GEN|39|3|Qui optime noverat esse Dominum cum eo et omnia, quae gereret, ab eo dirigi in manu illius.
GEN|39|4|Invenitque loseph gratiam coram domino suo et ministrabat ei. Et factum est, postquam praeposuit eum domui suae et omnia, quae possidebat, tradidit in manum eius,
GEN|39|5|benedixit Dominus domui Aegyptii propter Ioseph, et benedictio Domini erat in omni possessione eius tam in aedibus quam in agris.
GEN|39|6|Et reliquit omnia, quae possidebat, in manu Ioseph nec cum eo quidquam aliud noverat nisi panem, quo vescebatur. Erat autem Ioseph pulchra facie et decorus aspectu.
GEN|39|7|Post haec ergo iniecit uxor domini eius oculos suos in Ioseph et ait: " Dormi mecum ".
GEN|39|8|Qui nequaquam acquiescens dixit ad eam: " Ecce dominus meus, omnibus mihi traditis, non curat de ulla re in domo sua,
GEN|39|9|nec quisquam maior est in domo hac quam ego, et nihil mihi subtraxit praeter te, quae uxor eius es. Quomodo ergo possum malum hoc magnum facere et peccare in Deum? ".
GEN|39|10|Huiuscemodi verbis per singulos dies et mulier molesta erat adulescenti, et ille recusabat stuprum.
GEN|39|11|Accidit autem quadam die, ut intraret Ioseph domum et opus suum absque arbitris faceret;
GEN|39|12|illa, apprehensa lacinia vestimenti eius, dixit: " Dormi mecum ". Qui, relicto in manu illius pallio, fugit et egressus est foras.
GEN|39|13|Cumque vidisset illum mulier vestem reliquisse in manibus suis et fugisse foras,
GEN|39|14|vocavit homines domus suae et ait ad eos: " En introduxit virum Hebraeum, ut illuderet nobis; ingressus est ad me, ut coiret mecum. Cumque ego succlamassem,
GEN|39|15|et audisset vocem meam, reliquit pallium, quod tenebam, et fugit foras.
GEN|39|16|Retentum pallium ostendit marito revertenti domum
GEN|39|17|et secundum verba haec locuta est: " Ingressus est ad me servus Hebraeus, quem adduxisti, ut illuderet mihi;
GEN|39|18|cumque audisset me clamare, reliquit pallium, quod tenebam, et fugit foras ".
GEN|39|19|Dominus, auditis his verbis coniugis, iratus est valde;
GEN|39|20|tradiditque Ioseph in carcerem, ubi vincti regis custodiebantur. Et erat ibi clausus.
GEN|39|21|Fuit autem Dominus cum Ioseph et misertus illius dedit ei gratiam in conspectu principis carceris.
GEN|39|22|Qui tradidit in manu Ioseph universos vinctos, qui in custodia tenebantur, et, quidquid ibi faciendum erat, ipse faciebat,
GEN|39|23|nec princeps carceris spectabat quidquid in manu eius erat: Dominus enim erat cum illo et omnia opera eius dirigebat.
GEN|40|1|His ita gestis, accidit ut peccarent pincerna regis Aegypti et pistor domino suo.
GEN|40|2|Iratusque pharao contra duos eunuchos, praepositum pincernarum et praepositum pistorum,
GEN|40|3|misit eos in carcerem principis satellitum, in quo erat vinctus et Ioseph.
GEN|40|4|Et princeps satellitum tradidit eos Ioseph, qui ministrabat eis. Aliquantulum temporis illi in custodia tenebantur.
GEN|40|5|Videruntque ambo somnium nocte una iuxta interpretationem congruam sibi.
GEN|40|6|Ad quos cum introisset Ioseph mane et vidisset eos tristes,
GEN|40|7|sciscitatus est eos dicens: " Cur tristior est hodie solito facies vestra? ".
GEN|40|8|Qui responderunt: " Somnium vidimus, et non est qui interpretetur nobis. Dixitque ad eos Ioseph: " Numquid non Dei est interpretatio? Referte mihi quid videritis ".
GEN|40|9|Narravit praepositus pincernarum somnium suum: " Videbam coram me vitem,
GEN|40|10|in qua erant tres propagines, crescere paulatim in gemmas et post flores uvas maturescere;
GEN|40|11|calicemque pharaonis in manu mea. Tuli ergo uvas et expressi in calicem, quem tenebam, et tradidi poculum pharaoni ".
GEN|40|12|Respondit Ioseph: " Haec est interpretatio somnii: tres propagines, tres adhuc dies sunt,
GEN|40|13|post quos elevabit pharao caput tuum et restituet te in gradum pristinum; dabisque ei calicem iuxta officium tuum, sicut facere ante consueveras.
GEN|40|14|Tantum memento mei, cum tibi bene fuerit, et facias mecum misericordiam, ut suggeras pharaoni, ut educat me de isto carcere;
GEN|40|15|quia furto sublatus sum de terra Hebraeorum et hic innocens in lacum missus sum ".
GEN|40|16|Videns pistorum magister quod somnium in bonum dissolvisset, ait: " Et ego vidi somnium, quod tria canistra farinae haberem super caput meum;
GEN|40|17|et in uno canistro, quod erat excelsius, portare me ex omnibus cibis pharaonis, qui fiunt arte pistoria, avesque comedere eos ".
GEN|40|18|Respondit Ioseph: " Haec est interpretatio somnii: tria canistra, tres adhuc dies sunt,
GEN|40|19|post quos auferet pharao caput tuum ac suspendet te in patibulo, et comedent volucres carnes tuas ".
GEN|40|20|Exinde dies tertius natalicius pharaonis erat; qui faciens grande convivium pueris suis elevavit caput magistri pincernarum et caput pistorum principis in medio puerorum suorum;
GEN|40|21|restituitque alterum in locum suum, ut porrigeret ei poculum,
GEN|40|22|alterum suspendit in patibulo, sicut interpretatus erat eis Ioseph.
GEN|40|23|Attamen praepositus pincernarum non est recordatus Ioseph, sed oblitus est interpretis sui.
GEN|41|1|Post duos annos vidit pharao somnium. Putabat se stare super fluvium,
GEN|41|2|de quo ascendebant septem boves pulchrae et crassae et pascebantur in locis palustribus.
GEN|41|3|Aliae quoque septem emergebant post illas de flumine foedae confectaeque macie et stabant in ipsa amnis ripa;
GEN|41|4|devoraveruntque septem boves pulchras et crassas. Expergefactus pharao
GEN|41|5|rursum dormivit et vidit alterum somnium. Septem spicae pullulabant in culmo uno plenae atque formosae.
GEN|41|6|Aliae quoque totidem spicae tenues et percussae vento urente oriebantur
GEN|41|7|devorantes omnem priorum pulchritudinem. Evigilavit pharao, et ecce erat somnium!
GEN|41|8|Et, facto mane, pavore perterritus misit ad omnes coniectores Aegypti cunctosque sapientes suos; et accersitis narravit somnium, nec erat qui interpretaretur.
GEN|41|9|Tunc demum reminiscens pincernarum magister ait: " Confiteor peccatum meum.
GEN|41|10|Iratus rex servis suis me et magistrum pistorum retrudi iussit in carcerem principis satellitum,
GEN|41|11|ubi una nocte uterque vidimus somnium praesagum futurorum.
GEN|41|12|Erat ibi puer Hebraeus eiusdem ducis satellitum famulus, cui narrantes somnia
GEN|41|13|audivimus quidquid postea rei probavit eventus. Ego enim redditus sum officio meo, et ille suspensus est in patibulo ".
GEN|41|14|Protinus ad regis imperium eductum de carcere Ioseph totonderunt ac, veste mutata, obtulerunt ei.
GEN|41|15|Cui ille ait: " Vidi somnia, nec est qui edisserat; quae audivi te sapientissime conicere ".
GEN|41|16|Respondit Ioseph: " Absque me Deus respondebit prospera pharaoni! ".
GEN|41|17|Narravit ergo pharao, quod viderat: " Putabam me stare super ripam fluminis
GEN|41|18|et septem boves de amne conscendere pulchras nimis et obesis carnibus, quae in pastu paludis virecta carpebant.
GEN|41|19|Et ecce has sequebantur aliae septem boves in tantum deformes et macilentae, ut numquam tales in terra Aegypti viderim;
GEN|41|20|quae, devoratis et consumptis prioribus,
GEN|41|21|nullum saturitatis dedere vestigium; sed simili macie et squalore torpebant. Evigilans, rursus sopore depressus,
GEN|41|22|vidi somnium: Septem spicae pullulabant in culmo uno plenae atque pulcherrimae.
GEN|41|23|Aliae quoque septem tenues et percussae vento urente oriebantur e stipula;
GEN|41|24|quae priorum pulchritudinem devoraverunt. Narravi coniectoribus somnium, et nemo est qui edisserat ".
GEN|41|25|Respondit Ioseph: " Somnium regis unum est: quae facturus est, Deus ostendit pharaoni.
GEN|41|26|Septem boves pulchrae et septem spicae plenae septem ubertatis anni sunt; eandemque vim somnii comprehendunt.
GEN|41|27|Septem quoque boves tenues atque macilentae, quae ascenderunt post eas, et septem spicae tenues et vento urente percussae septem anni sunt venturae famis,
GEN|41|28|qui hoc ordine complebuntur:
GEN|41|29|ecce septem anni venient fertilitatis magnae in universa terra Aegypti;
GEN|41|30|quos sequentur septem anni alii tantae sterilitatis, ut oblivioni tradatur cuncta retro abundantia. Consumptura est enim fames omnem terram,
GEN|41|31|et ubertatis magnitudinem perditura est inopiae magnitudo.
GEN|41|32|Quod autem vidisti secundo ad eandem rem pertinens somnium, firmitatis indicium est, eo quod fiat sermo Dei et velocius a Deo impleatur.
GEN|41|33|Nunc ergo provideat rex virum intellegentem et sapientem et praeficiat eum terrae Aegypti
GEN|41|34|constituatque praepositos per cunctas regiones et quintam partem fructuum per septem annos fertilitatis,
GEN|41|35|qui iam nunc futuri sunt, congreget in horrea; et omne frumentum sub pharaonis potestate condatur serveturque in urbibus;
GEN|41|36|et paretur futurae septem annorum fami, quae pressura est Aegyptum, et non consumetur terra inopia ".
GEN|41|37|Placuit pharaoni consilium et cunctis ministris eius.
GEN|41|38|Locutusque est ad eos: " Num invenire poterimus talem virum, qui spiritu Dei plenus sit? ".
GEN|41|39|Dixit ergo ad Ioseph: " Quia ostendit tibi Deus omnia, quae locutus es, numquid sapientiorem et consimilem tui invenire potero?
GEN|41|40|Tu eris super domum meam, et ad tui oris imperium cunctus populus meus oboediet; uno tantum regni solio te praecedam ".
GEN|41|41|Dixitque rursus pharao ad Ioseph: " Ecce, constitui te super universam terram Aegypti ".
GEN|41|42|Tulitque anulum de manu sua et dedit eum in manu eius; vestivitque eum stola byssina et collo torquem auream circumposuit.
GEN|41|43|Fecitque eum ascendere super currum suum secundum, clamante praecone: " Abrech! ", ut omnes coram eo genuflecterent et praepositum esse scirent universae terrae Aegypti.
GEN|41|44|Dixit quoque rex ad Ioseph: " Ego sum pharao; absque tuo imperio non movebit quisquam manum aut pedem in omni terra Aegypti ".
GEN|41|45|Vertitque nomen eius et vocavit eum lingua Aegyptiaca Saphaneth Phanec quod interpretatur Salvator mundi) deditque illi uxorem Aseneth filiam Putiphare sacerdotis Heliopoleos.Egressus est itaque Ioseph ad terram Aegypti
GEN|41|46|­ triginta autem annorum erat quando stetit in conspectu regis pharaonis ­ et circuivit omnes regiones Aegypti.
GEN|41|47|Venitque fertilitas septem annorum, et segetes congregavit in horrea Aegypti
GEN|41|48|condens in singulis urbibus frumentum camporum in circuitu.
GEN|41|49|Tantaque fuit abundantia tritici, ut arenae maris coaequaretur, et copia mensuram excederet.
GEN|41|50|Nati sunt autem Ioseph filii duo, antequam veniret fames, quos ei peperit Aseneth filia Putiphare sacerdotis Heliopoleos.
GEN|41|51|Vocavitque nomen primogeniti Manasses dicens: " Oblivisci me fecit Deus omnium laborum meorum et domus patris mei ".
GEN|41|52|Nomen quoque secundi appellavit Ephraim dicens: " Crescere me fecit Deus in terra paupertatis meae ".
GEN|41|53|Igitur, transactis septem annis ubertatis, qui fuerant in Aegypto,
GEN|41|54|coeperunt venire septem anni inopiae, quos praedixerat Ioseph, et in universo orbe fames praevaluit; in cuncta autem terra Aegypti erat panis.
GEN|41|55|Qua esuriente, clamavit populus ad pharaonem alimenta petens. Quibus ille respondit: " Ite ad Ioseph et, quidquid vobis dixerit, facite ".
GEN|41|56|Et invaluit fames in omni terra Aegypti; aperuitque Ioseph universa horrea et vendebat Aegyptiis; nam et illos oppresserat fames.
GEN|41|57|Omnesque provinciae veniebant in Aegyptum, ut emerent escas apud Ioseph, quia inopia invaluerat in universa terra.
GEN|42|1|Audiens autem Iacob quod alimenta venderentur in Ae gypto, dixit filiis suis: " Quare aspicitis vos invicem?
GEN|42|2|Audivi quod triticum venumdetur in Aegypto; descendite et emite nobis necessaria, ut possimus vivere et non consumamur inopia ".
GEN|42|3|Descenderunt igitur fratres Ioseph decem, ut emerent frumenta in Aegypto,
GEN|42|4|Beniamin fratre Ioseph domi retento a Iacob, qui dixerat fratribus eius: Ne forte in itinere quidquam patiatur mali ".
GEN|42|5|Et ingressi sunt filii Israel terram Aegypti cum aliis, qui pergebant ad emendum. Erat autem fames in terra Chanaan.
GEN|42|6|Et Ioseph erat princeps in terra Aegypti, atque ad eius nutum frumenta populis vendebantur. Cumque venissent et adorassent eum fratres sui proni in terram,
GEN|42|7|et agnovisset eos, quasi ad alienos durius loquebatur interrogans eos: " Unde venistis? ". Qui responderunt: " De terra Chanaan, ut emamus victui necessaria ".
GEN|42|8|Et tamen fratres ipse cognoscens non est cognitus ab eis.
GEN|42|9|Recordatusque somniorum, quae aliquando viderat, ait ad eos: " Exploratores estis; ut videatis infirmiora terrae, venistis! ".
GEN|42|10|Qui dixerunt: " Non est ita, domine; sed servi tui venerunt, ut emerent cibos.
GEN|42|11|Omnes filii unius viri sumus; sinceri sumus, nec quidquam famuli tui machinantur mali ".
GEN|42|12|Quibus ille respondit: " Aliter est; immunita terrae huius considerare venistis! ".
GEN|42|13|At illi: " Duodecim, inquiunt, servi tui fratres sumus filii viri unius in terra Chanaan; minimus cum patre nostro est, alius non est super ".
GEN|42|14|" Hoc est, ait, quod locutus sum: exploratores estis!
GEN|42|15|Iam nunc experimentum vestri capiam: per salutem pharaonis, non egrediemini hinc, donec veniat frater vester minimus!
GEN|42|16|Mittite ex vobis unum, et adducat eum; vos autem eritis in vinculis, donec probentur, quae dixistis, utrum vera an falsa sint. Alioquin, per salutem pharaonis, exploratores estis! ".
GEN|42|17|Tradidit ergo illos custodiae tribus diebus.
GEN|42|18|Die autem tertio eductis de carcere, ait: " Facite, quae dixi, et vivetis; Deum enim timeo.
GEN|42|19|Si sinceri estis, frater vester unus ligetur in carcere; vos autem abite et ferte frumenta, quae emistis, in domos vestras,
GEN|42|20|et fratrem vestrum minimum ad me adducite, ut possim vestros probare sermones, et non moriamini ".Fecerunt, ut dixerat,
GEN|42|21|et locuti sunt ad invicem: " Merito haec patimur, quia peccavimus in fratrem nostrum videntes angustiam animae illius, cum deprecaretur nos, et non audivimus. Idcirco venit super nos ista tribulatio ".
GEN|42|22|Et Ruben ait: " Numquid non dixi vobis: Nolite peccare in puerum? Et non audistis me. En sanguis eius exquiritur ".
GEN|42|23|Nesciebant autem quod intellegeret Ioseph, eo quod per interpretem loquebatur ad eos.
GEN|42|24|Avertitque se parumper et flevit; et reversus locutus est ad eos.
GEN|42|25|Tollensque Simeon et ligans, illis praesentibus, iussit ministris, ut implerent eorum saccos tritico et reponerent pecunias singulorum in sacculis suis, datis supra cibariis in viam. Qui fecerunt ita.
GEN|42|26|At illi portantes frumenta in asinis suis profecti sunt.
GEN|42|27|Apertoque unus sacco, ut daret iumento pabulum in deversorio, contemplatus pecuniam in ore sacculi
GEN|42|28|dixit fratribus suis: " Reddita est mihi pecunia: en habetur in sacco!. Et obstupefacti turbatique mutuo dixerunt: " Quidnam est hoc, quod fecit nobis Deus? ".
GEN|42|29|Veneruntque ad Iacob patrem suum in terram Chanaan; et narraverunt ei omnia, quae accidissent sibi, dicentes:
GEN|42|30|" Locutus est nobis dominus terrae dure et putavit nos exploratores esse provinciae ".
GEN|42|31|Cui respondimus: " Sinceri sumus, nec ullas molimur insidias;
GEN|42|32|duodecim fratres uno patre geniti sumus, unus non est super, minimus cum patre nostro est in terra Chanaan.
GEN|42|33|Et dixit nobis vir, dominus terrae: "Sic probabo quod sinceri sitis: fratrem vestrum unum dimittite apud me et cibaria domibus vestris necessaria sumite et abite;
GEN|42|34|fratremque vestrum minimum adducite ad me, ut sciam quod non sitis exploratores et istum, qui tenetur in vinculis, recipere possitis ac deinceps peragrandi terram habeatis licentiam" ".
GEN|42|35|His dictis, cum frumenta effunderent, singuli reppererunt in ore saccorum ligatas pecunias; exterritisque simul omnibus,
GEN|42|36|dixit pater Iacob: " Absque liberis me esse fecistis: Ioseph non est super, Simeon tenetur in vinculis, et Beniamin auferetis. In me haec omnia mala reciderunt ".
GEN|42|37|Cui respondit Ruben: " Duos filios meos interfice, si non reduxero illum tibi; trade illum in manu mea, et ego eum tibi restituam ".
GEN|42|38|At ille: " Non descendet, inquit, filius meus vobiscum. Frater mortuus est, et ipse solus remansit; si quid ei adversi acciderit in via, deducetis canos meos cum dolore ad inferos ".
GEN|43|1|Interim fames omnem terram vehementer premebat;
GEN|43|2|consumptisque cibis, quos ex Aegypto detulerant, dixit Iacob ad filios suos: " Revertimini et emite nobis pauxillum escarum ".
GEN|43|3|Respondit Iudas: " Denuntiavit nobis vir ille sub attestatione iurisiurandi dicens: "Non videbitis faciem meam, nisi fratrem vestrum minimum adduxeritis vobiscum".
GEN|43|4|Si ergo vis eum mittere nobiscum, pergemus pariter et ememus tibi necessaria;
GEN|43|5|sin autem non vis, non ibimus. Vir enim, ut saepe diximus, denuntiavit nobis dicens: "Non videbitis faciem meam absque fratre vestro minimo" ".
GEN|43|6|Dixit eis Israel: " Cur in meam hoc fecistis miseriam, ut indicaretis ei et alium habere vos fratrem? ".
GEN|43|7|At illi responderunt: " Interrogavit nos homo per ordinem nostram progeniem: si pater viveret, si haberemus fratrem; et nos respondimus ei consequenter iuxta id, quod fuerat sciscitatus. Numquid scire poteramus quod dicturus esset: "Adducite fratrem vestrum vobiscum?" ".
GEN|43|8|Iudas quoque dixit patri suo Israel: " Mitte puerum mecum, ut proficiscamur et possimus vivere, ne moriamur nos et tu et parvuli nostri.
GEN|43|9|Ego spondeo pro puero; de manu mea require illum. Nisi reduxero et reddidero eum tibi, ero peccati reus in te omni tempore.
GEN|43|10|Si non intercessisset dilatio, iam vice altera venissemus ".
GEN|43|11|Igitur Israel pater eorum dixit ad eos: " Si sic necesse est, facite, quod vultis; sumite de optimis terrae fructibus in vasis vestris et deferte viro munera: modicum resinae et mellis et tragacanthum et ladanum, pistacias terebinthi et amygdalas.
GEN|43|12|Pecuniam quoque duplicem ferte vobiscum et illam, quam invenistis in sacculis, reportate, ne forte errore factum sit;
GEN|43|13|sed et fratrem vestrum tollite et ite ad virum.
GEN|43|14|Deus autem meus omnipotens faciat vobis eum placabilem, et remittat vobiscum fratrem vestrum, quem tenet, et hunc Beniamin. Ego autem quasi orbatus absque liberis ero ".
GEN|43|15|Tulerunt ergo viri munera et pecuniam duplicem et Beniamin descenderuntque in Aegyptum; et steterunt coram Ioseph.
GEN|43|16|Quos cum ille vidisset et Beniamin simul, praecepit dispensatori domus suae dicens: " Introduc viros domum et occide victimas et instrue convivium, quoniam mecum sunt comesturi meridie ".
GEN|43|17|Fecit ille, quod sibi fuerat imperatum, et introduxit viros in domum Ioseph.
GEN|43|18|Ibique exterriti dixerunt mutuo: " Propter pecuniam, quam rettulimus prius in saccis nostris, introducti sumus, ut irruant in nos et violenter subiciant servituti et nos et asinos nostros ".
GEN|43|19|Quam ob rem in ipsis foribus accedentes ad dispensatorem domus
GEN|43|20|locuti sunt: " Oramus, domine, ut audias nos. Iam ante descendimus, ut emeremus escas;
GEN|43|21|quibus emptis, cum venissemus ad deversorium, aperuimus saccos nostros et invenimus pecuniam in ore saccorum; quam nunc eodem pondere reportavimus.
GEN|43|22|Sed et aliud attulimus argentum, ut emamus, quae nobis necessaria sunt. Non est in nostra conscientia, quis posuerit argentum in marsupiis nostris.
GEN|43|23|At ille respondit: " Pax vobiscum, nolite timere. Deus vester et Deus patris vestri dedit vobis thesauros in saccis vestris; nam pecuniam, quam dedistis mihi, probatam ego habeo ". Eduxitque ad eos Simeon.
GEN|43|24|Et introductis domum attulit aquam, et laverunt pedes suos; deditque pabulum asinis eorum.
GEN|43|25|Illi vero parabant munera, donec ingrederetur Ioseph meridie; audierant enim quod ibi comesturi essent panem.
GEN|43|26|Igitur ingressus est Ioseph domum suam, obtuleruntque ei munera tenentes in manibus suis; et adoraverunt proni in terram.
GEN|43|27|At ille, clementer resalutatis eis, interrogavit eos dicens: " Salvusne est pater vester senex, de quo dixeratis mihi? Adhuc vivit? ".
GEN|43|28|Qui responderunt: " Sospes est servus tuus pater noster, adhuc vivit ". Et incurvati adoraverunt eum.
GEN|43|29|Attollens autem Ioseph oculos vidit Beniamin fratrem suum uterinum et ait: " Iste est frater vester parvulus, de quo dixeratis mihi? ". Et rursum: " Deus, inquit, misereatur tui, fili mi ".
GEN|43|30|Festinavitque, quia commota fuerant viscera eius super fratre suo, et erumpebant lacrimae; et introiens cubiculum flevit.
GEN|43|31|Rursumque, lota facie, egressus continuit se et ait: " Ponite panes ".
GEN|43|32|Quibus appositis, seorsum Ioseph et seorsum fratribus, Aegyptiis quoque, qui vescebantur simul, seorsum ­ illicitum est enim Aegyptiis comedere cum Hebraeis, et profanum putant huiuscemodi convivium ­
GEN|43|33|sederunt coram eo, primogenitus iuxta primogenita sua et minimus iuxta aetatem suam. Et mirabantur nimis,
GEN|43|34|sumptis partibus, quas ab eo acceperant; maiorque pars venit Beniamin, ita ut quinque partibus excederet. Biberuntque et inebriati sunt cum eo.
GEN|44|1|Praecepit autem Ioseph dispensatori domus suae dicens: " Imple saccos eorum frumento, quantum possunt capere, et pone pecuniam singulorum in summitate sacci.
GEN|44|2|Scyphum autem meum argenteum et pretium, quod dedit tritici, pone in ore sacci iunioris ". Factumque est ita.
GEN|44|3|Et, orto mane, dimissi sunt cum asinis suis.
GEN|44|4|Iamque urbem exierant et processerant paululum, tunc Ioseph, arcessito dispensatore domus: " Surge, inquit, et persequere viros; et apprehensis dicito: "Quare reddidistis malum pro bono? Cur furati estis mihi scyphum argenteum?
GEN|44|5|Nonne ipse est, in quo bibit dominus meus et in quo augurari solet? Pessimam rem fecistis!" ".
GEN|44|6|Fecit ille, ut iusserat, et apprehensis per ordinem locutus est.
GEN|44|7|Qui responderunt: " Quare sic loquitur dominus noster? Absit a servis tuis, ut tantum flagitii commiserimus.
GEN|44|8|Pecuniam, quam invenimus in summitate saccorum, reportavimus ad te de terra Chanaan; et quomodo consequens est, ut furati simus de domo domini tui aurum vel argentum?
GEN|44|9|Apud quemcumque fuerit inventum servorum tuorum, quod quaeris, moriatur; et nos erimus servi domini nostri ".
GEN|44|10|Qui dixit eis: " Fiat iuxta vestram sententiam: apud quemcumque fuerit inventum, ipse sit servus meus; vos autem eritis innoxii ".
GEN|44|11|Itaque festinato deponentes in terram saccos aperuerunt singuli.
GEN|44|12|Quos scrutatus incipiens a maiore usque ad minimum invenit scyphum in sacco Beniamin.
GEN|44|13|At illi, scissis vestibus, oneratisque rursum asinis, reversi sunt in oppidum.
GEN|44|14|Et Iudas cum fratribus ingressus est ad Ioseph ­ necdum enim de loco abierat ­ omnesque ante eum pariter in terram corruerunt.
GEN|44|15|Quibus ille ait: " Cur sic agere voluistis? An ignoratis quod non sit similis mei in augurandi scientia? ".
GEN|44|16|Cui Iudas: " Quid respondebimus, inquit, domino meo? Vel quid loquemur aut iuste poterimus obtendere? Deus invenit iniquitatem servorum tuorum; en omnes servi sumus domini mei, et nos et apud quem inventus est scyphus.
GEN|44|17|Respondit Ioseph: " Absit a me, ut sic agam! Qui furatus est scyphum, ipse sit servus meus; vos autem abite liberi ad patrem vestrum ".
GEN|44|18|Accedens autem propius Iudas confidenter ait: " Oro, domine mi, loquatur servus tuus verbum in auribus tuis, et ne irascaris famulo tuo; tu es enim sicut pharao!
GEN|44|19|Dominus meus interrogavit prius servos suos: "Habetis patrem aut fratrem?".
GEN|44|20|Et nos respondimus domino meo: "Est nobis pater senex et puer parvulus, qui in senectute illius natus est, cuius uterinus frater mortuus est; et ipse solus superest a matre sua, pater vero tenere diligit eum" ".
GEN|44|21|Dixistique servis tuis: "Adducite eum ad me, et ponam oculos meos super illum".
GEN|44|22|Suggessimus domino meo: "Non potest puer relinquere patrem suum; si enim illum dimiserit, morietur".
GEN|44|23|Et dixisti servis tuis: "Nisi venerit frater vester minimus vobiscum, non videbitis amplius faciem meam".
GEN|44|24|Cum ergo ascendissemus ad famulum tuum patrem nostrum, narravimus ei omnia, quae locutus est dominus meus,
GEN|44|25|et dixit pater noster: "Revertimini et emite nobis parum tritici".
GEN|44|26|Cui diximus: "Ire non possumus. Si frater noster minimus descenderit nobiscum, proficiscemur simul; alioquin, illo absente, non poterimus videre faciem viri".
GEN|44|27|Ad quae servus tuus pater meus respondit: "Vos scitis quod duos genuerit mihi uxor mea.
GEN|44|28|Egressus est unus a me, et dixi: Bestia devoravit eum! Et hucusque non comparet.
GEN|44|29|Si tuleritis et istum a facie mea, et aliquid ei in via contigerit, deducetis canos meos cum maerore ad inferos".
GEN|44|30|Igitur, si intravero ad servum tuum patrem meum, et puer defuerit ­ cum anima illius ex huius anima pendeat ­
GEN|44|31|videritque eum non esse nobiscum, morietur; et deducent famuli tui canos eius cum dolore ad inferos.
GEN|44|32|Servus tuus pro puero patri meo spopondit: Nisi reduxero eum, peccati reus ero in patrem meum omni tempore.
GEN|44|33|Manebo itaque servus tuus pro puero in ministerio domini mei, et puer ascendat cum fratribus suis.
GEN|44|34|Non enim possum redire ad patrem meum, absente puero, ne calamitatis, quae oppressura est patrem meum, testis assistam ".
GEN|45|1|Non se poterat ultra cohibere Ioseph omnibus coram astantibus, unde clamavit: " Egredimini, cuncti, foras! ". Et nemo aderat cum eo, quando manifestavit se fratribus suis.
GEN|45|2|Elevavitque vocem cum fletu, quam audierunt Aegyptii omnisque domus pharaonis.
GEN|45|3|Et dixit Ioseph fratribus suis: " Ego sum Ioseph! Adhuc pater meus vivit? ". Nec poterant respondere fratres nimio terrore perterriti.
GEN|45|4|Ad quos ille clementer: " Accedite, inquit, ad me ". Et cum accessissent prope: " Ego sum, ait, Ioseph frater vester, quem vendidistis in Aegyptum.
GEN|45|5|Nolite contristari, neque vobis durum esse videatur quod vendidistis me in his regionibus. Pro salute enim vestra misit me Deus ante vos in Aegyptum.
GEN|45|6|Biennium est enim quod coepit fames esse in terra, et adhuc quinque anni restant, quibus nec arari poterit nec meti.
GEN|45|7|Praemisitque me Deus, ut reservemini super terram, et servetur vita vestra in salvationem magnam.
GEN|45|8|Non vestro consilio, sed Dei voluntate huc missus sum, qui fecit me quasi patrem pharaonis et dominum universae domus eius ac principem in omni terra Aegypti.
GEN|45|9|Festinate et ascendite ad patrem meum et dicetis ei: "Haec mandat filius tuus Ioseph: Deus fecit me dominum universae terrae Aegypti; descende ad me, ne moreris.
GEN|45|10|Et habitabis in terra Gessen; erisque iuxta me tu et filii tui et filii filiorum tuorum, oves tuae et armenta tua et universa, quae possides.
GEN|45|11|Ibique te pascam ­ adhuc enim quinque anni residui sunt famis ­ ne et tu pereas et domus tua et omnia, quae possides".
GEN|45|12|En oculi vestri et oculi fratris mei Beniamin vident quia os meum est, quod loquitur ad vos.
GEN|45|13|Nuntiate patri meo universam gloriam meam in Aegypto et cuncta, quae vidistis. Festinate et adducite eum ad me ".
GEN|45|14|Cumque amplexatus recidisset in collum Beniamin fratris sui, flevit, illo quoque similiter flente, super collum eius.
GEN|45|15|Osculatusque est Ioseph omnes fratres suos et ploravit super singulos. Post quae ausi sunt loqui ad eum.
GEN|45|16|Auditumque est et celebri sermone vulgatum in aula regis: " Venerunt fratres Ioseph! ". Et gavisus est pharao atque omnis familia eius.
GEN|45|17|Dixitque ad Ioseph, ut imperaret fratribus suis dicens: " Onerantes iumenta ite in terram Chanaan
GEN|45|18|et tollite inde patrem vestrum et cognationem et venite ad me; et ego dabo vobis omnia bona Aegypti, ut comedatis medullam terrae.
GEN|45|19|Praecipe etiam: tollite plaustra de terra Aegypti ad subvectionem parvulorum vestrorum ac coniugum et tollite patrem vestrum et properate quantocius venientes.
GEN|45|20|Nec doleatis super supellectilem vestram, quia omnes opes Aegypti vestrae erunt ".
GEN|45|21|Feceruntque filii Israel, ut eis mandatum fuerat. Quibus dedit Ioseph plaustra secundum pharaonis imperium et cibaria in itinere.
GEN|45|22|Singulis quoque proferri iussit vestimentum mutatorium; Beniamin vero dedit trecentos argenteos cum quinque
GEN|45|23|vestimentis mutatoriis. Patri suo misit similiter asinos decem, qui subveherent ex omnibus divitiis Aegypti, et totidem asinas triticum et panem et cibum pro itinere portantes.
GEN|45|24|Dimisit ergo fratres suos et proficiscentibus ait: " Ne irascamini in via! ".
GEN|45|25|Qui ascendentes ex Aegypto venerunt in terram Chanaan ad patrem suum Iacob
GEN|45|26|et nuntiaverunt ei dicentes: " Ioseph vivit et ipse dominatur in omni terra Aegypti! ". At cor eius frigidum mansit; non enim credebat eis.
GEN|45|27|Tunc referebant omnia verba Ioseph, quae dixerat eis. Cumque vidisset plaustra et universa, quae miserat ad adducendum eum, revixit spiritus eius,
GEN|45|28|et ait: " Sufficit mihi, si adhuc Ioseph filius meus vivit. Vadam et videbo illum, antequam moriar ".
GEN|46|1|Profectusque Israel cum omnibus, quae habebat, venit Bersabee et, mactatis ibi victimis Deo patris sui Isaac,
GEN|46|2|audivit eum per visionem noctis vocantem se: " Iacob, Iacob! ". Cui respondit: " Ecce adsum! ".
GEN|46|3|Ait illi: " Ego sum Deus, Deus patris tui. Noli timere descendere in Aegyptum, quia in gentem magnam faciam te ibi.
GEN|46|4|Ego descendam tecum illuc et ego inde adducam te revertentem; Ioseph quoque ponet manus suas super oculos tuos ".
GEN|46|5|Surrexit igitur Iacob a Bersabee, tuleruntque eum filii cum parvulis et uxoribus suis in plaustris, quae miserat pharao ad portandum senem,
GEN|46|6|sumpserunt quoque omnia, quae possederant in terra Chanaan; veneruntque in Aegyptum Iacob et omne semen eius,
GEN|46|7|filii eius et nepotes, filiae et cuncta simul progenies.
GEN|46|8|Haec sunt autem nomina filiorum Israel, qui ingressi sunt in Aegyptum, ipse cum liberis suis.Primogenitus Ruben.
GEN|46|9|Filii Ruben: Henoch et Phallu et Hesron et Charmi.
GEN|46|10|Filii Simeon: Iamuel et Iamin et Ahod et Iachin et Sohar et Saul filius Chananitidis.
GEN|46|11|Filii Levi: Gerson et Caath et Merari.
GEN|46|12|Filii Iudae: Her et Onan et Sela et Phares et Zara. Mortui sunt autem Her et Onan in terra Chanaan. Natique sunt filii Phares: Esrom et Hamul.
GEN|46|13|Filii Issachar: Thola et Phua et Iasub et Semron.
GEN|46|14|Filii Zabulon: Sared et Elon et Iahelel.
GEN|46|15|Hi filii Liae, quos genuit in Paddanaram, cum Dina filia sua. Omnes animae filiorum eius et filiarum triginta tres.
GEN|46|16|Filii Gad: Sephon et Haggi, Suni et Esebon, Heri et Arodi et Areli.
GEN|46|17|Filii Aser: Iemna et lesua et Isui et Beria, Sara quoque soror eorum. Filii Beria: Heber et Melchiel.
GEN|46|18|Hi filii Zelphae, quam dedit Laban Liae filiae suae; et hos genuit Iacob: sedecim animas.
GEN|46|19|Filii Rachel uxoris Iacob: Ioseph et Beniamin.
GEN|46|20|Natique sunt Ioseph filii in terra Aegypti, quos genuit ei Aseneth filia Putiphare sacerdotis Heliopoleos: Manasses et Ephraim.
GEN|46|21|Filii Beniamin: Bela et Bochor et Asbel, Gera et Naaman et Echi et Ros, Mophim et Huphim et Ared.
GEN|46|22|Hi filii Rachel, quos genuit Iacob: omnes animae quattuordecim.
GEN|46|23|Filii Dan: Husim.
GEN|46|24|Filii Nephthali: Iasiel et Guni et Ieser et Sellem.
GEN|46|25|Hi filii Bilhae, quam dedit Laban Racheli filiae suae; et hos genuit Iacob: omnes animae septem.
GEN|46|26|Cunctae animae, quae ingressae sunt cum Iacob in Aegyptum et egressae de femore illius, absque uxoribus filiorum eius, sexaginta sex.
GEN|46|27|Filii autem Ioseph, qui nati sunt ei in terra Aegypti, animae duae. Omnes animae domus Iacob, quae ingressae sunt in Aegyptum, fuere septuaginta.
GEN|46|28|Misit autem Iudam ante se ad Ioseph, ut nuntiaret et occurreret in Gessen.
GEN|46|29|Et venerunt in terram Gessen. Iunctoque Ioseph curru suo, ascendit obviam patri suo in Gessen; vidensque eum irruit super collum eius et inter amplexus diu flevit.
GEN|46|30|Dixitque Israel ad Ioseph: " Iam laetus moriar, quia vidi faciem tuam et superstitem te relinquo ".
GEN|46|31|Et ille locutus est ad fratres suos et ad omnem domum patris sui: " Ascendam et nuntiabo pharaoni dicamque ei: Fratres mei et domus patris mei, qui erant in terra Chanaan, venerunt ad me.
GEN|46|32|Et sunt viri pastores ovium curamque habent alendorum gregum; pecora sua et armenta et omnia, quae habere potuerunt, adduxerunt secum.
GEN|46|33|Cumque vocaverit vos et dixerit: "Quod est opus vestrum?".
GEN|46|34|Respondebitis: "Viri pastores sumus servi tui ab infantia nostra usque in praesens et nos et patres nostri". Haec autem dicetis, ut habitare possitis in terra Gessen, quia detestantur Aegyptii omnes pastores ovium.
GEN|47|1|Ingressus ergo Ioseph nun tiavit pharaoni dicens: " Pater meus et fratres, oves eorum et armenta et cuncta, quae possident, venerunt de terra Chanaan; et ecce consistunt in terra Gessen ".
GEN|47|2|Ex omnibus fratribus suis quinque viros statuit coram rege,
GEN|47|3|quos ille interrogavit: " Quid habetis operis? ". Responderunt: " Pastores ovium sumus servi tui et nos et patres nostri ".
GEN|47|4|Dixeruntque ad pharaonem: " Ad peregrinandum in terra venimus, quoniam non est herba gregibus servorum tuorum, ingravescente fame, in terra Chanaan petimusque, ut esse nos iubeas servos tuos in terra Gessen ".
GEN|47|5|Dixit itaque rex ad Ioseph: " Pater tuus et fratres tui venerunt ad te.
GEN|47|6|Terra Aegypti in conspectu tuo est; in optimo loco fac eos habitare et trade eis terram Gessen. Quod si nosti in eis esse viros industrios, constitue illos magistros pecorum meorum ".
GEN|47|7|Post haec introduxit Ioseph patrem suum ad regem et statuit eum coram eo, qui benedicens illi
GEN|47|8|et interrogatus ab eo: " Quot sunt dies annorum vitae tuae? ",
GEN|47|9|respondit: " Dies peregrinationis meae centum triginta annorum sunt, parvi et mali; et non pervenerunt usque ad dies patrum meorum, quibus peregrinati sunt ".
GEN|47|10|Et benedicto rege, egressus est foras.
GEN|47|11|Ioseph vero patri et fratribus suis dedit possessionem in Aegypto in optimo terrae loco, in terra Ramesses, ut praeceperat pharao;
GEN|47|12|et alebat eos omnemque domum patris sui praebens cibaria singulis.
GEN|47|13|In tota terra panis deerat, et oppresserat fames terram valde, defecitque terra Aegypti et terra Chanaan prae fame.
GEN|47|14|E quibus omnem pecuniam congregavit pro venditione frumenti et intulit eam in aerarium regis.
GEN|47|15|Cumque defecisset emptoribus pretium, venit cuncta Aegyptus ad Ioseph dicens: " Da nobis panes! Quare morimur coram te, deficiente pecunia? ".
GEN|47|16|Quibus ille respondit: " Adducite pecora vestra, et dabo vobis pro eis cibos, si pretium non habetis ".
GEN|47|17|Quae cum adduxissent, dedit eis alimenta pro equis et ovibus et bobus et asinis; sustentavitque eos illo anno pro commutatione pecorum.
GEN|47|18|Venerunt quoque anno secundo et dixerunt ei: " Non celamus dominum nostrum quod, deficiente pecunia, pecora transierunt ad dominum nostrum; nec clam te est quod absque corporibus et terra nihil habeamus.
GEN|47|19|Cur ergo moriemur, te vidente, et nos et terra nostra? Eme nos et terram nostram in servitutem regiam et praebe semina, ne, pereunte cultore, redigatur terra in solitudinem ".
GEN|47|20|Emit igitur Ioseph omnem terram Aegypti, vendentibus singulis possessiones suas prae magnitudine famis. Subiecitque eam pharaoni
GEN|47|21|et cunctos populos eius redegit ei in servitutem, a novissimis terminis Aegypti usque ad extremos fines eius.
GEN|47|22|Terram autem sacerdotum non emit, qui cibariis a rege statutis fruebantur, et idcirco non sunt compulsi vendere possessiones suas.
GEN|47|23|Dixit ergo Ioseph ad populos: " En, ut cernitis, et vos et terram vestram pharao possidet; accipite semina et serite agros,
GEN|47|24|ut fruges habere possitis. Quintam partem regi dabitis; quattuor reliquas permitto vobis in sementem et in cibum familiis et liberis vestris ".
GEN|47|25|Qui responderunt: " Tu salvasti nos! Respiciat nos tantum dominus noster, et laeti serviemus regi ".
GEN|47|26|Ex eo tempore usque in praesentem diem in universa terra Aegypti regibus quinta pars solvitur; et factum est a Ioseph in legem absque terra sacerdotali, quae libera ab hac condicione est.
GEN|47|27|Habitavit ergo Israel in Aegypto, id est in terra Gessen, et possedit eam; auctusque est et multiplicatus nimis.
GEN|47|28|Et vixit Iacob in terra Aegypti decem et septem annis; factique sunt omnes dies vitae illius centum quadraginta septem annorum.
GEN|47|29|Cumque appropinquare cerneret diem mortis suae, vocavit filium suum Ioseph et dixit ad eum: " Si inveni gratiam in conspectu tuo, pone manum tuam sub femore meo et facies mihi misericordiam et veritatem, ut non sepelias me in Aegypto,
GEN|47|30|sed dormiam cum patribus meis, et auferas me de terra hac condasque in sepulcro maiorum meorum ". Cui respondit Ioseph: " Ego faciam, quod iussisti ".
GEN|47|31|Et ille: " Iura ergo, inquit, mihi! ". Quo iurante, adoravit Israel conversus ad lectuli caput.
GEN|48|1|His ita transactis, nuntiatum est Ioseph quod aegrotaret pater suus. Et assumpsit secum duos filios Manasse et Ephraim.
GEN|48|2|Dictumque est seni: " Ecce filius tuus Ioseph venit ad te ". Qui confortatus sedit in lectulo
GEN|48|3|et ingresso ad se ait: " Deus omnipotens apparuit mihi in Luza, quae est in terra Chanaan, benedixitque mihi
GEN|48|4|et ait: "Ego te augebo et multiplicabo et faciam te in multitudinem populorum; daboque tibi terram hanc et semini tuo post te in possessionem sempiternam".
GEN|48|5|Duo ergo filii tui, qui nati sunt tibi in terra Aegypti, antequam huc venirem ad te, mei erunt: Ephraim et Manasses sicut Ruben et Simeon reputabuntur mihi.
GEN|48|6|Reliquos autem, quos genueris post eos, tui erunt et nomine fratrum suorum vocabuntur in possessionibus suis.
GEN|48|7|Mihi enim, quando veniebam de Paddanaram, mortua est Rachel mater tua in terra Chanaan in ipso itinere, cum adhuc esset spatium aliquod usque ad Ephratham, et sepelivi eam iuxta viam Ephrathae, quae alio nomine appellatur Bethlehem ".
GEN|48|8|Videns autem filios eius dixit ad eum: " Qui sunt isti? ".
GEN|48|9|Respondit: " Filii mei sunt, quos donavit mihi Deus in hoc loco ". " Adduc, inquit, eos ad me, ut benedicam illis! ".
GEN|48|10|Oculi enim Israel caligabant prae nimia senectute, et clare videre non poterat. Applicitosque ad se deosculatus et circumplexus eos
GEN|48|11|dixit ad filium suum: " Non sum fraudatus aspectu tuo; insuper ostendit mihi Deus semen tuum ".
GEN|48|12|Cumque tulisset eos Ioseph de gremio patris, adoravit pronus in terram.
GEN|48|13|Et posuit Ephraim ad dexteram suam, id est ad sinistram Israel, Manassen vero in sinistra sua, ad dexteram scilicet patris; applicuitque ambos ad eum.
GEN|48|14|Qui extendens manum dexteram, posuit super caput Ephraim minoris fratris, sinistram autem super caput Manasse, qui maior natu erat, commutans manus.
GEN|48|15|Benedixitque Iacob Ioseph et ait: Deus, in cuius conspectu ambulaveruntpatres mei Abraham et Isaac,Deus, qui pascit me ab adulescentia meausque in praesentem diem,
GEN|48|16|Angelus, qui eruit me de cunctis malis,benedicat pueris istis!Et invocetur super eos nomen meum,nomina quoque patrum meorum Abraham et Isaac,et crescant in multitudinemsuper terram! ".
GEN|48|17|Videns autem Ioseph quod posuisset pater suus dexteram manum super caput Ephraim, graviter accepit et apprehensam manum patris levare conatus est de capite Ephraim et transferre super caput Manasse.
GEN|48|18|Dixitque ad patrem: " Non ita convenit, pater, quia hic est primogenitus; pone dexteram tuam super caput eius! ".
GEN|48|19|Qui renuens ait: " Scio, fili mi, scio; et iste quidem erit in populos et multiplicabitur, sed frater eius minor maior erit illo, et semen illius crescet in plenitudinem gentium ".
GEN|48|20|Benedixitque eis in die illo dicens: In te benedicet Israel atque dicet: "Faciat te Deus sicut Ephraim et sicut Manasse!" ".Constituitque Ephraim ante Manassen.
GEN|48|21|Et ait ad Ioseph filium suum: " En ego morior, et erit Deus vobiscum reducetque vos ad terram patrum vestrorum.
GEN|48|22|Do tibi partem unam extra fratres tuos, quam tuli de manu Amorraei in gladio et arcu meo ".
GEN|49|1|Vocavit autem Iacob filios suos et ait eis: " Congrega mini, ut annuntiem, quae ventura sunt vobis in diebus novissimis.
GEN|49|2|Congregamini et audite, filii Iacob,audite Israel patrem vestrum!
GEN|49|3|Ruben primogenitus meus,tu fortitudo mea et principium roboris mei;prior in dignitate, maior in robore!
GEN|49|4|Ebulliens sicut aqua non excellas,quia ascendisti cubile patris tuiet maculasti stratum meum.
GEN|49|5|Simeon et Levi fratres,vasa violentiae arma eorum.
GEN|49|6|In consilium eorum ne veniat anima mea,et in coetu illorum non sit gloria mea;quia in furore suo occiderunt virumet in voluntate sua subnervaverunt tauros.
GEN|49|7|Maledictus furor eorum, quia pertinax,et indignatio eorum, quia dura!Dividam eos in Iacobet dispergam eos in Israel.
GEN|49|8|Iuda, te laudabunt fratres tui;manus tua in cervicibus inimicorum tuorum;adorabunt te filii patris tui.
GEN|49|9|Catulus leonis Iuda:a praeda, fili mi, ascendisti;requiescens accubuit ut leoet quasi leaena; quis suscitabit eum?
GEN|49|10|Non auferetur sceptrum de Iudaet baculus ducis de pedibus eius,donec veniat ille, cuius est,et cui erit oboedientia gentium;
GEN|49|11|ligans ad vineam pullum suumet ad vitem filium asinae suae,lavabit in vino stolam suamet in sanguine uvae pallium suum;
GEN|49|12|nigriores sunt oculi eius vinoet dentes eius lacte candidiores.
GEN|49|13|Zabulon in litore maris habitabitet in statione navium,pertingens usque ad Sidonem.
GEN|49|14|Issachar asinus fortis,accubans inter caulas
GEN|49|15|vidit requiem quod esset bona,et terram quod optima;et supposuit umerum suum ad portandumfactusque est tributis serviens.
GEN|49|16|Dan iudicabit populum suumsicut una tribuum Israel.
GEN|49|17|Fiat Dan coluber in via,cerastes in semita,mordens calcanea equi,ut cadat ascensor eius retro.
GEN|49|18|Salutare tuum exspectabo, Domine!
GEN|49|19|Gad, latrones aggredientur eum,ipse autem aggredietur calcaneum eorum.
GEN|49|20|Aser, pinguis panis eius,et praebebit delicias regales.
GEN|49|21|Nephthali cerva emissa,dans cornua pulchra.
GEN|49|22|Arbor fructifera Ioseph,arbor fructifera super fontem:rami transcendunt murum.
GEN|49|23|Sed exasperaverunt eum et iurgati sunt,et adversati sunt illi habentes iacula.
GEN|49|24|Et confractus est arcus eorum,et dissoluti sunt nervi brachiorum eorumper manus Potentis Iacob,per nomen Pastoris, Lapidis Israel.
GEN|49|25|Deus patris tui erit adiutor tuus,et Omnipotens benedicet tibibenedictionibus caeli desuper,benedictionibus abyssi iacentisdeorsum,benedictionibus uberum et vulvae.
GEN|49|26|Benedictiones patris tui confortatae suntsuper benedictiones montium aeternorum,desiderium collium antiquorum;fiant in capite Iosephet in vertice nazaraei inter fratres suos.
GEN|49|27|Beniamin lupus rapax;mane comedet praedamet vespere dividet spolia ".
GEN|49|28|Omnes hi in tribubus Israel duodecim. Haec locutus est eis pater suus benedixitque singulis benedictionibus propriis.
GEN|49|29|Et praecepit eis dicens: " Ego congregor ad populum meum; sepelite me cum patribus meis in spelunca Machpela, quae est in agro Ephron Hetthaei
GEN|49|30|contra Mambre in terra Chanaan, quam emit Abraham cum agro ab Ephron Hetthaeo in possessionem sepulcri;
GEN|49|31|ibi sepelierunt eum et Saram uxorem eius, ibi sepultus est Isaac cum Rebecca coniuge sua, ibi et Lia condita iacet ".
GEN|49|32|Finitisque mandatis, quibus filios instruebat, collegit pedes suos super lectulum et obiit; appositusque est ad populum suum.
GEN|50|1|Ioseph ruit super faciem patris flens et deosculans eum.
GEN|50|2|Praecepitque servis suis medicis, ut aromatibus condirent patrem.
GEN|50|3|Quibus iussa explentibus, transierunt quadraginta dies; iste quippe mos erat cadaverum conditorum. Flevitque eum Aegyptus septuaginta diebus.
GEN|50|4|Et, expleto planctus tempore, locutus est Ioseph ad familiam pharaonis: Si inveni gratiam in conspectu vestro, loquimini in auribus pharaonis,
GEN|50|5|eo quod pater meus adiuraverit me dicens: "En morior; in sepulcro meo, quod fodi mihi in terra Chanaan, sepelies me"; ascendam nunc et sepeliam patrem meum ac revertar ".
GEN|50|6|Dixitque ei pharao: " Ascende et sepeli patrem tuum, sicut adiuratus es.
GEN|50|7|Quo ascendente, ierunt cum eo omnes servi pharaonis, senes domus eius cunctique maiores natu terrae Aegypti,
GEN|50|8|domus Ioseph cum fratribus suis, absque parvulis et gregibus atque armentis, quae dereliquerant in terra Gessen.
GEN|50|9|Habuit quoque in comitatu currus et equites; et facta est turba non modica.
GEN|50|10|Veneruntque ad Gorenatad (id est Aream rhamni), quae sita est trans Iordanem; ubi celebrantes exsequias planctu magno atque vehementi impleverunt septem dies.
GEN|50|11|Quod cum vidissent habitatores terrae Chanaan, dixerunt: " Planctus magnus est iste Aegyptiis "; et idcirco vocatum est nomen loci illius Abelmesraim (id est Planctus Aegypti).
GEN|50|12|Fecerunt ergo filii Iacob, sicut praeceperat eis;
GEN|50|13|et portantes eum in terram Chanaan sepelierunt eum in spelunca Machpela, quam emerat Abraham cum agro in possessionem sepulcri ab Ephron Hetthaeo contra faciem Mambre.
GEN|50|14|Reversusque est Ioseph in Aegyptum cum fratribus suis et omni comitatu, sepulto patre.
GEN|50|15|Quo mortuo, timentes fratres eius et mutuo colloquentes: " Ne forte memor sit iniuriae, quam passus est, et reddat nobis omne malum, quod fecimus ",
GEN|50|16|mandaverunt ei dicentes: " Pater tuus praecepit nobis, antequam moreretur,
GEN|50|17|ut haec tibi verbis illius diceremus: "Obsecro, ut obliviscaris sceleris fratrum tuorum et peccati atque malitiae, quam exercuerunt in te". Nos quoque oramus, ut servis Dei patris tui dimittas iniquitatem hanc. Quibus auditis, flevit Ioseph.
GEN|50|18|Veneruntque ad eum fratres sui et proni coram eo dixerunt: " Servi tui sumus ".
GEN|50|19|Quibus ille respondit: " Nolite timere. Num Dei possumus resistere voluntati?
GEN|50|20|Vos cogitastis de me malum; sed Deus vertit illud in bonum, ut exaltaret me, sicut in praesentiarum cernitis, et salvos faceret multos populos.
GEN|50|21|Nolite timere: ego pascam vos et parvulos vestros ". Consolatusque est eos et blande ac leniter est locutus.
GEN|50|22|Et habitavit in Aegypto cum omni domo patris sui; vixitque centum decem annis
GEN|50|23|et vidit Ephraim filios usque ad tertiam generationem; filii quoque Machir filii Manasse nati sunt in genibus Ioseph.
GEN|50|24|Quibus transactis, locutus est fratribus suis: " Post mortem meam Deus visitabit vos et ascendere vos faciet de terra ista ad terram, quam iuravit Abraham, Isaac et Iacob ".
GEN|50|25|Cumque adiurasset eos atque dixisset: " Deus visitabit vos; asportate ossa mea vobiscum de loco isto ",
GEN|50|26|mortuus est, expletis centum decem vitae suae annis. Et conditus aromatibus repositus est in loculo in Aegypto.
EXOD|1|1|Haec sunt nomina filiorum Is rael, qui ingressi sunt Aegyp tum cum Iacob; singuli cum domibus suis introierunt:
EXOD|1|2|Ruben, Simeon, Levi, Iuda,
EXOD|1|3|Issachar, Zabulon et Beniamin,
EXOD|1|4|Dan et Nephthali, Gad et Aser.
EXOD|1|5|Erant igitur omnes animae eorum, qui egressi sunt de femore Iacob, septuaginta; Ioseph autem in Aegypto erat.
EXOD|1|6|Quo mortuo et universis fratribus eius omnique cognatione illa,
EXOD|1|7|filii Israel creverunt et pullulantes multiplicati sunt ac roborati nimis impleverunt terram.
EXOD|1|8|Surrexit interea rex novus super Aegyptum, qui ignorabat Ioseph;
EXOD|1|9|et ait ad populum suum: " Ecce, populus filiorum Israel multus et fortior nobis est;
EXOD|1|10|venite, prudenter agamus cum eo, ne forte multiplicetur et, si ingruerit contra nos bellum, addatur inimicis nostris, expugnatisque nobis, egrediatur de terra ".
EXOD|1|11|Praeposuit itaque eis magistros operum, ut affligerent eos oneribus; aedificaveruntque urbes promptuarias pharaoni, Phithom et Ramesses.
EXOD|1|12|Quantoque opprimebant eos, tanto magis multiplicabantur et crescebant.
EXOD|1|13|Formidaveruntque filios Israel Aegyptii et in servitutem redegerunt eos
EXOD|1|14|atque ad amaritudinem perducebant vitam eorum operibus duris luti et lateris omnique famulatu, quo in terrae operibus premebantur.
EXOD|1|15|Dixit autem rex Aegypti obstetricibus Hebraeorum, quarum una vocabatur Sephra, altera Phua,
EXOD|1|16|praecipiens eis: " Quando obstetricabitis Hebraeas, et partus tempus advenerit, si masculus fuerit, interficite eum; si femina, reservate ".
EXOD|1|17|Timuerunt autem obstetrices Deum et non fecerunt iuxta praeceptum regis Aegypti, sed conservabant mares.
EXOD|1|18|Quibus ad se accersitis rex ait: " Quidnam est hoc, quod facere voluistis, ut pueros servaretis? ".
EXOD|1|19|Quae responderunt: " Non sunt Hebraeae sicut Aegyptiae mulieres; ipsae enim robustae sunt et, priusquam veniamus ad eas, pariunt ".
EXOD|1|20|Bene ergo fecit Deus obstetricibus, et crevit populus confortatusque est nimis;
EXOD|1|21|et, quia timuerunt obstetrices Deum, aedificavit illis domos.
EXOD|1|22|Praecepit ergo pharao omni populo suo dicens: " Quidquid masculini sexus natum fuerit, in flumen proicite; quidquid feminei, reservate ".
EXOD|2|1|Egressus est vir de domo Levi et accepit uxorem stirpis suae;
EXOD|2|2|quae concepit et peperit filium et videns eum elegantem abscondit tribus mensibus.
EXOD|2|3|Cumque iam celare non posset, sumpsit fiscellam scirpeam et linivit eam bitumine ac pice; posuitque intus infantulum et exposuit eum in carecto ripae fluminis,
EXOD|2|4|stante procul sorore eius et considerante eventum rei.
EXOD|2|5|Ecce autem descendebat filia pharaonis, ut lavaretur in flumine, et puellae eius gradiebantur per crepidinem alvei. Quae cum vidisset fiscellam in papyrione, misit unam e famulabus suis; et allatam
EXOD|2|6|aperiens cernensque in ea parvulum vagientem, miserta eius ait: " De infantibus Hebraeorum est hic ".
EXOD|2|7|Cui soror pueri: " Vis, inquit, ut vadam et vocem tibi mulierem Hebraeam, quae nutrire possit tibi infantulum? ".
EXOD|2|8|Respondit: " Vade ". Perrexit puella et vocavit matrem infantis.
EXOD|2|9|Ad quam locuta filia pharaonis: " Accipe, ait, puerum istum et nutri mihi; ego dabo tibi mercedem tuam ". Suscepit mulier et nutrivit puerum adultumque tradidit filiae pharaonis.
EXOD|2|10|Quem illa adoptavit in locum filii vocavitque nomen eius Moysen dicens: " Quia de aqua tuli eum ".
EXOD|2|11|In diebus illis, postquam creverat, Moyses egressus est ad fratres suos; viditque afflictionem eorum et virum Aegyptium percutientem quendam de Hebraeis fratribus suis.
EXOD|2|12|Cumque circumspexisset huc atque illuc et nullum adesse vidisset, percussum Aegyptium abscondit sabulo.
EXOD|2|13|Et egressus die altero conspexit duos Hebraeos rixantes dixitque ei, qui faciebat iniuriam: " Quare percutis proximum tuum? ".
EXOD|2|14|Qui respondit: " Quis te constituit principem et iudicem super nos? Num occidere me tu vis, sicut occidisti Aegyptium? ". Timuit Moyses et ait: " Quomodo palam factum est verbum istud? ".
EXOD|2|15|Audivitque pharao sermonem hunc et quaerebat occidere Moysen. Qui fugiens de conspectu eius moratus est in terra Madian; venit ergo in terram Madian et sedit iuxta puteum.
EXOD|2|16|Erant autem sacerdoti Madian septem filiae, quae venerunt ad hauriendam aquam; et impletis canalibus adaquare cupiebant greges patris sui.
EXOD|2|17|Supervenere pastores et eiecerunt eas: surrexitque Moyses et, defensis puellis, adaquavit oves earum.
EXOD|2|18|Quae cum revertissent ad Raguel patrem suum, dixit ad eas: " Cur velocius venistis solito? ".
EXOD|2|19|Responderunt: " Vir Aegyptius liberavit nos de manu pastorum; insuper et hausit aquam nobis potumque dedit ovibus ".
EXOD|2|20|At ille: " Ubi est? ", inquit. " Quare dimisistis hominem? Vocate eum, ut comedat panem ".
EXOD|2|21|Consensit ergo Moyses habitare cum eo accepitque Sephoram filiam eius uxorem.
EXOD|2|22|Quae peperit ei filium, quem vocavit Gersam dicens: " Advena sum in terra aliena ".
EXOD|2|23|Post multum vero temporis mortuus est rex Aegypti; et ingemiscentes filii Israel propter opera vociferati sunt, ascenditque clamor eorum ad Deum ab operibus.
EXOD|2|24|Et audivit gemitum eorum ac recordatus est foederis, quod pepigit cum Abraham, Isaac et Iacob;
EXOD|2|25|et respexit Dominus filios Israel et apparuit eis.
EXOD|3|1|Moyses autem pascebat oves Iethro soceri sui sacerdotis Ma dian; cumque minasset gregem ultra desertum, venit ad montem Dei Horeb.
EXOD|3|2|Apparuitque ei angelus Domini in flamma ignis de medio rubi; et videbat quod rubus arderet et non combureretur.
EXOD|3|3|Dixit ergo Moyses: " Vadam et videbo visionem hanc magnam, quare non comburatur rubus ".
EXOD|3|4|Cernens autem Dominus quod pergeret ad videndum, vocavit eum Deus de medio rubi et ait: " Moyses, Moyses ". Qui respondit: " Adsum ".
EXOD|3|5|At ille: " Ne appropies, inquit, huc; solve calceamentum de pedibus tuis; locus enim, in quo stas, terra sancta est ".
EXOD|3|6|Et ait: " Ego sum Deus patris tui, Deus Abraham, Deus Isaac et Deus Iacob ". Abscondit Moyses faciem suam; non enim audebat aspicere contra Deum.
EXOD|3|7|Cui ait Dominus: " Vidi afflictionem populi mei in Aegypto et clamorem eius audivi propter duritiam exactorum eorum.
EXOD|3|8|Et sciens dolorem eius descendi, ut liberem eum de manibus Aegyptiorum et educam de terra illa in terram bonam et spatiosam, in terram, quae fluit lacte et melle, ad loca Chananaei et Hetthaei et Amorraei et Pherezaei et Hevaei et Iebusaei.
EXOD|3|9|Clamor ergo filiorum Israel venit ad me, vidique afflictionem eorum, qua ab Aegyptiis opprimuntur;
EXOD|3|10|sed veni, mittam te ad pharaonem, ut educas populum meum, filios Israel, de Aegypto ".
EXOD|3|11|Dixitque Moyses ad Deum: " Quis sum ego, ut vadam ad pharaonem et educam filios Israel de Aegypto? ".
EXOD|3|12|Qui dixit ei: " Ego ero tecum; et hoc habebis signum quod miserim te: cum eduxeris populum de Aegypto, servietis Deo super montem istum ".
EXOD|3|13|Ait Moyses ad Deum: " Ecce, ego vadam ad filios Israel et dicam eis: Deus patrum vestrorum misit me ad vos. Si dixerint mihi: "Quod est nomen eius?" quid dicam eis? ".
EXOD|3|14|Dixit Deus ad Moysen: " Ego sum qui sum ". Ait: " Sic dices filiis Israel: Qui sum misit me ad vos ".
EXOD|3|15|Dixitque iterum Deus ad Moysen: " Haec dices filiis Israel: Dominus, Deus patrum vestrorum, Deus Abraham, Deus Isaac et Deus lacob, misit me ad vos; hoc nomen mihi est in aeternum, et hoc memoriale meum in generationem et generationem.
EXOD|3|16|Vade et congrega seniores Israel et dices ad eos: Dominus, Deus patrum vestrorum, apparuit mihi, Deus Abraham, Deus Isaac et Deus Iacob, dicens: Visitans visitavi vos et vidi omnia, quae acciderunt vobis in Aegypto;
EXOD|3|17|et dixi: Educam vos de afflictione Aegypti in terram Chananaei et Hetthaei et Amorraei et Pherezaei et Hevaei et Iebusaei, ad terram fluentem lacte et melle.
EXOD|3|18|Et audient vocem tuam; ingredierisque tu et seniores Israel ad regem Aegypti, et dicetis ad eum: Dominus, Deus Hebraeorum, occurrit nobis; et nunc eamus viam trium dierum in solitudinem, ut immolemus Domino Deo nostro.
EXOD|3|19|Sed ego scio quod non dimittet vos rex Aegypti, ut eatis, nisi per manum validam.
EXOD|3|20|Extendam enim manum meam et percutiam Aegyptum in cunctis mirabilibus meis, quae facturus sum in medio eius; post haec dimittet vos.
EXOD|3|21|Daboque gratiam populo huic coram Aegyptiis, et, cum egrediemini, non exibitis vacui.
EXOD|3|22|Sed postulabit mulier a vicina sua et ab hospita sua vasa argentea et aurea ac vestes; ponetisque eas super filios et filias vestras et spoliabitis Aegyptum ".
EXOD|4|1|Respondens Moyses ait: " Quid autem, si non credent mihi ne que audient vocem meam, sed dicent: "Non apparuit tibi Dominus?" ".
EXOD|4|2|Dixit ergo ad eum: " Quid est quod tenes in manu tua? ". Respondit: " Virga ".
EXOD|4|3|Dixitque Dominus: " Proice eam in terram! ". Proiecit, et versa est in serpentem, ita ut fugeret Moyses.
EXOD|4|4|Dixitque Dominus: " Extende manum tuam et apprehende caudam eius! ". Extendit et tenuit, versaque est in virgam.
EXOD|4|5|" Ut credant, inquit, quod apparuerit tibi Dominus, Deus patrum suorum, Deus Abraham, Deus Isaac et Deus Iacob ".
EXOD|4|6|Dixitque Dominus rursum: " Mitte manum tuam in sinum tuum! ". Quam cum misisset in sinum, protulit leprosam instar nivis.
EXOD|4|7|" Retrahe, ait, manum tuam in sinum tuum! ". Retraxit et protulit iterum, et erat similis carni reliquae.
EXOD|4|8|" Si non crediderint, inquit, tibi, neque audierint sermonem signi prioris, credent verbo signi sequentis.
EXOD|4|9|Quod si nec duobus quidem his signis crediderint neque audierint vocem tuam, sume aquam fluminis et effunde eam super aridam, et, quidquid hauseris de fluvio, vertetur in sanguinem ".
EXOD|4|10|Ait Moyses: " Obsecro, Domine, non sum eloquens ab heri et nudiustertius et ex quo locutus es ad servum tuum, nam impeditioris et tardioris linguae sum ".
EXOD|4|11|Dixit Dominus ad eum: " Quis fecit os hominis? Aut quis fabricatus est mutum vel surdum vel videntem vel caecum? Nonne ego?
EXOD|4|12|Perge igitur, et ego ero in ore tuo; doceboque te quid loquaris ".
EXOD|4|13|At ille: " Obsecro, inquit, Domine, mitte quem missurus es ".
EXOD|4|14|Iratus Dominus in Moysen ait: " Aaron, frater tuus Levites, scio quod eloquens sit; ecce ipse egreditur in occursum tuum vidensque te laetabitur corde.
EXOD|4|15|Loquere ad eum et pone verba mea in ore eius; et ego ero in ore tuo et in ore illius et ostendam vobis quid agere debeatis.
EXOD|4|16|Ipse loquetur pro te ad populum et erit os tuum; tu autem eris ei ut Deus.
EXOD|4|17|Virgam quoque hanc sume in manu tua, in qua facturus es signa ".
EXOD|4|18|Abiit Moyses et reversus est ad Iethro socerum suum dixitque ei: " Vadam, quaeso, et revertar ad fratres meos in Aegyptum, ut videam, si adhuc vivant ". Cui ait Iethro: " Vade in pace ".
EXOD|4|19|Dixit ergo Dominus ad Moysen in Madian: " Vade, revertere in Aegyptum; mortui sunt enim omnes, qui quaerebant animam tuam ".
EXOD|4|20|Tulit Moyses uxorem suam et filios suos et imposuit eos super asinum; reversusque est in Aegyptum portans virgam Dei in manu sua.
EXOD|4|21|Dixitque ei Dominus revertenti in Aegyptum: " Vide, ut omnia ostenta, quae posui in manu tua, facias coram pharaone; ego indurabo cor eius, et non dimittet populum.
EXOD|4|22|Dicesque ad eum: Haec dicit Dominus: Filius meus primogenitus Israel.
EXOD|4|23|Dico tibi: Dimitte filium meum, ut serviat mihi; si autem non vis dimittere eum, ecce ego interficiam filium tuum primogenitum ".
EXOD|4|24|Cumque esset in itinere, in deversorio, occurrit ei Dominus et volebat occidere eum.
EXOD|4|25|Tulit ilico Sephora acutissimam petram et circumcidit praeputium filii sui; tetigitque pedes eius et ait: " Sponsus sanguinum tu mihi es ".
EXOD|4|26|Et dimisit eum, postquam dixerat: " Sponsus sanguinum ", ob circumcisionem.
EXOD|4|27|Dixit autem Dominus ad Aaron: " Vade in occursum Moysi in desertum ". Qui perrexit obviam ei in montem Dei et osculatus est eum.
EXOD|4|28|Narravitque Moyses Aaron omnia verba Domini, quibus miserat eum, et signa, quae mandaverat.
EXOD|4|29|Veneruntque simul et congregaverunt cunctos seniores filiorum Israel.
EXOD|4|30|Locutusque est Aaron omnia verba, quae dixerat Dominus ad Moysen, et fecit signa coram populo.
EXOD|4|31|Et credidit populus, audieruntque quod visitasset Dominus filios Israel et quod respexisset afflictionem eorum; et proni adoraverunt.
EXOD|5|1|Post haec ingressi sunt Moyses et Aaron et dixerunt pharaoni: " Haec dicit Dominus, Deus Israel: Dimitte populum meum, ut sacrificet mihi in deserto ".
EXOD|5|2|At ille responclit: " Quis est Dominus, ut audiam vocem eius et dimittam Israel? Nescio Dominum et Israel non dimittam ".
EXOD|5|3|Dixeruntque: " Deus Hebraeorum occurrit nobis; eamus, quaeso, viam trium dierum in solitudinem et sacrificemus Domino Deo nostro, ne forte accidat nobis pestis aut gladius ".
EXOD|5|4|Ait ad eos rex Aegypti: " Quare, Moyses et Aaron, sollicitatis populum ab operibus suis? Ite ad onera vestra ".
EXOD|5|5|Dixitque pharao: " Multus nimis iam est populus terrae; videtis quod turba succreverit; quanto magis si dederitis eis requiem ab operibus? ".
EXOD|5|6|Praecepit ergo in die illo exactoribus populi et praefectis eius dicens:
EXOD|5|7|" Nequaquam ultra dabitis paleas populo ad conficiendos lateres sicut prius, sed ipsi vadant et colligant stipulas.
EXOD|5|8|Et mensuram laterum, quam prius faciebant, imponetis super eos; nec minuetis quidquam. Vacant enim et idcirco vociferantur dicentes: "Eamus et sacrificemus Deo nostro".
EXOD|5|9|Opprimantur operibus et expleant ea, ut non acquiescant verbis mendacibus ".
EXOD|5|10|Igitur egressi exactores populi et praefecti eius dixerunt ad populum: " Sic dicit pharao: "Non do vobis paleas.
EXOD|5|11|Ite et colligite, sicubi invenire poteritis, nec minuetur quid quam de opere vestro" ".
EXOD|5|12|Dispersusque est populus per omnem terram Aegypti ad colligendas paleas.
EXOD|5|13|Exactores quoque instabant dicentes: " Complete opus vestrum cotidie, ut prius facere solebatis, quando dabantur vobis paleae ".
EXOD|5|14|Flagellatique sunt praefecti filiorum Israel, quos constituerant super eos exactores pharaonis dicentes: " Quare non implestis mensuram laterum sicut prius, nec heri nec hodie? ".
EXOD|5|15|Veneruntque praefecti filiorum Israel et vociferati sunt ad pharaonem dicentes: " Cur ita agis contra servos tuos?
EXOD|5|16|Paleae non dantur nobis, et lateres similiter imperantur; en famuli tui flagellis caedimur, et populus tuus est in culpa ".
EXOD|5|17|Qui ait: " Vacatis otio et idcirco dicitis: "Eamus et sacrificemus Domino".
EXOD|5|18|Ite ergo et operamini; paleae non dabuntur vobis, et reddetis consuetum numerum laterum ".
EXOD|5|19|Videbantque se praefecti filiorum Israel in malo, eo quod diceretur eis: " Non minuetur quidquam de lateribus per singulos dies ";
EXOD|5|20|occurreruntque Moysi et Aaron, qui stabant ex adverso egredientibus a pharaone,
EXOD|5|21|et dixerunt ad eos: " Videat Dominus et iudicet, quoniam foetere fecistis odorem nostrum coram pharaone et servis eius; et praebuistis ei gladium, ut occideret nos ".
EXOD|5|22|Reversusque est Moyses ad Dominum et ait: " Domine, cur afflixisti populum istum? Quare misisti me?
EXOD|5|23|Ex eo enim quo ingressus sum ad pharaonem, ut loquerer in nomine tuo, afflixit populum tuum; et non liberasti eos ".
EXOD|6|1|Dixitque Dominus ad Moysen: " Nunc videbis quae facturus sim pharaoni; per manum enim fortem dimittet eos et in manu robusta eiciet illos de terra sua ".
EXOD|6|2|Locutusque est Dominus ad Moysen dicens: " Ego Dominus,
EXOD|6|3|qui apparui Abraham, Isaac et Iacob ut Deus omnipotens; et nomen meum Dominum non indicavi eis.
EXOD|6|4|Pepigique cum eis foedus, ut darem illis terram Chanaan, terram peregrinationis eorum, in qua fuerunt advenae.
EXOD|6|5|Ego audivi gemitum filiorum Israel, quia Aegyptii oppresserunt eos, et recordatus sum pacti mei.
EXOD|6|6|Ideo dic filiis Israel: Ego Dominus, qui educam vos de ergastulo Aegyptiorum; et eruam de servitute ac redimam in brachio excelso et iudiciis magnis.
EXOD|6|7|Et assumam vos mihi in populum et ero vester Deus; et scietis quod ego sum Dominus Deus vester, qui eduxerim vos de ergastulo Aegyptiorum
EXOD|6|8|et induxerim in terram, super quam levavi manum meam, ut darem eam Abraham, Isaac et Iacob; daboque illam vobis possidendam, ego Dominus ".
EXOD|6|9|Narravit ergo Moyses omnia filiis Israel; qui non acquieverunt ei propter angustiam spiritus et opus durissimum.
EXOD|6|10|Locutusque est Dominus ad Moysen dicens:
EXOD|6|11|" Ingredere et loquere ad pharaonem regem Aegypti, ut dimittat filios Israel de terra sua ".
EXOD|6|12|Respondit Moyses coram Domino: " Ecce, filii Israel non audiunt me, et quomodo audiet me pharao, praesertim cum incircumcisus sim labiis? ".
EXOD|6|13|Locutusque est Dominus ad Moysen et Aaron et dedit mandatum ad filios Israel et ad pharaonem regem Aegypti, ut educerent filios Israel de terra Aegypti.
EXOD|6|14|Isti sunt principes domorum per familias suas.Filii Ruben primogeniti Israelis: Henoch et Phallu, Hesron et Charmi; hae cognationes Ruben.
EXOD|6|15|Filii Simeon: Iamuel et Iamin et Ahod et Iachin et Sohar er Saul filius Chananitidis; hae progenies Simeon.
EXOD|6|16|Et haec nomina filiorum Levi per cognationes suas: Gerson et Caath et Merari; anni autem vitae Levi fuerunt centum triginta septem.
EXOD|6|17|Filii Gerson: Lobni et Semei per cognationes suas.
EXOD|6|18|Filii Caath: Amram et Isaar et Hebron et Oziel; anni quoque vitae Caath centum triginta tres.
EXOD|6|19|Filii Merari: Moholi et Musi; hae cognationes Levi per familias suas.
EXOD|6|20|Accepit autem Amram uxorem Iochabed amitam suam, quae peperit ei Aaron et Moysen; fueruntque anni vitae Amram centum triginta septem.
EXOD|6|21|Filii quoque Isaar: Core et Napheg et Zechri.
EXOD|6|22|Filii quoque Oziel: Misael et Elisaphan et Sethri.
EXOD|6|23|Accepit autem Aaron uxorem Elisabeth filiam Aminadab sororem Naasson, quae peperit ei Nadab et Abiu et Eleazar et Ithamar.
EXOD|6|24|Filii quoque Core: Asir et Elcana et Abiasaph; hae sunt cognationes Coritarum.
EXOD|6|25|At vero Eleazar filius Aaron accepit uxorem de filiabus Phutiel, quae peperit ei Phinees; hi sunt principes familiarum Leviticarum per cognationes suas.
EXOD|6|26|Iste est Aaron et Moyses, quibus praecepit Dominus, ut educerent filios Israel de terra Aegypti per turmas suas.
EXOD|6|27|Hi sunt qui loquuntur ad pharaonem regem Aegypti, ut educant filios Israel de Aegypto; iste est Moyses et Aaron
EXOD|6|28|in die, qua locutus est Dominus ad Moysen in terra Aegypti.
EXOD|6|29|Et locutus est Dominus ad Moysen dicens: " Ego Dominus; loquere ad pharaonem regem Aegypti omnia, quae ego loquor tibi ".
EXOD|6|30|Et ait Moyses coram Domino: " En incircumcisus labiis sum. Quomodo audiet me pharao? ".
EXOD|7|1|Dixitque Dominus ad Moysen: " Ecce constitui te deum pha raonis, et Aaron frater tuus erit propheta tuus.
EXOD|7|2|Tu loqueris omnia, quae mando tibi; et ille loquetur ad pharaonem, ut dimittat filios Israel de terra sua.
EXOD|7|3|Sed ego indurabo cor eius et multiplicabo signa et ostenta mea in terra Aegypti.
EXOD|7|4|Et non audiet vos; immittamque manum meam super Aegyptum et educam exercitum et populum meum, filios Israel, de terra Aegypti per iudicia maxima.
EXOD|7|5|Et scient Aegyptii quia ego sum Dominus, qui extenderim manum meam super Aegyptum et eduxerim filios Israel de medio eorum ".
EXOD|7|6|Fecit itaque Moyses et Aaron, sicut praeceperat Dominus; ita egerunt.
EXOD|7|7|Erat autem Moyses octoginta annorum, et Aaron octoginta trium, quando locuti sunt ad pharaonem.
EXOD|7|8|Dixitque Dominus ad Moysen et Aaron:
EXOD|7|9|" Cum dixerit vobis pharao: "Ostendite signum", dices ad Aaron: Tolle virgam tuam et proice eam coram pharaone, ac vertetur in colubrum ".
EXOD|7|10|Ingressi itaque Moyses et Aaron ad pharaonem fecerunt, sicut praeceperat Dominus; proiecitque Aaron virgam coram pharaone et servis eius, quae versa est in colubrum.
EXOD|7|11|Vocavit autem pharao sapientes et maleficos, et fecerunt etiam ipsi magi Aegypti per incantationes suas similiter.
EXOD|7|12|Proieceruntque singuli virgas suas, quae versae sunt in colubros; sed devoravit virga Aaron virgas eorum.
EXOD|7|13|Induratumque est cor pharaonis, et non audivit eos, sicut dixerat Dominus.
EXOD|7|14|Dixit autem Dominus ad Moysen: " Ingravatum est cor pharaonis: non vult dimittere populum.
EXOD|7|15|Vade ad eum mane. Ecce egredietur ad aquas; et stabis in occursum eius super ripam fluminis. Et virgam, quae conversa est in serpentem, tolles in manu tua
EXOD|7|16|dicesque ad eum: Dominus, Deus Hebraeorum, misit me ad te dicens: Dimitte populum meum, ut sacrificet mihi in deserto; et usque ad praesens audire noluisti.
EXOD|7|17|Haec igitur dicit Dominus: In hoc scies quod sim Dominus: ecce percutiam virga, quae in manu mea est, aquam fluminis; et vertetur in sanguinem.
EXOD|7|18|Pisces quoque, qui sunt in fluvio, morientur, et computrescent aquae, et taedebit Aegyptios bibere aquam fluminis ".
EXOD|7|19|Dixit quoque Dominus ad Moysen: " Dic ad Aaron: Tolle virgam tuam et extende manum tuam super aquas Aegypti, super fluvios eorum et rivos ac paludes et omnes lacus aquarum, ut vertantur in sanguinem; et sit cruor in omni terra Aegypti, tam in ligneis vasis quam in saxeis ".
EXOD|7|20|Feceruntque ita Moyses et Aaron, sicut praeceperat Dominus. Et elevans virgam percussit aquam fluminis coram pharaone et servis eius; quae versa est in sanguinem.
EXOD|7|21|Et pisces, qui erant in flumine, mortui sunt, computruitque fluvius, et non poterant Aegyptii bibere aquam fluminis; et fuit sanguis in tota terra Aegypti.
EXOD|7|22|Feceruntque similiter malefici Aegyptiorum incantationibus suis; et induratum est cor pharaonis, nec audivit eos, sicut dixerat Dominus.
EXOD|7|23|Avertitque se et ingressus est domum suam nec ad hoc apposuit cor suum.
EXOD|7|24|Foderunt autem omnes Aegyptii per circuitum fluminis aquam, ut biberent; non enim poterant bibere de aqua fluminis.
EXOD|7|25|Impletique sunt septem dies, postquam percussit Dominus fluvium.
EXOD|7|26|Dixit quoque Dominus ad Moysen: " Ingredere ad pharaonem et dices ad eum: Haec dicit Dominus: Dimitte populum meum, ut sacrificet mihi.
EXOD|7|27|Sin autem nolueris dimittere, ecce ego percutiam omnes terminos tuos ranis.
EXOD|7|28|Et ebulliet fluvius ranas, quae ascendent et ingredientur domum tuam et cubiculum lectuli tui et super stratum tuum et in domos servorum tuorum et in populum tuum et in furnos tuos et in pistrina tua;
EXOD|7|29|et ad te et ad populum tuum et ad omnes servos tuos intrabunt ranae ".
EXOD|8|1|Dixitque Dominus ad Moysen: " Dic ad Aaron: Extende ma num tuam cum baculo tuo super fluvios, super rivos ac paludes et educ ranas super terram Aegypti ".
EXOD|8|2|Et extendit Aaron manum super aquas Aegypti, et ascenderunt ranae operueruntque terram Aegypti.
EXOD|8|3|Fecerunt autem et malefici per incantationes suas similiter eduxeruntque ranas super terram Aegypti.
EXOD|8|4|Vocavit autem pharao Moysen et Aaron et dixit: " Orate Dominum, ut auferat ranas a me et a populo meo, et dimittam populum, ut sacrificet Domino ".
EXOD|8|5|Dixitque Moyses ad pharaonem: " Constitue mihi, quando deprecer pro te et pro servis et pro populo tuo, ut abigantur ranae a te et a domo tua et tantum in flumine remaneant ".
EXOD|8|6|Qui respondit: " Cras ". At ille: " Iuxta verbum, inquit, tuum faciam, ut scias quoniam non est sicut Dominus Deus noster.
EXOD|8|7|Et recedent ranae a te et a domo tua et a servis tuis et a populo tuo; tantum in flumine remanebunt ".
EXOD|8|8|Egressique sunt Moyses et Aaron a pharaone; et clamavit Moyses ad Dominum pro sponsione ranarum, quam condixerat pharaoni.
EXOD|8|9|Fecitque Dominus iuxta verbum Moysi, et mortuae sunt ranae de domibus et de villis et de agris;
EXOD|8|10|congregaveruntque eas in immensos aggeres, et computruit terra.
EXOD|8|11|Videns autem pharao quod data esset requies, ingravavit cor suum et non audivit eos, sicut dixerat Dominus.
EXOD|8|12|Dixitque Dominus ad Moysen: " Loquere ad Aaron: Extende virgam tuam et percute pulverem terrae, et sint scinifes in universa terra Aegypti ".
EXOD|8|13|Feceruntque ita; et extendit Aaron manum virgam tenens percussitque pulverem terrae. Et facti sunt scinifes in hominibus et in iumentis; omnis pulvis terrae versus est in scinifes per totam terram Aegypti.
EXOD|8|14|Feceruntque similiter malefici incantationibus suis, ut educerent scinifes; et non potuerunt. Erantque scinifes tam in hominibus quam in iumentis;
EXOD|8|15|et dixerunt malefici ad pharaonem: " Digitus Dei est hic ". Induratumque est cor pharaonis et non audivit eos, sicut praeceperat Dominus.
EXOD|8|16|Dixit quoque Dominus ad Moysen: " Consurge diluculo et sta coram pharaone. Egredietur enim ad aquas, et dices ad eum: Haec dicit Dominus: Dimitte populum meum, ut sacrificet mihi.
EXOD|8|17|Quod si non dimiseris eum, ecce ego immittam in te et in servos tuos et in populum tuum et in domos tuas omne genus muscarum; et implebuntur domus Aegyptiorum muscis et etiam humus, in qua fuerint.
EXOD|8|18|Et segregabo in die illa terram Gessen, in qua populus meus est, ut non sint ibi muscae, et scias quoniam ego Dominus in medio terrae;
EXOD|8|19|ponamque divi sionem inter populum meum et populum tuum; cras erit signum istud ".
EXOD|8|20|Fecitque Dominus ita; et venit musca gravissima in domos pharaonis et servorum eius et in omnem terram Aegypti, corruptaque est terra ab huiuscemodi muscis.
EXOD|8|21|Vocavitque pharao Moysen et Aaron et ait eis: " Ite, sacrificate Deo vestro in terra ".
EXOD|8|22|Et ait Moyses: " Non potest ita fieri: abominationes enim Aegyptiorum immolabimus Domino Deo nostro; quod si mactaverimus ea, quae colunt Aegyptii, coram eis, lapidibus nos obruent.
EXOD|8|23|Viam trium dierum pergemus in solitudinem et sacrificabimus Domino Deo nostro, sicut praecepit nobis ".
EXOD|8|24|Dixitque pharao: " Ego dimittam vos, ut sacrificetis Domino Deo vestro in deserto, verumtamen longius ne abeatis; rogate pro me ".
EXOD|8|25|Et ait Moyses: " Egressus a te, orabo Dominum, et recedet musca a pharaone et a servis suis et a populo eius cras; verumtamen noli ultra fallere, ut non dimittas populum sacrificare Domino ".
EXOD|8|26|Egressusque Moyses a pharaone oravit Dominum;
EXOD|8|27|qui fecit iuxta verbum illius et abstulit muscas a pharaone et a servis suis et a populo eius; non superfuit ne una quidem.
EXOD|8|28|Et ingravatum est cor pharaonis, ita ut ne hac quidem vice dimitteret populum.
EXOD|9|1|Dixit autem Dominus ad Moysen: " Ingredere ad pharaonem et loquere ad eum: Haec dicit Dominus, Deus Hebraeorum: Dimitte populum meum, ut sacrificet mihi.
EXOD|9|2|Quod si adhuc renuis et retines eos,
EXOD|9|3|ecce manus Domini erit super possessionem tuam in agris, super equos et asinos et camelos et boves et oves, pestis valde gravis;
EXOD|9|4|et distinguet Dominus inter possessiones Israel et possessiones Aegyptiorum, ut nihil omnino pereat ex his, quae pertinent ad filios Israel.
EXOD|9|5|Constituitque Dominus tempus dicens: Cras faciet Dominus verbum istud in terra ".
EXOD|9|6|Fecit ergo Dominus verbum hoc altera die, mortuaque sunt omnia animantia Aegyptiorum; de animalibus vero filiorum Israel nihil omnino periit.
EXOD|9|7|Et misit pharao ad videndum; nec erat quidquam mortuum de his, quae possidebat Israel. Ingravatumque est cor pharaonis, et non dimisit populum.
EXOD|9|8|Et dixit Dominus ad Moysen et Aaron: " Tollite plenas manus cineris de camino, et spargat illum Moyses in caelum coram pharaone;
EXOD|9|9|sitque pulvis super omnem terram Aegypti; erunt enim in hominibus et iumentis ulcera et vesicae turgentes in universa terra Aegypti ".
EXOD|9|10|Tuleruntque cinerem de camino et steterunt coram pharaone, et sparsit illum Moyses in caelum; factaque sunt ulcera vesicarum turgentium in hominibus et iumentis.
EXOD|9|11|Nec poterant malefici stare coram Moyse propter ulcera, quae in illis erant et in omni terra Aegypti.
EXOD|9|12|Induravitque Dominus cor pharaonis, et non audivit eos, sicut locutus est Dominus ad Moysen.
EXOD|9|13|Dixitque Dominus ad Moysen: " Mane consurge et sta coram pharaone et dices ad eum: Haec dicit Dominus, Deus Hebraeorum: Dimitte populum meum, ut sacrificet mihi;
EXOD|9|14|quia in hac vice mittam omnes plagas meas super cor tuum et super servos tuos et super populum tuum, ut scias quod non sit similis mei in omni terra.
EXOD|9|15|Nunc enim extendens manum si percussissem te et populum tuum peste, perisses de terra.
EXOD|9|16|Idcirco autem servavi te, ut ostendam in te fortitudinem meam, et narretur nomen meum in omni terra.
EXOD|9|17|Adhuc retines populum meum et non vis dimittere eum?
EXOD|9|18|En pluam cras, hac ipsa hora, grandinem multam nimis, qualis non fuit in Aegypto a die, qua fundata est, usque in praesens tempus.
EXOD|9|19|Mitte ergo iam nunc et congrega iumenta tua et omnia, quae habes in agro; homines enim et iumenta universa, quae inventa fuerint foris nec congregata de agris, cadet super ea grando, et morientur ".
EXOD|9|20|Qui timuit verbum Domini de servis pharaonis, fecit confugere servos suos et iumenta in domos;
EXOD|9|21|qui autem neglexit sermonem Domini, dimisit servos suos et iumenta in agris.
EXOD|9|22|Et dixit Dominus ad Moysen: " Extende manum tuam in caelum, ut fiat grando in universa terra Aegypti super homines et super iumenta et super omnem herbam agri in terra Aegypti ".
EXOD|9|23|Extenditque Moyses virgam in caelum, et Dominus dedit tonitrua et grandinem ac discurrentia fulgura super terram; pluitque Dominus grandinem super terram Aegypti.
EXOD|9|24|Et grando et ignis immixta pariter ferebantur; tantaeque fuit magnitudinis, quanta ante numquam apparuit in universa terra Aegypti, ex quo gens illa condita est.
EXOD|9|25|Et percussit grando in omni terra Aegypti cuncta, quae fuerunt in agris, ab homine usque ad iumentum; cunctamque herbam agri percussit grando et omne lignum regionis confregit.
EXOD|9|26|Tantum in terra Gessen, ubi erant filii Israel, grando non cecidit.
EXOD|9|27|Misitque pharao et vocavit Moysen et Aaron dicens ad eos: " Nunc peccavi; Dominus iustus, ego et populus meus rei.
EXOD|9|28|Orate Dominum, ut desinant tonitrua Dei et grando, et dimittam vos, et nequaquam hic ultra manebitis ".
EXOD|9|29|Ait Moyses: " Cum egressus fuero de urbe, extendam palmas meas ad Dominum; et cessabunt tonitrua, et grando non erit, ut scias quia Domini est terra.
EXOD|9|30|Novi autem quod et tu et servi tui necdum timeatis Dominum Deum ".
EXOD|9|31|Linum ergo et hordeum laesum est, eo quod hordeum iam spicas et linum iam folliculos germinaret;
EXOD|9|32|triticum autem et far non sunt laesa, quia serotina erant.
EXOD|9|33|Egressusque Moyses a pharaone ex urbe tetendit manus ad Dominum; et cessaverunt tonitrua et grando, nec ultra effundebatur pluvia super terram. 34 Videns autem pharao quod cessasset pluvia et grando et tonitrua, auxit peccatum; 35 et ingravatum est cor eius et servorum illius et induratum nimis; nec dimisit filios Israel, sicut dixerat Dominus per manum Moysi.
EXOD|10|1|Et dixit Dominus ad Moy sen: " Ingredere ad pharao nem: ego enim induravi cor eius et servorum illius, ut faciam signa mea haec in medio eorum,
EXOD|10|2|et narres in auribus filii tui et nepotum tuorum, quotiens contriverim Aegyptios et signa mea fecerim in eis; et sciatis quia ego Dominus ".
EXOD|10|3|Introierunt ergo Moyses et Aaron ad pharaonem et dixerunt ei: " Haec dicit Dominus, Deus Hebraeorum: Usquequo non vis subici mihi? Dimitte populum meum, ut sacrificet mihi.
EXOD|10|4|Sin autem resistis et non vis dimittere eum, ecce ego inducam cras locustam in fines tuos,
EXOD|10|5|quae operiat superficiem terrae, ne quidquam eius appareat, sed comedatur, quod residuum fuerit grandini; corrodet enim omnia ligna, quae germinant in agris.
EXOD|10|6|Et implebunt domos tuas et servorum tuorum et omnium Aegyptiorum, quantam non viderunt patres tui et avi, ex quo orti sunt super terram usque in praesentem diem ". Avertitque se et egressus est a pharaone.
EXOD|10|7|Dixerunt autem servi pharaonis ad eum: " Usquequo patiemur hoc scandalum? Dimitte homines, ut sacrificent Domino Deo suo; nonne vides quod perierit Aegyptus? ".
EXOD|10|8|Revocaveruntque Moysen et Aaron ad pharaonem, qui dixit eis: " Ite, sacrificate Domino Deo vestro. Quinam sunt qui ituri sunt? ".
EXOD|10|9|Ait Moyses: " Cum parvulis nostris et senioribus pergemus, cum filiis et filiabus, cum ovibus et armentis; est enim sollemnitas Domini nobis ".
EXOD|10|10|Et respondit eis: " Sic Dominus sit vobiscum, quomodo ego dimittam vos et parvulos vestros. Cui dubium est quod pessime cogitetis?
EXOD|10|11|Non fiet ita, sed ite tantum viri et sacrificate Domino; hoc enim et ipsi petistis ". Statimque eiecti sunt de conspectu pharaonis.
EXOD|10|12|Dixit autem Dominus ad Moysen: " Extende manum tuam super terram Aegypti, ut veniat locusta et ascendat super eam et devoret omnem herbam, quidquid residuum fuerit grandini ".
EXOD|10|13|Et extendit Moyses virgam super terram Aegypti, et Dominus induxit ventum urentem tota die illa et nocte. Et mane facto, ventus urens levavit locustas;
EXOD|10|14|quae ascenderunt super universam terram Aegypti et sederunt in cunctis finibus Aegyptiorum innumerabiles, quales ante illud tempus non fuerant nec postea futurae sunt.
EXOD|10|15|Operueruntque universam superficiem terrae, et obscurata est terra. Devoraverunt igitur omnem herbam terrae et, quidquid pomorum in arboribus fuit, quae grando dimiserat; nihilque omnino virens relictum est in lignis et in herbis terrae in cuncta Aegypto.
EXOD|10|16|Quam ob rem festinus pharao vocavit Moysen et Aaron et dixit eis: " Peccavi in Dominum Deum vestrum et in vos.
EXOD|10|17|Sed nunc dimittite peccatum mihi tantum hac vice et rogate Dominum Deum vestrum, ut auferat a me saltem mortem istam ".
EXOD|10|18|Egressusque Moyses de conspectu pharaonis oravit Dominum,
EXOD|10|19|qui flare fecit ventum ab occidente vehementissimum et arreptam locustam proiecit in mare Rubrum; non remansit ne una quidem in cunctis finibus Aegypti.
EXOD|10|20|Et induravit Dominus cor pharaonis, nec dimisit filios Israel.
EXOD|10|21|Dixit autem Dominus ad Moysen: " Extende manum tuam in caelum, et sint tenebrae super terram Aegypti tam densae ut palpari queant ".
EXOD|10|22|Extenditque Moyses manum in caelum, et factae sunt tenebrae horribiles in universa terra Aegypti tribus diebus.
EXOD|10|23|Nemo vidit fratrem suum nec movit se de loco, in quo erat. Ubicumque autem habitabant filii Israel, lux erat.
EXOD|10|24|Vocavitque pharao Moysen et Aaron et dixit eis: " Ite, sacrificate Domino; oves tantum vestrae et armenta remaneant, parvuli vestri eant vobiscum ".
EXOD|10|25|Ait Moyses: " Etiamsi tu hostias et holocausta dares nobis, quae offeramus Domino Deo nostro,
EXOD|10|26|tamen et greges nostri pergent nobiscum; non remanebit ex eis ungula, quoniam ex ipsis sumemus, quae necessaria sunt in cultum Domini Dei nostri; praesertim cum ignoremus quid debeat immolari, donec ad ipsum locum perveniamus ".
EXOD|10|27|Induravit autem Dominus cor pharaonis, et noluit dimittere eos.
EXOD|10|28|Dixitque pharao ad eum: " Recede a me. Cave, ne ultra videas faciem meam; quocumque die apparueris mihi, morieris ".
EXOD|10|29|Respondit Moyses: " Ita fiet, ut locutus es; non videbo ultra faciem tuam ".
EXOD|11|1|Et dixit Dominus ad Moy sen: " Adhuc una plaga tan gam pharaonem et Aegyptum, et post haec dimittet vos utique, immo et exire compellet.
EXOD|11|2|Dices ergo omni plebi, ut postulet vir ab amico suo et mulier a vicina sua vasa argentea et aurea;
EXOD|11|3|dabit autem Dominus gratiam populo coram Aegyptiis ". Fuitque Moyses vir magnus valde in terra Aegypti coram servis pharaonis et omni populo.
EXOD|11|4|Et ait Moyses: " Haec dicit Dominus: Media nocte egrediar in Aegyptum;
EXOD|11|5|et morietur omne primogenitum in terra Aegyptiorum, a primogenito pharaonis, qui sedet in solio eius, usque ad primogenitum ancillae, quae est ad molam, et omnia primogenita iumentorum.
EXOD|11|6|Eritque clamor magnus in universa terra Aegypti, qualis nec ante fuit nec postea futurus est.
EXOD|11|7|Apud omnes autem filios Israel non mutiet canis contra hominem et pecus, ut sciatis quanto miraculo dividat Dominus Aegyptios et Israel.
EXOD|11|8|Descendentque omnes servi tui isti ad me et adorabunt me dicentes: "Egredere tu et omnis populus, qui sequitur te". Post haec egrediar ". Et exivit a pharaone iratus nimis.
EXOD|11|9|Dixit autem Dominus ad Moysen: " Non audiet vos pharao, ut multa signa fiant in terra Aegypti ".
EXOD|11|10|Moyses autem et Aaron fecerunt omnia ostenta haec coram pharaone; et induravit Dominus cor pharaonis, nec dimisit filios Israel de terra sua.
EXOD|12|1|Dixit Dominus ad Moysen et Aaron in terra Aegypti:
EXOD|12|2|" Mensis iste vobis principium mensium, primus erit in mensibus anni.
EXOD|12|3|Loquimini ad universum coetum filiorum Israel et dicite eis: Decima die mensis huius tollat unusquisque agnum per familias et domos suas.
EXOD|12|4|Sin autem minor est numerus, ut sufficere possit ad vescendum agnum, assumet vicinum suum, qui iunctus est domui suae, iuxta numerum animarum, quae sufficere possunt ad esum agni.
EXOD|12|5|Erit autem vobis agnus absque macula, masculus, anniculus; quem de agnis vel haedis tolletis
EXOD|12|6|et servabitis eum usque ad quartam decimam diem mensis huius; immolabitque eum universa congregatio filiorum Israel ad vesperam.
EXOD|12|7|Et sument de sanguine eius ac ponent super utrumque postem et in superliminaribus domorum, in quibus comedent illum;
EXOD|12|8|et edent carnes nocte illa assas igni et azymos panes cum lactucis amaris.
EXOD|12|9|Non comedetis ex eo crudum quid nec coctum aqua, sed tantum assum igni; caput cum pedibus eius et intestinis vorabitis.
EXOD|12|10|Nec remanebit quidquam ex eo usque mane; si quid residuum fuerit, igne comburetis.
EXOD|12|11|Sic autem comedetis illum: renes vestros accingetis, calceamenta habebitis in pedibus, tenentes baculos in manibus, et comedetis festinanter; est enim Pascha (id est Transitus) Domini!
EXOD|12|12|Et transibo per terram Aegypti nocte illa percutiamque omne primogenitum in terra Aegypti ab homine usque ad pecus; et in cunctis diis Aegypti faciam iudicia, ego Dominus.
EXOD|12|13|Erit autem sanguis vobis in signum in aedibus, in quibus eritis; et videbo sanguinem et transibo vos, nec erit in vobis plaga disperdens, quando percussero terram Aegypti.
EXOD|12|14|Habebitis autem hanc diem in monumentum et celebrabitis eam sollemnem Domino in generationibus vestris cultu sempiterno.
EXOD|12|15|Septem diebus azyma comedetis. Iam in die primo non erit fermentum in domibus vestris; quicumque comederit fermentatum, a primo die usque ad diem septimum, peribit anima illa de Israel.
EXOD|12|16|Dies prima erit sancta atque sollemnis, et dies septima eadem festivitate venerabilis. Nihil operis facietis in eis, exceptis his, quae ad vescendum pertinent.
EXOD|12|17|Et observabitis azyma, in eadem enim ipsa die eduxi exercitum vestrum de terra Aegypti; et custodietis diem istum in generationes vestras ritu perpetuo.
EXOD|12|18|Primo mense, quarta decima die mensis ad vesperam comedetis azyma; usque ad diem vicesimam primam eiusdem mensis ad vesperam.
EXOD|12|19|Septem diebus fermentum non invenietur in domibus vestris. Qui comederit fermentatum, peribit anima eius de coetu Israel, tam de advenis quam de indigenis terrae.
EXOD|12|20|Omne fermentatum non comedetis; in cunctis habitaculis vestris edetis azyma ".
EXOD|12|21|Vocavit autem Moyses omnes seniores filiorum Israel et dixit ad eos: " Ite tollentes animal per familias vestras et immolate Pascha.
EXOD|12|22|Fasciculumque hyssopi tingite in sanguine, qui est in pelvi, et aspergite ex eo superliminare et utrumque postem. Nullus vestrum egrediatur ostium domus suae usque mane.
EXOD|12|23|Transibit enim Dominus percutiens Aegyptios; cumque viderit sanguinem in superliminari et in utroque poste, transcendet ostium et non sinet percussorem ingredi domos vestras et laedere.
EXOD|12|24|Custodite verbum istud legitimum tibi et filiis tuis usque in aeternum.
EXOD|12|25|Cumque introieritis terram, quam Dominus daturus est vobis, ut pollicitus est, observabitis caeremonias istas;
EXOD|12|26|et, cum dixerint vobis filii vestri: "Quae est ista religio?",
EXOD|12|27|dicetis eis: "Victima Paschae Domino est, quando transivit super domos filiorum Israel in Aegypto percutiens Aegyptios et domos nostras liberans" ". Incurvatusque populus adoravit;
EXOD|12|28|et egressi filii Israel fecerunt, sicut praeceperat Dominus Moysi et Aaron.
EXOD|12|29|Factum est autem in noctis medio, percussit Dominus omne primogenitum in terra Aegypti, a primogenito pharaonis, qui in solio eius sedebat, usque ad primogenitum captivi, qui erat in carcere, et omne primogenitum iumentorum.
EXOD|12|30|Surrexitque pharao nocte et omnes servi eius cunctaque Aegyptus, et ortus est clamor magnus in Aegypto, neque enim erat domus, in qua non iaceret mortuus.
EXOD|12|31|Vocatisque pharao Moyse et Aaron nocte, ait: " Surgite, egredimini a populo meo, vos et filii Israel; ite, immolate Domino, sicut dicitis.
EXOD|12|32|Oves vestras et armenta assumite, ut petieratis, et abeuntes benedicite mihi ".
EXOD|12|33|Urgebantque Aegyptii populum de terra exire velociter dicentes: " Omnes moriemur ".
EXOD|12|34|Tulit igitur populus conspersam farinam, antequam fermentaretur; et ligans pistrina in palliis suis posuit super umeros suos.
EXOD|12|35|Feceruntque filii Israel, sicut praeceperat Moyses, et petierunt ab Aegyptiis vasa argentea et aurea vestemque plurimam.
EXOD|12|36|Dominus autem dedit gratiam populo coram Aegyptiis, ut commodarent eis; et spoliaverunt Aegyptios.
EXOD|12|37|Profectique sunt filii Israel de Ramesse in Succoth, sescenta fere milia peditum virorum absque parvulis.
EXOD|12|38|Sed et vulgus promiscuum innumerabile ascendit cum eis, oves et armenta, animantia multa nimis.
EXOD|12|39|Coxeruntque farinam, quam dudum de Aegypto conspersam tulerant, et fecerunt subcinericios panes azymos; neque enim poterant fermentari, cogentibus exire Aegyptiis et nullam facere sinentibus moram; nec pulmenti quidquam occurrerant praeparare.
EXOD|12|40|Habitatio autem filiorum Israel, qua manserant in Aegypto, fuit quadringentorum triginta annorum.
EXOD|12|41|Quibus expletis, eadem die egressus est omnis exercitus Domini de terra Aegypti.
EXOD|12|42|Nox ista vigiliarum Domino, quando eduxit eos de terra Aegypti: hanc observare debent Domino omnes filii Israel in generationibus suis.
EXOD|12|43|Dixitque Dominus ad Moysen et Aaron: " Haec est religio Paschae: Omnis alienigena non comedet ex eo;
EXOD|12|44|omnis autem servus empticius circumcidetur et sic comedet;
EXOD|12|45|advena et mercennarius non edent ex eo.
EXOD|12|46|In una domo comedetur, nec efferetis de carnibus eius foras nec os illius confringetis.
EXOD|12|47|Omnis coetus filiorum Israel faciet illud.
EXOD|12|48|Quod si quis peregrinorum in vestram voluerit transire coloniam et facere Pascha Domini, circumcidetur prius omne masculinum eius, et tunc rite celebrabit eritque sicut indigena terrae; si quis autem circumcisus non fuerit, non vescetur ex eo.
EXOD|12|49|Eadem lex erit indigenae et colono, qui peregrinatur apud vos ".
EXOD|12|50|Feceruntque omnes filii Israel, sicut praeceperat Dominus Moysi et Aaron;
EXOD|12|51|et in eadem die eduxit Dominus filios Israel de terra Aegypti per turmas suas.
EXOD|13|1|Locutusque est Dominus ad Moysen dicens:
EXOD|13|2|" Sanctifica mihi omne primogenitum, quod aperit vulvam in filiis Israel, tam de hominibus quam de iumentis: mea sunt enim omnia ".
EXOD|13|3|Et ait Moyses ad populum: " Mementote diei huius, in qua egressi estis de Aegypto et de domo servitutis, quoniam in manu forti eduxit vos Dominus de loco isto, ut non comedatis fermentatum panem.
EXOD|13|4|Hodie egredimini, mense Abib (id est novarum Frugum).
EXOD|13|5|Cumque introduxerit te Dominus in terram Chananaei et Hetthaei et Amorraei et Hevaei et Iebusaei, quam iuravit patribus tuis, ut daret tibi, terram fluentem lacte et melle; celebrabis hunc morem sacrorum mense isto.
EXOD|13|6|Septem diebus vesceris azymis, et in die septimo erit sollemnitas Domini.
EXOD|13|7|Azyma comedetis septem diebus: non apparebit apud te aliquid fermentatum nec in cunctis finibus tuis.
EXOD|13|8|Narrabisque filio tuo in die illo dicens: "Propter hoc, quod fecit mihi Dominus, quando egressus sum de Aegypto".
EXOD|13|9|Et erit quasi signum in manu tua et quasi monumentum inter oculos tuos, ut lex Domini semper sit in ore tuo; in manu enim forti eduxit te Dominus de Aegypto.
EXOD|13|10|Custodies huiuscemodi cultum statuto tempore a diebus in dies.
EXOD|13|11|Cumque introduxerit te Dominus in terram Chananaei, sicut iuravit tibi et patribus tuis, et dederit tibi eam,
EXOD|13|12|separabis omne, quod aperit vulvam, Domino et quod primitivum est in pecoribus tuis; quidquid habueris masculini sexus, consecrabis Domino.
EXOD|13|13|Primogenitum asini mutabis ove; quod, si non redemeris, interficies. Omne autem primogenitum hominis de filiis tuis pretio redimes.
EXOD|13|14|Cumque interrogaverit te filius tuus cras dicens: "Quid est hoc?", respondebis ei: "In manu forti eduxit nos Dominus de Aegypto, de domo servitutis.
EXOD|13|15|Nam, cum induratus esset pharao et nollet nos dimittere, occidit Dominus omne primogenitum in terra Aegypti, a primogenito hominis usque ad primogenitum iumentorum; idcirco immolo Domino omne, quod aperit vulvam, masculini sexus, et omnia primogenita filiorum meorum redimo".
EXOD|13|16|Erit igitur quasi signum in manu tua et quasi appensum quid ob recordationem inter oculos tuos, eo quod in manu forti eduxit nos Dominus de Aegypto ".
EXOD|13|17|Igitur cum emisisset pharao populum, non eos duxit Deus per viam terrae Philisthim, quae vicina est, reputans ne forte paeniteret populum, si vidisset adversum se bella consurgere, et reverteretur in Aegyptum,
EXOD|13|18|sed circumduxit per viam deserti, quae est iuxta mare Rubrum. Et armati ascenderunt filii Israel de terra Aegypti.
EXOD|13|19|Tulit quoque Moyses ossa Ioseph secum, eo quod adiurasset filios Israel dicens: " Visitabit vos Deus; efferte ossa mea hinc vobiscum ".
EXOD|13|20|Profectique de Succoth castrametati sunt in Etham, in extremis finibus solitudinis.
EXOD|13|21|Dominus autem praecedebat eos ad ostendendam viam per diem in columna nubis et per noctem in columna ignis, ut dux esset itineris utroque tempore.
EXOD|13|22|Nunquam defuit columna nubis per diem, nec columna ignis per noctem, coram populo.
EXOD|14|1|Locutus est autem Dominus ad Moysen dicens:
EXOD|14|2|" Lo quere filiis Israel: Reversi castrametentur e regione Phihahiroth, quae est inter Magdolum et mare contra Beelsephon; in conspectu eius castra ponetis super mare.
EXOD|14|3|Dicturusque est pharao super filiis Israel: "Errant in terra, conclusit eos desertum".
EXOD|14|4|Et indurabo cor eius, ac persequetur eos, et glorificabor in pharaone et in omni exercitu eius; scientque Aegyptii quia ego sum Dominus ". Feceruntque ita.
EXOD|14|5|Et nuntiatum est regi Aegyptiorum quod fugisset populus; immutatumque est cor pharaonis et servorum eius super populo, et dixerunt: " Quid hoc fecimus, ut dimitteremus Israel, ne servirent nobis? ".
EXOD|14|6|Iunxit ergo currum et omnem populum suum assumpsit secum;
EXOD|14|7|tulitque sescentos currus electos et quidquid in Aegypto curruum fuit et bellatores in singulis curribus.
EXOD|14|8|Induravitque Dominus cor pharaonis regis Aegypti, et persecutus est filios Israel; at illi egressi erant in manu excelsa.
EXOD|14|9|Cumque persequerentur Aegyptii vestigia praecedentium, reppererunt eos in castris super mare; omnes equi et currus pharaonis, equites et exercitus eius erant in Phihahiroth contra Beelsephon.
EXOD|14|10|Cumque appropinquasset pharao, levantes filii Israel oculos viderunt Aegyptios post se et timuerunt valde clamaveruntque ad Dominum
EXOD|14|11|et dixerunt ad Moysen: " Forsitan non erant sepulcra in Aegypto? Ideo tulisti nos, ut moreremur in solitudine. Quid hoc fecisti, ut educeres nos ex Aegypto?
EXOD|14|12|Nonne iste est sermo, quem loquebamur ad te in Aegypto dicentes: Recede a nobis, ut serviamus Aegyptiis? Multo enim melius erat servire eis quam mori in solitudine ".
EXOD|14|13|Et ait Moyses ad populum: " Nolite timere; state et videte salutem Domini, quam facturus est vobis hodie; Aegyptios enim, quos nunc videtis, nequaquam ultra videbitis usque in sempiternum.
EXOD|14|14|Dominus pugnabit pro vobis, et vos silebitis ".
EXOD|14|15|Dixitque Dominus ad Moysen: " Quid clamas ad me? Loquere filiis Israel, ut proficiscantur.
EXOD|14|16|Tu autem eleva virgam tuam et extende manum tuam super mare et divide illud, ut gradiantur filii Israel in medio mari per siccum.
EXOD|14|17|Ego autem indurabo cor Aegyptiorum, ut persequantur eos; et glorificabor in pharaone et in omni exercitu eius, in curribus et in equitibus illius.
EXOD|14|18|Et scient Aegyptii quia ego sum Dominus, cum glorificatus fuero in pharaone, in curribus atque in equitibus eius ".
EXOD|14|19|Tollensque se angelus Dei, qui praecedebat castra Israel, abiit post eos; et cum eo pariter columna nubis, priora dimittens, post tergum.
EXOD|14|20|Stetit inter castra Aegyptiorum et castra Israel; et erat nubes tenebrosa et illuminans noctem, ita ut ad se invicem toto noctis tempore accedere non valerent.
EXOD|14|21|Cumque extendisset Moyses manum super mare, reppulit illud Dominus, flante vento vehementi et urente tota nocte, et vertit in siccum; divisaque est aqua.
EXOD|14|22|Et ingressi sunt filii Israel per medium maris sicci; erat enim aqua quasi murus a dextra eorum et laeva.
EXOD|14|23|Persequentesque Aegyptii ingressi sunt post eos, omnis equitatus pharaonis, currus eius et equites per medium maris.
EXOD|14|24|Iamque advenerat vigilia matutina, et ecce respiciens Dominus super castra Aegyptiorum per columnam ignis et nubis perturbavit exercitum eorum;
EXOD|14|25|et impedivit rotas curruum, ita ut difficile moverentur. Dixerunt ergo Aegyptii: " Fugiamus Israelem! Dominus enim pugnat pro eis contra nos ".
EXOD|14|26|Et ait Dominus ad Moysen: " Extende manum tuam super mare, ut revertantur aquae ad Aegyptios super currus et equites eorum ".
EXOD|14|27|Cumque extendisset Moyses manum contra mare, reversum est primo diluculo ad priorem locum; fugientibusque Aegyptiis occurrerunt aquae, et involvit eos Dominus in mediis fluctibus.
EXOD|14|28|Reversaeque sunt aquae et operuerunt currus et equites cuncti exercitus pharaonis, qui sequentes ingressi fuerant mare; ne unus quidem superfuit ex eis.
EXOD|14|29|Filii autem Israel perrexerunt per medium sicci maris, et aquae eis erant quasi pro muro a dextris et a sinistris.
EXOD|14|30|Liberavitque Dominus in die illo Israel de manu Aegyptiorum. Et viderunt Aegyptios mortuos super litus maris
EXOD|14|31|et manum magnam, quam exercuerat Dominus contra eos; timuitque populus Dominum et crediderunt Domino et Moysi servo eius.
EXOD|15|1|Tunc cecinit Moyses et filii Israel carmen hoc Domino, et dixerunt:" Cantemus Domino,gloriose enim magnificatus est:equum et ascensorem eiusdeiecit in mare!
EXOD|15|2|Fortitudo mea et robur meum Dominus,et factus est mihi in salutem.Iste Deus meus,et glorificabo eum;Deus patris mei,et exaltabo eum!
EXOD|15|3|Dominus quasi vir pugnator;Dominus nomen eius!
EXOD|15|4|Currus pharaonis et exercitum eiusproiecit in mare;electi bellatores eiussubmersi sunt in mari Rubro.
EXOD|15|5|Abyssi operuerunt eos,descenderunt in profundum quasi lapis.
EXOD|15|6|Dextera tua, Domine,magnifice in fortitudine,dextera tua, Domine,percussit inimicum.
EXOD|15|7|Et in multitudine gloriae tuaedeposuisti adversarios tuos;misisti iram tuam,quae devoravit eos sicut stipulam.
EXOD|15|8|Et in spiritu furoris tuicongregatae sunt aquae;stetit ut aggerunda fluens,coagulatae sunt abyssiin medio mari.
EXOD|15|9|Dixit inimicus:"Persequar, comprehendam,dividam spolia,implebitur anima mea;evaginabo gladium meum,interficiet eos manus mea!".
EXOD|15|10|Flavit spiritus tuus,et operuit eos mare;submersi sunt quasi plumbumin aquis vehementibus.
EXOD|15|11|Quis similis tuiin diis, Domine?Quis similis tui,magnificus in sanctitate,terribilis atque laudabilis,faciens mirabilia?
EXOD|15|12|Extendisti manum tuam,devoravit eos terra.
EXOD|15|13|Dux fuisti in misericordia tuapopulo, quem redemisti,et portasti eum in fortitudine tuaad habitaculum sanctum tuum.
EXOD|15|14|Attenderunt populi et commoti sunt,dolores obtinuerunt habitatores Philisthaeae.
EXOD|15|15|Tunc conturbati sunt principes Edom,potentes Moab obtinuit tremor,obriguerunt omnes habitatores Chanaan.
EXOD|15|16|Irruit super eosformido et pavor;in magnitudine brachii tuifiunt immobiles quasi lapis,donec pertranseat populus tuus, Domine,donec pertranseat populus tuus iste,quem possedisti.
EXOD|15|17|Introduces eos et plantabisin monte hereditatis tuae,firmissimo habitaculo tuo,quod operatus es, Domine,sanctuario, Domine,quod firmaverunt manus tuae.
EXOD|15|18|Dominus regnabitin aeternum et ultra! ".
EXOD|15|19|Ingressi sunt enim equi pharaonis cum curribus et equitibus eius in mare, et reduxit super eos Dominus aquas maris; filii autem Israel ambu laverunt per siccum in medio eius.
EXOD|15|20|Sumpsit ergo Maria prophetissa soror Aaron tympanum in manu sua; egressaeque sunt omnes mulieres post eam cum tympanis et choris,
EXOD|15|21|quibus praecinebat dicens:" Cantemus Domino,gloriose enim magnificatus est:equum et ascensorem eiusdeiecit in mare! ".
EXOD|15|22|Tulit autem Moyses Israel de mari Rubro, et egressi sunt in desertum Sur; ambulaveruntque tribus diebus per solitudinem et non inveniebant aquam.
EXOD|15|23|Et venerunt in Mara nec poterant bibere aquas de Mara, eo quod essent amarae; unde vocatum est nomen eius Mara (id est Amaritudo).
EXOD|15|24|Et murmuravit populus contra Moysen dicens: " Quid bibemus? ".
EXOD|15|25|At ille clamavit ad Dominum, qui ostendit ei lignum; quod cum misisset in aquas, in dulcedinem versae sunt. Ibi constituit ei praecepta atque iudicia et ibi tentavit eum
EXOD|15|26|dicens: " Si audieris vocem Domini Dei tui et, quod rectum est coram eo, feceris et oboedieris mandatis eius custodierisque omnia praecepta illius, cunctum languorem, quem posui in Aegypto, non inducam super te: Ego enim Dominus sanator tuus ".
EXOD|15|27|Venerunt autem in Elim, ubi erant duodecim fontes aquarum et septuaginta palmae; et castrametati sunt iuxta aquas.
EXOD|16|1|Profectique sunt de Elim, et venit omnis congregatio filio rum Israel in desertum Sin, quod est inter Elim et Sinai, quinto decimo die mensis secundi postquam egressi sunt de terra Aegypti.
EXOD|16|2|Et murmuravit omnis congregatio filiorum Israel contra Moysen et Aaron in solitudine,
EXOD|16|3|dixeruntque filii Israel ad eos: " Utinam mortui essemus per manum Domini in terra Aegypti, quando sedebamus super ollas carnium et comedebamus panem in saturitate. Cur eduxistis nos in desertum istud, ut occideretis omnem coetum fame? ".
EXOD|16|4|Dixit autem Dominus ad Moysen: " Ecce ego pluam vobis panes de caelo; egrediatur populus et colligat, quae sufficiunt per singulos dies, ut tentem eum, utrum ambulet in lege mea an non.
EXOD|16|5|Die autem sexta parabunt quod intulerint, et duplum erit quam colligere solebant per singulos dies ".
EXOD|16|6|Dixeruntque Moyses et Aaron ad omnes filios Israel:" Vespere scietisquod Dominus eduxerit vosde terra Aegypti;
EXOD|16|7|et mane videbitisgloriam Domini.Audivit enim murmur vestrum contra Dominum. Nos vero quid sumus, quia mussitatis contra nos? ".
EXOD|16|8|Et ait Moyses:" Dabit Dominus vobisvespere carnes edereet mane panes in saturitate,eo quod audierit murmurationes vestras, quibus murmurati estis contra eum. Nos enim quid sumus? Nec contra nos est murmur vestrum, sed contra Dominum ".
EXOD|16|9|Dixitque Moyses ad Aaron: " Dic universae congregationi filiorum Israel: Accedite coram Domino; audivit enim murmur ve strum ".
EXOD|16|10|Cumque loqueretur Aaron ad omnem coetum filiorum Israel, respexerunt ad solitudinem, et ecce gloria Domini apparuit in nube.
EXOD|16|11|Locutus est autem Dominus ad Moysen dicens:
EXOD|16|12|" Audivi murmurationes filiorum Israel. Loquere ad eos: Vespere comedetis carnes et mane saturabimini panibus scietisque quod ego sum Dominus Deus vester ".
EXOD|16|13|Factum est ergo vespere, et ascendens coturnix operuit castra; mane quoque ros iacuit per circuitum castrorum.
EXOD|16|14|Cumque operuisset superficiem deserti, apparuit minutum et squamatum in similitudinem pruinae super terram.
EXOD|16|15|Quod cum vidissent filii Israel, dixerunt ad invicem: " Manhu? " (quod significat: " Quid est hoc? "). Ignorabant enim quid esset. Quibus ait Moyses: " Iste est panis, quem dedit Dominus vobis ad vescendum.
EXOD|16|16|Hic est sermo, quem praecepit Dominus: "Colligat ex eo unusquisque quantum sufficiat ad vescendum; gomor per singula capita iuxta numerum animarum vestrarum, quae habitant in tabernaculo, sic tolletis" ".
EXOD|16|17|Feceruntque ita filii Israel; et collegerunt alius plus, alius minus.
EXOD|16|18|Et mensi sunt ad mensuram gomor; nec qui plus collegerat, habuit amplius, nec qui minus paraverat, repperit minus, sed singuli, iuxta id quod edere poterant, congregaverunt.
EXOD|16|19|Dixitque Moyses ad eos: " Nullus relinquat ex eo in mane ".
EXOD|16|20|Qui non audierunt eum, sed dimiserunt quidam ex eis usque mane, et scatere coepit vermibus atque computruit; et iratus est contra eos Moyses.
EXOD|16|21|Colligebant autem mane singuli, quantum sufficere poterat ad vescendum; cumque incaluisset sol, liquefiebat.
EXOD|16|22|In die autem sexta collegerunt cibos duplices, id est duo gomor per singulos homines. Venerunt autem omnes principes congregationis et narraverunt Moysi.
EXOD|16|23|Qui ait eis: " Hoc est quod locutus est Dominus: Requies, sabbatum sanctum Domino cras; quodcumque torrendum est, torrete et, quae coquenda sunt, coquite; quidquid autem reliquum fuerit, reponite usque in mane ".
EXOD|16|24|Feceruntque ita, ut praeceperat Moyses, et non computruit, neque vermis inventus est in eo.
EXOD|16|25|Dixitque Moyses: " Comedite illud hodie, quia sabbatum est Domino; non invenietur hodie in agro.
EXOD|16|26|Sex diebus colligite; in die autem septimo sabbatum est Domino, idcirco non invenietur in eo ".
EXOD|16|27|Venitque septima dies; et egressi de populo, ut colligerent, non invenerunt.
EXOD|16|28|Dixit autem Dominus ad Moysen: " Usquequo non vultis custodire mandata mea et legem meam?
EXOD|16|29|Videte quod Dominus dederit vobis sabbatum et propter hoc die sexta tribuit vobis cibos duplices; maneat unusquisque apud semetipsum, nullus egrediatur de loco suo die septimo ".
EXOD|16|30|Et sabbatizavit populus die septimo.
EXOD|16|31|Appellavitque domus Israel nomen eius Man: quod erat quasi semen coriandri album, gustusque eius quasi similae cum melle.
EXOD|16|32|Dixit autem Moyses: " Iste est sermo, quem praecepit Dominus: "Imple gomor ex eo, et custodiatur in generationes vestras, ut noverint panem, quo alui vos in solitudine, quando educti estis de terra Aegypti" ".
EXOD|16|33|Dixitque Moyses ad Aaron: " Sume vas unum et mitte ibi man, quantum potest capere gomor; et repone coram Domino ad servandum in generationes vestras ".
EXOD|16|34|Sicut praecepit Dominus Moysi, posuit illud Aaron coram testimonio reservandum.
EXOD|16|35|Filii autem Israel comederunt man quadraginta annis, donec venirent in terram habitabilem; hoc cibo aliti sunt, usquequo tangerent fines terrae Chanaan.
EXOD|16|36|Gomor autem decima pars est ephi.
EXOD|17|1|Igitur profecta omnis congregatio filiorum Israel de deserto Sin per mansiones suas iuxta sermonem Domini, castrametati sunt in Raphidim, ubi non erat aqua ad bibendum populo.
EXOD|17|2|Qui iurgatus contra Moysen ait: " Da nobis aquam, ut bibamus ". Quibus respondit Moyses: " Quid iurgamini contra me? Cur tentatis Dominum? ".
EXOD|17|3|Sitivit ergo ibi populus prae aquae penuria et murmuravit contra Moysen dicens: " Cur fecisti nos exire de Aegypto, ut occideres nos et liberos nostros ac iumenta siti? ".
EXOD|17|4|Clamavit autem Moyses ad Dominum dicens: " Quid faciam populo huic? Adhuc paululum et lapidabunt me ".
EXOD|17|5|Et ait Dominus ad Moysen: " Antecede populum et sume tecum de senioribus Israel, et virgam, qua percussisti fluvium, tolle in manu tua et vade.
EXOD|17|6|En ego stabo coram te ibi super petram Horeb; percutiesque petram, et exibit ex ea aqua, ut bibat populus ". Fecit Moyses ita coram senioribus Israel.
EXOD|17|7|Et vocavit nomen loci illius Massa et Meriba, propter iurgium filiorum Israel et quia tentaverunt Dominum dicentes: " Estne Dominus in nobis an non? ".
EXOD|17|8|Venit autem Amalec et pugnabat contra Israel in Raphidim.
EXOD|17|9|Dixitque Moyses ad Iosue: " Elige nobis viros et egressus pugna contra Amalec; cras ego stabo in vertice collis habens virgam Dei in manu mea ".
EXOD|17|10|Fecit Iosue, ut locutus erat ei Moyses, et pugnavit contra Amalec; Moyses autem et Aaron et Hur ascenderunt super verticem collis.
EXOD|17|11|Cumque levaret Moyses manus, vincebat Israel; sin autem remisisset, superabat Amalec.
EXOD|17|12|Manus autem Moysi erant graves; sumentes igitur lapidem posuerunt subter eum, in quo sedit; Aaron autem et Hur sustentabant manus eius ex utraque parte. Et factum est ut manus eius non lassarentur usque ad occasum solis.
EXOD|17|13|Vicitque Iosue Amalec et populum eius in ore gladii.
EXOD|17|14|Dixit autem Dominus ad Moysen: " Scribe hoc ob monumentum in libro et trade auribus Iosue; delebo enim memoriam Amalec sub caelo ".
EXOD|17|15|Aedificavitque Moyses altare et vocavit nomen eius Dominus Nissi "Dominus vexillum meum)
EXOD|17|16|dicens:" Quia manus contra solium Domini:bellum Domino erit contra Amalec a generatione in generationem ".
EXOD|18|1|Cumque audisset Iethro sacerdos Madian socer Moysi omnia, quae fecerat Deus Moysi et Israel populo suo, eo quod eduxisset Dominus Israel de Aegypto,
EXOD|18|2|tulit Sephoram uxorem Moysi, quam remiserat,
EXOD|18|3|et duos filios eius, quorum unus vocabatur Gersam, dicente patre: " Advena fui in terra aliena ",
EXOD|18|4|alter vero Eliezer: " Deus enim, ait, patris mei adiutor meus, et eruit me de gladio pharaonis ".
EXOD|18|5|Venit ergo Iethro socer Moysi et filii eius et uxor eius ad Moysen in desertum, ubi erat castrametatus iuxta montem Dei;
EXOD|18|6|et mandavit Moysi dicens: " Ego socer tuus Iethro venio ad te et uxor tua et duo filii tui cum ea ".
EXOD|18|7|Qui egressus in occursum soceri sui adoravit et osculatus est eum, salutaveruntque se mutuo verbis pacificis. Cumque intrasset tabernaculum,
EXOD|18|8|narravit Moyses socero suo cuncta, quae fecerat Dominus pharaoni et Aegyptiis propter Israel, universumque laborem, qui accidisset eis in itinere, et quod liberaverat eos Dominus.
EXOD|18|9|Laetatusque est Iethro super omnibus bonis, quae fecerat Dominus Israel, eo quod eruisset eum de manu Aegyptiorum,
EXOD|18|10|et ait: " Benedictus Dominus, qui liberavit vos de manu Aegyptiorum et de manu pharaonis.
EXOD|18|11|Nunc cognovi quia magnus Dominus super omnes deos, eo quod eruerit populum de manu Aegyptiorum, qui superbe egerunt contra illos ".
EXOD|18|12|Obtulit ergo Iethro socer Moysi holocausta et hostias Deo; veneruntque Aaron et omnes seniores Israel, ut comederent panem cum eo coram Deo.
EXOD|18|13|Altero autem die sedit Moyses, ut iudicaret populum, qui assistebat Moysi de mane usque ad vesperam.
EXOD|18|14|Quod cum vidisset socer eius, omnia scilicet, quae agebat in populo, ait: " Quid est hoc, quod facis in plebe? Cur solus sedes, et omnis populus praestolatur de mane usque ad vesperam? ".
EXOD|18|15|Cui respondit Moyses: " Venit ad me populus quaerens sententiam Dei.
EXOD|18|16|Cumque acciderit eis aliqua disceptatio, veniunt ad me, ut iudicem inter eos et ostendam praecepta Dei et leges eius ".
EXOD|18|17|At ille: " Non bonam, inquit, rem facis.
EXOD|18|18|Consumeris et tu et populus iste, qui tecum est. Ultra vires tuas est negotium; solus illud non poteris sustinere.
EXOD|18|19|Sed audi verba mea atque consilia, et erit Deus tecum: Esto tu populo in his, quae ad Deum pertinent, ut referas causas ad Deum
EXOD|18|20|ostendasque populo praecepta et leges viamque, per quam ingredi debeant, et opus, quod facere debeant.
EXOD|18|21|Provide autem de omni plebe viros strenuos et timentes Deum, in quibus sit veritas, et qui oderint avaritiam, et constitue ex eis tribunos et centuriones et quinquagenarios et decanos,
EXOD|18|22|qui iudicent populum omni tempore. Quidquid autem maius fuerit, referant ad te, et ipsi minora tantummodo iudicent; leviusque sit tibi, partito cum aliis onere.
EXOD|18|23|Si hoc feceris, implebis imperium Dei et praecepta eius poteris sustentare, et omnis hic populus revertetur ad loca sua cum pace ".
EXOD|18|24|Quibus auditis, Moyses fecit omnia, quae ille suggesserat;
EXOD|18|25|et, electis viris strenuis de cuncto Israel, constituit eos principes populi, tribunos et centuriones et quinquagenarios et decanos,
EXOD|18|26|qui iudicabant plebem omni tempore. Quidquid autem gravius erat, referebant ad eum, faciliora tantummodo iudicantes.
EXOD|18|27|Dimisitque socerum suum, qui reversus abiit in terram suam.
EXOD|19|1|Mense tertio egressionis Israel de terra Aegypti, in die hac venerunt in solitudinem Sinai.
EXOD|19|2|Nam profecti de Raphidim et pervenientes usque in desertum Sinai, castrametati sunt in eodem loco,ibique Israel fixit tentoria e regione montis.
EXOD|19|3|Moyses autem ascendit ad Deum, vocavitque eum Dominus de monte et ait:" Haec dices domui Iacobet annuntiabis filiis Israel:
EXOD|19|4|Vos ipsi vidistis, quae fecerim Aegyptiis,quomodo portaverim vos super alas aquilarumet adduxerim ad me.
EXOD|19|5|Si ergo audieritis vocem meamet custodieritis pactum meum,eritis mihi in peculium de cunctis populis;mea est enim omnis terra.
EXOD|19|6|Et vos eritis mihi regnum sacerdotumet gens sancta.Haec sunt verba, quae loqueris ad filios Israel ".
EXOD|19|7|Venit Moyses et, convocatis maioribus natu populi, exposuit omnes sermones, quos mandaverat Dominus.
EXOD|19|8|Responditque universus populus simul: " Cuncta, quae locutus est Dominus, faciemus ". Cumque rettulisset Moyses verba populi ad Dominum,
EXOD|19|9|ait ei Dominus: " Ecce ego veniam ad te in caligine nubis, ut audiat me populus loquentem ad te et tibi quoque credat in perpetuum ".Nuntiavit ergo Moyses verba populi ad Dominum,
EXOD|19|10|qui dixit ei: " Vade ad populum et sanctifica illos hodie et cras; laventque vestimenta sua
EXOD|19|11|et sint parati in diem tertium. In die enim tertio descendet Dominus coram omni plebe super montem Sinai.
EXOD|19|12|Constituesque terminos populo per circuitum et dices: Cavete, ne ascendatis in montem nec tangatis fines illius; omnis, qui tetigerit montem, morte morietur.
EXOD|19|13|Manus non tanget eum, sed lapidibus opprimetur aut confodietur iaculis; sive iumentum fuerit, sive homo, non vivet. Cum coeperit clangere bucina, tunc ascendant in montem ".
EXOD|19|14|Descenditque Moyses de monte ad populum et sanctificavit eum; cumque lavissent vestimenta sua,
EXOD|19|15|ait ad eos: " Estote parati in diem tertium; ne appropinquetis uxoribus vestris ".
EXOD|19|16|Iamque advenerat tertius dies, et mane inclaruerat; et ecce coeperunt audiri tonitrua ac micare fulgura et nubes densissima operire montem, clangorque bucinae vehementius perstrepebat; et timuit populus, qui erat in castris.
EXOD|19|17|Cumque eduxisset eos Moyses in occursum Dei de loco castrorum, steterunt ad radices montis.
EXOD|19|18|Totus autem mons Sinai fumabat, eo quod descendisset Dominus super eum in igne, et ascenderet fumus ex eo quasi de fornace. Et tremuit omnis mons vehementer.
EXOD|19|19|Et sonitus bucinae paulatim crescebat in maius; Moyses loquebatur, et Deus respondebat ei cum voce.
EXOD|19|20|Descenditque Dominus super montem Sinai in ipso montis vertice et vocavit Moysen in cacumen eius. Quo cum ascendisset,
EXOD|19|21|dixit ad eum: " Descende et contestare populum, ne velit transcendere terminos ad videndum Dominum, et pereat ex eis plurima multitudo.
EXOD|19|22|Sacerdotes quoque, qui accedunt ad Dominum, sanctificentur, ne percutiat eos ".
EXOD|19|23|Dixitque Moyses ad Dominum: " Non poterit vulgus ascendere in montem Sinai, tu enim testificatus es et iussisti dicens: "Pone terminos circa montem et sanctifica illum" ".
EXOD|19|24|Cui ait Dominus: " Vade, descende; ascendesque tu et Aaron tecum, sacerdotes autem et populus ne transeant terminos nec ascendant ad Dominum, ne interficiat illos ".
EXOD|19|25|Descenditque Moyses ad populum et omnia narravit eis.
EXOD|20|1|Locutusque est Deus cunctos sermones hos:
EXOD|20|2|" Ego sum Dominus Deus tuus, qui eduxi te de terra Aegypti, de domo servitutis.
EXOD|20|3|Non habebis deos alienos coram me.
EXOD|20|4|Non facies tibi sculptile neque omnem similitudinem eorum, quae sunt in caelo desuper et quae in terra deorsum et quae in aquis sub terra.
EXOD|20|5|Non adorabis ea neque coles, quia ego sum Dominus Deus tuus, Deus zelotes, visitans iniquitatem patrum in filiis in tertiam et quartam generationem eorum, qui oderunt me,
EXOD|20|6|et faciens misericordiam in milia his, qui diligunt me et custodiunt praecepta mea.
EXOD|20|7|Non assumes nomen Domini Dei tui in vanum, nec enim habebit insontem Dominus eum, qui assumpserit nomen Domini Dei sui frustra.
EXOD|20|8|Memento, ut diem sabbati sanctifices.
EXOD|20|9|Sex diebus operaberis et facies omnia opera tua;
EXOD|20|10|septimus autem dies sabbatum Domino Deo tuo est; non facies omne opus tu et filius tuus et filia tua, servus tuus et ancilla tua, iumentum tuum et advena, qui est intra portas tuas.
EXOD|20|11|Sex enim diebus fecit Dominus caelum et terram et mare et omnia, quae in eis sunt, et requievit in die septimo; idcirco benedixit Dominus diei sabbati et sanctificavit eum.
EXOD|20|12|Honora patrem tuum et matrem tuam, ut sis longaevus super terram, quam Dominus Deus tuus dabit tibi.
EXOD|20|13|Non occides.
EXOD|20|14|Non moechaberis.
EXOD|20|15|Non furtum facies.
EXOD|20|16|Non loqueris contra proximum tuum falsum testimonium.
EXOD|20|17|Non concupisces domum proximi tui: non desiderabis uxorem eius, non servum, non ancillam, non bovem, non asinum nec omnia, quae illius sunt ".
EXOD|20|18|Cunctus autem populus videbat voces et lampades et sonitum bucinae montemque fumantem; et perterriti ac pavore concussi steterunt procul
EXOD|20|19|dicentes Moysi: " Loquere tu nobis, et audiemus; non loquatur nobis Deus, ne moriamur ".
EXOD|20|20|Et ait Moyses ad populum: " Nolite timere; ut enim probaret vos, venit Deus, et ut timor illius esset in vobis, ne peccaretis ".
EXOD|20|21|Stetitque populus de longe; Moyses autem accessit ad caliginem, in qua erat Deus.
EXOD|20|22|Dixit praeterea Dominus ad Moysen: " Haec dices filiis Israel: Vos vidistis quod de caelo locutus sim vobis.
EXOD|20|23|Non facietis praeter me deos argenteos nec deos aureos facietis vobis.
EXOD|20|24|Altare de terra facietis mihi et offeretis super eo holocausta et pacifica vestra, oves vestras et boves; in omni loco, in quo memoriam fecero nominis mei, veniam ad te et benedicam tibi.
EXOD|20|25|Quod si altare lapideum feceris mihi, non aedificabis illud de sectis lapidibus; si enim levaveris cultrum super eo, polluetur.
EXOD|20|26|Non ascendes per gradus ad altare meum, ne reveletur turpitudo tua.
EXOD|21|1|Haec sunt iudicia, quae propones eis:
EXOD|21|2|Si emeris servum Hebraeum, sex annis serviet tibi; in septimo egredietur liber gratis.
EXOD|21|3|Si solus intraverit, solus exeat; si habens uxorem, et uxor egredietur simul.
EXOD|21|4|Sin autem dominus dederit illi uxorem, et pepererit filios et filias, mulier et liberi eius erunt domini sui; ipse vero exibit solus.
EXOD|21|5|Quod si dixerit servus: "Diligo dominum meum et uxorem ac liberos, non egrediar liber",
EXOD|21|6|afferet eum dominus ad Deum et applicabit eum ad ostium vel postes perforabitque aurem eius subula; et erit ei servus in saeculum.
EXOD|21|7|Si quis vendiderit filiam suam in famulam, non egredietur sicut servi exire consueverunt.
EXOD|21|8|Si displicuerit oculis domini sui, cui tradita fuerat, faciat eam redimi; populo autem alieno vendendi non habebit potestatem, quia fraudavit eam.
EXOD|21|9|Sin autem filio suo desponderit eam, iuxta morem filiarum faciet illi.
EXOD|21|10|Quod si alteram sibi acceperit, cibum et vestimentum et concubitum non negabit.
EXOD|21|11|Si tria ista non fecerit ei, egredietur gratis absque pretio.
EXOD|21|12|Qui percusserit hominem, et ille mortuus fuerit, morte moriatur.
EXOD|21|13|Qui autem non est insidiatus, sed Deus illum tradidit in manus eius, constituam tibi locum, in quem fugere debeat.
EXOD|21|14|Si quis de industria occiderit proximum suum et per insidias, ab altari meo evelles eum, ut moriatur.
EXOD|21|15|Qui percusserit patrem suum aut matrem, morte moriatur.
EXOD|21|16|Qui furatus fuerit hominem sive vendiderit eum sive inventus fuerit in manu eius, morte moriatur.
EXOD|21|17|Qui maledixerit patri suo vel matri, morte moriatur.
EXOD|21|18|Si rixati fuerint viri, et percusserit alter proximum suum lapide vel pugno, et ille mortuus non fuerit, sed iacuerit in lectulo,
EXOD|21|19|si surrexerit et ambulaverit foris super baculum suum, impunitus erit, qui percusserit, ita tamen, ut operas eius deperditas et impensas pro medela restituat.
EXOD|21|20|Qui percusserit servum suum vel ancillam virga, et mortui fuerint in manibus eius, ultioni subiacetur.
EXOD|21|21|Sin autem uno die vel duobus supervixerit, non subiacebit poenae, quia pecunia illius est.
EXOD|21|22|Si rixati fuerint viri, et percusserit quis mulierem praegnantem et abortivum quidem fecerit, sed aliud quid adversi non acciderit, subiacebit damno, quantum maritus mulieris expetierit, et arbitri iudicaverint.
EXOD|21|23|Sin autem quid adversi acciderit, reddet animam pro anima,
EXOD|21|24|oculum pro oculo, dentem pro dente, manum pro manu, pedem pro pede,
EXOD|21|25|adustionem pro adustione, vulnus pro vulnere, livorem pro livore.
EXOD|21|26|Si percusserit quispiam oculum servi sui aut ancillae et luscos eos fecerit, dimittet eos liberos pro oculo.
EXOD|21|27|Dentem quoque si excusserit servo vel ancillae suae, dimittet eos liberos pro dente.
EXOD|21|28|Si bos cornu percusserit virum aut mulierem, et mortui fuerint, lapidibus obruetur, et non comedentur carnes eius; dominus autem bovis innocens erit.
EXOD|21|29|Quod si bos cornupeta fuerit ab heri et nudiustertius, et contestati sunt dominum eius, nec recluserit eum, occideritque virum aut mulierem: et bos lapidibus obruetur, et dominum illius occident.
EXOD|21|30|Quod si pretium ei fuerit impositum, dabit pro anima sua, quidquid fuerit postulatus.
EXOD|21|31|Filium quoque vel filiam si cornu percusserit, simili sententiae subiacebit.
EXOD|21|32|Si servum vel ancillam invaserit, triginta siclos argenti dabit domino; bos vero lapidibus opprimetur.
EXOD|21|33|Si quis aperuerit cisternam vel foderit et non operuerit eam, cedideritque bos vel asinus in eam,
EXOD|21|34|dominus cisternae reddet pretium iumentorum; quod autem mortuum est, ipsius erit.
EXOD|21|35|Si bos alienus bovem alterius vulneraverit, et ille mortuus fuerit, vendent bovem vivum et divident pretium; cadaver autem mortui inter se dispertient.
EXOD|21|36|Sin autem notum erat quod bos cornupeta esset ab heri et nudiustertius, et non custodivit eum dominus suus, reddet bovem pro bove et cadaver integrum accipiet.
EXOD|21|37|Si quis furatus fuerit bovem aut ovem et occiderit vel vendiderit, quinque boves pro uno bove restituet et quattuor oves pro una ove.
EXOD|22|1|Si effringens fur domum sive suffodiens fuerit inventus et, accepto vulnere, mortuus fuerit, percussor non erit reus sanguinis.
EXOD|22|2|Quod si orto sole hoc fecerit, erit reus sanguinis. Fur plene restituet. Si non habuerit, quod reddat, venumdabitur pro furto.
EXOD|22|3|Si inventum fuerit apud eum, quod furatus est, vivens sive bos sive asinus sive ovis, duplum restituet.
EXOD|22|4|Si quispiam depasci permiserit agrum vel vineam et dimiserit iumentum suum, ut depascatur agrum alienum, restituet plene ex agro suo secundum fruges eius; si autem totum agrum depastum fuerit, quidquid optimum habuerit in agro suo vel in vinea, restituet.
EXOD|22|5|Si egressus ignis invenerit spinas et comprehenderit acervos frugum sive stantes segetes sive agrum, reddet damnum, qui ignem succenderit.
EXOD|22|6|Si quis commendaverit amico pecuniam aut vasa in custodiam, et ab eo, qui susceperat, furto ablata fuerint, si invenitur fur, duplum reddet.
EXOD|22|7|Si latet fur, dominus domus applicabitur ad Deum et iurabit quod non extenderit manum in rem proximi sui.
EXOD|22|8|In omni causa fraudis tam de bove quam de asino et ove ac vestimento et, quidquid damnum inferre potest, si quis dixerit: " Hoc est! ", ad Deum utriusque causa perveniet, et, quem Deus condemnaverit, duplum restituet proximo suo.
EXOD|22|9|Si quis commendaverit proximo suo asinum, bovem, ovem vel omne iumentum ad custodiam, et mortuum fuerit aut fractum vel captum ab hostibus, nullusque hoc viderit,
EXOD|22|10|iusiurandum per Dominum erit in medio quod non extenderit manum ad rem proximi sui; suscipietque dominus iuramentum, et ille reddere non cogetur.
EXOD|22|11|Quod si furto ablatum fuerit, restituet damnum domino;
EXOD|22|12|si dilaceratum a bestia, deferat, quod occisum est, in testimonium et non restituet.
EXOD|22|13|Qui a proximo suo quidquam horum mutuo postulaverit, et fractum aut mortuum fuerit, domino non praesente, reddere compelletur.
EXOD|22|14|Quod si impraesentiarum dominus fuerit, non restituet. Si mercennarius est, venit in mercedem operis sui.
EXOD|22|15|Si seduxerit quis virginem necdum desponsatam dormieritque cum ea, pretio acquiret eam sibi uxorem.
EXOD|22|16|Si pater virginis eam dare noluerit, appendet ei pecuniam iuxta pretium pro virginibus dandum.
EXOD|22|17|Maleficam non patieris vivere.
EXOD|22|18|Qui coierit cum iumento, morte moriatur.
EXOD|22|19|Qui immolat diis, occidetur, praeter Domino soli.
EXOD|22|20|Advenam non opprimes neque affliges eum; advenae enim et ipsi fuistis in terra Aegypti.
EXOD|22|21|Viduae et pupillo non nocebitis.
EXOD|22|22|Si laeseritis eos, vociferabuntur ad me, et ego audiam clamorem eorum;
EXOD|22|23|et indignabitur furor meus, percutiamque vos gladio, et erunt uxores vestrae viduae et filii vestri pupilli.
EXOD|22|24|Si pecuniam mutuam dederis in populo meo pauperi, qui habitat tecum, non eris ei quasi creditor; non imponetis ei usuram.
EXOD|22|25|Si pignus a proximo tuo acceperis pallium, ante solis occasum reddes ei;
EXOD|22|26|ipsum enim est solum, quo operitur, indumentum carnis eius, nec habet aliud, in quo dormiat; si clamaverit ad me, exaudiam eum, quia misericors sum.
EXOD|22|27|Deo non detrahes et principi populi tui non maledices.
EXOD|22|28|Abundantiam areae tuae et torcularis tui non tardabis reddere.Primogenitum filiorum tuorum dabis mihi.
EXOD|22|29|De bobus quoque et ovibus similiter facies: septem diebus sit cum matre sua, die octavo reddes illum mihi.
EXOD|22|30|Viri sancti eritis mihi; carnem animalis in agro dilacerati non comedetis, sed proicietis canibus.
EXOD|23|1|Non suscipies famam falsam nec iunges manum tuam cum impio, ut dicas falsum testimonium.
EXOD|23|2|Non sequeris turbam ad faciendum malum; nec in iudicio plurimorum acquiesces sententiae, ut a vero devies.
EXOD|23|3|Pauperis quoque non misereberis in iudicio.
EXOD|23|4|Si occurreris bovi inimici tui aut asino erranti, reduc ad eum.
EXOD|23|5|Si videris asinum odientis te iacere sub onere suo, non pertransibis, sed sublevabis cum eo.
EXOD|23|6|Non pervertes iudicium pauperis in lite eius.
EXOD|23|7|Mendacium fugies. Insontem et iustum non occides, quia aversor impium.
EXOD|23|8|Nec accipies munera, quae excaecant etiam prudentes et subvertunt verba iustorum.
EXOD|23|9|Peregrinum non opprimes; scitis enim advenarum animas, quia et ipsi peregrini fuistis in terra Aegypti.
EXOD|23|10|Sex annis seminabis terram tuam et congregabis fruges eius.
EXOD|23|11|Anno autem septimo dimittes eam et requiescere facies, ut comedant pauperes populi tui; et quidquid reliquum fuerit, edant bestiae agri. Ita facies in vinea et in oliveto tuo.
EXOD|23|12|Sex diebus operaberis; septima die cessabis, ut requiescat bos et asinus tuus, et refrigeretur filius ancillae tuae et advena.
EXOD|23|13|Omnia, quae dixi vobis, custodite, et nomen externorum deorum non invocabitis, neque audietur ex ore tuo.
EXOD|23|14|Tribus vicibus per singulos annos mihi festa celebrabitis.
EXOD|23|15|Sollemnitatem Azymorum custodies: septem diebus comedes azyma, sicut praecepi tibi, tempore statuto mensis Abib, quando egressus es de Aegypto.Non apparebis in conspectu meo vacuus.
EXOD|23|16|Et sollemnitatem Messis primitivorum operis tui, quaecumque seminaveris in agro; sollemnitatem quoque Collectae in exitu anni, quando congregaveris omnes fruges tuas de agro.
EXOD|23|17|Ter in anno apparebit omne masculinum tuum coram Domino Deo.
EXOD|23|18|Non immolabis super fermento sanguinem victimae meae, nec remanebit adeps sollemnitatis meae usque mane.
EXOD|23|19|Primitias primarum frugum terrae tuae deferes in domum Domini Dei tui.Non coques haedum in lacte matris suae.
EXOD|23|20|Ecce ego mittam angelum, qui praecedat te et custodiat in via et introducat ad locum, quem paravi.
EXOD|23|21|Observa eum et audi vocem eius nec contemnendum putes; quia non dimittet, cum peccaveritis, quia est nomen meum in illo.
EXOD|23|22|Quod si audieris vocem eius et feceris omnia, quae loquor, inimicus ero inimicis tuis et affligam affligentes te.
EXOD|23|23|Praecedet enim te angelus meus et introducet te ad Amorraeum et Hetthaeum et Pherezaeum Chananaeumque et Hevaeum et Iebusaeum, quos ego conteram.
EXOD|23|24|Non adorabis deos eorum nec coles eos; non facies secundum opera eorum, sed destrues eos et confringes lapides eorum.
EXOD|23|25|Servietisque Domino Deo vestro, ut benedicam panibus tuis et aquis et auferam infirmitatem de medio tui.
EXOD|23|26|Non erit abortiens nec sterilis in terra tua; numerum dierum tuorum implebo.
EXOD|23|27|Terrorem meum mittam in praecursum tuum et perturbabo omnem populum, ad quem ingre dieris; cunctorumque inimicorum tuorum coram te terga vertam
EXOD|23|28|emittens crabrones prius, qui fugabunt Hevaeum et Chananaeum et Hetthaeum, antequam introeas.
EXOD|23|29|Non eiciam eos a facie tua anno uno, ne terra in solitudinem redigatur, et multiplicentur contra te bestiae agri.
EXOD|23|30|Paulatim expellam eos de conspectu tuo, donec augearis et possideas terram.
EXOD|23|31|Ponam autem terminos tuos a mari Rubro usque ad mare Palaestinorum et a deserto usque ad Fluvium. Tradam manibus vestris habitatores terrae et eiciam eos de conspectu vestro.
EXOD|23|32|Non inibis cum eis foedus nec cum diis eorum.
EXOD|23|33|Non habitent in terra tua, ne peccare te faciant in me, si servieris diis eorum; quod tibi certo erit in scandalum ".
EXOD|24|1|Moysi quoque dixit: " Ascende ad Dominum, tu et Aa ron, Nadab et Abiu et septuaginta senes ex Israel, et adorabitis procul.
EXOD|24|2|Solusque Moyses ascendet ad Dominum, et illi non appropinquabunt, nec populus ascendet cum eo ".
EXOD|24|3|Venit ergo Moyses et narravit plebi omnia verba Domini atque iudicia; responditque omnis populus una voce: " Omnia verba Domini, quae locutus est, faciemus ".
EXOD|24|4|Scripsit autem Moyses universos sermones Domini; et mane consurgens aedificavit altare ad radices montis et duodecim lapides per duodecim tribus Israel.
EXOD|24|5|Misitque iuvenes de filiis Israel, et obtulerunt holocausta; immolaveruntque victimas pacificas Domino vitulos.
EXOD|24|6|Tulit itaque Moyses dimidiam partem sanguinis et misit in crateras; partem autem residuam respersit super altare.
EXOD|24|7|Assumensque volumen foederis legit, audiente populo, qui dixerunt: " Omnia, quae locutus est Dominus, faciemus et erimus oboedientes ".
EXOD|24|8|Ille vero sumptum sanguinem respersit in populum et ait: " Hic est sanguis foederis, quod pepigit Dominus vobiscum super cunctis sermonibus his ".
EXOD|24|9|Ascenderuntque Moyses et Aaron, Nadab et Abiu et septuaginta de senioribus Israel.
EXOD|24|10|Et viderunt Deum Israel, et sub pedibus eius quasi opus lapidis sapphirini et quasi ipsum caelum, cum serenum est.
EXOD|24|11|Nec in electos filiorum Israel misit manum suam; videruntque Deum et comederunt ac biberunt.
EXOD|24|12|Dixit autem Dominus ad Moysen: " Ascende ad me in montem et esto ibi; daboque tibi tabulas lapideas et legem ac mandata, quae scripsi, ut doceas eos ".
EXOD|24|13|Surrexerunt Moyses et Iosue minister eius; ascendensque Moyses in montem Dei
EXOD|24|14|senioribus ait: " Exspectate hic, donec revertamur ad vos. Habetis Aaron et Hur vobiscum; si quid natum fuerit quaestionis, referetis ad eos ".
EXOD|24|15|Cumque ascendisset Moyses in montem, operuit nubes montem;
EXOD|24|16|et habitavit gloria Domini super Sinai tegens illum nube sex diebus; septimo autem die vocavit eum de medio caliginis.
EXOD|24|17|Erat autem species gloriae Domini quasi ignis ardens super verticem montis in conspectu filiorum Israel.
EXOD|24|18|Ingressusque Moyses medium nebulae ascendit in montem; et fuit ibi quadraginta diebus et quadraginta noctibus.
EXOD|25|1|Locutusque est Dominus ad Moysen dicens:
EXOD|25|2|" Loquere filiis Israel, ut tollant mihi donaria; ab omni homine, qui offert ultroneus, accipietis ea.
EXOD|25|3|Haec sunt autem, quae accipere debetis: aurum et argentum et aes,
EXOD|25|4|hyacinthum et purpuram coccumque et byssum, pilos caprarum
EXOD|25|5|et pelles arietum rubricatas pellesque delphini et ligna acaciae,
EXOD|25|6|oleum ad luminaria concinnanda, aromata in unguentum et in thymiama boni odoris,
EXOD|25|7|lapides onychinos et gemmas ad ornandum ephod ac pectorale.
EXOD|25|8|Facientque mihi sanctuarium, et habitabo in medio eorum.
EXOD|25|9|Iuxta omnem similitudinem habitaculi, quam ostendam tibi, et omnium vasorum in cultum eius: sicque facietis illud.
EXOD|25|10|Arcam de lignis acaciae compingent; cuius longitudo habeat duos semis cubitos, latitudo cubitum et dimidium, altitudo cubitum similiter ac semissem.
EXOD|25|11|Et deaurabis eam auro mundissimo intus et foris; faciesque supra coronam auream per circuitum
EXOD|25|12|et conflabis ei quattuor circulos aureos, quos pones in quattuor arcae pedibus: duo circuli sint in latere uno et duo in altero.
EXOD|25|13|Facies quoque vectes de lignis acaciae et operies eos auro;
EXOD|25|14|inducesque per circulos, qui sunt in arcae lateribus, ut portetur in eis;
EXOD|25|15|qui semper erunt in circulis nec umquam extrahentur ab eis.
EXOD|25|16|Ponesque in arcam testimonium, quod dabo tibi.
EXOD|25|17|Facies et propitiatorium de auro mundissimo; duos cubitos et dimidium tenebit longitudo eius, et cubitum ac semissem latitudo.
EXOD|25|18|Duos quoque cherubim aureos et productiles facies ex utraque parte propitiatorii,
EXOD|25|19|cherub unus sit in latere uno et alter in altero; ex propitiatorio facies cherubim in utraque parte eius.
EXOD|25|20|Expandent alas sursum et operient alis suis propitiatorium; respicientque se mutuo, versis vultibus in propitiatorium,
EXOD|25|21|quo operienda est arca, in qua pones testimonium, quod dabo tibi.
EXOD|25|22|Et conveniam te ibi et loquar ad te supra propitiatorium de medio duorum cherubim, qui erunt super arcam testimonii, cuncta, quae mandabo per te filiis Israel.
EXOD|25|23|Facies et mensam de lignis acaciae habentem duos cubitos longitudinis et in latitudine cubitum et in altitudine cubitum ac semissem.
EXOD|25|24|Et inaurabis eam auro purissimo; faciesque illi coronam auream per circuitum.
EXOD|25|25|Facies quoque ei limbum altum quattuor digitis per circuitum et super illum coronam auream.
EXOD|25|26|Quattuor quoque circulos aureos praeparabis et pones eos in quattuor angulis eiusdem mensae per singulos pedes.
EXOD|25|27|Iuxta limbum erunt circuli aurei, ut mittantur vectes per eos, et possit mensa portari.
EXOD|25|28|Ipsosque vectes facies de lignis acaciae et circumdabis auro, et per ipsos subvehitur mensa.
EXOD|25|29|Parabis et acetabula ac phialas, vasa et cyathos, in quibus offerenda sunt libamina, ex auro purissimo.
EXOD|25|30|Et pones super mensam panes propositionis in conspectu meo semper.
EXOD|25|31|Facies et candelabrum ductile de auro mundissimo: basis et hastile eius, scyphi et sphaerulae ac flores in unum efformentur.
EXOD|25|32|Sex calami egredientur de lateribus, tres ex uno latere et tres ex altero.
EXOD|25|33|Tres scyphi quasi in nucis modum in calamo uno sphaerulaeque simul et flores; et tres similiter scyphi instar nucis in calamo altero sphaerulaeque simul et flores: hoc erit opus sex calamorum, qui producendi sunt de hastili.
EXOD|25|34|In ipso autem hastili candelabri erunt quattuor scyphi in nucis modum sphaerulaeque et flores.
EXOD|25|35|Singulae sphaerulae sub binis calamis per tria loca, qui simul sex fiunt, procedentes de hastili uno.
EXOD|25|36|Sphaerulae igitur et calami unum cum ipso erunt, totum ductile de auro purissimo.
EXOD|25|37|Facies et lucernas septem et pones eas super candelabrum, ut luceant in locum ex adverso.
EXOD|25|38|Emunctoria quoque et vasa, in quibus emuncta condantur, fient de auro purissimo.
EXOD|25|39|Omne pondus candelabri cum universis vasis suis habebit talentum auri purissimi.
EXOD|25|40|Inspice et fac secundum exemplar, quod tibi in monte monstratum est.
EXOD|26|1|Habitaculum vero ita facies: decem cortinas de bysso re torta et hyacintho ac purpura coccoque cum cherubim opere polymito facies.
EXOD|26|2|Longitudo cortinae unius habebit viginti octo cubitos, latitudo quattuor cubitorum erit. Unius mensurae fient universae cortinae.
EXOD|26|3|Quinque cortinae sibi iungentur mutuo, et aliae quinque nexu simili cohaerebunt.
EXOD|26|4|Ansulas hyacinthinas in latere facies cortinae unius in extremitate iuncturae et similiter facies in latere cortinae extremae in iunctura altera.
EXOD|26|5|Quinquaginta ansulas facies in cortina una et quinquaginta ansulas facies in summitate cortinae, quae est in iunctura altera, ita insertas, ut ansa contra ansam veniat.
EXOD|26|6|Facies et quinquaginta fibulas aureas, quibus cortinarum vela iungenda sunt, ut unum habitaculum fiat.
EXOD|26|7|Facies et saga cilicina undecim pro tabernaculo super habitaculum.
EXOD|26|8|Longitudo sagi unius habebit triginta cubitos et latitudo quattuor; aequa erit mensura sagorum omnium.
EXOD|26|9|E quibus quinque iunges seorsum et sex sibi mutuo copulabis, ita ut sextum sagum in fronte tecti duplices.
EXOD|26|10|Facies et quinquaginta ansas in ora sagi ultimi iuncturae unius et quinquaginta ansas in ora sagi iuncturae alterius.
EXOD|26|11|Facies et quinquaginta fibulas aeneas, quibus iungantur ansae, ut unum ex omnibus tabernaculum fiat.
EXOD|26|12|Quod autem superfuerit in sagis, quae parantur tecto, id est unum sagum, quod amplius est, ex medietate eius operies posteriora habitaculi;
EXOD|26|13|et cubitus ex una parte pendebit, et alter ex altera, qui plus est in longitudine sagorum tabernaculi utrumque latus habitaculi protegens.
EXOD|26|14|Facies et operimentum aliud pro tabernaculo de pellibus arietum rubricatis et super hoc rursum aliud operimentum de pellibus delphini.
EXOD|26|15|Facies et tabulas stantes habitaculi de lignis acaciae,
EXOD|26|16|quae singulae denos cubitos in longitudine habeant et in latitudine singulos ac semissem.
EXOD|26|17|In tabula una duo pedes fient, quibus tabula alteri tabulae conectatur; atque in hunc modum cunctae tabulae habitaculi parabuntur.
EXOD|26|18|Quarum viginti erunt in latere meridiano, quod vergit ad austrum;
EXOD|26|19|quibus quadraginta bases argenteas fundes, ut binae bases singulis pedibus singularum tabularum subiciantur.
EXOD|26|20|In latere quoque secundo habitaculi, quod vergit ad aquilonem, viginti tabulae erunt,
EXOD|26|21|quadraginta habentes bases argenteas; binae bases singulis tabulis supponentur.
EXOD|26|22|Ad occidentalem vero plagam in tergo habitaculi facies sex tabulas;
EXOD|26|23|et rursum alias duas, quae in angulis erigantur, post tergum habitaculi.
EXOD|26|24|Eruntque geminae a deorsum usque sursum in compaginem unam; ita erit duabus istis, pro duabus angulis erunt.
EXOD|26|25|Et erunt simul tabulae octo, bases earum argenteae sedecim, duabus basibus per unam tabulam supputatis.
EXOD|26|26|Facies et vectes de lignis acaciae, quinque ad continendas tabulas in uno latere habitaculi
EXOD|26|27|et quinque alios in altero et eiusdem numeri in tergo ad occidentalem plagam;
EXOD|26|28|vectis autem medius transibit per medias tabulas a summo usque ad summum.
EXOD|26|29|Ipsasque tabulas deaurabis et fundes eis anulos aureos, per quos vectes tabulata contineant, quos operies laminis aureis.
EXOD|26|30|Et eriges habitaculum iuxta exemplar, quod tibi in monte monstratum est.
EXOD|26|31|Facies et velum de hyacintho et purpura coccoque et bysso retorta, opere polymito, cum cherubim intextis.
EXOD|26|32|Quod appendes in quattuor columnis de lignis acaciae, quae ipsae quidem deauratae erunt et habebunt uncos aureos, sed bases argenteas.
EXOD|26|33|Inseres autem velum subter fibulas, intra quod pones arcam testimonii et quo sanctum et sanctum sanctorum dividentur.
EXOD|26|34|Pones et propitiatorium super arcam testimonii in sancto sanctorum
EXOD|26|35|mensamque extra velum et contra mensam candelabrum in latere habitaculi meridiano; mensa enim stabit in parte aquilonis.
EXOD|26|36|Facies et velum in introitu tabernaculi de hyacintho et purpura coccoque et bysso retorta opere plumarii.
EXOD|26|37|Et quinque columnas deaurabis lignorum acaciae, ante quas ducetur velum, quarum erunt unci aurei et bases aeneae.
EXOD|27|1|Facies et altare de lignis acaciae, quod habebit quinque cubitos in longitudine et totidem in latitudine, id est quadrum, et tres cubitos in altitudine.
EXOD|27|2|Cornua autem per quattuor angulos ex ipso erunt, et operies illud aere.
EXOD|27|3|Faciesque in usus eius lebetes ad suscipiendos cineres et vatilla et pateras atque fuscinulas et ignium receptacula; omnia vasa ex aere fabricabis.
EXOD|27|4|Craticulamque facies ei in modum retis aeneam, per cuius quattuor angulos erunt quattuor anuli aenei,
EXOD|27|5|et pones eam subter marginem altaris; eritque craticula usque ad altaris medium.
EXOD|27|6|Facies et vectes altaris de lignis acaciae duos, quos operies laminis aeneis,
EXOD|27|7|et induces per anulos; eruntque ex utroque latere altaris ad portandum.
EXOD|27|8|Cavum ex tabulis facies illud; sicut tibi in monte monstratum est, sic facient.
EXOD|27|9|Facies et atrium habitaculi, in cuius plaga australi contra meridiem erunt tentoria de bysso retorta: centum cubitos unum latus tenebit in longitudine
EXOD|27|10|et columnas viginti et bases totidem aeneas et uncos columnarum anulosque earum argenteos.
EXOD|27|11|Similiter in latere aquilonis: per longum erunt tentoria centum cubitorum, columnae viginti et bases aeneae eiusdem numeri et unci columnarum anulique earum argentei.
EXOD|27|12|In latitudine vero atrii, quae respicit ad occidentem, erunt tentoria per quinquaginta cubitos et columnae decem basesque totidem.
EXOD|27|13|In ea quoque atrii latitudine, quae respicit ad orientem, quinquaginta cubiti erunt,
EXOD|27|14|in quibus quindecim cubitorum tentoria lateri uno deputabuntur columnaeque tres et bases totidem;
EXOD|27|15|et in latere altero erunt tentoria, cubitos obtinentia quindecim, columnae tres et bases totidem.
EXOD|27|16|In introitu vero atrii fiet velum cubitorum viginti, ex hyacintho et purpura coccoque et bysso retorta opere plumarii; columnas habebit quattuor cum basibus totidem.
EXOD|27|17|Omnes columnae atrii per circuitum cinctae erunt anulis argenteis, et unci earum erunt argentei et bases aeneae.
EXOD|27|18|In longitudine occupabit atrium cubitos centum, in latitudine quinquaginta, altitudo quinque cubitorum erit; fietque de bysso retorta, et habebit bases aeneas.
EXOD|27|19|Cuncta vasa habitaculi in omnes usus eius et omnes paxillos eius et omnes paxillos atrii ex aere facies.
EXOD|27|20|Praecipe filiis Israel, ut afferant tibi oleum de arboribus olivarum purissimum piloque contusum, ut ardeat lucerna semper
EXOD|27|21|in tabernaculo conventus, extra velum, quod oppansum est testimonio. Et parabunt eam Aaron et filii eius, ut a vespere usque mane luceat coram Domino. Perpetuus erit cultus per successiones eorum a filiis Israel.
EXOD|28|1|Applica quoque ad te Aaron fratrem tuum cum filiis suis de medio filiorum Israel, ut sacerdotio fungantur mihi: Aaron, Nadab et Abiu, Eleazar et Ithamar.
EXOD|28|2|Faciesque vestes sanctas Aaron fratri tuo in gloriam et decorem;
EXOD|28|3|et loqueris cunctis sapientibus corde, quos replevi spiritu prudentiae, ut faciant vestes Aaron, in quibus sanctificatus ministret mihi.
EXOD|28|4|Haec autem erunt vestimenta, quae facient: pectorale et ephod, tunicam et subuculam textam, tiaram et balteum. Facient vestimenta sancta Aaron fratri tuo et filiis eius, ut sacerdotio fungantur mihi;
EXOD|28|5|accipientque aurum et hyacinthum et purpuram coccumque et byssum.
EXOD|28|6|Facient autem ephod de auro et hyacintho ac purpura coccoque bysso retorta opere polymito.
EXOD|28|7|Duas fascias umerales habebit et in utroque latere summitatum suarum copulabitur cum eis.
EXOD|28|8|Et balteus super ephod ad constringendum, eiusdem operis et unum cum eo, erit ex auro et hyacintho et purpura coccoque et bysso retorta.
EXOD|28|9|Sumesque duos lapides onychinos et sculpes in eis nomina filiorum Israel:
EXOD|28|10|sex nomina in lapide uno et sex reliqua in altero, iuxta ordinem nativitatis eorum.
EXOD|28|11|Opere sculptoris et caelatura gemmarii sculpes eos nominibus filiorum Israel, inclusos textura aurea;
EXOD|28|12|et pones duos lapides super fascias umerales ephod, lapides memorialis filiorum Israel. Portabitque Aaron nomina eorum coram Domino super utrumque umerum ob recordationem.
EXOD|28|13|Facies ergo margines textas ex auro
EXOD|28|14|et duas catenulas ex auro purissimo quasi funiculos opus tortile et inseres catenulas tortas marginibus.
EXOD|28|15|Pectorale quoque iudicii facies opere polymito, iuxta texturam ephod, ex auro, hyacintho et purpura coccoque et bysso retorta.
EXOD|28|16|Quadrangulum erit et duplex; mensuram palmi habebit tam in longitudine quam in latitudine.
EXOD|28|17|Ponesque in eo quattuor ordines lapidum: in primo versu erit lapis sardius et topazius et smaragdus;
EXOD|28|18|in secundo carbunculus, sapphirus et iaspis;
EXOD|28|19|in tertio hyacinthus, achates et amethystus;
EXOD|28|20|in quarto chrysolithus, onychinus et beryllus. Inclusi auro erunt per ordines suos.
EXOD|28|21|Habebuntque nomina filiorum Israel: duodecim nominibus caelabuntur, singuli lapides nominibus singulorum per duodecim tribus.
EXOD|28|22|Facies in pectorali catenas quasi funiculos, opus tortile, ex auro purissimo;
EXOD|28|23|et duos anulos aureos, quos pones in utraque pectoralis summitate;
EXOD|28|24|catenasque aureas iunges anulis, qui sunt in marginalibus eius;
EXOD|28|25|et ipsarum catenarum extrema duobus copulabis marginibus in fasciis umeralibus ephod in parte eius anteriore.
EXOD|28|26|Facies et duos anulos aureos, quos pones in summitatibus pectoralis in ora interiore, quae respicit ephod.
EXOD|28|27|Necnon et alios duos anulos aureos, qui ponendi sunt in utraque fascia umerali ephod deorsum, versus partem anteriorem eius iuxta iuncturam eius supra balteum ephod,
EXOD|28|28|et stringatur pectorale anulis suis cum anulis ephod vitta hyacinthina, ut maneat supra balteum ephod, et a se invicem pectorale et ephod nequeant separari.
EXOD|28|29|Portabitque Aaron nomina filiorum Israel in pectorali iudicii super cor suum, quando ingredietur sanctuarium: memoriale coram Domino in aeternum.
EXOD|28|30|Pones autem in pectorali iudicii Urim et Tummim, quae erunt super cor Aaron, quando ingredietur coram Domino; et gestabit iudicium filiorum Israel super cor suum in conspectu Domini semper.
EXOD|28|31|Facies et pallium ephod totum hyacinthinum,
EXOD|28|32|in cuius medio supra erit capitium et ora per gyrum eius textilis, sicut in capitio loricae, ne rumpatur.
EXOD|28|33|Deorsum vero, ad pedes eiusdem pallii per circuitum, quasi mala punica facies ex hyacintho et purpura et cocco, mixtis in medio tintinnabulis aureis;
EXOD|28|34|ita ut sit tintinnabulum aureum inter singula mala punica.
EXOD|28|35|Et vestietur eo Aaron in officio ministerii, ut audiatur sonitus, quando ingreditur et egreditur sanctuarium in conspectu Domini, et non moriatur.
EXOD|28|36|Facies et laminam de auro purissimo, in qua sculpes opere caelatoris: "Sanctum Domino".
EXOD|28|37|Ligabisque eam vitta hyacinthina, et erit super tiaram
EXOD|28|38|super frontem Aaron. Portabitque Aaron iniquitatem contra sancta, quae sanctificabunt filii Israel in cunctis muneribus et donariis suis. Eritque lamina semper in fronte eius, ut placatus eis sit Dominus.
EXOD|28|39|Texesque tunicam bysso et tiaram byssinam facies et balteum opere plumarii.
EXOD|28|40|Porro filiis Aaron tunicas lineas parabis et balteos ac mitras in gloriam et decorem;
EXOD|28|41|vestiesque his omnibus Aaron fratrem tuum et filios eius cum eo. Et unges eos et implebis manus eorum sanctificabisque illos, ut sacerdotio fungantur mihi.
EXOD|28|42|Facies eis et feminalia linea, ut operiant carnem turpitudinis suae a renibus usque ad femora;
EXOD|28|43|et utentur eis Aaron et filii eius, quando ingredientur tabernaculum conventus, vel quando appropinquant ad altare, ut ministrent in sanctuario, ne iniquitatis rei moriantur: legitimum sempiternum erit Aaron et semini eius post eum.
EXOD|29|1|Sed et hoc facies eis, ut mihi in sacerdotio consecrentur: tolle vitulum unum de armento et arietes duos immaculatos
EXOD|29|2|panesque azymos et crustulas absque fermento, quae conspersa sint oleo, lagana quoque azyma oleo lita; de simila triticea cuncta facies
EXOD|29|3|et posita in canistro offeres, vitulum quoque et duos arietes.
EXOD|29|4|Aaron ac filios eius applicabis ad ostium tabernaculi conventus. Cumque laveris patrem cum filiis suis aqua,
EXOD|29|5|indues Aaron vestimentis suis, id est subucula et tunica ephod et ephod et pectorali, quod constringes ei cingulo ephod;
EXOD|29|6|et pones tiaram in capite eius et diadema sanctum super tiaram
EXOD|29|7|et oleum unctionis fundes super caput eius; atque hoc ritu consecrabitur.
EXOD|29|8|Filios quoque illius applicabis et indues tunicis lineis cingesque balteo
EXOD|29|9|et impones eis mitras; eruntque sacerdotes mihi iure perpetuo.Postquam impleveris manus Aaron et filiorum eius,
EXOD|29|10|applicabis et vitulum coram tabernaculo conventus; imponentque Aaron et filii eius manus super caput illius,
EXOD|29|11|et mactabis eum in conspectu Domini, iuxta ostium tabernaculi conventus.
EXOD|29|12|Sumptumque de sanguine vituli, pones super cornua altaris digito tuo, reliquum autem sanguinem fundes iuxta basim eius.
EXOD|29|13|Sumes et adipem totum, qui operit intestina, et reticulum iecoris ac duos renes et adipem, qui super eos est, et offeres comburens super altare;
EXOD|29|14|carnes vero vituli et corium et fimum combures foris extra castra, eo quod pro peccato sit.
EXOD|29|15|Unum quoque arietem sumes, super cuius caput ponent Aaron et filii eius manus;
EXOD|29|16|quem cum mactaveris, tolles sanguinem eius et fundes super altare per circuitum.
EXOD|29|17|Ipsum autem arietem secabis in frusta lotaque intestina eius ac pedes pones super concisas carnes et super caput illius.
EXOD|29|18|Et adolebis totum arietem super altare: holocaustum est Domino, odor suavissimus, incensum est Domino.
EXOD|29|19|Tolles quoque arietem alterum, super cuius caput Aaron et filii eius ponent manus;
EXOD|29|20|quem cum immolaveris, sumes de sanguine ipsius et pones super extremum auriculae dextrae Aaron et filiorum eius et super pollices manus eorum ac pedis dextri; fundesque sanguinem super altare per circuitum.
EXOD|29|21|Cumque tuleris de sanguine, qui est super altare, et de oleo unctionis, asperges Aaron et vestes eius, filios et vestimenta eorum cum ipso. Et sanctus erit ipse et vestimenta eius et filii eius et vestimenta eorum cum ipso.
EXOD|29|22|Tollesque adipem de ariete et caudam et arvinam, quae operit intestina, ac reticulum iecoris et duos renes atque adipem, qui super eos est, armumque dextrum, eo quod sit aries consecrationis,
EXOD|29|23|tortamque panis unam, crustulam unam conspersam oleo, laganum unum de canistro azymorum, quod positum est in conspectu Domini;
EXOD|29|24|ponesque omnia super manus Aaron et filiorum eius, ut agitent ea coram Domino.
EXOD|29|25|Suscipiesque universa de manibus eorum et incendes in altari super holocausto in odorem suavissimum in conspectu Domini; quia incensum est Domino.
EXOD|29|26|Sumes quoque pectusculum de ariete, quo initiatus est Aaron, elevabisque illud coram Domino; et cedet in partem tuam.
EXOD|29|27|Sanctificabisque pectusculum elevatum et armum oblatum, quem de ariete separasti,
EXOD|29|28|quo initiatus est Aaron et filii eius; cedentque in partem Aaron et filiorum eius iure perpetuo a filiis Israel; quia oblatio est et oblatio erit a filiis Israel de victimis eorum pacificis, oblatio eorum Domino.
EXOD|29|29|Vestem autem sanctam, qua utetur Aaron, habebunt filii eius post eum, ut ungantur in ea, et impleantur in ea manus eorum.
EXOD|29|30|Septem diebus utetur illa, qui pontifex pro eo fuerit constitutus de filiis eius, qui ingredietur tabernaculum conventus, ut ministret in sanctuario.
EXOD|29|31|Arietem autem consecrationis tolles et coques carnes eius in loco sancto.
EXOD|29|32|Et vescetur Aaron et filii eius carnibus arietis et panibus, qui sunt in canistro, in vestibulo tabernaculi conventus.
EXOD|29|33|Et comedent ea, quibus expiatio facta fuerit ad implendum manus eorum, ad sanctificandum eos. Alienigena non vescetur ex eis, quia sancta sunt.
EXOD|29|34|Quod si remanserit de carnibus consecrationis sive de panibus usque mane, combures reliquias igni; non comedentur, quia sancta sunt.
EXOD|29|35|Omnia, quae praecepi tibi, facies super Aaron et filiis eius. Septem diebus consecrabis manus eorum
EXOD|29|36|et vitulum pro peccato offeres per singulos dies ad expiandum. Mundabisque altare expians illud et unges illud in sanctificationem.
EXOD|29|37|Septem diebus expiabis altare et sanctificabis; et erit sanctum sanctorum: omnis, qui tetigerit illud, sanctificabitur.
EXOD|29|38|Hoc est quod facies in altari: agnos anniculos duos per singulos dies iugiter,
EXOD|29|39|unum agnum mane et alterum vespere;
EXOD|29|40|decimam partem similae conspersae oleo tunso, quod habeat mensuram quartam partem hin, et vinum ad libandum eiusdem mensurae in agno uno.
EXOD|29|41|Alterum vero agnum offeres ad vesperam iuxta ritum matutinae oblationis et libationis in odorem suavitatis, incensum Domino,
EXOD|29|42|holocaustum perpetuum in generationes vestras, ad ostium tabernaculi conventus coram Domino, ubi conveniam vos, ut loquar ad te.
EXOD|29|43|Ibi conveniam filios Israel, et sanctificabitur locus in gloria mea.
EXOD|29|44|Sanctificabo et tabernaculum conventus cum altari et Aaron cum filiis eius, ut sacerdotio fungantur mihi.
EXOD|29|45|Et habitabo in medio filiorum Israel eroque eis Deus;
EXOD|29|46|et scient quia ego Dominus Deus eorum, qui eduxi eos de terra Aegypti, ut manerem inter illos: ego Dominus Deus ipsorum.
EXOD|30|1|Facies quoque altare ad adolendum thymiama de lignis acaciae
EXOD|30|2|habens cubitum longitudinis et alterum latitudinis, id est quadrangulum, et duos cubitos in altitudine; cornua ex ipso procedent.
EXOD|30|3|Vestiesque illud auro purissimo, tam craticulam eius quam parietes per circuitum et cornua. Faciesque ei coronam aureolam per gyrum
EXOD|30|4|et duos anulos aureos sub corona in duobus lateribus, ut mittantur in eos vectes, et altare portetur.
EXOD|30|5|Ipsos quoque vectes facies de lignis acaciae et inaurabis.
EXOD|30|6|Ponesque altare contra velum, quod ante arcam pendet testimonii, coram propitiatorio, quo tegitur testimonium, ubi conveniam ad te.
EXOD|30|7|Et adolebit incensum super eo Aaron suave fragrans mane. Quando componet lucernas, incendet illud;
EXOD|30|8|et quando collocabit eas ad vesperum, uret thymiama sempiternum coram Domino in generationes vestras.
EXOD|30|9|Non offeretis super eo thymiama compositionis alterius nec holocaustum nec oblationem, nec libabitis libamina.
EXOD|30|10|Et expiabit Aaron super cornua eius semel per annum in sanguine sacrificii pro peccato; et placabit super eo in generationibus vestris: sanctum sanctorum erit Domino ".
EXOD|30|11|Locutusque est Dominus ad Moysen dicens:
EXOD|30|12|" Quando tuleris summam filiorum Israel iuxta numerum, dabunt singuli pretium expiationis pro animabus suis Domino; et non erit plaga in eis, cum fuerint recensiti.
EXOD|30|13|Hoc autem dabit omnis, qui transit ad censum, dimidium sicli iuxta mensuram sanctuarii ­ siclus viginti obolos habet ­; media pars sicli offeretur Domino.
EXOD|30|14|Qui habetur in numero a viginti annis et supra, dabit pretium;
EXOD|30|15|dives non addet ad medium sicli, et pauper nihil minuet, quando dabitis oblationem Domino in expiationem animarum vestrarum.
EXOD|30|16|Susceptamque expiationis pecuniam, quae collata est a filiis Israel, trades in usus tabernaculi conventus, ut sit monumentum eorum coram Domino et propitietur animabus illorum ".
EXOD|30|17|Locutusque est Dominus ad Moysen dicens:
EXOD|30|18|" Facies et labrum aeneum cum basi aenea ad lavandum; ponesque illud inter tabernaculum conventus et altare. Et, missa aqua,
EXOD|30|19|lavabunt in eo Aaron et filii eius manus suas ac pedes.
EXOD|30|20|Quando ingressuri sunt tabernaculum conventus, lavabunt se aqua, ne moriantur; vel quando accessuri sunt ad altare, ut ministrent, ut adoleant victimam Domino.
EXOD|30|21|Et lavabunt manus et pedes, ne moriantur: legitimum sempiternum erit, ipsi et semini eius per successiones ".
EXOD|30|22|Locutusque est Dominus ad Moysen
EXOD|30|23|dicens: " Sume tibi aromata prima myrrhae electae quingentos siclos et cinnamomi boni odoris medium, id est ducentos quinquaginta siclos, calami suave olentis similiter ducentos quinquaginta,
EXOD|30|24|casiae autem quingentos siclos, in pondere sanctuarii, olei de olivetis mensuram hin.
EXOD|30|25|Faciesque unctionis oleum sanctum, unguentum compositum opere unguentarii; unctionis oleum sanctum erit.
EXOD|30|26|Et unges ex eo tabernaculum conventus et arcam testamenti
EXOD|30|27|mensamque cum vasis suis, candelabrum et utensilia eius, altaria thymiamatis
EXOD|30|28|et holocausti et universam supellectilem, quae ad cultum eorum pertinet, et labrum cum basi sua.
EXOD|30|29|Sanctificabisque omnia, et erunt sancta sanctorum: qui tetigerit ea, sanctificabitur.
EXOD|30|30|Aaron et filios eius unges sanctificabisque eos, ut sacerdotio fungantur mihi.
EXOD|30|31|Filiis quoque Israel dices: Hoc oleum unctionis sanctum erit mihi in generationes vestras.
EXOD|30|32|Caro hominis non ungetur ex eo, et iuxta compositionem eius non facietis aliud, quia sanctum est et sanctum erit vobis.
EXOD|30|33|Homo quicumque tale composuerit et dederit ex eo super alienum, exterminabitur de populo suo ".
EXOD|30|34|Dixitque Dominus ad Moysen: " Sume tibi aromata, stacten et onycha, galbanum boni odoris et tus lucidissimum; aequalis ponderis erunt omnia.
EXOD|30|35|Faciesque thymiama compositum opere unguentarii, sale conditum et purum et sanctum.
EXOD|30|36|Cumque in tenuissimum pulverem ex parte contuderis, pones ex eo coram testimonio in tabernaculo conventus, in quo conveniam ad te: sanctum sanctorum erit vobis thymiama.
EXOD|30|37|Talem compositionem non facietis in usus vestros, quia tibi sanctum erit pro Domino;
EXOD|30|38|homo quicumque fecerit simile, ut odore illius perfruatur, peribit de populis suis ".
EXOD|31|1|Locutusque est Dominus ad Moysen dicens:
EXOD|31|2|" Ecce voca vi ex nomine Beseleel filium Uri filii Hur de tribu Iudae
EXOD|31|3|et implevi eum spiritu Dei, sapientia et intellegentia et scientia in omni opere
EXOD|31|4|ad excogitandum, quidquid fabrefieri potest ex auro et argento et aere,
EXOD|31|5|ad scindendum et includendum gemmas et ad sculpendum ligna, ad faciendum omne opus;
EXOD|31|6|dedique ei socium Ooliab filium Achisamech de tribu Dan et in corde omnis eruditi posui sapientiam, ut faciant cuncta, quae praecepi tibi:
EXOD|31|7|tabernaculum conventus et arcam testimonii et propitiatorium, quod super eam est, et cuncta vasa tabernaculi
EXOD|31|8|mensamque et vasa eius, candelabrum purissimum cum vasis suis et altaria thymiamatis
EXOD|31|9|et holocausti et omnia vasa eorum, labrum cum basi sua
EXOD|31|10|et vestes textas et vestes sanctas Aaron sacerdoti et vestes filiorum eius, ut fungantur officio suo in sacris,
EXOD|31|11|oleum unctionis et thymiama aromatum in sanctuario: omnia, quae praecepi tibi, facient ".
EXOD|31|12|Et locutus est Dominus ad Moysen dicens:
EXOD|31|13|" Loquere filiis Israel et dices ad eos: Videte ut sabbatum meum custodiatis, quia signum est inter me et vos in generationibus vestris, ut sciatis quia ego Dominus, qui sanctifico vos.
EXOD|31|14|Custodite sabbatum, sanctum est enim vobis. Qui polluerit illud, morte morietur; qui fecerit in eo opus, peribit anima illius de medio populi sui.
EXOD|31|15|Sex diebus facietis opus; in die septimo sabbatum est, requies sancta Domino: omnis, qui fecerit opus in hac die, morietur.
EXOD|31|16|Custodiant filii Israel sabbatum et celebrent illud in generationibus suis: pactum est sempiternum
EXOD|31|17|inter me et filios Israel signumque perpetuum; sex enim diebus fecit Dominus caelum et terram et in septimo ab opere cessavit et respiravit ".
EXOD|31|18|Deditque Dominus Moysi, completis huiuscemodi sermonibus in monte Sinai, duas tabulas testimonii lapideas scriptas digito Dei.
EXOD|32|1|Videns autem populus quod moram faceret descendendi de monte Moyses, congregatus ad Aaron dixit: " Surge, fac nobis deos, qui nos praecedant; Moysi enim, huic viro, qui nos eduxit de terra Aegypti, ignoramus quid acciderit ".
EXOD|32|2|Dixitque ad eos Aaron: " Tollite inaures aureas de uxorum filiorumque et filiarum vestrarum auribus et afferte ad me ".
EXOD|32|3|Fecitque omnis populus, quae iusserat, deferens inaures ad Aaron.
EXOD|32|4|Quas cum ille accepisset, formavit stilo imaginem et fecit ex eis vitulum conflatilem. Dixeruntque: " Hi sunt dii tui, Israel, qui te eduxerunt de terra Aegypti! ".
EXOD|32|5|Quod cum vidisset Aaron, aedificavit altare coram eo et praeconis voce clamavit dicens: " Cras sollemnitas Domini est ".
EXOD|32|6|Surgen tesque mane altero die obtulerunt holocausta et hostias pacificas; et sedit populus manducare et bibere et surrexerunt ludere.
EXOD|32|7|Locutus est autem Dominus ad Moysen: " Vade, descende; peccavit populus tuus, quem eduxisti de terra Aegypti.
EXOD|32|8|Recesserunt cito de via, quam praecepi eis, feceruntque sibi vitulum conflatilem et adoraverunt atque immolantes ei hostias dixerunt: "Isti sunt dii tui, Israel, qui te eduxerunt de terra Aegypti!" ".
EXOD|32|9|Rursumque ait Dominus ad Moysen: " Cerno quod populus iste durae cervicis sit;
EXOD|32|10|dimitte me, ut irascatur furor meus contra eos et deleam eos faciamque te in gentem magnam ".
EXOD|32|11|Moyses autem orabat Dominum Deum suum dicens: " Cur, Domine, irascitur furor tuus contra populum tuum, quem eduxisti de terra Aegypti in fortitudine magna et in manu robusta?
EXOD|32|12|Ne, quaeso, dicant Aegyptii: "Callide eduxit eos, ut interficeret in montibus et deleret e terra". Quiescat ira tua, et esto placabilis super nequitia populi tui.
EXOD|32|13|Recordare Abraham, Isaac et Israel servorum tuorum, quibus iurasti per temetipsum dicens: "Multiplicabo semen vestrum sicut stellas caeli; et universam terram hanc, de qua locutus sum, dabo semini vestro, et possidebitis eam semper" ".
EXOD|32|14|Placatusque est Dominus, ne faceret malum, quod locutus fuerat adversus populum suum.
EXOD|32|15|Et reversus est Moyses de monte portans duas tabulas testimonii in manu sua scriptas ex utraque parte
EXOD|32|16|et factas opere Dei; scriptura quoque Dei erat sculpta in tabulis.
EXOD|32|17|Audiens autem Iosue tumultum populi vociferantis dixit ad Moysen: " Ululatus pugnae auditur in castris ".
EXOD|32|18|Qui respondit:" Non est clamor vincentiumneque clamor fugientium,sed clamorem cantantiumego audio ".
EXOD|32|19|Cumque appropinquasset ad castra, vidit vitulum et choros; iratusque valde proiecit de manu tabulas et confregit eas ad radices montis.
EXOD|32|20|Arripiensque vitulum, quem fecerant, combussit et contrivit usque ad pulverem, quem sparsit in aquam et dedit ex eo potum filiis Israel.
EXOD|32|21|Dixitque ad Aaron: " Quid tibi fecit hic populus, ut induceres super eum peccatum maximum? ".
EXOD|32|22|Cui ille respondit: " Ne indignetur dominus meus; tu enim nosti populum istum, quod pronus sit ad malum.
EXOD|32|23|Dixerunt mihi: "Fac nobis deos, qui nos praecedant; huic enim Moysi, qui nos eduxit de terra Aegypti, nescimus quid acciderit".
EXOD|32|24|Quibus ego dixi: Quis vestrum habet aurum? Abstulerunt et dederunt mihi, et proieci illud in ignem; egressusque est hic vitulus ".
EXOD|32|25|Vidit ergo Moyses populum quod esset effrenatus; relaxaverat enim ei Aaron frenum in ludibrium hostium eorum.
EXOD|32|26|Et stans in porta castrorum ait: " Si quis est Domini, iungatur mihi! ". Congregatique sunt ad eum omnes filii Levi.
EXOD|32|27|Quibus ait: " Haec dicit Dominus, Deus Israel: Ponat unusquisque gladium super femur suum. Ite et redite de porta usque ad portam per medium castrorum, et occidat unusquisque fratrem et amicum et proximum suum ".
EXOD|32|28|Fecerunt filii Levi iuxta sermonem Moysi; cecideruntque de populo in die illa quasi tria milia hominum.
EXOD|32|29|Et ait Moyses: " Implestis manus vestras hodie Domino unusquisque in filio et in fratre suo, ut detur vobis benedictio ".
EXOD|32|30|Facto autem altero die, locutus est Moyses ad populum: " Peccastis peccatum maximum; ascendam ad Dominum, si quo modo quivero eum deprecari pro scelere vestro ".
EXOD|32|31|Reversusque ad Dominum ait: " Obsecro, peccavit populus iste peccatum maximum, feceruntque sibi deos aureos; aut dimitte eis hanc noxam
EXOD|32|32|aut, si non facis, dele me de libro tuo, quem scripsisti ".
EXOD|32|33|Cui respondit Dominus: " Qui peccaverit mihi, delebo eum de libro meo.
EXOD|32|34|Tu autem vade et duc populum istum, quo locutus sum tibi: angelus meus praecedet te; ego autem in die ultionis visitabo et hoc peccatum eorum ".
EXOD|32|35|Percussit ergo Dominus populum pro reatu vituli, quem fecerat Aaron.
EXOD|33|1|Locutusque est Dominus ad Moysen: " Vade, ascende de loco isto, tu et populus tuus, quem eduxisti de terra Aegypti, in terram, quam iuravi Abraham, Isaac et Iacob dicens: Semini tuo dabo eam.
EXOD|33|2|Et mittam praecursorem tui angelum et eiciam Chananaeum et Amorraeum et Hetthaeum et Pherezaeum et Hevaeum et Iebusaeum,
EXOD|33|3|et intres in terram fluentem lacte et melle. Non enim ascendam tecum, quia populus durae cervicis es, ne forte disperdam te in via ".
EXOD|33|4|Audiens populus sermonem hunc pessimum luxit, et nullus ex more indutus est cultu suo.
EXOD|33|5|Dixitque Dominus ad Moysen: " Loquere filiis Israel: Populus durae cervicis es; uno momento, si ascendam in medio tui, delebo te. Nunc autem depone ornatum tuum, ut sciam quid faciam tibi ".
EXOD|33|6|Deposuerunt ergo filii Israel ornatum suum a monte Horeb.
EXOD|33|7|Moyses autem tollens tabernaculum tetendit ei extra castra procul; vocavitque nomen eius Tabernaculum conventus. Et omnis, qui quaerebat Dominum, egrediebatur ad tabernaculum conventus extra castra.
EXOD|33|8|Cumque egrederetur Moyses ad tabernaculum, surgebat universa plebs, et stabat unusquisque in ostio papilionis sui; aspiciebantque tergum Moysi, donec ingrederetur tabernaculum.
EXOD|33|9|Ingresso autem illo tabernaculum, descendebat columna nubis et stabat ad ostium; loquebaturque cum Moyse,
EXOD|33|10|cernentibus universis quod columna nubis staret ad ostium tabernaculi. Stabantque ipsi et adorabant per fores tabernaculorum suorum.
EXOD|33|11|Loquebatur autem Dominus ad Moysen facie ad faciem, sicut solet loqui homo ad amicum suum. Cumque ille reverteretur in castra, minister eius Iosue filius Nun puer non recedebat de medio tabernaculi.
EXOD|33|12|Dixit autem Moyses ad Dominum: " Praecipis, ut educam populum istum, et non indicas mihi, quem missurus es mecum; cum dixeris: "Novi te ex nomine, et invenisti gratiam coram me".
EXOD|33|13|Si ergo inveni gratiam in conspectu tuo, ostende mihi viam tuam, ut sciam te et inveniam gratiam ante oculos tuos; respice quia populus tuus est natio haec ".
EXOD|33|14|Dixitque Dominus: " Facies mea ibit, et requiem dabo tibi ".
EXOD|33|15|Et ait Moyses: " Si non tu ipse eas, ne educas nos de loco isto;
EXOD|33|16|in quo enim scietur me et populum tuum invenisse gratiam in conspectu tuo, nisi ambulaveris nobiscum, ut glorificemur ego et populus tuus prae omnibus populis, qui habitant super terram? ".
EXOD|33|17|Dixitque Dominus ad Moysen: " Et verbum istud, quod locutus es, faciam; invenisti enim gratiam coram me, et teipsum novi ex nomine ".
EXOD|33|18|Qui ait: " Ostende mihi gloriam tuam ".
EXOD|33|19|Respondit: " Ego ostendam omne bonum tibi et vocabo in nomine Domini coram te; et miserebor, cui voluero, et clemens ero, in quem mihi placuerit ".
EXOD|33|20|Rursumque ait: " Non poteris videre faciem meam; non enim videbit me homo et vivet ".
EXOD|33|21|Et iterum: " Ecce, inquit, est locus apud me, stabis super petram;
EXOD|33|22|cumque transibit gloria mea, ponam te in foramine petrae et protegam dextera mea, donec transeam;
EXOD|33|23|tollamque manum meam, et videbis posteriora mea; faciem autem meam videre non poteris ".
EXOD|34|1|Dixitque Dominus ad Moy sen: " Praecide tibi duas ta bulas lapideas instar priorum, et scribam super eas verba, quae habuerunt tabulae, quas fregisti.
EXOD|34|2|Esto paratus mane, ut ascendas statim in montem Sinai; stabisque mihi super verticem montis.
EXOD|34|3|Nullus ascendat tecum, nec videatur quispiam per totum montem; oves quoque et boves non pascantur e contra ".
EXOD|34|4|Excidit ergo duas tabulas lapideas, quales antea fuerant; et de nocte consurgens ascendit in montem Sinai, sicut praeceperat ei Dominus, portans secum tabulas.
EXOD|34|5|Cumque descendisset Dominus per nubem, stetit cum eo vocans in nomine Domini.
EXOD|34|6|Et transiens coram eo clamavit: " Dominus, Dominus Deus, misericors et clemens, patiens et multae miserationis ac verax,
EXOD|34|7|qui custodit misericordiam in milia, qui aufert iniquitatem et scelera atque peccata, nihil autem impunitum sinit, qui reddit iniquitatem patrum in filiis ac nepotibus in tertiam et quartam progeniem ".
EXOD|34|8|Festinusque Moyses curvatus est pronus in terram et adorans
EXOD|34|9|ait: " Si inveni gratiam in conspectu tuo, Domine, obsecro, ut gradiaris nobiscum; populus quidem durae cervicis est, sed tu auferes iniquitates nostras atque peccata nosque possidebis ".
EXOD|34|10|Respondit Dominus: " Ego inibo pactum coram universo populo tuo; mirabilia faciam, quae numquam visa sunt super totam terram nec in ullis gentibus, ut cernat cunctus populus, in cuius es medio, opus Domini terribile, quod facturus sum tecum.
EXOD|34|11|Observa cuncta, quae hodie mando tibi: ego ipse eiciam ante faciem tuam Amorraeum et Chananaeum et Hetthaeum, Pherezaeum quoque et Hevaeum et Iebusaeum.
EXOD|34|12|Cave, ne umquam cum habitatoribus terrae, quam intraveris, iungas amicitias, quae tibi sint in ruinam;
EXOD|34|13|sed aras eorum destrue, confringe lapides palosque succide.
EXOD|34|14|Noli adorare deum alienum: Dominus Zelotes nomen eius, Deus est aemulator.
EXOD|34|15|Ne ineas pactum cum hominibus illarum regionum, ne, cum fornicati fuerint cum diis suis et sacrificaverint eis, vocet te quispiam, et comedas de immolatis.
EXOD|34|16|Nec uxorem de filiabus eorum accipies filiis tuis, ne, postquam ipsae fuerint fornicatae cum diis suis, fornicari faciant et filios tuos in deos suos.
EXOD|34|17|Deos conflatiles non facies tibi.
EXOD|34|18|Sollemnitatem Azymorum custodies: septem diebus vesceris azymis, sicut praecepi tibi, in tempore constituto mensis Abib; mense enim verni temporis egressus es de Aegypto.
EXOD|34|19|Omne, quod aperit vulvam generis masculini, meum erit; de cuncto grege tuo tam de bobus quam de ovibus meum erit.
EXOD|34|20|Primogenitum asini redimes ove, sin autem nec pretium pro eo dederis, franges cervicem eius. Primogenitum filiorum tuorum redimes; nec apparebis in conspectu meo vacuus.
EXOD|34|21|Sex diebus operaberis, die septimo cessabis etiam arare et metere.
EXOD|34|22|Sollemnitatem Hebdomadarum facies tibi in primitiis frugum messis tuae triticeae et sollemnitatem Collectae, quando, redeunte anni tempore, cuncta conduntur.
EXOD|34|23|Tribus temporibus anni apparebit omne masculinum tuum in conspectu omnipotentis Domini, Dei Israel.
EXOD|34|24|Cum enim tulero gentes a facie tua et dilatavero terminos tuos, nullus insidiabitur terrae tuae, ascendente te et apparente in conspectu Domini Dei tui ter in anno.
EXOD|34|25|Non immolabis super fermento sanguinem hostiae meae; neque residebit mane de victima sollemnitatis Paschae.
EXOD|34|26|Primitias frugum terrae tuae afferes in domum Domini Dei tui.Non coques haedum in lacte matris suae ".
EXOD|34|27|Dixitque Dominus ad Moysen: " Scribe tibi verba haec, quibus et tecum et cum Israel pepigi foedus ".
EXOD|34|28|Fuit ergo ibi cum Domino quadraginta dies et quadraginta noctes; panem non comedit et aquam non bibit et scripsit in tabulis verba foederis, decem verba.
EXOD|34|29|Cumque descenderet Moyses de monte Sinai, tenebat duas tabulas testimonii et ignorabat quod resplenderet cutis faciei suae ex consortio sermonis Domini.
EXOD|34|30|Videntes autem Aaron et filii Israel resplendere cutem faciei Moysi, timuerunt prope accedere;
EXOD|34|31|vocatique ab eo reversi sunt tam Aaron quam principes synagogae. Et postquam locutus est ad eos,
EXOD|34|32|venerunt ad eum etiam omnes filii Israel; quibus praecepit cuncta, quae audierat a Domino in monte Sinai.
EXOD|34|33|Impletisque sermonibus, posuit velamen super faciem suam,
EXOD|34|34|quod ingressus ad Dominum et loquens cum eo auferebat, donec exiret; et tunc loquebatur ad filios Israel omnia, quae sibi fuerant imperata.
EXOD|34|35|Qui videbant cutem faciei Moysi resplendere, sed operiebat ille rursus faciem suam, donec ingressus loqueretur cum eo.
EXOD|35|1|Igitur, congregato omni coetu filiorum Israel, dixit ad eos: " Haec sunt, quae iussit Dominus fieri:
EXOD|35|2|sex diebus facietis opus, septimus dies erit vobis sanctus, sabbatum et requies Domino; qui fecerit opus in eo, occidetur.
EXOD|35|3|Non succendetis ignem in omnibus habitaculis vestris per diem sabbati ".
EXOD|35|4|Et ait Moyses ad omnem coetum filiorum Israel: " Iste est sermo, quem praecepit Dominus dicens:
EXOD|35|5|"Separate apud vos donaria Domino". Omnis voluntarius et proni animi offerat ea Domino: aurum et argentum et aes,
EXOD|35|6|hyacinthum et purpuram coccumque et byssum, pilos caprarum
EXOD|35|7|et pelles arietum rubricatas et pelles delphini, ligna acaciae
EXOD|35|8|et oleum ad luminaria concinnanda et aromata, ut conficiatur unguentum et thymiama suavissimum,
EXOD|35|9|lapides onychinos et gemmas ad ornatum ephod et pectoralis.
EXOD|35|10|Quisquis vestrum sapiens est, veniat et faciat, quod Dominus imperavit,
EXOD|35|11|habitaculum scilicet et tentorium eius atque operimentum, fibulas et tabulata cum vectibus, columnas et bases;
EXOD|35|12|arcam et vectes, propitiatorium et velum, quod ante illud oppanditur;
EXOD|35|13|mensam cum vectibus et vasis et propositionis panibus;
EXOD|35|14|candelabrum ad luminaria sustentanda, vasa illius et lucernas et oleum ad nutrimenta luminarium;
EXOD|35|15|altare thymiamatis et vectes et oleum unctionis et thymiama ex aromatibus; velum ad ostium habitaculi;
EXOD|35|16|altare holocausti et craticulam eius aeneam cum vectibus et vasis suis, labrum et basim eius;
EXOD|35|17|cortinas atrii cum columnis et basibus, velum in foribus atrii;
EXOD|35|18|paxillos habitaculi et atrii cum funiculis suis;
EXOD|35|19|vestimenta texta, quorum usus est in ministerio sanctuarii, vestes sanctas Aaron pontificis ac vestes filiorum eius, ut sacerdotio fungantur mihi ".
EXOD|35|20|Egressus est omnis coetus filiorum Israel de conspectu Moysi,
EXOD|35|21|et venit, quisquis erat mentis promptissimae, et attulit sponte sua donaria Domino ad faciendum opus tabernaculi conventus et quidquid ad cultum et ad vestes sanctas necessarium erat.
EXOD|35|22|Viri cum mulieribus, omnes voluntarii praebuerunt fibulas et inaures, anulos et dextralia; omne vas aureum in donaria Domini separatum est.
EXOD|35|23|Si quis habebat hyacinthum et purpuram coccumque, byssum et pilos caprarum, pelles arietum rubricatas et pelles delphini,
EXOD|35|24|argenti aerisque metalla, obtulerunt Domino lignaque acaciae in varios usus.
EXOD|35|25|Sed et mulieres eruditae dederunt, quae neverant, hyacinthum, purpuram et coccum ac byssum
EXOD|35|26|et pilos caprarum, sponte propria cuncta tribuentes.
EXOD|35|27|Principes vero obtulerunt lapides onychinos et gemmas ad ephod et pectorale
EXOD|35|28|aromataque et oleum ad luminaria concinnanda et ad praeparandum unguentum ac thymiama odoris suavissimi componendum.
EXOD|35|29|Omnes viri et mulieres mente prompta obtulerunt donaria, ut fierent opera, quae iusserat Dominus per manum Moysi. Cuncti filii Israel voluntaria Domino dedicaverunt.
EXOD|35|30|Dixitque Moyses ad filios Israel: " Ecce vocavit Dominus ex nomine Beseleel filium Uri filii Hur de tribu Iudae;
EXOD|35|31|implevitque eum spiritu Dei, sapientia et intellegentia et scientia ad omne opus,
EXOD|35|32|ad excogitandum et faciendum opus in auro et argento et aere,
EXOD|35|33|ad scindendum et includendum gemmas et ad sculpendum ligna, quidquid fabre adinveniri potest.
EXOD|35|34|Dedit quoque in corde eius, ut alios doceret, ipsi et Ooliab filio Achisamech de tribu Dan.
EXOD|35|35|Ambos implevit sapientia, ut faciant opera fabri polymitarii ac plumarii de hyacintho ac purpura coccoque et bysso et textoris, facientes omne opus ac nova quaeque reperientes ".
EXOD|36|1|Fecit ergo Beseleel et Ooliab et omnis vir sapiens, quibus dedit Dominus sapientiam et intellectum, ut scirent fabre operari, quae in usus sanctuarii necessaria sunt et quae praecepit Dominus.
EXOD|36|2|Cumque vocasset Moyses Beseleel et Ooliab et omnem eruditum virum, cui dederat Dominus sapientiam, omnes, qui sponte sua obtulerant se ad faciendum opus,
EXOD|36|3|acceperunt ab ipso universa donaria, quae attulerant filii Israel ad faciendum opus in cultum sanctuarii. Ipsi autem cotidie mane donaria ei offerebant.
EXOD|36|4|Unde omnes sapientes artifices venerunt singuli de opere suo pro sanctuario
EXOD|36|5|et dixerunt Moysi: " Plus offert populus quam necessarium est operi, quod Dominus iussit facere ".
EXOD|36|6|Iussit ergo Moyses praeconis voce per castra clamari: " Nec vir nec mulier quidquam offerat ultra pro omni opere sanctuario ". Sicque cessatum est a muneribus offerendis,
EXOD|36|7|eo quod oblata sufficerent et superabundarent.
EXOD|36|8|Feceruntque omnes corde sapientes inter artifices habitaculi cortinas decem de bysso retorta et hyacintho et purpura coccoque, cum cherubim intextis arte polymita;
EXOD|36|9|quarum una habebat in longitudine viginti octo cubitos et in latitudine quattuor: una mensura erat omnium cortinarum.
EXOD|36|10|Coniunxitque cortinas quinque alteram alteri et alias quinque sibi invicem copulavit.
EXOD|36|11|Fecit et ansas hyacinthinas in ora cortinae unius in extremitate iuncturae et in ora cortinae extremae in iunctura altera similiter.
EXOD|36|12|Quinquagenas ansas fecit pro utraque cortina, ut contra se invicem venirent ansae et mutuo iungerentur.
EXOD|36|13|Unde et quinquaginta fudit fibulas aureas, quae morderent cortinarum ansas, et fieret unum habitaculum.
EXOD|36|14|Fecit et saga undecim de pilis caprarum pro tentorio super habitaculum;
EXOD|36|15|unum sagum in longitudine habebat cubitos triginta et in latitudine cubitos quattuor: unius mensurae erant omnia saga.
EXOD|36|16|Quorum quinque iunxit seorsum et sex alia separatim.
EXOD|36|17|Fecitque ansas quinquaginta in ora sagi ultimi iuncturae unius et quinquaginta in ora sagi iuncturae alterius, ut sibi invicem iungerentur;
EXOD|36|18|et fecit fibulas aeneas quinquaginta, quibus necteretur tentorium, ut esset unum.
EXOD|36|19|Fecit et opertorium tentorio de pellibus arietum rubricatis aliudque desuper velamentum de pellibus delphini.
EXOD|36|20|Fecit et tabulas habitaculi de lignis acaciae stantes.
EXOD|36|21|Decem cubitorum erat longitudo tabulae unius, et unum ac semis cubitum latitudo retinebat.
EXOD|36|22|Bini pedes erant per singulas tabulas, ut altera alteri iungeretur: sic fecit in omnibus tabulis habitaculi.
EXOD|36|23|E quibus viginti ad plagam meridianam erant contra austrum
EXOD|36|24|cum quadraginta basibus argenteis. Duae bases sub singulis tabulis ponebantur pro duabus pedibus.
EXOD|36|25|Ad plagam quoque habitaculi, quae respicit ad aquilonem, fecit viginti tabulas
EXOD|36|26|cum quadraginta basibus argenteis: duas bases per singulas tabulas.
EXOD|36|27|Contra occidentem vero, id est ad eam partem habitaculi quae mare respicit, fecit sex tabulas
EXOD|36|28|et duas alias per singulos angulos habitaculi retro;
EXOD|36|29|quae gemellae erant a deorsum usque sursum in unam compaginem. Ita fecit duas tabulas in duobus angulis,
EXOD|36|30|ut octo essent simul tabulae et haberent bases argenteas sedecim: binas scilicet bases sub singulis tabulis.
EXOD|36|31|Fecit et vectes de lignis acaciae quinque ad continendas tabulas unius lateris habitaculi
EXOD|36|32|et quinque alios ad alterius lateris coaptandas tabulas; et extra hos quinque alios vectes ad occidentalem plagam habitaculi contra mare.
EXOD|36|33|Fecit autem vectem medium, qui per medias tabulas ab una extremitate usque ad alteram perveniret.
EXOD|36|34|Ipsa autem tabulata deauravit. Et anulos eorum fecit aureos, per quos vectes induci possent; quos et ipsos laminis aureis operuit.
EXOD|36|35|Fecit et velum de hyacintho et purpura coccoque ac bysso retorta, opere polymitario, cum cherubim intextis;
EXOD|36|36|et quattuor columnas de lignis acaciae, quas cum uncis suis deauravit, fusis basibus earum argenteis.
EXOD|36|37|Fecit et velum in introitu tabernaculi ex hyacintho, purpura, cocco byssoque retorta opere plumarii;
EXOD|36|38|et columnas quinque cum uncis suis. Et operuit auro capita et anulos earum basesque earum fudit aeneas.
EXOD|37|1|Fecit autem Beseleel et ar cam de lignis acaciae haben tem duos semis cubitos in longitudine et cubitum ac semissem in latitudine, altitudo quoque unius cubiti fuit et dimidii; vestivitque eam auro purissimo intus ac foris.
EXOD|37|2|Et fecit illi coronam auream per gyrum,
EXOD|37|3|conflans quattuor anulos aureos in quattuor pedibus eius; duos anulos in latere uno et duos in altero.
EXOD|37|4|Vectes quoque fecit de lignis acaciae, quos vestivit auro
EXOD|37|5|et quos misit in anulos, qui erant in lateribus arcae, ad portandum eam.
EXOD|37|6|Fecit et propitiatorium de auro mundissimo: duorum cubitorum et dimidii in longitudine et cubiti ac semis in latitudine.
EXOD|37|7|Duos etiam cherubim ex auro ductili fecit ex utraque parte propitiatorii:
EXOD|37|8|cherub unum ex summitate unius partis et cherub alterum ex summitate partis alterius; duos cherubim ex singulis summitatibus propitiatorii
EXOD|37|9|extendentes alas sursum et tegentes alis suis propitiatorium seque mutuo et illud respicientes.
EXOD|37|10|Fecit et mensam de lignis acaciae in longitudine duorum cubitorum et in latitudine unius cubiti, quae habebat in altitudine cubitum ac semissem;
EXOD|37|11|circumdeditque eam auro mundissimo et fecit illi coronam auream per gyrum.
EXOD|37|12|Fecit ei quoque limbum aureum quattuor digitorum per circuitum et super illum coronam auream.
EXOD|37|13|Fudit et quattuor circulos aureos, quos posuit in quattuor angulis per singulos pedes mensae
EXOD|37|14|iuxta limbum; misitque in eos vectes, ut possit mensa portari.
EXOD|37|15|Ipsos quoque vectes fecit de lignis acaciae et circumdedit eos auro;
EXOD|37|16|et vasa ad diversos usus mensae, acetabula, phialas et cyathos et crateras ex auro puro, in quibus offerenda sunt libamina.
EXOD|37|17|Fecit et candelabrum ductile de auro mundissimo, basim et hastile eius; scyphi sphaerulaeque ac flores unum cum ipso erant:
EXOD|37|18|sex in utroque latere, tres calami ex parte una et tres ex altera;
EXOD|37|19|tres scyphi in nucis modum in calamo uno sphaerulaeque simul et flores et tres scyphi instar nucis in calamo altero sphaerulaeque simul et flores. Aequum erat opus sex calamorum, qui procedebant de hastili candelabri.
EXOD|37|20|In ipso autem hastili erant quattuor scyphi in nucis modum sphaerulaeque et flores;
EXOD|37|21|singulae sphaerulae sub binis calamis per loca tria, qui simul sex fiunt calami procedentes de hastili uno.
EXOD|37|22|Sphaerulae igitur et calami unum cum ipso erant, totum ductile ex auro purissimo.
EXOD|37|23|Fecit et lucernas septem cum emunctoriis suis et vasa, ubi emuncta condantur, de auro mundissimo.
EXOD|37|24|Talentum auri purissimi appendebat candelabrum cum omnibus vasis suis.
EXOD|37|25|Fecit et altare thymiamatis de lignis acaciae habens per quadrum singulos cubitos et in altitudine duos; e cuius angulis procedebant cornua.
EXOD|37|26|Vestivitque illud auro purissimo cum craticula ac parietibus et cornibus.
EXOD|37|27|Fecitque ei coronam aureolam per gyrum et binos anulos aureos sub corona in duobus lateribus, ut mittantur in eos vectes, et possit altare portari.
EXOD|37|28|Ipsos autem vectes fecit de lignis acaciae et operuit laminis aureis.
EXOD|37|29|Composuit et oleum ad sanctificationis unguentum et thymiama de aromatibus mundissimis opere pigmentarii.
EXOD|38|1|Fecit et altare holocausti de lignis acaciae quinque cubi torum per quadrum et trium in altitudine,
EXOD|38|2|cuius cornua de angulis procedebant; operuitque illud laminis aeneis.
EXOD|38|3|Et in usus eius paravit ex aere vasa diversa: lebetes, vatilla et pateras, fuscinulas et ignium receptacula.
EXOD|38|4|Craticulamque eius in modum retis fecit aeneam subter marginem altaris ab imo usque ad medium eius,
EXOD|38|5|fusis quattuor anulis per totidem craticulae summitates, ad immittendos vectes ad portandum.
EXOD|38|6|Quos et ipsos fecit de lignis acaciae et operuit laminis aeneis;
EXOD|38|7|induxitque in circulos, qui in lateribus altaris eminebant. Ipsum autem altare non erat solidum, sed cavum ex tabulis et intus vacuum.
EXOD|38|8|Fecit et labrum aeneum cum basi sua de speculis mulierum, quae excubabant in ostio tabernaculi conventus.
EXOD|38|9|Fecit et atrium, in cuius australi plaga erant tentoria de bysso retorta cubitorum centum;
EXOD|38|10|columnae aeneae viginti cum basibus suis; unci columnarum et anuli earum argentei.
EXOD|38|11|Aeque ad septentrionalem plagam tentoria, columnae basesque et unci anulique columnarum eiusdem mensurae et operis ac metalli erant.
EXOD|38|12|In ea vero plaga, quae ad occidentem respicit, fuerunt tentoria cubitorum quinquaginta, columnae decem cum basibus suis; et unci columnarum anulique earum argentei.
EXOD|38|13|Porro contra orientem quinquaginta cubitorum paravit tentoria,
EXOD|38|14|e quibus quindecim cubitos columnarum trium cum basibus suis unum tenebat latus;
EXOD|38|15|et in parte altera ­ quia inter utraque introitum tabernaculi fecit ­ quindecim aeque cubitorum erant tentoria columnaeque tres et bases totidem.
EXOD|38|16|Cuncta atrii tentoria in circuitu ex bysso retorta texuerat.
EXOD|38|17|Bases columnarum fuere aeneae, unci autem earum et anuli earum argentei et capita earum vestivit argento et omnes columnas atrii cinxit anulis argenteis.
EXOD|38|18|Et in introitu eius opere plumario fecit velum ex hyacintho, purpura, cocco ac bysso retorta; quod habebat viginti cubitos in longitudine, altitudo vero quinque cubitorum erat iuxta mensuram, quam cuncta atrii tentoria habebant.
EXOD|38|19|Columnae autem in ingressu fuere quattuor cum basibus aeneis, uncis argenteis; capitaque et anulos earum vestivit argento.
EXOD|38|20|Paxillos quoque habitaculi et atrii per gyrum fecit aeneos.
EXOD|38|21|Hic est census habitaculi, habitaculi testimonii, qui recensitus est iuxta praeceptum Moysi ministerio Levitarum per manum Ithamar filii Aaron sacerdotis.
EXOD|38|22|Beseleel filius Uri filii Hur de tribu Iudae fecit cuncta, quae praeceperat Dominus Moysi,
EXOD|38|23|iuncto sibi socio Ooliab filio Achisamech de tribu Dan fabro et polymitario atque plumario ex hyacintho, purpura, cocco et bysso.
EXOD|38|24|Omne aurum, quod expensum est in opere sanctuarii et quod oblatum est in donariis, viginti novem talentorum fuit et septingentorum triginta siclorum ad mensuram sicli sanctuarii.
EXOD|38|25|Argentum autem eorum, qui in congregatione recensiti sunt, centum talentorum fuit et mille septingentorum et septuaginta quinque siclorum ad mensuram sicli sanctuarii.
EXOD|38|26|Beca, id est dimidium sicli iuxta mensuram sicli sanctuarii, dedit quisquis transit ad censum a viginti annis et supra, de sescentis tribus milibus et quingentis quinquaginta armatorum.
EXOD|38|27|De talentis centum argenti conflatae sunt bases sanctuarii et veli, singulis talentis per bases singulas supputatis.
EXOD|38|28|De mille autem septingentis et septuaginta quinque siclis fecit uncos columnarum et vestivit capita earum et cinxit eas argento.
EXOD|38|29|Aeris quoque oblata sunt septuaginta talenta et duo milia et quadringenti sicli,
EXOD|38|30|ex quibus fecit bases in introitu tabernaculi conventus et altare aeneum cum craticula sua omniaque vasa, quae ad usum eius pertinent,
EXOD|38|31|et bases atrii tam in circuitu quam in ingressu eius et omnes paxillos habitaculi atque atrii per gyrum.
EXOD|39|1|De hyacintho vero et purpura, cocco ac bysso fecerunt vestes textas pro ministerio sanctuarii. Et fecerunt vestes sacras Aaron, sicut praecepit Dominus Moysi.
EXOD|39|2|Fecerunt igitur ephod de auro, hyacintho et purpura coccoque et bysso retorta
EXOD|39|3|opere polymitario tundentes bratteas aureas et extenuantes in fila, ut possent torqueri cum priorum colorum subtegmine.
EXOD|39|4|Fasciasque umerales fecerunt ei, cum quibus in utroque latere summitatum suarum copulabatur,
EXOD|39|5|et balteum, quo constringebatur ephod, eiusdem operis et unum cum eo ex auro, et hyacintho et purpura coccoque et bysso retorta, sicut praeceperat Dominus Moysi.
EXOD|39|6|Paraverunt et duos lapides onychinos, inclusos texturis aureis et sculptos arte gemmaria nominibus filiorum Israel;
EXOD|39|7|posueruntque eos in fasciis umeralibus ephod, lapides memorialis filiorum Israel, sicut praeceperat Dominus Moysi.
EXOD|39|8|Fecerunt et pectorale opere polymito iuxta opus ephod ex auro, hyacintho, purpura coccoque et bysso retorta,
EXOD|39|9|quadrangulum duplex mensurae palmi.
EXOD|39|10|Et posuerunt in eo gemmarum ordines quattuor: in primo versu erat sardius, topazius, smaragdus;
EXOD|39|11|in secundo carbunculus, sapphirus et iaspis;
EXOD|39|12|in tertio hyacinthus, achates et amethystus;
EXOD|39|13|in quarto chrysolithus, onychinus et beryllus: inclusi textura aurea per ordines suos.
EXOD|39|14|Ipsique lapides duodecim sculpti erant nominibus duodecim tribuum Israel, singuli per nomina singulorum.
EXOD|39|15|Fecerunt in pectorali catenulas quasi funiculos opus tortile de auro purissimo
EXOD|39|16|et duos margines aureos totidemque anulos aureos. Porro duos anulos posuerunt in utraque summitate pectoralis;
EXOD|39|17|duos funiculos aureos inseruerunt anulis, qui in pectoralis angulis eminebant.
EXOD|39|18|Duas summitates amborum funiculorum colligaverunt duobus marginibus in fasciis umeralibus ephod in parte eius anteriore.
EXOD|39|19|Et fecerunt duos anulos aureos et posuerunt super duas summitates pectoralis in eius margine interiore contra ephod, sicut praecepit Dominus Moysi.
EXOD|39|20|Feceruntque duos anulos aureos, quos posuerunt in duabus fasciis umeralibus ephod deorsum in latere eius anteriore secus iuncturam eius super balteum ephod.
EXOD|39|21|Et strinxerunt pectorale anulis eius ad anulos ephod vitta hyacinthina, ut esset super balteum ephod, ne amoveretur ab ephod, sicut praecepit Dominus Moysi.
EXOD|39|22|Fecerunt quoque pallium ephod opere textili totum hyacinthinum
EXOD|39|23|et capitium in medio eius supra oramque per gyrum sicut in capitio loricae;
EXOD|39|24|deorsum autem ad pedes mala punica ex hyacintho, purpura, cocco ac bysso retorta
EXOD|39|25|et tintinnabula de auro purissimo, quae posuerunt inter malogranata in inferiore parte pallii per gyrum,
EXOD|39|26|ut sit tintinnabulum inter singula mala punica, quibus ornatus incedebat pontifex, quando ministerio fungebatur, sicut praeceperat Dominus Moysi.
EXOD|39|27|Fecerunt et tunicas byssinas opere textili Aaron et filiis eius
EXOD|39|28|et tiaram et ornatum mitrarum ex bysso, feminalia quoque linea ex bysso retorta,
EXOD|39|29|cingulum vero de bysso retorta, hyacintho, purpura ac cocco, arte plumaria, sicut praeceperat Dominus Moysi.
EXOD|39|30|Fecerunt et laminam diadema sanctitatis de auro purissimo; scripseruntque in ea opere caelatoris: " Sanctum Domino ";
EXOD|39|31|et strinxerunt eam desuper cum tiara vitta hyacinthina, sicut praeceperat Dominus Moysi.
EXOD|39|32|Perfectum est igitur omne opus habitaculi et tabernaculi conventus; feceruntque filii Israel cuncta, quae praeceperat Dominus Moysi: sic fecerunt.
EXOD|39|33|Et obtulerunt habitaculum et tabernaculum et universam supellectilem, fibulas, tabulas, vectes, columnas ac bases,
EXOD|39|34|opertorium de pellibus arietum rubricatis et operimentum de pellibus delphini, velum,
EXOD|39|35|arcam testimonii, vectes, propitiatorium,
EXOD|39|36|mensam cum vasis suis et propositionis panibus,
EXOD|39|37|candelabrum ex auro puro, lucernas in ordine earum et utensilia earum cum oleo candelabri,
EXOD|39|38|altare aureum et unguentum et thymiama ex aromatibus et velum in introitu tabernaculi,
EXOD|39|39|altare aeneum, craticulam aeneam, vectes et vasa eius omnia, labrum cum basi sua,
EXOD|39|40|tentoria atrii et columnas cum basibus suis, velum in introitu atrii funiculosque illius et paxillos. Nihil ex vasis defuit, quae in ministerium habitaculi in tabernaculo conventus iussa sunt fieri.
EXOD|39|41|Vestes quoque textas, quibus sacerdotes utuntur in sanctuario, et vestes sacras Aaron sacerdotis et vestes filiorum eius
EXOD|39|42|obtulerunt filii Israel, sicut praeceperat Dominus Moysi.
EXOD|39|43|Quae postquam Moyses cuncta vidit completa, benedixit eis.
EXOD|40|1|Locutusque est Dominus ad Moysen dicens:
EXOD|40|2|" Mense pri mo, die prima mensis eriges habitaculum, tabernaculum conventus,
EXOD|40|3|et pones in eo arcam testimonii, abscondes illam velo;
EXOD|40|4|et, illata mensa, pones super eam, quae rite praecepta sunt. Candelabrum stabit cum lucernis suis
EXOD|40|5|et altare aureum, in quo adoletur incensum, coram arca testimonii. Velum in introitu habitaculi pones,
EXOD|40|6|et ante tabernaculum conventus altare holocausti,
EXOD|40|7|et labrum inter altare et tabernaculum conventus et implebis illud aqua.
EXOD|40|8|Circumdabisque atrium tentoriis et pones velum in porta eius.
EXOD|40|9|Et, assumpto unctionis oleo, unges habitaculum et omnia, quae in eo sunt, et consecrabis illud cum vasis suis, et erit sanctum.
EXOD|40|10|Unges quoque altare holocausti et omnia vasa eius et consecrabis altare, et erit sanctum sanctorum.
EXOD|40|11|Et unges labrum cum basi sua et consecrabis illud.
EXOD|40|12|Applicabisque Aaron et filios eius ad fores tabernaculi conventus; et lotos aqua
EXOD|40|13|indues Aaron sanctis vestibus, unges et consecrabis eum, ut mihi sacerdotio fungatur;
EXOD|40|14|filios eius applicabis et vesties eos tunicis
EXOD|40|15|et unges eos, sicut unxisti patrem eorum, ut mihi sacerdotio fungantur, et unctio eorum erit eis in sacerdotium sempiternum in generationibus eorum ".
EXOD|40|16|Fecitque Moyses omnia, quae praeceperat ei Dominus: sic fecit.
EXOD|40|17|Igitur mense primo anni secundi, prima die mensis collocatum est habitaculum.
EXOD|40|18|Erexitque Moyses illud et posuit bases ac tabulas et vectes statuitque columnas
EXOD|40|19|et expandit tentorium super habitaculum, imposito desuper operimento, sicut Dominus imperaverat Moysi.
EXOD|40|20|Sumpsit et posuit testimonium in arca et, subditis infra vectibus, posuit propitiatorium desuper.
EXOD|40|21|Cumque intulisset arcam in habitaculum, appendit ante eam velum, sicut iusserat Dominus Moysi.
EXOD|40|22|Posuit et mensam in tabernaculo conventus ad plagam septentrionalem extra velum,
EXOD|40|23|ordinatis coram propositionis panibus, sicut praeceperat Dominus Moysi.
EXOD|40|24|Posuit et candelabrum in tabernaculo conventus e regione mensae in parte australi,
EXOD|40|25|locatis per ordinem lucernis, sicut praeceperat Dominus Moysi.
EXOD|40|26|Posuit et altare aureum in tabernaculo conventus coram propitiatorio
EXOD|40|27|et adolevit super eo incensum aromatum, sicut iusserat Dominus Moysi.
EXOD|40|28|Posuit et velum in introitu habitaculi
EXOD|40|29|et altare holocausti in vestibulo habitaculi, tabernaculi conventus, offerens in eo holocaustum et sacrificium, sicut Dominus imperaverat Moysi.
EXOD|40|30|Labrum quoque statuit inter tabernaculum conventus et altare implens illud aqua;
EXOD|40|31|laveruntque Moyses et Aaron ac filii eius manus suas et pedes,
EXOD|40|32|cum ingrederentur tabernaculum conventus et accederent ad altare, sicut praeceperat Dominus Moysi.
EXOD|40|33|Erexit et atrium per gyrum habitaculi et altaris, ducto in introitu eius velo. Sic complevit opus.
EXOD|40|34|Et operuit nubes tabernaculum conventus, et gloria Domini implevit habitaculum.
EXOD|40|35|Nec poterat Moyses ingredi tabernaculum conventus, quia habitavit nubes super illud, et gloria Domini replevit habitaculum.
EXOD|40|36|Si quando nubes de tabernaculo ascendebat, proficiscebantur filii Israel in omnibus stationibus suis;
EXOD|40|37|si autem non ascendebat nubes, non proficiscebantur usque in diem, quo levabatur.
EXOD|40|38|Nubes quippe Domini incubabat per diem habitaculo, et ignis in nocte, ante oculos universae domus Israel per cunctas mansiones suas." "
LEV|1|1|Vocavit autem Moysen et locu tus est ei Dominus de tabernacu lo conventus dicens:
LEV|1|2|" Loquere filiis Israel et dices ad eos: Homo, qui obtulerit ex vobis hostiam Domino de animalibus domesticis, de bobus et pecoribus offerens victimas,
LEV|1|3|si holocaustum fuerit eius oblatio de armento, masculum immaculatum offeret ad ostium tabernaculi conventus ad placandum sibi Dominum;
LEV|1|4|ponetque manum super caput hostiae, et acceptabilis erit atque in expiationem eius proficiens.
LEV|1|5|Immolabitque vitulum coram Domino, et offerent filii Aaron sacerdotes sanguinem eius aspergentes per altaris circuitum, quod est ante ostium tabernaculi conventus.
LEV|1|6|Detracta pelle, hostiam offerens in frusta concidet;
LEV|1|7|et filii Aaron sacerdotis ponent in altari ignem, strueque lignorum super ignem composita,
LEV|1|8|membra, quae caesa sunt, desuper ordinabunt, caput videlicet et adipem.
LEV|1|9|Intestina autem et crura offerens lavabit aqua adolebitque ea sacerdos super altare in holocaustum, incensum suavissimi odoris Domino.
LEV|1|10|Quod si de pecoribus eius oblatio est, de ovibus sive de capris holocaustum, masculum absque macula offeret;
LEV|1|11|immolabitque ad latus altaris, quod respicit ad aquilonem, coram Domino. Sanguinem vero illius aspergent contra altare filii Aaron sacerdotes per circuitum;
LEV|1|12|dividetque offerens membra, caput et adipem, et sacerdos imponet ea super ligna, quibus subest ignis in altari.
LEV|1|13|Intestina vero et crura lavabit offerens aqua, et oblata omnia adolebit sacerdos super altare: holocaustum est et incensum odoris suavissimi Domino.
LEV|1|14|Sin autem de avibus holocausti oblatio fuerit Domino, offeret de turturibus aut pullis columbae oblationem suam.
LEV|1|15|Et sacerdos afferet eam ad altare; retortum ad collum caput adolebit in altari, sanguisque eius exprimetur contra parietem altaris.
LEV|1|16|Vesiculam vero gutturis et plumas proiciet offerens prope altare ad orientalem plagam in loco, in quo cineres effundi solent;
LEV|1|17|confringetque eam inter alas, quas non secabit, et adolebit eam sacerdos super altare, lignis super ignem positis: holocaustum est et incensum suavissimi odoris Domino.
LEV|2|1|Anima cum obtulerit oblationem sacrificii farinae Domino, simila erit eius oblatio, fundetque super eam oleum et ponet tus
LEV|2|2|ac deferet ad filios Aaron sacerdotes, tolletque ex eo pugillum plenum similae et olei ac totum tus, et sacerdos adolebit memoriale super altare, incensum odoris suavissimi Domino.
LEV|2|3|Quod autem reliquum fuerit de sacrificio, erit Aaron et filiorum eius: sanctum sanctorum de incensis Domini.
LEV|2|4|Cum autem obtuleris sacrificium similae coctum in clibano: de simila erunt panes, scilicet absque fermento conspersi oleo et lagana azyma oleo lita;
LEV|2|5|si oblatio tua fuerit de sartagine, simila erit, conspersa oleo et absque fermento;
LEV|2|6|divides eam minutatim et fundes super eam oleum: oblatio similae est.
LEV|2|7|Sin autem de frixorio fuerit sacrificium, aeque simila oleo conspergetur.
LEV|2|8|Et deferes oblationem ex his Domino factam tradens manibus sacerdotis,
LEV|2|9|qui afferet eam ad altare, tollet memoriale de sacrificio et adolebit super altare: incensum odoris suavissimi Domino.
LEV|2|10|Quidquid autem reliquum est, erit Aaron et filiorum eius: sanctum sanctorum de incensis Domini.
LEV|2|11|Omnis oblatio similae, quam offeretis Domino, absque fermento fiet, quia nihil fermenti ac mellis adolebitis incensum Domino.
LEV|2|12|Primitias tantum eorum offeretis tamquam munera Domino; super altare vero non ponentur in odorem suavitatis.
LEV|2|13|Quidquid obtuleris sacrificii, similae sale condies nec auferes sal foederis Dei tui de sacrificio tuo: in omni oblatione tua offeres sal.
LEV|2|14|Sin autem obtuleris munus primarum frugum tuarum Domino, spicas tostas igni et grana fracta farris recentis offeres in sacrificium primarum frugum tuarum
LEV|2|15|fundens supra oleum et tus imponens: similae oblatio est.
LEV|2|16|De qua adolebit sacerdos tamquam memoriale partem farris fracti et olei ac totum tus.
LEV|3|1|Quod si hostia pacificorum fue rit eius oblatio et de bobus vo luerit offerre marem sive feminam, immaculata offeret coram Domino.
LEV|3|2|Ponetque manum super caput victimae suae, quam immolabit ad ostium tabernaculi conventus, fundentque filii Aaron sacerdotes sanguinem per circuitum altaris
LEV|3|3|et offerent de hostia pacificorum tamquam incensum Domino adipem, qui operit vitalia, et quidquid pinguedinis eis adhaeret,
LEV|3|4|duos renes cum adipe, quo teguntur iuxta ilia, et reticulum iecoris, quem iuxta renes, auferet.
LEV|3|5|Adolebuntque ea filii Aaron in altari super holocausto, quod est super lignis et igne: incensum suavissimi odoris Domino.
LEV|3|6|Si vero de pecoribus fuerit Domino eius oblatio, pacificorum scilicet hostia, sive masculum sive feminam obtulerit, immaculata erunt.
LEV|3|7|Si agnum obtulerit coram Domino,
LEV|3|8|ponet manum super caput victimae suae, quam immolabit coram tabernaculo conventus; fundentque filii Aaron sanguinem eius per altaris circuitum;
LEV|3|9|et offeret de pacificorum hostia incensum Domino adipem et caudam totam, quam iuxta tergum, auferet, et pinguedinem, quae operit ventrem, atque universum adipem, qui vitalibus adhaeret,
LEV|3|10|et utrumque renunculum cum adipe, qui est iuxta ilia, reticulumque iecoris, quem iuxta renunculos, auferet.
LEV|3|11|Et adolebit ea sacerdos super altare: panis et incensum Domino.
LEV|3|12|Si capra fuerit eius oblatio, offeret eam coram Domino,
LEV|3|13|ponet manum suam super caput eius immolabitque eam coram tabernaculo conventus. Et fundent filii Aaron sanguinem eius per altaris circuitum,
LEV|3|14|tolletque ex ea oblationem suam, incensum Domino, adipem scilicet, qui operit ventrem, et universum, qui vitalibus adhaeret,
LEV|3|15|duos renunculos cum adipe, qui est super eos iuxta ilia, et reticulum iecoris, quem iuxta renunculos, auferet;
LEV|3|16|adolebitque ea sacerdos super altare: panis et incensum suavissimi odoris omnis adeps Domino.
LEV|3|17|Iure perpetuo in generationibus et cunctis habitaculis vestris, nec adipem nec sanguinem omnino comedetis ".
LEV|4|1|Locutusque est Dominus ad Moysen dicens:
LEV|4|2|" Loquere filiis Israel: Anima cum peccaverit per ignorantiam et de universis mandatis Domini, quae praecepit ut non fierent, quippiam fecerit,
LEV|4|3|si sacerdos, qui est unctus, peccaverit, delinquere faciens populum, offeret pro peccato suo vitulum immaculatum Domino sacrificium pro peccato;
LEV|4|4|et adducet illum ad ostium tabernaculi conventus coram Domino ponetque manum super caput eius et immolabit eum coram Domino.
LEV|4|5|Hauriet quoque sacerdos unctus de sanguine vituli inferens illum in tabernaculum conventus;
LEV|4|6|cumque intinxerit digitum in sanguinem, asperget eo septies coram Domino contra velum sanctuarii;
LEV|4|7|ponetque de eodem sanguine super cornua altaris thymiamatis gratissimi coram Domino, quod est in tabernaculo conventus; omnem autem reliquum sanguinem fundet in basim altaris holocausti in introitu tabernaculi.
LEV|4|8|Et omnem adipem vituli pro peccato auferet tam eum, qui operit vitalia, quam omnem, qui vitalibus adhaeret,
LEV|4|9|duos renunculos et adipem, qui est super eos iuxta ilia, et reticulum iecoris, quem iuxta renunculos, auferet,
LEV|4|10|sicut aufertur de vitulo hostiae pacificorum; et adolebit ea sacerdos super altare holocausti.
LEV|4|11|Pellem vero et omnes carnes cum capite et pedibus et intestinis et fimo,
LEV|4|12|totum vitulum efferet extra castra in locum mundum, ubi cineres effundi solent; incendetque eum super lignorum struem igne: in loco effusorum cinerum cremabitur.
LEV|4|13|Quod si omnis coetus Israel ignoraverit, et res abscondita fuerit ab oculis congregationis, feceritque quod contra mandatum Domini est et deliquerit,
LEV|4|14|et postea intellexerit peccatum suum, offeret congregatio vitulum pro peccato adducetque eum ad ostium tabernaculi conventus.
LEV|4|15|Et ponent seniores coetus populi manus super caput eius coram Domino, immolatoque vitulo in conspectu Domini,
LEV|4|16|inferet sacerdos, qui unctus est, de sanguine eius in tabernaculum conventus,
LEV|4|17|tincto digito aspergens septies contra velum;
LEV|4|18|ponetque de eodem sanguine in cornibus altaris, quod est coram Domino in tabernaculo conventus. Reliquum autem sanguinem fundet iuxta basim altaris holocaustorum, quod est in ostio tabernaculi conventus;
LEV|4|19|omnemque eius adipem tollet et adolebit super altare.
LEV|4|20|Sic faciens et de hoc vitulo quomodo fecit de vitulo pro peccato; sic faciet ei. Expiante eos sacerdote, propitius erit Dominus.
LEV|4|21|Ipsum autem vitulum efferet extra castra atque comburet sicut et priorem vitulum: sacrificium pro peccato est congregationis.
LEV|4|22|Si peccaverit princeps et fecerit unum ex omnibus per ignorantiam, quod Domini Dei sui lege prohibetur, deliqueritque,
LEV|4|23|aut indicatum ei fuerit peccatum suum, offeret hostiam Domino hircum de capris immaculatum
LEV|4|24|ponetque manum suam super caput eius et immolabit eum in loco, ubi solet mactari holocaustum coram Domino: sacrificium pro peccato est.
LEV|4|25|Et tinguat sacerdos digitum in sanguine hostiae pro peccato ponetque super cornua altaris holocausti et reliquum fundet ad basim eius.
LEV|4|26|Adipem vero adolebit supra, sicut in victimis pacificorum fieri solet; expiabitque eum a peccato eius, ac dimittetur ei.
LEV|4|27|Quod si peccaverit anima per ignorantiam de populo terrae, ut faciat quidquam ex his, quae Domini lege prohibentur, atque delinquat,
LEV|4|28|aut indicatum ei fuerit peccatum suum, offeret capram immaculatam;
LEV|4|29|ponetque manum super caput hostiae pro peccato et immolabit eam in loco holocausti.
LEV|4|30|Tolletque sacerdos de sanguine in digito suo et ponet super cornua altaris holocausti et reliquum fundet ad basim eius.
LEV|4|31|Omnem autem auferens adipem, sicut auferri solet de victimis pacificorum, adolebit super altare in odorem suavitatis Domino, expiabitque eum, et propitius erit Dominus.
LEV|4|32|Sin autem de ovibus obtulerit victimam pro peccato, adducet agnam immaculatam;
LEV|4|33|ponet manum super caput eius et immolabit eam in loco, ubi solent holocaustorum caedi hostiae.
LEV|4|34|Sumetque sacerdos de sanguine eius digito suo et ponens super cornua altaris holocausti reliquum fundet ad basim eius.
LEV|4|35|Omnem quoque auferens adipem, sicut auferri solet adeps agni, qui immolatur pro pacificis, cremabit in altari super incensis Domini; expiabitque eum et peccatum eius, et dimittetur illi.
LEV|5|1|Si peccaverit anima et audiverit vocem iurantis testisque fuerit, quod aut ipse vidit aut comperit, si non indicaverit, iniquitatem portabit;
LEV|5|2|vel si anima tetigerit aliquid immundum, sive cadaver bestiae sit aut iumenti vel reptilis, et absconditum fuerit ab eo, ipse immundus et reus erit;
LEV|5|3|aut si tetigerit quidquam de immunditia hominis iuxta omnem impuritatem, qua pollui solet, absconditumque fuerit ab eo, sed ipse cognoverit postea, subiacebit delicto;
LEV|5|4|aut si anima temere iuraverit et protulerit labiis suis, ut vel male quid faceret vel bene iuxta omnia, quae homines temere iurant, absconditumque fuerit ab eo, sed ipse postea intellexerit, delicto subiacebit;
LEV|5|5|si ergo reus factus fuerit uno ex istis, confiteatur peccatum suum
LEV|5|6|et offerat Domino sacrificium delicti pro peccato suo agnam de gregibus sive capram ut sacrificium pro peccato; expiabitque eum sacerdos a peccato eius.
LEV|5|7|Sin autem non potuerit offerre pecus, offerat ut sacrificium pro delicto duos turtures vel duos pullos columbarum Domino: unum in sacrificium pro peccato et alterum in holocaustum;
LEV|5|8|dabitque eos sacerdoti, qui primum offerens ut sacrificium pro peccato retorquebit caput eius ad pennulas, ita ut collo haereat et non penitus abrumpatur;
LEV|5|9|et asperget de sanguine eius parietem altaris; quidquid autem reliquum fuerit, faciet destillare ad fundamentum eius: sacrificium pro peccato est.
LEV|5|10|Alterum vero adolebit holocaustum, ut fieri solet; expiabitque eum sacerdos a peccato eius, et dimittetur ei.
LEV|5|11|Quod si non quiverit manus eius offerre duos turtures aut duos pullos columbarum, offeret pro peccato suo similae partem ephi decimam in sacrificium pro peccato; non mittet in eam oleum, nec turis aliquid imponet, quia sacrificium pro peccato est.
LEV|5|12|Tradetque eam sacerdoti, qui, plenum ex toto pugillum in memoriale hauriens, cremabit in altari super incensis Domini: sacrificium pro peccato est.
LEV|5|13|Et expiabit eum sacerdos et peccatum eius in uno ex his casibus, et propitius erit Dominus. Reliquam vero partem sacerdos habebit sicut in oblatione similae ".
LEV|5|14|Locutus est Dominus ad Moysen dicens:
LEV|5|15|" Anima, si praevaricans per errorem in his, quae Domino sunt sanctificata, peccaverit, offeret sacrificium pro delicto arietem immaculatum de gregibus iuxta aestimationem argenti siclorum pondere sanctuarii in paenitentiam;
LEV|5|16|ipsumque, quod intulit damni, restituet et quintam partem ponet supra tradens sacerdoti, qui expiabit eum offerens arietem, et dimittetur ei.
LEV|5|17|Anima, si peccaverit per ignorantiam feceritque unum ex his, quae Domini lege prohibentur, et peccati rea portaverit iniquitatem suam,
LEV|5|18|offeret arietem immaculatum de gregibus iuxta aestimationem sacerdoti, qui expiabit eum ab eo, quod nesciens fecerit, et dimittetur ei:
LEV|5|19|sacrificium pro delicto est, delinquens deliquit in Dominum ".
LEV|5|20|Locutus est Dominus ad Moysen dicens:
LEV|5|21|" Anima, quae peccaverit et, contempto Domino, negaverit proximo suo depositum, quod fidei eius creditum fuerat, vel vi aliquid extorserit aut calumniam fecerit,
LEV|5|22|sive rem perditam invenerit et infitians insuper peierarit in uno ex omnibus, in quibus peccare solent homines,
LEV|5|23|si quis sic peccaverit et deliquerit, reddet omnia, quae per rapinam vel calumniam abstulerit vel deposita retinuerit vel perdita invenerit
LEV|5|24|vel de quibus peierarit, et restituet integra et quintam insuper addet partem domino, cui damnum intulerat, in die sacrificii pro delicto.
LEV|5|25|Sacrificium pro delicto offeret Domino: arietem immaculatum de grege iuxta aestimationem;
LEV|5|26|qui expiabit eum coram Domino, et dimittetur illi pro singulis, quae faciendo peccaverit ".
LEV|6|1|Locutus est Dominus ad Moysen dicens:
LEV|6|2|" Praecipe Aaron et filiis eius: Haec est lex holocausti: cremabitur in foco altaris tota nocte usque mane; ignis altaris in eo ardebit.
LEV|6|3|Vestietur sacerdos tunica et feminalibus lineis super verecunda sua; tolletque cineres, quos vorans ignis exussit, et ponet iuxta altare.
LEV|6|4|Porro spoliabitur prioribus vestimentis; indutusque aliis efferet cineres extra castra in locum mundum.
LEV|6|5|Ignis autem in altari semper ardebit, non exstinguetur, quem nutriet sacerdos subiciens ligna mane per singulos dies et, imposito holocausto, desuper adolebit adipes pacificorum.
LEV|6|6|Ignis est iste perpetuus, qui numquam deficiet in altari.
LEV|6|7|Haec est lex sacrificii similae, quod offerent filii Aaron coram Domino et coram altare:
LEV|6|8|tollet sacerdos ex eo pugillum similae, quae conspersa est oleo, et totum tus, quod super similam positum est; adolebitque illud in altari in odorem suavissimum, memoriale Domino.
LEV|6|9|Reliquam autem partem similae comedet Aaron cum filiis suis, et panis absque fermento comedetur in loco sancto; in atrio tabernaculi conventus comedent illam.
LEV|6|10|Ideo autem non coquetur fermentata, quia ut partem eorum dedi illam ex incensis meis: sanctum sanctorum est, sicut sacrificium pro peccato atque pro delicto;
LEV|6|11|mares tantum stirpis Aaron comedent illud. Legitimum sempiternum est in generationibus vestris de incensis Domini; omnis, qui tetigerit illa, sanctificabitur ".
LEV|6|12|Et locutus est Dominus ad Moysen dicens:
LEV|6|13|" Haec est oblatio Aaron et filiorum eius, quam offerre debent Domino in die unctionis ipsius: decimam partem ephi offerent similae in sacrificio sempiterno medium eius mane et medium vespere;
LEV|6|14|quae in sartagine oleo conspersa frigetur. Afferes eam calidam et offeres divisam minutatim, sacrificium in odorem suavissimum Domino.
LEV|6|15|Sacerdos unctus, qui patri iure successerit, faciet illud. Legitimum sempiternum: Domino tota cremabitur;
LEV|6|16|omne enim sacrificium similae sacerdotum igne consumetur, nec quisquam comedet ex eo ".
LEV|6|17|Locutus est Dominus ad Moysen dicens:
LEV|6|18|" Loquere Aaron et filiis eius: Ista est lex sacrificii pro peccato: in loco, ubi mactatur holocaustum, mactabitur coram Domino: sanctum sanctorum est.
LEV|6|19|Sacerdos, qui offert, comedet illud in loco sancto, in atrio tabernaculi conventus.
LEV|6|20|Quidquid tetigerit carnes eius, sanctificabitur: si de sanguine illius vestis fuerit aspersa, lavabitur in loco sancto;
LEV|6|21|vas autem fictile, in quo coctum est, confringetur; quod si vas aeneum fuerit, defricabitur et lavabitur aqua.
LEV|6|22|Omnis masculus de genere sacerdotali vescetur carnibus eius, quia sanctum sanctorum est.
LEV|6|23|Omne autem sacrificium pro peccato, de cuius sanguine infertur in tabernaculum conventus ad expiandum in sanctuario, non comedetur, sed comburetur igni.
LEV|7|1|Haec quoque est lex sacrificii pro delicto: sanctum sanctorum est,
LEV|7|2|idcirco, ubi immolatur holocaustum, mactabitur et victima pro delicto; sanguis eius per gyrum fundetur altaris.
LEV|7|3|Omnemque adipem offeret ex ea, caudam scilicet et adipem, qui operit vitalia,
LEV|7|4|duos renunculos et pinguedinem, quae super eos iuxta ilia est, reticulumque iecoris, quem iuxta renunculos, auferet;
LEV|7|5|et adolebit ea sacerdos super altare ut incensum Domino: sacrificium pro delicto est.
LEV|7|6|Omnis masculus de sacerdotali genere in loco sancto vescetur his carnibus, quia sanctum sanctorum est.
LEV|7|7|Sicut sacrificium pro peccato, ita et sacrificium pro delicto, utriusque hostiae lex una est; ad sacerdotem, qui eam obtulerit, pertinebit.
LEV|7|8|Sacerdos, qui offert holocaustum cuiusdam viri, habebit pellem victimae,
LEV|7|9|et omne sacrificium similae, quod coquitur in clibano, et, quidquid in frixorio vel in sartagine praeparatur, eius erit sacerdotis, a quo offertur;
LEV|7|10|et omne sacrificium similae sive oleo conspersum sive aridum fuerit, cunctis filiis Aaron aequa mensura per singulos dividetur.
LEV|7|11|Haec est lex hostiae pacificorum quae offertur Domino;
LEV|7|12|si pro gratiarum actione fuerit oblatio, offerent panes absque fermento conspersos oleo et lagana azyma uncta oleo coctamque similam ut collyridas olei admixtione conspersas,
LEV|7|13|panes quoque fermentatos cum hostia pacificorum pro gratiarum actione,
LEV|7|14|ex quibus unus offeretur munus Domino et erit sacerdotis, qui fundet hostiae sanguinem.
LEV|7|15|Cuius carnes eadem comedentur die, nec remanebit ex eis quidquam usque mane.
LEV|7|16|Si voto vel sponte quisquam obtulerit hostiam, eadem similiter edetur die; sed et si quid in crastinum remanserit, vesci licitum est;
LEV|7|17|quidquid autem tertius invenerit dies, ignis absumet.
LEV|7|18|Si quis de carnibus victimae pacificorum die tertio comederit, irrita fiet oblatio nec proderit offerenti; quin potius, quaecumque anima tali se edulio contaminarit, praevaricationis rea erit.
LEV|7|19|Caro, quae aliquid tetigerit immundum, non comedetur, sed comburetur igni; ceterum carne, qui fuerit mundus, vescetur.
LEV|7|20|Anima polluta, quae ederit de carnibus hostiae pacificorum, quae oblata est Domino, peribit de populis suis;
LEV|7|21|et, quae tetigerit immunditiam hominis vel iumenti, sive omnis rei abominabilis, quae polluere potest, et comederit de huiuscemodi carnibus, interibit de populis suis ".
LEV|7|22|Locutusque est Dominus ad Moysen dicens:
LEV|7|23|" Loquere filiis Israel: Adipem bovis et ovis et caprae non comedetis.
LEV|7|24|Adipem cadaveris morticini et eius animalis, quod a bestia laceratum est, habebitis in usus varios, sed non comedetis.
LEV|7|25|Si quis adipem, qui offertur in incensum Domini, comederit, peribit de populo suo.
LEV|7|26|Sanguinem quoque omnis animalis non sumetis in cibo, tam de avibus quam de pecoribus;
LEV|7|27|omnis anima, quae ederit sanguinem, peribit de populis suis ".
LEV|7|28|Locutus est Dominus ad Moysen dicens:
LEV|7|29|" Loquere filiis Israel: Qui offert victimam pacificorum Domino, afferat oblationem suam Domino de victima pacificorum.
LEV|7|30|Tenebit manibus incensa Domini, adipem scilicet et pectusculum afferet; pectusculum, ut elevetur coram Domino.
LEV|7|31|Et sacerdos adolebit adipem super altare; pectusculum autem erit Aaron et filiorum eius.
LEV|7|32|Armus quoque dexter de pacificorum hostiis cedet in munus sacerdotis.
LEV|7|33|Qui de filiis Aaron obtulerit sanguinem et adipem victimae pacificorum, ipse habebit armum dextrum in portione sua;
LEV|7|34|pectusculum enim elationis et armum donationis tuli a filiis Israel de hostiis eorum pacificis et dedi Aaron sacerdoti ac filiis eius, lege perpetua, ab omni populo Israel ".
LEV|7|35|Haec est portio Aaron et filiorum eius de incensis Domini die, qua applicavit eos, ut sacerdotio fungerentur;
LEV|7|36|et quae praecepit dari eis Dominus a filiis Israel die, qua unxit eos, religione perpetua in generationibus eorum.
LEV|7|37|Ista est lex holocausti et oblationis similae et sacrificii pro peccato atque delicto et pro consecratione et pacificorum victimis,
LEV|7|38|quam constituit Dominus Moysi in monte Sinai, quando mandavit filiis Israel, ut offerrent oblationes suas Domino in deserto Sinai.
LEV|8|1|Locutusque est Dominus ad Moysen dicens:
LEV|8|2|" Tolle Aaron cum filiis suis, vestes eorum et unctionis oleum, vitulum pro peccato, duos arietes, canistrum cum azymis;
LEV|8|3|et congregabis omnem coetum ad ostium tabernaculi conventus ".
LEV|8|4|Fecit Moyses, ut Dominus imperarat; congregatoque omni coetu ante fores tabernaculi conventus,
LEV|8|5|ait: " Iste est sermo, quem iussit Dominus fieri ".
LEV|8|6|Statimque applicavit Aaron et filios eius. Cumque lavisset eos aqua,
LEV|8|7|vestivit pontificem subucula linea accingens eum balteo et induens tunica hyacinthina et desuper ephod imposuit,
LEV|8|8|quod astrinxit cingulo ephod firmiter; et imposuit ei pectorale, in quo dedit Urim et Tummim.
LEV|8|9|Cidari quoque texit caput et super eam contra frontem posuit laminam auream, diadema sanctum, sicut praeceperat Dominus Moysi.
LEV|8|10|Tulit et unctionis oleum, quo levit habitaculum cum omni supellectili sua et sanctificavit ea.
LEV|8|11|Cumque de eo aspersisset altare septem vicibus, unxit illud et omnia vasa eius labrumque cum basi sua sanctificavit oleo.
LEV|8|12|Quod fundens super caput Aaron, unxit eum et consecravit;
LEV|8|13|filios quoque eius applicatos vestivit subuculis lineis et cinxit balteo imposuitque mitras, ut iusserat Dominus Moysi.
LEV|8|14|Adduxit et vitulum pro peccato; cumque super caput eius posuissent Aaron et filii eius manus suas,
LEV|8|15|immolavit eum; et hauriens Moyses sanguinem tincto digito tetigit cornua altaris per gyrum et mundavit illud; fuditque reliquum sanguinem ad fundamenta eius et sanctificavit illud expiando.
LEV|8|16|Adipem autem, qui erat super vitalia, et reticulum iecoris duosque renunculos cum arvinulis suis adolevit super altare;
LEV|8|17|vitulum cum pelle, carnibus et fimo cremans extra castra, sicut praeceperat Dominus Moysi.
LEV|8|18|Attulit et arietem in holocaustum, super cuius caput cum imposuissent Aaron et filii eius manus suas,
LEV|8|19|immolavit eum et fudit sanguinem eius per altaris circuitum.
LEV|8|20|Ipsumque arietem in frusta concidens, caput eius et artus et adipem adolevit igni;
LEV|8|21|lotis prius intestinis et pedibus, totumque simul arietem adolevit super altare, eo quod esset holocaustum suavissimi odoris, incensum Domino, sicut praeceperat Dominus Moysi.
LEV|8|22|Attulit et arietem secundum in consecrationem sacerdotum; posueruntque super caput illius Aaron et filii eius manus suas.
LEV|8|23|Quem cum immolasset Moyses, sumens de sanguine tetigit extremum auriculae dextrae Aaron et pollicem manus eius dextrae, similiter et pedis.
LEV|8|24|Applicavit et filios Aaron; cumque de sanguine arietis immolati tetigisset extremum auriculae singulorum dextrae et pollices manus ac pedis dextri, reliquum fudit super altare per circuitum.
LEV|8|25|Tulitque adipem et caudam omnemque pinguedinem, quae operit intestina reticulumque iecoris, et duos renes cum adipibus suis et armo dextro.
LEV|8|26|Tollens autem de canistro azymorum, quod erat coram Domino, panem absque fermento et collyridam conspersam oleo laganumque posuit super adipes et armum dextrum,
LEV|8|27|tradens simul omnia super manus Aaron et filiorum eius. Qui, postquam levaverunt ea coram Domino,
LEV|8|28|rursum suscepta de manibus eorum adolevit in altari super holocausto, eo quod illa essent consecrationis oblatio, in odorem suavitatis: incensum erat Domino.
LEV|8|29|Tulit et pectusculum elevans illud coram Domino de ariete consecrationis in partem suam, sicut praeceperat Dominus Moysi.
LEV|8|30|Assumensque de unguento et sanguine, qui erat in altari, aspersit super Aaron et vestimenta eius et super filios illius ac vestes eorum.
LEV|8|31|Cumque sanctificasset eos in vestitu suo, praecepit eis dicens: " Coquite carnes ante fores tabernaculi et ibi comedite eas; panes quoque consecrationis edite, qui positi sunt in canistro, sicut mihi praeceptum est: "Aaron et filii eius comedent eos;
LEV|8|32|quidquid autem reliquum fuerit de carne et panibus, ignis absumet".
LEV|8|33|De ostio quoque tabernaculi conventus non exibitis septem diebus usque ad diem, quo complebitur tempus consecrationis vestrae; septem enim diebus finitur consecratio.
LEV|8|34|Sicut et impraesentiarum factum est, praecepit Dominus, ut fieret in expiationem eorum.
LEV|8|35|Die ac nocte manebitis in ostio tabernaculi conventus observantes observationem Domini, ne moriamini: sic enim mihi praeceptum est ".
LEV|8|36|Feceruntque Aaron et filii eius cuncta, quae locutus est Dominus per manum Moysi.
LEV|9|1|Facto autem octavo die, vocavit Moyses Aaron et filios eius ac maiores natu Israel dixitque ad Aaron:
LEV|9|2|" Tolle de armento vitulum pro peccato et arietem in holocaustum, utrumque immaculatum, et affer illos coram Domino.
LEV|9|3|Et ad filios Israel loqueris: "Tollite hircum pro peccato et vitulum atque agnum anniculos et sine macula in holocaustum,
LEV|9|4|bovem et arietem pro pacificis, et immolate eos coram Domino, et sacrificium similae oleo conspersae: hodie enim Dominus apparebit vobis" ".
LEV|9|5|Tulerunt ergo cuncta, quae iusserat Moyses, ad ostium tabernaculi conventus; ubi, cum omnis coetus accessisset et staret coram Domino,
LEV|9|6|ait Moyses: " Iste est sermo, quem praecepit Dominus: facite, et apparebit vobis gloria eius ".
LEV|9|7|Dixit et ad Aaron: " Accede ad altare et immola pro peccato tuo; offer holocaustum et expia te et populum. Et fac hostiam populi et expia eum, sicut praecepit Dominus ".
LEV|9|8|Statimque Aaron accedens ad altare immolavit vitulum pro peccato suo,
LEV|9|9|cuius sanguinem obtulerunt ei filii sui; in quo tinguens digitum tetigit cornua altaris et fudit residuum ad basim eius.
LEV|9|10|Adipemque et renunculos ac reticulum iecoris, quae sunt de sacrificio pro peccato, adolevit super altare, sicut praeceperat Dominus Moysi.
LEV|9|11|Carnes vero et pellem eius extra castra combussit igni.
LEV|9|12|Immolavit et holocausti victimam; obtuleruntque ei filii sui sanguinem eius, quem fudit per altaris circuitum.
LEV|9|13|Ipsam etiam hostiam in frusta concisam cum capite ei obtulerunt, quae omnia super altare cremavit igni;
LEV|9|14|lavit quoque aqua intestina cruraque et adolevit super holocausto in altari.
LEV|9|15|Et applicavit oblationem populi sumensque hircum pro peccato populi mactavit et obtulit in expiationem sicut priorem;
LEV|9|16|fecit quoque holocaustum secundum ritum
LEV|9|17|et addens sacrificium similae implevit manum ex illa et adolevit super altare praeter holocaustum matutinum.
LEV|9|18|Immolavit et bovem atque arietem, hostias pacificas populi; obtuleruntque ei filii sui sanguinem, quem fudit super altare in circuitu.
LEV|9|19|Adipes autem bovis et caudam arietis renunculosque cum adipibus suis et reticulum iecoris
LEV|9|20|posuerunt super pectora; cumque cremati essent adipes in altari,
LEV|9|21|pectora eorum et armos dextros Aaron elevavit coram Domino, sicut praeceperat Moyses.
LEV|9|22|Et elevans Aaron manus ad populum benedixit eis. Sicque, completis hostiis pro peccato et holocaustis et pacificis, descendit.
LEV|9|23|Ingressi autem Moyses et Aaron tabernaculum conventus et deinceps egressi benedixerunt populo. Apparuitque gloria Domini omni populo;
LEV|9|24|et ecce egressus ignis a Domino devoravit holocaustum et adipes, qui erant super altare. Quod cum vidissent turbae, exultaverunt ruentes in facies suas.
LEV|10|1|Arreptisque Nadab et Abiu filii Aaron turibulis, posue runt ignem et incensum desuper offerentes coram Domino ignem alienum, qui eis praeceptus non erat.
LEV|10|2|Egressusque ignis a Domino devoravit eos, et mortui sunt coram Domino.
LEV|10|3|Dixitque Moyses ad Aaron: " Hoc est, quod locutus est Dominus: "Sanctificabor in his, qui appropinquant mihi, et in conspectu omnis populi glorificabor" ". Quod audiens tacuit Aaron.
LEV|10|4|Vocatis autem Moyses Misael et Elisaphan filiis Oziel patrui Aaron, ait ad eos: " Ite et tollite fratres vestros de conspectu sanctuarii et asportate extra castra ".
LEV|10|5|Confestimque pergentes tulerunt eos, sicut iacebant vestitos subuculis suis, foras, ut sibi fuerat imperatum.
LEV|10|6|Locutus est Moyses ad Aaron et ad Eleazar atque Ithamar filios eius: " Comas vestras nolite excutere et vestimenta nolite scindere, ne moriamini, et super omnem coetum oriatur indignatio. Fratres vestri, omnis domus Israel, plangant incendium, quod Dominus suscitavit.
LEV|10|7|Vos autem non egredimini fores tabernaculi conventus, alioquin peribitis; oleum quippe unctionis Domini est super vos ". Qui fecerunt omnia iuxta praeceptum Moysi.
LEV|10|8|Dixit quoque Dominus ad Aaron:
LEV|10|9|" Vinum et omne, quod inebriare potest, non bibetis tu et filii tui, quando intratis tabernaculum conventus, ne moriamini ­ praeceptum est sempiternum in generationes vestras ­
LEV|10|10|et ut habeatis scientiam discernendi inter sanctum et profanum, inter pollutum et mundum,
LEV|10|11|doceatisque filios Israel omnia legitima mea, quae locutus est Dominus ad eos per manum Moysi ".
LEV|10|12|Locutusque est Moyses ad Aaron et ad Eleazar atque Ithamar filios eius, qui residui erant: " Tollite oblationem similae, quae remansit de incensis Domini, et comedite illam absque fermento iuxta altare, quia sanctum sanctorum est.
LEV|10|13|Comedetis autem in loco sancto, quia data est tibi et filiis tuis de incensis Domini, sicut praeceptum est mihi.
LEV|10|14|Pectusculum quoque elationis et armum donationis edetis in loco mundissimo, tu et filii tui ac filiae tuae tecum; tibi enim ac liberis tuis reposita sunt de hostiis pacificis filiorum Israel.
LEV|10|15|Armum et pectus cum incensis adipum afferent ad elationem coram Domino, et pertineant ad te et ad filios tuos lege perpetua, sicut praecepit Dominus ".
LEV|10|16|De hirco autem pro peccato cum quaereret Moyses, exustum repperit; iratusque contra Eleazar et Ithamar filios Aaron, qui remanserant, ait:
LEV|10|17|" Cur non comedistis sacrificium pro peccato in loco sancto? Quod sanctum sanctorum est, et datum vobis, ut portetis iniquitatem coetus in expiationem eorum in conspectu Domini;
LEV|10|18|praesertim cum de sanguine illius non sit illatum intra sancta, comedere eam debuistis in sanctuario, sicut praeceptum est mihi ".
LEV|10|19|Respondit Aaron: " Oblata est hodie victima pro peccato et holocaustum eorum coram Domino; mihi autem accidit, quod vides. Quomodo potui comedere eam et placere Domino? ".
LEV|10|20|Quod cum audisset Moyses, recepit satisfactionem.
LEV|11|1|Locutus est Dominus ad Moysen et Aaron dicens:
LEV|11|2|" Dicite filiis Israel: Haec sunt animalia, quae comedere debetis de cunctis animantibus terrae.
LEV|11|3|Omne, quod habet plene divisam ungulam et ruminat in pecoribus, comedetis.
LEV|11|4|Haec autem non comedetis ex ruminantibus vel dividentibus ungulam: camelum, quia ruminat quidem, sed non dividit ungulam, inter immunda reputabis;
LEV|11|5|hyracem, qui ruminat ungulamque non dividit, immundus est;
LEV|11|6|leporem quoque, nam et ipse ruminat, sed ungulam non dividit;
LEV|11|7|et suem, qui, cum ungulam plene dividat, non ruminat.
LEV|11|8|Horum carnibus non vescemini nec cadavera contingetis, quia immunda sunt vobis.
LEV|11|9|Haec sunt, quae gignuntur in aquis et vesci licitum est: omne, quod habet pinnulas et squamas, tam in mari quam in fluminibus et torrentibus, comedetis.
LEV|11|10|Quidquid autem pinnulas et squamas non habet, reptilium vel quorumlibet aliorum animalium, quae in aquis moventur, abominabile vobis
LEV|11|11|et execrandum erit; carnes eorum non comedetis et morticina vitabitis.
LEV|11|12|Cuncta, quae non habent pinnulas et squamas in aquis, polluta erunt vobis.
LEV|11|13|Haec sunt, quae de avibus comedere non debetis, et vitanda sunt vobis: aquilam et grypem et haliaeetum,
LEV|11|14|milvum ac vulturem iuxta genus suum
LEV|11|15|et omne corvini generis,
LEV|11|16|struthionem et noctuam et larum et accipitrem iuxta genus suum,
LEV|11|17|bubonem et mergulum et ibin,
LEV|11|18|cycnum et nyctocoracem et porphyrionem,
LEV|11|19|erodionem et charadrion iuxta genus suum, upupam quoque et vespertilionem.
LEV|11|20|Omne de volucribus, quod reptat super quattuor pedes, abominabile erit vobis.
LEV|11|21|Quidquid autem ambulat quidem super quattuor pedes, sed habet longiora retro crura, per quae salit super terram,
LEV|11|22|comedere debetis; ut est bruchus in genere suo et attacus atque ophiomachus ac locusta, singula iuxta genus suum.
LEV|11|23|Quidquid autem ex volucribus reptantibus quattuor tantum habet pedes, execrabile erit vobis.
LEV|11|24|Et quicumque morticina eorum tetigerit, polluetur et erit immundus usque ad vesperum.
LEV|11|25|Et si necesse fuerit, ut portet quippiam horum mortuum, lavabit vestimenta sua et immundus erit usque ad solis occasum.
LEV|11|26|Omne animal, quod habet quidem ungulam, sed non dividit eam nec ruminat, immundum erit vobis; et, qui tetigerit illud, contaminabitur.
LEV|11|27|Quod ambulat super plantas pedum ex cunctis animantibus, quae incedunt quadrupedia, immundum erit; qui tetigerit morticina eorum, polluetur usque ad vesperum.
LEV|11|28|Et, qui portaverit huiuscemodi cadavera, lavabit vestimenta sua et immundus erit usque ad vesperum; quia omnia haec immunda sunt vobis.
LEV|11|29|Haec quoque inter polluta reputabuntur de his, quae reptant in terra: mustela et mus et lacerta iuxta genus suum,
LEV|11|30|mygale et testudo et stellio et talpa et chamaeleon:
LEV|11|31|omnia haec immunda sunt.Qui tetigerit morticina eorum, immundus erit usque ad vesperum;
LEV|11|32|et super quod ceciderit quidquam de morticinis eorum, polluetur tam vas ligneum et vestimentum quam pelles et cilicia, et in quocumque fit opus; tinguentur aqua et polluta erunt usque ad vesperum et postea munda.
LEV|11|33|Vas autem fictile, in quo horum quidquam intro ceciderit, polluetur et frangendum est.
LEV|11|34|Omnis cibus, quem comedetis, si fusa fuerit exinde super eum aqua, immundus erit; et omne liquens, quod bibitur de tali vase, immundum erit.
LEV|11|35|Et quidquid de morticinis istiusmodi ceciderit super illud, immundum erit; sive clibani sive chytropodes destruentur: immundi sunt et immundi erunt vobis.
LEV|11|36|Fontes tamen et cisternae et omnis aquarum congregatio munda erit. Qui vero morticinum eorum tetigerit, polluetur.
LEV|11|37|Si ceciderint super sementem, non polluent eam;
LEV|11|38|sin autem quispiam aqua sementem perfuderit, et postea morticinis tacta fuerit, immunda erit vobis.
LEV|11|39|Si mortuum fuerit animal, quod licet vobis comedere, qui cadaver eius tetigerit, immundus erit usque ad vesperum;
LEV|11|40|et, qui comederit ex eo quippiam sive portaverit cadaver eius, lavabit vestimenta sua et immundus erit usque ad vesperum.
LEV|11|41|Omne, quod reptat super terram, abominabile erit nec assumetur in cibum.
LEV|11|42|Quidquid super pectus et quidquid quadrupes graditur, vel multos habet pedes sive per humum trahitur, non comedetis, quia abominabile est.
LEV|11|43|Nolite contaminare animas vestras nec tangatis quidquam eorum, ne immundi sitis.
LEV|11|44|Ego enim sum Dominus Deus vester; sanctificamini et sancti estote, quoniam et ego sanctus sum. Ne polluatis animas vestras in omni reptili, quod movetur super terram.
LEV|11|45|Ego enim sum Dominus, qui eduxi vos de terra Aegypti, ut essem vobis in Deum: sancti eritis, quia et ego sanctus sum.
LEV|11|46|Ista est lex animantium et volucrum et omnis animae viventis, quae movetur in aqua et reptat in terra,
LEV|11|47|ut differentias noveritis mundi et immundi, et sciatis quid comedere et quid respuere debeatis ".
LEV|12|1|Locutus est Dominus ad Moysen dicens:
LEV|12|2|" Loquere fi liis Israel et dices ad eos: Mulier, si, suscepto semine, pepererit masculum, immunda erit septem diebus iuxta dies separationis menstruae,
LEV|12|3|et die octavo circumcidetur infantulus;
LEV|12|4|ipsa vero triginta tribus diebus manebit in sanguine purificationis suae; omne sanctum non tanget nec ingredietur sanctuarium, donec impleantur dies purificationis eius.
LEV|12|5|Sin autem feminam pepererit, immunda erit duabus hebdomadibus iuxta ritum fluxus menstrui, et sexaginta ac sex diebus manebit in sanguine purificationis suae.
LEV|12|6|Cumque expleti fuerint dies purificationis suae pro filio sive pro filia, deferet agnum anniculum in holocaustum et pullum columbae sive turturem pro peccato ad ostium tabernaculi conventus et tradet sacerdoti.
LEV|12|7|Qui offeret illa coram Domino et expiabit eam; et sic mundabitur a profluvio sanguinis sui: ista est lex parientis masculum aut feminam.
LEV|12|8|Quod si non invenerit manus eius, nec potuerit offerre agnum, sumet duos turtures vel duos pullos columbae, unum in holocaustum et alterum pro peccato; expiabitque eam sacerdos, et sic mundabitur ".
LEV|13|1|Locutus est Dominus ad Moysen et Aaron dicens:
LEV|13|2|" Homo, in cuius carne et cute ortus fuerit tumor sive pustula aut quasi lucens quippiam, id est plaga leprae, adducetur ad Aaron sacerdotem vel ad unum quemlibet filiorum eius sacerdotum.
LEV|13|3|Qui cum viderit plagam in cute et pilos in album mutatos colorem ipsamque speciem plagae humiliorem cute et carne reliqua: plaga leprae est; quod cum viderit sacerdos, eum immundum esse decernet.
LEV|13|4|Sin autem lucens candor fuerit in cute nec humilior carne reliqua, et pili coloris pristini, recludet eum sacerdos septem diebus.
LEV|13|5|Et considerabit eum die septimo: et, siquidem plaga ultra non creverit nec transierit in cute priores terminos, rursum recludet eum septem diebus aliis.
LEV|13|6|Et die septimo contemplabitur eum iterum: si obscurior fuerit plaga et non creverit in cute, eum mundum esse decernet, quia scabies est. Lavabitque homo vestimenta sua et mundus erit.
LEV|13|7|Quod si, postquam a sacerdote visus est et redditus munditiae, iterum scabies creverit, adducetur ad eum;
LEV|13|8|et, si viderit ita esse, immunditiae condemnabitur: est lepra.
LEV|13|9|Plaga leprae si fuerit in homine, adducetur ad sacerdotem,
LEV|13|10|et videbit eum. Cumque tumor albus in cute fuerit et capillorum mutaverit aspectum in album, caro quoque viva creverit in tumore,
LEV|13|11|lepra vetustissima iudicabitur atque inolita cuti. Contaminabit itaque eum sacerdos et non recludet, quia perspicue immunditia est.
LEV|13|12|Sin autem effloruerit discurrens lepra in cute et operuerit omnem cutem a capite usque ad pedes, quidquid sub aspectu oculorum cadit,
LEV|13|13|considerabit eum sacerdos et teneri lepra mundissima iudicabit, eo quod omnis in candorem versa sit, et idcirco homo mundus erit.
LEV|13|14|Quando vero caro vivens in eo apparuerit, immundus erit.
LEV|13|15|Quod cum sacerdos viderit, inter immundos reputabit; caro enim viva immunda est: lepra est.
LEV|13|16|Quod si rursum versa fuerit in alborem, veniet ad sacerdotem,
LEV|13|17|qui cum hoc consideraverit, eum mundum esse decernet.
LEV|13|18|Caro et cutis, in qua ulcus natum est et sanatum,
LEV|13|19|et in loco ulceris tumor apparuerit albus sive macula subrufa, ostendet se homo sacerdoti.
LEV|13|20|Qui cum viderit locum maculae humiliorem carne reliqua et pilos versos in candorem, contaminabit eum: plaga enim leprae orta est in ulcere.
LEV|13|21|Quod si pilus coloris est pristini et cicatrix subobscura et vicina carne non est humilior, recludet eum septem diebus.
LEV|13|22|Et, siquidem creverit, adiudicabit eum leprae;
LEV|13|23|sin autem steterit in loco suo macula nec creverit, ulceris est cicatrix, et sacerdos eum mundum esse decernet.
LEV|13|24|Vel si alicuius cutem ignis exusserit, et locus exustionis subrufam sive albam habuerit maculam,
LEV|13|25|considerabit eam sacerdos; et ecce pilus versus est in alborem, et locus eius reliqua cute humilior, contaminabit eum, quia plaga leprae in cicatrice orta est.
LEV|13|26|Quod si pilorum color non fuerit immutatus, nec humilior macula carne reliqua, et ipsa leprae species fuerit subobscura, recludet eum septem diebus.
LEV|13|27|Et die septimo contemplabitur eum; si creverit in cute macula, contaminabit eum: plaga est leprae;
LEV|13|28|sin autem in loco suo macula steterit non satis clara, tumor combustionis est, et idcirco mundabit eum, quia cicatrix est combusturae.
LEV|13|29|Vir sive mulier, in cuius capite vel barba germinarit plaga, videbit eam sacerdos.
LEV|13|30|Et, siquidem humilior fuerit locus carne reliqua, et capillus flavus solitoque subtilior, contaminabit eos, quia scabies est, lepra capitis vel barbae.
LEV|13|31|Sin autem viderit plagam scabiei aequalem vicinae carni nec capillum nigrum in ea, recludet eos septem diebus.
LEV|13|32|Et die septimo intuebitur plagam: si non creverit scabies, nec capillus flavus fuerit in ea, et locus plagae carni reliquae aequalis,
LEV|13|33|radetur homo absque loco maculae, et includet eum sacerdos septem diebus aliis.
LEV|13|34|Si die septimo visa fuerit stetisse plaga in loco suo nec humilior carne reliqua, mundabit eum sacerdos; lotisque vestibus mundus erit.
LEV|13|35|Sin autem post emundationem rursus creverit scabies in cute,
LEV|13|36|non quaeret amplius utrum capillus in flavum colorem sit commutatus, quia aperte immundus est.
LEV|13|37|Porro si steterit macula, et capilli nigri fuerint, noverit hominem esse sanatum et confidenter eum pronuntiet mundum.
LEV|13|38|Vir et mulier, in cuius cute maculae, maculae albae apparuerint,
LEV|13|39|intuebitur eos sacerdos. Si deprehenderit subobscurum alborem lucere in cute, sciat impetiginem ortam esse in cute; mundus est.
LEV|13|40|Vir, de cuius capite capilli fluunt, calvus ac mundus est;
LEV|13|41|et, si a fronte ceciderint pili, recalvaster et mundus est.
LEV|13|42|Sin autem in calvitio sive in recalvatione plaga alba vel subrufa fuerit exorta, lepra est capitis.
LEV|13|43|Sacerdos eum videbit, et ecce tumor plagae subrufus secundum aspectum leprae cutis carnis.
LEV|13|44|Vir maculatus est lepra, et sacerdos omnino decernet eum esse immundum; plaga est in capite eius.
LEV|13|45|Leprosus hac plaga percussus habebit vestimenta dissuta, comam capitis excussam, barbam contectam; clamabit: "Immundus! Immundus!".
LEV|13|46|Omni tempore, quo leprosus est immundus, immundus est et solus habitabit extra castra.
LEV|13|47|Si in veste lanea sive linea lepra fuerit,
LEV|13|48|in stamine sive subtemine lineo vel laneo aut in pelle vel quolibet ex pelle confecto,
LEV|13|49|si macula pallida aut rufa fuerit, lepra reputabitur ostendeturque sacerdoti.
LEV|13|50|Qui considerabit macula infectum et recludet septem diebus;
LEV|13|51|et die septimo rursus aspiciens, si crevisse deprehenderit, lepra maligna est; pollutum iudicabit vestimentum et omne, in quo fuerit inventa,
LEV|13|52|et idcirco comburetur flammis.
LEV|13|53|Quod si eam viderit non crevisse,
LEV|13|54|praecipiet, et lavabunt id, in quo plaga est; recludetque illud septem diebus aliis.
LEV|13|55|Et cum viderit post lavationem faciem quidem pristinam non mutatam, nec tamen crevisse plagam, immunda est res, et igne combures eam, eo quod infusa sit plaga in superficie rei vel in parte aversa.
LEV|13|56|Sin autem obscurior fuerit locus plagae, postquam res est lota, sacerdos abrumpet eum et a solido dividet.
LEV|13|57|Quod si macula ultra apparuerit in his rebus, quae prius immaculata erant, lepra volatilis et vaga, igne combures illas.
LEV|13|58|Quas vero laveris et a quibus cessaverit plaga, illas lavabis secundo, et mundae erunt.
LEV|13|59|Ista est lex leprae vestimenti lanei et linei, staminis atque subteminis, omnisque supellectilis pelliceae, quomodo mundari debeat vel contaminari ".
LEV|14|1|Locutusque est Dominus ad Moysen dicens:
LEV|14|2|" Hic est ri tus leprosi, quando mundandus est: adducetur ad sacerdotem,
LEV|14|3|qui egressus e castris, cum invenerit lepram esse sanatam,
LEV|14|4|praecipiet, ut sumant pro eo, qui purificatur, duas aves vivas, mundas et lignum cedrinum vermiculumque et hyssopum.
LEV|14|5|Et unam ex avibus immolari iubebit in vase fictili super aquas viventes.
LEV|14|6|Aliam autem vivam cum ligno cedrino et cocco et hyssopo tinguet in sanguine avis super aquas viventes immolatae,
LEV|14|7|quo asperget illum, qui a lepra mundandus est, septies, ut iure purgetur; et dimittet avem vivam, ut in agrum avolet.
LEV|14|8|Cumque laverit homo vestimenta sua, radet omnes pilos corporis, et lavabitur aqua; purificatusque ingredietur castra, ita dumtaxat ut maneat extra tabernaculum suum septem diebus.
LEV|14|9|Et die septimo radet capillos capitis barbamque et supercilia ac totius corporis pilos et lavabit vestimenta carnemque suam aqua, et mundus erit.
LEV|14|10|Die octavo assumet duos agnos immaculatos et ovem anniculam absque macula et tres decimas ephi similae in sacrificium, quae conspersa sit oleo, et log olei.
LEV|14|11|Cumque sacerdos purificans hominem statuerit eum et haec omnia coram Domino in ostio tabernaculi conventus,
LEV|14|12|tollet agnum unum et offeret eum in sacrificium pro delicto, oleique log et, elevatis ante Dominum omnibus,
LEV|14|13|immolabit agnum, ubi immolari solet hostia pro peccato et holocaustum, id est in loco sancto. Sicut enim pro peccato ita et pro delicto ad sacerdotem pertinet sacrificium: sanctum sanctorum est.
LEV|14|14|Assumensque sacerdos de sanguine hostiae pro delicto ponet super extremum auriculae dextrae eius, qui mundatur, et super pollices manus dextrae et pedis;
LEV|14|15|et de olei log mittet in manum suam sinistram
LEV|14|16|tinguetque digitum dextrum in eo et asperget septies coram Domino.
LEV|14|17|Quod autem reliquum est olei in laeva manu, fundet super extremum auriculae dextrae eius, qui mundatur, et super pollices manus ac pedis dextri et super sanguinem sacrificii pro delicto
LEV|14|18|et super caput eius, qui mundatur; expiabitque eum coram Domino
LEV|14|19|et faciet sacrificium pro peccato. Tunc immolabit holocaustum
LEV|14|20|et ponet illud in altari cum sacrificio similae, et homo rite mundabitur.
LEV|14|21|Quod si pauper est, et non potest manus eius invenire, quae dicta sunt, assumet agnum pro delicto ad elationem, ut expiet eum sacerdos, decimamque partem similae conspersae oleo in sacrificium et olei log
LEV|14|22|duosque turtures sive duos pullos columbae, quos manus eius invenire poterit, unum pro peccato et alterum in holocaustum.
LEV|14|23|Offeretque ea die octavo purificationis suae sacerdoti ad ostium tabernaculi conventus coram Domino.
LEV|14|24|Qui suscipiens agnum pro delicto et log olei levabit simul coram Domino;
LEV|14|25|immolatoque agno pro delicto, de sanguine eius ponet super extremum auriculae dextrae illius, qui mundatur, et super pollices manus eius ac pedis dextri;
LEV|14|26|olei vero partem mittet in manum suam sinistram.
LEV|14|27|In quo tinguens digitum dextrae manus asperget septies coram Domino;
LEV|14|28|tangetque extremum auriculae dextrae illius, qui mundatur, et pollices manus ac pedis dextri super locum sanguinis, qui effusus est pro delicto.
LEV|14|29|Reliquam autem partem olei, quae est in sinistra manu, mittet super caput hominis, qui purificatur, in expiationem eius coram Domino;
LEV|14|30|et turtures sive pullos columbae, quos manus illius invenerit, offeret,
LEV|14|31|unum pro delicto et alterum in holocaustum cum sacrificio similae, et sic expiabit eum sacerdos coram Domino.
LEV|14|32|Hoc est sacrificium leprosi, qui habere non potest omnia in emundationem sui ".
LEV|14|33|Locutus est Dominus ad Moysen et Aaron dicens:
LEV|14|34|" Cum ingressi fueritis terram Chanaan, quam ego dabo vobis in possessionem, si fuerit plaga leprae in aedibus terrae possessionis vestrae,
LEV|14|35|ibit, cuius est domus, nuntians sacerdoti et dicet: "Quasi plaga videtur mihi esse in domo mea".
LEV|14|36|At ille praecipiet, ut efferant universa de domo, priusquam ingrediatur eam, et videat plagam, ne immunda fiant omnia, quae in domo sunt. Intrabitque postea, ut consideret domum;
LEV|14|37|et, cum viderit in parietibus illius quasi valliculas pallore sive rubore deformes et humiliores superficie reliqua,
LEV|14|38|egredietur ostium domus et statim claudet eam septem diebus.
LEV|14|39|Reversusque die septimo considerabit eam; si invenerit crevisse plagam,
LEV|14|40|iubebit erui lapides, in quibus plaga est, et proici eos extra civitatem in loco immundo;
LEV|14|41|domum autem ipsam radi intrinsecus per circuitum et spargi pulverem rasurae extra urbem in locum immundum
LEV|14|42|lapidesque alios reponi pro his, qui ablati fuerint, et luto alio liniri domum.
LEV|14|43|Sin autem plaga rursum effloruerit in domo, postquam eruti sunt lapides et pulvis erasus et alia terra lita,
LEV|14|44|et ingressus sacerdos viderit crevisse plagam in domo: lepra est maligna et domus immunda.
LEV|14|45|Quam statim destruent et lapides eius ac ligna atque universum pulverem domus proicient extra oppidum in loco immundo.
LEV|14|46|Qui intraverit domum, quando clausa est, immundus erit usque ad vesperum;
LEV|14|47|et, qui dormierit in ea vel comederit quippiam, lavabit vestimenta sua.
LEV|14|48|Quod si introiens sacerdos viderit plagam non crevisse in domo, postquam denuo lita est, mundam eam esse decernet, reddita sanitate.
LEV|14|49|Et in purificationem eius sumet duas aves lignumque cedrinum et vermiculum atque hyssopum
LEV|14|50|et, immolata una avi in vase fictili super aquas vivas,
LEV|14|51|tollet lignum cedrinum et hyssopum et coccum et avem vivam et intinguet omnia in sanguine avis immolatae atque in aquis viventibus et asperget domum septies;
LEV|14|52|purificabitque eam tam in sanguine avis quam in aquis viventibus et in avi viva lignoque cedrino et hyssopo atque vermiculo;
LEV|14|53|cumque dimiserit avem avolare extra urbem in agrum libere, expiabit domum, et erit munda.
LEV|14|54|Ista est lex omnis leprae et scabiei,
LEV|14|55|leprae vestium et domorum,
LEV|14|56|tumoris et pustulae et lucentis maculae,
LEV|14|57|ut possit sciri quo tempore immundum quid vel mundum sit ".
LEV|15|1|Locutus est Dominus ad Moysen et Aaron dicens:
LEV|15|2|" Loquimini filiis Israel et dicite eis: Vir, si patitur fluxum seminis, immundus erit.
LEV|15|3|Et tunc iudicabitur huic vitio subiacere: sive emiserit caro eius fluxum suum vel occluserit se a fluxu.
LEV|15|4|Omne stratum, in quo iacuerit, immundum erit, et ubicumque sederit.
LEV|15|5|Si quis hominum tetigerit lectum eius, lavabit vestimenta sua, et ipse lotus aqua immundus erit usque ad vesperum.
LEV|15|6|Si sederit, ubi ille sederat, et ipse lavabit vestimenta sua et lotus aqua immundus erit usque ad vesperum.
LEV|15|7|Qui tetigerit carnem eius, lavabit vestimenta sua et ipse lotus aqua immundus erit usque ad vesperum.
LEV|15|8|Si salivam huiuscemodi homo iecerit super eum, qui mundus est, hic lavabit vestem suam et lotus aqua immundus erit usque ad vesperum.
LEV|15|9|Sagma, super quo sederit, immundum erit;
LEV|15|10|et quicumque tetigerit omne, quod sub eo fuerit, qui fluxum seminis patitur, pollutus erit usque ad vesperum. Qui portaverit horum aliquid, lavabit vestem suam et ipse lotus aqua immundus erit usque ad vesperum.
LEV|15|11|Omnis, quem tetigerit, qui fluxum patitur, non lotis ante manibus, lavabit vestimenta sua et lotus aqua immundus erit usque ad vesperum.
LEV|15|12|Vas fictile, quod tetigerit, confringetur; vas autem ligneum lavabitur aqua.
LEV|15|13|Si sanatus fuerit, qui huiuscemodi sustinet passionem, numerabit septem dies ad emundationem sui et, lotis vestibus ac toto corpore in aquis viventibus, erit mundus.
LEV|15|14|Die autem octavo sumet duos turtures aut duos pullos columbae et veniet in conspectu Domini ad ostium tabernaculi conventus dabitque eos sacerdoti.
LEV|15|15|Qui faciet unum in sacrificium pro peccato et alterum in holocaustum; expiabitque eum coram Domino et emundabitur a fluxu seminis sui.
LEV|15|16|Vir, de quo egreditur semen, lavabit aqua omne corpus suum et immundus erit usque ad vesperum.
LEV|15|17|Vestem et pellem, super quam fuerit semen effusum, lavabitur aqua et immunda erit usque ad vesperum.
LEV|15|18|Si cum muliere coierit vir, lavabunt se aqua et immundi erunt usque ad vesperum.
LEV|15|19|Mulier, quae redeunte mense patitur fluxum sanguinis, septem diebus separabitur. Omnis, qui tetigerit eam, immundus erit usque ad vesperum;
LEV|15|20|et in quo iacuerit vel sederit diebus separationis suae, polluetur.
LEV|15|21|Qui tetigerit lectum eius, lavabit vestimenta sua et ipse lotus aqua immundus erit usque ad vesperum.
LEV|15|22|Omne vas, super quo illa sederit, quisquis attigerit, lavabit vestimenta sua et ipse lotus aqua pollutus erit usque ad vesperum.
LEV|15|23|Et quicumque tetigerit omne, quod fuerit super lectum vel supellectilem, in qua illa sederit, immundus erit usque ad vesperum.
LEV|15|24|Si coierit cum ea vir tempore sanguinis menstrualis, immundus erit septem diebus, et omne stratum, in quo dormierit, polluetur.
LEV|15|25|Mulier, quae patitur multis diebus fluxum sanguinis non in tempore menstruali vel quae post menstruum sanguinem fluere non cessat, quamdiu huic subiacet passioni, immunda erit quasi sit in tempore menstruo.
LEV|15|26|Omne stratum, in quo dormierit, et vas, in quo sederit, pollutum erit.
LEV|15|27|Quicumque tetigerit ea, polluetur; lavabit vestimenta sua et ipse lotus aqua immundus erit usque ad vesperum.
LEV|15|28|Si steterit sanguis et fluere cessarit, numerabit septem dies et deinde munda erit.
LEV|15|29|Et octavo die assumet pro se duos turtures vel duos pullos columbae afferetque sacerdoti ad ostium tabernaculi conventus.
LEV|15|30|Qui unum faciet in sacrificium pro peccato et alterum in holocaustum; expiabitque eam coram Domino a fluxu immunditiae eius.
LEV|15|31|Docebitis ergo filios Israel, ut caveant immunditiam, ne moriantur in sordibus suis, cum polluerint habitaculum meum, quod est inter eos.
LEV|15|32|Ista est lex eius, qui patitur fluxum seminis et de quo egreditur semen et polluitur,
LEV|15|33|et quae menstruis temporibus separatur vel quae iugi fluit sanguine, et hominis, qui dormierit cum immunda ".
LEV|16|1|Locutusque est Dominus ad Moysen post mortem duum filiorum Aaron, quando appropinquantes in conspectum Domini interfecti sunt,
LEV|16|2|et praecepit ei dicens: " Loquere ad Aaron fratrem tuum, ne omni tempore ingrediatur sanctuarium, quod est intra velum coram propitiatorio, quo tegitur arca, ut non moriatur, quia in nube apparebo super propitiatorium;
LEV|16|3|sed hoc modo ingrediatur: vitulum offeret pro peccato et arietem in holocaustum;
LEV|16|4|subucula linea sancta vestietur, feminalibus lineis verecunda celabit, accingetur zona linea, cidarim lineam imponet capiti. Haec enim vestimenta sunt sancta, quibus cunctis, cum lotus fuerit, induetur.
LEV|16|5|Suscipietque a coetu filiorum Israel duos hircos in sacrificium pro peccato et unum arietem in holocaustum.
LEV|16|6|Cumque obtulerit vitulum in sacrificium suum pro peccato et expiaverit se et domum suam,
LEV|16|7|duos hircos stare faciet coram Domino in ostio tabernaculi conventus,
LEV|16|8|mittens super utrumque sortem, unam Domino et alteram Azazel.
LEV|16|9|Cuius sors exierit Domino, offeret illum pro peccato;
LEV|16|10|cuius autem in Azazel, statuet eum vivum coram Domino in expiationem, ut emittat illum ad Azazel in solitudinem.
LEV|16|11|Afferet ergo Aaron vitulum pro peccato et expians se et domum suam immolabit eum;
LEV|16|12|assumptoque turibulo, quod de prunis altaris coram Domino impleverit, et hauriens manu compositum thymiama in incensum ultra velum intrabit in sancta,
LEV|16|13|ut, positis super ignem aromatibus coram Domino, nebula eorum et vapor operiat propitiatorium, quod est super testimonium, et non moriatur.
LEV|16|14|Tollet quoque de sanguine vituli et asperget digito septies contra frontem propitiatorii.
LEV|16|15|Cumque mactaverit hircum pro peccato populi, inferet sanguinem eius intra velum, sicut praeceptum est de sanguine vituli, ut aspergat e regione propitiatorii
LEV|16|16|et expiet sanctuarium ab immunditiis filiorum Israel et a praevaricationibus eorum cunctisque peccatis. Iuxta hunc ritum faciet tabernaculo conventus, quod fixum est inter eos in medio sordium habitationis eorum.
LEV|16|17|Nullus hominum sit in tabernaculo conventus, quando pontifex ingreditur sanctuarium, ut expiet se et domum suam et universam congregationem Israel, donec egrediatur.
LEV|16|18|Cum autem exierit ad altare, quod coram Domino est, expiabit illud et sumptum sanguinem vituli atque hirci fundet super cornua eius per gyrum;
LEV|16|19|aspergensque de sanguine digito septies mundabit sanctificabitque illud ab immunditiis filiorum Israel.
LEV|16|20|Et postquam compleverit expiationem sanctuarii et tabernaculi conventus et altaris, tunc afferat hircum viventem;
LEV|16|21|et, posita utraque manu super caput eius, confiteatur Aaron super eum omnes iniquitates filiorum Israel et universa delicta atque peccata eorum; quae ponens super caput eius emittet illum per hominem paratum in desertum.
LEV|16|22|Cumque portaverit hircus super se omnes iniquitates eorum in terram solitariam et dimissus fuerit in desertum,
LEV|16|23|ingredietur Aaron in tabernaculum conventus; et, depositis vestibus lineis, quibus prius indutus erat, cum intraret sanctuarium, relictisque ibi,
LEV|16|24|lavabit carnem suam aqua in loco sancto indueturque vestimentis suis. Et postquam egressus obtulerit holocaustum suum ac plebis, expiabit se et populum;
LEV|16|25|et adipem sacrificii pro peccato adolebit super altare.
LEV|16|26|Ille vero, qui dimiserit caprum emissarium ad Azazel, lavabit vestimenta sua et corpus aqua et postea ingredietur in castra.
LEV|16|27|Vitulum autem et hircum, qui pro peccato fuerant immolati, et quorum sanguis illatus est, ut in sanctuario expiatio compleretur, asportabunt foras castra et comburent igni tam pelles quam carnes eorum et fimum;
LEV|16|28|et quicumque combusserit ea, lavabit vestimenta sua et carnem aqua et postea ingredietur in castra.
LEV|16|29|Eritque hoc vobis legitimum sempiternum: mense septimo, decima die mensis affligetis animas vestras nullumque facietis opus sive indigena sive advena, qui peregrinatur inter vos.
LEV|16|30|In hac die expiatio erit vestri atque mundatio; ab omnibus peccatis vestris coram Domino mundabimini.
LEV|16|31|Sabbatum requietionis est vobis, et affligetis animas vestras religione perpetua.
LEV|16|32|Expiabit autem sacerdos, qui unctus fuerit, et cuius initiatae manus, ut sacerdotio fungatur pro patre suo; indueturque vestimentis lineis, vestibus sanctis,
LEV|16|33|et expiabit sanctuarium sanctissimum et tabernaculum conventus atque altare, sacerdotes quoque et universum populum congregationis.
LEV|16|34|Eritque hoc vobis legitimum sempiternum, ut expietis filios Israel a cunctis peccatis eorum semel in anno ".Fecit igitur, sicut praeceperat Dominus Moysi.
LEV|17|1|Et locutus est Dominus ad Moysen dicens:
LEV|17|2|" Loquere Aaron et filiis eius et cunctis filiis Israel et dices ad eos: Iste est sermo, quem mandavit Dominus dicens:
LEV|17|3|Homo quilibet de domo Israel, si occiderit bovem aut ovem sive capram in castris vel extra castra
LEV|17|4|et non attulerit ad ostium tabernaculi conventus in oblationem Domino coram habitaculo Domini, sanguinis reus erit; sanguinem fudit et peribit de medio populi sui.
LEV|17|5|Ideo offerre debent sacerdoti filii Israel hostias suas, quas occidunt in agro, ut afferant Domino ante ostium tabernaculi conventus et immolent eas hostias pacificas Domino.
LEV|17|6|Fundetque sacerdos sanguinem super altare Domini ad ostium tabernaculi conventus et adolebit adipem in odorem suavitatis Domino;
LEV|17|7|et nequaquam ultra immolabunt hostias suas daemonibus, cum quibus fornicati sunt: legitimum sempiternum erit hoc illis et posteris eorum ".
LEV|17|8|Et ad ipsos dices: " Homo de domo Israel et de advenis, qui peregrinantur apud vos, qui obtulerit holocaustum sive sacrificium
LEV|17|9|et ad ostium tabernaculi conventus non adduxerit victimam, ut offeratur Domino, interibit de populo suo.
LEV|17|10|Homo quilibet de domo Israel et de advenis, qui peregrinantur inter eos, si comederit sanguinem, confirmabo faciem meam contra talem animam et disperdam eam de populo suo.
LEV|17|11|Quia anima carnis in sanguine est, et ego dedi illum vobis, ut super altare in eo expietis pro animabus vestris, quia sanguis ipse per animam expiat.
LEV|17|12|Idcirco dixi filiis Israel: Omnis anima ex vobis non comedet sanguinem, nec ex advenis, qui peregrinantur inter vos.
LEV|17|13|Homo quicumque de filiis Israel et de advenis, qui peregrinantur apud vos, si venatione ceperit feram vel avem, quibus vesci licitum est, fundat sanguinem eius et operiat illum terra.
LEV|17|14|Anima enim omnis carnis, sanguis est anima eius, unde dixi filiis Israel: Sanguinem universae carnis non comedetis, quia anima omnis carnis sanguis eius est; et, quicumque comederit illum, interibit.
LEV|17|15|Anima, quae comederit morticinum vel captum a bestia, tam de indigenis quam de advenis, lavabit vestes suas et semetipsum aqua, et contaminatus erit usque ad vesperum; et hoc ordine mundus fiet.
LEV|17|16|Quod si non laverit vestimenta sua nec corpus, portabit iniquitatem suam ".
LEV|18|1|Locutus est Dominus ad Moysen dicens:
LEV|18|2|" Loquere fi liis Israel et dices ad eos: Ego Dominus Deus vester.
LEV|18|3|Iuxta consuetudinem terrae Aegypti, in qua habitastis, non facietis; et iuxta morem regionis Chanaan, ad quam ego introducturus sum vos, non agetis nec in legitimis eorum ambulabitis.
LEV|18|4|Facietis iudicia mea et praecepta mea servabitis et ambulabitis in eis. Ego Dominus Deus vester.
LEV|18|5|Custodite leges meas atque iudicia; quae faciens homo vivet in eis. Ego Dominus.
LEV|18|6|Omnis homo ad consanguineum suum non accedet, ut revelet turpitudinem eius. Ego Dominus.
LEV|18|7|Turpitudinem patris et turpitudinem matris tuae non discooperies: mater tua est, non revelabis turpitudinem eius.
LEV|18|8|Turpitudinem uxoris patris tui non discooperies, turpitudo enim patris tui est.
LEV|18|9|Turpitudinem sororis tuae ex patre sive ex matre, quae domi vel foris genita est, non revelabis.
LEV|18|10|Turpitudinem filiae filii tui vel neptis ex filia non revelabis, quia turpitudo tua est.
LEV|18|11|Turpitudinem filiae uxoris patris tui, quam peperit patri tuo et est soror tua, non revelabis.
LEV|18|12|Turpitudinem sororis patris tui non discooperies, quia caro est patris tui.
LEV|18|13|Turpitudinem sororis matris tuae non revelabis, eo quod caro sit matris tuae.
LEV|18|14|Turpitudinem patrui tui non revelabis nec accedes ad uxorem eius, quae tibi affinitate coniungitur.
LEV|18|15|Turpitudinem nurus tuae non revelabis, quia uxor filii tui est, nec discooperies ignominiam eius.
LEV|18|16|Turpitudinem uxoris fratris tui non revelabis, quia turpitudo fratris tui est.
LEV|18|17|Turpitudinem mulieris et filiae eius non revelabis. Filiam filii eius et filiam filiae illius non sumes, ut reveles ignominiam eius, quia caro illius sunt: nefas est.
LEV|18|18|Sororem uxoris tuae aemulam illius non accipies nec revelabis turpitudinem eius, adhuc illa vivente.
LEV|18|19|Ad mulierem, quae patitur menstrua, non accedes nec revelabis foeditatem eius.
LEV|18|20|Cum uxore proximi tui non coibis nec seminis commixtione maculaberis.
LEV|18|21|De semine tuo non dabis, ut consecretur idolo Moloch, nec pollues nomen Dei tui. Ego Dominus.
LEV|18|22|Cum masculo non commisceberis coitu femineo: abominatio est.
LEV|18|23|Cum omni pecore non coibis nec maculaberis cum eo. Mulier non succumbet iumento nec miscebitur ei, quia scelus est.
LEV|18|24|Ne polluamini in omnibus his, quibus contaminatae sunt universae gentes, quas ego eiciam ante conspectum vestrum
LEV|18|25|et quibus polluta est terra, cuius ego scelera visitavi, et evomuit habitatores suos.
LEV|18|26|Vos autem custodite legitima mea atque iudicia et non faciatis ex omnibus abominationibus istis tam indigena quam colonus, qui peregrinatur apud vos.
LEV|18|27|Omnes enim execrationes istas fecerunt accolae terrae, qui fuerunt ante vos, et polluerunt eam.
LEV|18|28|Cavete ergo, ne et vos similiter evomat, cum pollueritis eam, sicut evomuit gentem, quae fuit ante vos.
LEV|18|29|Omnis enim anima, quae fecerit de abominationibus his quippiam, peribit de medio populi sui.
LEV|18|30|Custodite mandata mea. Nolite facere legitima abominabilia, quae fecerunt hi, qui fuerunt ante vos, et ne polluamini in eis. Ego Dominus Deus vester ".
LEV|19|1|Locutus est Dominus ad Moysen dicens:
LEV|19|2|" Loquere ad omnem coetum filiorum Israel et dices ad eos: Sancti estote, quia sanctus sum ego, Dominus Deus vester.
LEV|19|3|Unusquisque matrem et patrem suum timeat. Sabbata mea custodite. Ego Dominus Deus vester.
LEV|19|4|Nolite converti ad idola nec deos conflatiles faciatis vobis. Ego Dominus Deus vester.
LEV|19|5|Si immolaveritis hostiam pacificorum Domino, immolabitis eam ita ut sit vobis placabilis.
LEV|19|6|Eo die, quo fuerit immolata, comedetur et die altero; quidquid autem residuum fuerit in diem tertium, igne comburetur.
LEV|19|7|Si quid post biduum comestum fuerit, profanum erit neque acceptabile.
LEV|19|8|Qui manducaverit illud, portabit iniquitatem suam, quia sanctum Domini polluit, et peribit anima illa de populo suo.
LEV|19|9|Cum messueris segetes terrae tuae, non tondebis usque ad marginem agri tui nec remanentes spicas colliges.
LEV|19|10|Neque in vinea tua racemos et grana decidentia congregabis, sed pauperibus et peregrinis carpenda dimittes. Ego Dominus Deus vester.
LEV|19|11|Non facietis furtum. Non mentiemini, nec decipiet unusquisque proximum suum.
LEV|19|12|Non periurabis in nomine meo nec pollues nomen Dei tui. Ego Dominus.
LEV|19|13|Non facies calumniam proximo tuo nec spoliabis eum. Non morabitur merces mercennarii apud te usque mane.
LEV|19|14|Non maledices surdo nec coram caeco pones offendiculum; sed timebis Deum tuum. Ego Dominus.
LEV|19|15|Non facietis, quod iniquum est in iudicio. Non consideres personam pauperis nec honores vultum potentis. Iuste iudica proximo tuo.
LEV|19|16|Non eris criminator et susurro in populo tuo. Non stabis contra sanguinem proximi tui. Ego Dominus.
LEV|19|17|Ne oderis fratrem tuum in corde tuo; argue eum, ne habeas super illo peccatum.
LEV|19|18|Non quaeres ultionem nec irasceris civibus tuis. Diliges proximum tuum sicut teipsum. Ego Dominus.
LEV|19|19|Leges meas custodite.Iumenta tua non facies coire cum alterius generis animantibus. Agrum tuum non seres diverso semine. Veste, quae ex duobus texta est, non indueris.
LEV|19|20|Homo, si dormierit cum muliere coitu seminis, quae sit ancilla destinata viro et tamen pretio non redempta nec libertate donata, vapulabunt ambo et non morientur, quia non fuit libera.
LEV|19|21|Et in sacrificium suum pro delicto offeret Domino ad ostium tabernaculi conventus arietem;
LEV|19|22|expiabitque eum sacerdos ariete a peccato eius coram Domino, et dimittetur ei peccatum, quod peccavit.
LEV|19|23|Quando ingressi fueritis terram et plantaveritis omnimoda ligna pomifera, non auferetis praeputia eorum, id est poma, quae germinant; tribus annis erunt vobis immunda ut praeputia, nec edetis ex eis.
LEV|19|24|Quarto anno omnis fructus eorum sanctificabitur laudabilis Domino.
LEV|19|25|Quinto autem anno comedetis fructus eorum, ut augeatur vobis proventus eorum. Ego Dominus Deus vester.
LEV|19|26|Non comedetis cum sanguine.Non augurabimini nec observabitis omina.
LEV|19|27|Neque in rotundum attondebitis marginem comae nec truncabis barbam.
LEV|19|28|Et super mortuo non incidetis carnem vestram neque figuras aliquas in cute incidetis vobis. Ego Dominus.
LEV|19|29|Ne polluas et prostituas filiam tuam, ne contaminetur terra et impleatur piaculo.
LEV|19|30|Sabbata mea custodite et sanctuarium meum metuite. Ego Dominus.
LEV|19|31|Non declinetis ad pythones nec ab hariolis aliquid sciscitemini, ut polluamini per eos. Ego Dominus Deus vester.
LEV|19|32|Coram cano capite consurge et honora personam senis; et time Deum tuum. Ego Dominus.
LEV|19|33|Si habitaverit tecum advena in terra vestra, non opprimetis eum;
LEV|19|34|sed sit inter vos quasi indigena, et diliges eum sicut teipsum: fuistis enim et vos advenae in terra Aegypti. Ego Dominus Deus vester.
LEV|19|35|Nolite facere iniquum aliquid in iudicio, in regula, in pondere, in mensura.
LEV|19|36|Statera iusta, aequa pondera, iustum ephi aequumque hin sint vobis. Ego Dominus Deus vester, qui eduxi vos de terra Aegypti.
LEV|19|37|Custodite omnia praecepta mea et universa iudicia et facite ea. Ego Dominus ".
LEV|20|1|Locutusque est Dominus ad Moysen dicens:
LEV|20|2|" Haec lo queris filiis Israel: Homo de filiis Israel et de advenis, qui habitant in Israel, si dederit de semine suo idolo Moloch, morte moriatur: populus terrae lapidabit eum.
LEV|20|3|Et ego ponam faciem meam contra illum; succidamque eum de medio populi sui, eo quod dederit de semine suo Moloch et contaminaverit sanctuarium meum ac polluerit nomen sanctum meum.
LEV|20|4|Quod si clauserit populus terrae oculos suos, ne videat hominem illum, qui dederit de semine suo Moloch, nec voluerit eum occidere,
LEV|20|5|ponam ego faciem meam super hominem illum et cognationem eius succidamque et ipsum et omnes, qui consenserunt ei, ut fornicarentur cum Moloch, de medio populi sui.
LEV|20|6|Anima, quae declinaverit ad pythones et hariolos et fornicata fuerit cum eis, ponam faciem meam contra eam et interficiam illam de medio populi sui.
LEV|20|7|Sanctificamini et estote sancti, quia ego Dominus Deus vester.
LEV|20|8|Custodite praecepta mea et facite ea. Ego Dominus, qui sanctifico vos.
LEV|20|9|Qui maledixerit patri suo et matri, morte moriatur; qui patri matrique maledixit, sanguis eius sit super eum.
LEV|20|10|Si moechatus quis fuerit cum uxore alterius et adulterium perpetrarit cum coniuge proximi sui, morte moriantur et moechus et adultera.
LEV|20|11|Qui dormierit cum noverca sua et revelaverit ignominiam patris sui, morte moriantur ambo: sanguis eorum sit super eos.
LEV|20|12|Si quis dormierit cum nuru sua, uterque moriatur, quia scelus operati sunt: sanguis eorum sit super eos.
LEV|20|13|Qui dormierit cum masculo coitu femineo, uterque operatus est nefas, morte moriantur: sit sanguis eorum super eos.
LEV|20|14|Qui supra uxorem filiam duxerit matrem eius, scelus operatus est: vivus ardebit cum eis, nec permanebit tantum nefas in medio vestri.
LEV|20|15|Qui cum iumento et pecore coierit, morte moriatur; pecus quoque occidite.
LEV|20|16|Mulier, quae succubuerit cuilibet iumento, simul interficies illam cum eo, morte moriantur: sanguis eorum sit super eos.
LEV|20|17|Qui acceperit sororem suam filiam patris sui vel filiam matris suae et viderit turpitudinem eius, illaque conspexerit fratris ignominiam, nefaria res est; occidentur in conspectu populi sui, eo quod turpitudinem sororis suae revelaverit, portabit iniquitatem suam.
LEV|20|18|Qui coierit cum muliere in fluxu menstruo et revelaverit turpitudinem eius ­ fontem eius nudavit, ipsaque aperuit fontem sanguinis sui ­ interficientur ambo de medio populi sui.
LEV|20|19|Turpitudinem materterae et amitae tuae non discooperies; qui hoc fecerit, ignominiam carnis suae nudavit; portabunt ambo iniquitatem suam.
LEV|20|20|Qui coierit cum uxore patrui vel avunculi sui et revelaverit ignominiam cognationis suae, portabunt ambo peccatum suum: absque liberis morientur.
LEV|20|21|Qui duxerit uxorem fratris sui, immunditia est, turpitudinem fratris sui revelavit: absque liberis erunt.
LEV|20|22|Custodite omnes leges meas atque omnia iudicia et facite ea, ne et vos evomat terra, quam intraturi estis et habitaturi.
LEV|20|23|Nolite ambulare in legitimis nationum, quas ego expulsurus sum ante vos. Omnia enim haec fecerunt, et abominatus sum eas
LEV|20|24|locutusque sum vobis: Vos possidebitis terram eorum, et ego dabo eam vobis in hereditatem, terram fluentem lacte et melle. Ego Dominus Deus vester, qui separavi vos a ceteris populis.
LEV|20|25|Separate ergo et vos iumentum mundum ab immundo et avem immundam a munda, ne polluatis animas vestras in pecore et in avibus et cunctis, quae moventur in terra, et quae vobis separavi tamquam immunda.
LEV|20|26|Eritis mihi sancti, quia sanctus sum ego Dominus et separavi vos a ceteris populis, ut essetis mei.
LEV|20|27|Vir sive mulier, in quibus pythonicus vel divinationis fuerit spiritus, morte moriantur; lapidibus obruent eos: sanguis eorum sit super illos ".
LEV|21|1|Dixit quoque Dominus ad Moysen: " Loquere ad sacer dotes filios Aaron et dices eis: Ne contaminetur sacerdos in mortibus civium suorum,
LEV|21|2|nisi tantum in consanguineis propinquis, id est super matre et patre et filio ac filia, fratre quoque
LEV|21|3|et sorore virgine propinqua, quae non est nupta viro; in ipsa contaminabitur.
LEV|21|4|Non contaminabitur ut maritus in cognatis suis, ne profanetur.
LEV|21|5|Non radent caput nec barbam neque in carne sua facient incisuras.
LEV|21|6|Sancti erunt Deo suo et non polluent nomen eius: incensa enim Domini et panem Dei sui offerunt et ideo sancti erunt.
LEV|21|7|Scortum et oppressam non ducent uxorem nec eam, quae repudiata est a marito, quia consecratus est Deo suo.
LEV|21|8|Et sanctificabis eum, quia panem Dei sui offert. Sit ergo sanctus tibi, quia ego sanctus sum, Dominus, qui sanctifico vos.
LEV|21|9|Sacerdotis filia, si profanaverit se stupro, profanat nomen patris sui; flammis exuretur.
LEV|21|10|Sacerdos maximus inter fratres suos, super cuius caput fusum est unctionis oleum, et cuius manus in sacerdotio consecratae sunt, vestitusque est sanctis vestibus, comam suam non excutiet, vestimenta non scindet
LEV|21|11|et ad omnem mortuum non ingredietur omnino; super patre quoque suo et matre non contaminabitur.
LEV|21|12|Nec egredietur de sanctuario, ne polluat sanctuarium Domini, quia consecratus est oleo unctionis Dei sui. Ego Dominus.
LEV|21|13|Virginem ducet uxorem;
LEV|21|14|viduam et repudiatam et oppressam atque meretricem non accipiet, sed virginem de cognatis suis ducet uxorem.
LEV|21|15|Ne profanet stirpem suam inter cognatos suos, quia ego Dominus, qui sanctifico eum ".
LEV|21|16|Locutusque est Dominus ad Moysen dicens:
LEV|21|17|" Loquere ad Aaron: Homo de semine tuo in generationibus suis, qui habuerit maculam, non accedet, ut offerat panem Dei sui;
LEV|21|18|quia quicumque habuerit maculam, non accedet: si caecus fuerit vel claudus, si mutilo naso vel deformis,
LEV|21|19|si fracto pede vel manu,
LEV|21|20|si gibbus, si pusillus, si albuginem habens in oculo, si iugem scabiem, si impetiginem in corpore vel contritos testiculos.
LEV|21|21|Omnis, qui habuerit maculam de semine Aaron sacerdotis, non accedet offerre incensa Domini nec panem Dei sui.
LEV|21|22|Vescetur tamen pane Dei sui de sanctissimis et de sanctis.
LEV|21|23|Sed ad velum non ingrediatur nec accedat ad altare, quia maculam habet et contaminare non debet sanctuaria mea, quia ego Dominus, qui sanctifico ea ".
LEV|21|24|Locutus est ergo Moyses ad Aaron et filios eius et ad omnem Israel.
LEV|22|1|Locutus quoque est Dominus ad Moysen dicens:
LEV|22|2|" Loquere ad Aaron et ad filios eius, ut caveant ab his, quae consecrata sunt filiorum Israel, et non contaminent nomen sanctum meum, quae ipsi offerunt mihi. Ego Dominus.
LEV|22|3|Dic ad eos pro posteris vestris: Omnis homo, qui accesserit de omni stirpe vestra ad sancta, quae consecraverunt filii Israel Domino, in immunditia sua, peribit coram me. Ego Dominus.
LEV|22|4|Homo de semine Aaron, qui fuerit leprosus aut patiens fluxum, non vescetur de his, quae sanctificata sunt, donec sanetur. Qui tetigerit omne, quod immundum est ex mor tuo, vel vir, ex quo egreditur semen,
LEV|22|5|et qui tangit reptile, quo polluitur, vel hominem, quo polluitur qualibet immunditia illius,
LEV|22|6|immundus erit usque ad vesperum et non vescetur his, quae sanctificata sunt; sed cum laverit carnem suam aqua,
LEV|22|7|et occubuerit sol, tunc mundatus vescetur de sanctificatis, quia cibus illius est.
LEV|22|8|Morticinum et dilaceratum a bestia non comedent, nec polluentur in eis. Ego Dominus.
LEV|22|9|Custodient praeceptum meum, ut non habeant super illo peccatum et propterea moriantur, cum polluerint illud; ego Dominus, qui sanctifico eos.
LEV|22|10|Omnis alienigena non comedet de sanctificatis, inquilinus sacerdotis et mercennarius non vescentur ex eis.
LEV|22|11|Quem autem sacerdos emerit, et qui vernaculus domus eius fuerit, hi comedent ex eis.
LEV|22|12|Si filia sacerdotis cuilibet ex populo nupta fuerit, de muneribus, quae sanctificata sunt, non vescetur;
LEV|22|13|sin autem vidua vel repudiata et absque liberis reversa fuerit ad domum patris sui, sicut puella consueverat, aletur cibo patris sui. Omnis alienigena comedendi ex eo non habet potestatem.
LEV|22|14|Qui comederit de sanctificatis per ignorantiam, addet quintam partem cum eo, quod comedit, et dabit sacerdoti sanctificatum.
LEV|22|15|Nec contaminabunt sanctificata filiorum Israel, quae tamquam munus offerunt Domino,
LEV|22|16|ne inducant super eos iniquitatem delicti, cum illi sanctificata sua comederint. Ego Dominus, qui sanctifico ".
LEV|22|17|Locutus est Dominus ad Moysen dicens:
LEV|22|18|" Loquere ad Aaron et filios eius et ad omnes filios Israel dicesque ad eos: Homo de domo Israel et de advenis, qui habitant apud vos, qui obtulerit oblationem suam vel vota solvens vel sponte offerens, quidquid illud obtulerit in holocaustum Domino,
LEV|22|19|in beneplacitum pro vobis offeratur masculus immaculatus ex bobus et ex ovibus et ex capris;
LEV|22|20|si maculam habuerit, non offeretis, quia non erit vobis acceptabile.
LEV|22|21|Homo, qui obtulerit victimam pacificorum Domino, vel vota solvens vel sponte offerens tam de bobus quam de ovibus immaculatum offeret, ut acceptabile sit; omnis macula non erit in eo.
LEV|22|22|Si caecum fuerit, si fractum, si mutilum, si verrucam habens aut scabiem vel impetiginem, non offeretis ea Domino nec in incensum dabitis ex eis super altare Domino.
LEV|22|23|Bovem et ovem deformem et debilem voluntarie offerre potes; votum autem ex his solvi non potest.
LEV|22|24|Omne animal, quod vel contritis vel tusis vel sectis ablatisque testiculis est, non offeretis Domino, et in terra vestra hoc omnino ne faciatis.
LEV|22|25|De manu alienigenae non offeretis cibum Dei vestri ex omnibus his animalibus, quia corrupta et maculata sunt omnia; non erunt in beneplacitum pro vobis ".
LEV|22|26|Locutusque est Dominus ad Moysen dicens:
LEV|22|27|" Bos, ovis et capra, cum genita fuerint, septem diebus erunt sub ubere matris suae; die autem octavo et deinceps erunt acceptabile munus incensi Domino.
LEV|22|28|Sive illa bos sive ovis non immolabuntur una die cum fetibus suis.
LEV|22|29|Si sacrificaveritis hostiam pro gratiarum actione Domino, sacrificabitis, ut possit esse placabilis.
LEV|22|30|Eodem die comedetis eam; non remanebit quidquam in mane alterius diei. Ego Dominus.
LEV|22|31|Custodite mandata mea et facite ea. Ego Dominus.
LEV|22|32|Ne polluatis nomen meum sanctum, ut sanctificer in medio filiorum Israel. Ego Dominus, qui sanctifico vos
LEV|22|33|et eduxi de terra Aegypti, ut essem vobis in Deum. Ego Dominus ".
LEV|23|1|Locutus est Dominus ad Moysen dicens:
LEV|23|2|" Loquere filiis Israel et dices ad eos: Hae sunt feriae Domini, quas vocabitis conventus sanctos; hae sunt feriae meae.
LEV|23|3|Sex diebus facietis opus; dies septimus sabbatum requiei est, conventus sanctus; omne opus non facietis; sabbatum est Domino in cunctis habitationibus vestris.
LEV|23|4|Hae sunt ergo feriae Domini, conventus sancti, quas celebrare debetis temporibus suis.
LEV|23|5|Mense primo, quarta decima die mensis, ad vesperum Pascha Domini est.
LEV|23|6|Et quinta decima die mensis huius sollemnitas Azymorum Domini est. Septem diebus azyma comedetis.
LEV|23|7|Die primo erit vobis conventus sanctus; omne opus servile non facietis in eo,
LEV|23|8|sed offeretis incensum Domino septem diebus. Die autem septimo erit conventus sanctus, nullumque servile opus facietis in eo ".
LEV|23|9|Locutusque est Dominus ad Moysen dicens:
LEV|23|10|" Loquere filiis Israel et dices ad eos: Cum ingressi fueritis terram, quam ego dabo vobis, et messueritis segetem, feretis manipulum spicarum primitias messis vestrae ad sacerdotem,
LEV|23|11|qui elevabit fasciculum coram Domino, ut acceptabile sit pro vobis; altero die sabbati sanctificabit illum.
LEV|23|12|Atque in eodem die, quo manipulum consecrabitis, facietis agnum immaculatum anniculum in holocaustum Domino,
LEV|23|13|et oblationem cum eo duas decimas similae conspersae oleo in incensum Domino odoremque suavissimum et libamentum eius vini quartam partem hin.
LEV|23|14|Panem et grana tosta farrem recentem non comedetis ex segete usque ad diem, qua offeretis ex ea munus Deo vestro. Praeceptum est sempiternum generationibus vestris in cunctis habitaculis vestris.
LEV|23|15|Numerabitis vobis ab altero die sabbati, in quo obtulistis manipulum elationis, septem hebdomadas plenas
LEV|23|16|usque ad alteram diem expletionis hebdomadae septimae, id est quinquaginta dies; et sic offeretis oblationem novam Domino
LEV|23|17|ex habitaculis vestris panes elationis duos de duabus decimis similae fermentatae, quos coquetis in primitias Domino;
LEV|23|18|offeretisque cum panibus septem agnos immaculatos anniculos et vitulum de armento unum et arietes duos, et erunt holocaustum Domino cum oblatione similae et libamentis suis in odorem suavissimum Domino.
LEV|23|19|Facietis et hircum in sacrificium pro peccato duosque agnos anniculos, hostias pacificorum.
LEV|23|20|Cumque elevaverit eos sacerdos cum panibus primitiarum coram Domino, cum duobus agnis sanctum erunt Domino in usum sacerdotis.
LEV|23|21|Et vocabitis hoc ipso die conventum, conventus sanctus erit vobis; omne opus servile non facietis in eo. Legitimum sempiternum erit in cunctis habitaculis generationibus vestris.
LEV|23|22|Cum autem metatis segetem terrae vestrae, non secabis eam usque ad oram agri nec remanentes spicas colliges, sed pauperibus et peregrinis dimittes eas. Ego Dominus Deus vester ".
LEV|23|23|Locutusque est Dominus ad Moysen dicens:
LEV|23|24|" Loquere filiis Israel: Mense septimo, prima die mensis, erit vobis requies, memoriale, clangentibus tubis, conventus sanctus.
LEV|23|25|Omne opus servile non facietis in eo et offeretis incensum Domino ".
LEV|23|26|Locutusque est Dominus ad Moysen dicens:
LEV|23|27|" Attamen decimo die mensis huius septimi dies Expiationum est, conventus sanctus erit vobis; affligetisque animas vestras in eo et offeretis incensum Domino.
LEV|23|28|Omne opus non facietis in tempore diei huius, quia dies expiationum est in expiationem vestram coram Domino Deo vestro.
LEV|23|29|Omnis anima, quae afflicta non fuerit die hoc, peribit de populis suis;
LEV|23|30|et,quae operis quippiam fecerit die hac, delebo eam de populo suo.
LEV|23|31|Nihil ergo operis facietis in eo: legitimum sempiternum erit vestris generationibus in cunctis habitationibus vestris.
LEV|23|32|Sabbatum requietionis est vobis, et affligetis animas vestras; die nono mensis a vespero usque ad vesperum servabitis sabbatum vestrum ".
LEV|23|33|Et locutus est Dominus ad Moysen dicens:
LEV|23|34|" Loquere filiis Israel: Quinto decimo die mensis huius septimi erit festum Tabernaculorum septem diebus Domino.
LEV|23|35|Die primo conventus sanctus, omne opus servile non facietis in eo;
LEV|23|36|septem diebus offeretis incensum Domino. Die octavo conventus sanctus erit vobis et offeretis incensum Domino; est enim coetus: omne opus servile non facietis.
LEV|23|37|Hae sunt feriae Domini, quas vocabitis conventus sanctos, offeretisque in eis incensum Domino, holocausta et oblationes similae, sacrificia et libamenta iuxta ritum uniuscuiusque diei;
LEV|23|38|praeter sabbata Domini donaque vestra et omnia, quae offeretis ex voto vel quae sponte tribuetis Domino.
LEV|23|39|Sed quinto decimo die mensis septimi, quando congregaveritis omnes fructus terrae, celebrabitis festum Domini septem diebus; die primo et die octavo erit requies.
LEV|23|40|Sumetisque vobis die primo fructus arboris pulcherrimos spatulasque palmarum et ramos ligni densarum frondium et salices de torrente et laetabimini coram Domino Deo vestro.
LEV|23|41|Celebrabitisque sollemnitatem eius septem diebus per annum: legitimum sempiternum erit generationibus vestris. Mense septimo festum celebrabitis
LEV|23|42|et habitabitis in umbraculis septem diebus; omnis, qui de genere est Israel, manebit in tabernaculis,
LEV|23|43|ut discant posteri vestri quod in tabernaculis habitare fecerim filios Israel, cum educerem eos de terra Aegypti. Ego Dominus Deus vester ".
LEV|23|44|Locutusque est Moyses super sollemnitatibus Domini ad filios Israel.
LEV|24|1|Et locutus est Dominus ad Moysen dicens:
LEV|24|2|" Praecipe fi liis Israel, ut afferant tibi oleum de olivis purissimum ac lucidum ad concinnandas lucernas candelabri iugiter.
LEV|24|3|Extra velum testimonii in tabernaculo conventus parabit illud Aaron a vespere usque ad mane coram Domino iugiter, ritu perpetuo in generationibus vestris.
LEV|24|4|Super candelabro mundissimo parabit lucernas semper in conspectu Domini.
LEV|24|5|Accipies quoque similam et coques ex ea duodecim panes, qui singuli habebunt duas decimas,
LEV|24|6|quorum senos altrinsecus super mensam purissimam coram Domino statues.
LEV|24|7|Et pones super ambas strues tus lucidissimum, ut sit panis in memoriale, incensum Domino.
LEV|24|8|Per singula sabbata mutabuntur coram Domino suscepti a filiis Israel; foedus sempiternum.
LEV|24|9|Eruntque Aaron et filiorum eius, ut comedant eos in loco sancto, quia sanctum sanctorum est ei de incensis Domini; iure perpetuo ".
LEV|24|10|Ecce autem egressus filius mulieris Israelitis, quem pepererat de viro Aegyptio inter filios Israel, iurgatus est in castris cum viro Israelita.
LEV|24|11|Cumque blasphemasset nomen et maledixisset ei, adductus est ad Moysen; vocabatur autem mater eius Salomith filia Dabri de tribu Dan.
LEV|24|12|Miseruntque eum in custodiam, donec nossent quid iuberet Dominus.
LEV|24|13|Qui locutus est ad Moysen dicens:
LEV|24|14|" Educ blasphemum extra castra, et ponant omnes, qui audierunt, manus suas super caput eius, et lapidet eum coetus universus.
LEV|24|15|Et ad filios Israel loqueris:Homo, qui maledixerit Deo suo, portabit peccatum suum;
LEV|24|16|et, qui blasphemaverit nomen Domini, morte moriatur: lapidibus opprimet eum omnis coetus, sive ille peregrinus sive civis fuerit. Qui blasphemaverit nomen Domini, morte moriatur.
LEV|24|17|Qui percusserit et occiderit hominem, morte moriatur.
LEV|24|18|Qui percusserit animal, reddet vicarium, id est animam pro anima.
LEV|24|19|Qui irrogaverit maculam cuilibet civium suorum, sicut fecit, sic fiet ei:
LEV|24|20|fracturam pro fractura, oculum pro oculo, dentem pro dente restituet; qualem inflixerit maculam, talem sustinere cogetur.
LEV|24|21|Qui percusserit iumentum, reddet aliud. Qui percusserit hominem, morietur.
LEV|24|22|Aequum iudicium sit inter vos, sive peregrinus sive civis peccaverit; quia ego sum Dominus Deus vester ".
LEV|24|23|Locutusque est Moyses ad filios Israel, et eduxerunt eum, qui blasphemaverat, extra castra, ac lapidibus oppresserunt. Feceruntque filii Israel, sicut praeceperat Dominus Moysi.
LEV|25|1|Locutusque est Dominus ad Moysen in monte Sinai di cens:
LEV|25|2|" Loquere filiis Israel et dices ad eos: Quando ingressi fueritis terram, quam ego dabo vobis, sabbatizet terra sabbatum Domino.
LEV|25|3|Sex annis seres agrum tuum et sex annis putabis vineam tuam colligesque fructus eius;
LEV|25|4|septimo autem anno, sabbatum requietionis erit terrae, sabbatum Domino: agrum tuum non seres et vineam tuam non putabis.
LEV|25|5|Quae sponte gignit humus, non metes et uvas vineae tuae non putatae non colliges quasi vindemiam; annus enim requietionis erit terrae.
LEV|25|6|Et erit sabbatum terrae vobis in cibum: tibi et servo tuo, ancillae et mercennario tuo et advenis, qui peregrinantur apud te,
LEV|25|7|iumentis tuis et animalibus, quae in terra tua sunt, omnia, quae nascuntur, praebebunt cibum.
LEV|25|8|Numerabis quoque tibi septem hebdomadas annorum, id est septem septies, quae simul faciunt annos quadraginta novem;
LEV|25|9|et clanges bucina mense septimo, decima die mensis expiationis die clangetis tuba in universa terra vestra.
LEV|25|10|Sanctificabitisque annum quinquagesimum et vocabitis remissionem in terra cunctis habitatoribus eius: ipse est enim iobeleus. Revertemini unusquisque ad possessionem suam, et unusquisque rediet ad familiam pristinam.
LEV|25|11|Iobeleus erit vobis quinquagesimus annus. Non seretis neque metetis sponte in agro nascentia neque vineas non putatas vindemiabitis
LEV|25|12|ob sanctificationem iobelei; sed de agro statim ablatas comedetis fruges.
LEV|25|13|Hoc anno iobelei rediet unusquisque vestrum ad possessionem suam.
LEV|25|14|Quando vendes quippiam civi tuo vel emes ab eo, ne contristet unusquisque fratrem suum; sed iuxta numerum annorum post iobeleum emes ab eo,
LEV|25|15|et iuxta supputationem annorum frugum vendet tibi.
LEV|25|16|Quanto plures anni remanserint post iobeleum, tanto crescet et pretium; et quanto minus temporis numeraveris, tanto minoris et emptio constabit: tempus enim frugum vendet tibi.
LEV|25|17|Nolite affligere contribules vestros, sed timeas Deum tuum, quia ego Dominus Deus vester.
LEV|25|18|Facite praecepta mea et iudicia, custodite et implete ea, ut habitare possitis in terra absque ullo pavore,
LEV|25|19|et gignat vobis humus fructus suos, quibus vescamini usque ad saturitatem, et habitabitis super terram, nullius impetum formidantes.
LEV|25|20|Quod si dixeritis: "Quid comedemus anno septimo, si non seruerimus neque collegerimus fruges nostras?".
LEV|25|21|Dabo benedictionem meam vobis anno sexto, et faciet fructus trium annorum,
LEV|25|22|seretisque anno octavo et comedetis veteres fruges usque ad nonum annum; donec nova nascantur, edetis vetera.
LEV|25|23|Terra quoque non veniet in perpetuum, quia mea est, et vos advenae et coloni mei estis.
LEV|25|24|Unde cuncta regio possessionis vestrae sub redemptionis condicione a vobis vendetur.
LEV|25|25|Si attenuatus frater tuus vendiderit partem possessionis suae, veniet ut redemptor propinquus eius, et redimet, quod ille vendiderat.
LEV|25|26|Sin autem non habuerit redemptorem et ipse pretium ad redimendum potuerit invenire,
LEV|25|27|computabuntur fructus ex eo tempore, quo vendidit; et, quod reliquum est, reddet emptori sicque recipiet possessionem suam.
LEV|25|28|Quod si non invenerit manus eius, ut reddat pretium, habebit emptor, quod emerat, usque ad annum iobeleum. In ipso enim omnis venditio rediet ad dominum et ad possessorem pristinum.
LEV|25|29|Qui vendiderit domum intra urbis muros, habebit licentiam redimendi, donec unus impleatur annus.
LEV|25|30|Si non redemerit, et anni circulus fuerit evolutus, emptor possidebit eam et posteri eius in perpetuum; et redimi non poterit, etiam in iobeleo.
LEV|25|31|Sin autem in villa fuerit domus, quae muros non habet, agrorum iure vendetur: potest redimi et in iobeleo revertetur ad dominum.
LEV|25|32|Aedes Levitarum, quae in urbibus possessionis eorum sunt, semper possunt ab eis redimi.
LEV|25|33|Si autem quis redemerit a Levitis, domus et urbs in iobeleo revertentur ad dominos; quia domus urbium leviticarum pro possessionibus eorum sunt inter filios Israel.
LEV|25|34|Suburbana autem pascua eorum non venient, quia possessio sempiterna est eis.
LEV|25|35|Si attenuatus fuerit frater tuus, et infirma manus eius apud te, suscipies eum quasi advenam et peregrinum, et vivet tecum.
LEV|25|36|Ne accipias usuras ab eo nec amplius quam dedisti: time Deum tuum, ut vivere possit frater tuus apud te.
LEV|25|37|Pecuniam tuam non dabis ei ad usuram nec plus aequo exiges pro cibo tuo.
LEV|25|38|Ego Dominus Deus vester, qui eduxi vos de terra Aegypti, ut darem vobis terram Chanaan et essem vester Deus.
LEV|25|39|Si paupertate compulsus vendiderit se tibi frater tuus, non eum opprimes servitute servorum,
LEV|25|40|sed quasi mercennarius et colonus erit tecum. Usque ad annum iobeleum operabitur apud te
LEV|25|41|et postea egredietur cum liberis suis et revertetur ad cognationem suam et ad possessionem patrum suorum.
LEV|25|42|Mei enim servi sunt, et ego eduxi eos de terra Aegypti: non venient condicione servorum;
LEV|25|43|ne affligas eum per po tentiam, sed metuito Deum tuum.
LEV|25|44|Servus et ancilla sint tibi de nationibus, quae in circuitu vestro sunt; de illis emetis servum et ancillam.
LEV|25|45|De filiis quoque advenarum, qui peregrinantur apud vos, emetis et de cognatione eorum, quae est apud vos et quam genuerint in terra vestra, hos habebitis in possessionem
LEV|25|46|et hereditario iure transmittetis ad posteros ac possidebitis in aeternum ut servos; fratres autem vestros filios Israel ne opprimatis cum potentia.
LEV|25|47|Si invaluerit apud vos manus advenae atque peregrini, et attenuatus frater tuus vendiderit se ei aut cuiquam de stirpe eius,
LEV|25|48|post venditionem potest redimi. Unus ex fratribus suis redimet eum
LEV|25|49|et patruus et patruelis et consanguineus et affinis. Sin autem et ipse potuerit, redimat se,
LEV|25|50|supputatis dumtaxat cum emptore annis a tempore venditionis suae usque ad annum iobeleum, et pecunia, qua venditus fuerat, iuxta annorum numerum et rationem mercennarii supputata.
LEV|25|51|Si plures fuerint anni, qui remanent usque ad iobeleum, secundum hos reddet et pretium redemptionis de pecunia emptionis;
LEV|25|52|si pauci, ponet rationem cum eo; iuxta annorum numerum reddet emptori, quod reliquum est annorum,
LEV|25|53|quibus ante servivit, mercedibus mercennarii imputatis. Non affliget eum violenter in conspectu tuo.
LEV|25|54|Quod si per haec redimi non potuerit, anno iobeleo egredietur cum liberis suis:
LEV|25|55|mei sunt enim servi filii Israel, quos eduxi de terra Aegypti. Ego Dominus Deus vester ".
LEV|26|1|" Non facietis vobis idolum et sculptile nec lapidem eri getis nec imaginem sculptam in petra ponetis in terra vestra, ut adoretis eam. Ego enim sum Dominus Deus vester.
LEV|26|2|Custodite sabbata mea et pavete sanctuarium meum. Ego Dominus.
LEV|26|3|Si in praeceptis meis ambulaveritis et mandata mea custodieritis et feceritis ea,
LEV|26|4|dabo vobis pluvias temporibus suis, et terra gignet germen suum, et pomis arbores replebuntur.
LEV|26|5|Apprehendet messium tritura vindemiam, et vindemia occupabit sementem; et comedetis panem vestrum in saturitatem et absque pavore habitabitis in terra vestra.
LEV|26|6|Dabo pacem in finibus vestris, dormietis, et non erit qui exterreat. Auferam malas bestias, et gladius non transibit per terminos vestros.
LEV|26|7|Persequemini inimicos vestros, et corruent coram vobis gladio.
LEV|26|8|Persequentur quinque de vestris centum alienos, et centum ex vobis decem milia; cadent inimici vestri in conspectu vestro gladio.
LEV|26|9|Respiciam vos et crescere faciam; multiplicabimini, et firmabo pactum meum vobiscum.
LEV|26|10|Comedetis vetusta congregata priorum messium; et vetera, novis supervenientibus, proicietis.
LEV|26|11|Ponam habitaculum meum in medio vestri, et non abominabitur vos anima mea.
LEV|26|12|Ambulabo inter vos et ero vester Deus, vosque eritis populus meus.
LEV|26|13|Ego Dominus Deus vester, qui eduxi vos de terra Aegyptiorum, ne serviretis eis, et qui confregi vectes iugi vestri, ut incederetis erecti.
LEV|26|14|Quod si non audieritis me nec feceritis omnia mandata haec,
LEV|26|15|si spreveritis leges meas, et iudicia mea contempserit anima vestra, ut non faciatis omnia, quae a me constituta sunt, et ad irritum perducatis pactum meum,
LEV|26|16|ego quoque haec faciam vobis: visitabo vos in terrore repentino, in tabe et ardore, qui conficiant oculos et consumant animam, frustra seretis sementem, quae ab hostibus devorabitur.
LEV|26|17|Ponam faciem meam contra vos, et corruetis coram hostibus vestris et subiciemini his, qui oderunt vos, et fugietis, nemine persequente.
LEV|26|18|Sin autem nec sic oboedieritis mihi, addam correptiones vestras septuplum propter peccata vestra
LEV|26|19|et conteram superbiam duritiae vestrae. Daboque caelum vobis desuper sicut ferrum et terram aeneam.
LEV|26|20|Consumetur incassum robur vestrum: non proferet terra germen, nec arbores poma praebebunt.
LEV|26|21|Si ambulaveritis ex adverso mihi nec volueritis audire me, addam plagas vestras usque in septuplum propter peccata vestra;
LEV|26|22|emittamque in vos bestias agri, quae absque liberis vos faciant et deleant pecora vestra et ad paucitatem vos redigant, desertaeque fiant viae vestrae.
LEV|26|23|Quod si nec sic volueritis recipere disciplinam, sed ambulaveritis ex adverso mihi,
LEV|26|24|ego quoque contra vos adversus incedam et percutiam vos septies propter peccata vestra.
LEV|26|25|inducamque super vos gladium ultorem foederis mei; cumque confugeritis in urbes vestras, mittam pestilentiam in medio vestri, et trademini hostium manibus.
LEV|26|26|Postquam confregero vobis baculum panis, coquent decem mulieres in uno clibano panem vestrum et reddent eum ad pondus, et comedetis et non saturabimini.
LEV|26|27|Sin autem nec per haec audieritis me, sed ambulaveritis contra me,
LEV|26|28|et ego incedam adversus vos in furore contrario; et corripiam vos septem plagis propter peccata vestra,
LEV|26|29|ita ut comedatis carnes filiorum et filiarum vestrarum.
LEV|26|30|Destruam excelsa vestra et thymiamateria confringam et ponam cadavera vestra super cadavera idolorum vestrorum, et abominabitur vos anima mea,
LEV|26|31|in tantum ut urbes vestras redigam in solitudinem et deserta faciam sanctuaria vestra nec recipiam ultra odorem suavissimum.
LEV|26|32|Disperdamque terram vestram; et stupebunt super ea inimici vestri, cum habitatores illius fuerint.
LEV|26|33|Vos autem dispergam in gentes et evaginabo post vos gladium; eritque terra vestra deserta et civitates dirutae.
LEV|26|34|Tunc placebunt terrae sabbata sua cunctis diebus solitudinis suae; quando fueritis in terra hostili, sabbatizabit et sabbata sua supplebit.
LEV|26|35|Cunctis diebus solitudinis sabbatizabit, eo quod non requieverit in sabbatis vestris, quando habitabatis in ea.
LEV|26|36|Et, qui de vobis remanserint, dabo pavorem in cordibus eorum in regionibus hostium; terrebit eos sonitus folii volantis, et ita fugient quasi gladium; cadent, nullo persequente.
LEV|26|37|Et corruent singuli super fratres suos quasi bella fugientes, nemine persequente. Nemo vestrum inimicis audebit resistere.
LEV|26|38|Peribitis inter gentes, et hostilis vos terra consumet.
LEV|26|39|Quod si et de vobis aliqui remanserint, tabescent in iniquitatibus suis in terris inimicorum vestrorum et propter peccata patrum suorum cum ipsis tabescent.
LEV|26|40|Et confitebuntur iniquitates suas et maiorum suorum, quibus praevaricati sunt in me et ambulaverunt ex adverso mihi,
LEV|26|41|ut et ego ambularem contra eos et inducerem illos in terram hostilem; vel tunc humiliabitur incircumcisum cor eorum, et tunc expiabunt pro impietatibus suis.
LEV|26|42|Et recordabor foederis mei, quod pepigi cum Iacob et Isaac et Abraham. Terrae quoque memor ero,
LEV|26|43|quae, cum relicta fuerit ab eis, complacebit sibi in sabbatis suis patiens solitudinem propter illos. Ipsi vero expiabunt pro peccatis suis, eo quod abiecerint iudicia mea et leges meas despexerint.
LEV|26|44|Et tamen, etiam cum essent in terra hostili, non penitus abieci eos neque sic despexi, ut consumerentur, et irritum facerem pactum meum cum eis. Ego enim sum Dominus, Deus eorum.
LEV|26|45|Et recordabor eis foederis cum maioribus, quos eduxi de terra Aegypti in conspectu gentium, ut essem Deus eorum. Ego Dominus ".
LEV|26|46|Haec sunt iudicia atque praecepta et leges, quas dedit Dominus inter se et inter filios Israel in monte Sinai per manum Moysi.
LEV|27|1|Locutusque est Dominus ad Moysen dicens:
LEV|27|2|" Loquere fi liis Israel et dices ad eos: Homo, qui votum fecerit et spoponderit Deo animas, sub aestimatione dabit pretium:
LEV|27|3|si fuerit masculus a vicesimo usque ad sexagesimum annum, dabit quinquaginta siclos argenti ad mensuram sanctuarii;
LEV|27|4|si mulier, triginta.
LEV|27|5|A quinto autem anno usque ad vicesimum masculus dabit viginti siclos, femina decem;
LEV|27|6|ab uno mense usque ad annum quintum pro masculo dabuntur quinque sicli, pro femina tres;
LEV|27|7|sexagenarius et ultra masculus dabit quindecim siclos, femina decem.
LEV|27|8|Si pauper fuerit et aestimationem reddere non valebit, sistet eum coram sacerdote, et quantum ille aestimaverit et viderit posse reddere, tantum dabit.
LEV|27|9|Animal autem, quod immolari potest Domino, si quis voverit, sanctum erit
LEV|27|10|et mutari non poterit, id est nec melius malo nec peius bono. Quod si mutaverit, et ipsum quod mutatum est et illud pro quo mutatum est, consecratum erit Domino.
LEV|27|11|Animal immundum, quod immolari Domino non potest, si quis voverit, adducetur ante sacerdotem,
LEV|27|12|qui diiudicans utrum bonum an malum sit, sicut statuet pretium, sic erit.
LEV|27|13|Quod si redimere illud voluerit is qui offert, addet supra aestimationem quintam partem.
LEV|27|14|Homo si voverit domum suam et sanctificaverit Domino, considerabit eam sacerdos utrum bona an mala sit, et iuxta pretium, quod ab eo fuerit constitutum, stabit.
LEV|27|15|Sin autem ille, qui voverat, voluerit redimere eam, dabit quintam partem aestimationis supra et habebit domum.
LEV|27|16|Quod si agrum possessionis suae voverit et consecraverit Domino, iuxta mensuram sementis aestimabitur pretium: si triginta homer hordei seritur terra, quinquaginta siclis aestimabitur argenti.
LEV|27|17|Si statim ab anno iobelei voverit agrum, quanto valere potest, tanto aestimabitur.
LEV|27|18|Sin autem post aliquantum temporis, supputabit ei sacerdos pecuniam iuxta annorum, qui reliqui sunt, numerum usque ad iobeleum, et detrahetur ex pretio.
LEV|27|19|Quod si voluerit redimere agrum ille, qui voverat, addet quintam partem aestimatae pecuniae et possidebit eum.
LEV|27|20|Sin autem noluerit redimere, sed alteri cuilibet vendiderit, ultra redimi non poterit;
LEV|27|21|sed, cum iobelei venerit dies, sanctum erit Domino sicut ager anathematis; sacerdotis erit possessio eius.
LEV|27|22|Quod si agrum emptum, qui non est de possessione maiorum, sanctificare voluerit Domino,
LEV|27|23|supputabit ei sacerdos iuxta annorum numerum usque ad iobeleum pretium, quod dabit ille, qui voverat, in ipso die ut sanctum Domino.
LEV|27|24|In anno autem iobelei revertetur ager ad priorem dominum, qui vendiderat eum et habuerat in sortem possessionis suae.
LEV|27|25|Omnis aestimatio siclo sanctuarii ponderabitur; siclus viginti gera habet.
LEV|27|26|Primogenita, quae de animalibus ad Dominum pertinent, nemo sanctificare poterit et vovere: sive bos sive ovis fuerit, Domini sunt.
LEV|27|27|Quod si immundum est animal, redimet, qui obtulit, iuxta aestimationem et addet quintam partem pretii; si redimere noluerit, vendetur quanto fuerit.
LEV|27|28|Omne anathema, quod aliquis vir consecrat Domino de omni possessione sua, sive homo fuerit sive animal sive ager, non veniet nec redimi poterit; quidquid semel fuerit consecratum, sanctum sanctorum erit Domino.
LEV|27|29|Et omnis homo, qui ut anathema offertur, non redimetur, sed morte morietur.
LEV|27|30|Omnes decimae terrae sive de frugibus sive de pomis arborum Domini sunt, sanctum Domino.
LEV|27|31|Si quis autem voluerit redimere aliquid de decimis suis, addet quintam partem.
LEV|27|32|Omnes decimae boves et oves et caprae, quae sub pastoris virga transeunt, quidquid decimum venerit, erit sanctum Domino.
LEV|27|33|Non discernetur inter bonum et malum nec altero commutabitur; si quis mutaverit, et quod mutatum est et pro quo mutatum est, sanctum erit et non redimetur ".
LEV|27|34|Haec sunt praecepta, quae mandavit Dominus Moysi ad filios Israel in monte Sinai.
NUM|1|1|Locutusque est Dominus ad Moysen in deserto Sinai in ta bernaculo conventus, prima die mensis secundi, anno altero egressionis eorum ex Aegypto, dicens:
NUM|1|2|" Tollite summam universae congregationis filiorum Israel per cognationes et domos suas et nomina singulorum, quidquid sexus est masculini
NUM|1|3|a vicesimo anno et supra omnium ex Israel, qui possunt ad bella procedere, et numerabitis eos per turmas suas, tu et Aaron.
NUM|1|4|Eritque vobiscum vir per tribum, princeps domus patrum suorum,
NUM|1|5|quorum ista sunt nomina: de Ruben Elisur filius Sedeur;
NUM|1|6|de Simeon Salamiel filius Surisaddai;
NUM|1|7|de Iuda Naasson filius Aminadab;
NUM|1|8|de Issachar Nathanael filius Suar;
NUM|1|9|de Zabulon Eliab filius Helon.
NUM|1|10|Filiorum autem Ioseph: de Ephraim Elisama filius Ammiud; de Manasse Gamaliel filius Phadassur.
NUM|1|11|De Beniamin Abidan filius Gedeonis;
NUM|1|12|de Dan Ahiezer filius Ammisaddai;
NUM|1|13|de Aser Phegiel filius Ochran;
NUM|1|14|de Gad Eliasaph filius Deuel;
NUM|1|15|de Nephthali Ahira filius Enan ".
NUM|1|16|Hi viri nobilissimi congregationis principes tribuum patrum suorum et capita milium Israel.
NUM|1|17|Quos tulerunt Moyses et Aaron nominatim designatos
NUM|1|18|et omnem congregationem congregaverunt primo die mensis secundi recensentes eos per cognationes et domos patrum eorum, per nomina singulorum a vicesimo anno et supra per capita,
NUM|1|19|sicut praeceperat Dominus Moysi. Numeratique sunt in deserto Sinai.
NUM|1|20|De Ruben primogenito Israelis generationes per familias ac domos patrum suorum, per nomina capitum singulorum omne quod sexus est masculini a vicesimo anno et supra procedentium ad bellum.
NUM|1|21|Recensiti tribus Ruben quadraginta sex milia quingenti.
NUM|1|22|De filiis Simeon generationes per familias ac domos cognationum suarum recensiti sunt per nomina et capita singulorum omne quod sexus est masculini a vicesimo anno et supra procedentium ad bellum.
NUM|1|23|Recensiti tribus Simeon quinquaginta novem milia trecenti.
NUM|1|24|De filiis Gad generationes per familias ac domos cognationum suarum recensiti sunt per nomina singulorum a viginti annis et supra omnes, qui ad bella procederent,
NUM|1|25|quadraginta quinque milia sescenti quinquaginta.
NUM|1|26|De filiis Iudae generationes per familias ac domos cognationum suarum per nomina singulorum a vicesimo anno et supra omnes, qui poterant ad bella procedere,
NUM|1|27|recensiti sunt septuaginta quattuor milia sescenti.
NUM|1|28|De filiis Issachar generationes per familias ac domos cognationum suarum per nomina singulorum a vicesimo anno et supra omnes, qui ad bella procederent,
NUM|1|29|recensiti sunt quinquaginta quattuor milia quadringenti.
NUM|1|30|De filiis Zabulon generationes per familias ac domos cognationum suarum recensiti sunt per nomina singulorum a vicesimo anno et supra omnes, qui poterant ad bella procedere,
NUM|1|31|quinquaginta septem milia quadringenti.
NUM|1|32|De filiis Ioseph filiorum Ephraim generationes per familias ac domos cognationum suarum recensiti sunt per nomina singulorum a vicesimo anno et supra omnes, qui poterant ad bella procedere,
NUM|1|33|quadraginta milia quingenti.
NUM|1|34|Porro filiorum Manasse generationes per familias ac domos cognationum suarum recensiti sunt per nomina singulorum a viginti annis et supra omnes, qui poterant ad bella procedere,
NUM|1|35|triginta duo milia ducenti.
NUM|1|36|De filiis Beniamin generationes per familias ac domos cognationum suarum recensiti sunt nominibus singulorum a vicesimo anno et supra omnes, qui poterant ad bella procedere,
NUM|1|37|triginta quinque milia quadringenti.
NUM|1|38|De filiis Dan generationes per familias ac domos cognationum suarum recensiti sunt nominibus singulorum a vicesimo anno et supra omnes, qui poterant ad bella procedere,
NUM|1|39|sexaginta duo milia septingenti.
NUM|1|40|De filiis Aser generationes per familias ac domos cognationum suarum recensiti sunt per nomina singulorum a vicesimo anno et supra omnes, qui poterant ad bella procedere,
NUM|1|41|quadraginta milia et mille quingenti.
NUM|1|42|De filiis Nephthali generationes per familias ac domos cognationum suarum recensiti sunt nominibus singulorum a vicesimo anno et supra omnes, qui poterant ad bella procedere,
NUM|1|43|quinquaginta tria milia quadringenti.
NUM|1|44|Hi sunt quos numeraverunt Moyses et Aaron et duodecim principes Israel, singuli per domos patrum suorum.
NUM|1|45|Fueruntque omnis numerus filiorum Israel per domos patrum suorum a vicesimo anno et supra, qui poterant ad bella procedere,
NUM|1|46|sescenta tria milia virorum quingenti quinquaginta.
NUM|1|47|Levitae autem in tribu patrum suorum non sunt numerati cum eis.
NUM|1|48|Locutusque est Dominus ad Moysen dicens:
NUM|1|49|" Tribum Levi noli numerare neque pones summam eorum cum filiis Israel,
NUM|1|50|sed constitue eos super habitaculum testimonii et cuncta vasa eius et quidquid ad caeremonias pertinet. Ipsi portabunt habitaculum et omnia utensilia eius et erunt in ministerio ac per gyrum habitaculi metabuntur.
NUM|1|51|Cum proficiscendum fuerit, deponent Levitae habitaculum; cum castrametandum, erigent; quisquis externorum accesserit, occidetur.
NUM|1|52|Metabuntur autem castra filii Israel, unusquisque per turmas et cuneos atque exercitum suum.
NUM|1|53|Porro Levitae per gyrum habitaculi testimonii figent tentoria, ne fiat indignatio super congregationem filiorum Israel, et excubabunt in custodiis habitaculi testimonii ".
NUM|1|54|Fecerunt ergo filii Israel iuxta omnia, quae praeceperat Dominus Moysi.
NUM|2|1|Locutusque est Dominus ad Moysen et Aaron dicens:
NUM|2|2|" Singuli per turmas, signa atque vexilla et domos patrum suorum castrametabuntur filii Israel per gyrum tabernaculi conventus.
NUM|2|3|Ad orientem Iudas figet tentoria per turmas exercitus sui, fuitque princeps filiorum eius Naasson filius Aminadab;
NUM|2|4|et eius summa pugnantium septuaginta quattuor milia sescenti.
NUM|2|5|Iuxta eum castrametabuntur de tribu Issachar, quorum princeps fuit Nathanael filius Suar;
NUM|2|6|et omnis numerus pugnatorum eius quinquaginta quattuor milia quadringenti.
NUM|2|7|In tribu Zabulon princeps fuit Eliab filius Helon;
NUM|2|8|et numerus exercitus pugnatorum eius quinquaginta septem milia quadringenti.
NUM|2|9|Universi, qui in castris Iudae annumerati sunt, fuerunt centum octoginta sex milia quadringenti, et per turmas suas primi egredientur.
NUM|2|10|Vexillum castrorum Ruben ad meridianam plagam erit, secundum exercitus eorum; princeps Elisur filius Sedeur;
NUM|2|11|et cunctus exercitus pugnatorum eius, qui numerati sunt, quadraginta sex milia quingenti.
NUM|2|12|Iuxta eum castrametabuntur de tribu Simeon, quorum princeps fuit Salamiel filius Surisaddai;
NUM|2|13|et cunctus exercitus pugnatorum eius, qui numerati sunt, quinquaginta novem milia trecenti.
NUM|2|14|In tribu Gad princeps fuit Eliasaph filius Deuel;
NUM|2|15|et cunctus exercitus pugnatorum eius, qui numerati sunt, quadraginta quinque milia sescenti quinquaginta.
NUM|2|16|Omnes, qui recensiti sunt in castris Ruben, centum quinquaginta milia et mille quadringenti quinquaginta, per turmas suas in secundo loco proficiscentur.
NUM|2|17|Levabitur deinde tabernaculum conventus, castra Levitarum in medio castrorum, quomodo erigetur ita et deponetur; singuli per loca et vexilla sua proficiscentur.
NUM|2|18|Ad occidentalem plagam erit vexillum castrorum filiorum Ephraim per turmas suas, quorum princeps fuit Elisama filius Ammiud;
NUM|2|19|cunctus exercitus pugnatorum eius, qui numerati sunt, quadraginta milia quingenti.
NUM|2|20|Et cum eis tribus filiorum Manasse, quorum princeps fuit Gamaliel filius Phadassur;
NUM|2|21|cunctusque exercitus pugnatorum eius, qui numerati sunt, triginta duo milia ducenti.
NUM|2|22|In tribu filiorum Beniamin princeps fuit Abidan filius Gedeonis;
NUM|2|23|et cunctus exercitus pugnatorum eius, qui recensiti sunt, triginta quinque milia quadringenti.
NUM|2|24|Omnes, qui numerati sunt in castris Ephraim, centum octo milia centum, per turmas suas tertii proficiscentur.
NUM|2|25|Ad aquilonis partem stabit vexillum castrorum filiorum Dan secundum exercitus suos, quorum princeps fuit Ahiezer filius Ammisaddai;
NUM|2|26|cunctus exercitus pugnatorum eius, qui numerati sunt, sexaginta duo milia septingenti.
NUM|2|27|Iuxta eum figet tentoria tribus Aser, quorum princeps fuit Phegiel filius Ochran;
NUM|2|28|cunctus exercitus pugnatorum eius, qui numerati sunt, quadraginta milia et mille quingenti.
NUM|2|29|De tribu filiorum Nephthali princeps fuit Ahira filius Enan;
NUM|2|30|cunctus exercitus pugnatorum eius quinquaginta tria milia quadringenti.
NUM|2|31|Omnes, qui numerati sunt in castris Dan, fuerunt centum quinquaginta septem milia sescenti, et novissimi proficiscentur secundum vexilla sua ".
NUM|2|32|Hic numerus filiorum Israel, per domos patrum suorum omnes recensiti secundum exercitus suos, sescenta tria milia quingenti quinquaginta.
NUM|2|33|Levitae autem non sunt numerati inter filios Israel; sic enim praeceperat Dominus Moysi.
NUM|2|34|Feceruntque filii Israel iuxta omnia, quae mandaverat Dominus: castrametati sunt per vexilla sua et profecti per tribus ad domos patrum suorum.
NUM|3|1|Hae sunt generationes Aaron et Moysi in die, qua locutus est Dominus ad Moysen in monte Sinai.
NUM|3|2|Et haec nomina filiorum Aaron: primogenitus eius Nadab, deinde Abiu et Eleazar et Ithamar.
NUM|3|3|Haec nomina filiorum Aaron sacerdotum, qui uncti sunt et quorum repletae manus, ut sacerdotio fungerentur.
NUM|3|4|Mortui sunt enim Nadab et Abiu, cum offerrent ignem alienum in conspectu Domini in deserto Sinai, absque liberis; functique sunt sacerdotio Eleazar et Ithamar coram Aaron patre suo.
NUM|3|5|Locutusque est Dominus ad Moysen dicens:
NUM|3|6|" Applica tribum Levi et fac stare in conspectu Aaron sacerdotis, ut ministrent ei
NUM|3|7|et observent, quidquid ad eum pertinet et ad totam congregationem coram tabernaculo conventus, servientes in ministerio habitaculi,
NUM|3|8|et custodiant vasa tabernaculi conventus explentes officia filiorum Israel, servientes in ministerio habitaculi.
NUM|3|9|Dabisque dono Levitas Aaron et filiis eius, quibus traditi sunt a filiis Israel;
NUM|3|10|Aaron autem et filios eius constitues super cultum sacerdotii. Externus, qui ad ministrandum accesserit, morietur ".
NUM|3|11|Locutusque est Dominus ad Moysen dicens:
NUM|3|12|" Ecce ego tuli Levitas a filiis Israel pro omni primogenito, qui aperit vulvam in filiis Israel; eruntque Levitae mei.
NUM|3|13|Meum est enim omne primogenitum: ex quo percussi omnes primogenitos in terra Aegypti, sanctificavi mihi, quidquid primum nascitur in Israel ab homine usque ad pecus; mei sunt. Ego Dominus ".
NUM|3|14|Locutusque est Dominus ad Moysen in deserto Sinai dicens:
NUM|3|15|" Numera filios Levi per domos patrum suorum et familias omnem masculum ab uno mense et supra ".
NUM|3|16|Numeravit eos Moyses, ut praeceperat Dominus,
NUM|3|17|et inventi sunt filii Levi per nomina sua Gerson et Caath et Merari.
NUM|3|18|Haec sunt nomina filiorum Gerson secundum familias suas: Lobni et Semei;
NUM|3|19|filii Caath secundum familias suas: Amram et Isaar, Hebron et Oziel;
NUM|3|20|filii Merari secundum familias suas: Moholi et Musi. Hae sunt familiae Levi per domos patrum suorum.
NUM|3|21|De Gerson fuere familiae duae Lobnitica et Semeitica,
NUM|3|22|quarum numeratus est omnis populus sexus masculini ab uno mense et supra septem milia quingenti.
NUM|3|23|Hi post habitaculum metabantur ad occidentem
NUM|3|24|sub principe Eliasaph filio Lael;
NUM|3|25|et habebant excubias in tabernaculo conventus, ipsum habitaculum et tabernaculum, operimentum eius, velum, quod trahitur ante fores tabernaculi conventus,
NUM|3|26|et cortinas atrii, velum quoque, quod appenditur in introitu atrii, quod est circa habitaculum et circa altare, et funes ad omne opus eius.
NUM|3|27|Caath habet familias: Amramitas et Isaaritas et Hebronitas et Ozielitas; hae sunt familiae Caathitarum.
NUM|3|28|Omnes generis masculini ab uno mense et supra octo milia sescenti habebant excubias sanctuarii.
NUM|3|29|Familiae filiorum Caath castrametabantur ad latus habitaculi ad meridianam plagam,
NUM|3|30|princepsque eorum erat Elisaphan filius Oziel.
NUM|3|31|Et custodiebant arcam mensamque et candelabrum, altaria et vasa sanctuarii, in quibus ministratur, et velum cunctamque huiuscemodi supellectilem.
NUM|3|32|Princeps autem principum Levitarum Eleazar filius Aaron sacerdotis erat super excubitores custodiae sanctuarii.
NUM|3|33|At vero de Merari erant familiae Moholitae et Musitae.
NUM|3|34|Omnes generis masculini ab uno mense et supra sex milia ducenti;
NUM|3|35|princeps familiarum Merari Suriel filius Abihail. In plaga septentrionali ad latus habitaculi castrametabantur;
NUM|3|36|erant sub custodia eorum tabulae habitaculi et vectes et columnae ac bases earum et cuncta vasa eius et omnia, quae ad cultum huiuscemodi pertinent,
NUM|3|37|columnaeque atrii per circuitum cum basibus suis et paxilli cum funibus.
NUM|3|38|Castrametabantur ante habitaculum, ad orientalem plagam ante tabernaculum conventus ad orientem, Moyses et Aaron cum filiis suis habentes custodiam sanctuarii in medio filiorum Israel. Quisquis alienus accesserit, morietur.
NUM|3|39|Omnes Levitae, quos numeravit Moyses iuxta praeceptum Domini per familias suas in genere masculino a mense uno et supra, fuerunt viginti duo milia.
NUM|3|40|Et ait Dominus ad Moysen: " Numera omnes primogenitos sexus masculini de filiis Israel ab uno mense et supra et habebis summam eorum;
NUM|3|41|tollesque Levitas mihi pro omni primogenito filiorum Israel ­ ego sum Dominus ­ et pecora eorum pro universis primogenitis pecorum filiorum Israel ".
NUM|3|42|Recensuit Moyses, sicut praeceperat Dominus, omnes primogenitos filiorum Israel,
NUM|3|43|et fuerunt omnes masculi per nomina sua a mense uno et supra viginti duo milia ducenti septuaginta tres.
NUM|3|44|Locutusque est Dominus ad Moysen dicens:
NUM|3|45|" Tolle Levitas pro omnibus primogenitis filiorum Israel et pecora Levitarum pro pecoribus corum; eruntque Levitae mei. Ego sum Dominus.
NUM|3|46|In pretio autem ducentorum septuaginta trium, qui excedunt numerum Levitarum de primogenitis filiorum Israel,
NUM|3|47|accipies quinque siclos per singula capita, ad mensuram sanctuarii. Siclus habet viginti obolos.
NUM|3|48|Dabisque pecuniam Aaron et filiis eius pretium eorum, qui supra sunt ".
NUM|3|49|Tulit igitur Moyses pecuniam eorum, qui excesserant numerum eorum, qui redempti erant a Levitis;
NUM|3|50|a primogenitis filiorum Israel tulit pecuniam mille trecentorum sexaginta quinque siclorum iuxta pondus sanctuarii.
NUM|3|51|Et dedit eam Aaron et filiis eius iuxta verbum, quod praeceperat sibi Dominus.
NUM|4|1|Locutusque est Dominus ad Moysen et Aaron dicens:
NUM|4|2|" Tolle summam filiorum Caath de medio Levitarum per familias et domos suas
NUM|4|3|a tricesimo anno et supra usque ad quinquagesimum annum omnium, qui ingrediuntur, ut stent et ministrent in tabernaculo conventus.
NUM|4|4|Hic est cultus filiorum Caath in tabernaculo conventus: sanctum sanctorum.
NUM|4|5|Ingredientur Aaron et filii eius, quando movenda sunt castra, et deponent velum, quod pendet ante fores, involventque eo arcam testimonii;
NUM|4|6|et operient rursum velamine pellium delphini extendentque desuper pallium totum hyacinthinum et inducent vectes.
NUM|4|7|Mensam quoque propositionis involvent hyacinthino pallio et ponent cum ea acetabula et phialas, cyathos et crateras ad liba fundenda; panes semper in ea erunt.
NUM|4|8|Extendentque desuper pallium coccineum, quod rursum operient velamento pellium delphini et inducent vectes.
NUM|4|9|Sument et pallium hyacinthinum, quo operient candelabrum cum lucernis et forcipibus suis et emunctoriis et cunctis vasis olei, quae ad concinnandas lucernas necessaria sunt;
NUM|4|10|et super omnia ponent operimentum pellium delphini et ponent super feretrum.
NUM|4|11|Nec non et altare aureum involvent hyacinthino vestimento et extendent desuper operimentum pellium delphini et inducent vectes.
NUM|4|12|Omnia vasa, quibus ministratur in sanctuario, involvent hyacinthino pallio; et extendent desuper operimentum pellium delphini ponentque super feretrum.
NUM|4|13|Sed et altare mundabunt cinere et involvent illud purpureo vestimento;
NUM|4|14|ponentque super illud omnia vasa, quibus in ministerio eius utuntur, id est ignium receptacula, fuscinulas ac vatilla et pateras. Cuncta vasa altaris operient simul velamine pellium delphini et inducent vectes.
NUM|4|15|Cumque involverint Aaron et filii eius sanctuarium et omnia vasa eius in commotione castrorum, tunc intrabunt filii Caath, ut portent involuta, et non tangent sanctuarium, ne moriantur. Ista sunt onera filiorum Caath in tabernaculo conventus.
NUM|4|16|Ad curam Eleazari filii Aaron sacerdotis pertinet oleum ad concinnandas lucernas et gratissimum incensum et oblatio, quae semper offertur, et oleum unctionis et quidquid ad cultum habitaculi pertinet omniumque vasorum, quae in sanctuario sunt ".
NUM|4|17|Locutusque est Dominus ad Moysen et Aaron dicens:
NUM|4|18|" Nolite perdere populum Caath de medio Levitarum,
NUM|4|19|sed hoc facite eis, ut vivant et non moriantur, quando appropinquant ad sancta sanctorum: Aaron et filii eius intrabunt ipsique disponent opera singulorum et divident quid portare quis debeat.
NUM|4|20|Non intrabunt ad videndum, nec puncto quidem, sanctuarium; alioquin morientur ".
NUM|4|21|Locutusque est Dominus ad Moysen dicens:
NUM|4|22|" Tolle summam etiam filiorum Gerson per domos ac familias et cognationes suas;
NUM|4|23|a triginta annis et supra usque ad annos quinquaginta numera omnes, qui ingrediuntur et ministrant in tabernaculo conventus.
NUM|4|24|Hoc est officium familiarum Gersonitarum,
NUM|4|25|ut portent cortinas habitaculi, tabernaculum conventus, operimentum eius et super illud velamen delphini velumque, quod pendet in introitu tabernaculi conventus,
NUM|4|26|cortinas atrii et velum in introitu atrii, quod est circa habitaculum et altare, funiculos et vasa ministerii, omnia, quae facta sunt, ut eis laborent.
NUM|4|27|Iubente Aaron et filiis eius, portabunt filii Gerson, et scient singuli cui debeant oneri mancipari.
NUM|4|28|Hic est cultus familiarum Gersonitarum in tabernaculo conventus; eruntque sub manu Ithamar filii Aaron sacerdotis.
NUM|4|29|Filios quoque Merari per familias et domos patrum suorum recensebis
NUM|4|30|a triginta annis et supra usque ad annos quinquaginta, omnes, qui ingrediuntur ad officium ministerii sui et cultum tabernaculi conventus.
NUM|4|31|Haec sunt onera eorum: portabunt tabulas habitaculi et vectes eius, columnas ac bases earum,
NUM|4|32|columnas quoque atrii per circuitum cum basibus et paxillis et funibus suis; omnia vasa et supellectilem ad numerum accipient sicque portabunt.
NUM|4|33|Hoc est officium familiarum Meraritarum et ministerium in tabernaculo conventus; eruntque sub manu Ithamar filii Aaron sacerdotis ".
NUM|4|34|Recensuerunt igitur Moyses et Aaron et principes synagogae filios Caath per cognationes et domos patrum suorum
NUM|4|35|a triginta annis et supra usque ad annum quinquagesimum, omnes, qui ingrediuntur ad ministerium tabernaculi conventus;
NUM|4|36|et inventi sunt duo milia septingenti quinquaginta.
NUM|4|37|Hic est numerus familiarum Caath, qui ministrant in tabernaculo conventus: hos numeravit Moyses et Aaron iuxta sermonem Domini per manum Moysi.
NUM|4|38|Numerati sunt et filii Gerson per cognationes et domos patrum suorum
NUM|4|39|a triginta annis et supra usque ad quinquagesimum annum, omnes, qui ingrediuntur, ut ministrent in tabernaculo conventus;
NUM|4|40|et inventi sunt secundum familias et domus patrum suorum duo milia sescenti triginta.
NUM|4|41|Hic est numerus Gersonitarum, omnes, qui ministrant in tabernaculo conventus, quos numeraverunt Moy ses et Aaron iuxta verbum Domini.
NUM|4|42|Numeratae sunt et familiae filiorum Merari per cognationes et domos patrum suorum
NUM|4|43|a triginta annis et supra usque ad annum quinquagesimum, omnes, qui ingrediuntur ad explendos ritus tabernaculi conventus;
NUM|4|44|et inventi sunt tria milia ducenti.
NUM|4|45|Hic est numerus familiarum filiorum Merari, quos recensuerunt Moyses et Aaron iuxta imperium Domini per manum Moysi.
NUM|4|46|Omnes, qui recensiti sunt de Levitis et quos recenseri fecit ad nomen Moyses et Aaron et principes Israel per cognationes et domos patrum suorum
NUM|4|47|a triginta annis et supra usque ad annum quinquagesimum ingredientes ad ministerium tabernaculi et onera portanda in tabernaculo conventus,
NUM|4|48|fuerunt simul octo milia quingenti octoginta. 49 Iuxta verbum Domini per manum Moysi recensuit eos unumquemque iuxta officium et onera sua, sicut praeceperat ei Dominus.
NUM|5|1|Locutusque est Dominus ad Moysen dicens:
NUM|5|2|" Praecipe filiis Israel, ut eiciant de castris omnem leprosum et qui semine fluit pollutusque est super mortuo.
NUM|5|3|Tam masculum quam feminam eicite de castris, ne contaminent ea, cum habitaverim cum eis ".
NUM|5|4|Feceruntque ita filii Israel et eiecerunt eos extra castra, sicut locutus erat Dominus Moysi.
NUM|5|5|Locutusque est Dominus ad Moysen dicens:
NUM|5|6|" Loquere ad filios Israel: Vir sive mulier, cum fecerint ex omnibus peccatis, quae solent hominibus accidere, et fraude transgressi fuerint mandatum Domini, ille homo reus erit;
NUM|5|7|et confitebuntur peccatum suum et reddent ipsum caput quintamque partem desuper ei, in quem peccaverint.
NUM|5|8|Sin autem non fuerit qui recipiat, dabunt Domino, et erit sacerdotis, praeter arietem, qui offertur pro expiatione, ut sit placabilis hostia.
NUM|5|9|Omnis quoque praelibatio rerum sacrarum, quas offerunt filii Israel, ad sacerdotem pertinet;
NUM|5|10|et, quidquid in sanctuarium offertur a singulis et traditur manibus sacerdotis, ipsius erit ".
NUM|5|11|Locutusque est Dominus ad Moysen dicens:
NUM|5|12|" Loquere ad filios Israel et dices ad eos: Vir, cuius uxor erraverit maritumque decipiens
NUM|5|13|dormierit cum altero viro, et hoc maritus deprehendere non quiverit, sed latet quod impuram se reddiderit et testibus argui non potest, quia non est inventa in stupro,
NUM|5|14|si spiritus zelotypiae concitaverit virum contra uxorem suam, quae vel polluta est vel falsa suspicione appetitur,
NUM|5|15|adducet eam ad sacerdotem et offeret oblationem pro illa decimam partem ephi farinae hordeaceae. Non fundet super eam oleum nec imponet tus, quia sacrificium zelotypiae est et oblatio investigans adulterium.
NUM|5|16|Afferet igitur eam sacerdos et statuet coram Domino;
NUM|5|17|assumetque aquam sanctam in vase fictili et pauxillum terrae de pavimento habitaculi mittet in eam.
NUM|5|18|Cumque posuerit sacerdos mulierem in conspectu Domini, discooperiet caput eius et ponet super manus illius sacrificium recordationis, oblationem zelotypiae; ipse autem tenebit aquas amarissimas, in quibus cum exsecratione maledicta congessit.
NUM|5|19|Adiurabitque eam et dicet: "Si non dormivit vir alienus tecum, et si non declinasti a viro tuo et non polluta es, deserto mariti toro, non te nocebunt aquae istae amarissimae, in quas maledicta congessi.
NUM|5|20|Sin autem declinasti a viro tuo atque polluta es et concubuisti cum altero viro",
NUM|5|21|adiurabit eam sacerdos iuramento maledictionis: "Det te Dominus in maledictionem, iuramentum in medio populi tui; putrescere faciat femur tuum, et tumens uterus tuus disrumpatur;
NUM|5|22|ingrediantur aquae maledictae in ventrem tuum, et utero tumescente putrescat femur!". Et respondebit mulier: "Amen, amen".
NUM|5|23|Scribetque sacerdos in libello ista maledicta et delebit ea aquis amarissimis
NUM|5|24|et dabit ei bibere aquas amaras, in quas maledicta congessit, et ingredientur in eam aquae maledictionis, quae amarae fient;
NUM|5|25|tollet sacerdos de manu eius sacrificium zelotypiae et agitabit illud coram Domino imponetque illud super altare;
NUM|5|26|pugillum sacrificii tollat de eo, quod offertur in memoriale, et incendat super altare; et deinde potum det mulieri aquas amarissimas.
NUM|5|27|Quas cum biberit, si polluta est et, contempto viro, adulterii rea, pertransibunt eam aquae maledictionis et, inflato ventre, computrescet femur; eritque mulier in maledictionem omni populo eius.
NUM|5|28|Quod si polluta non fuerit sed munda, erit innoxia et faciet liberos ".
NUM|5|29|Ista est lex zelotypiae, si declinaverit mulier a viro suo et si polluta fuerit,
NUM|5|30|maritusque zelotypiae spiritu concitatus adduxerit eam in conspectu Domini, et fecerit ei sacerdos iuxta omnia, quae scripta sunt;
NUM|5|31|maritus absque culpa erit, et illa recipiet iniquitatem suam.
NUM|6|1|Locutusque est Dominus ad Moysen dicens:
NUM|6|2|" Loquere ad filios Israel et dices ad eos: Vir sive mulier cum fecerint votum, ut sanctificentur et se voluerint Domino consecrare,
NUM|6|3|a vino et omni quod inebriare potest abstinebunt; acetum ex vino et ex qualibet alia potione et, quidquid de uva exprimitur, non bibent; uvas recentes siccasque non comedent
NUM|6|4|cunctis diebus, quibus ex voto Domino consecrantur: quidquid ex vinea esse potest ab uva acerba usque ad pellicula non comedent.
NUM|6|5|Omni tempore separationis suae novacula non transibit per caput eius usque ad completum tempus, quo Domino consecratur; sanctus erit crescente caesarie capitis eius.
NUM|6|6|Omni tempore consecrationis suae ad mortuum non ingredietur;
NUM|6|7|nec super patris quidem et matris et fratris sororisque funere contaminabitur, quia consecratio Dei sui super caput eius est.
NUM|6|8|Omnibus diebus separationis suae sanctus erit Domino.
NUM|6|9|Sin autem mortuus fuerit subito quispiam coram eo, polluetur caput consecrationis eius; quod radet ilico in eadem die purgationis suae, id est die septima.
NUM|6|10|In octava autem die offeret duos turtures vel duos pullos columbae sacerdoti in introitu tabernaculi conventus,
NUM|6|11|facietque sacerdos unum pro peccato et alterum in holocaustum et expiabit pro eo, quia peccavit super mortuo, sanctificabitque caput eius in die illo
NUM|6|12|et consecrabit Domino dies separationis suae offerens agnum anniculum pro delicto; ita tamen, ut dies priores irriti fiant, quoniam polluta est consecratio eius.
NUM|6|13|Ista est lex consecrationis, cum dies, quos ex voto decreverat, complebuntur: adducent eum ad ostium tabernaculi conventus,
NUM|6|14|et offeret oblationem suam Domino agnum anniculum immaculatum in holocaustum et ovem anniculam immaculatam pro peccato et arietem immaculatum hostiam pacificam,
NUM|6|15|canistrum quoque panum azymorum, qui permixti sint oleo, et lagana absque fermento uncta oleo ac oblationem et libamina singulorum.
NUM|6|16|Quae offeret sacerdos coram Domino et faciet tam pro peccato quam in holocaustum;
NUM|6|17|arietem vero immolabit hostiam pacificam Domino offerens simul canistrum azymorum; facietque oblationem eius et libamenta.
NUM|6|18|Tunc radet nazaraeus ante ostium tabernaculi conventus caesariem consecrationis suae tolletque capillos suos et ponet super ignem, qui est suppositus sacrificio pacificorum,
NUM|6|19|et sumet sacerdos armum coctum arietis tortamque absque fermento unam de canistro et laganum azymum unum et tradet in manus nazaraei, postquam rasum fuerit caput eius;
NUM|6|20|et agitabit in conspectu Domini, et sanctificata sacerdotis erunt sicut pectusculum, quod agitari, et femur, quod praelevari iussum est. Post haec potest bibere nazaraeus vinum ".
NUM|6|21|Ista est lex nazaraei, cum voverit oblationem suam Domino tempore consecrationis suae, exceptis his, quae invenerit manus eius. Iuxta quod devoverat, ita faciet secundum legem consecrationis suae.
NUM|6|22|Locutusque est Dominus ad Moysen dicens:
NUM|6|23|" Loquere Aaron et filiis eius: Sic benedicetis filiis Israel et dicetis eis:
NUM|6|24|"Benedicat tibi Dominus et custodiat te!
NUM|6|25|Illuminet Dominus faciem suam super te et misereatur tui!
NUM|6|26|Convertat Dominus vultum suum ad te et det tibi pacem!".
NUM|6|27|Invocabuntque nomen meum super filios Israel, et ego benedicam eis ".
NUM|7|1|Factum est autem in die, qua complevit Moyses habitaculum et erexit illud unxitque et sanctificavit cum omnibus vasis suis, altare similiter et omnia vasa eius,
NUM|7|2|obtulerunt principes Israel et capita familiarum, qui erant per singulas tribus praefecti eorum, qui numerati fuerant,
NUM|7|3|munera coram Domino sex plaustra tecta cum duodecim bobus. Unum plaustrum obtulere duo duces et unum bovem singuli; obtuleruntque ea in conspectu habitaculi.
NUM|7|4|Ait autem Dominus ad Moysen:
NUM|7|5|" Suscipe ab eis, ut serviant in ministerio tabernaculi conventus, et trades ea Levitis iuxta ordinem ministerii sui ".
NUM|7|6|Itaque cum suscepisset Moyses plaustra et boves, tradidit eos Levitis.
NUM|7|7|Duo plaustra et quattuor boves dedit filiis Gerson, iuxta id quod habebant necessarium.
NUM|7|8|Quattuor alia plaustra et octo boves dedit filiis Merari, secundum offficia sua sub manu Ithamar filii Aaron sacerdotis.
NUM|7|9|Filiis autem Caath non dedit plaustra et boves, quia in sanctuario serviunt et onera propriis portant umeris.
NUM|7|10|Igitur obtulerunt duces in dedicationem altaris die, qua unctum est, oblationem suam ante altare.
NUM|7|11|Dixitque Dominus ad Moysen: " Singuli duces per singulos dies offerant munera in dedicationem altaris ".
NUM|7|12|Primo die obtulit oblationem suam Naasson filius Aminadab de tribu Iudae.
NUM|7|13|Fueruntque in ea scutula argentea pondo centum triginta siclorum, phiala argentea habens septuaginta siclos iuxta pondus sanctuarii, utraque plena simila conspersa oleo in sacrificium,
NUM|7|14|acetabulum ex decem siclis aureis plenum incenso,
NUM|7|15|bos de armento et aries et agnus anniculus in holocaustum
NUM|7|16|hircusque pro peccato;
NUM|7|17|et in sacrificio pacificorum boves duo, arietes quinque, hirci quinque, agni anniculi quinque: haec est oblatio Naasson filii Aminadab.
NUM|7|18|Secundo die obtulit Nathanael filius Suar dux de tribu Issachar
NUM|7|19|scutulam argenteam appendentem centum triginta siclos, phialam argenteam habentem septuaginta siclos iuxta pondus sanctuarii, utramque plenam simila conspersa oleo in sacrificium,
NUM|7|20|acetabulum aureum habens decem siclos plenum incenso,
NUM|7|21|bovem de armento et arietem et agnum anniculum in holocaustum
NUM|7|22|hircumque pro peccato;
NUM|7|23|et in sacrificio pacificorum boves duos, arietes quinque, hircos quinque, agnos anniculos quinque: haec fuit oblatio Nathanael filii Suar.
NUM|7|24|Tertio die princeps filiorum Zabulon Eliab filius Helon
NUM|7|25|obtulit scutulam argenteam appendentem centum triginta siclos, phialam argenteam habentem septuaginta siclos ad pondus sanctuarii, utramque plenam simila conspersa oleo in sacrificium,
NUM|7|26|acetabulum aureum appendens decem siclos plenum incenso,
NUM|7|27|bovem de armento et arietem et agnum anniculum in holocaustum
NUM|7|28|hircumque pro peccato;
NUM|7|29|et in sacrificio pacificorum boves duos, arietes quinque, hircos quinque, agnos anniculos quinque: haec est oblatio Eliab filii Helon.
NUM|7|30|Die quarto princeps filiorum Ruben Elisur filius Sedeur
NUM|7|31|obtulit scutulam argenteam appendentem centum triginta siclos, phialam argenteam habentem septuaginta siclos ad pondus sanctuarii, utramque plenam simila conspersa oleo in sacrificium,
NUM|7|32|acetabulum aureum appendens decem siclos plenum incenso,
NUM|7|33|bovem de armento et arietem et agnum anniculum in holocaustum
NUM|7|34|hircumque pro peccato;
NUM|7|35|et in hostias pacificorum boves duos, arietes quinque, hircos quinque, agnos anniculos quinque: haec fuit oblatio Elisur filii Sedeur.
NUM|7|36|Die quinto princeps filiorum Simeon Salamiel filius Surisaddai
NUM|7|37|obtulit scutulam argenteam appendentem centum triginta siclos, phialam argenteam habentem septuaginta siclos ad pondus sanctuarii, utramque plenam simila conspersa oleo in sacrificium,
NUM|7|38|acetabulum aureum appendens decem siclos plenum incenso,
NUM|7|39|bovem de armento et arietem et agnum anniculum in holocaustum,
NUM|7|40|hircumque pro peccato;
NUM|7|41|et in hostias pacificorum boves duos, arietes quinque, hircos quinque, agnos anniculos quinque: haec fuit oblatio Salamiel filii Surisaddai.
NUM|7|42|Die sexto princeps filiorum Gad Eliasaph filius Deuel
NUM|7|43|obtulit scutulam argenteam appendentem centum triginta siclos, phialam argenteam habentem septuaginta siclos ad pondus sanctuarii, utramque plenam simila conspersa oleo in sacrificium,
NUM|7|44|acetabulum aureum appendens decem siclos plenum incenso,
NUM|7|45|bovem de armento et arietem et agnum anniculum in holocaustum,
NUM|7|46|hircumque pro peccato;
NUM|7|47|et in hostias pacificorum boves duos, arietes quinque, hircos quinque, agnos anniculos quinque: haec fuit oblatio Eliasaph filii Deuel.
NUM|7|48|Die septimo princeps filiorum Ephraim Elisama filius Ammiud
NUM|7|49|obtulit scutulam argenteam appendentem centum triginta siclos, phialam argenteam habentem septuaginta siclos ad pondus sanctuarii, utramque plenam simila conspersa oleo in sacrificium,
NUM|7|50|acetabulum aureum appendens decem siclos plenum incenso,
NUM|7|51|bovem de armento et arietem et agnum anniculum in holocaustum,
NUM|7|52|hircumque pro peccato;
NUM|7|53|et in hostias pacificorum boves duos, arietes quinque, hircos quinque, agnos anniculos quinque: haec fuit oblatio Elisama filii Ammiud.
NUM|7|54|Die octavo princeps filiorum Manasse Gamaliel filius Phadassur
NUM|7|55|obtulit scutulam argenteam appendentem centum triginta siclos, phialam argenteam habentem septuaginta siclos ad pondus sanctuarii, utramque plenam simila conspersa oleo in sacrificium,
NUM|7|56|acetabulum aureum appendens decem siclos plenum incenso,
NUM|7|57|bovem de armento et arietem et agnum anniculum in holocaustum
NUM|7|58|hircumque pro peccato;
NUM|7|59|et in hostias pacificorum boves duos, arietes quinque, hircos quinque, agnos anniculos quinque: haec fuit oblatio Gamaliel filii Phadassur.
NUM|7|60|Die nono princeps filiorum Beniamin Abidan filius Gedeonis
NUM|7|61|obtulit scutulam argenteam appendentem centum triginta siclos, phialam argenteam habentem septuaginta siclos ad pondus sanctuarii, utramque plenam simila conspersa oleo in sacrificium,
NUM|7|62|et acetabulum aureum appendens decem siclos plenum incenso,
NUM|7|63|bovem de armento et arietem et agnum anniculum in holocaustum
NUM|7|64|hircumque pro peccato;
NUM|7|65|et in hostias pacificorum boves duos, arietes quinque, hircos quinque, agnos anniculos quinque: haec fuit oblatio Abidan filii Gedeonis.
NUM|7|66|Die decimo princeps filiorum Dan Ahiezer filius Ammisaddai
NUM|7|67|obtulit scutulam argenteam appendentem centum triginta siclos, phialam argenteam habentem septuaginta siclos ad pondus sanctuarii, utramque plenam simila conspersa oleo in sacrificium,
NUM|7|68|acetabulum aureum appendens decem siclos plenum incenso,
NUM|7|69|bovem de armento et arietem et agnum anniculum in holocaustum
NUM|7|70|hircumque pro peccato;
NUM|7|71|et in hostias pacificorum boves duos, arietes quinque, hircos quinque, agnos anniculos quinque: haec fuit oblatio Ahiezer filii Ammisaddai.
NUM|7|72|Die undecimo princeps filiorum Aser Phegiel filius Ochran
NUM|7|73|obtulit scutulam argenteam appendentem centum triginta siclos, phialam argenteam habentem septuaginta siclos ad pondus sanctuarii, utramque plenam simila conspersa oleo in sacrificium,
NUM|7|74|acetabulum aureum appendens decem siclos plenum incenso,
NUM|7|75|bovem de armento et arietem et agnum anniculum in holocaustum
NUM|7|76|hircumque pro peccato;
NUM|7|77|et in hostias pacificorum boves duos, arietes quinque, hircos quinque, agnos anniculos quinque: haec fuit oblatio Phegiel filii Ochran.
NUM|7|78|Die duodecimo princeps filiorum Nephthali Ahira filius Enan
NUM|7|79|obtulit scutulam argenteam appendentem centum triginta siclos, phialam argenteam habentem septuaginta siclos ad pondus sanctuarii, utramque plenam simila oleo conspersa in sacrificium,
NUM|7|80|acetabulum aureum appendens decem siclos plenum incenso,
NUM|7|81|bovem de armento et arietem et agnum anniculum in holocaustum
NUM|7|82|hircumque pro peccato;
NUM|7|83|et in hostias pacificorum boves duos, arietes quinque, hircos quinque, agnos anniculos quinque: haec fuit oblatio Ahira filii Enan.
NUM|7|84|Haec in dedicatione altaris oblata sunt a principibus Israel in die, qua consecratum est: scutulae argenteae duodecim, phialae argenteae duodecim, acetabula duodecim,
NUM|7|85|ita ut centum triginta siclos argenti haberet una scutella, et septuaginta siclos haberet una phiala, id est in commune vasorum omnium ex argento sicli duo milia quadringenti pondere sanctuarii;
NUM|7|86|acetabula aurea duodecim plena incenso denos siclos appendentia pondere sanctuarii, id est simul auri sicli centum viginti;
NUM|7|87|omnes boves de armento in holocaustum duodecim, arietes duodecim, agni anniculi duodecim et libamenta eorum; hirci duodecim pro peccato.
NUM|7|88|In hostias pacificorum omnes boves viginti quattuor, arietes sexaginta, hirci sexaginta, agni anniculi sexaginta: haec oblata sunt in dedicatione altaris, quando unctum est.
NUM|7|89|Cumque ingrederetur Moyses tabernaculum testimonii, ut consuleret oraculum, audiebat vocem loquentis ad se de propitiatorio, quod erat super arcam testimonii inter duos cherubim, unde et loquebatur ei.
NUM|8|1|Locutusque est Dominus ad Moysen dicens:
NUM|8|2|" Loquere Aa ron et dices ad eum: Cum posueris lucernas, contra eam partem, quam candelabrum respicit, lucere debebunt septem lucernae ".
NUM|8|3|Fecitque sic Aaron et posuit lucernas super candelabrum, ut praeceperat Dominus Moysi.
NUM|8|4|Haec autem erat factura candelabri: ex auro ductili, tam medius stipes quam flores eius. Iuxta exemplum, quod ostendit Dominus Moysi, ita operatus est candelabrum.
NUM|8|5|Et locutus est Dominus ad Moysen dicens:
NUM|8|6|" Tolle Levitas de medio filiorum Israel et purificabis eos
NUM|8|7|iuxta hunc ritum. Aspergantur aqua lustrationis et radant omnes pilos carnis suae, lavabunt vestimenta sua et mundabunt se.
NUM|8|8|Tollent bovem de armentis et oblationem eius similam oleo conspersam; bovem autem alterum de armento tu accipies pro peccato
NUM|8|9|et applicabis Levitas coram tabernaculo conventus, convocata omni multitudine filiorum Israel.
NUM|8|10|Cumque Levitae fuerint coram Domino, ponent filii Israel manus suas super eos,
NUM|8|11|et agitabit Aaron Levitas munus in conspectu Domini a filiis Israel, ut serviant in ministerio eius.
NUM|8|12|Levitae quoque ponent manus suas super capita boum, e quibus unum facies pro peccato et alterum in holocaustum Domini, ut expies eos.
NUM|8|13|Statuesque Levitas in conspectu Aaron et filiorum eius et agitabis eos Domino
NUM|8|14|ac separabis de medio filiorum Israel, ut sint mei;
NUM|8|15|et postea ingredientur, ut serviant tabernaculo conventus.Sicque purificabis et agitabis eos,
NUM|8|16|quoniam dono donati sunt mihi e medio filiorum Israel; pro primogenitis, quae aperiunt omnem vulvam in Israel, accepi eos.
NUM|8|17|Mea sunt enim omnia primogenita filiorum Israel, tam ex hominibus quam ex iumentis. Ex die, quo percussi omne primogenitum in terra Aegypti, sanctificavi eos mihi.
NUM|8|18|Et tuli Levitas pro cunctis primogenitis filiorum Israel
NUM|8|19|tradidique eos dono Aaron et filiis eius de medio filiorum Israel, ut serviant mihi pro Israel in tabernaculo conventus et expient pro eis, ne sit in populo plaga, si ausi fuerint accedere ad sanctuarium ".
NUM|8|20|Feceruntque Moyses et Aaron et omnis congregatio filiorum Israel super Levitis, quae praeceperat Dominus Moysi.
NUM|8|21|Purificatique sunt et laverunt vestimenta sua, agitavitque eos Aaron in conspectu Domini et expiavit eos, ut purificati
NUM|8|22|ingrederentur ad officia sua in tabernaculo conventus coram Aaron et filiis eius; sicut praeceperat Dominus Moysi de Levitis, ita factum est.
NUM|8|23|Locutusque est Dominus ad Moysen dicens:
NUM|8|24|" Haec est lex Levitarum: a viginti quinque annis et supra ingredientur, ut ministrent in tabernaculo conventus;
NUM|8|25|cumque quinquagesimum annum aetatis impleverint, servire cessabunt
NUM|8|26|eruntque ministri fratrum suorum in tabernaculo conventus, ut custodiant, quae sibi fuerint commendata; opera autem ipsa non faciant. Sic dispones Levitis in custodiis suis ".
NUM|9|1|Locutus est Dominus ad Moy sen in deserto Sinai anno secun do, postquam egressi sunt de terra Aegypti, mense primo dicens:
NUM|9|2|" Faciant filii Israel Pascha in tempore suo
NUM|9|3|quarta decima die mensis huius ad vesperam iuxta omnia praecepta et iustificationes eius ".
NUM|9|4|Praecepitque Moyses filiis Israel, ut facerent Pascha.
NUM|9|5|Qui fecerunt tempore suo quarta decima die mensis ad vesperam in deserto Sinai; iuxta omnia, quae mandaverat Dominus Moysi, fecerunt filii Israel.
NUM|9|6|Ecce autem quidam immundi super animam hominis, qui non poterant facere Pascha in die illo, accedentes ad Moysen et Aaron
NUM|9|7|dixerunt ei: " Immundi sumus super animam hominis; quare fraudamur, ut non valeamus oblationem offerre Domino in tempore suo inter filios Israel? ".
NUM|9|8|Quibus respondit Moyses: " State, ut consulam quid praecipiat Dominus de vobis ".
NUM|9|9|Locutusque est Dominus ad Moysen dicens:
NUM|9|10|" Loquere filiis Israel: Homo, qui fuerit immundus super anima, sive in via procul in gente vestra, faciat Pascha Domino
NUM|9|11|in mense secundo quarta decima die mensis ad vesperam; cum azymis et lactucis agrestibus comedent illud,
NUM|9|12|non relinquent ex eo quippiam usque mane et os eius non confringent: omnem ritum Pascha observabunt.
NUM|9|13|Si quis autem et mundus est et in itinere non fuit et tamen non fecit Pascha, exterminabitur anima illa de populis suis, quia sacrificium Domino non obtulit tempore suo: peccatum suum ipse portabit.
NUM|9|14|Peregrinus quoque et advena, si fuerint apud vos, facient Pascha Domino iuxta praecepta et iustificationes eius; praeceptum idem erit apud vos tam advenae quam indigenae ".
NUM|9|15|Igitur die, qua erectum est habitaculum, operuit nubes habitaculum, tabernaculum testimonii; a vespere autem super habitaculum erat quasi species ignis usque mane.
NUM|9|16|Sic fiebat iugiter: per diem operiebat illud nubes, et per noctem quasi species ignis.
NUM|9|17|Cumque ablata fuisset nubes, quae tabernaculum protegebat, tunc proficiscebantur filii Israel; et in loco, ubi stetisset nubes, ibi castrametabantur.
NUM|9|18|Ad imperium Domini proficiscebantur et ad imperium illius castrametabantur. Cunctis diebus, quibus stabat nubes super habitaculum, manebant in eodem loco.
NUM|9|19|Et si evenisset ut multo tempore maneret super illud, erant filii Israel in excubiis Domini et non proficiscebantur;
NUM|9|20|si diebus paucis fuisset nubes super habitaculum, ad imperium Domini erigebant tentoria et ad imperium illius deponebant.
NUM|9|21|Si fuisset nubes a vespere usque mane et statim diluculo habitaculum reliquisset, proficiscebantur; et si post diem et noctem recessisset, dissipabant tentoria.
NUM|9|22|Si vero biduo aut uno mense vel longiore tempore fuisset super habitaculum, manebant filii Israel in eodem loco et non proficiscebantur. Statim autem ut recessisset, movebant castra.
NUM|9|23|Per verbum Domini figebant tentoria et per verbum illius proficiscebantur; erantque in excubiis Domini iuxta imperium eius per manum Moysi.
NUM|10|1|Locutusque est Dominus ad Moysen dicens:
NUM|10|2|" Fac tibi duas tubas argenteas ductiles, quibus convocare possis congregationem, quando movenda sunt castra.
NUM|10|3|Cumque increpueris tubis, congregabitur ad te omnis turba ad ostium tabernaculi conventus.
NUM|10|4|Si semel clangueris, venient ad te principes et capita congregationis Israel;
NUM|10|5|si autem prolixior clangor increpuerit, movebunt castra primi, qui sunt ad orientalem plagam;
NUM|10|6|in secundo autem sonitu et pari ululatu tubae levabunt tentoria, qui habitant ad meridiem, et iuxta hunc modum reliqui facient, ululantibus tubis in profectionem.
NUM|10|7|Quando autem congregandus est populus, simplex tubarum clangor erit, et non ululabunt.
NUM|10|8|Filii autem Aaron sacerdotes clangent tubis. Eritque hoc vobis legitimum sempiternum in generationibus vestris.
NUM|10|9|Si exieritis ad bellum in terra vestra contra hostes, qui dimicant adversum vos, clangetis ululantibus tubis; et erit recordatio vestri coram Domino Deo vestro, ut eruamini de manibus inimicorum vestrorum.
NUM|10|10|Si quando habebitis epulum et dies festos et calendas, canetis tubis super holocaustis vestris et pacificis victimis, ut sint vobis in recordationem Dei vestri. Ego Dominus Deus vester ".
NUM|10|11|Anno secundo, mense secundo, vicesima die mensis elevata est nubes de habitaculo testimonii;
NUM|10|12|profectique sunt filii Israel per migrationes suas de deserto Sinai, et recubuit nubes in solitudine Pharan.
NUM|10|13|Moveruntque castra prima vice, iuxta imperium Domini in manu Moysi.
NUM|10|14|Elevatum est primum vexillum castrorum filiorum Iudae per turmas suas, quorum princeps erat Naasson filius Aminadab;
NUM|10|15|et super turmam tribus filiorum Issachar fuit princeps Nathanael filius Suar;
NUM|10|16|et super turmam tribus Zabulon erat princeps Eliab filius Helon.
NUM|10|17|Depositumque est habitaculum, quod portantes egressi sunt filii Gerson et Merari.
NUM|10|18|Profectum est vexillum castrorum filiorum Ruben per turmas suas, et super turbam suam princeps erat Elisur filius Sedeur.
NUM|10|19|Super turmam autem tribus filiorum Simeon princeps fuit Salamiel filius Surisaddai.
NUM|10|20|Porro super turmam tribus filiorum Gad erat princeps Eliasaph filius Deuel.
NUM|10|21|Profectique sunt et Caathitae portantes sanctuarium. Et erectum est habitaculum, antequam venirent.
NUM|10|22|Elevatum est vexillum castrorum filiorum Ephraim per turmas suas, in quorum exercitu princeps erat Elisama filius Ammiud.
NUM|10|23|Et super turmam tribus filiorum Manasse princeps fuit Gamaliel filius Phadassur;
NUM|10|24|et super turmam tribus filiorum Beniamin erat dux Abidan filius Gedeonis.
NUM|10|25|Novissime elevatum est vexillum castrorum filiorum Dan per turmas suas, in quorum exercitu princeps fuit Ahiezer filius Ammisaddai.
NUM|10|26|Et super turmam tribus filiorum Aser erat princeps Phegiel filius Ochran;
NUM|10|27|et super turmam tribus filiorum Nephthali princeps fuit Ahira filius Enan.
NUM|10|28|Hae sunt profectiones filiorum Israel per turmas suas, quando egrediebantur.
NUM|10|29|Dixitque Moyses Hobab filio Raguel Madianitae cognato suo: " Proficiscimur ad locum, quem Dominus daturus est nobis; veni nobiscum, ut benefaciamus tibi, quia Dominus bona promisit Israeli ".
NUM|10|30|Cui ille respondit: " Non vadam tecum, sed revertar in terram meam, in qua natus sum ".
NUM|10|31|Et ille: " Noli, inquit, nos relinquere; tu enim nosti in quibus locis per desertum castra ponere debeamus, et eris ductor noster.
NUM|10|32|Cumque nobiscum veneris, quidquid optimum fuerit ex opibus, quas nobis traditurus est Dominus, dabimus tibi ".
NUM|10|33|Profecti sunt ergo de monte Domini viam trium dierum; arcaque foederis Domini praecedebat eos per dies tres providens castrorum locum.
NUM|10|34|Nubes quoque Domini super eos erat per diem, cum incederent.
NUM|10|35|Cumque elevaretur arca, dicebat Moyses: " Surge, Domine, et dissipentur inimici tui; et fugiant, qui oderunt te, a facie tua ".
NUM|10|36|Cum autem deponeretur, aiebat: " Revertere, Domine, ad multitudinem exercitus Israel ".
NUM|11|1|Ortum est murmur populi, quasi dolentium pro labore, contra Dominum. Quod cum audisset Dominus, iratus est, et accensus in eos ignis Domini devoravit extremam castrorum partem.
NUM|11|2|Cumque clamasset populus ad Moysen, oravit Moyses ad Dominum, et absorptus est ignis.
NUM|11|3|Vocaverunt nomen loci illius Tabera, eo quod incensus fuisset contra eos ignis Domini.
NUM|11|4|Vulgus autem promiscuum, quod erat in medio eius, flagravit desiderio, et sedentes fleverunt pariter filii Israel et dixerunt: " Quis dabit nobis ad vescendum carnes?
NUM|11|5|Recordamur piscium, quos comedebamus in Aegypto gratis; in mentem nobis veniunt cucumeres et pepones porrique et cepae et alia.
NUM|11|6|Guttur nostrum aridum est; nihil aliud respiciunt oculi nostri nisi man ".
NUM|11|7|Erat autem man quasi semen coriandri aspectus bdellii.
NUM|11|8|Circuibatque populus et colligens illud frangebat mola sive terebat in mortario coquens in olla et faciens ex eo tortulas saporis quasi panis oleati.
NUM|11|9|Cumque descenderet nocte super castra ros, descendebat pariter et man.
NUM|11|10|Audivit ergo Moyses flentem populum per familias, singulos per ostia tentorii sui. Iratusque est furor Domini valde; quod Moysi intoleranda res visa est,
NUM|11|11|et ait ad Dominum: " Cur afflixisti servum tuum? Quare non invenio gratiam coram te? Et cur imposuisti pondus universi populi huius super me?
NUM|11|12|Numquid ego concepi omnem hunc populum vel genui eum, ut dicas mihi: "Porta eum in sinu tuo, sicut portare solet nutrix infantulum, et defer in terram, pro qua iurasti patribus eorum?".
NUM|11|13|Unde mihi carnes, ut dem universo populo isti? Flent contra me dicentes: "Da nobis carnes, ut comedamus!".
NUM|11|14|Non possum ego solus sustinere omnem hunc populum, quia nimis gravis est mihi.
NUM|11|15|Si hoc modo agis mecum, obsecro ut interficias me, si inveni gratiam in oculis tuis, ne videam amplius mala mea! ".
NUM|11|16|Et dixit Dominus ad Moysen: " Congrega mihi septuaginta viros de senibus Israel, quos tu nosti quod senes populi sint ac magistri, et duces eos ad ostium tabernaculi conventus, stabuntque ibi tecum.
NUM|11|17|Et descendam et loquar tibi et auferam de spiritu tuo tradamque eis, ut sustentent tecum onus populi, et non tu solus graveris.
NUM|11|18|Populo quoque dices: Sanctificamini, cras comedetis carnes; ego enim audivi vos flere: "Quis dabit nobis escas carnium? Bene nobis erat in Aegypto". Et dabit vobis Dominus carnes, et comedetis
NUM|11|19|non uno die nec duobus vel quinque aut decem nec viginti quidem,
NUM|11|20|sed usque ad mensem dierum, donec exeat per nares vestras et vertatur in nauseam, eo quod reppuleritis Dominum, qui in medio vestri est, et fleveritis coram eo dicentes: "Quare egressi sumus ex Aegypto?" ".
NUM|11|21|Et ait Moyses: " Populus, in cuius medio sum, sescenta milia peditum sunt, et tu dicis: "Dabo eis esum carnium mense integro!".
NUM|11|22|Numquid ovium et boum multitudo caedetur, ut possit sufficere ad cibum? Vel omnes pisces maris in unum congregabuntur, ut eos satient? ".
NUM|11|23|Cui respondit Dominus: " Numquid manus Domini abbreviata est? Iam nunc videbis utrum meus sermo opere compleatur an non ".
NUM|11|24|Venit igitur Moyses et narravit populo verba Domini congregans septuaginta viros de senibus Israel, quos stare fecit circa tabernaculum.
NUM|11|25|Descenditque Dominus per nubem et locutus est ad eum auferens de spiritu, qui erat in Moyse, et dans septuaginta viris senibus. Cumque requievisset in eis spiritus, prophetaverunt nec ultra fecerunt.
NUM|11|26|Remanserant autem in castris duo viri, quorum unus vocabatur Eldad et alter Medad, super quos requievit spiritus; nam et ipsi descripti fuerant et non exierant ad tabernaculum. Cumque prophetarent in castris,
NUM|11|27|cucurrit puer et nuntiavit Moysi dicens: " Eldad et Medad prophetant in castris ".
NUM|11|28|Statim Iosue filius Nun minister Moysi et electus eius a iuventute sua ait: " Domine mi Moyses, prohibe eos! ".
NUM|11|29|At ille: " Quid, inquit, aemularis pro me? Quis tribuat, ut omnis populus prophetet, et det eis Dominus spiritum suum? ".
NUM|11|30|Reversusque est Moyses et maiores natu Israel in castra.
NUM|11|31|Ventus autem egrediens a Domino arreptas trans mare coturnices detulit et demisit in castra itinere, quantum uno die confici potest, ex omni parte castrorum per circuitum; volabantque in aere duobus cubitis altitudine super terram.
NUM|11|32|Surgens ergo populus toto die illo et nocte ac die altero congregavit coturnicum, qui parum, decem choros; et extenderunt eas per gyrum castrorum.
NUM|11|33|Adhuc carnes erant in dentibus eorum, nec defecerat huiuscemodi cibus, et ecce furor Domini concitatus in populum percussit eum plaga magna nimis.
NUM|11|34|Vocatusque est ille locus Cibrottaava; ibi enim sepelierunt populum, qui desideraverat.
NUM|11|35|Egressi autem de Cibrottaava, venerunt in Aseroth et manserunt ibi.
NUM|12|1|Locutaque est Maria et Aaron contra Moysen propter uxorem eius Aethiopissam
NUM|12|2|et dixerunt: " Num per solum Moysen locutus est Dominus? Nonne et per nos similiter est locutus? ". Quod cum audisset Dominus
NUM|12|3|­ erat enim Moyses vir humillimus super omnes homines, qui morabantur in terra ­
NUM|12|4|statim locutus est ad eum et ad Aaron et Mariam: " Egredimini vos tantum tres ad tabernaculum conventus ". Cumque fuissent egressi,
NUM|12|5|descendit Dominus in columna nubis et stetit in introitu tabernaculi vocans Aaron et Mariam. Qui cum issent,
NUM|12|6|dixit ad eos:" Audite sermones meos!Si quis fuerit inter vos propheta Domini,in visione apparebo eivel per somnium loquar ad illum.
NUM|12|7|At non talis servus meus Moyses,qui in omni domo mea fidelissimus est!
NUM|12|8|Ore enim ad os loquor ei,et palam et non per aenigmata et figurasDominum videt!Quare ergo non timuistis detrahereservo meo Moysi? ".
NUM|12|9|Iratusque contra eos abiit,
NUM|12|10|nubes quoque recessit, quae erat super tabernaculum; et ecce Maria apparuit candens lepra quasi nix.Cumque respexisset eam Aaron et vidisset perfusam lepra,
NUM|12|11|ait ad Moysen: " Obsecro, domine mi, ne imponas nobis hoc peccatum, quod stulte commisimus,
NUM|12|12|ne fiat haec quasi mortua et ut abortivum, quod proicitur de vulva matris suae; ecce iam medium carnis eius devoratum est a lepra ".
NUM|12|13|Clamavitque Moyses ad Dominum dicens: " Deus, obsecro, sana eam! ".
NUM|12|14|Cui respondit Dominus: " Si pater eius spuisset in faciem illius, nonne debuerat saltem septem diebus rubore suffundi? Separetur septem diebus extra castra et postea revocabitur ".
NUM|12|15|Exclusa est itaque Maria extra castra septem diebus, et populus non est motus de loco illo, donec revocata est Maria.
NUM|12|16|Profectusque est populus de Aseroth, fixis tentoriis in deserto Pharan.
NUM|13|1|Ibi locutus est Dominus ad Moysen dicens:
NUM|13|2|" Mitte vi ros, qui considerent terram Chanaan, quam daturus sum filiis Israel, singulos de singulis tribubus ex principibus ".
NUM|13|3|Fecit Moyses quod Dominus imperaverat, de deserto Pharan mittens principes viros, quorum ista sunt nomina:
NUM|13|4|de tribu Ruben Sammua filium Zacchur,
NUM|13|5|de tribu Simeon Saphat filium Hori,
NUM|13|6|de tribu Iudae Chaleb filium Iephonne,
NUM|13|7|de tribu Issachar Igal filium Ioseph,
NUM|13|8|de tribu Ephraim Osee filium Nun,
NUM|13|9|de tribu Beniamin Phalti filium Raphu,
NUM|13|10|de tribu Zabulon Geddiel filium Sodi,
NUM|13|11|de tribu Ioseph, tribu Manasse, Gaddi filium Susi,
NUM|13|12|de tribu Dan Ammiel filium Gemalli,
NUM|13|13|de tribu Aser Sthur filium Michael,
NUM|13|14|de tribu Nephthali Nahabi filium Vaphsi,
NUM|13|15|de tribu Gad Guel filium Machi.
NUM|13|16|Haec sunt nomina virorum, quos misit Moyses ad considerandam terram. Vocavitque Osee filium Nun Iosue.
NUM|13|17|Misit ergo eos Moyses ad considerandam terram Chanaan et dixit ad eos: " Ascendite per Nageb. Cumque veneritis ad montes,
NUM|13|18|considerate terram, qualis sit, et populum, qui habitator est eius, utrum fortis sit an infirmus, si pauci numero an plures;
NUM|13|19|ipsa terra bona an mala, urbes quales, absque muris an muratae;
NUM|13|20|humus pinguis an sterilis, nemorosa an absque arboribus. Confortamini et afferte nobis de fructibus terrae ". Erat autem tempus, quando iam praecoquae uvae vesci possunt.
NUM|13|21|Cumque ascendissent, exploraverunt terram a deserto Sin usque Rohob in introitu Emath.
NUM|13|22|Ascenderuntque ad Nageb et venerunt in Hebron, ubi erant Ahiman et Sesai et Tholmai filii Enac. Nam Hebron septem annis ante Tanim urbem Aegypti condita est.
NUM|13|23|Pergentesque usque ad Nehelescol absciderunt palmitem cum uva sua, quem portaverunt in vecte duo viri. De malis quoque granatis et de ficis loci illius tulerunt,
NUM|13|24|qui appellatus est Nehelescol, eo quod botrum portassent inde filii Israel.
NUM|13|25|Reversique exploratores terrae post quadraginta dies, omni regione circuita,
NUM|13|26|venerunt ad Moysen et Aaron et ad omnem coetum filiorum Israel in desertum Pharan, quod est in Cades. Locutique eis et omni congregationi ostenderunt fructus terrae
NUM|13|27|et narraverunt dicentes: " Venimus in terram, ad quam misisti nos, quae re vera fluit lacte et melle, ut ex his fructibus cognosci potest.
NUM|13|28|Sed cultores fortissimos habet et urbes grandes atque muratas. Stirpem Enac vidimus ibi;
NUM|13|29|Amalec habitat in Nageb, Hetthaeus et Iebusaeus et Amorraeus in montanis, Chananaeus vero moratur iuxta mare et circa fluenta Iordanis ".
NUM|13|30|Inter haec Chaleb compescens murmur populi, qui oriebatur contra Moysen, ait: " Ascendamus et possideamus terram, quoniam poterimus obtinere eam ".
NUM|13|31|Alii vero, qui fuerant cum eo, dicebant: " Nequaquam ad hunc populum valemus ascendere, quia fortior nobis est ".
NUM|13|32|Detraxeruntque terrae, quam inspexerant, apud filios Israel dicentes: " Terra, quam lustravimus, devorat habitatores suos; populus, quem aspeximus, procerae staturae est;
NUM|13|33|ibi vidimus gigantes, filios Enac de genere giganteo, quibus comparati quasi locustae videbamur ".
NUM|14|1|Igitur vociferans omnis tur ba flevit nocte illa,
NUM|14|2|et mur murati sunt contra Moysen et Aaron cuncti filii Israel dicentes: " Utinam mortui essemus in Aegypto vel in hac vasta solitudine!
NUM|14|3|Cur inducit nos Dominus in terram istam, ut cadamus gladio, et uxores ac liberi nostri ducantur captivi? Nonne melius est reverti in Aegyptum? ".
NUM|14|4|Dixeruntque alter ad alterum: " Constituamus nobis ducem et revertamur in Aegyptum! ".
NUM|14|5|Quo audito, Moyses et Aaron ceciderunt proni in terram coram omni congregatione filiorum Israel.
NUM|14|6|At vero Iosue filius Nun et Chaleb filius Iephonne, qui et ipsi lustraverant terram, sciderunt vestimenta sua
NUM|14|7|et ad omnem congregationem filiorum Israel locuti sunt: " Terra, quam circuivimus, valde bona est.
NUM|14|8|Si propitius fuerit Dominus, inducet nos in eam et tradet humum lacte et melle manantem.
NUM|14|9|Nolite rebelles esse contra Dominum neque timeatis populum terrae huius, quia sicut panem ita eos possumus devorare. Recessit ab eis omne praesidium; Dominus nobiscum est, nolite metuere ".
NUM|14|10|Cumque clamaret omnis congregatio et lapidibus eos vellet opprimere, apparuit gloria Domini super tabernaculum conventus cunctis filiis Israel,
NUM|14|11|et dixit Dominus ad Moysen: " Usquequo detrahet mihi populus iste? Quousque non credent mihi in omnibus signis, quae feci coram eis?
NUM|14|12|Feriam igitur eos pestilentia atque consumam; te autem faciam in gentem magnam et fortiorem quam haec est ".
NUM|14|13|Et ait Moyses ad Dominum:? Audient Aegyptii, de quorum medio eduxisti populum istum in virtute tua,
NUM|14|14|et dicent ad habitatores terrae huius, quia audierunt quod tu, Domine, in populo isto sis et facie videaris ad faciem, et nubes tua protegat illos, et in columna nubis praecedas eos per diem et in columna ignis per noctem.
NUM|14|15|Et occidisti hunc populum quasi unum hominem, et dicent gentes, quae audierunt auditum tuum:
NUM|14|16|"Non poterat Dominus introducere populum in terram, pro qua iuraverat, idcirco occidit eos in solitudine!".
NUM|14|17|Magnificetur ergo fortitudo Domini, sicut iurasti dicens:
NUM|14|18|"Dominus patiens et multae misericordiae, auferens iniquitatem et scelera nullumque innoxium derelinquens, qui visitas peccata patrum in filios in tertiam et quartam generationem".
NUM|14|19|Dimitte obsecro peccatum populi huius secundum magnitudinem misericordiae tuae, sicut propitius fuisti populo huic de Aegypto usque ad locum istum ".
NUM|14|20|Dixitque Dominus: " Dimisi iuxta verbum tuum.
NUM|14|21|Vivo ego, et implebit gloria Domini universam terram!
NUM|14|22|Attamen omnes homines, qui viderunt maiestatem meam et signa, quae feci in Aegypto et in solitudine, et tentaverunt me iam per decem vices nec oboedierunt voci meae,
NUM|14|23|non videbunt terram, pro qua iuravi patribus eorum; nec quisquam ex illis, qui detraxit mihi, intuebitur eam.
NUM|14|24|Servum meum Chaleb, qui plenus alio spiritu secutus est me, inducam in terram hanc, quam circuivit, et semen eius possidebit eam.
NUM|14|25|Quoniam Amalecites et Chananaeus habitant in vallibus, cras movete castra et revertimini in solitudinem per viam maris Rubri ".
NUM|14|26|Locutusque est Dominus ad Moysen et Aaron dicens:
NUM|14|27|" Usquequo congregatio haec pessima murmurat contra me? Querelas filiorum Israel audivi.
NUM|14|28|Dic ergo eis: Vivo ego, ait Dominus, sicut locuti estis, audiente me, sic faciam vobis!
NUM|14|29|In solitudine hac iacebunt cadavera vestra. Omnes, qui numerati estis a viginti annis et supra et murmurastis contra me,
NUM|14|30|non intrabitis terram, super quam levavi manum meam, ut habitare vos facerem, praeter Chaleb filium Iephonne et Iosue filium Nun.
NUM|14|31|Parvulos autem vestros, de quibus dixistis quod praedae hostibus forent, introducam, ut videant terram, quae vobis displicuit.
NUM|14|32|Vestra cadavera iacebunt in solitudine hac;
NUM|14|33|filii vestri erunt pastores in deserto annis quadraginta et portabunt fornicationem vestram, donec consumantur cadavera vestra in deserto.
NUM|14|34|Iuxta numerum quadraginta dierum, quibus considerastis terram ­ annus pro die imputabitur ­ quadraginta annis portabitis iniquitates vestras et scietis ultionem meam.
NUM|14|35|Ego Dominus locutus sum, ita faciam omni congregationi huic pessimae, quae consurrexit adversum me: in solitudine hac deficiet et morietur ".
NUM|14|36|Igitur omnes viri, quos miserat Moyses ad contemplandam terram et qui reversi murmurare fecerant contra eum omnem congregationem detrahentes terrae quod esset mala,
NUM|14|37|mortui sunt atque percussi in conspectu Domini.
NUM|14|38|Iosue autem filius Nun et Chaleb filius Iephonne vixerunt ex omnibus, qui perrexerant ad considerandam terram.
NUM|14|39|Locutusque est Moyses universa verba haec ad omnes filios Israel, et luxit populus nimis.
NUM|14|40|Et ecce mane primo surgentes ascenderunt verticem montis atque dixerunt: " Parati sumus ascendere ad locum, de quo Dominus locutus est, quia peccavimus ".
NUM|14|41|Quibus Moyses: " Cur, inquit, transgredimini verbum Domini, quod vobis non cedet in prosperum?
NUM|14|42|Nolite ascendere, non enim est Dominus vobiscum, ne corruatis coram inimicis vestris!
NUM|14|43|Amalecites et Chananaeus ante vos sunt, quorum gladio corruetis, eo quod nolueritis acquiescere Domino, nec erit Dominus vobiscum ".
NUM|14|44|At illi contenebrati ascenderunt in verticem montis; arca autem foederis Domini et Moyses non recesserunt de castris.
NUM|14|45|Descenditque Amalecites et Chananaeus, qui habitabat in monte, et percutiens eos atque concidens persecutus est eos usque Horma.
NUM|15|1|Locutus est Dominus ad Moysen dicens:
NUM|15|2|" Loquere ad filios Israel et dices ad eos: Cum ingressi fueritis terram habitationis vestrae, quam ego dabo vobis,
NUM|15|3|et feceritis oblationem Domino in holocaustum aut victimam vota solventes vel sponte offerentes munera aut in sollemnitatibus vestris adolentes odorem suavitatis Domino de bobus sive de ovibus,
NUM|15|4|offeret, quicumque immolaverit victimam, sacrificium similae decimam partem ephi conspersae oleo, quod mensuram habebit quartam partem hin,
NUM|15|5|et vinum ad liba fundenda eiusdem mensurae dabit in holocaustum sive in victimam per agnos singulos.
NUM|15|6|Per arietes erit sacrificium similae duarum decimarum, quae conspersa sit oleo tertiae partis hin;
NUM|15|7|et vinum ad libamentum tertiae partis eiusdem mensurae offeret in odorem suavitatis Domino.
NUM|15|8|Quando vero de bobus feceris holocaustum aut hostiam, ut impleas votum vel pacificas victimas,
NUM|15|9|dabis per singulos boves similae tres decimas conspersae oleo, quod habeat medium mensurae hin,
NUM|15|10|et vinum ad liba fundenda eiusdem mensurae in oblationem suavissimi odoris Domino.
NUM|15|11|Sic facies per singulos boves et arietes et agnos et capras.
NUM|15|12|Secundum numerum victimarum quas offeretis, ita facietis singulis secundum numerum earum.
NUM|15|13|Omnis indigena eodem ritu offeret sacrificium ignis in odorem suavitatis Domino.
NUM|15|14|Et omnis peregrinus, qui habitat vobiscum vel qui commoratur in medio vestri in omnibus generationibus vestris, offeret sacrificium ignis in odorem suavitatis Domino eodem modo sicut et vos.
NUM|15|15|Unum praeceptum erit tam vobis quam advenis pro omnibus generationibus vestris coram Domino.
NUM|15|16|Una lex erit atque unum iudicium tam vobis quam advenis, qui vobiscum commorantur ".
NUM|15|17|Locutus est Dominus ad Moysen dicens:
NUM|15|18|" Loquere filiis Israel et dices ad eos: Cum veneritis in terram, quam dabo vobis,
NUM|15|19|et comederitis de panibus regionis illius, separabitis donaria Domino
NUM|15|20|de pulmento placentam. Sicut de areis donaria separatis,
NUM|15|21|ita et de pulmentis dabitis ea Domino.
NUM|15|22|Quod si per ignorantiam praeterieritis quidquam horum, quae locutus est Dominus ad Moysen
NUM|15|23|et mandavit per eum ad vos a die, qua coepit iubere et ultra ad generationes vestras,
NUM|15|24|si longe ab oculis congregationis, offeret congregatio vitulum de armento, holocaustum in odorem placabilem Domino et oblationem ac liba eius, ut caeremoniae postulant, hircumque pro peccato.
NUM|15|25|Et expiabit sacerdos pro omni congregatione filiorum Israel, et dimittetur eis, quoniam non sponte peccaverunt, nihilominus offerentes sacrificium ignis Domino pro se et pro peccato atque errore suo.
NUM|15|26|Et dimittetur universae plebi filiorum Israel et advenis, qui peregrinantur inter eos, quoniam culpa est omnis populi per ignorantiam.
NUM|15|27|Quod si anima una nesciens peccaverit, offeret capram anniculam pro peccato suo.
NUM|15|28|Et expiabit pro ea sacerdos, quod inscia peccaverit coram Domino; expiabit pro ea, et dimittetur illi.
NUM|15|29|Tam indigenis quam advenis una lex erit omnium, qui peccaverint ignorantes.
NUM|15|30|Anima vero, quae per superbiam aliquid commiserit, sive civis sit ille sive peregrinus, quoniam adversus Dominum rebellis fuit, peribit de populo suo.
NUM|15|31|Verbum enim Domini contempsit et praeceptum illius fecit irritum; idcirco delebitur et portabit iniquitatem suam ".
NUM|15|32|Factum est autem, cum essent filii Israel in solitudine et invenissent hominem colligentem ligna in die sabbati,
NUM|15|33|obtulerunt eum Moysi et Aaron et universae congregationi,
NUM|15|34|qui recluserunt eum in carcerem nescientes quid super eo facere deberent.
NUM|15|35|Dixitque Dominus ad Moysen: " Morte moriatur homo iste; obruat eum lapidibus omnis turba extra castra ".
NUM|15|36|Cumque eduxissent eum foras, obruerunt lapidibus; et mortuus est, sicut praeceperat Dominus.
NUM|15|37|Dixit quoque Dominus ad Moysen:
NUM|15|38|" Loquere filiis Israel et dices ad eos, ut faciant sibi fimbrias per angulos palliorum ponentes in eis vittas hyacinthinas.
NUM|15|39|Quas cum videbitis, recordabimini omnium mandatorum Domini eaque facietis nec sequamini cogitationes vestras et oculos per res varias fornicantes,
NUM|15|40|sed magis memores omnium praeceptorum meorum faciatis ea sitisque sancti Deo vestro.
NUM|15|41|Ego Dominus Deus vester, qui eduxi vos de terra Aegypti, ut essem Deus vester. Ego Dominus Deus vester ".
NUM|16|1|Ecce autem Core filius Isaar filii Caath filii Levi et Dathan atque Abiram filii Eliab, Hon quoque filius Pheleth de filiis Ruben
NUM|16|2|surrexerunt contra Moysen aliique filiorum Israel ducenti quinquaginta viri proceres synagogae vocati ad concilium, viri famosi.
NUM|16|3|Cumque stetissent adversum Moysen et Aaron, dixerunt: " Sufficiat vobis quia omnis congregatio sanctorum est, et in ipsis est Dominus! Cur elevamini super congregationem Domini? ".
NUM|16|4|Quod cum audisset Moyses, cecidit pronus in faciem
NUM|16|5|locutusque ad Core et ad omne concilium: " Mane, inquit, notum faciet Dominus qui ad se pertineant et qui sint sancti, et sanctos applicabit sibi; et, quos elegerit, appropinquare sibi faciet.
NUM|16|6|Hoc igitur facite: tollat unusquisque turibulum suum, tu, Core, et omne concilium tuum;
NUM|16|7|et hausto cras igne, ponite desuper thymiama coram Domino; et, quemcumque elegerit, ipse erit sanctus. Sufficiat vobis, filii Levi! ".
NUM|16|8|Dixitque rursum ad Core: " Audite, filii Levi.
NUM|16|9|Num parum vobis est quod separavit vos Deus Israel ab omni congregatione et iunxit sibi, ut serviretis ei in cultu habitaculi Domini et staretis coram frequentia populi et ministraretis pro ea?
NUM|16|10|Idcirco ad se fecit accedere te et omnes fratres tuos filios Levi, ut vobis etiam sacerdotium vindicetis,
NUM|16|11|et omne concilium tuum stet contra Dominum? Quid est enim Aaron, ut murmuretis contra eum? ".
NUM|16|12|Misit ergo Moyses, ut vocaret Dathan et Abiram filios Eliab, qui responderunt: " Non venimus!
NUM|16|13|Numquid parum est tibi quod eduxisti nos de terra, quae lacte et melle manabat, ut occideres in deserto, nisi et dominatus fueris nostri?
NUM|16|14|Revera non induxisti nos in terram, quae fluit rivis lactis et mellis, nec dedisti nobis possessiones agrorum et vinearum! An et oculos illorum hominum vis eruere? Non venimus! ".
NUM|16|15|Iratusque Moyses valde ait ad Dominum: " Ne respicias sacrificia eorum; tu scis quod ne asellum quidem umquam acceperim ab eis nec afflixerim quempiam eorum ".
NUM|16|16|Dixitque ad Core: " Tu et omne concilium tuum state seorsum coram Domino, et Aaron die crastino separatim.
NUM|16|17|Tollite singuli turibula vestra et ponite super ea incensum offerentes Domino ducenta quinquaginta turibula; tu et Aaron teneatis unusquisque turibulum suum ".
NUM|16|18|Quod cum fecissent, stantibus Moyse et Aaron,
NUM|16|19|et coacervasset Core adversum eos omne concilium ad ostium tabernaculi conventus, apparuit cunctis gloria Dornini.
NUM|16|20|Locutusque Dominus ad Moysen et Aaron ait:
NUM|16|21|" Separamini de medio congregationis huius, ut eos repente disperdam ".
NUM|16|22|Qui ceciderunt proni in faciem atque dixerunt: " Deus, Deus spirituum universae carnis; num, uno peccante, contra omnes ira tua desaeviet? ".
NUM|16|23|Et ait Dominus ad Moysen:
NUM|16|24|" Praecipe universo populo, ut separetur ab habitaculis Core et Dathan et Abiram ".
NUM|16|25|Surrexitque Moyses et abiit ad Dathan et Abiram et, sequentibus eum senioribus Israel,
NUM|16|26|dixit ad turbam: " Recedite ab habitaculis hominum impiorum et nolite tangere, quae ad eos pertinent, ne involvamini in peccatis eorum ".
NUM|16|27|Cumque recessissent a tentoriis eorum per circuitum, Dathan et Abiram egressi stabant in introitu papilionum suorum cum uxoribus et filiis et parvulis.
NUM|16|28|Et ait Moyses: " In hoc scietis quod Dominus miserit me, ut facerem universa, quae cernitis, et non ex proprio ea corde protulerim:
NUM|16|29|si consueta hominum morte interierint, et visitaverit eos plaga, qua et ceteri visitari solent, non misit me Dominus.
NUM|16|30|Sin autem novam rem fecerit Dominus, ut aperiens terra os suum deglutiat eos et omnia, quae ad illos pertinent, descenderintque viventes in infernum, scietis quod blasphemaverint Dominum ".
NUM|16|31|Confestim igitur, ut cessavit loqui, dirupta est terra sub pedibus eorum
NUM|16|32|et aperiens os suum devoravit illos cum domibus suis et omnibus hominibus Core et universa substantia eorum;
NUM|16|33|descenderuntque vivi in infernum operti humo et perierunt de medio congregationis.
NUM|16|34|At vero omnis Israel, qui stabat per gyrum, fugit ad clamorem pereuntium dicens: " Ne forte et nos terra deglutiat ".
NUM|16|35|Sed et ignis egressus a Domino interfecit ducentos quinquaginta viros, qui offerebant incensum.
NUM|17|1|Locutusque est Dominus ad Moysen dicens:
NUM|17|2|" Praecipe Eleazaro filio Aaron sacerdoti, ut tollat turibula, quae iacent in incendio, et ignem huc illucque dispergat, quoniam sanctificata sunt
NUM|17|3|in mortibus peccatorum; producatque ea in laminas et affigat altari, eo quod attulerunt ea Domino, et sanctificata sunt, ut sint pro signo filiis Israel ".
NUM|17|4|Tulit ergo Eleazar sacerdos turibula aenea, in quibus obtulerant hi, quos incendium devoravit, et produxit ea in laminas affigens altari,
NUM|17|5|ut haberent postea filii Israel, quibus commonerentur, ne quis accedat alienigena et, qui non est de semine Aaron, ad offerendum incensum Domino, ne patiatur sicut passus est Core et omnis congregatio eius, loquente Domino ad Moysen.
NUM|17|6|Murmuravit autem omnis congregatio filiorum Israel sequenti die contra Moysen et Aaron dicens: " Vos interfecistis populum Domini ".
NUM|17|7|Cumque oriretur seditio contra Moysen et Aaron, converterunt se ad tabernaculum conventus; quod operuit nubes, et apparuit gloria Domini.
NUM|17|8|Moyses et Aaron venerunt ante tabernaculum conventus.
NUM|17|9|Dixitque Dominus ad Moysen:
NUM|17|10|" Recedite de medio congregationis huius, nam extemplo delebo eos ". Et ceciderunt in faciem suam.
NUM|17|11|Dixit Moyses ad Aaron: " Tolle turibulum et, hausto igne de altari, mitte incensum desuper pergens cito ad populum, ut expies pro eis; iam enim egressa est ira a Domino, et plaga desaevit ".
NUM|17|12|Quod cum fecisset Aaron et cucurrisset ad mediam congregationem, quam iam vastabat plaga, obtulit thymiama et expiavit pro populo;
NUM|17|13|et stetit inter mortuos ac viventes, et plaga cessavit.
NUM|17|14|Fuerunt autem, qui percussi sunt, quattuordecim milia hominum et septingenti, absque his, qui perierant in seditione Core.
NUM|17|15|Reversusque est Aaron ad Moysen ad ostium tabernaculi conventus, postquam quievit interitus.
NUM|17|16|Et locutus est Dominus ad Moysen dicens:
NUM|17|17|" Loquere ad filios Israel et accipe ab eis virgas singulas per cognationes suas, a cunctis principibus tribuum virgas duodecim, et uniuscuiusque nomen superscribes virgae suae.
NUM|17|18|Nomen autem Aaron scribes in virga Levi, et una virga cunctas seorsum familias continebit.
NUM|17|19|Ponesque eas in tabernaculo conventus coram testimonio, ubi conveniam cum vobis.
NUM|17|20|Quem ex his elegero, germinabit virga eius; et cohibebo a me querimonias filiorum Israel, quibus contra vos murmurant ".
NUM|17|21|Locutusque est Moyses ad filios Israel, et dederunt ei omnes principes virgas per singulas tribus; fueruntque virgae duodecim, et virga Aaron in medio earum.
NUM|17|22|Quas cum posuisset Moyses coram Domino in tabernaculo testimonii,
NUM|17|23|sequenti die regressus invenit germinasse virgam Aaron in domo Levi; et turgentibus gemmis eruperant flores, qui, foliis dilatatis, in amygdalas deformati sunt.
NUM|17|24|Protulit ergo Moyses omnes virgas de conspectu Domini ad cunctos filios Israel; videruntque et receperunt singuli virgas suas.
NUM|17|25|Dixitque Dominus ad Moysen: " Refer virgam Aaron coram testimonio, ut servetur ibi in signum rebellium filiorum Israel, et quiescant querelae eorum a me, ne moriantur ".
NUM|17|26|Fecitque Moyses, sicut praeceperat Dominus.
NUM|17|27|Dixerunt autem filii Israel ad Moysen: " Ecce consumpti sumus, perimus, omnes perimus!
NUM|17|28|Quicumque accedit ad habitaculum Domini, moritur. Num usque ad internecionem cuncti delendi sumus? ".
NUM|18|1|Dixitque Dominus ad Aaron: " Tu et filii tui et domus patris tui tecum portabitis iniquitatem sanctuarii; et tu et filii tui simul sustinebitis peccata sacerdotii vestri.
NUM|18|2|Sed et fratres tuos de tribu Levi, tribum patris tui sume tecum, praestoque sint et ministrent tibi; tu autem et filii tui ministrabitis in tabernaculo testimonii.
NUM|18|3|Excubabuntque Levitae ad praecepta tua et ad cuncta opera tabernaculi, ita dumtaxat ut ad vasa sanctuarii et ad altare non accedant, ne et illi moriantur, et vos pereatis simul.
NUM|18|4|Sint autem tecum et excubent in custodiis tabernaculi conventus et in omni ministerio eius; alienigena non miscebitur vobis.
NUM|18|5|Excubate in ministerio sanctuarii et in ministerio altaris, ne oriatur amplius indignatio super filios Israel.
NUM|18|6|Ego sumpsi fratres vestros Levitas de medio filiorum Israel et tradidi donum Domino, ut serviant in ministeriis tabernaculi conventus.
NUM|18|7|Tu autem et filii tui custodite sacerdotium vestrum et omnia, quae ad cultum altaris pertinent et intra velum sunt, administrabitis. Ministerium do vobis sacerdotium in donum; si quis externus accesserit, occidetur ".
NUM|18|8|Locutusque est Dominus ad Aaron: " Ecce dedi tibi custodiam praelibationum mearum. Omnia, quae sanctificantur a filiis Israel, tradidi tibi et filiis tuis pro officio sacerdotali, legitima sempiterna.
NUM|18|9|Haec ergo accipies de sanctis sanctorum, exceptis his, quae comburuntur: omnis oblatio et sacrificium pro peccato atque delicto, quod redditur mihi, sanctum sanctorum tuum erit et filiorum tuorum.
NUM|18|10|In sanctuario comedes illud; mares tantum edent ex eo, quia consecratum est tibi.
NUM|18|11|Praelibationem donorum, quae elevando obtulerint filii Israel, tibi dedi et filiis tuis ac filiabus tuis iure perpetuo: qui mundus est in domo tua, vescetur eis.
NUM|18|12|Omnem medullam olei et vini ac frumenti quidquid offerunt primitiarum Domino, tibi dedi.
NUM|18|13|Universa frugum initia, quas gignit humus et Domino deportantur, cedent in usus tuos: qui mundus est in domo tua, vescetur eis.
NUM|18|14|Omne, quod ex voto reddiderint filii Israel, tuum erit.
NUM|18|15|Quidquid primum erumpit e vulva cunctae carnis, quod offerunt Domino, sive ex hominibus sive de pecoribus fuerit, tui iuris erit; ita dumtaxat, ut hominis primogenitum et omne animal, quod immundum est, redimi facias.
NUM|18|16|Cuius redemptio erit post unum mensem siclis argenti quinque pondere sanctuarii. Siclus viginti obolos habet.
NUM|18|17|Primogenitum autem bovis vel ovis vel caprae non facies redimi, quia sanctificata sunt Domino; sanguinem tantum eorum fundes super altare et adipes adolebis in suavissimum odorem Domino.
NUM|18|18|Carnes vero eorum in usum tuum cedent, sicut pectusculum elevatum et armus dexter tua erunt.
NUM|18|19|Omnes praelibationes sanctas, quas offerunt filii Israel Domino, tibi dedi et filiis ac filiabus tuis iure perpetuo: pactum salis est sempiternum coram Domino tibi ac filiis tuis ".
NUM|18|20|Dixitque Dominus ad Aaron: " In terra eorum nihil possidebitis nec habebitis partem inter eos: Ego pars et hereditas tua in medio filiorum Israel.
NUM|18|21|Filiis autem Levi dedi omnes decimas Israelis in possessionem pro ministerio, quo serviunt mihi in tabernaculo conventus,
NUM|18|22|ut non accedant ultra filii Israel ad tabernaculum conventus nec committant peccatum mortiferum.
NUM|18|23|Solis filiis Levi mihi in tabernaculo conventus servientibus et portantibus peccata populi; legitimum sempiternum erit in generationibus vestris, et in medio filiorum Israel nihil aliud possidebunt.
NUM|18|24|Decimas, quas filii Israel in praelibationem elevant Domino, dedi Levitis in possessionem. Propterea dixi eis: In medio filiorum Israel non habebitis possessionem ".
NUM|18|25|Locutusque est Dominus ad Moysen dicens:
NUM|18|26|" Praecipe Levitis atque denuntia: Cum acceperitis a filiis Israel decimas, quas dedi vobis, praelibationem earum elevabitis Domino, id est decimam partem decimae,
NUM|18|27|ut reputetur vobis in praelibationem tam de areis quam de torcularibus.
NUM|18|28|Sic de universis, quorum accipitis primitias a filiis Israel, elevate Domino: date Aaron sacerdoti.
NUM|18|29|Omnia, quae offeretis ex decimis, in donaria Domini separabitis: optima et electa erunt.
NUM|18|30|Dicesque ad eos: Si praeclara et meliora quaeque obtuleritis ex decimis, reputabitur vobis quasi de area et torculari dederitis fructus;
NUM|18|31|et comedetis eas in omnibus locis vestris, tam vos quam familiae vestrae, quia pretium est pro ministerio, quo servitis in tabernaculo conventus.
NUM|18|32|Et non peccabitis super hoc egregia vobis et pinguia reservantes, ne polluatis oblationes filiorum Israel et moriamini ".
NUM|19|1|Locutusque est Dominus ad Moysen et Aaron dicens:
NUM|19|2|" Ista est religio legis, quam constituit Dominus. Praecipe filiis Israel, ut adducant ad te vaccam rufam aetatis integrae, in qua nulla sit macula, nec portaverit iugum.
NUM|19|3|Tradetisque eam Eleazaro sacerdoti, quae educta extra castra mactabitur in conspectu eius;
NUM|19|4|et tinguens digitum in sanguine eius asperget contra fores tabernaculi conventus septem vicibus,
NUM|19|5|combureturque in conspectu eius, tam pelle et carnibus eius quam sanguine et fimo flammae traditis.
NUM|19|6|Lignum quoque cedrinum et hyssopum coccumque sacerdos mittet in flammam, quae vaccam vorat.
NUM|19|7|Et tunc demum, lotis vestibus et corpore suo, ingredietur in castra commaculatusque erit usque ad vesperum.
NUM|19|8|Sed et ille, qui combusserit eam, lavabit vestimenta sua et corpus, et immundus erit usque ad vesperum.
NUM|19|9|Colliget autem vir mundus cineres vaccae et effundet eos extra castra in loco purissimo, ut sint congregationi filiorum Israel in custodiam pro aqua aspersionis.
NUM|19|10|Cumque laverit, qui vaccae portaverat cineres, vestimenta sua, immundus erit usque ad vesperum. Habebunt hoc filii Israel et advenae, qui habitant inter eos, sanctum iure perpetuo.
NUM|19|11|Qui tetigerit cadaver hominis et propter hoc septem diebus fuerit immundus,
NUM|19|12|aspergetur ex hac aqua die tertio et septimo et sic mundabitur. Si die tertio aspersus non fuerit, septimo non erit mundus.
NUM|19|13|Omnis, qui tetigerit humanae animae morticinum et aspersus hac commixtione non fuerit, polluet habitaculum Domini et peribit ex Israel, quia aqua expiationis non est aspersus: immundus erit, et manebit spurcitia eius super eum.
NUM|19|14|Ista est lex hominis, qui moritur in tabernaculo: omnes, qui ingrediuntur tentorium illius, et universa vasa, quae ibi sunt, polluta erunt septem diebus.
NUM|19|15|Vas, quod non habuerit operculum nec ligaturam desuper, immundum erit.
NUM|19|16|Si quis in agro tetigerit cadaver hominis gladio occisi aut per se mortui sive os illius vel sepulcrum, immundus erit septem diebus.
NUM|19|17|Tollentque de cineribus combustionis peccati et mittent aquas vivas super eos in vas;
NUM|19|18|in quibus cum homo mundus tinxerit hyssopum, asperget ex eo omne tentorium et cunctam supellectilem et homines, qui ibi fuerint, et super eum, qui tetigerit ossa vel occisum hominem aut per se mortuum aut sepultum.
NUM|19|19|Atque hoc modo mundus lustrabit immundum tertio et septimo die; expiatusque die septimo lavabit et se et vestimenta sua et mundus erit ad vesperum.
NUM|19|20|Si quis hoc ritu non fuerit expiatus, peribit anima illius de medio ecclesiae, quia sanctuarium Domini polluit et non est aqua lustrationis aspersus; immundus est.
NUM|19|21|Erit vobis praeceptum legitimum sempiternum. Ipse quoque, qui aspergit aqua lustrali, lavabit vestimenta sua; omnis, qui tetigerit aquas expiationis, immundus erit usque ad vesperum.
NUM|19|22|Quidquid tetigerit immundus, immundum erit, et anima, quae horum quippiam tetigerit, immunda erit usque ad vesperum ".
NUM|20|1|Veneruntque filii Israel et omnis congregatio in de sertum Sin mense primo, et mansit populus in Cades. Mortuaque est ibi Maria et sepulta in eodem loco.
NUM|20|2|Cumque indigeret aqua populus, convenerunt adversum Moysen et Aaron
NUM|20|3|et versi in seditionem dixerunt: " Utinam perissemus inter fratres nostros coram Domino!
NUM|20|4|Cur eduxistis ecclesiam Domini in solitudinem, ut et nos et nostra iumenta moriamur?
NUM|20|5|Quare nos fecistis ascendere de Aegypto et adduxistis in locum istum pessimum, qui seri non potest, qui nec ficum gignit nec vineas nec malogranata, insuper et aquam non habet ad bibendum? ".
NUM|20|6|Venitque Moyses et Aaron, relicta congregatione, ad introitum tabernaculi conventus corrueruntque proni in terram, et apparuit gloria Domini super eos.
NUM|20|7|Locutusque est Dominus ad Moysen dicens:
NUM|20|8|" Tolle virgam et congrega populum, tu et Aaron frater tuus; et loquimini ad petram coram eis, et illa dabit aquas. Cumque eduxeris aquam de petra, potabis congregationem et iumenta eius ".
NUM|20|9|Tulit igitur Moyses virgam, quae erat in conspectu Domini, sicut praeceperat ei.
NUM|20|10|Et congregaverunt Moyses et Aaron populum ante petram, dixitque eis: " Audite, rebelles; num de petra hac vobis aquam poterimus eicere? ".
NUM|20|11|Cumque elevasset Moyses manum percutiens virga bis silicem, egressae sunt aquae largissimae, ita ut populus biberet et iumenta.
NUM|20|12|Dixitque Dominus ad Moysen et Aaron: " Quia non credidistis mihi, ut sanctificaretis me coram filiis Israel, non introducetis hos populos in terram, quam dabo eis ".
NUM|20|13|Hae sunt aquae Meriba, ubi iurgati sunt filii Israel contra Dominum, et sanctificatus est in eis.
NUM|20|14|Misit nuntios Moyses de Cades ad regem Edom, qui dicerent: " Haec mandat frater tuus Israel: Nosti omnem laborem, qui apprehendit nos,
NUM|20|15|quomodo descenderint patres nostri in Aegyptum, et habitaverimus ibi multo tempore, afflixerintque nos Aegyptii et patres nostros,
NUM|20|16|et quomodo clamaverimus ad Dominum, et exaudierit nos miseritque angelum, qui eduxerit nos de Aegypto. Ecce nos in urbe Cades, quae est in extremis finibus tuis, positi
NUM|20|17|obsecramus, ut nobis transire liceat per terram tuam: non ibimus per agros nec per vineas, non bibemus aquas de puteis tuis; sed gradiemur via regia, nec ad dexteram nec ad sinistram declinantes, donec transeamus terminos tuos ".
NUM|20|18|Cui respondit Edom: " Non transibis per me, alioquin armatus occurram tibi ".
NUM|20|19|Dixeruntque filii Israel: " Per tritam gradiemur viam et, si biberimus aquas tuas ego et pecora mea, dabo, quod iustum est: nulla erit in pretio difficultas; tantum velociter transeamus ".
NUM|20|20|At ille respondit: " Non transibis! ". Statimque egressus est obvius cum infinita multitudine et manu forti
NUM|20|21|nec voluit acquiescere Israeli, ut concederet transitum per fines suos; quam ob rem divertit ab eo Israel.
NUM|20|22|Cumque castra movissent de Cades, venerunt in montem Hor,
NUM|20|23|ubi locutus est Dominus ad Moysen et Aaron in monte Hor, qui est in finibus terrae Edom:
NUM|20|24|" Congregabitur, inquit, Aaron ad populum suum. Non enim intrabit terram, quam dedi filiis Israel, eo quod rebelles fuistis ori meo ad aquas Meriba.
NUM|20|25|Tolle Aaron et Eleazarum filium eius cum eo et duces eos in montem Hor.
NUM|20|26|Cumque nudaveris patrem veste sua, indues ea Eleazarum filium eius: Aaron colligetur et morietur ibi ".
NUM|20|27|Fecit Moyses, ut praeceperat Dominus, et ascenderunt in montem Hor coram omni congregatione.
NUM|20|28|Cumque Aaron spoliasset vestibus suis, induit eis Eleazarum filium eius. Illo mortuo in montis supercilio, descendit cum Eleazaro.
NUM|20|29|Omnis autem congregatio videns occubuisse Aaron flevit super eo triginta diebus tota domus Israel.
NUM|21|1|Quod cum audisset Chana naeus rex Arad, qui habita bat in Nageb, venisse scilicet Israel per viam Atarim, pugnavit contra illum et duxit ex eo captivos.
NUM|21|2|At Israel voto se Domino obligans ait: " Si tradideris populum istum in manu mea, delebo urbes eius ".
NUM|21|3|Exaudivitque Dominus preces Israel et tradidit Chananaeum, quem ille interfecit, subversis urbibus eius, et vocavit nomen loci illius Horma.
NUM|21|4|Profecti sunt autem et de monte Hor per viam, quae ducit ad mare Rubrum, ut circumirent terram Edom. Et taedere coepit populum itineris.
NUM|21|5|Locutusque contra Deum et Moysen ait: " Cur eduxisti nos de Aegypto, ut moreremur in solitudine? Deest panis, non sunt aquae; anima nostra iam nauseat super cibo isto levissimo ".
NUM|21|6|Quam ob rem misit Dominus in populum ignitos serpentes, qui mordebant populum, et mortuus est populus multus ex Israel.
NUM|21|7|Et venerunt ad Moysen atque dixerunt: " Peccavimus, quia locuti sumus contra Dominum et te; ora, ut tollat a nobis serpentes ". Oravitque Moyses pro populo.
NUM|21|8|Et locutus est Dominus ad eum: " Fac serpentem ignitum et pone eum pro signo: qui percussus aspexerit eum, vivet ".
NUM|21|9|Fecit ergo Moyses serpentem aeneum et posuit eum pro signo; quem cum percussi aspicerent, sanabantur.
NUM|21|10|Profectique filii Israel castrametati sunt in Oboth,
NUM|21|11|unde egressi fixere tentoria in Ieabarim, in solitudine, quae respicit Moab contra orientalem plagam.
NUM|21|12|Et inde moventes venerunt ad torrentem Zared;
NUM|21|13|quem relinquentes castrametati sunt ultra Arnon, qui est in deserto, quod prominet de finibus Amorraei. Siquidem Arnon terminus est Moab dividens Moabitas et Amorraeos.
NUM|21|14|Unde dicitur in libro bellorum Domini:" Vaheb in Suphaet torrentes Arnon.
NUM|21|15|Scopuli torrentium inclinati suntin habitationem Aret recumbunt in finibus Moabitarum ".
NUM|21|16|Ex eo loco in Beer. Hic est puteus, super quo locutus est Dominus ad Moysen: " Congrega populum, et dabo ei aquam ".
NUM|21|17|Tunc cecinit Israel carmen istud:" Ascendat puteus. Concinite ei.
NUM|21|18|Puteus, quem foderunt principeset paraverunt duces populiin sceptris et in baculis suis ".De solitudine in Matthana;
NUM|21|19|de Matthana in Nahaliel; de Nahaliel in Bamoth;
NUM|21|20|de Bamoth in vallem, quae est in regione Moab in vertice Phasga, qui respicit contra desertum.
NUM|21|21|Misit autem Israel nuntios ad Sehon regem Amorraeorum dicens:
NUM|21|22|" Obsecro, ut transire mihi liceat per terram tuam: non declinabimus in agros et vineas, non bibemus aquas ex puteis. Via regia gradiemur, donec transeamus terminos tuos ".
NUM|21|23|Qui concedere noluit, ut transiret Israel per fines suos; quin potius, populo congregato, egressus est obviam in desertum et venit in Iasa pugnavitque contra Israel.
NUM|21|24|A quo percussus est in ore gladii, et possessa est terra eius ab Arnon usque Iaboc et filios Ammon; quia forti praesidio tenebantur termini Ammonitarum.
NUM|21|25|Tulit ergo Israel omnes civitates eius et habitavit in urbibus Amorraei, in Hesebon scilicet et viculis eius.
NUM|21|26|Hesebon enim erat urbs Sehon regis Amorraei, qui pugnavit contra primum regem Moab et tulit omnem terram, quae dicionis illius fuerat usque Arnon.
NUM|21|27|Idcirco dicitur in proverbio:" Venite in Hesebon!Aedificetur et construatur civitas Sehon!
NUM|21|28|Ignis egressus est de Hesebon,flamma de oppido Sehonet devoravit Ar Moabitarumet deglutivit excelsa Arnon.
NUM|21|29|Vae tibi, Moab;peristi, popule Chamos!Dedit filios eius in fugamet filias in captivitatemregi Amorraeorum Sehon.
NUM|21|30|Iecimus sagittas in eos,disperiit Hesebon usque Dibon.Vastavimus usque Nopheet usque Medaba ".
NUM|21|31|Habitavit itaque Israel in terra Amorraei.
NUM|21|32|Misitque Moyses, qui explorarent Iazer, cuius ceperunt viculos et expulerunt Amorraeos, qui erant ibi.
NUM|21|33|Verteruntque se et ascenderunt per viam Basan, et occurrit eis Og rex Basan cum omni populo suo pugnaturus in Edrai.
NUM|21|34|Dixitque Dominus ad Moysen: " Ne timeas eum, quia in manu tua tradidi illum et omnem populum ac terram eius, faciesque illi, sicut fecisti Sehon regi Amorraeorum habitatori Hesebon ".
NUM|21|35|Percusserunt igitur et hunc cum filiis suis universumque populum eius usque ad internecionem; et possederunt terram illius.
NUM|22|1|Profectique castrametati sunt filii Israel in campestri bus Moab, ubi trans Iordanem Iericho sita est.
NUM|22|2|Videns autem Balac filius Sephor omnia, quae fecerat Israel Amorraeo,
NUM|22|3|valde metuit Moab populum, quia multus erat. Et cum pertimeret Moab filios Israel,
NUM|22|4|dixit ad maiores natu Madian: " Nunc carpet haec congregatio omnem regionem per circuitum, quomodo solet bos herbas campi carpere ".Balac filius Sephor erat eo tempore rex in Moab.
NUM|22|5|Misit ergo nuntios ad Balaam filium Beor in Phethor, quae est super flumen in terra filiorum Ammau, ut vocarent eum et dicerent: " Ecce egressus est populus ex Aegypto, qui operuit superficiem terrae sedens contra me.
NUM|22|6|Veni igitur et maledic populo huic, quia fortior me est; si quo modo possim percutere et eicere eum de terra mea. Novi enim quod benedictus sit, cui benedixeris, et maledictus, in quem maledicta congesseris ".
NUM|22|7|Perrexeruntque seniores Moab et maiores natu Madian habentes divinationis pretium in manibus. Cumque venissent ad Balaam et narrassent ei omnia verba Balac,
NUM|22|8|ille respondit: " Manete hic nocte, et respondebo quidquid mihi dixerit Dominus ". Manentibus illis apud Balaam,
NUM|22|9|venit Deus et ait ad eum: " Quid sibi volunt homines isti apud te? ".
NUM|22|10|Respondit: " Balac filius Sephor rex Moabitarum misit ad me
NUM|22|11|dicens: "Ecce populus, qui egressus est de Aegypto, operuit superficiem terrae; veni et maledic ei pro me, si quo modo possim pugnans abigere eum".
NUM|22|12|Dixitque Deus ad Balaam: "Noli ire cum eis neque maledicas populo, quia benedictus est ".
NUM|22|13|Qui mane consurgens dixit ad principes: " Ite in terram vestram, quia prohibuit me Dominus venire vobiscum ".
NUM|22|14|Reversi principes dixerunt ad Balac: " Noluit Balaam venire nobiscum ".
NUM|22|15|Rursum ille multo plures et nobiliores, quam ante miserat, misit.
NUM|22|16|Qui cum venissent ad Balaam, dixerunt: " Sic dicit Balac filius Sephor: "Ne cuncteris venire ad me;
NUM|22|17|paratus sum honorare te et, quidquid volueris, dabo tibi. Veni et maledic pro me populo isti" ".
NUM|22|18|Respondit Balaam: " Si dederit mihi Balac plenam domum suam argenti et auri, non potero transgredi verbum Domini Dei mei, ut vel plus vel minus loquar.
NUM|22|19|Obsecro, ut hic maneatis etiam hac nocte, et scire queam quid mihi rursum respondeat Dominus ".
NUM|22|20|Venit ergo Deus ad Balaam nocte et ait ei: " Si vocare te venerunt homines isti, surge et vade cum eis, ita dumtaxat, ut, quod tibi praecepero, facias ".
NUM|22|21|Surrexit Balaam mane et, strata asina sua, profectus est cum eis.
NUM|22|22|Et iratus est Deus, cum profectus esset; stetitque angelus Domini in via contra Balaam, ut adversaretur ei, qui insidebat asinae et duos pueros habebat secum.
NUM|22|23|Cernens asina angelum Domini stantem in via, evaginato gladio in manu sua, avertit se de itinere et ibat per agrum. Quam cum verberaret Balaam et vellet ad semitam reducere,
NUM|22|24|stetit angelus Domini in angustiis duarum maceriarum, quibus vineae cingebantur.
NUM|22|25|Quem videns asina iunxit se parieti et attrivit sedentis pedem. At ille iterum verberabat eam;
NUM|22|26|et angelus Domini iterum transiens ad locum angustum, ubi nec ad dexteram nec ad sinistram poterat deviare, obvius stetit.
NUM|22|27|Cumque vidisset asina stantem angelum Domini, concidit sub pedibus sedentis; qui iratus vehementius caedebat fuste latera eius.
NUM|22|28|Aperuitque Dominus os asinae, et locuta est: " Quid feci tibi? Cur percutis me ecce iam tertio? ".
NUM|22|29|Respondit Balaam: " Quia illusisti mihi. Utinam haberem gladium, ut te interficerem! ".
NUM|22|30|Dixit asina: " Nonne animal tuum sum, cui semper sedere consuevisti usque in praesentem diem? Dic quid simile umquam fecerim tibi ". At ille ait: " Numquam ".
NUM|22|31|Protinus aperuit Dominus oculos Balaam, et vidit angelum Domini stantem in via, evaginato gladio in manu eius; adoravitque eum pronus in terram.
NUM|22|32|Cui angelus Domini: " Cur, inquit, tertio verberas asinam tuam? Ego veni, ut adversarer tibi, quia perversa est via tua mihique contraria.
NUM|22|33|Et videns me asina declinavit ter a me; nisi declinasset, te occidissem et illam vivam reliquissem ".
NUM|22|34|Dixit Balaam: " Peccavi nesciens quod tu stares contra me in via; et nunc, si displicet tibi, revertar ".
NUM|22|35|Ait angelus Domini: " Vade cum istis et cave, ne aliud, quam praecepero tibi, loquaris ". Ivit igitur cum principibus Balac.
NUM|22|36|Quod cum audisset Balac, venisse scilicet Balaam, egressus est in occursum eius in Irmoab, quod situm est in extremis finibus Arnon;
NUM|22|37|dixitque ad Balaam: " Nonne misi nuntios, ut vocarem te? Cur non statim venisti ad me? An quia honorare te nequeo? ".
NUM|22|38|Cui ille respondit: " Ecce adsum; numquid loqui potero aliud, nisi quod Deus posuerit in ore meo? ".
NUM|22|39|Perrexerunt ergo simul et venerunt in Cariathusoth.
NUM|22|40|Cumque occidisset Balac boves et oves, misit ad Balaam et principes, qui cum eo erant.
NUM|22|41|Mane autem facto, duxit eum ad excelsa Baal et intuitus est extremam partem populi.
NUM|23|1|Dixitque Balaam ad Balac: " Aedifica mihi hic septem aras et para totidem vitulos eiusdemque numeri arietes ".
NUM|23|2|Cumque fecisset iuxta sermonem Balaam, imposuerunt vitulum et arietem super aram.
NUM|23|3|Dixitque Balaam ad Balac: " Sta paulisper iuxta holocaustum tuum, donec vadam, si forte occurrat mihi Dominus; et, quodcumque imperaverit, loquar tibi ". Cumque abiisset in collem nudum,
NUM|23|4|occurrit illi Deus. Locutusque ad eum Balaam: " Septem, inquit, aras erexi et imposui vitulum et arietem desuper ".
NUM|23|5|Dominus autem posuit verbum in ore eius et ait: " Revertere ad Balac et haec loqueris ".
NUM|23|6|Reversus invenit stantem Balac iuxta holocaustum suum et omnes principes Moabitarum;
NUM|23|7|assumptaque parabola sua, dixit:" De Aram adduxit me Balac,rex Moabitarum de montibus orientis:"Veni, inquit, et maledic pro me Iacob;propera et detestare Israel!".
NUM|23|8|Quomodo maledicam, cui non maledixit Deus?Qua ratione detester, quem Dominus non detestatur?
NUM|23|9|De summis silicibus video eumet de collibus considero illum:populus solus habitabitet inter gentes non reputabitur.
NUM|23|10|Et quis dinumerare possit pulverem Iacobet quis numeravit arenam Israel?Moriatur anima mea morte iustorum,et fiant novissima mea horum similia ".
NUM|23|11|Dixitque Balac ad Balaam: " Quid est hoc, quod agis? Ut malediceres inimicis meis, vocavi te, et tu e contrario benedicis eis! ".
NUM|23|12|Cui ille respondit: " Num aliud possum loqui, nisi quod iusserit Dominus? ".
NUM|23|13|Dixit ergo Balac: " Veni mecum in alterum locum, unde partem Israel videas et totum videre non possis; inde maledicito ei ".
NUM|23|14|Cumque duxisset eum in campum speculatorum super verticem montis Phasga, aedificavit septem aras imposuitque supra vitulum atque arietem.
NUM|23|15|Et dixit Balaam ad Balac: " Sta hic iuxta holocaustum tuum, donec ego obvius pergam ".
NUM|23|16|Cui cum Dominus occurrisset posuissetque verbum in ore eius, ait: " Revertere ad Balac et haec loqueris ei ".
NUM|23|17|Reversus invenit eum stantem iuxta holocaustum suum et principes Moabitarum cum eo. Ad quem Balac: " Quid, inquit, locutus est Dominus? ".
NUM|23|18|At ille, assumpta parabola sua, ait:" Surge, Balac, et ausculta;audi, fili Sephor.
NUM|23|19|Non est Deus quasi homo, ut mentiatur,nec ut filius hominis, ut mutetur.Numquid dixit et non faciet?Locutus est et non implebit?
NUM|23|20|Ad benedicendum adductus sum,benedictionem prohibere non valeo.
NUM|23|21|Non conspicitur malum in Iacob,nec videtur calamitas in Israel.Dominus Deus eius cum eo est,et clangor regis in illo.
NUM|23|22|Deus eduxit illum de Aegypto,sicut cornua bubali est ei.
NUM|23|23|Non est augurium in Iacob,nec divinatio in Israel.Temporibus suis dicetur Iacob et Israeliquid operatus sit Deus.
NUM|23|24|Ecce populus ut leaena consurget,et quasi leo erigetur;non accubabit, donec devoret praedamet occisorum sanguinem bibat ".
NUM|23|25|Dixitque Balac ad Balaam: " Nec maledicas ei, nec benedicas! ".
NUM|23|26|Et ille ait: " Nonne dixi tibi quod, quidquid mihi Dominus imperaret, hoc facerem? ".
NUM|23|27|Et ait Balac ad eum: " Veni, et ducam te ad alîum locum, si forte placeat Deo, ut inde maledicas ei ".
NUM|23|28|Cumque duxisset eum super verticem montis Phegor, qui respicit solitudinem,
NUM|23|29|dixit ei Balaam: " Aedifica mihi hic septem aras et para totidem vitulos eiusdemque numeri arietes ".
NUM|23|30|Fecit Balac, ut Balaam dixerat, imposuitque vitulos et arietes per singulas aras.
NUM|24|1|Cumque vidisset Balaam quod placeret Domino, ut be nediceret Israeli, nequaquam abiit, ut ante perrexerat, ut augurium quaereret; sed dirigens contra desertum vultum suum
NUM|24|2|et elevans oculos vidit Israel commorantem per tribus suas et, irruente in se spiritu Dei,
NUM|24|3|assumpta parabola sua, ait:" Dixit Balaam filius Beor,dixit homo, cuius apertus est oculus,
NUM|24|4|dixit auditor sermonum Dei,qui visionem Omnipotentis intuitus est,qui cadit, et sic aperiuntur oculi eius.
NUM|24|5|Quam pulchra tabernacula tua, Iacob,et tentoria tua, Israel!
NUM|24|6|Ut valles dilatantur,ut horti iuxta fluvios irrigui,ut aloe, quam plantavit Dominus,quasi cedri prope aquas.
NUM|24|7|Fluet aqua de situlis eius,et semen illius erit in aquis multis. Extolletur super Agag rex eius,et elevabitur regnum illius.
NUM|24|8|Deus eduxit illum de Aegypto,sicut cornua bubali est ei.Devorabit gentes, hostes suos,ossaque eorum confringetet perforabit sagittis.
NUM|24|9|Accubans dormit ut leo,et quasi leaena, quis suscitare illum audebit?Qui benedixerit tibi, erit et ipse benedictus;qui maledixerit tibi, maledictus erit! ".
NUM|24|10|Iratusque Balac contra Balaam, complosis manibus, ait: " Ad maledicendum inimicis meis vocavi te, quibus iam tertio benedixisti!
NUM|24|11|Revertere nunc ad locum tuum! Decreveram quidem magnifice honorare te, sed Dominus privavit te honore disposito ".
NUM|24|12|Respondit Balaam ad Balac: " Nonne iam nuntiis tuis, quos misisti ad me, dixi:
NUM|24|13|Si dederit mihi Balac plenam domum suam argenti et auri, non potero praeterire sermonem Domini, ut vel boni quid vel mali proferam ex corde meo, sed, quidquid Dominus dixerit, hoc loquar?
NUM|24|14|Et nunc, pergens ad populum meum dabo consilium, quid populus hic populo tuo faciat extremo tempore ".
NUM|24|15|Sumpta igitur parabola sua, rursum ait:" Dixit Balaam filius Beor,dixit homo, cuius apertus est oculus,
NUM|24|16|dixit auditor sermonum Dei,qui novit doctrinam Altissimiet visiones Omnipotentis videt,qui cadens apertos habet oculos.
NUM|24|17|Video eum, sed non modo;intueor illum, sed non prope.Oritur stella ex Iacob,et consurgit virga de Israel;et percutit tempora Moabet verticem omnium filiorum Seth.
NUM|24|18|Et erit Idumaea possessio eius,et hereditas eius Seir, inimicus eius; Israel vero fortiter aget.
NUM|24|19|De Iacob erit, qui domineturet perdat reliquias civitatis ".
NUM|24|20|Cumque vidisset Amalec, assumens parabolam suam ait:" Principium gentium Amalec,cuius extrema perdentur ".
NUM|24|21|Vidit quoque Cinaeum et, assumpta parabola sua, ait:" Robustum quidem est habitaculum tuum,et in petra positus nidus tuus.
NUM|24|22|Erit in combustionem Cain,donec Assur capiat te ".
NUM|24|23|Assumptaque parabola sua, iterum locutus est:" Heu! Quis vivet,quando ista faciet Deus?
NUM|24|24|Venient naves de Cetthim,superabunt Assyrios vastabuntque Heber;et ad extremum etiam ipsi peribunt ".Surrexitque Balaam et reversus est in locum suum; Balac quoque via, qua venerat, rediit.
NUM|25|1|Morabatur autem Israel in Settim, et incepit populus fornicari cum filiabus Moab,
NUM|25|2|quae vocaverunt populum ad sacrificia deorum suorum. Et illi comederunt et adoraverunt deos earum;
NUM|25|3|et adhaesit Israel Baalphegor. Et iratus Dominus
NUM|25|4|ait ad Moysen: " Tolle cunctos principes populi et suspende eos coram Domino contra solem in patibulis, ut avertatur furor meus ab Israel ".
NUM|25|5|Dixitque Moyses ad iudices Israel: " Occidat unusquisque proximos suos, qui adhaeserunt Baalphegor ".
NUM|25|6|Et ecce unus de filiis Israel intravit coram fratribus suis ad Madianitin, vidente Moyse et omni turba filiorum Israel, qui flebant ante fores tabernaculi conventus.
NUM|25|7|Quod cum vidisset Phinees filius Eleazari filii Aaron sacerdotis, surrexit de medio congregationis et, arrepta lancea,
NUM|25|8|ingressus est post virum Israelitem in cubiculum et perfodit ambos simul, virum scilicet et mulierem, in locis genitalibus; cessavitque plaga a filiis Israel.
NUM|25|9|Et occisi sunt viginti quattuor milia hominum.
NUM|25|10|Dixitque Dominus ad Moysen:
NUM|25|11|" Phinees filius Eleazari filii Aaron sacerdotis avertit iram meam a filiis Israel, quia zelo meo commotus est in medio eorum, ut non ipse delerem filios Israel in zelo meo.
NUM|25|12|Idcirco loquere ad eum: Ecce do ei pacem foederis mei,
NUM|25|13|et erit tam ipsi quam semini eius pactum sacerdotii sempiternum, quia zelatus est pro Deo suo et expiavit scelus filiorum Israel ".
NUM|25|14|Erat autem nomen viri Israelitae, qui occisus est cum Madianitide, Zamri filius Salu dux de cognatione et tribu Simeonis;
NUM|25|15|porro mulier Madianitis, quae pariter interfecta est, vocabatur Cozbi filia Sur principis tribus in Madian.
NUM|25|16|Locutusque est Dominus ad Moysen dicens:
NUM|25|17|" Pugnate contra Madianitas et percutite eos,
NUM|25|18|quia ipsi hostiliter egerunt contra vos et decepere insidiis per idolum Phegor et in negotio Cozbi filiae ducis Madian sororis eorum, quae percussa est in die plagae pro sacrilegio Phegor ".
NUM|26|1|Post hanc plagam dixit Do minus ad Moysen et Eleaza rum filium Aaron sacerdotem:
NUM|26|2|" Numerate summam totius congregationis filiorum Israel a viginti annis et supra per domos et cognationes suas, cunctos, qui possunt ad bella procedere ".
NUM|26|3|Locuti sunt itaque Moyses et Eleazar sacerdos in campestribus Moab super Iordanem contra Iericho ad eos, qui erant
NUM|26|4|a viginti annis et supra, sicut Dominus imperaverat Moysi.Filiorum Israel, qui egressi sunt de terra Aegypti, iste est numerus.
NUM|26|5|Ruben primogenitus Israel. Huius filius Henoch, a quo familia Henochitarum, et Phallu, a quo familia Phalluitarum,
NUM|26|6|et Hesron, a quo familia Hesronitarum, et Charmi, a quo familia Charmitarum.
NUM|26|7|Hae sunt familiae de stirpe Ruben, quarum numerus inventus est quadraginta tria milia et septingenti triginta.
NUM|26|8|Filius Phallu: Eliab.
NUM|26|9|Huius filii: Namuel et Dathan et Abiram. Isti sunt Dathan et Abiram principes populi, qui surrexerunt contra Moysen et Aaron in seditione Core, quando adversus Dominum rebellaverunt,
NUM|26|10|et aperiens terra os suum devoravit eos et Core, morientibus plurimis, quando combussit ignis ducentos quinquaginta viros; et facti sunt in signum.
NUM|26|11|Core pereunte, filii illius non perierunt.
NUM|26|12|Filii Simeon per cognationes suas: Namuel, ab hoc familia Namuelitarum; Iamin, ab hoc familia Iaminitarum; Iachin, ab hoc familia Iachinitarum;
NUM|26|13|Zara, ab hoc familia Zaraitarum; Saul, ab hoc familia Saulitarum.
NUM|26|14|Hae sunt familiae de stirpe Simeon, quarum omnis numerus fuit viginti duo milia ducenti.
NUM|26|15|Filii Gad per cognationes suas: Sephon, ab hoc familia Sephonitarum; Haggi, ab hoc familia Haggitarum; Suni, ab hoc familia Sunitarum;
NUM|26|16|Ozni, ab hoc familia Oznitarum; Heri, ab hoc familia Heritarum;
NUM|26|17|Arodi, ab hoc familia Aroditarum; Areli, ab hoc familia Arelitarum.
NUM|26|18|Istae sunt familiae Gad, quarum omnis numerus fuit quadraginta milia quingenti.
NUM|26|19|Filii Iudae Her et Onan, qui ambo mortui sunt in terra Chanaan.
NUM|26|20|Fueruntque filii Iudae per cognationes suas: Sela, a quo familia Selanitarum; Phares, a quo familia Pharesitarum; Zara, a quo familia Zaraitarum.
NUM|26|21|Porro filii Phares: Esrom, a quo familia Esromitarum; et Hamul, a quo familia Hamulitarum.
NUM|26|22|Istae sunt familiae Iudae, quarum omnis numerus fuit septuaginta sex milia quingenti.
NUM|26|23|Filii Issachar per cognationes suas: Thola, a quo familia Tholaitarum; Phua, a quo familia Phuaitarum;
NUM|26|24|Iasub, a quo familia Iasubitarum; Semron, a quo familia Semronitarum.
NUM|26|25|Hae sunt cognationes Issachar, quarum numerus fuit sexaginta quattuor milia trecenti.
NUM|26|26|Filii Zabulon per cognationes suas: Sared, a quo familia Sareditarum; Elon, a quo familia Elonitarum; Iahelel, a quo familia Iahelelitarum.
NUM|26|27|Hae sunt cognationes Zabulon, quarum numerus fuit sexaginta milia quingenti.
NUM|26|28|Filii Ioseph per cognationes suas: Manasse et Ephraim.
NUM|26|29|De Manasse ortus est Machir, a quo familia Machiritarum; Machir genuit Galaad, a quo familia Galaaditarum.
NUM|26|30|Galaad habuit filios: Iezer, a quo familia Iezeritarum; et Helec, a quo familia Helecitarum;
NUM|26|31|et Asriel, a quo familia Asrielitarum; et Sechem, a quo familia Sechemitarum;
NUM|26|32|et Semida, a quo familia Semidaitarum; et Hepher, a quo familia Hepheritarum.
NUM|26|33|Fuit autem Hepher pater Salphaad, qui filios non habebat sed tantum filias, quarum ista sunt nomina: Maala et Noa et Hegla et Melcha et Thersa.
NUM|26|34|Hae sunt familiae Manasse, et numerus earum quinquaginta duo milia septingenti.
NUM|26|35|Filii autem Ephraim per cognationes suas fuerunt hi: Suthala, a quo familia Suthalaitarum; Becher, a quo familia Becheritarum; Thehen, a quo familia Thehenitarum.
NUM|26|36|Porro filius Suthala fuit Heran, a quo familia Heranitarum.
NUM|26|37|Hae sunt cognationes filiorum Ephraim, quarum numerus fuit triginta duo milia quingenti. Isti sunt filii Ioseph per familias suas.
NUM|26|38|Filii Beniamin in cognationibus suis: Bela, a quo familia Belaitarum; Asbel, a quo familia Asbelitarum; Ahiram, a quo familia Ahiramitarum;
NUM|26|39|Supham, a quo familia Suphamitarum; Hupham, a quo familia Huphamitarum.
NUM|26|40|Filii Bela: Ared et Naaman; de Ared familia Areditarum, de Naaman familia Naamanitarum.
NUM|26|41|Hi sunt filii Beniamin per cognationes suas, quorum numerus fuit quadraginta quinque milia sescenti.
NUM|26|42|Filii Dan per cognationes suas: Suham, a quo familia Suhamitarum. Hae sunt cognationes Dan per familias suas:
NUM|26|43|omnes fuere Suhamitae, quorum numerus erat sexaginta quattuor milia quadringenti.
NUM|26|44|Filii Aser per cognationes suas: Iemna, a quo familia Iemnaitarum; Isui, a quo familia Isuitarum; Beria, a quo familia Beriaitarum.
NUM|26|45|Filii Beria: Heber, a quo familia Heberitarum, et Melchiel a quo familia Melchielitarum.
NUM|26|46|Nomen autem filiae Aser fuit Sara.
NUM|26|47|Hae cognationes filiorum Aser, et numerus eorum quinquaginta tria milia quadringenti.
NUM|26|48|Filii Nephthali per cognationes suas: Iasiel, a quo familia Iasielitarum; Guni, a quo familia Gunitarum;
NUM|26|49|Ieser, a quo familia Ieseritarum; Sellem, a quo familia Sellemitarum.
NUM|26|50|Hae sunt cognationes filiorum Nephthali per familias suas, quorum numerus quadraginta quinque milia quadringenti.
NUM|26|51|Ista est summa filiorum Israel qui recensiti sunt: sescenta milia et mille septingenti triginta.
NUM|26|52|Locutusque est Dominus ad Moysen dicens:
NUM|26|53|" Istis dividetur terra iuxta numerum vocabulorum in possessiones suas.
NUM|26|54|Pluribus maiorem partem dabis et paucioribus minorem: singulis, sicut nunc recensiti sunt, tradetur possessio;
NUM|26|55|ita dumtaxat, ut sors terram dividat. Secundum numerum tribuum patrum suorum hereditabunt.
NUM|26|56|Quidquid sorte contigerit, hoc vel plures accipiant vel pauciores.
NUM|26|57|Hic quoque est numerus filiorum Levi per familias suas: Gerson, a quo familia Gersonitarum; Caath, a quo familia Caathitarum; Merari, a quo familia Meraritarum.
NUM|26|58|Hae sunt familiae Levi: familia Lobni, familia Hebroni, familia Moholi, familia Musi, familia Core. At vero Caath genuit Amram,
NUM|26|59|qui habuit uxorem Iochabed filiam Levi, quae nata est ei in Aegypto. Haec genuit Amram viro suo filios, Aaron et Moysen et Mariam sororem eorum.
NUM|26|60|De Aaron orti sunt Nadab et Abiu et Eleazar et Ithamar,
NUM|26|61|quorum Nadab et Abiu mortui sunt, cum obtulissent ignem alienum coram Domino.
NUM|26|62|Fueruntque omnes, qui numerati sunt, viginti tria milia generis masculini ab uno mense et supra; quia non sunt recensiti inter filios Israel, nec eis cum ceteris data possessio est.
NUM|26|63|Hic est numerus filiorum Israel, qui descripti sunt a Moyse et Eleazaro sacerdote in campestribus Moab supra Iordanem contra Iericho;
NUM|26|64|inter quos nullus fuit eorum, qui ante numerati sunt a Moyse et Aaron in deserto Sinai:
NUM|26|65|praedixerat enim Dominus quod omnes morerentur in solitudine; nullusque remansit ex eis, nisi Chaleb filius Iephonne et Iosue filius Nun.
NUM|27|1|Accesserunt autem filiae Sal phaad filii Hepher filii Ga laad filii Machir filii Manasse, e cognationibus Manasse, qui fuit filius Ioseph, quarum sunt nomina: Maala et Noa et Hegla et Melcha et Thersa.
NUM|27|2|Steteruntque coram Moyse et Eleazaro sacerdote et principibus et cuncta congregatione ad ostium tabernaculi conventus atque dixerunt:
NUM|27|3|" Pater noster mortuus est in deserto, nec fuit in seditione, quae concitata est contra Dominum sub Core, sed in peccato suo mortuus est; hic non habuit mares filios.
NUM|27|4|Cur tollitur nomen illius de familia sua, quia non habuit filium? Date nobis possessionem inter fratres patris nostri ".
NUM|27|5|Rettulitque Moyses causam earum ad iudicium Domini,
NUM|27|6|qui dixit ad eum:
NUM|27|7|" Iustam rem postulant filiae Salphaad. Da eis possessionem inter fratres patris sui, et ei in hereditatem succedant.
NUM|27|8|Ad filios autem Israel loqueris haec: Homo cum mortuus fuerit absque filio, ad filiam eius transibit hereditas;
NUM|27|9|si filiam non habuerit, habebit successores fratres suos.
NUM|27|10|Quod si et fratres non fuerint, dabitis hereditatem fratribus patris eius.
NUM|27|11|Sin autem nec patruos habuerit, dabitur hereditas illi, qui ei proximus est e cognatione sua; possidebitque eam. Eritque hoc filiis Israel sanctum lege perpetua, sicut praecepit Dominus Moysi ".
NUM|27|12|Dixit quoque Dominus ad Moysen: " Ascende in montem istum Abarim et contemplare inde terram, quam daturus sum filiis Israel.
NUM|27|13|Cumque videris eam, ibis et tu ad populum tuum, sicut ivit frater tuus Aaron,
NUM|27|14|quia offendistis me in deserto Sin in contradictione congregationis, nec sanctificare me voluistis coram ea super aquas ". Hae sunt aquae Meribathcades deserti Sin.
NUM|27|15|Cui respondit Moyses:
NUM|27|16|" Provideat Dominus, Deus spirituum omnis carnis, hominem, qui sit super congregationem hanc
NUM|27|17|et possit exire et intrare ante eos et educere eos vel introducere, ne sit populus Domini sicut oves absque pastore ".
NUM|27|18|Dixitque Dominus ad eum: " Tolle Iosue filium Nun, virum in quo est spiritus; et pone manum tuam super eum,
NUM|27|19|quem statues coram Eleazaro sacerdote et omni congregatione et dabis ei praecepta, cunctis videntibus,
NUM|27|20|et partem gloriae tuae, ut audiat eum omnis synagoga filiorum Israel.
NUM|27|21|Stabit coram Eleazaro sacerdote, qui pro eo iudicium Urim consulet Dominum. Ad verbum eius egredietur et ingredietur ipse et omnes filii Israel cum eo, cuncta congregatio ".
NUM|27|22|Fecit Moyses, ut praeceperat Dominus. Cumque tulisset Iosue, statuit eum coram Eleazaro sacerdote et omni frequentia populi;
NUM|27|23|et, impositis capiti eius manibus, constituit eum, sicut mandaverat Dominus per manum Moysi.
NUM|28|1|Dixit quoque Dominus ad Moysen:
NUM|28|2|" Praecipe filiis Is rael et dices ad eos: Oblationem meam et panem meum, sacrificium ignis in odorem suavissimum offerte per tempora sua.
NUM|28|3|Hoc est sacrificium ignis, quod offerre debetis: agnos anniculos immaculatos duos cotidie in holocaustum sempiternum;
NUM|28|4|unum offeretis mane et alterum ad vesperam;
NUM|28|5|decimam partem ephi similae in oblationem, quae conspersa sit oleo purissimo et habeat quartam partem hin.
NUM|28|6|Holocaustum iuge est, quod obtulistis in monte Sinai in odorem suavissimum, sacrificium ignis Domino;
NUM|28|7|et libabitis vini quartam partem hin per agnos singulos; in sanctuario effundetis libamen potus inebriantis Domino.
NUM|28|8|Alterumque agnum similiter offeretis ad vesperam, iuxta ritum sacrificii matutini: sacrificium ignis in odorem suavissimum Domino.
NUM|28|9|Die autem sabbati offeretis duos agnos anniculos immaculatos et duas decimas similae oleo conspersae et libamentum eius.
NUM|28|10|Est holocaustum sabbati per singula sabbata, praeter holocaustum sempiternum et libamentum eius.
NUM|28|11|In calendis autem offeretis holocaustum Domino vitulos de armento duos, arietem unum, agnos anniculos septem immaculatos
NUM|28|12|et tres decimas similae oleo conspersae in oblatione per singulos vitulos et duas decimas similae oleo conspersae per singulos arietes,
NUM|28|13|et decimam unam similae oleo conspersae in oblatione per agnos singulos: holocaustum in odorem suavissimum, sacrificium ignis Domino.
NUM|28|14|Libamenta autem eorum ista erunt: media pars hin vini per singulos vitulos, tertia per arietem, quarta per agnum. Hoc erit holocaustum per omnes menses, qui sibi anno vertente succedunt.
NUM|28|15|Hircus quoque offeretur Domino pro peccato, praeter holocaustum sempiternum cum libamentis suis.
NUM|28|16|Mense autem primo, quarta decima die mensis Pascha Domini erit,
NUM|28|17|et quinta decima die sollemnitas. Septem diebus vescemini azymis,
NUM|28|18|quarum die prima conventus sanctus erit; omne opus servile non facietis in ea.
NUM|28|19|Offeretisque sacrificium ignis, holocaustum Domino: vitulos de armento duos, arietem unum, agnos anniculos immaculatos septem;
NUM|28|20|et oblationem singulorum ex simila, quae conspersa sit oleo, tres decimas per singulos vitulos et duas decimas per arietem
NUM|28|21|et decimam unam per agnos singulos, id est per septem agnos;
NUM|28|22|et hircum pro peccato unum, ut expietur pro vobis,
NUM|28|23|praeter holocaustum matutinum, quod semper offeretis.
NUM|28|24|Ita facietis per singulos dies septem dierum: panem, sacrificium ignis in odorem suavissimum Domino praeter holocaustum iuge et libationem eius.
NUM|28|25|Die quoque septimo conventus sanctus erit vobis; omne opus servile non facietis in eo.
NUM|28|26|Die etiam primitivorum, quando offeretis oblationem novam Domino, in sollemnitate Hebdomadarum, conventus sanctus erit vobis; omne opus servile non facietis in ea.
NUM|28|27|Offeretisque holocaustum in odorem suavissimum Domino: vitulos de armento duos, arietem unum et agnos anniculos immaculatos septem,
NUM|28|28|atque in oblatione eorum similae oleo conspersae, tres decimas per singulos vitulos, per arietem duas,
NUM|28|29|per agnos decimam unam, qui simul sunt agni septem;
NUM|28|30|hircum quoque, qui mactatur pro expiatione,
NUM|28|31|praeter holocaustum sempiternum et oblationem eius. Immaculata offeretis omnia cum libationibus suis.
NUM|29|1|Mensis etiam septimi prima die conventus sanctus erit vo bis; omne opus servile non facietis in ea, quia dies clangoris est et tubarum.
NUM|29|2|Offeretisque holocaustum in odorem suavissimum Domino: vitulum de armento unum, arietem unum et agnos anniculos immaculatos septem;
NUM|29|3|et in oblationibus eorum similae oleo conspersae tres decimas per vitulum, duas decimas per arietem,
NUM|29|4|unam decimam per agnum, qui simul sunt agni septem;
NUM|29|5|et hircum pro peccato, qui offertur in expiationem vestram,
NUM|29|6|praeter holocaustum calendarum cum oblatione et holocaustum sempiternum cum oblatione et libationibus solitis in odorem suavissimum, sacrificium ignis Domino.
NUM|29|7|Decima quoque die mensis huius septimi erit vobis conventus sanctus, et affligetis animas vestras; omne opus servile non facietis.
NUM|29|8|Offeretisque holocaustum Domino in odorem suavissimum: vitulum de armento unum, arietem unum, agnos anniculos immaculatos septem;
NUM|29|9|et in oblatione eorum similae oleo conspersae tres decimas per vitulum, duas decimas per arietem,
NUM|29|10|decimam unam per agnos singulos, qui sunt simul septem agni;
NUM|29|11|et hircum pro peccato, absque his, quae offerri pro delicto solent in expiationem et holocaustum sempiternum cum oblatione et libaminibus eorum.
NUM|29|12|Quinta decima vero die mensis septimi conventus sanctus erit; omne opus servile non facietis in ea, sed celebrabitis sollemnitatem Domino septem diebus
NUM|29|13|offeretisque holocaustum in odorem suavissimum Domino: vitulos de armento tredecim, arietes duos, agnos anniculos immaculatos quattuordecim;
NUM|29|14|et in oblatione eorum similae oleo conspersae tres decimas per vitulos singulos, qui sunt simul vituli tredecim, et duas decimas arieti uno, id est simul arietibus duobus,
NUM|29|15|et decimam unam agnis singulis, qui sunt simul agni quattuordecim;
NUM|29|16|et hircum pro peccato absque holocausto sempiterno et oblatione et libamine eius.
NUM|29|17|In die altero offeretis vitulos de armento duodecim, arietes duos, agnos anniculos immaculatos quattuordecim;
NUM|29|18|oblationemque et libamina singulorum per vitulos et arietes et agnos iuxta numerum eorum rite celebrabitis,
NUM|29|19|et hircum pro peccato absque holocausto sempiterno oblationeque et libamine eorum.
NUM|29|20|Die tertio offeretis vitulos undecim, arietes duos, agnos anniculos imma culatos quattuordecim,
NUM|29|21|oblationem et libamina singulorum per vitulos et arietes et agnos iuxta numerum eorum rite celebrabitis,
NUM|29|22|et hircum pro peccato absque holocausto sempiterno oblationeque et libamine eius.
NUM|29|23|Die quarto offeretis vitulos decem, arietes duos, agnos anniculos immaculatos quattuordecim,
NUM|29|24|oblationem et libamina singulorum per vitulos et arietes et agnos iuxta numerum eorum rite celebrabitis,
NUM|29|25|et hircum pro peccato absque holocausto sempiterno, oblatione eius et libamine.
NUM|29|26|Die quinto offeretis vitulos novem, arietes duos, agnos anniculos immaculatos quattuordecim,
NUM|29|27|oblationem et libamina singulorum per vitulos et arietes et agnos iuxta numerum eorum rite celebrabitis,
NUM|29|28|et hircum pro peccato absque holocausto sempiterno, oblatione eius et libamine.
NUM|29|29|Die sexto offeretis vitulos octo, arietes duos, agnos anniculos immaculatos quattuordecim,
NUM|29|30|oblationem et libamina singulorum per vitulos et arietes et agnos iuxta numerum eorum rite celebrabitis,
NUM|29|31|et hircum pro peccato absque holocausto sempiterno, oblatione eius et libamine.
NUM|29|32|Die septimo offeretis vitulos septem et arietes duos, agnos anniculos immaculatos quattuordecim,
NUM|29|33|oblationem et libamina singulorum per vitulos et arietes et agnos iuxta numerum eorum rite celebrabitis,
NUM|29|34|et hircum pro peccato absque holocausto sempiterno, oblatione eius et libamine.
NUM|29|35|Die octavo erit conventus sollemnis, omne opus servile non facietis
NUM|29|36|offerentes holocaustum in odorem suavissimum Domino: vitulum unum, arietem unum, agnos anniculos immaculatos septem,
NUM|29|37|oblationem et libamina singulorum per vitulum et arietem et agnos iuxta numerum eorum rite celebrabitis,
NUM|29|38|et hircum pro peccato absque holocausto sempiterno, oblatione eius et libamine.
NUM|29|39|Haec offeretis Domino in sollemnitatibus vestris, praeter vota et oblationes spontaneas in holocaustis, in oblationibus, in libaminibus et in hostiis pacificis ".
NUM|30|1|Narravitque Moyses filiis Israel omnia, quae ei Dominus imperarat,
NUM|30|2|et locutus est ad principes tribuum filiorum Israel: " Iste est sermo, quem praecepit Dominus:
NUM|30|3|Si quis virorum votum Domino voverit aut se constrinxerit iuramento, non faciet irritum verbum suum, sed omne, quod promisit, implebit.
NUM|30|4|Mulier, si quippiam voverit Domino aut se constrinxerit iuramento, quae est in domo patris sui et in aetate adhuc puellari,
NUM|30|5|si cognoverit pater votum, quod pollicita est, aut iuramentum, quo ligavit animam suam, et tacuerit, voti rea erit; quidquid pollicita est aut iuravit, opere complebit.
NUM|30|6|Sin autem, quo die audierit contradixerit pater, et vota et iuramenta eius irrita erunt; et propitius erit ei Dominus, eo quod contradixerit pater.
NUM|30|7|Si maritum habuerit et voverit aliquid, aut semel de ore eius verbum egrediens animam eius ligaverit iuramento,
NUM|30|8|quo die audierit vir eius et non contradixerit, voti rea erit reddetque, quodcumque promiserat.
NUM|30|9|Sin autem, quo die audierit contradixerit, irritas facit pollicitationes eius verbaque, quibus obstrinxerat animam suam; et propitius erit ei Dominus.
NUM|30|10|Vidua et repudiata, quidquid voverint, reddent.
NUM|30|11|Uxor in domo viri cum se voto constrinxerit aut iuramento,
NUM|30|12|si audierit vir et tacuerit nec contradixerit sponsioni, reddet, quodcumque promiserat.
NUM|30|13|Sin autem extemplo contradixerit, non tenebitur promissionis rea, quia maritus contradixit, et Dominus ei propitius erit.
NUM|30|14|Si voverit aut iuramento se constrinxerit, ut per ieiunium affligat animam suam, in arbitrio viri erit, ut faciat sive non faciat.
NUM|30|15|Quod si audiens vir tacuerit et de die in diem distulerit sententiam, quidquid voverat atque promiserat, reddet, quia, quo die audierat, tacuit.
NUM|30|16|Sin autem contradixerit, postquam rescivit, portabit ipse iniquitatem eius ".
NUM|30|17|Istae sunt leges, quas constituit Dominus Moysi inter virum et uxorem, inter patrem et filiam, quae in puellari adhuc aetate manet in parentis domo.
NUM|31|1|Locutusque est Dominus ad Moysen dicens:
NUM|31|2|" Ulciscere filios Israel de Madianitis et sic colligeris ad populum tuum ".
NUM|31|3|Statimque Moyses: " Armate, inquit, ex vobis viros ad pugnam, qui possint ultionem Domini expetere de Madianitis.
NUM|31|4|Mille viri de singulis tribubus eligantur ex Israel, qui mittantur ad bellum ".
NUM|31|5|Dederuntque millenos de singulis tribubus, id est duodecim milia expeditorum ad pugnam,
NUM|31|6|quos misit Moyses cum Phinees filio Eleazari sacerdotis. Vasa quoque sancta et tubas ad clangendum tradidit ei.
NUM|31|7|Cumque pugnassent contra Madianitas, sicut praeceperat Dominus Moysi, omnes mares occiderunt
NUM|31|8|et reges eorum Evi et Recem et Sur et Hur et Rebe, quinque principes gentis, Balaam quoque filium Beor interfecerunt gladio;
NUM|31|9|ceperuntque mulieres eorum et parvulos. Omniaque pecora et cunctam supellectilem, quidquid habere potuerant, depopulati sunt:
NUM|31|10|tam urbes quam viculos et castra flamma consumpsit;
NUM|31|11|et tulerunt praedam et universa, quae ceperant, tam ex hominibus quam ex iumentis,
NUM|31|12|et adduxerunt captivos, spolia et praedam ad Moysen et Eleazarum sacerdotem et ad omnem congregationem filiorum Israel ad castra in campestribus Moab iuxta Iordanem contra Iericho.
NUM|31|13|Egressi sunt autem Moyses et Eleazar sacerdos et omnes principes synagogae in occursum eorum extra castra.
NUM|31|14|Iratusque Moyses principibus exercitus, tribunis et centurionibus, qui venerant de bello,
NUM|31|15|ait: " Cur omnes feminas reservastis?
NUM|31|16|Nonne istae sunt, quae deceperunt filios Israel ad suggestionem Balaam et praevaricari vos fecerunt in Dominum super peccato Phegor, unde et percussus est populus Domini?
NUM|31|17|Ergo cunctos interficite parvulos generis masculini et omnes mulieres, quae noverunt viros in coitu, iugulate;
NUM|31|18|puellas autem et omnes feminas virgines reservate vobis.
NUM|31|19|Et vos manete extra castra septem diebus; qui occiderit hominem vel occisum tetigerit, lustrabitur die tertio et septimo, vos et captivi vestri.
NUM|31|20|Et de omni praeda, sive vestimentum fuerit sive aliquid in utensilia praeparatum de caprarum pellibus et pilis et ligno, lustrabitis ".
NUM|31|21|Eleazar quoque sacerdos ad viros exercitus, qui pugnaverant, sic locutus est: " Hoc est praeceptum legis, quod mandavit Dominus Moysi:
NUM|31|22|Aurum et argentum et aes et ferrum et stannum et plumbum,
NUM|31|23|omne, quod potest transire per flammas, igne purgabitur; quidquid autem ignem non potest sustinere, aqua expiationis sanctificabitur.
NUM|31|24|Et lavabitis vestimenta vestra die septimo, et purificati postea castra intrabitis ".
NUM|31|25|Dixit quoque Dominus ad Moysen:
NUM|31|26|" Tollite summam eorum, quae capta sunt, ab homine usque ad pecus, tu et Eleazar sacerdos et principes familiarum;
NUM|31|27|dividesque ex aequo praedam inter eos, qui pugnaverunt egressique sunt ad bellum, et inter omnem congregationem.
NUM|31|28|Et separabis partem Domino ab his, qui pugnaverunt et fuerunt in bello, unam animam de quingentis tam ex hominibus quam ex bobus et asinis et ovibus
NUM|31|29|et dabis eam Eleazaro sacerdoti, quia praelibatio Domini sunt.
NUM|31|30|Ex media quoque parte filiorum Israel accipies quinquagesimum caput hominum et boum et asinorum et ovium cunctorum animantium et dabis ea Levitis, qui excubant in custodiis habitaculi Domini ".
NUM|31|31|Feceruntque Moyses et Eleazar sacerdos, sicut praeceperat Dominus.
NUM|31|32|Fuit autem praeda, quae supererat, quam exercitus ceperat, ovium sescenta septuaginta quinque milia,
NUM|31|33|boum septuaginta duo milia,
NUM|31|34|asinorum sexaginta milia et mille,
NUM|31|35|animae hominum sexus feminei, quae non cognoverant viros, triginta duo milia.
NUM|31|36|Dataque est media pars his, qui in proelio fuerant, ovium trecenta triginta septem milia quingentae,
NUM|31|37|e quibus in partem Domini supputatae sunt oves sescentae septuaginta quinque,
NUM|31|38|et de bobus triginta sex milibus, boves septuaginta et duo,
NUM|31|39|de asinis triginta milibus quingentis, asini sexaginta unus,
NUM|31|40|de animabus hominum sedecim milibus, cesserunt in partem Domini triginta duae animae.
NUM|31|41|Tradiditque Moyses tributum praelibationis Domini Eleazaro sacerdoti, sicut fuerat ei imperatum.
NUM|31|42|Ex media vero parte filiorum Israel, quam separaverat a parte eorum, qui in proelio fuerant,
NUM|31|43|de hac media parte, quae contigerat congregationi, id est de ovibus trecentis triginta septem milibus quingentis
NUM|31|44|et de bobus triginta sex milibus
NUM|31|45|et de asinis triginta milibus quingentis
NUM|31|46|et de hominibus sedecim milibus,
NUM|31|47|tulit Moyses quinquagesimum caput et dedit Levitis, qui excubabant in habitaculo Domini, sicut praeceperat Dominus.
NUM|31|48|Cumque accessissent principes exercitus ad Moysen, tribuni centurionesque, dixerunt:
NUM|31|49|" Nos servi tui recensuimus numerum pugnatorum, quos habuimus sub manu nostra, et ne unus quidem defuit.
NUM|31|50|Ob hanc causam offerimus in donariis Domini singuli, quod auri potuimus invenire, periscelidas et armillas, anulos et inaures ac muraenulas, ad placandum pro nobis Dominum ".
NUM|31|51|Susceperuntque Moyses et Eleazar sacerdos aurum in diversis speciebus;
NUM|31|52|omne aurum, quod elevaverunt Domino, pondo sedecim milia septingentos quinquaginta siclos, a tribunis et centurionibus.
NUM|31|53|Unusquisque enim, quod in praeda rapuerat, suum erat.
NUM|31|54|Et susceptum intulerunt in tabernaculum conventus in monumentum filiorum Israel coram Domino.
NUM|32|1|Filii autem Ruben et Gad habebant pecora multa, et erat illis in iumentis infinita substantia. Cumque vidissent Iazer et Galaad aptas animalibus alendis terras,
NUM|32|2|venerunt ad Moysen et ad Eleazarum sacerdotem et principes congregationis atque dixerunt:
NUM|32|3|" Ataroth et Dibon et Iazer et Nemra, Hesebon et Eleale et Sabam et Nabo et Beon,
NUM|32|4|terra, quam percussit Dominus in conspectu congregationis Israel, regio uberrima est ad pastum animalium, et nos servi tui habemus iumenta plurima ".
NUM|32|5|Dixeruntque: " Si invenimus gratiam coram te, detur haec terra famulis tuis in possessionem, nec facias nos transire Iordanem ".
NUM|32|6|Quibus respondit Moyses: " Numquid fratres vestri ibunt ad pugnam, et vos hic sedebitis?
NUM|32|7|Cur subvertitis mentes filiorum Israel, ne transire audeant in terram, quam eis daturus est Dominus?
NUM|32|8|Nonne ita egerunt patres vestri, quando misi de Cadesbarne ad explorandam terram?
NUM|32|9|Cumque venissent usque ad Nehelescol, lustrata omni regione, subverterunt cor filiorum Israel, ut non intrarent terram, quam eis Dominus dedit.
NUM|32|10|Qui iratus iuravit dicens:
NUM|32|11|"Non videbunt homines isti, qui ascenderunt ex Aegypto, a viginti annis et supra, terram, quam sub iuramento pollicitus sum Abraham, Isaac et Iacob; nam noluerunt sequi me,
NUM|32|12|praeter Chaleb filium Iephonne Cenezaeum et Iosue filium Nun: isti secuti sunt Dominum!".
NUM|32|13|Iratusque Dominus adversum Israel circumduxit eum per desertum quadraginta annis, donec consumeretur universa generatio, quae fecerat malum in conspectu eius.
NUM|32|14|Et ecce, inquit, vos surrexistis pro patribus vestris progenies hominum peccatorum, ut augeretis furorem irae Domini contra Israel.
NUM|32|15|Quod si nolueritis sequi eum, in solitudine iterum populum hunc circumducet, et vos causa eritis necis omnium ".
NUM|32|16|At illi prope accedentes dixerunt: " Caulas ovium fabricabimus pro iumentis nostris, parvulis quoque nostris urbes;
NUM|32|17|nos autem ipsi armati et accincti pergemus ad proelium ante filios Israel, donec introducamus eos ad loca sua. Parvuli nostri erunt in urbibus muratis propter habitatorum insidias.
NUM|32|18|Non revertemur in domos nostras usque dum possideant filii Israel hereditatem suam;
NUM|32|19|nec quidquam quaeremus trans Iordanem et ultra, quia iam habemus nostram hereditatem in orientali eius plaga ".
NUM|32|20|Quibus Moyses ait: " Si feceritis quod promittitis, si expediti perrexeritis coram Domino ad pugnam,
NUM|32|21|et omnis vir bellator armatus Iordanem transierit, donec expulerit Dominus inimicos suos ante se,
NUM|32|22|et subiecta ei omni terra redieritis in terram hanc, tunc eritis inculpabiles apud Dominum et apud Israel et obtinebitis terram hanc in hereditatem coram Domino.
NUM|32|23|Sin autem, quod dicitis, non feceritis, nulli dubium est quin peccetis in Dominum; et scitote quoniam peccatum vestrum apprehendet vos.
NUM|32|24|Aedificate ergo urbes parvulis vestris et caulas ovibus et, quod polliciti estis, implete ".
NUM|32|25|Dixeruntque filii Gad et Ruben ad Moysen: " Servi tui sumus, faciemus, quod iubet dominus noster:
NUM|32|26|parvulos nostros, mulieres, pecora ac iumenta remanebunt ibi in urbibus Galaad;
NUM|32|27|famuli autem tui, omnes expediti pergent coram Domino ad bellum, sicut tu, domine, loqueris ".
NUM|32|28|Praecepit ergo Moyses Eleazaro sacerdoti et Iosue filio Nun et principibus familiarum per tribus filiorum Israel et dixit ad eos:
NUM|32|29|" Si transierint filii Gad et filii Ruben vobiscum Iordanem omnes armati ad bellum coram Domino, et vobis fuerit terra subiecta, date eis Galaad in possessionem.
NUM|32|30|Sin autem noluerint transire armati vobiscum in terram Chanaan, inter vos habitandi accipiant loca ".
NUM|32|31|Responderuntque filii Gad et filii Ruben: " Sicut locutus est Dominus servis suis, ita faciemus.
NUM|32|32|Ipsi armati pergemus coram Domino in terram Chanaan; et possidebimus hereditatem nostram trans Iordanem ".
NUM|32|33|Dedit itaque Moyses filiis Gad et Ruben et dimidiae tribui Manasse filii Ioseph regnum Sehon regis Amorraei et regnum Og regis Basan, terram cum urbibus suis et terminis, urbes terrae per circuitum.
NUM|32|34|Igitur exstruxerunt filii Gad Dibon et Ataroth et Aroer
NUM|32|35|et Atrothsophan et Iazer et Iegbaa
NUM|32|36|et Bethnemra et Betharan, urbes munitas, et caulas pecoribus suis.
NUM|32|37|Filii vero Ruben aedificaverunt Hesebon et Eleale et Cariathaim
NUM|32|38|et Nabo et Baalmeon, versis nominibus, Sabama quoque, imponentes vocabula urbibus, quas exstruxerant.
NUM|32|39|Porro filii Machir filii Manasse perrexerunt in Galaad et ceperunt eam, expulso Amorraeo habitatore eius.
NUM|32|40|Dedit ergo Moyses terram Galaad Machir filio Manasse, qui habitavit in ea.
NUM|32|41|Iair autem filius Manasse abiit et occupavit vicos eius, quos appellavit Havoth Iair (id est villas Iair).
NUM|32|42|Nobe quoque perrexit et apprehendit Canath cum viculis suis vocavitque eam ex nomine suo Nobe.
NUM|33|1|Hae sunt mansiones filiorum Israel, qui egressi sunt de Ae gypto per turmas suas in manu Moysi et Aaron,
NUM|33|2|quas descripsit Moyses iuxta castrorum loca, quae Domini iussione mutabant.
NUM|33|3|Profecti igitur de Ramesse mense primo, quinta decima die mensis primi, altera die Paschae, filii Israel in manu excelsa, videntibus cunctis Aegyptiis
NUM|33|4|et sepelientibus primogenitos, quos percusserat Dominus, nam et in diis eorum exercuerat ultionem,
NUM|33|5|castrametati sunt in Succoth.
NUM|33|6|Et de Succoth venerunt in Etham, quae est in extremis finibus solitudinis.
NUM|33|7|Inde egressi venerunt contra Phihahiroth, quae respicit Beelsephon, et castrametati sunt ante Magdolum.
NUM|33|8|Profectique de Phihahiroth transierunt per medium mare in solitudinem, et ambulantes tribus diebus per desertum Etham castrametati sunt in Mara.
NUM|33|9|Profectique de Mara venerunt in Elim, ubi erant duodecim fontes aquarum et palmae septuaginta; ibique castrametati sunt.
NUM|33|10|Sed et inde egressi fixerunt tentoria super mare Rubrum. Profectique de mari Rubro
NUM|33|11|castrametati sunt in deserto Sin;
NUM|33|12|unde egressi venerunt in Daphca.
NUM|33|13|Profectique de Daphca castrametati sunt in Alus.
NUM|33|14|Egressique de Alus in Raphidim fixere tentoria, ubi populo defuit aqua ad bibendum;
NUM|33|15|profectique de Raphidim castrametati sunt in deserto Sinai.
NUM|33|16|Sed et de solitudine Sinai egressi venerunt ad Cibrottaava;
NUM|33|17|profectique de Cibrottaava castrametati sunt in Aseroth.
NUM|33|18|Et de Aseroth venerunt in Rethma;
NUM|33|19|profectique de Rethma castrametati sunt in Remmonphares.
NUM|33|20|Unde egressi venerunt in Lebna;
NUM|33|21|de Lebna castrametati sunt in Ressa;
NUM|33|22|egressique de Ressa venerunt in Ceelatha,
NUM|33|23|unde profecti castrametati sunt in monte Sepher.
NUM|33|24|Egressi de monte Sepher venerunt in Arada;
NUM|33|25|inde proficiscentes castrametati sunt in Maceloth;
NUM|33|26|profectique de Maceloth venerunt in Thahath;
NUM|33|27|de Thahath castrametati sunt in Thare.
NUM|33|28|Unde egressi fixere tentoria in Methca
NUM|33|29|et de Methca castrametati sunt in Hesmona;
NUM|33|30|profectique de Hesmona venerunt in Moseroth.
NUM|33|31|Et de Moseroth castrametati sunt in Beneiacan;
NUM|33|32|profectique de Beneiacan venerunt in montem Gadgad;
NUM|33|33|unde profecti castrametati sunt in Ietebatha.
NUM|33|34|Et de Ietebatha venerunt in Ebrona;
NUM|33|35|egressique de Ebrona castrametati sunt in Asiongaber.
NUM|33|36|Inde profecti venerunt in desertum Sin, hoc est Cades.
NUM|33|37|Egressique de Cades castrametati sunt in monte Hor in extremis finibus terrae Edom.
NUM|33|38|Ascenditque Aaron sacerdos in montem Hor, iubente Domino, et ibi mortuus est anno quadragesimo egressionis filiorum Israel ex Aegypto, mense quinto, prima die mensis,
NUM|33|39|cum esset annorum centum viginti trium.
NUM|33|40|Audivitque Chananaeus rex Arad, qui habitabat in Nageb, in terra Chanaan, venisse filios Israel.
NUM|33|41|Et profecti de monte Hor castrametati sunt in Salmona;
NUM|33|42|unde egressi venerunt in Phinon.
NUM|33|43|Profectique de Phinon castrametati sunt in Oboth;
NUM|33|44|et de Oboth venerunt in Ieabarim, quae est in finibus Moabitarum.
NUM|33|45|Profectique de Ieabarim fixere tentoria in Dibongad;
NUM|33|46|unde egressi castrametati sunt in Elmondeblathaim.
NUM|33|47|Egressique de Elmondeblathaim venerunt ad montes Abarim contra Nabo.
NUM|33|48|Profectique de montibus Abarim transierunt ad campestria Moab supra Iordanem contra Iericho;
NUM|33|49|ibique castrametati sunt de Bethiesimoth usque ad Abelsettim in campestribus Moab.
NUM|33|50|Ubi locutus est Dominus ad Moysen:
NUM|33|51|" Praecipe filiis Israel et dic ad eos: Quando transieritis Iordanem intrantes terram Chanaan,
NUM|33|52|disperdite cunctos habitatores terrae ante vos, confringite omnes imagines eorum et omnes statuas comminuite atque omnia excelsa vastate.
NUM|33|53|Possidebitis terram et habitabitis in ea. Ego enim dedi vobis illam in possessionem,
NUM|33|54|quam dividetis inter tribus vestras. Maiori dabitis latiorem et minori angustiorem; singulis, ut sors ceciderit, ita tribuetur hereditas; per tribus et familias possessio dividetur.
NUM|33|55|Sin autem nolueritis expellere habitatores terrae, qui remanserint, erunt vobis quasi spinae in oculis vestris et sudes in lateribus, et adversabuntur vobis in terra habitationis vestrae;
NUM|33|56|et, quidquid illis cogitaveram facere, vobis faciam ".
NUM|34|1|Locutusque est Dominus ad Moysen dicens:
NUM|34|2|" Praecipe fi liis Israel et dices ad eos: Cum ingressi fueritis terram hanc Chanaan, et in possessionem vobis sorte ceciderit, his finibus terminabitur.
NUM|34|3|Pars meridiana incipiet a solitudine Sin, quae est iuxta Edom, et habebit terminos contra orientem mare Salsissimum.
NUM|34|4|Qui circuibunt australem plagam per ascensum Acrabbim (id est Scorpionum), ita ut transeant in Sin et perveniant ad meridiem Cadesbarne, unde egredientur ad Asaraddar et tendent usque ad Asemona.
NUM|34|5|Ibitque per gyrum terminus ab Asemona usque ad torrentem Aegypti, et maris Magni litore finietur.
NUM|34|6|Plaga autem occidentalis a mari Magno incipiet et ipso fine claudetur.
NUM|34|7|Porro ad septentrionalem plagam a mari Magno termini incipient pervenientes usque ad montem Hor,
NUM|34|8|a quo venient in introitum Emath usque ad terminos Sedada.
NUM|34|9|Ibuntque confinia usque ad Zephrona et Asarenon. Hi erunt termini in parte aquilonis.
NUM|34|10|Inde metabuntur fines contra orientalem plagam de Asarenon usque Sephama;
NUM|34|11|et de Sephama descendent termini in Rebla ad orientem Ain; inde descendent et pervenient ad latus maris Chenereth in oriente
NUM|34|12|et tendent usque ad Iordanem, et ad ultimum Salsissimo claudentur mari.Hanc habebitis terram per fines suos in circuitu ".
NUM|34|13|Praecepitque Moyses filiis Israel dicens: " Haec erit terra, quam possidebitis sorte et quam iussit Dominus dari novem tribubus et dimidiae tribui.
NUM|34|14|Tribus enim filiorum Ruben per familias suas et tribus filiorum Gad iuxta cognationum numerum media quoque tribus Manasse,
NUM|34|15|id est duae semis tribus, acceperunt partem suam trans Iordanem contra Iericho ad orientalem plagam ".
NUM|34|16|Et ait Dominus ad Moysen:
NUM|34|17|" Haec sunt nomina virorum, qui terram vobis divident: Eleazar sacerdos et Iosue filius Nun
NUM|34|18|et singuli principes de tribubus singulis,
NUM|34|19|quorum ista sunt vocabula: de tribu Iudae Chaleb filius Iephonne;
NUM|34|20|de tribu Simeon Samuel filius Ammiud;
NUM|34|21|de tribu Beniamin Elidad filius Chaselon;
NUM|34|22|de tribu filiorum Dan Bocci filius Iogli.
NUM|34|23|Filiorum Ioseph: de tribu Manasse Hanniel filius Ephod,
NUM|34|24|de tribu Ephraim Camuel filius Sephtan.
NUM|34|25|De tribu Zabulon Elisaphan filius Pharnach;
NUM|34|26|de tribu Issachar dux Phaltiel filius Ozan;
NUM|34|27|de tribu Aser Ahiud filius Salomi;
NUM|34|28|de tribu Nephthali Phedael filius Ammiud ".
NUM|34|29|Hi sunt, quibus praecepit Dominus, ut dividerent filiis Israel terram Chanaan.
NUM|35|1|Haec quoque locutus est Do minus ad Moysen in campe stribus Moab supra Iordanem contra Iericho:
NUM|35|2|" Praecipe filiis Israel, ut dent Levitis de possessionibus suis urbes ad habitandum et suburbana earum per circuitum,
NUM|35|3|ut ipsi in oppidis maneant, et suburbana sint pecoribus ac substantiae et omnibus animalibus eorum;
NUM|35|4|quae a muris civitatum forinsecus per circuitum mille cubitos spatio tendentur.
NUM|35|5|Et mensurabitis extra civitatem contra orientem duo milia cubitorum, et contra meridiem similiter duo milia, ad mare quoque, quod respicit ad occidentem, eadem mensura erit, et septentrionalis plaga aequali termino finietur; eruntque urbes in medio et foris suburbana.
NUM|35|6|De ipsis autem oppidis, quae Levitis dabitis, sex erunt in fugitivorum auxilia separata, ut fugiat ad ea, qui nesciens fuderit sanguinem; et, exceptis his, alia quadraginta duo oppida dabitis,
NUM|35|7|id est simul quadraginta octo cum suburbanis suis.
NUM|35|8|Ipsaeque urbes, quas dabitis de possessionibus filiorum Israel, ab his, qui plus habent, plures auferetis, et, qui minus, pauciores; singuli iuxta mensuram hereditatis suae dabunt oppida Levitis ".
NUM|35|9|Ait Dominus ad Moysen:
NUM|35|10|" Loquere filiis Israel et dices ad eos: Quando transgressi fueritis Iordanem in terram Chanaan,
NUM|35|11|eligetis urbes, quae esse debeant in praesidia fugitivorum, qui nolentes sanguinem fuderint;
NUM|35|12|erunt vobis urbes refugii contra ultorem, et occisor non morietur, donec stet in conspectu congregationis, et causa illius iudicetur.
NUM|35|13|De ipsis autem sex urbibus, quae ad fugitivorum subsidia separantur,
NUM|35|14|tres erunt trans Iordanem et tres in terra Chanaan,
NUM|35|15|tam filiis Israel quam advenis atque peregrinis, ut confugiat ad eas sex, qui nolens sanguinem fuderit.
NUM|35|16|Si quis ferro percusserit, et mortuus fuerit, qui percussus est, reus erit homicidii et ipse morietur.
NUM|35|17|Si lapidem mortiferum iecerit, et ictus occiderit, similiter punietur.
NUM|35|18|Si ligno mortifero percusserit eum et interfecerit, homicida est; ipse morte punietur.
NUM|35|19|Ultor sanguinis homicidam interficiet: statim ut apprehenderit eum, interficiet.
NUM|35|20|Si per odium quis hominem impulerit vel iecerit quippiam in eum per insidias
NUM|35|21|aut, cum esset inimicus, manu percusserit, et ille mortuus fuerit, percussor homicidii reus erit: ultor sanguinis statim ut invenerit eum, iugulabit.
NUM|35|22|Quod si fortuitu et absque odio eum percusserit vel quidpiam in eum iecerit absque insidiis,
NUM|35|23|vel quemlibet lapidem mortiferum in eum devolverit, cum eum non vidisset, et ille mortuus est, quamvis eum non oderit nec quaesierit ei malum,
NUM|35|24|iudicabit congregatio inter percussorem et ultorem sanguinis secundum has regulas
NUM|35|25|et liberabit occisorem de manu ultoris sanguinis et reducet in civitatem refugii, ad quam confugerat, manebitque ibi, donec sacerdos magnus, qui oleo sancto unctus est, moriatur.
NUM|35|26|Si interfector extra fines civitatis refugii, in quam confugerat, exierit,
NUM|35|27|et invenerit eum ultor sanguinis ibi et interfecerit, absque noxa erit, qui eum occiderit;
NUM|35|28|debuerat enim profugus usque ad mortem pontificis in civitate refugii residere. Postquam autem ille obierit, homicida revertetur in terram suam.
NUM|35|29|Haec erunt vobis in legitima iudicii pro generationibus vestris, in cunctis habitationibus vestris.
NUM|35|30|Homicida sub testibus occidetur; ad unius testimonium nullus ad mortem condemnabitur.
NUM|35|31|Non accipietis pretium pro eo, qui reus est sanguinis, sed morietur.
NUM|35|32|Neque accipietis pretium, ut fugiat in civitatem refugii sui, ut revertatur et habitet in terra ante mortem sacerdotis.
NUM|35|33|Non polluetis terram habitationis vestrae, quia sanguis polluit terram, nec aliter expiari potest nisi per eius sanguinem, qui alterius sanguinem fuderit.
NUM|35|34|Non maculabitis terram habitationis vestrae, me commorante vobiscum. Ego enim sum Dominus, qui habito inter filios Israel ".
NUM|36|1|Accesserunt autem et princi pes familiarum tribus filio rum Galaad filii Machir filii Manasse de stirpe filiorum Ioseph; locutique sunt Moysi coram principibus familiarum Israel
NUM|36|2|atque dixerunt: " Tibi domino nostro praecepit Dominus, ut terram sorte divideres filiis Israel et ut filiabus Salphaad fratris nostri dares hereditatem debitam patri;
NUM|36|3|quas si alterius tribus homines uxores acceperint, sequetur possessio sua, et translata ad aliam tribum de nostra hereditate minuetur.
NUM|36|4|Atque ita fiet, ut cum iobeleus advenerit, addetur possessio earum possessioni tribus, ad quam pertinent, et a possessione tribus patrum nostrorum auferetur ".
NUM|36|5|Respondit Moyses filiis Israel et, Domino praecipiente, ait: " Recte tribus filiorum Ioseph locuta est,
NUM|36|6|et haec lex super filiabus Salphaad a Domino promulgata est: Nubant, quibus volunt, tantum ut suae tribus hominibus,
NUM|36|7|ne commisceatur possessio filiorum Israel de tribu in tribum; filii Israel adhaerebunt possessioni tribus patrum suorum,
NUM|36|8|et cunctae filiae heredes e filiis Israel maritos e cognatione tribus patrum suorum accipient, ut hereditas permaneat in familiis,
NUM|36|9|nec commisceatur possessio de tribu in tribum alteram, sed filii Israel adhaerebunt possessioni tribuum suarum ".
NUM|36|10|Sicut mandavit Dominus Moysi, sic fecerunt filiae Salphaad
NUM|36|11|et nupserunt Maala et Thersa et Hegla et Melcha et Noa filiis patruorum suorum
NUM|36|12|de familiis Manasse, qui fuit filius Ioseph; et possessio, quae illis fuerat attributa, mansit in tribu et familia patris earum.
NUM|36|13|Haec sunt mandata atque iudicia, quae mandavit Dominus per manum Moysi ad filios Israel in campestribus Moab supra Iordanem contra Iericho.
DEUT|1|1|Haec sunt verba, quae locutus est Moyses ad omnem Israel trans Iordanem in solitudine, in Araba contra Suph, inter Pharan et Thophel et Laban et Aseroth et Dizahab.
DEUT|1|2|Undecim dies de Horeb per viam montis Seir usque Cadesbarne.
DEUT|1|3|Quadragesimo anno, undecimo mense, prima die mensis locutus est Moyses ad filios Israel omnia, quae praeceperat illi Dominus ut diceret eis.
DEUT|1|4|Postquam percussit Sehon regem Amorraeorum, qui habitavit in Hesebon, et Og regem Basan, qui mansit in Astharoth et in Edrai,
DEUT|1|5|trans Iordanem in terra Moab coepitque Moyses explanare legem hanc et dicere:
DEUT|1|6|" Dominus Deus noster locutus est ad nos in Horeb dicens: "Sufficit vobis quod in hoc monte mansistis;
DEUT|1|7|convertimini et proficiscimini et venite ad montem Amorraeorum et ad omnes vicinos eius: in Araba atque montanis et in Sephela et in Nageb et iuxta litus maris, in terram Chananaeorum et in Libanum usque ad flumen magnum Euphraten.
DEUT|1|8|En, inquit, tradidi vobis terram: ingredimini et possidete eam, super qua iuravit Dominus patribus vestris, Abraham, Isaac et Iacob, ut daret illam eis et semini eorum post eos".
DEUT|1|9|Dixique vobis illo in tempore: Non possum solus sustinere vos;
DEUT|1|10|Dominus Deus vester multiplicavit vos, et estis hodie sicut stellae caeli plurimi.
DEUT|1|11|Dominus, Deus patrum vestrorum, addat ad hunc numerum multa milia et benedicat vobis, sicut locutus est vobis.
DEUT|1|12|Non valeo solus vestra negotia sustinere et pondus ac iurgia;
DEUT|1|13|date vobis viros sapientes et gnaros, et quorum conversatio sit probata in tribubus vestris, ut ponam eos vobis principes.
DEUT|1|14|Tunc respondistis mihi: "Bona res est, quam vis facere".
DEUT|1|15|Tulique principes de tribubus vestris viros sapientes et probatos et constitui eos principes super vos: tribunos et centuriones et quinquagenarios ac decanos et praefectos operum pro tribubus vestris.
DEUT|1|16|Praecepique iudicibus vestris in tempore illo: Audite causam fratrum vestrorum et, quod iustum est, iudicate, sive civis sit ille sive peregrinus.
DEUT|1|17|Non accipietis personam in iudicio; ita parvum audietis ut magnum nec timebitis cuiusquam personam, quia Dei iudicium est. Quod si difficile vobis aliquid visum fuerit, referte ad me, et ego audiam.
DEUT|1|18|Praecepique vobis in tempore illo omnia, quae facere deberetis.
DEUT|1|19|Profecti autem de Horeb transivimus per totam illam eremum maximam et terribilem, quam vidistis, per viam montis Amorraei, sicut praeceperat Dominus Deus noster nobis. Cumque venissemus in Cadesbarne,
DEUT|1|20|dixi vobis: Venistis ad montem Amorraei, quem Dominus Deus noster daturus est nobis.
DEUT|1|21|Vide terram, quam Dominus Deus tuus dat tibi: ascende et posside eam, sicut locutus est tibi Dominus, Deus patrum tuorum; noli metuere nec quidquam paveas.
DEUT|1|22|Et accessistis ad me vos omnes atque dixistis: "Mittamus viros ante nos, qui considerent terram et renuntient de itinere, per quod debeamus ascendere, et de civitatibus, ad quas pergere".
DEUT|1|23|Cumque mihi sermo placuisset, misi ex vobis duodecim viros singulos de tribubus suis.
DEUT|1|24|Qui cum perrexissent et ascendissent in montana, venerunt usque ad Nehelescol et, considerata terra,
DEUT|1|25|sumentes de fructibus eius attulerunt ad nos atque dixerunt: "Bona est terra, quam Dominus Deus noster daturus est nobis".
DEUT|1|26|Et noluistis ascendere, sed increduli ad sermonem Domini Dei vestri
DEUT|1|27|murmurastis in tabernaculis vestris atque dixistis: "Odit nos Dominus et idcirco eduxit nos de terra Aegypti, ut traderet nos in manu Amorraei atque deleret.
DEUT|1|28|Quo ascendemus? Fratres nostri terruerunt cor nostrum dicentes: Maxima multitudo est et nobis in statura procerior; urbes magnae et ad caelum usque munitae; etiam filios Enacim vidimus ibi".
DEUT|1|29|Et dixi vobis: Nolite metuere nec timeatis eos.
DEUT|1|30|Dominus Deus, qui ductor est vester, ipse pro vobis pugnabit, sicut fecit in Aegypto, vobis videntibus.
DEUT|1|31|Et in solitudine - ipse vidisti - portavit te Dominus Deus tuus, ut solet homo gestare parvulum filium suum, in omni via, per quam ambulastis, donec veniretis ad locum istum.
DEUT|1|32|Et nec sic quidem credidistis Domino Deo vestro,
DEUT|1|33|qui praecessit vos in via, et metatus est locum, in quo tentoria figere deberetis, nocte ostendens vobis iter per ignem et die per columnam nubis.
DEUT|1|34|Cumque audisset Dominus vocem sermonum vestrorum, iratus iuravit et ait:
DEUT|1|35|"Non videbit quispiam de viris generationis huius pessimae terram bonam, quam sub iuramento pollicitus sum patribus vestris,
DEUT|1|36|praeter Chaleb filium Iephonne: ipse enim videbit eam, et ipsi dabo terram, quam calcavit, et filiis eius, quia adimplevit ut sequeretur Dominum".
DEUT|1|37|Mihi quoque iratus Dominus propter vos dixit: "Nec tu ingredieris illuc;
DEUT|1|38|sed Iosue filius Nun minister tuus ipse intrabit illuc. Hunc robora, et ipse terram sorte dividat Israeli.
DEUT|1|39|Parvuli vestri, de quibus dixistis quod captivi ducerentur, et filii, qui hodie boni ac mali ignorant distantiam, ipsi ingredientur; et ipsis dabo terram, et possidebunt eam.
DEUT|1|40|Vos autem revertimini et abite in solitudinem per viam maris Rubri".
DEUT|1|41|Et respondistis mihi: "Peccavimus Domino; nos ascendemus atque pugnabimus, sicut praecepit nobis Dominus Deus noster". Cumque instructi armis pergeretis in montem,
DEUT|1|42|ait mihi Dominus: "Dic ad eos: Nolite ascendere neque pugnetis, non enim sum vobiscum, ne cadatis coram inimicis vestris".
DEUT|1|43|Locutus sum, et non audistis, sed adversantes imperio Domini et tumentes superbia ascendistis in montem.
DEUT|1|44|Itaque egressus Amorraeus, qui habitat in monte illo, obviam vobis, persecutus est vos, sicut solent apes persequi, et cecidit vos de Seir usque Horma.
DEUT|1|45|Cumque reversi ploraretis coram Domino, non audivit vos nec voci vestrae voluit acquiescere.
DEUT|1|46|Sedistis ergo in Cades multo illo tempore, dum ibi mansistis.
DEUT|2|1|Profectique inde venimus in solitudinem per viam maris Ru bri, sicut mihi dixerat Dominus; et circuivimus montem Seir longo tempore.
DEUT|2|2|Dixitque Dominus ad me:
DEUT|2|3|"Sufficit vobis circuire montem istum; ite contra aquilonem.
DEUT|2|4|Et populo praecipe dicens: Transibitis per terminos fratrum vestrorum filiorum Esau, qui habitant in Seir, et timebunt vos.
DEUT|2|5|Cavete ergo diligenter, ne moveamini contra eos; neque enim dabo vobis de terra eorum, quantum potest unius pedis calcare vestigium, quia in possessionem Esau dedi montem Seir.
DEUT|2|6|Cibos emetis ab eis pecunia et comedetis; etiam aquam emptam haurietis et bibetis.
DEUT|2|7|Dominus Deus tuus benedixit tibi in omni opere manuum tuarum; novit iter tuum, quomodo transieris solitudinem hanc magnam per quadraginta annos habitans tecum Dominus Deus tuus, et nihil tibi defuit".
DEUT|2|8|Cumque transissemus fratres nostros filios Esau, qui habitabant in Seir, per viam Arabae de Ailath et de Asiongaber, vertimus nos et venimus per iter, quod ducit in desertum Moab.
DEUT|2|9|Dixitque Dominus ad me: "Non pugnes contra Moabitas nec ineas adversus eos proelium; non enim dabo tibi quidquam de terra eorum, quia filiis Lot tradidi Ar in possessionem.
DEUT|2|10|- Emim primi fuerunt habitatores eius, populus magnus et multus et tam excelsus ut Enacim;
DEUT|2|11|ipsi quoque Raphaim reputabantur sicut Enacim; denique Moabitae appellant eos Emim.
DEUT|2|12|In Seir autem prius habitaverunt Horim; quibus expulsis atque deletis, habitaverunt filii Esau pro eis, sicut fecit Israel in terra possessionis suae, quam dedit eis Dominus C.
DEUT|2|13|Surgite ergo et transite torrentem Zared". Et transivimus torrentem Zared.
DEUT|2|14|Tempus autem, quo ambulavimus de Cadesbarne usque ad transitum torrentis Zared, triginta octo annorum fuit, donec consumeretur omnis generatio hominum bellatorum de castris, sicut iuraverat eis Dominus,
DEUT|2|15|cuius manus fuit adversum eos, ut interirent de castrorum medio.
DEUT|2|16|Postquam autem universi ceciderunt pugnatores de medio populi,
DEUT|2|17|locutus est Dominus ad me dicens:
DEUT|2|18|"Tu transibis hodie terminos Moab, urbem nomine Ar;
DEUT|2|19|et accedens in vicina filiorum Ammon, cave, ne pugnes contra eos nec movearis ad proelium; non enim dabo tibi de terra filiorum Ammon, quia filiis Lot dedi eam in possessionem.
DEUT|2|20|- Terra Raphaim reputata est et ipsa olim habitaverunt Raphaim in ea, quos Ammonitae vocant Zomzommim,
DEUT|2|21|populus magnus et multus et procerae longitudinis sicut Enacim, quos delevit Dominus a facie eorum et fecit illos habitare pro eis,
DEUT|2|22|sicut fecerat filiis Esau, qui habitant in Seir, delens Horim et terram eorum illis tradens, quam possident usque in praesens.
DEUT|2|23|Hevaeos quoque, qui habitabant in villis usque Gazam, Caphtorim, qui egressi de Caphtor deleverunt eos et habitaverunt pro illis C.
DEUT|2|24|Surgite! Proficiscimini et transite torrentem Arnon: ecce tradidi in manu tua Sehon regem Hesebon Amorraeum; et terram eius incipe possidere et committe adversus eum proelium.
DEUT|2|25|Hodie incipiam mittere terrorem atque formidinem tuam in populos, qui habitant sub omni caelo, ut, audito nomine tuo, paveant et contremiscant coram te".
DEUT|2|26|Misi ergo nuntios de solitudine Cademoth ad Sehon regem Hesebon verbis pacificis dicens:
DEUT|2|27|Transibo per terram tuam, publica gradiar via, non declinabo neque ad dexteram neque ad sinistram;
DEUT|2|28|alimenta pretio vende mihi, ut vescar, aquam pecunia tribue mihi, et sic bibam; tantum est ut mihi concedas transitum,
DEUT|2|29|sicut fecerunt mihi filii Esau, qui habitant in Seir, et Moabitae, qui morantur in Ar, donec veniam ad Iordanem et transeam in terram, quam Dominus Deus noster daturus est nobis.
DEUT|2|30|Noluitque Sehon rex Hesebon dare nobis transitum, quia induraverat Dominus Deus tuus spiritum eius et obfirmaverat cor illius, ut traderetur in manus tuas, sicut est in praesenti die.
DEUT|2|31|Dixitque Dominus ad me: "Ecce coepi tradere tibi Sehon et terram eius. Incipe possidere eam!".
DEUT|2|32|Egressusque est Sehon obviam nobis cum omni populo suo ad proelium in Iasa,
DEUT|2|33|et tradidit eum Dominus Deus noster nobis; percussimusque eum cum filiis suis et omni populo suo.
DEUT|2|34|Cunctasque urbes eius in tempore illo cepimus et percussimus anathemate singulas civitates cum viris ac mulieribus et parvulis; neminem reliquimus in eis superstitem,
DEUT|2|35|absque iumentis, quae in partem venere praedantium, et spoliis urbium, quas cepimus.
DEUT|2|36|Ab Aroer, quae est super ripam torrentis Arnon, et oppido, quod in valle situm est, usque Galaad non fuit civitas, quae nostras effugeret manus: omnia tradidit Dominus Deus noster nobis,
DEUT|2|37|absque terra filiorum Ammon, ad quam non accessisti, cunctis, quae adiacent torrenti Iaboc, et urbibus montanis universisque locis, a quibus nos prohibuit Dominus Deus noster.
DEUT|3|1|Itaque conversi ascendimus per iter Basan; egressusque est Og rex Basan in occursum nobis cum omni populo suo ad bellandum in Edrai.
DEUT|3|2|Dixitque Dominus ad me: "Ne timeas eum, quia in manu tua tradidi eum cum omni populo ac terra sua; faciesque ei, sicut fecisti Sehon regi Amorraeorum, qui habitavit in Hesebon".
DEUT|3|3|Tradidit ergo Dominus Deus noster in manibus nostris etiam Og regem Basan et universum populum eius; percussimusque eos usque ad internecionem.
DEUT|3|4|Et cepimus cunctas civitates eius in illo tempore. Non fuit oppidum, quod nos effugeret: sexaginta urbes, omnem regionem Argob, regnum Og in Basan.
DEUT|3|5|Cunctae urbes erant munitae muris altissimis portisque et vectibus, absque oppidis innumeris, quae non habebant muros.
DEUT|3|6|Et percussimus eos anathemate, sicut feceramus Sehon regi Hesebon, disperdentes omnem civitatem virosque ac mulieres et parvulos;
DEUT|3|7|iumenta autem et spolia urbium diripuimus.
DEUT|3|8|Tulimusque illo in tempore terram de manu duorum regum Amorraeorum, qui erant trans Iordanem, a torrente Arnon usque ad montem Hermon
DEUT|3|9|- Sidonii vocant Hermon Sarion et Amorraei Sanir -
DEUT|3|10|omnes civitates, quae sitae sunt in planitie, et universam terram Galaad et Basan usque Salcha et Edrai, civitates regni Og in Basan.
DEUT|3|11|- Solus quippe Og rex Basan remanserat de residuis Raphaim. Monstratur lectus eius ferreus. Nonne est in Rabba filiorum Ammon? Novem cubitos habet longitudinis et quattuor latitudinis ad mensuram cubiti virilis manus C.
DEUT|3|12|Terramque hanc possedimus in tempore illo ab Aroer, quae est super ripam torrentis Arnon, usque ad mediam partem montis Galaad; et civitates illius dedi Ruben et Gad.
DEUT|3|13|Reliquam autem partem Galaad et omnem Basan, regnum Og, tradidi mediae tribui Manasse, omnem regionem Argob. Cuncta Basan vocatur terra Raphaim.
DEUT|3|14|Iair filius Manasse possedit omnem regionem Argob usque ad terminos Gesuri et Maachathi; vocavitque ea ex nomine suo Basan Havoth Iair (id est villas Iair) usque in praesentem diem.
DEUT|3|15|Machir quoque dedi Galaad.
DEUT|3|16|Et tribubus Ruben et Gad dedi de terra Galaad usque ad torrentem Arnon, medium torrentis et confinium usque ad torrentem Iaboc, qui est terminus filiorum Ammon;
DEUT|3|17|et Arabam atque Iordanem et terminos a Chenereth usque ad mare Arabae, quod est mare Salis, ad radices montis Phasga contra orientem.
DEUT|3|18|Praecepique vobis in tempore illo dicens: Dominus Deus vester dedit vobis terram hanc in hereditatem; expediti praecedite fratres vestros filios Israel, omnes viri robusti,
DEUT|3|19|absque uxoribus et parvulis ac iumentis. Novi enim quod plura habeatis pecora, et in urbibus remanere debebunt, quas tradidi vobis,
DEUT|3|20|donec requiem tribuat Dominus fratribus vestris, sicut vobis tribuit, et possideant etiam ipsi terram, quam Dominus Deus vester daturus est eis trans Iordanem; tunc revertetur unusquisque in possessionem suam, quam dedi vobis.
DEUT|3|21|Iosue quoque in tempore illo praecepi dicens: Oculi tui viderunt, quae fecit Dominus Deus vester duobus his regibus; sic faciet omnibus regnis, ad quae transiturus es.
DEUT|3|22|Ne timeas eos: Dominus enim Deus vester pugnabit pro vobis.
DEUT|3|23|Precatusque sum Dominum in tempore illo dicens:
DEUT|3|24|Domine Deus, tu coepisti ostendere servo tuo magnitudinem tuam manumque fortissimam; neque enim est alius Deus vel in caelo vel in terra, qui possit facere opera tua et comparari fortitudini tuae.
DEUT|3|25|Transeam igitur et videam terram hanc optimam trans Iordanem et montem istum egregium et Libanum.
DEUT|3|26|Iratusque est Dominus mihi propter vos nec exaudivit me, sed dixit mihi: "Sufficit tibi; nequaquam ultra loquaris de hac re ad me.
DEUT|3|27|Ascende cacumen Phasgae et oculos tuos circumfer ad occidentem et aquilonem austrumque et orientem et aspice; nec enim transibis Iordanem istum.
DEUT|3|28|Praecipe Iosue et corrobora eum atque conforta, quia ipse praecedet populum istum et dividet eis terram, quam visurus es".
DEUT|3|29|Mansimusque in valle contra Bethphegor.
DEUT|4|1|Et nunc, Israel, audi praecepta et iudicia, quae ego doceo vos, ut facientes ea vivatis et ingredientes possideatis terram, quam Dominus, Deus patrum vestrorum, daturus est vobis.
DEUT|4|2|Non addetis ad verbum, quod vobis loquor, neque auferetis ex eo; custodite mandata Domini Dei vestri, quae ego praecipio vobis.
DEUT|4|3|Oculi vestri viderunt omnia, quae fecit Dominus contra Baalphegor, quomodo contriverit omnes cultores eius de medio vestri;
DEUT|4|4|vos autem, qui adhaeretis Domino Deo vestro, vivitis universi usque in praesentem diem.
DEUT|4|5|En docui vos praecepta atque iudicia, sicut mandavit mihi Dominus Deus meus, ut faceretis ea in terra, quam possessuri estis,
DEUT|4|6|et observaretis et impleretis opere. Haec est enim vestra sapientia et intellectus coram populis, ut audientes universa praecepta haec dicant: En populus sapiens et intellegens, gens magna haec!".
DEUT|4|7|Quae est enim alia natio tam grandis, quae habeat deos appropinquantes sibi, sicut Dominus Deus noster adest cunctis obsecrationibus nostris?
DEUT|4|8|Et quae est alia gens sic inclita, ut habeat praecepta iustaque iudicia, sicut est universa lex haec, quam ego proponam hodie ante oculos vestros?
DEUT|4|9|Custodi igitur temetipsum et animam tuam sollicite, ne obliviscaris verborum, quae viderunt oculi tui, et ne excidant de corde tuo cunctis diebus vitae tuae. Docebis ea filios ac nepotes tuos
DEUT|4|10|die, in quo stetisti coram Domino Deo tuo in Horeb, quando Dominus locutus est mihi: "Congrega ad me populum, ut audiant sermones meos et discant timere me omni tempore, quo vivunt in terra, doceantque filios suos".
DEUT|4|11|Et accessistis et stetistis ad radices montis, qui ardebat usque ad caelum, erantque in eo tenebrae, nubes et caligo.
DEUT|4|12|Locutusque est Dominus ad vos de medio ignis; vocem verborum audistis et formam penitus non vidistis.
DEUT|4|13|Et ostendit vobis pactum suum, quod praecepit, ut faceretis, et decem verba, quae scripsit in duabus tabulis lapideis.
DEUT|4|14|Mihique mandavit in illo tempore, ut docerem vos praecepta et iudicia, quae facere deberetis in terra, quam possessuri estis.
DEUT|4|15|Custodite igitur sollicite animas vestras. Non vidistis aliquam similitudinem in die, qua locutus est vobis Dominus in Horeb de medio ignis;
DEUT|4|16|ne forte corrupti faciatis vobis sculptam similitudinem, imaginem masculi vel feminae,
DEUT|4|17|similitudinem omnium iumentorum, quae sunt super terram, vel avium sub caelo volantium
DEUT|4|18|atque reptilium, quae moventur in terra, sive piscium, qui sub terra morantur in aquis;
DEUT|4|19|et ne forte oculis elevatis ad caelum videas solem et lunam et astra, omnem exercitum caeli, et errore deceptus adores ea et colas, quae attribuit Dominus Deus tuus cunctis gentibus, quae sub caelo sunt.
DEUT|4|20|Vos autem tulit Dominus et eduxit de fornace ferrea Aegypti, ut haberet populum hereditarium, sicut est in praesenti die.
DEUT|4|21|Iratusque est Dominus contra me propter sermones vestros et iuravit, ut non transirem Iordanem nec ingrederer terram optimam, quam Dominus Deus tuus daturus est tibi in haereditatem.
DEUT|4|22|Ecce morior in hac humo, non transibo Iordanem; vos transibitis et possidebitis terram egregiam hanc.
DEUT|4|23|Cavete, ne quando obliviscamini pacti Domini Dei vestri, quod pepigit vobiscum, et faciatis vobis sculptam similitudinem omnium, quae fieri Dominus Deus tuus prohibuit;
DEUT|4|24|quia Dominus Deus tuus ignis consumens est, Deus aemulator.
DEUT|4|25|Si genueris filios ac nepotes, et morati fueritis in terra corruptique feceritis aliquam similitudinem sculptam patrantes malum coram Domino Deo tuo, ut eum ad iracundiam provocetis,
DEUT|4|26|testes invoco contra vos hodie caelum et terram, cito perituros vos esse de terra, quam, transito Iordane, possessuri estis: non habitabitis in ea longo tempore, sed delebit vos Dominus
DEUT|4|27|atque disperget in gentes, et remanebitis pauci in nationibus, ad quas vos ducturus est Dominus.
DEUT|4|28|Ibique servietis diis, qui hominum manu fabricati sunt, ligno et lapidi, qui non vident nec audiunt nec comedunt nec odorantur.
DEUT|4|29|Cumque quaesieris ibi Dominum Deum tuum, invenies eum, si tamen toto corde quaesieris eum et tota anima tua.
DEUT|4|30|Postquam in tribulatione tua te invenerint omnia, quae praedicta sunt, novissimo tempore reverteris ad Dominum Deum tuum et audies vocem eius;
DEUT|4|31|quia Deus misericors Dominus Deus tuus est, non dimittet te nec omnino delebit neque obliviscetur pacti, in quo iuravit patribus tuis.
DEUT|4|32|Interroga de diebus antiquis, qui fuerunt ante te ex die, quo creavit Deus hominem super terram, et a summo caeli usque ad summum eius, si facta est aliquando huiuscemodi res magna, aut umquam cognitum est,
DEUT|4|33|num audivit populus vocem Dei loquentis de medio ignis, sicut tu audisti et vixisti?
DEUT|4|34|Aut tentavit Deus, ut ingrederetur et tolleret sibi gentem de medio nationis per tentationes, signa atque portenta, per pugnam et robustam manum extentumque brachium et terrores magnos, iuxta omnia, quae fecit pro vobis Dominus Deus vester in Aegypto, videntibus oculis tuis?
DEUT|4|35|Tibi monstratum est, ut scires quoniam Dominus ipse est Deus, et non est alius praeter eum.
DEUT|4|36|De caelo te fecit audire vocem suam, ut doceret te, et in terra ostendit tibi ignem suum maximum; et audisti verba illius de medio ignis,
DEUT|4|37|quia dilexit patres tuos et elegit semen eorum post eos. Eduxitque te vultu suo in virtute sua magna ex Aegypto,
DEUT|4|38|ut expelleret nationes maiores et fortiores te in introitu tuo et introduceret te daretque tibi terram earum in possessionem, sicut cernis in praesenti die.
DEUT|4|39|Scito ergo hodie et cogitato in corde tuo quod Dominus ipse sit Deus in caelo sursum et in terra deorsum, et non sit alius.
DEUT|4|40|Custodi praecepta eius atque mandata, quae ego praecipio tibi hodie, ut bene sit tibi et filiis tuis post te, et permaneas multo tempore super terram, quam Dominus Deus tuus daturus est tibi ".
DEUT|4|41|Tunc separavit Moyses tres civitates trans Iordanem ad orientalem plagam,
DEUT|4|42|ut confugiat ad eas, qui occiderit nolens proximum suum, nec fuerit inimicus ante unum et alterum diem, et ad harum aliquam urbium possit evadere et vivat:
DEUT|4|43|Bosor in solitudine, quae sita est in terra campestri, pro tribu Ruben, et Ramoth in Galaad pro tribu Gad et Golan in Basan pro tribu Manasse.
DEUT|4|44|Ista est lex, quam proposuit Moyses coram filiis Israel;
DEUT|4|45|haec testimonia et praecepta atque iudicia, quae locutus est ad filios Israel, quando egressi sunt de Aegypto,
DEUT|4|46|trans Iordanem in valle contra Bethphegor, in terra Sehon regis Amorraei, qui habitavit in Hesebon, quem percussit Moyses et filii Israel egressi ex Aegypto.
DEUT|4|47|Et possederunt terram eius et terram Og regis Basan, duorum regum Amorraeorum, qui erant trans Iordanem ad solis ortum,
DEUT|4|48|ab Aroer, quae sita est super ripam torrentis Arnon, usque ad montem Sion, qui est Hermon,
DEUT|4|49|omnem Arabam trans Iordanem ad orientalem plagam usque ad mare Arabae et usque ad radices montis Phasga.
DEUT|5|1|Vocavitque Moyses omnem Israelem et dixit ad eos: " Audi, Israel, praecepta atque iudicia, quae ego loquor in auribus vestris hodie; discite ea et opere complete.
DEUT|5|2|Dominus Deus noster pepigit nobiscum foedus in Horeb.
DEUT|5|3|Non cum patribus nostris iniit pactum hoc sed nobiscum, qui in praesentiarum hic sumus, omnibus nobis, qui vivimus.
DEUT|5|4|Facie ad faciem locutus est vobis in monte de medio ignis;
DEUT|5|5|ego sequester et medius fui inter Dominum et vos in tempore illo, ut annuntiarem vobis verba eius; timuistis enim ignem et non ascendistis in montem. Et ait:
DEUT|5|6|"Ego Dominus Deus tuus, qui eduxi te de terra Aegypti, de domo servitutis.
DEUT|5|7|Non habebis deos alienos in conspectu meo.
DEUT|5|8|Non facies tibi sculptile nec similitudinem omnium, quae in caelo sunt desuper et quae in terra deorsum et quae versantur in aquis sub terra.
DEUT|5|9|Non adorabis ea et non coles: Ego enim sum Dominus Deus tuus, Deus aemulator, reddens iniquitatem patrum super filios in tertiam et quartam generationem his, qui oderunt me,
DEUT|5|10|et faciens misericordiam in multa milia diligentibus me et custodientibus praecepta mea.
DEUT|5|11|Non usurpabis nomen Domini Dei tui frustra, quia non erit impunitus, qui super re vana nomen eius assumpserit.
DEUT|5|12|Observa diem sabbati, ut sanctifices eum, sicut praecepit tibi Dominus Deus tuus.
DEUT|5|13|Sex diebus operaberis et facies omnia opera tua.
DEUT|5|14|Septimus dies sabbatum est Domino Deo tuo. Non facies in eo quidquam operis tu et filius tuus et filia, servus et ancilla et bos et asinus et omne iumentum tuum et peregrinus tuus, qui est intra portas tuas, ut requiescat servus tuus et ancilla tua sicut et tu.
DEUT|5|15|Memento quod et ipse servieris in Aegypto, et eduxerit te inde Dominus Deus tuus in manu forti et brachio extento: idcirco praecepit tibi, ut observares diem sabbati.
DEUT|5|16|Honora patrem tuum et matrem, sicut praecepit tibi Dominus Deus tuus, ut longo vivas tempore et bene sit tibi in terra, quam Dominus Deus tuus daturus est tibi.
DEUT|5|17|Non occides.
DEUT|5|18|Neque moechaberis.
DEUT|5|19|Furtumque non facies.
DEUT|5|20|Nec loqueris contra proximum tuum falsum testimonium.
DEUT|5|21|Nec concupisces uxorem proximi tui. Nec desiderabis domum proximi tui, non agrum, non servum, non ancillam, non bovem, non asinum et universa, quae illius sunt".
DEUT|5|22|Haec verba locutus est Dominus ad omnem multitudinem vestram in monte, de medio ignis et nubis et caliginis voce magna nihil addens amplius; et scripsit ea in duabus tabulis lapideis, quas tradidit mihi.
DEUT|5|23|Vos autem, postquam audistis vocem de medio tenebrarum et montem ardere vidistis, accessistis ad me omnes principes tribuum et maiores natu
DEUT|5|24|atque dixistis: "Ecce ostendit nobis Dominus Deus noster maiestatem et magnitudinem suam; vocem eius audivimus de medio ignis et probavimus hodie quod, loquente Deo cum homine, vixerit homo.
DEUT|5|25|Nunc autem cur moriemur, et devorabit nos ignis hic maximus? Si enim audierimus ultra vocem Domini Dei nostri, moriemur.
DEUT|5|26|Quid est omnis caro, ut audiat vocem Dei viventis, qui de medio ignis loquitur, sicut nos audivimus, et possit vivere?
DEUT|5|27|Tu magis accede et audi cuncta, quae dixerit Dominus Deus noster, et tu loqueris ad nos cuncta, quae dixerit Dominus Deus noster tibi, et nos audientes faciemus ea".
DEUT|5|28|Quod cum audisset Dominus, ait ad me: "Audivi vocem verborum populi huius, quae locuti sunt tibi: bene omnia sunt locuti.
DEUT|5|29|Quis det talem eos habere mentem, ut timeant me et custodiant universa mandata mea in omni tempore, ut bene sit eis et filiis eorum in sempiternum?
DEUT|5|30|Vade et dic eis: Revertimini in tentoria vestra.
DEUT|5|31|Tu vero, hic sta mecum, et loquar tibi omnia mandata et praecepta atque iudicia, quae docebis eos, ut faciant ea in terra, quam dabo illis in possessionem".
DEUT|5|32|Custodite igitur et facite, quae praecepit Dominus Deus vester vobis; non declinabitis neque ad dexteram neque ad sinistram,
DEUT|5|33|sed per totam viam, quam praecepit Dominus Deus vester, ambulabitis, ut vivatis, et bene sit vobis, et protelentur dies in terra possessionis vestrae.
DEUT|6|1|Haec sunt mandata et praecep ta atque iudicia, quae mandavit Dominus Deus vester, ut docerem vos, et faciatis ea in terra, ad quam transgredimini possidendam;
DEUT|6|2|ut timeas Dominum Deum tuum et custodias omnia praecepta et mandata eius, quae ego praecipio tibi et filiis ac nepotibus tuis, cunctis diebus vitae tuae, ut prolongentur dies tui.
DEUT|6|3|Audi, Israel, et observa, ut facias, et bene sit tibi, et multipliceris amplius, sicut pollicitus est Dominus, Deus patrum tuorum, tibi terram lacte et melle manantem.
DEUT|6|4|Audi, Israel: Dominus Deus noster Dominus unus est.
DEUT|6|5|Diliges Dominum Deum tuum ex toto corde tuo et ex tota anima tua et ex tota fortitudine tua.
DEUT|6|6|Eruntque verba haec, quae ego praecipio tibi hodie, in corde tuo,
DEUT|6|7|et inculcabis ea filiis tuis et loqueris ea sedens in domo tua et ambulans in itinere, decumbens atque consurgens;
DEUT|6|8|et ligabis ea quasi signum in manu tua, eruntque quasi appensum quid inter oculos tuos,
DEUT|6|9|scribesque ea in postibus domus tuae et in portis tuis.
DEUT|6|10|Cumque introduxerit te Dominus Deus tuus in terram, pro qua iuravit patribus tuis Abraham, Isaac et Iacob, ut daret tibi, civitates magnas et optimas, quas non aedificasti,
DEUT|6|11|domos plenas cunctarum opum, quas non implevisti, cisternas, quas non fodisti, vineta et oliveta, quae non plantasti, et comederis et saturatus fueris,
DEUT|6|12|cave diligenter, ne obliviscaris Domini, qui eduxit te de terra Aegypti, de domo servitutis:
DEUT|6|13|Dominum Deum tuum timebis et ipsi servies ac per nomen illius iurabis.
DEUT|6|14|Non ibitis post deos alienos, de diis gentium, quae in circuitu vestro sunt,
DEUT|6|15|quoniam Deus aemulator Dominus Deus tuus in medio tui; ne quando irascatur furor Domini Dei tui contra te et auferat te de superficie terrae.
DEUT|6|16|Non tentabitis Dominum Deum vestrum, sicut tentastis in Massa.
DEUT|6|17|Custodite mandata Domini Dei vestri ac testimonia et praecepta, quae praecepit tibi;
DEUT|6|18|et fac, quod rectum est et bonum in conspectu Domini, ut bene sit tibi, et ingressus possideas terram optimam, de qua iuravit Dominus patribus tuis,
DEUT|6|19|ut deleret omnes inimicos tuos coram te, sicut locutus est Dominus.
DEUT|6|20|Cumque interrogaverit te filius tuus cras dicens: "Quid sibi volunt testimonia haec et praecepta atque iudicia, quae praecepit Dominus Deus noster vobis?",
DEUT|6|21|dices ei: "Servi eramus pharaonis in Aegypto, et eduxit nos Dominus de Aegypto in manu forti
DEUT|6|22|fecitque signa atque prodigia magna et pessima in Aegypto contra pharaonem et omnem domum illius in conspectu nostro;
DEUT|6|23|et eduxit nos inde, ut introductis daret terram, super qua iuravit patribus nostris.
DEUT|6|24|Praecepitque nobis Dominus, ut faciamus omnia praecepta haec et timeamus Dominum Deum nostrum, et bene sit nobis cunctis diebus vitae nostrae, sicut est hodie.
DEUT|6|25|Eritque iustitia nobis, si custodierimus et fecerimus omnia mandata haec coram Domino Deo nostro, sicut mandavit nobis".
DEUT|7|1|Cum introduxerit te Dominus Deus tuus in terram, quam pos sessurus ingredieris, et deleverit gentes multas coram te, Hetthaeum et Gergesaeum et Amorraeum, Chananaeum et Pherezaeum et Hevaeum et Iebusaeum, septem gentes multo maioris numeri quam tu es et robustiores te,
DEUT|7|2|tradideritque eas Dominus Deus tuus tibi, percuties eas usque ad internecionem. Non inibis cum eis foedus nec misereberis earum
DEUT|7|3|neque sociabis cum eis coniugia; filiam tuam non dabis filio eius nec filiam illius accipies filio tuo,
DEUT|7|4|quia seducet filium tuum, ne sequatur me et ut serviat diis alienis, irasceturque furor Domini contra vos et delebit te cito.
DEUT|7|5|Quin potius haec facietis eis: aras eorum subvertite et confringite lapides et palos lucosque succidite et sculptilia comburite;
DEUT|7|6|quia populus sanctus es Domino Deo tuo. Te elegit Dominus Deus tuus, ut sis ei populus peculiaris de cunctis populis, qui sunt super terram.
DEUT|7|7|Non quia cunctas gentes numero vincebatis, vobis iunctus est Dominus et elegit vos, cum omnibus sitis populis pauciores,
DEUT|7|8|sed quia dilexit vos Dominus et custodivit iuramentum, quod iuravit patribus vestris, eduxit vos in manu forti et redemit te de domo servitutis, de manu pharaonis regis Aegypti.
DEUT|7|9|Et scies quia Dominus Deus tuus ipse est Deus, Deus fidelis, custodiens pactum et misericordiam diligentibus se et his, qui custodiunt mandata eius, in mille generationes
DEUT|7|10|et reddens odientibus se protinus, ita ut disperdat eos et ultra non differat, protinus eis restituens, quod merentur.
DEUT|7|11|Custodi ergo mandata et praecepta atque iudicia, quae ego mando tibi hodie, ut facias.
DEUT|7|12|Si audieritis haec iudicia et custodieritis ea et feceritis, custodiet et Dominus Deus tuus tibi pactum et misericordiam, quam iuravit patribus tuis,
DEUT|7|13|et diliget te et benedicet tibi ac multiplicabit te benedicetque fructui ventris tui et fructui terrae tuae, frumento tuo atque vindemiae, oleo et partui armentorum et incremento ovium tuarum super terram, pro qua iuravit patribus tuis, ut daret eam tibi.
DEUT|7|14|Benedictus eris prae omnibus populis. Non erit apud te sterilis utriusque sexus, tam in hominibus quam in gregibus tuis.
DEUT|7|15|Auferet Dominus a te omnem languorem; et infirmitates Aegypti pessimas, quas novisti, non inferet tibi, sed cunctis hostibus tuis.
DEUT|7|16|Devorabis omnes populos, quos Dominus Deus tuus daturus est tibi; non parcet eis oculus tuus, nec servies diis eorum, ne sint in ruinam tui.
DEUT|7|17|Si dixeris in corde tuo: "Plures sunt gentes istae quam ego; quomodo potero delere eas?",
DEUT|7|18|noli metuere eas, sed recordare, quae fecerit Dominus Deus tuus pharaoni et cunctis Aegyptiis,
DEUT|7|19|plagas maximas, quas viderunt oculi tui, et signa atque portenta manumque robustam et extentum brachium, ut educeret te Dominus Deus tuus; sic faciet cunctis populis, quos metuis.
DEUT|7|20|Insuper et crabrones mittet Dominus Deus tuus in eos, donec deleat omnes atque disperdat, qui te fugerint et latere potuerint.
DEUT|7|21|Non timebis eos, quia Dominus Deus tuus in medio tui est, Deus magnus et terribilis.
DEUT|7|22|Ipse consumet nationes has in conspectu tuo paulatim atque per partes. Non poteris delere eas cito, ne multiplicentur contra te bestiae terrae.
DEUT|7|23|Dabitque eos Dominus Deus tuus in conspectu tuo et conturbabit illos conturbatione magna, donec penitus deleantur.
DEUT|7|24|Tradetque reges eorum in manus tuas, et disperdes nomina eorum sub caelo; nullus poterit resistere tibi, donec conteras eos.
DEUT|7|25|Sculptilia eorum igne combures; non concupisces argentum et aurum, quibus vestita sunt, neque assumes ex eis tibi quidquam, ne offendas propterea, quia abominatio est Domini Dei tui.
DEUT|7|26|Nec inferes abominationem in domum tuam, ne fias anathema sicut et illa est; quasi spurcitiam detestaberis et velut inquinamentum ac sordes abominationi habebis, quia anathema est.
DEUT|8|1|Omne mandatum, quod ego praecipio tibi hodie, cave dili genter ut facias, ut possitis vivere et multiplicemini ingressique possideatis terram, pro qua iuravit Dominus patribus vestris.
DEUT|8|2|Et recordaberis cuncti itineris, per quod adduxit te Dominus Deus tuus his quadraginta annis per desertum, ut affligeret te atque tentaret, et nota fierent, quae in tuo animo versabantur, utrum custodires mandata illius an non.
DEUT|8|3|Afflixit te penuria et dedit tibi cibum manna, quem ignorabas tu et patres tui, ut ostenderet tibi quod non in solo pane vivat homo, sed in omni verbo, quod egreditur de ore Domini.
DEUT|8|4|Vestimentum tuum, quo operiebaris, nequaquam defecit, et pes tuus non intumuit his quadraginta annis.
DEUT|8|5|Recogites ergo in corde tuo quia, sicut erudit homo filium suum, sic Dominus Deus tuus erudivit te,
DEUT|8|6|ut custodias mandata Domini Dei tui et ambules in viis eius et timeas eum.
DEUT|8|7|Dominus enim Deus tuus introducet te in terram bonam, terram rivorum aquarum et fontium, in cuius campis et montibus erumpunt fluviorum abyssi,
DEUT|8|8|terram frumenti, hordei ac vinearum, in qua ficus et malogranata et oliveta nascuntur, terram olei ac mellis,
DEUT|8|9|ubi absque ulla penuria comedes panem tuum et rerum omnium abundantia perfrueris; cuius lapides ferrum sunt, et de montibus eius aeris metalla fodiuntur;
DEUT|8|10|ut, cum comederis et satiatus fueris, benedicas Domino Deo tuo pro terra optima, quam dedit tibi.
DEUT|8|11|Observa et cave, ne quando obliviscaris Domini Dei tui et neglegas mandata eius atque iudicia et praecepta, quae ego praecipio tibi hodie;
DEUT|8|12|ne, postquam comederis et satiatus fueris, domos pulchras aedificaveris et habitaveris in eis
DEUT|8|13|habuerisque armenta et ovium greges multos, argenti et auri cunctarumque rerum copiam,
DEUT|8|14|elevetur cor tuum, et obliviscaris Domini Dei tui, qui eduxit te de terra Aegypti, de domo servitutis,
DEUT|8|15|et ductor tuus fuit in solitudine magna atque terribili, in qua erat serpens adurens et scorpio ac terra arida et nullae omnino aquae; qui eduxit tibi rivos de petra durissima
DEUT|8|16|et cibavit te manna in solitudine, quod nescierunt patres tui, et, postquam afflixit ac probavit te, ad extremum misertus est tui,
DEUT|8|17|ne diceres in corde tuo: "Fortitudo mea et robur manus meae haec mihi omnia praestiterunt";
DEUT|8|18|sed recorderis Domini Dei tui, quod ipse vires tibi praebuerit, ut consequereris prosperitatem, ut impleret pactum suum, super quo iuravit patribus tuis, sicut praesens indicat dies.
DEUT|8|19|Sin autem oblitus Domini Dei tui secutus fueris deos alienos coluerisque illos et adoraveris, ecce nunc testificor vobis quod omnino dispereatis:
DEUT|8|20|sicut gentes, quas delevit Dominus in introitu vestro, ita et vos peribitis, si inoboedientes fueritis voci Domini Dei vestri.
DEUT|9|1|Audi, Israel: Tu transgredieris hodie Iordanem, ut possideas nationes maximas et fortiores te, civitates ingentes et ad caelum usque muratas,
DEUT|9|2|populum magnum atque sublimem, filios Enacim, quos ipse nosti et audisti, quibus nullus potest ex adverso resistere.
DEUT|9|3|Scies ergo hodie quod Dominus Deus tuus ipse transibit ante te ignis devorans, qui conteret eos atque subiciet ante faciem tuam, ut velociter expellas et deleas eos, sicut locutus est tibi.
DEUT|9|4|Ne dicas in corde tuo, cum deleverit eos Dominus Deus tuus in conspectu tuo: "Propter iustitiam meam introduxit me Dominus, ut terram hanc possiderem", cum propter impietates nationum istarum expellat eas Dominus ante te.
DEUT|9|5|Neque enim propter iustitiam tuam et aequitatem cordis tui ingredieris, ut possideas terras earum, sed quia illae egerunt impie, introeunte te, Dominus Deus tuus expellet eos ante te, et ut compleat verbum suum Dominus, quod sub iuramento pollicitus est patribus tuis, Abraham, Isaac et Iacob.
DEUT|9|6|Scito igitur quod non propter iustitiam tuam Dominus Deus tuus dederit tibi terram hanc optimam in possessionem, cum durissimae cervicis sis populus.
DEUT|9|7|Memento et ne obliviscaris quomodo ad iracundiam provocaveris Dominum Deum tuum in solitudine; ex eo die, quo egressus es ex Aegypto, usque ad locum istum adversum Dominum contendistis.
DEUT|9|8|Nam et in Horeb provocastis eum, et iratus delere vos voluit,
DEUT|9|9|quando ascendi in montem, ut acciperem tabulas lapideas, tabulas pacti, quod pepigit vobiscum Dominus, et perseveravi in monte quadraginta diebus ac noctibus panem non comedens et aquam non bibens.
DEUT|9|10|Deditque mihi Dominus duas tabulas lapideas scriptas digito Dei et continentes omnia verba, quae vobis locutus est in monte de medio ignis, quando contio populi congregata est.
DEUT|9|11|Cumque transissent quadraginta dies et totidem noctes, dedit mihi Dominus duas tabulas lapideas, tabulas foederis,
DEUT|9|12|dixitque mihi: "Surge et descende hinc cito, quia peccavit populus tuus, quem eduxisti de Aegypto: deseruerunt velociter viam, quam praecepi eis, feceruntque sibi conflatile".
DEUT|9|13|Rursumque ait Dominus ad me: "Cerno quod populus iste durae cervicis sit;
DEUT|9|14|dimitte me, ut conteram eos et deleam nomen eorum sub caelo et faciam te in gentem, quae hac fortior et maior sit".
DEUT|9|15|Cumque reversus de monte ardente descenderem et duas tabulas foederis utraque tenerem manu
DEUT|9|16|vidissemque vos peccasse Domino Deo vestro et fecisse vobis vitulum conflatilem ac deseruisse velociter viam eius, quam Dominus vobis praeceperat,
DEUT|9|17|arripui duas tabulas et proieci eas de manibus meis confregique eas in conspectu vestro;
DEUT|9|18|et procidi ante Dominum, sicut prius quadraginta diebus et noctibus panem non comedens et aquam non bibens propter omnia peccata vestra, quae gessistis contra Dominum et eum ad iracundiam provocastis;
DEUT|9|19|timui enim indignationem et iram illius, qua adversum vos concitatus delere vos voluit. Et exaudivit me Dominus etiam hac vice.
DEUT|9|20|Adversum Aaron quoque vehementer iratus voluit eum conterere; et pro illo similiter tunc deprecatus sum.
DEUT|9|21|Peccatum autem vestrum, quod feceratis, id est vitulum, arripiens igne combussi et in frusta comminuens omninoque in pulverem redigens proieci in torrentem, qui de monte descendit.
DEUT|9|22|In Tabera quoque et in Massa et in Cibrottaava provocastis Dominum;
DEUT|9|23|et quando misit Dominus vos de Cadesbarne dicens: "Ascendite et possidete terram, quam dedi vobis", contempsistis imperium Domini Dei vestri et non credidistis ei neque vocem eius audire voluistis;
DEUT|9|24|semper fuistis rebelles contra Dominum a die, qua nosse vos coepi.
DEUT|9|25|Et iacui coram Domino quadraginta diebus ac noctibus, quibus eum suppliciter deprecabar, ne deleret vos, ut fuerat comminatus.
DEUT|9|26|Et orans dixi: Domine Deus, ne disperdas populum tuum et hereditatem tuam, quam redemisti in magnitudine tua, quos eduxisti de Aegypto in manu forti.
DEUT|9|27|Recordare servorum tuorum Abraham, Isaac et Iacob; ne aspicias duritiam populi huius et impietatem atque peccatum,
DEUT|9|28|ne forte dicant habitatores terrae, de qua eduxisti nos: "Non poterat Dominus introducere eos in terram, quam pollicitus est eis, et oderat illos; idcirco eduxit, ut interficeret eos in solitudine".
DEUT|9|29|Attamen ipsi sunt populus tuus et hereditas tua, quos eduxisti in fortitudine tua magna et in brachio tuo extento.
DEUT|10|1|In tempore illo dixit Dominus ad me: "Dola tibi duas tabulas lapideas, sicut priores fuerunt, et ascende ad me in montem faciesque tibi arcam ligneam.
DEUT|10|2|Et scribam in tabulis verba, quae fuerunt in his, quas ante confregisti, ponesque eas in arca".
DEUT|10|3|Feci igitur arcam de lignis acaciae; cumque dolassem duas tabulas lapideas instar priorum, ascendi in montem habens eas in manibus.
DEUT|10|4|Scripsitque in tabulis iuxta id quod prius scripserat, verba decem, quae locutus est Dominus ad vos in monte de medio ignis, quando populus congregatus est, et dedit eas mihi.
DEUT|10|5|Reversusque de monte descendi et posui tabulas in arcam, quam feceram; quae hucusque ibi sunt, sicut mihi praecepit Dominus.
DEUT|10|6|Filii autem Israel castra moverunt ex Berothbeneiacan in Mosera, ubi Aaron mortuus ac sepultus est; pro quo sacerdotio functus est Eleazar filius eius.
DEUT|10|7|Inde venerunt in Gadgad; de quo loco profecti castrametati sunt in Ietebatha, in terra torrentium aquarum.
DEUT|10|8|Eo tempore separavit Dominus tribum Levi, ut portaret arcam foederis Domini et staret coram eo in ministerio ac benediceret in nomine illius usque in praesentem diem.
DEUT|10|9|Quam ob rem non habuit Levi partem neque hereditatem cum fratribus suis, quia ipse Dominus hereditas eius est, sicut promisit ei Dominus Deus tuus.
DEUT|10|10|Ego autem steti in monte sicut prius quadraginta diebus ac noctibus, exaudivitque me Dominus etiam hac vice et te perdere noluit.
DEUT|10|11|Dixitque mihi: "Surge, vade et praecede populum, ut ingrediatur et possideat terram, quam iuravi patribus eorum, ut traderem eis".
DEUT|10|12|Et nunc, Israel, quid Dominus Deus tuus petit a te, nisi ut timeas Dominum Deum tuum et ambules in viis eius et diligas eum ac servias Domino Deo tuo in toto corde tuo et in tota anima tua
DEUT|10|13|custodiasque mandata Domini et praecepta eius, quae ego hodie praecipio, ut bene sit tibi?
DEUT|10|14|En Domini Dei tui caelum est et caelum caeli, terra et omnia, quae in ea sunt;
DEUT|10|15|et tamen patribus tuis conglutinatus est Dominus et amavit eos elegitque semen eorum post eos, id est vos, de cunctis gentibus, sicut hodie comprobatur.
DEUT|10|16|Circumcidite igitur praeputium cordis vestri et cervicem vestram, ne induretis amplius,
DEUT|10|17|quia Dominus Deus vester ipse est Deus deorum et Dominus dominantium, Deus magnus, potens et terribilis, qui personam non accipit nec munera,
DEUT|10|18|facit iudicium pupillo et viduae, amat peregrinum et dat ei victum atque vestitum.
DEUT|10|19|Et vos ergo, amate peregrinos, quia et ipsi fuistis advenae in terra Aegypti.
DEUT|10|20|Dominum Deum tuum timebis et ei servies, ipsi adhaerebis iurabisque in nomine illius.
DEUT|10|21|Ipse est laus tua et Deus tuus, qui fecit tibi haec magnalia et terribilia, quae viderunt oculi tui.
DEUT|10|22|In septuaginta animabus descenderunt patres tui in Aegyptum; et ecce nunc multiplicavit te Dominus Deus tuus sicut astra caeli.
DEUT|11|1|Ama itaque Dominum Deum tuum et custodi obser vationem eius et praecepta, iudicia atque mandata omni tempore.
DEUT|11|2|Cognoscite hodie, quae ignorant filii vestri, qui non viderunt disciplinam Domini Dei vestri, magnalia eius et robustam manum extentumque brachium,
DEUT|11|3|signa et opera, quae fecit in medio Aegypti pharaoni regi et universae terrae eius
DEUT|11|4|omnique exercitui Aegyptiorum et equis ac curribus; quomodo operuerint eos aquae maris Rubri, cum vos persequerentur, et deleverit eos Dominus usque in praesentem diem;
DEUT|11|5|vobisque, quae fecerit in solitudine, donec veniretis ad hunc locum;
DEUT|11|6|et Dathan atque Abiram filiis Eliab, qui fuit filius Ruben, quos aperto ore suo terra absorbuit cum domibus et tabernaculis et universa substantia eorum, quam habebant in medio Israel.
DEUT|11|7|Oculi vestri viderunt omnia opera Domini magna, quae fecit,
DEUT|11|8|ut custodiatis universa mandata, quae ego hodie praecipio vobis, ut roboremini et possitis introire et possidere terram, ad quam ingredimini,
DEUT|11|9|multoque in ea vivatis tempore, quam sub iuramento pollicitus est Dominus patribus vestris et semini eorum, lacte et melle manantem.
DEUT|11|10|Terra enim, ad quam ingredieris possidendam, non est sicut terra Aegypti, de qua existis, ubi, iacto semine, in hortorum morem aquae pede ducuntur irriguae;
DEUT|11|11|sed montuosa est et campestris, de caelo exspectans pluvias,
DEUT|11|12|quam Dominus Deus tuus semper invisit, et oculi illius in ea sunt a principio anni usque ad finem eius.
DEUT|11|13|Si ergo oboedieritis mandatis meis, quae hodie praecipio vobis, ut diligatis Dominum Deum vestrum et serviatis ei in toto corde vestro et in tota anima vestra,
DEUT|11|14|dabo pluviam terrae vestrae temporaneam et serotinam in tempore suo, ut colligas frumentum et vinum et oleum,
DEUT|11|15|et dabit fenum ex agris ad pascenda iumenta, et ut ipse comedas ac satureris.
DEUT|11|16|Cavete, ne decipiatur cor vestrum, et recedatis a Domino serviatisque diis alienis et adoretis eos,
DEUT|11|17|iratusque Dominus contra vos claudat caelum, et pluviae non descendant, nec terra det fructum suum, pereatisque velociter de terra optima, quam Dominus daturus est vobis.
DEUT|11|18|Ponite haec verba mea in cordibus et in animis vestris et ligate ea pro signo in manibus et inter oculos vestros collocate quasi appensum quid.
DEUT|11|19|Docete ea filios vestros, de illis loquendo, quando sederis in domo tua et ambulaveris in via et accubueris atque surrexeris.
DEUT|11|20|Scribes ea super postes domus tuae et portas tuas,
DEUT|11|21|ut multiplicentur dies tui et filiorum tuorum in terra, quam iuravit Dominus patribus tuis, ut daret eis, quamdiu caelum imminet terrae.
DEUT|11|22|Si enim custodieritis omnia mandata haec, quae ego praecipio vobis, et feceritis ea, ut diligatis Dominum Deum vestrum et ambuletis in omnibus viis eius adhaerentes ei,
DEUT|11|23|disperdet Dominus omnes gentes istas ante faciem vestram, et possidebitis eas, quae maiores et fortiores vobis sunt;
DEUT|11|24|omnis locus, quem calcaverit pes vester, vester erit. A deserto et a Libano, a flumine magno Euphrate usque ad mare occidentale erunt termini vestri.
DEUT|11|25|Nullus stabit contra vos; terrorem vestrum et formidinem dabit Dominus Deus vester super omnem terram, quam calcaturi estis, sicut locutus est vobis.
DEUT|11|26|En propono in conspectu vestro hodie benedictionem et maledictionem:
DEUT|11|27|benedictionem, si oboedieritis mandatis Domini Dei vestri, quae ego hodie praecipio vobis;
DEUT|11|28|maledictionem, si non oboedieritis mandatis Domini Dei vestri, sed recesseritis de via, quam ego nunc ostendo vobis, et ambulaveritis post deos alienos, quos ignoratis.
DEUT|11|29|Cum introduxerit te Dominus Deus tuus in terram, ad quam pergis habitandam, pones benedictionem super montem Garizim, maledictionem super montem Hebal,
DEUT|11|30|qui sunt trans Iordanem, post viam quae vergit ad solis occubitum in terra Chananaei, qui habitat in Araba contra Galgalam, quae est iuxta Quercus Moreh.
DEUT|11|31|Vos enim transibitis Iordanem, ut possideatis terram, quam Dominus Deus vester daturus est vobis, et habitetis in illa.
DEUT|11|32|Videte ergo ut impleatis omnia praecepta atque iudicia, quae ego hodie ponam in conspectu vestro.
DEUT|12|1|Haec sunt praecepta atque iudicia, quae facere debetis in terra, quam Dominus, Deus patrum tuorum, daturus est tibi, ut possideas eam cunctis diebus, quibus super humum gradieris.
DEUT|12|2|Subvertite omnia loca, in quibus coluerunt gentes, quas possessuri estis, deos suos super montes excelsos et colles et subter omne lignum frondosum.
DEUT|12|3|Dissipate aras eorum et confringite lapides, palos igne comburite et idola comminuite, disperdite nomina eorum de locis illis.
DEUT|12|4|Non facietis ita Domino Deo vestro.
DEUT|12|5|Sed ad locum, quem elegerit Dominus Deus vester de cunctis tribubus vestris, ut ponat nomen suum ibi et habitet in eo, venietis
DEUT|12|6|et offeretis in illo loco holocausta et victimas vestras, decimas et donaria manuum vestrarum et vota atque dona, primogenita boum et ovium.
DEUT|12|7|Et comedetis ibi in conspectu Domini Dei vestri ac laetabimini in cunctis, ad quae miseritis manum vos et domus vestrae, in quibus benedixerit vobis Dominus Deus vester.
DEUT|12|8|Non facietis secundum omnia, quae nos hic facimus hodie, singuli, quod sibi rectum videtur;
DEUT|12|9|neque enim usque in praesens tempus venistis ad requiem et possessionem, quam Dominus Deus vester daturus est vobis.
DEUT|12|10|Transibitis Iordanem et habitabitis in terra, quam Dominus Deus vester daturus est vobis, ut requiescatis a cunctis hostibus per circuitum et absque ullo timore habitetis
DEUT|12|11|in loco, quem elegerit Dominus Deus vester, ut habitet nomen eius in eo. Illuc omnia, quae praecipio, conferetis: holocausta et hostias ac decimas et donaria manuum vestrarum et, quidquid praecipuum est in muneribus, quae vovebitis Domino.
DEUT|12|12|Ibi laetabimini coram Domino Deo vestro vos, filii ac filiae vestrae, famuli et famulae atque Levites, qui in urbibus vestris commoratur; neque enim habet partem et possessionem inter vos.
DEUT|12|13|Cave, ne offeras holocausta tua in omni loco, quem videris,
DEUT|12|14|sed in eo, quem elegerit Dominus in una tribuum tuarum, offeres holocausta et ibi facies quaecumque praecipio tibi.
DEUT|12|15|Sin autem comedere volueris, et te esus carnium delectaverit, occide et comede carnem iuxta benedictionem Domini Dei tui, quam dedit tibi in omnibus urbibus tuis; sive immundus sive mundus comedet illam, sicut capream et cervum,
DEUT|12|16|absque esu dumtaxat sanguinis, quem super terram quasi aquam effundes.
DEUT|12|17|Non poteris comedere in oppidis tuis decimam frumenti et vini et olei tui, primogenita armentorum et pecorum et omnia, quae voveris et sponte offerre volueris, et primitiva manuum tuarum.
DEUT|12|18|Sed coram Domino Deo tuo comedes ea in loco, quem elegerit Dominus Deus tuus, tu et filius tuus ac filia tua, servus et famula atque Levites, qui manet in urbibus tuis; et laetaberis coram Domino Deo tuo in cunctis, ad quae extenderis manum tuam.
DEUT|12|19|Cave, ne derelinquas Levitem omni tempore, quo versaris in terra tua.
DEUT|12|20|Quando dilataverit Dominus Deus tuus terminos tuos, sicut locutus est tibi, et volueris vesci carnibus, quas desiderat anima tua, comedes carnem secundum omne desiderium animae tuae;
DEUT|12|21|locus autem, quem elegerit Dominus Deus tuus, ut sit nomen eius ibi, si procul fuerit, occides de armentis et pecoribus, quae dederit tibi Dominus, sicut praecepi tibi, et comedes in oppidis tuis, ut tibi placet.
DEUT|12|22|Sicut comeditur caprea et cervus, ita vesceris eis; et mundus et immundus in commune vescentur.
DEUT|12|23|Hoc solum cave, ne sanguinem comedas; sanguis enim eorum anima est, et idcirco non debes animam comedere cum carnibus.
DEUT|12|24|Non comedes eum, sed super terram fundes quasi aquam;
DEUT|12|25|non comedes eum, ut bene sit tibi et filiis tuis post te, cum feceris, quod placet in conspectu Domini.
DEUT|12|26|Quae autem sanctificaveris et voveris Domino, tolles et venies ad locum, quem elegerit Dominus,
DEUT|12|27|et offeres holocausta tua, carnem et sanguinem super altare Domini Dei tui; sanguis hostiarum tuarum fundetur in altari, carnibus autem ipse vesceris.
DEUT|12|28|Observa et audi omnia, quae ego praecipio tibi, ut bene sit tibi et filiis tuis post te in sempiternum, cum feceris, quod bonum est et placitum in conspectu Domini Dei tui.
DEUT|12|29|Quando disperdiderit Dominus Deus tuus ante faciem tuam gentes, ad quas ingredieris possidendas, et possederis eas atque habitaveris in terra earum,
DEUT|12|30|cave, ne irretiaris per eas, postquam te fuerint introeunte subversae, et requiras caeremonias earum dicens: "Sicut coluerunt gentes istae deos suos, ita et ego colam".
DEUT|12|31|Non facies similiter Domino Deo tuo; omnes enim abominationes, quas aversatur Dominus, fecerunt diis suis offerentes etiam filios et filias et comburentes igne.
DEUT|13|1|Quod praecipio vobis, hoc custodite et facite, nec addas quidquam nec minuas.
DEUT|13|2|Si surrexerit in medio tui prophetes aut, qui somnium vidisse se dicat, et dederit tibi signum vel portentum,
DEUT|13|3|et evenerit, quod locutus est, et dixerit tibi: "Eamus et sequamur deos alienos, quos ignoras, et serviamus eis",
DEUT|13|4|non audies verba prophetae illius aut somniatoris, quia tentat vos Dominus Deus vester, ut sciat utrum diligatis eum an non in toto corde et in tota anima vestra.
DEUT|13|5|Dominum Deum vestrum sequimini et ipsum timete et mandata illius custodite et audite vocem eius; ipsi servietis et ipsi adhaerebitis.
DEUT|13|6|Propheta autem ille aut fictor somniorum interficietur, quia locutus est, ut vos averteret a Domino Deo vestro, qui eduxit vos de terra Aegypti et redemit te de domo servitutis; ut errare te faceret de via, quam tibi praecepit Dominus Deus tuus; et auferes malum de medio tui.
DEUT|13|7|Si tibi voluerit persuadere frater tuus filius matris tuae aut filius tuus vel filia sive uxor, quae est in sinu tuo, aut amicus, quem diligis ut animam tuam, clam dicens: "Eamus et serviamus diis alienis", quos ignorasti tu et patres tui,
DEUT|13|8|de diis cunctarum in circuitu gentium, quae iuxta vel procul sunt ab initio usque ad finem terrae,
DEUT|13|9|non acquiescas ei nec audias, neque parcat ei oculus tuus, ut miserearis et occultes eum,
DEUT|13|10|sed interficies. Sit primum manus tua super eum, et postea omnis populus mittat manum:
DEUT|13|11|lapidibus obrutus necabitur, quia voluit te abstrahere a Domino Deo tuo, qui eduxit te de terra Aegypti, de domo servitutis,
DEUT|13|12|ut omnis Israel audiens timeat, et nequaquam ultra faciat quippiam huius rei simile in medio tui.
DEUT|13|13|Si audieris in una urbium tuarum, quas Dominus Deus tuus dabit tibi ad habitandum, dicentes aliquos:
DEUT|13|14|"Egressi sunt filii Belial de medio tui et averterunt habitatores urbis suae atque dixerunt: Eamus et serviamus diis alienis", quos ignorastis,
DEUT|13|15|quaere sollicite et, diligenter rei veritate perspecta, si inveneris certum esse, quod dicitur, et abominationem hanc opere perpetratam in medio tui,
DEUT|13|16|percuties habitatores urbis illius in ore gladii et delebis eam ac omnia, quae in illa sunt.
DEUT|13|17|Quidquid etiam supellectilis fuerit, congregabis in medio platearum eius et cum ipsa civitate succendes, ita ut universa consumas Domino Deo tuo, et sit tumulus sempiternus: non aedificabitur amplius.
DEUT|13|18|Et non adhaerebit de illo anathemate quidquam in manu tua, ut avertatur Dominus ab ira furoris sui et misereatur tui multiplicetque te, sicut iuravit patribus tuis,
DEUT|13|19|quando audieris vocem Domini Dei tui custodiens omnia mandata eius, quae ego praecipio tibi hodie, ut facias quod placitum est in conspectu Domini Dei tui.
DEUT|14|1|Filii estote Domini Dei ve stri; non vos incidetis nec fa cietis calvitium inter oculos vestros super mortuo,
DEUT|14|2|quoniam populus sanctus es Domino Deo tuo, et te elegit, ut sis ei in populum peculiarem de cunctis gentibus, quae sunt super terram.
DEUT|14|3|Ne comedatis quidquid abominabile est.
DEUT|14|4|Hoc est animal, quod comedere potestis: bovem et ovem et capram,
DEUT|14|5|cervum et capream, bubalum, tragelaphum, pygargum, orygem, rupicapram.
DEUT|14|6|Omne animal inter pecora, quod findit ungulam plene in duas partes et ruminat, comedetis;
DEUT|14|7|de his autem, quae ruminant et ungulam non findunt, haec comedere non debetis: camelum, leporem, hyracem, quia ruminant et non dividunt ungulam, immunda erunt vobis.
DEUT|14|8|Sus quoque, quoniam dividit ungulam et non ruminat, immunda erit vobis: carnibus eorum non vescemini et cadavera non tangetis.
DEUT|14|9|Haec comedetis ex omnibus, quae morantur in aquis: quae habent pinnulas et squamas comedite;
DEUT|14|10|quae absque pinnulis et squamis sunt, ne comedatis, quia immunda sunt vobis.
DEUT|14|11|Omnes aves mundas comedite;
DEUT|14|12|has autem ne comedatis: aquilam scilicet et grypem et alietum,
DEUT|14|13|ixon et vulturem ac milvum iuxta genus suum
DEUT|14|14|et omne corvini generis,
DEUT|14|15|struthionem ac noctuam et larum atque accipitrem iuxta genus suum,
DEUT|14|16|bubonem ac cycnum et ibin
DEUT|14|17|ac mergulum, porphyrionem et nycticoracem,
DEUT|14|18|erodium et charadrium, singula in genere suo, upupam quoque et vespertilionem.
DEUT|14|19|Et omne, quod reptat et pinnulas habet, immundum erit vobis, nec comedetur.
DEUT|14|20|Omne volatile, quod mundum est, comedite.
DEUT|14|21|Quidquid morticinum est, ne vescamini ex eo; advenae, qui intra portas tuas est, da, ut comedat, aut vende peregrino: quia tu populus sanctus es Domino Deo tuo.Non coques haedum in lacte matris suae.
DEUT|14|22|Decimam partem separabis de cunctis frugibus seminis tui, quae nascuntur in terra per annos singulos;
DEUT|14|23|et comedes in conspectu Domini Dei tui in loco, quem elegerit, ut in eo nomen illius habitet, decimam frumenti tui et vini et olei et primogenita de armentis et ovibus tuis, ut discas timere Dominum Deum tuum omni tempore.
DEUT|14|24|Cum autem longior fuerit tibi via et locus, quem elegerit Dominus Deus tuus, ut ponat nomen suum ibi tibique benedixerit, nec potueris ad eum haec cuncta portare,
DEUT|14|25|vendes omnia et in pretium rediges; portabisque manu tua et proficisceris ad locum, quem elegerit Dominus Deus tuus,
DEUT|14|26|et emes ex eadem pecunia, quidquid tibi placuerit, sive ex armentis sive ex ovibus, vinum quoque et siceram et omne, quod desiderat anima tua; et comedes ibi coram Domino Deo tuo et epulaberis tu et domus tua
DEUT|14|27|et Levites, qui intra portas tuas est: cave, ne derelinquas eum, quia non habet partem nec possessionem tecum.
DEUT|14|28|Anno tertio separabis aliam decimam ex omnibus, quae nascuntur tibi eo tempore, et repones intra portas tuas;
DEUT|14|29|venietque Levites, qui non habet partem nec possessionem tecum, et peregrinus ac pupillus ac vidua, qui intra portas tuas sunt, et comedent et saturabuntur, ut benedicat tibi Dominus Deus tuus in cunctis operibus manuum tuarum, quae feceris.
DEUT|15|1|Septimo anno facies remis sionem,
DEUT|15|2|quae hoc ordine ce lebrabitur: cui debetur aliquid a proximo ac fratre suo, repetere non poterit, quia annus remissionis est Domino.
DEUT|15|3|A peregrino exiges; civem et propinquum repetendi, quod tuum est, non habebis potestatem.
DEUT|15|4|Sed omnino indigens non erit apud te, quia benedicet tibi Dominus Deus tuus in terra, quam traditurus est tibi in possessionem,
DEUT|15|5|si tamen audieris vocem Domini Dei tui et custodieris universum mandatum hoc, quod ego hodie praecipio tibi,
DEUT|15|6|quia Dominus Deus tuus benedicet tibi, ut pollicitus est. Fenerabis gentibus multis et ipse a nullo accipies mutuum; dominaberis nationibus plurimis, et tui nemo dominabitur.
DEUT|15|7|Si unus de fratribus tuis, qui morantur in una civitatum tuarum in terra, quam Dominus Deus tuus daturus est tibi, ad paupertatem venerit, non obdurabis cor tuum nec contrahes manum;
DEUT|15|8|sed aperies eam pauperi fratri tuo et dabis mutuum, quod eum indigere perspexeris.
DEUT|15|9|Cave, ne forte subrepat tibi impia cogitatio, et dicas in corde tuo: Appropinquat septimus annus remissionis", et avertas oculos tuos a paupere fratre tuo nolens ei, quod postulat, mutuum commodare, ne clamet contra te ad Dominum, et fiat tibi in peccatum.
DEUT|15|10|Sed dabis ei, nec contristabitur cor tuum in eius necessitatibus sublevandis, nam propter hoc benedicet tibi Dominus Deus tuus in omni opere tuo et in cunctis, ad quae manum miseris.
DEUT|15|11|Non deerunt pauperes in terra habitationis tuae; idcirco ego praecipio tibi, ut aperias manum fratri tuo egeno et pauperi, qui tecum versatur in terra tua.
DEUT|15|12|Cum tibi venditus fuerit frater tuus Hebraeus aut Hebraea et sex annis servierit tibi, in septimo anno dimittes eum liberum;
DEUT|15|13|et quem libertate donaveris, nequaquam vacuum abire patieris.
DEUT|15|14|Sed dabis ei viaticum de gregibus et de area et torculari tuo, quibus Dominus Deus tuus benedixerit tibi.
DEUT|15|15|Memento quod et ipse servieris in terra Aegypti, et liberaverit te Dominus Deus tuus; idcirco ego nunc hoc praecipio tibi.
DEUT|15|16|Sin autem dixerit: "Nolo egredi", eo quod diligat te et domum tuam et bene sibi apud te esse sentiat,
DEUT|15|17|assumes subulam et perforabis aurem eius in ianua domus tuae, et serviet tibi usque in aeternum. Ancillae quoque similiter facies.
DEUT|15|18|Non sit durum in oculis tuis dimittere eum liberum, quoniam iuxta mercedem mercennarii per sex annos servivit tibi, et benedicet tibi Dominus Deus tuus in cunctis operibus, quae egeris.
DEUT|15|19|De primogenitis, quae nascuntur in armentis et ovibus tuis, quidquid sexus est masculini, sanctificabis Domino Deo tuo; non operaberis in primogenito bovis et non tondebis primogenita ovium.
DEUT|15|20|In conspectu Domini Dei tui comedes ea per annos singulos in loco, quem elegerit Dominus, tu et domus tua.
DEUT|15|21|Sin autem habuerit maculam et vel claudum fuerit vel caecum aut in aliqua parte deforme vel debile, non immolabis illud Domino Deo tuo,
DEUT|15|22|sed intra portas tuas comedes illud; tam mundus quam immundus similiter vescentur eis, quasi caprea et cervo.
DEUT|15|23|Solum sanguinem eorum non comedes, sed effundes in terram quasi aquam.
DEUT|16|1|Observa mensem Abib, ut facias Pascha Domino Deo tuo; quoniam in isto mense Abib eduxit te Dominus Deus tuus de Aegypto nocte.
DEUT|16|2|Immolabisque Pascha Domino Deo tuo de ovibus et de bobus in loco, quem elegerit Dominus Deus tuus, ut habitet nomen eius ibi.
DEUT|16|3|Non comedes cum eo panem fermentatum; septem diebus comedes absque fermento afflictionis panem, quoniam festinanter egressus es de Aegypto, ut memineris diei egressionis tuae de Aegypto omnibus diebus vitae tuae.
DEUT|16|4|Non apparebit fermentum in omnibus terminis tuis septem diebus; et non manebit de carnibus eius, quod immolatum est vespere in die primo, usque mane.
DEUT|16|5|Non poteris immolare Pascha in qualibet urbium tuarum, quas Dominus Deus tuus daturus est tibi,
DEUT|16|6|sed in loco, quem elegerit Dominus Deus tuus, ut habitet nomen eius ibi, immolabis Pascha vespere ad solis occasum, quando egressus es de Aegypto.
DEUT|16|7|Et coques et comedes in loco, quem elegerit Dominus Deus tuus, maneque consurgens vades in tabernacula tua.
DEUT|16|8|Sex diebus comedes azyma et in die septimo, quia collecta est Domino Deo tuo, non facies opus.
DEUT|16|9|Septem hebdomadas numerabis tibi ab ea die, qua falcem in segetem miseris,
DEUT|16|10|et celebrabis diem festum Hebdomadarum Domino Deo tuo, oblationem spontaneam manus tuae, quam offeres iuxta benedictionem Domini Dei tui.
DEUT|16|11|Et epulaberis coram Domino Deo tuo tu, filius tuus et filia tua, servus tuus et ancilla tua et Levites, qui est intra portas tuas, advena ac pupillus et vidua, qui morantur tecum in loco, quem elegerit Dominus Deus tuus, ut habitet nomen eius ibi;
DEUT|16|12|et recordaberis quoniam servus fueris in Aegypto custodiesque ac facies, quae praecepta sunt.
DEUT|16|13|Sollemnitatem quoque Tabernaculorum celebrabis per septem dies, quando collegeris de area et torculari fruges tuas;
DEUT|16|14|et epulaberis in festivitate tua tu, filius tuus et filia, servus tuus et ancilla, Levites quoque et advena, pupillus ac vidua, qui intra portas tuas sunt.
DEUT|16|15|Septem diebus Domino Deo tuo festa celebrabis in loco, quem elegerit Dominus, quia benedicet tibi Dominus Deus tuus in cunctis frugibus tuis et in omni opere manuum tuarum, erisque totus in laetitia.
DEUT|16|16|Tribus vicibus per annum apparebit omne masculinum tuum in conspectu Domini Dei tui in loco, quem elegerit: in sollemnitate Azymorum et in sollemnitate Hebdomadarum et in sollemnitate Tabernaculorum. Non apparebit ante Dominum vacuus,
DEUT|16|17|sed offeret unusquisque secundum quod habuerit, iuxta benedictionem Domini Dei tui, quam dederit tibi.
DEUT|16|18|Iudices et praefectos operum constitues in omnibus portis tuis, quas Dominus Deus tuus dederit tibi per singulas tribus tuas, ut iudicent populum iusto iudicio.
DEUT|16|19|Non declinabis iudicium. Non accipies personam nec munera, quia munera excaecant oculos sapientum et mutant causas iustorum.
DEUT|16|20|Iustitiam, iustitiam persequeris, ut vivas et possideas terram, quam Dominus Deus tuus dederit tibi.
DEUT|16|21|Non plantabis tibi palum, omnem arborem iuxta altare Domini Dei tui, quod feceris tibi.
DEUT|16|22|Neque constitues lapidem, quem odit Dominus Deus tuus.
DEUT|17|1|Non immolabis Domino Deo tuo ovem et bovem, in quo est macula aut quippiam vitii, quia abominatio est Domino Deo tuo.
DEUT|17|2|Cum reperti fuerint apud te intra unam portarum tuarum, quas Dominus Deus tuus dabit tibi, vir aut mulier, qui faciant, quod malum est in conspectu Domini Dei tui, et transgrediantur pactum illius,
DEUT|17|3|ut vadant et serviant diis alienis et adorent eos, solem vel lunam vel omnem militiam caeli, quae non praecepi,
DEUT|17|4|et hoc tibi fuerit nuntiatum, audiensque inquisieris diligenter et verum esse reppereris, et abominatio haec facta est in Israel,
DEUT|17|5|educes virum vel mulierem, qui hanc rem sceleratissimam perpetrarunt, ad portas civitatis tuae, et lapidibus obruentur.
DEUT|17|6|In ore duorum aut trium testium peribit, qui interficietur; nemo occidatur uno contra se dicente testimonium.
DEUT|17|7|Manus testium prima erit ad interficiendum eum, et manus reliqui populi extrema mittetur, ut auferas malum de medio tui.
DEUT|17|8|Si intra portas tuas in litibus difficile et ambiguum apud te iudicium esse perspexeris inter sanguinem et sanguinem, causam et causam, plagam et plagam, surge et ascende ad locum, quem elegerit Dominus Deus tuus,
DEUT|17|9|veniesque ad sacerdotes levitici generis et ad iudicem, qui fuerit illo tempore; quaeresque ab eis, qui indicabunt tibi iudicii sententiam.
DEUT|17|10|Et facies quodcumque dixerint tibi de loco, quem elegerit Dominus, et observabis, ut facias omnia quae docuerint te
DEUT|17|11|iuxta mandatum, quod mandaverunt, et iuxta sententiam, quam dixerint tibi. Nec declinabis ad dexteram vel ad sinistram.
DEUT|17|12|Qui autem superbierit nolens oboedire sacerdotis imperio, qui eo tempore ministrat Domino Deo tuo, aut decreto iudicis, morietur homo ille, et auferes malum de Israel;
DEUT|17|13|cunctusque populus audiens timebit, ut nullus deinceps intumescat superbia.
DEUT|17|14|Cum ingressus fueris terram, quam Dominus Deus tuus dabit tibi, et possederis eam habitaverisque in illa et dixeris: "Constituam super me regem, sicut habent omnes per circuitum nationes",
DEUT|17|15|eum constitues super te regem, quem Dominus Deus tuus elegerit de numero fratrum tuorum. Non poteris alterius gentis hominem regem facere, qui non sit frater tuus.
DEUT|17|16|Tantummodo non multiplicabit sibi equos nec reducet populum in Aegyptum, ut equitatus numerum augeat, praesertim cum Dominus praeceperit vobis, ut nequaquam amplius per hanc viam revertamini.
DEUT|17|17|Neque habebit uxores plurimas, ne declinet cor eius, neque argenti et auri immensa pondera.
DEUT|17|18|Postquam autem sederit in solio regni sui, describet sibi exemplar legis huius in volumine accipiens illam a sacerdotibus leviticae tribus;
DEUT|17|19|et habebit secum legetque illud omnibus diebus vitae suae, ut discat timere Dominum Deum suum. et custodire verba legis huius et praecepta ista et quae in lege praecepta sunt.
DEUT|17|20|Nec elevetur cor eius in superbiam super fratres suos neque declinet a mandatis in partem dexteram vel sinistram, ut longo tempore regnet ipse et filii eius in medio Israel.
DEUT|18|1|Non habebunt sacerdotes le vitae, omnis tribus Levi, par tem et hereditatem cum reliquo Israel; de sacrificiis Domini et hereditate eius comedent
DEUT|18|2|et nihil accipient de possessione fratrum suorum: Dominus enim ipse est hereditas eorum, sicut locutus est illis.
DEUT|18|3|Hoc erit ius sacerdotum a populo, ab his qui offerunt victimas: sive bovem sive ovem immolaverint, dabunt sacerdoti armum et duas maxillas ac ventriculum,
DEUT|18|4|primitias frumenti, vini et olei et lanarum ex ovium tonsione.
DEUT|18|5|Ipsum enim elegit Dominus Deus tuus de cunctis tribubus tuis, ut stet et ministret in nomine Domini ipse et filii eius in sempiternum.
DEUT|18|6|Si exierit Levites de una urbium tuarum ex omni Israel, in qua ut advena habitat, et voluerit venire desiderans locum, quem elegerit Dominus,
DEUT|18|7|ministrabit in nomine Domini Dei sui, sicut omnes fratres eius levitae, qui stabunt ibi coram Domino.
DEUT|18|8|Partem ciborum eandem accipiet quam et ceteri, excepto eo, quod ex paterna ei successione debetur.
DEUT|18|9|Quando ingressus fueris terram, quam Dominus Deus tuus dabit tibi, cave, ne imitari velis abominationes illarum gentium.
DEUT|18|10|Nec inveniatur in te, qui filium suum aut filiam traducat per ignem, aut qui sortes sciscitetur et observet nubes atque auguria, nec sit maleficus
DEUT|18|11|nec incantator, nec qui pythones consulat nec divinos, aut quaerat a mortuis veritatem;
DEUT|18|12|omnia enim haec abominatur Dominus et propter istiusmodi scelera expellet eos in introitu tuo.
DEUT|18|13|Perfectus eris et absque macula cum Domino Deo tuo.
DEUT|18|14|Gentes istae, quarum possidebis terram, augures et divinos audiunt; tu autem a Domino Deo tuo aliter institutus es.
DEUT|18|15|Prophetam de gente tua et de fratribus tuis sicut me suscitabit tibi Dominus Deus tuus; ipsum audietis,
DEUT|18|16|ut petiisti a Domino Deo tuo in Horeb, quando contio congregata est, atque dixisti: "Ultra non audiam vocem Domini Dei mei et ignem hunc maximum amplius non videbo, ne moriar".
DEUT|18|17|Et ait Dominus mihi: "Bene omnia sunt locuti;
DEUT|18|18|prophetam suscitabo eis de medio fratrum suorum similem tui et ponam verba mea in ore eius, loqueturque ad eos omnia, quae praecepero illi.
DEUT|18|19|Qui autem verba mea, quae loquetur in nomine meo, audire noluerit, ego ultor exsistam.
DEUT|18|20|Propheta autem qui, arrogantia depravatus, voluerit loqui in nomine meo, quae ego non praecepi illi ut diceret, aut ex nomine alienorum deorum, interficietur".
DEUT|18|21|Quod si tacita cogitatione responderis: "Quomodo possum intellegere verbum, quod Dominus non est locutus?",
DEUT|18|22|hoc habebis signum: quod in nomine Domini propheta ille praedixerit, et non evenerit, hoc Dominus non est locutus, sed per tumorem animi sui propheta confinxit; et idcirco non timebis eum.
DEUT|19|1|Cum disperderit Dominus Deus tuus gentes, quarum ti bi traditurus est terram, et possederis eam habitaverisque in urbibus eius et in aedibus,
DEUT|19|2|tres civitates separabis tibi in medio terrae, quam Dominus Deus tuus dabit tibi in possessionem
DEUT|19|3|sternens diligenter viam; et in tres aequaliter partes totam terrae tuae provinciam divides, ut habeat e vicino, qui propter homicidium profugus est, quo possit evadere.
DEUT|19|4|Haec erit lex homicidae fugientis, cuius vita servanda est: qui percusserit proximum suum nesciens et qui heri et nudiustertius nullum contra eum habuisse odium comprobatur,
DEUT|19|5|sed abiisse cum eo simpliciter in silvam ad ligna caedenda, et in succisione lignorum securis fugerit manu, ferrumque lapsum de manubrio amicum eius percusserit et occiderit, hic ad unam supradictarum urbium confugiet et vivet;
DEUT|19|6|ne forsitan ultor sanguinis cordis calore stimulatus persequatur et apprehendat eum, si longior via fuerit, et percutiat eum, et moriatur, qui non est reus mortis, quia nullum contra eum, qui occisus est, odium prius habuisse monstratur.
DEUT|19|7|Idcirco praecipio tibi, ut tres civitates aequalis inter se spatii dividas.
DEUT|19|8|Cum autem dilataverit Dominus Deus tuus terminos tuos, sicut iuravit patribus tuis, et dederit tibi cunctam terram, quam eis pollicitus est
DEUT|19|9|- si tamen custodieris omne mandatum hoc et feceris, quae hodie praecipio tibi, ut diligas Dominum Deum tuum et ambules in viis eius omni tempore - addes tibi tres alias civitates et supradictarum trium urbium numerum duplicabis,
DEUT|19|10|ut non effundatur sanguis innoxius in medio terrae, quam Dominus Deus tuus dabit tibi possidendam, nec sis sanguinis reus.
DEUT|19|11|Si quis autem odio habens proximum suum insidiatus fuerit vitae eius surgensque percusserit illum, et mortuus fuerit, fugeritque ad unam de supradictis urbibus,
DEUT|19|12|mittent seniores civitatis eius et arripient eum de loco effugii tradentque in manu ultoris sanguinis, et morietur:
DEUT|19|13|non misereberis eius et auferes innoxium sanguinem de Israel, ut bene sit tibi.
DEUT|19|14|Non transferes terminos proximi tui, quos fixerunt priores in possessione tua, quam acceperis in terra, quam Dominus Deus tuus dabit tibi possidendam.
DEUT|19|15|Non stabit testis unus contra aliquem, quidquid illius peccatum vel facinus fuerit; sed in ore duorum aut trium testium stabit omne verbum.
DEUT|19|16|Si steterit testis mendax contra hominem accusans eum praevaricationis,
DEUT|19|17|stabunt ambo, quorum causa est, ante Dominum in conspectu sacerdotum et iudicum, qui fuerint in diebus illis.
DEUT|19|18|Cumque diligentissime perscrutantes iudices invenerint falsum testem dixisse contra fratrem suum mendacium,
DEUT|19|19|reddent ei, sicut fratri suo facere cogitavit, et auferes malum de medio tui,
DEUT|19|20|ut audientes ceteri timorem habeant et nequaquam ultra talia audeant facere in medio tui.
DEUT|19|21|Non misereberis eius, sed animam pro anima, oculum pro oculo, dentem pro dente, manum pro manu, pedem pro pede exiges.
DEUT|20|1|Si exieris ad bellum contra hostes tuos et videris equita tus et currus et maiorem, quam tu habes, adversarii exercitus multitudinem, non timebis eos, quia Dominus Deus tuus tecum est, qui eduxit te de terra Aegypti.
DEUT|20|2|Appropinquante autem iam proelio, stabit sacerdos ante aciem et sic loquetur ad populum:
DEUT|20|3|"Audi, Israel: Vos hodie contra inimicos vestros pugnam committitis; non pertimescat cor vestrum, nolite metuere, nolite cedere nec formidetis eos,
DEUT|20|4|quia Dominus Deus vester incedit vobiscum et pro vobis contra adversarios vestros dimicabit, ut eruat vos de periculo".
DEUT|20|5|Praefecti quoque per singulas turmas, audiente exercitu, proclamabunt: Quis est homo, qui aedificavit domum novam et non dedicavit eam? Vadat et revertatur in domum suam, ne forte moriatur in bello, et alius dedicet illam.
DEUT|20|6|Quis est homo, qui plantavit vineam et necdum vindemiavit eam? Vadat et revertatur in domum suam, ne forte moriatur in bello, et alius homo vindemiet illam.
DEUT|20|7|Quis est homo, qui despondit uxorem et non accepit eam? Vadat et revertatur in domum suam, ne forte moriatur in bello, et alius homo accipiat eam".
DEUT|20|8|His dictis, addent reliqua et loquentur ad populum: "Quis est homo formidulosus et corde pavido? Vadat et revertatur in domum suam, ne pavere faciat corda fratrum suorum, sicut ipse timore perterritus est".
DEUT|20|9|Cumque praefecti finem loquendi ad populum fecerint, constituantur duces exercitus in capite populi.
DEUT|20|10|Si quando accesseris ad expugnandam civitatem, offeres ei primum pacem;
DEUT|20|11|si receperit et aperuerit tibi portas, cunctus populus, qui in ea est, serviet tibi sub tributo.
DEUT|20|12|Sin autem foedus inire noluerit et coeperit contra te bellum, oppugnabis eam.
DEUT|20|13|Cumque tradiderit Dominus Deus tuus illam in manu tua, percuties omne, quod in ea generis masculini est, in ore gladii
DEUT|20|14|absque mulieribus et infantibus, iumentis et ceteris, quae in civitate sunt. Omnem praedam hanc diripies tibi et comedes de spoliis hostium tuorum, quae Dominus Deus tuus dederit tibi.
DEUT|20|15|Sic facies cunctis civitatibus, quae a te procul valde sunt et non sunt de gentium istarum urbibus, quas in possessionem accepturus es.
DEUT|20|16|De his autem civitatibus, quae dabuntur tibi, nullum omnino permittes vivere,
DEUT|20|17|sed interficies in ore gladii, Hetthaeum videlicet et Amorraeum et Chananaeum, Pherezaeum et Hevaeum et Iebusaeum, sicut praecepit tibi Dominus Deus tuus,
DEUT|20|18|ne forte doceant vos facere cunctas abominationes, quas ipsi operati sunt diis suis, et peccetis in Dominum Deum vestrum.
DEUT|20|19|Quando obsederis civitatem multo tempore et munitionibus circumdederis, ut expugnes eam, non immittes securim in arbores eius, de quibus vesci potes, nec succidas eas. Numquid homo est arbor campi, ut eam obsideas?
DEUT|20|20|Si qua autem ligna non sunt pomifera, succide illa et exstrue machinas, donec capias civitatem, quae contra te dimicat.
DEUT|21|1|Quando inventum fuerit in terra, quam Dominus Deus tuus daturus est tibi, hominis cadaver occisi, et ignoratur caedis reus,
DEUT|21|2|egredientur maiores natu et iudices tui et metientur a loco cadaveris singularum per circuitum spatia civitatum
DEUT|21|3|et, quam viciniorem ceteris esse perspexerint, seniores civitatis illius tollent vitulam de armento, quae non traxit iugum nec terram scidit vomere,
DEUT|21|4|et ducent eam ad torrentem perennem, ubi numquam aratum est nec seminatum, et caedent apud eum cervices vitulae;
DEUT|21|5|accedentque sacerdotes filii Levi, quos elegerit Dominus Deus tuus, ut ministrent ei et benedicant in nomine eius, et ad verbum eorum omnis causa et omnis percussio iudicetur.
DEUT|21|6|Et omnes maiores natu civitatis illius, qui prope interfectum sunt, lavabunt manus suas super vitulam, quae apud torrentem percussa est,
DEUT|21|7|et dicent: "Manus nostrae non effuderunt hunc sanguinem, nec oculi nostri viderunt;
DEUT|21|8|propitius esto populo tuo Israel, quem redemisti, Domine, et non reputes sanguinem innocentem in medio populi tui Israel". Et auferetur ab eis reatus sanguinis.
DEUT|21|9|Tu autem removebis innocentem cruorem, cum feceris, quod rectum est in oculis Domini.
DEUT|21|10|Si egressus fueris ad pugnam contra inimicos tuos, et tradiderit eos Dominus Deus tuus in manu tua, captivosque duxeris
DEUT|21|11|et videris in numero captivorum mulierem pulchram et adamaveris eam voluerisque habere uxorem,
DEUT|21|12|introduces eam in domum tuam. Quae radet caesariem et circumcidet ungues
DEUT|21|13|et deponet vestem captivitatis sedensque in domo tua flebit patrem et matrem suam uno mense; et postea intrabis ad eam sociaberisque illi, et erit uxor tua.
DEUT|21|14|Sin autem postea non sederit animo tuo, dimittes eam liberam; nec vendere poteris pecunia nec opprimere per potentiam, quia humiliasti eam.
DEUT|21|15|Si habuerit homo uxores duas, unam dilectam et alteram odiosam, genuerintque ei liberos, et fuerit filius odiosae primogenitus,
DEUT|21|16|volueritque substantiam inter filios suos dividere, non poterit filium dilectae facere primogenitum et praeferre filio odiosae,
DEUT|21|17|sed filium odiosae agnoscet primogenitum dabitque ei de cunctis, quae habuerit, duplicia; iste est enim principium roboris eius, et huic debentur primogenita.
DEUT|21|18|Si genuerit homo filium contumacem et protervum, qui non audiat patris aut matris imperium et coercitus oboedire contempserit,
DEUT|21|19|apprehendent eum et ducent ad seniores civitatis suae et ad portam iudicii
DEUT|21|20|dicentque ad eos: "Filius noster iste protervus et contumax est: monita nostra audire contemnit, comissationibus vacat et luxuriae atque conviviis potatorum".
DEUT|21|21|Lapidibus eum obruent viri civitatis, et morietur, ut auferatis malum de medio vestri, et universus Israel audiens pertimescat.
DEUT|21|22|Quando peccaverit homo, quod morte plectendum est, et occisum appenderis in patibulo,
DEUT|21|23|non permanebit cadaver eius in ligno; sed in eadem die sepelietur, quia maledictus a Deo est, qui pendet in ligno; et nequaquam contaminabis terram tuam, quam Dominus Deus tuus dederit tibi in possessionem.
DEUT|22|1|Non videbis bovem fratris tui aut ovem errantem et praeteribis, sed reduces fratri tuo;
DEUT|22|2|si autem non est prope frater tuus nec nosti eum, duces in domum tuam, et erunt apud te quamdiu quaerat ea frater tuus et recipiat.
DEUT|22|3|Similiter facies de asino et de vestimento et de omni re fratris tui, quae perierit: si inveneris eam, ne subtrahas te.
DEUT|22|4|Si videris asinum fratris tui aut bovem cecidisse in via, non subtrahes te, sed sublevabis cum eo.
DEUT|22|5|Non induetur mulier veste virili, nec vir utetur veste feminea: abominabilis enim apud Dominum Deum tuum est omnis, qui facit haec.
DEUT|22|6|Si ambulans per viam, in arbore vel in terra nidum avis inveneris et matrem pullis vel ovis desuper incubantem, non sumes eam de filiis,
DEUT|22|7|sed abire patieris matrem tenens filios, ut bene sit tibi, et longo vivas tempore.
DEUT|22|8|Cum aedificaveris domum novam, facies murum tecto tuo per circuitum, ne adducas sanguinem super domum tuam et sis reus, labente aliquo in praeceps ruente.
DEUT|22|9|Non seres vineam tuam altero semine, ne et sementis, quam sevisti, et quae nascuntur ex vinea, pariter sanctificentur.
DEUT|22|10|Non arabis in bove simul et asino.
DEUT|22|11|Non indueris vestimento, quod ex lana linoque contextum est.
DEUT|22|12|Funiculos facies per quattuor angulos pallii tui, quo operieris.
DEUT|22|13|Si duxerit vir uxorem et intraverit ad eam et postea odio habuerit eam
DEUT|22|14|imputaveritque ei obiciens ei nomen pessimum et dixerit: "Uxorem hanc accepi et ingressus ad eam non inveni virginem",
DEUT|22|15|tollent pater et mater eius et ferent secum signa virginitatis eius ad seniores urbis, qui in porta sunt,
DEUT|22|16|et dicet pater: "Filiam meam dedi huic uxorem, quam, quia odit,
DEUT|22|17|imponit ei nomen pessimum, ut dicat: Non inveni filiam tuam virginem; et ecce haec sunt signa virginitatis filiae meae". Expandent vestimentum coram se nioribus civitatis.
DEUT|22|18|Apprehendentque senes urbis illius virum et verberabunt illum
DEUT|22|19|condemnantes insuper centum siclis argenti, quos dabunt patri puellae, quoniam diffamavit nomen pessimum super virginem Israel; habebitque eam uxorem et non poterit dimittere eam omnibus diebus vitae suae.
DEUT|22|20|Quod si verum est, quod obicit, et non est in puella inventa virginitas,
DEUT|22|21|educent eam ad fores domus patris sui, et lapidibus obruent viri civitatis eius, et morietur, quoniam fecit nefas in Israel, ut fornicaretur in domo patris sui; et auferes malum de medio tui.
DEUT|22|22|Si inventus fuerit vir dormiens cum uxore alterius, uterque morietur, id est adulter et adultera; et auferes malum de Israel.
DEUT|22|23|Si puellam virginem desponsatam viro invenerit aliquis in civitate et concubuerit cum illa,
DEUT|22|24|educetis utrumque ad portam civitatis illius et lapidibus obruetis, et morientur: puella quia non clamavit, cum esset in civitate, vir quia humiliavit uxorem proximi sui; et auferes malum de medio tui.
DEUT|22|25|Sin autem in agro reppererit vir puellam, quae desponsata est, et apprehendens concubuerit cum illa, ipse morietur solus;
DEUT|22|26|puella nihil patietur nec est rea mortis, quoniam sicut vir consurgit contra fratrem suum et occidit eum, ita et puella perpessa est:
DEUT|22|27|sola erat in agro, clamavit puella desponsata, et nullus affuit, qui liberaret eam.
DEUT|22|28|Si invenerit vir puellam virginem, quae non habet sponsum, et apprehendens concubuerit cum ea, et res ad iudicium venerit,
DEUT|22|29|dabit, qui dormivit cum ea, patri puellae quinquaginta siclos argenti et habebit eam uxorem, quia humiliavit illam: non poterit dimittere eam cunctis diebus vitae suae.
DEUT|23|1|Non accipiet homo uxorem patris sui nec revelabit operi mentum eius.
DEUT|23|2|Non intrabit eunuchus, attritis vel amputatis testiculis et absciso veretro, ecclesiam Domini.
DEUT|23|3|Non ingredietur mamzer in ecclesiam Domini neque decima generatione.
DEUT|23|4|Ammonites et Moabites etiam in decima generatione non intrabunt ecclesiam Domini in aeternum,
DEUT|23|5|quia noluerunt vobis occurrere cum pane et aqua in via, quando egressi estis de Aegypto, et quia conduxerunt contra te Balaam filium Beor de Phethor in Aramnaharaim, ut malediceret tibi;
DEUT|23|6|et noluit Dominus Deus tuus audire Balaam vertitque tibi maledictionem eius in benedictionem, eo quod diligeret te.
DEUT|23|7|Non facies cum eis pacem nec quaeres eis bona cunctis diebus vitae tuae in sempiternum.
DEUT|23|8|Non abominaberis Idumaeum, quia frater tuus est, nec Aegyptium, quia advena fuisti in terra eius:
DEUT|23|9|qui nati fuerint ex eis tertia generatione, intrabunt ecclesiam Domini.
DEUT|23|10|Quando egressus fueris adversus hostes tuos in pugnam, custodies te ab omni re mala.
DEUT|23|11|Si fuerit apud te homo, qui nocturno pollutus sit somnio, egredietur extra castra et non revertetur,
DEUT|23|12|priusquam ad vesperam lavetur aqua; et ad solis occasum regredietur in castra.
DEUT|23|13|Habebis locum extra castra, ad quem egrediaris ad requisita naturae
DEUT|23|14|gerens paxillum in balteo; cumque sederis foris, fodies foveam et egesta humo operies.
DEUT|23|15|Dominus enim Deus tuus ambulat in medio castrorum tuorum, ut eruat te et tradat tibi inimicos tuos; sint castra tua sancta, et nihil in eis videat foeditatis nec derelinquat te.
DEUT|23|16|Non trades servum domino suo, qui ad te confugerit:
DEUT|23|17|habitabit tecum in medio tui in loco, quem elegerit in una urbium tuarum, quae placuerit ei, nec contristes eum.
DEUT|23|18|Non erit prostibulum sacrum de filiabus Israel, nec scortator sacer de filiis Israel.
DEUT|23|19|Non offeres mercedem prostibuli nec pretium canis in domo Domini Dei tui, quidquid illud est, quod voveris, quia abominatio est utrumque apud Dominum Deum tuum.
DEUT|23|20|Non fenerabis fratri tuo ad usuram pecuniam nec alimenta nec quamlibet aliam rem,
DEUT|23|21|sed alieno fenerabis. Fratri autem tuo absque usura id, quo indiget, commodabis, ut benedicat tibi Dominus Deus tuus in omni opere tuo in terra, ad quam ingredieris possidendam.
DEUT|23|22|Cum voveris votum Domino Deo tuo, non tardabis reddere; quia requiret illud Dominus Deus tuus a te, et reputabitur tibi in peccatum.
DEUT|23|23|Si nolueris polliceri, absque peccato eris;
DEUT|23|24|quod autem egressum est de labiis tuis, observabis et facies, sicut promisisti Domino Deo tuo: propria voluntate et ore tuo locutus es.
DEUT|23|25|Ingressus vineam proximi tui comede uvas, quantum tibi placuerit; in sporta autem ne efferas tecum.
DEUT|23|26|Si intraveris in segetem amici tui, franges spicas manu; falce autem non metes.
DEUT|24|1|Si acceperit homo uxorem et habuerit eam, et non invene rit gratiam ante oculos eius propter aliquam foeditatem, et scripserit libellum repudii dederitque in manu illius et dimiserit eam de domo sua,
DEUT|24|2|cumque egressa alterius uxor facta fuerit,
DEUT|24|3|et ille quoque oderit eam dederitque ei libellum repudii et dimiserit de domo sua, vel mortuus fuerit,
DEUT|24|4|non poterit prior maritus recipere eam in uxorem, quia polluta est; hoc esset abominatio coram Domino. Ne peccare facias terram tuam, quam Dominus Deus tuus tradiderit tibi possidendam.
DEUT|24|5|Cum acceperit homo nuper uxorem, non procedet ad bellum, nec ei quippiam necessitatis iniungetur publicae, sed vacabit liber domui suae, ut uno anno laetetur cum uxore sua.
DEUT|24|6|Non accipies loco pignoris molam vel superiorem lapidem molarem, quia animam suam apposuit tibi.
DEUT|24|7|Si deprehensus fuerit homo rapiens unum de fratribus suis de filiis Israel et, vendito eo, accipiens pretium, interficietur; et auferes malum de medio tui.
DEUT|24|8|Observa diligenter, si incurras plagam leprae, quaecumque docuerint vos sacerdotes levitici generis; quod praecepi eis, implete sollicite.
DEUT|24|9|Memento, quae fecerit Dominus Deus tuus Mariae in via, cum egrederemini de Aegypto.
DEUT|24|10|Cum mutuam dabis proximo tuo rem aliquam, non ingredieris domum eius, ut pignus auferas,
DEUT|24|11|sed stabis foris, et ille tibi pignus proferet, quod habuerit.
DEUT|24|12|Sin autem pauper est, non pernoctabit apud te pignus,
DEUT|24|13|sed statim reddes ei ad solis occasum, ut dormiens in vestimento suo benedicat tibi, et habeas iustitiam coram Domino Deo tuo.
DEUT|24|14|Non negabis mercedem indigentis et pauperis ex fratribus tuis sive advenis, qui tecum morantur in terra intra portas tuas,
DEUT|24|15|sed eadem die reddes ei pretium laboris sui ante solis occasum, quia pauper est, et illud desiderat anima sua; ne clamet contra te ad Dominum, et reputetur tibi in peccatum.
DEUT|24|16|Non occidentur patres pro filiis, nec filii pro patribus, sed unusquisque pro peccato suo morietur.
DEUT|24|17|Non pervertes iudicium advenae et pupilli nec auferes pignoris loco viduae vestimentum.
DEUT|24|18|Memento quod servieris in Aegypto, et eruerit te Dominus Deus tuus inde; idcirco praecipio tibi, ut facias hanc rem.
DEUT|24|19|Quando messueris segetem in agro tuo et oblitus manipulum reliqueris, non reverteris, ut tollas eum, sed advenam et pupillum et viduam auferre patieris, ut benedicat tibi Dominus Deus tuus in omni opere manuum tuarum.
DEUT|24|20|Si fruges collegeris olivarum, quidquid remanserit in arboribus, non reverteris, ut colligas, sed relinques advenae, pupillo ac viduae.
DEUT|24|21|Si vindemiaveris vineam tuam, non colliges remanentes racemos, sed cedent in usus advenae, pupilli ac viduae.
DEUT|24|22|Memento quod et tu servieris in Aegypto; et idcirco praecipio tibi, ut facias hanc rem.
DEUT|25|1|Si fuerit causa inter aliquos, et interpellaverint iudices, quem iustum esse perspexerint, illi iustitiae palmam dabunt; quem impium, condemnabunt impietatis.
DEUT|25|2|Sin autem iudex eum, qui peccavit, dignum viderit plagis, prosternet et coram se faciet verberari; pro mensura peccati erit et plagarum modus,
DEUT|25|3|ita dumtaxat, ut quadragenarium numerum non excedant, ne ultra percussus plagis multis et foede laceratus ante oculos tuos abeat frater tuus.
DEUT|25|4|Non ligabis os bovis terentis in area fruges tuas.
DEUT|25|5|Quando habitaverint fratres simul, et unus ex eis absque filio mortuus fuerit, uxor defuncti non nubet foras alteri, sed accipiet eam frater eius uxorem et suscitabit semen fratris sui;
DEUT|25|6|et primogenitum ex ea filium nomine illius appellabit, ut non deleatur nomen eius ex Israel.
DEUT|25|7|Sin autem noluerit accipere uxorem fratris sui, quae ei lege debetur, perget mulier ad portam civitatis et interpellabit maiores natu dicetque: Non vult frater viri mei suscitare nomen fratris sui in Israel nec me in coniugium sumere";
DEUT|25|8|statimque accersiri eum facient et interrogabunt. Si responderit: "Nolo eam uxorem accipere",
DEUT|25|9|accedet mulier ad eum coram senioribus et tollet calceamentum de pede eius spuetque in faciem illius et dicet: "Sic fit homini, qui non aedificat domum fratris sui".
DEUT|25|10|Et vocabitur nomen illius in Israel: "Domus discalceati".
DEUT|25|11|Si habuerint inter se iurgium viri, et unus contra alterum rixari coeperit, volensque uxor alterius eruere virum suum de manu fortioris, miserit manum et apprehenderit verenda eius,
DEUT|25|12|abscides manum illius nec flecteris super eam ulla misericordia.
DEUT|25|13|Non habebis in sacculo tuo diversa pondera maius et minus;
DEUT|25|14|nec erit in domo tua ephi maius et minus.
DEUT|25|15|Pondus habebis iustum et verum, et ephi iustum et verum erit tibi, ut multo vivas tempore super terram, quam Dominus Deus tuus dederit tibi.
DEUT|25|16|Abominatur enim Dominus tuus eum, qui facit haec, et aversatur omnem iniustitiam.
DEUT|25|17|Memento quae fecerit tibi Amalec in via, quando egrediebaris ex Aegypto;
DEUT|25|18|quomodo occurrerit tibi et omnes extremos agminis tui, qui lassi residebant, ceciderit, quando tu eras fame et labore confectus, et non timuerit Deum.
DEUT|25|19|Cum ergo Dominus Deus tuus dederit tibi requiem a cunctis per circuitum inimicis tuis in terra, quam tibi daturus est, delebis nomen Amalec sub caelo: cave, ne obliviscaris!
DEUT|26|1|Cumque intraveris terram, quam Dominus Deus tuus ti bi daturus est possidendam, et obtinueris eam atque habitaveris in illa,
DEUT|26|2|tolles primitias de cunctis frugibus agri, quas collegeris de terra tua, quam Dominus Deus tuus dabit tibi, et pones in cartallo pergesque ad locum, quem Dominus Deus tuus elegerit, ut ibi habitet nomen eius,
DEUT|26|3|accedesque ad sacerdotem, qui fuerit in diebus illis, et dices ad eum: Profiteor hodie coram Domino Deo tuo quod ingressus sim terram, pro qua iuravit patribus nostris, ut daret eam nobis".
DEUT|26|4|Suscipiensque sacerdos cartallum de manu tua ponet ante altare Domini Dei tui,
DEUT|26|5|et loqueris in conspectu Domini Dei tui: "Syrus vagus erat pater meus et descendit in Aegyptum et ibi peregrinatus est in paucissimo numero; crevitque in gentem magnam ac robustam et infinitae multitudinis.
DEUT|26|6|Afflixeruntque nos Aegyptii et persecuti sunt imponentes onera gravissima.
DEUT|26|7|Et clamavimus ad Dominum, Deum patrum nostrorum, qui exaudivit nos et respexit humilitatem nostram et laborem atque angustias,
DEUT|26|8|et eduxit nos Dominus de Aegypto in manu forti et brachio extento, in ingenti pavore, in signis atque portentis,
DEUT|26|9|et introduxit ad locum istum et tradidit nobis terram hanc lacte et melle manantem.
DEUT|26|10|Et ecce nunc attuli primitias frugum terrae, quam dedisti mihi, Domine". Et dimittes eas in conspectu Domini Dei tui et adorato Domino Deo tuo.
DEUT|26|11|Et epulaberis in omnibus bonis, quae Dominus Deus tuus dederit tibi et domui tuae, tu et Levites et advena, qui tecum est.
DEUT|26|12|Quando compleveris decimam cunctarum frugum tuarum, anno tertio, anno decimarum, et dederis Levitae et advenae et pupillo et viduae, ut comedant intra portas tuas et saturentur,
DEUT|26|13|loqueris in conspectu Domini Dei tui: "Abstuli, quod sanctificatum est, de domo mea et dedi illud Levitae et advenae, pupillo ac viduae, sicut iussisti mihi; non praeterivi mandata tua nec sum oblitus imperii tui,
DEUT|26|14|non comedi ex eis in luctu meo nec separavi ex eis in qualibet immunditia nec expendi ex his quidquam mortuo: oboedivi voci Domini Dei mei et feci omnia, sicut praecepisti mihi.
DEUT|26|15|Respice de habitaculo sancto tuo, de caelo, et benedic populo tuo Israel et terrae, quam dedisti nobis, sicut iurasti patribus nostris, terrae lacte et melle mananti".
DEUT|26|16|Hodie Dominus Deus tuus mandavit tibi, ut facias praecepta haec atque iudicia et custodias et impleas illa ex toto corde tuo et ex tota anima tua.
DEUT|26|17|Dominum elegisti hodie, ut sit tibi Deus, et ambules in viis eius et custodias praecepta illius et mandata atque iudicia et oboedias eius imperio;
DEUT|26|18|et Dominus elegit te hodie, ut sis ei populus peculiaris, sicut locutus est tibi, et custodias omnia mandata illius,
DEUT|26|19|et faciat te excelsiorem cunctis gentibus, quas creavit in laudem et nomen et gloriam suam, ut sis populus sanctus Domini Dei tui, sicut locutus est ".
DEUT|27|1|Praecepit autem Moyses et seniores Israel populo dicen tes: " Custodite omne mandatum, quod praecipio vobis hodie.
DEUT|27|2|Cumque transieritis Iordanem in terram, quam Dominus Deus tuus dabit tibi, eriges ingentes lapides et calce obduces eos,
DEUT|27|3|ut possis in eis scribere omnia verba legis huius, Iordane transmisso, ut introeas terram, quam Dominus Deus tuus dabit tibi, terram lacte et melle manantem, sicut locutus est Dominus, Deus patrum tuorum, tibi.
DEUT|27|4|Quando ergo transieritis Iordanem, erigite istos lapides, sicut ego hodie praecipio vobis, in monte Hebal, et obduces eos calce;
DEUT|27|5|et aedificabis ibi altare Domino Deo tuo de lapidibus, quos ferrum non tetigit,
DEUT|27|6|de saxis impolitis, et offeres super eo holocausta Domino Deo tuo.
DEUT|27|7|Et immolabis hostias pacificas comedesque ibi et epulaberis coram Domino Deo tuo;
DEUT|27|8|et scribes super lapides omnia verba legis huius plane et lucide ".
DEUT|27|9|Dixeruntque Moyses et sacerdotes levitici generis ad omnem Israelem: " Attende et audi, Israel: hodie factus es populus Domino Deo tuo;
DEUT|27|10|audies vocem eius et facies mandata atque praecepta, quae ego praecipio tibi ".
DEUT|27|11|Praecepitque Moyses populo in die illo dicens:
DEUT|27|12|" Hi stabunt ad benedicendum populo super montem Garizim, Iordane transmisso: Simeon, Levi, Iudas, Issachar, Ioseph et Beniamin.
DEUT|27|13|Et e regione isti stabunt ad maledicendum in monte Hebal: Ruben, Gad et Aser et Zabulon, Dan et Nephthali.
DEUT|27|14|Et pronunciabunt Levitae dicentque ad omnes viros Israel excelsa voce:
DEUT|27|15|"Maledictus homo, qui facit sculptile et conflatile, abominationem Domini, opus manuum artificum, ponetque illud in abscondito". Et respondebit omnis populus et dicet: "Amen".
DEUT|27|16|"Maledictus, qui contemnit patrem suum et matrem". Et dicet omnis populus: "Amen".
DEUT|27|17|"Maledictus, qui transfert terminos proximi sui". Et dicet omnis populus: "Amen".
DEUT|27|18|"Maledictus, qui errare facit caecum in itinere". Et dicet omnis populus: "Amen".
DEUT|27|19|"Maledictus, qui pervertit iudicium advenae, pupilli et viduae". Et dicet omnis populus: "Amen".
DEUT|27|20|"Maledictus, qui dormit cum uxore patris sui, quia revelat operimentum lectuli eius". Et dicet omnis populus: "Amen".
DEUT|27|21|"Maledictus, qui dormit cum omni iumento". Et dicet omnis populus: Amen".
DEUT|27|22|"Maledictus, qui dormit cum sorore sua, filia patris sui sive matris suae". Et dicet omnis populus: "Amen".
DEUT|27|23|"Maledictus, qui dormit cum socru sua". Et dicet omnis populus: "Amen".
DEUT|27|24|"Maledictus, qui clam percusserit proximum suum". Et dicet omnis populus: "Amen".
DEUT|27|25|"Maledictus, qui accipit munera, ut percutiat sanguinem innocentem". Et dicet omnis populus: "Amen".
DEUT|27|26|"Maledictus, qui non permanet in sermonibus legis huius nec eos opere perficit". Et dicet omnis populus: "Amen".
DEUT|28|1|Sin audieris vocem Domini Dei tui, ut facias atque custo dias omnia mandata eius, quae ego praecipio tibi hodie, faciet te Dominus Deus tuus excelsiorem cunctis gentibus, quae versantur in terra,
DEUT|28|2|venientque super te universae benedictiones istae et apprehendent te, si tamen vocem Domini Dei tui audieris.
DEUT|28|3|Benedictus tu in civitate et benedictus in agro.
DEUT|28|4|Benedictus fructus ventris tui et fructus terrae tuae fructusque iumentorum tuorum, partus armentorum tuorum et incrementum ovium tuarum.
DEUT|28|5|Benedictum canistrum et pistrinum tuum.
DEUT|28|6|Benedictus eris et ingrediens et egrediens.
DEUT|28|7|Dabit Dominus inimicos tuos, qui consurgunt adversum te, corruentes in conspectu tuo; per unam viam venient contra te et per septem fugient a facie tua.
DEUT|28|8|Emittet Dominus benedictionem super cellaria tua et super omnia opera manuum tuarum; benedicetque tibi in terra, quam Dominus Deus tuus dabit tibi.
DEUT|28|9|Suscitabit te Dominus sibi in populum sanctum, sicut iuravit tibi, si custodieris mandata Domini Dei tui et ambulaveris in viis eius.
DEUT|28|10|Videbuntque omnes terrarum populi quod nomen Domini invocatum sit super te, et timebunt te.
DEUT|28|11|Abundare te faciet Dominus omnibus bonis, fructu uteri tui et fructu iumentorum tuorum, fructu terrae tuae, quam iuravit Dominus patribus tuis, ut daret tibi.
DEUT|28|12|Aperiet Dominus tibi thesaurum suum optimum, caelum, ut tribuat pluviam terrae tuae in tempore suo; benedicatque cunctis operibus manuum tuarum; et fenerabis gentibus multis et ipse a nullo fenus accipies.
DEUT|28|13|Constituet te Dominus in caput et non in caudam, et eris semper supra et non subter, si audieris mandata Domini Dei tui, quae ego praecipio tibi hodie, et custodieris et feceris
DEUT|28|14|ac non declinaveris a verbis, quae ego praecipio vobis hodie, nec ad dexteram nec ad sinistram, nec secutus fueris deos alienos neque colueris eos.
DEUT|28|15|Quod si audire nolueris vocem Domini Dei tui, ut custodias et facias omnia mandata eius et praecepta, quae ego praecipio tibi hodie, venient super te omnes maledictiones istae et apprehendent te:
DEUT|28|16|Maledictus eris in civitate, maledictus in agro.
DEUT|28|17|Maledictum canistrum et pistrinum tuum.
DEUT|28|18|Maledictus fructus ventris tui et fructus terrae tuae, partus armentorum tuorum et incrementum ovium tuarum.
DEUT|28|19|Maledictus eris ingrediens et maledictus egrediens.
DEUT|28|20|Mittet Dominus super te maledictionem et conturbationem et increpationem in omnia opera tua, quae facies, donec conterat te et perdat velociter propter adinventiones tuas pessimas, in quibus reliquisti me.
DEUT|28|21|Adiunget Dominus tibi pestilentiam, donec consumat te de terra, ad quam ingredieris possidendam.
DEUT|28|22|Percutiet te Dominus consumptione, febri et inflammatione, ardore et aestu, uredine ac aurugine, et persequentur te, donec pereas.
DEUT|28|23|Et erit caelum, quod est supra caput tuum, aeneum, et terra, quam calcas, ferrea.
DEUT|28|24|Convertet Dominus imbrem terrae tuae in pulverem, et de caelo descendet super te cinis, donec conteraris.
DEUT|28|25|Tradet te Dominus corruentem ante hostes tuos: per unam viam egredieris contra eos et per septem fugies et eris in terrorem omnibus regnis terrae.
DEUT|28|26|Eritque cadaver tuum in escam cunctis volatilibus caeli et bestiis terrae, et non erit qui abigat.
DEUT|28|27|Percutiet te Dominus ulcere Aegypti et tumore, scabie quoque et prurigine, ita ut curari nequeas.
DEUT|28|28|Percutiet te Dominus amentia et caecitate ac stupore mentis;
DEUT|28|29|et palpabis in meridie, sicut palpare solet caecus in tenebris, et non diriges vias tuas. Omnique tempore eris oppressus et exspoliatus nec habebis, qui liberet te.
DEUT|28|30|Uxorem accipies, et alius dormiet cum ea. Domum aedificabis et non habitabis in ea. Plantabis vineam et non vindemiabis eam.
DEUT|28|31|Bos tuus mactabitur coram te, et non comedes ex eo. Asinus tuus rapietur in conspectu tuo et non reddetur tibi. Oves tuae dabuntur inimicis tuis, et non erit qui te adiuvet.
DEUT|28|32|Filii tui et filiae tuae tradentur alteri populo, videntibus oculis tuis et deficientibus ad conspectum eorum tota die, et non erit fortitudo in manu tua.
DEUT|28|33|Fructus terrae tuae et omnes labores tuos comedet populus, quem ignoras, et eris semper oppressus et confractus cunctis diebus
DEUT|28|34|et insanies in aspectu eorum, quae videbunt oculi tui.
DEUT|28|35|Percutiet te Dominus ulcere pessimo in genibus et in suris, sanarique non poteris a planta pedis usque ad verticem tuum.
DEUT|28|36|Ducet te Dominus et regem tuum, quem constitueris super te, in gentem, quam ignorasti tu et patres tui, et servies ibi diis alienis, ligno et lapidi;
DEUT|28|37|et eris in stuporem et in proverbium ac fabulam omnibus populis, ad quos te introduxerit Dominus.
DEUT|28|38|Sementem multam iacies in terram et modicum congregabis, quia locustae devorabunt omnia.
DEUT|28|39|Vineas plantabis et coles et vinum non bibes nec colliges ex ea quippiam, quoniam vastabitur vermibus.
DEUT|28|40|Olivas habebis in omnibus terminis tuis et non ungeris oleo, quia defluent et peribunt.
DEUT|28|41|Filios generabis et filias et non frueris eis, quoniam ducentur in captivitatem.
DEUT|28|42|Omnes arbores tuas et fruges terrae tuae locusta consumet.
DEUT|28|43|Advena, qui tecum versatur in terra, ascendet super te eritque sublimior; tu autem descendes et eris inferior.
DEUT|28|44|Ipse fenerabit tibi, et tu non fenerabis ei; ipse erit in caput, et tu eris in caudam.
DEUT|28|45|Et venient super te omnes maledictiones istae et persequentes apprehendent te, donec intereas, quia non audisti vocem Domini Dei tui nec servasti mandata eius et praecepta, quae praecepit tibi.
DEUT|28|46|Et erunt in te signa atque prodigia et in semine tuo usque in sempiternum.
DEUT|28|47|Eo quod non servieris Domino Deo tuo in gaudio cordisque laetitia propter rerum omnium abundantiam,
DEUT|28|48|servies inimico tuo, quem immittet Dominus tibi, in fame et siti et nuditate et omnium penuria, et ponet iugum ferreum super cervicem tuam, donec te conterat.
DEUT|28|49|Adducet Dominus super te gentem de longinquo et de extremis finibus terrae in similitudinem aquilae volantis cum impetu, cuius linguam intellegere non possis:
DEUT|28|50|gentem procacissimam, quae non deferat seni nec misereatur parvulo;
DEUT|28|51|et devoret fructum iumentorum tuorum ac fruges terrae tuae, donec intereas, et non relinquat tibi triticum, vinum et oleum, partum armentorum et incrementum ovium, donec te disperdat
DEUT|28|52|et obsideat te in cunctis urbibus tuis, donec destruantur muri tui firmi atque sublimes, in quibus habebas fiduciam in omni terra tua. Obsideberis intra portas tuas in omni terra tua, quam dabit tibi Dominus Deus tuus,
DEUT|28|53|et comedes fructum uteri tui, carnes filiorum tuorum et filiarum tuarum, quas dederit tibi Dominus Deus tuus, in obsidione et angustia, qua opprimet te hostis tuus.
DEUT|28|54|Homo tener in te et delicatus valde invidebit fratri suo et uxori, quae cubat in sinu suo, et residuis filiis suis, quos reservaverit,
DEUT|28|55|ne det uni ex eis de carnibus filiorum suorum, quas comedet, eo quod nihil aliud habeat in obsidione et angustia, qua oppresserit te inimicus tuus intra omnes portas tuas.
DEUT|28|56|Tenera mulier in te et delicata, quae non tentabat pedis vestigium figere in terram propter mollitiem et teneritudinem nimiam, invidebit viro suo, qui cubat in sinu eius, filio et filiae
DEUT|28|57|et illuviei secundarum, quae egrediuntur de medio feminum eius, et liberis, qui eadem hora nati sunt; comedet enim eos clam propter rerum omnium penuriam in obsidione et angustia, qua opprimet te inimicus tuus intra portas tuas.
DEUT|28|58|Nisi custodieris et feceris omnia verba legis huius, quae scripta sunt in hoc volumine, et timueris nomen gloriosum et terribile hoc, Dominum Deum tuum,
DEUT|28|59|augebit ultra modum Dominus plagas tuas et plagas seminis tui, plagas magnas et perseverantes, infirmitates pessimas et perpetuas,
DEUT|28|60|et convertet in te omnes afflictiones Aegypti, quas timuisti, et adhaerebunt tibi.
DEUT|28|61|Insuper universos languores et plagas, quae non sunt scriptae in volumine legis huius, inducet Dominus super te, donec te conterat;
DEUT|28|62|et remanebitis pauci numero, qui prius eratis sicut astra caeli prae multitudine, quoniam non audisti vocem Domini Dei tui.
DEUT|28|63|Et sicut ante laetatus est Dominus super vos bene vobis faciens vosque multiplicans, sic laetabitur super vos disperdens vos atque subvertens, ut auferamini de terra, ad quam ingredieris possidendam.
DEUT|28|64|Disperget te Dominus in omnes populos a summitate terrae usque ad terminos eius, et servies ibi diis alienis, quos et tu ignorasti et patres tui, lignis et lapidibus.
DEUT|28|65|In gentibus quoque illis non quiesces, neque erit requies vestigio pedis tui; dabit enim tibi Dominus ibi cor pavidum et deficientes oculos et animam consumptam maerore.
DEUT|28|66|Et erit vita tua quasi pendens ante te; timebis nocte et die et non credes vitae tuae.
DEUT|28|67|Mane dices: "Quis mihi det vesperum?"; et vespere: "Quis mihi det mane?", propter cordis tui formidinem, qua terreberis, et propter ea, quae tuis videbis oculis.
DEUT|28|68|Reducet te Dominus classibus in Aegyptum per viam, de qua dixi tibi, ut eam amplius non videres; ibi vendetis vos inimicis vestris in servos et ancillas, et non erit qui emat ".
DEUT|28|69|Haec sunt verba foederis, quod praecepit Dominus Moysi, ut feriret cum filiis Israel in terra Moab, praeter illud foedus, quod cum eis pepigit in Horeb.
DEUT|29|1|Vocavitque Moyses omnem Israel et dixit ad eos: " Vos vidistis universa, quae fecit Dominus coram vobis in terra Aegypti pharaoni et omnibus servis eius universaeque terrae illius,
DEUT|29|2|tentationes magnas, quas viderunt oculi tui, signa illa portentaque ingentia;
DEUT|29|3|et non dedit Dominus vobis cor intellegens et oculos videntes et aures, quae possint audire, usque in praesentem diem.
DEUT|29|4|Adduxi vos quadraginta annis per desertum; non sunt attrita vestimenta vestra, nec calceamenta pedum tuorum vetustate consumpta sunt,
DEUT|29|5|panem non comedistis, vinum et siceram non bibistis, ut sciretis quia ego sum Dominus Deus vester.
DEUT|29|6|Et venistis ad hunc locum, egressusque est Sehon rex Hesebon et Og rex Basan occurrentes nobis ad pugnam, et percussimus eos.
DEUT|29|7|Et tulimus terram eorum ac tradidimus possidendam Ruben et Gad et dimidiae tribui Manasse.
DEUT|29|8|Custodite ergo verba pacti huius et implete ea, ut prosperemini in universis, quae facitis.
DEUT|29|9|Vos statis hodie cuncti coram Domino Deo vestro, principes vestri ac tribus et maiores natu atque praefecti, omnis vir Israel,
DEUT|29|10|liberi et uxores vestrae et advena tuus, qui tecum moratur in castris, a lignorum caesoribus usque ad hos, qui hauriunt aquas tuas,
DEUT|29|11|ut transeas in foedere Domini Dei tui et in iure iurando, quod hodie Dominus Deus tuus percutit tecum,
DEUT|29|12|ut suscitet te sibi hodie in populum, et ipse sit Deus tuus, sicut locutus est tibi et sicut iuravit patribus tuis, Abraham, Isaac et Iacob.
DEUT|29|13|Nec vobis solis ego hoc foedus ferio et haec iuramenta confirmo,
DEUT|29|14|sed cunctis hic nobiscum hodie praesentibus coram Domino Deo nostro et illis, qui hodie hic nobiscum non adsunt.
DEUT|29|15|Vos enim nostis quomodo habitaverimus in terra Aegypti et quomodo transierimus per medium nationum, quas transeuntes
DEUT|29|16|vidistis abominationes et idola eorum, lignum et lapidem, argentum et aurum, quae colebant.
DEUT|29|17|Ne forte sit inter vos vir aut mulier, familia aut tribus, cuius cor aversum est hodie a Domino Deo nostro, ut vadat et serviat diis illarum gentium, et sit inter vos radix germinans fel et absinthium;
DEUT|29|18|cumque audierit verba iuramenti huius, benedicat sibi in corde suo dicens: "Pax erit mihi, etsi ambulabo in pravitate cordis mei", et absumat terram irriguam et sitientem.
DEUT|29|19|Dominus non ignoscet ei, sed tunc quam maxime furor eius fumabit et zelus contra hominem illum, et sedebunt super eum omnia maledicta, quae scripta sunt in hoc volumine, et delebit Dominus nomen eius sub caelo
DEUT|29|20|et consumet eum in perditionem ex omnibus tribubus Israel, iuxta maledictiones foederis, quae in hoc libro legis scriptae sunt.
DEUT|29|21|Dicetque sequens generatio, filii vestri, qui nascentur deinceps, et peregrini, qui de longe venerint, videntes plagas terrae illius et infirmitates, quibus eam afflixerit Dominus,
DEUT|29|22|sulphur et salem: combusta est omnis humus eius, ita ut ultra non seratur, nec virens quippiam germinet in exemplum subversionis Sodomae et Gomorrae, Adamae et Seboim, quas subvertit Dominus in ira et furore suo.
DEUT|29|23|Et dicent omnes gentes: "Quare sic fecit Dominus terrae huic? Quae est haec ira furoris immensa?".
DEUT|29|24|Et respondebunt: "Quia dereliquerunt pactum Domini, Dei patrum suorum, quod pepigit cum eis, quando eduxit eos de terra Aegypti,
DEUT|29|25|et servierunt diis alienis et adoraverunt eos, quos nesciebant et quibus non fuerant attributi;
DEUT|29|26|idcirco iratus est furor Domini contra terram istam, ut induceret super eam omnia maledicta, quae in hoc volumine scripta sunt,
DEUT|29|27|et eiecit eos de terra eorum in ira et furore et indignatione maxima proiecitque in terram alienam, sicut hodie comprobatur".
DEUT|29|28|Abscondita Domino Deo nostro, manifesta autem nobis et filiis nostris usque in sempiternum, ut faciamus universa verba legis huius.
DEUT|30|1|Cum ergo venerint super te omnes sermones isti, benedic tio et maledictio, quas proposui in conspectu tuo, et ductus paenitudine cordis tui in universis gentibus, in quas disperserit te Dominus Deus tuus,
DEUT|30|2|et reversus fueris ad eum et oboedieris eius imperiis secundum omnia, quae ego hodie praecipio tibi, cum filiis tuis in toto corde tuo et in tota anima tua,
DEUT|30|3|reducet Dominus Deus tuus captivitatem tuam ac miserebitur tui et rursum congregabit te de cunctis populis, in quos te ante dispersit.
DEUT|30|4|Si ad cardines caeli fueris dissipatus, inde te retrahet Dominus Deus tuus et assumet
DEUT|30|5|atque introducet in terram, quam possederunt patres tui, et obtinebis eam; et feliciorem et maioris numeri esse te faciet quam fuerunt patres tui.
DEUT|30|6|Circumcidet Dominus Deus tuus cor tuum et cor seminis tui, ut diligas Dominum Deum tuum in toto corde tuo et in tota anima tua, ut possis vivere.
DEUT|30|7|Omnes autem maledictiones has convertet super inimicos tuos et eos, qui oderunt te et persequuntur.
DEUT|30|8|Tu autem reverteris et audies vocem Domini faciesque universa mandata, quae ego praecipio tibi hodie;
DEUT|30|9|et abundare te faciet Dominus Deus tuus in cunctis operibus manuum tuarum, in subole uteri tui et in fructu iumentorum tuorum et in ubertate terrae tuae, in rerum omnium largitate; revertetur enim Dominus, ut gaudeat super te in omnibus bonis, sicut gavisus est in patribus tuis.
DEUT|30|10|Si tamen audieris vocem Domini Dei tui et custodieris mandata eius et praecepta, quae in hac lege conscripta sunt, et revertaris ad Dominum Deum tuum in toto corde tuo et in tota anima tua.
DEUT|30|11|Mandatum hoc, quod ego praecipio tibi hodie, non supra te est neque procul positum
DEUT|30|12|nec in caelo situm, ut possis dicere: "Quis nobis ad caelum valet ascendere, ut deferat illud ad nos, et audiamus atque opere compleamus?".
DEUT|30|13|Neque trans mare positum, ut causeris et dicas: "Quis nobis transfretare poterit mare et illud ad nos usque deferre, ut possimus audire et facere quod praeceptum est?".
DEUT|30|14|Sed iuxta te est sermo valde in ore tuo et in corde tuo, ut facias illum.
DEUT|30|15|Considera quod hodie proposuerim in conspectu tuo vitam et bonum, et e contrario mortem et malum.
DEUT|30|16|Si oboedieris mandatis Domini Dei tui, quae ego praecipio tibi hodie, ut diligas Dominum Deum tuum et ambules in viis eius et custodias mandata illius et praecepta atque iudicia, vives; ac multiplicabit te benedicetque tibi in terra, ad quam ingredieris possidendam.
DEUT|30|17|Sin autem aversum fuerit cor tuum, et audire nolueris atque errore deceptus adoraveris deos alienos et servieris eis,
DEUT|30|18|praedico vobis hodie quod pereatis et parvo tempore moremini in terra, ad quam, Iordane transmisso, ingredieris possidendam.
DEUT|30|19|Testes invoco hodie contra vos caelum et terram quod proposuerim vobis vitam et mortem, benedictionem et maledictionem. Elige ergo vitam, ut et tu vivas et semen tuum
DEUT|30|20|et diligas Dominum Deum tuum atque oboedias voci eius et illi adhaereas ipse est enim vita tua et longitudo dierum tuorum - ut habites in terra, pro qua iuravit Dominus patribus tuis, Abraham, Isaac et Iacob, ut daret eam illis ".
DEUT|31|1|Abiit itaque Moyses et locu tus est omnia verba haec ad universum Israel
DEUT|31|2|et dixit ad eos: " Centum viginti annorum sum hodie, non possum ultra egredi et ingredi, praesertim cum et Dominus dixerit mihi: "Non transibis Iordanem istum".
DEUT|31|3|Dominus Deus tuus ipse transibit ante te; ipse delebit gentes has in conspectu tuo, et possidebis eas, et Iosue transibit ante te, sicut locutus est Dominus.
DEUT|31|4|Facietque Dominus eis, sicut fecit Sehon et Og regibus Amorraeorum et terrae eorum delevitque eos.
DEUT|31|5|Cum ergo et hos tradiderit vobis, similiter facietis eis, sicut praecepi vobis.
DEUT|31|6|Viriliter agite et confortamini; nolite timere nec paveatis a conspectu eorum, quia Dominus Deus tuus ipse est ductor tuus et non dimittet nec derelinquet te ".
DEUT|31|7|Vocavitque Moyses Iosue et dixit ei coram omni Israel: " Confortare et esto robustus; tu enim introduces populum istum in terram, quam daturum se patribus eorum iuravit Dominus, et tu eam sorte divides eis.
DEUT|31|8|Et Dominus, qui ductor tuus est, ipse erit tecum, non dimittet nec derelinquet te; noli timere nec paveas ".
DEUT|31|9|Et scripsit Moyses legem hanc et tradidit eam sacerdotibus filiis Levi, qui portabant arcam foederis Domini, et cunctis senioribus Israel;
DEUT|31|10|praecepitque eis dicens: " Post septem annos, anno remissionis, in sollemnitate Tabernaculorum,
DEUT|31|11|convenientibus cunctis ex Israel, ut appareant in conspectu Domini Dei tui in loco, quem elegerit, leges verba legis huius coram omni Israel, audientibus eis;
DEUT|31|12|congrega populum tam viros quam mulieres, parvulos et advenas, qui sunt intra portas tuas, ut audientes discant et timeant Dominum Deum vestrum et custodiant impleantque omnes sermones legis huius;
DEUT|31|13|filii quoque eorum, qui nunc ignorant, audiant et discant timere Dominum Deum vestrum cunctis diebus, quibus versamini in terra, ad quam vos, Iordane transmisso, pergitis obtinendam ".
DEUT|31|14|Et ait Dominus ad Moysen: " Ecce prope sunt dies mortis tuae; voca Iosue, et state in tabernaculo conventus, ut praecipiam ei ". Abierunt ergo Moyses et Iosue et steterunt in tabernaculo conventus;
DEUT|31|15|apparuitque Dominus ibi in columna nubis, quae stetit in introitu tabernaculi.
DEUT|31|16|Dixitque Dominus ad Moysen: " Ecce tu dormies cum patribus tuis, et populus iste consurgens fornicabitur post deos alienos terrae, ad quam ingredietur; ibi derelinquet me et irritum faciet foedus, quod pepigi cum eo.
DEUT|31|17|Et irascetur furor meus contra eum in die illo, et derelinquam eos et abscondam faciem meam ab eis, et erit in devorationem; invenient eum mala multa et afflictiones, ita ut dicat in illo die: "Vere, quia non est Deus mecum, invenerunt me haec mala".
DEUT|31|18|Ego autem abscondam et celabo faciem meam in die illo, propter omnia mala, quae fecit, quia secutus est deos alienos.
DEUT|31|19|Nunc itaque scribite vobis canticum istud, et doce filios Israel, ut memoriter teneant et ore decantent, ut sit mihi carmen istud pro testimonio inter filios Israel.
DEUT|31|20|Introducam enim eum in terram, pro qua iuravi patribus eius, lacte et melle manantem. Cumque comederit et saturatus crassusque fuerit, avertetur ad deos alienos, et servient eis detrahentque mihi et irritum facient pactum meum.
DEUT|31|21|Postquam invenerint eum mala multa et afflictiones, respondebit ei canticum istud pro testimonio, quod nulla delebit oblivio ex ore seminis sui; scio enim cogitationes eius, quae facit hodie, antequam introducam eum in terram, quam ei pollicitus sum ".
DEUT|31|22|Scripsit ergo Moyses canticum istud in die illo et docuit filios Israel.
DEUT|31|23|Praecepitque Dominus Iosue filio Nun et ait: " Confortare et esto robustus; tu enim introduces filios Israel in terram, quam eis pollicitus sum, et ego ero tecum ".
DEUT|31|24|Postquam ergo scripsit Moyses verba legis huius in volumine atque complevit,
DEUT|31|25|praecepit Levitis, qui portabant arcam foederis Domini, dicens:
DEUT|31|26|" Tollite librum legis istum et ponite eum in latere arcae foederis Domini Dei vestri, ut sit ibi contra te in testimonium.
DEUT|31|27|Ego enim scio contentionem tuam et cervicem tuam durissimam. Adhuc vivente me vobiscum, semper contentiose egistis contra Dominum; quanto magis cum mortuus fuero?
DEUT|31|28|Congregate ad me omnes maiores natu per tribus vestras atque praefectos vestros, et loquar audientibus eis sermones istos et invocabo contra eos caelum et terram.
DEUT|31|29|Novi enim quod post mortem meam inique agetis et declinabitis de via, quam praecepi vobis, et occurrent vobis mala in extremo tempore, quando feceritis malum in conspectu Domini, ut irritetis eum per opera manuum vestrarum ".
DEUT|31|30|Locutus est ergo Moyses, audiente universo coetu Israel, verba carminis huius et ad finem usque complevit:
DEUT|32|1|" Audite, caeli, quae loquor; audiat terra verba oris mei!
DEUT|32|2|Stillet ut pluvia doctrina mea, fluat ut ros eloquium meumquasi imber super herbamet quasi stillae super gramina.
DEUT|32|3|Quia nomen Domini invocabo:date magnificentiam Deo nostro!
DEUT|32|4|Petra, perfecta sunt opera eius,quia omnes viae eius iustitia.Deus fidelis et absque ulla iniquitate,iustus et rectus.
DEUT|32|5|Peccaverunt ei non filii eius in sordibus suis,generatio prava atque perversa.
DEUT|32|6|Haeccine redditis Domino,popule stulte et insipiens?Numquid non ipse est pater tuus, qui possedit te,ipse fecit et stabilivit te?
DEUT|32|7|Memento dierum antiquorum,cogita generationes singulas;interroga patrem tuum, et annuntiabit tibi,maiores tuos, et dicent tibi.
DEUT|32|8|Quando dividebat Altissimus gentes,quando separabat filios Adam,constituit terminos populorumiuxta numerum filiorum Israel;
DEUT|32|9|pars autem Domini populus eius,Iacob funiculus hereditatis eius.
DEUT|32|10|Invenit eum in terra deserta,in loco horroris et ululatu solitudinis;circumdedit eum et attenditet custodivit quasi pupillam oculi sui.
DEUT|32|11|Sicut aquila provocans ad volandum pullos suoset super eos volitans expandit alas suaset assumpsit eumatque portavit super pennas suas.
DEUT|32|12|Dominus solus dux eius fuit,et non erat cum eo deus alienus.
DEUT|32|13|Constituit eum super excelsam terram,ut comederet fructus agrorum,ut sugeret mel de petraoleumque de saxo durissimo,
DEUT|32|14|butyrum de armento et lac de ovibus,cum adipe agnorum et arietumfiliorum Basan et hircorum,cum medulla tritici,et sanguinem uvae biberet meracissimum.
DEUT|32|15|Incrassatus est dilectus et recalcitravit;incrassatus, impinguatus, dilatatus dereliquit Deum factorem suumet recessit a Petra salutari suo.
DEUT|32|16|Provocaverunt eum in diis alieniset in abominationibus ad iracundiam concitaverunt.
DEUT|32|17|Immolaverunt daemonibus et non Deo,diis, quos ignorabant;novi recentesque venerunt,quos non coluerunt patres vestri.
DEUT|32|18|Petram, quae te genuit, dereliquisti,et oblitus es Domini creatoris tui.
DEUT|32|19|Vidit Dominus et sprevit,quia provocaverunt eum filii sui et filiae.
DEUT|32|20|Et ait: "Abscondam faciem meam ab eiset considerabo novissima eorum;generatio enim perversa est,et infideles filii.
DEUT|32|21|Ipsi me provocaverunt in eo, qui non erat Deus,et irritaverunt in vanitatibus suis;et ego provocabo eos in eo, qui non est populus,et in gente stulta irritabo illos.
DEUT|32|22|Ignis succensus est in furore meoet ardebit usque ad inferni profundissima;devorabitque terram cum germine suoet montium fundamenta comburet.
DEUT|32|23|Congregabo super eos malaet sagittas meas complebo in eis.
DEUT|32|24|Consumentur fame et devorabuntur febriet peste amarissima;dentes bestiarum immittam in eos, cum veneno serpentium in pulvere.
DEUT|32|25|Foris vastabit eos gladius,et intus pavor:iuvenem simul ac virginem,lactantem cum homine sene.
DEUT|32|26|Dixi: Disperdam eos,cessare faciam ex hominibus memoriam eorum!,
DEUT|32|27|sed arrogantiam inimicorum timui,ne superbirent hostes eorumet dicerent: >Manus nostra excelsa, et non Dominus fecit haec omnia!'.
DEUT|32|28|Gens enim absque consilio estet sine prudentia.
DEUT|32|29|Utinam saperent et intellegerent haecac novissima sua providerent!
DEUT|32|30|Quomodo persequatur unus mille,et duo fugent decem milia?Nonne ideo, quia Petra eorum vendidit eos,et Dominus tradidit illos?".
DEUT|32|31|Non enim est petra eorum ut Petra nostra,et inimici nostri sunt iudices.
DEUT|32|32|Vere de vinea Sodomorum vinea eorumet de suburbanis Gomorrae;uva eorum uva felliset botri amarissimi;
DEUT|32|33|fel draconum vinum eorumet venenum aspidum insanabile.
DEUT|32|34|Nonne haec condita sunt apud meet signata in thesauris meis?
DEUT|32|35|Mea est ultio, et ego retribuam in tempore,in quo labetur pes eorum!Iuxta est dies perditionis,et adesse festinat sors eorum.
DEUT|32|36|Iudicabit Dominus populum suumet in servis suis miserebitur;videbit quod infirmata sit manus,et defecerint clausi ac liberati.
DEUT|32|37|Et dicet: "Ubi sunt dii eorum,petra, in qua habebant fiduciam,
DEUT|32|38|de quorum victimis comedebant adipeset bibebant vinum libaminum?Surgant et opitulentur vobiset in necessitate vos protegant!
DEUT|32|39|Videte nunc quod ego sim solus,et non sit Deus praeter me.Ego occidam et ego vivere faciam;percutiam et ego sanabo;et non est qui de manu mea possit eruere.
DEUT|32|40|Levabo ad caelum manum meamet dicam: Vivo ego in aeternum!
DEUT|32|41|Si acuero ut fulgur gladium meum,et arripuerit iudicium manus mea,reddam ultionem hostibus meiset his, qui oderunt me, retribuam.
DEUT|32|42|Inebriabo sagittas meas sanguine,et gladius meus devorabit carnes:de cruore occisorum et captivorum,de capite ducum inimici!".
DEUT|32|43|Laudate, gentes, populum eius,quia sanguinem servorum suorum ulcisceturet vindictam retribuet in hostes suoset propitius erit terrae populi sui ".
DEUT|32|44|Venit ergo Moyses et locutus est omnia verba cantici huius in auribus populi, ipse et Iosue filius Nun;
DEUT|32|45|complevitque omnes sermones istos loquens ad universum Israel.
DEUT|32|46|Et dixit ad eos: " Ponite corda vestra in omnia verba, quae ego testificor vobis hodie, ut mandetis ea filiis vestris custodire et facere et implere universa verba legis huius;
DEUT|32|47|quia verbum non incassum vobis, sed est vita vestra: et in verbo hoc longo perseverabitis tempore in terra, ad quam, Iordane transmisso, ingredimini possidendam ".
DEUT|32|48|Locutusque est Dominus ad Moysen in eadem die dicens:
DEUT|32|49|" Ascende in montem istum Abarim, in montem Nabo, qui est in terra Moab contra Iericho, et vide terram Chanaan, quam ego tradam filiis Israel obtinendam.
DEUT|32|50|Et morere in monte, quem conscendens iungeris populo tuo, sicut mortuus est Aaron frater tuus in monte Hor et appositus populo suo.
DEUT|32|51|Quia praevaricati estis contra me in medio filiorum Israel ad aquas Meribathcades deserti Sin, quia non sanctificastis me inter filios Israel.
DEUT|32|52|E contra videbis terram et non ingredieris in eam, quam ego dabo filiis Israel ".
DEUT|33|1|Haec est benedictio, qua be nedixit Moyses homo Dei fi liis Israel ante mortem suam.
DEUT|33|2|Et ait: Dominus de Sinai venitet de Seir ortus est eis;apparuit de monte Pharanet venit in Meribathcadesde meridie eius in Asedoth.
DEUT|33|3|Vere diligit populos;omnes sancti eius in manu illius sunt;et, qui appropinquant pedibus tuis,accipient de doctrina tua.
DEUT|33|4|Legem praecepit nobis Moyses,hereditatem multitudinis Iacob.
DEUT|33|5|Et factus est apud dilectum rex,congregatis principibus populicum tribubus Israel ".
DEUT|33|6|" Vivat Ruben et non moriaturet sit parvus in numero ".
DEUT|33|7|Haec est Iudae benedictio: Audi, Domine, vocem Iudaeet ad populum suum introduc eum.Manus eius pugnabunt pro eo,et adiutor illius contra adversarios eius eris ".
DEUT|33|8|De Levi quoque ait: Tummim et Urim tuiviro sancto tuo,quem probasti in Massaet cum quo litigasti ad aquas Meriba.
DEUT|33|9|Qui dixit de patre suo et matre sua:Nescio vos";et fratres suos ignoravitet filios suos nescivit.Quia custodierunt eloquium tuumet pactum tuum servaverunt.
DEUT|33|10|Docebunt iudicia tua Iacobet legem tuam Israel;ponent thymiama in naribus tuiset holocaustum super altare tuum.
DEUT|33|11|Benedic, Domine, fortitudini eiuset opera manuum illius suscipe.Percute lumbos inimicorum eius;et, qui oderunt eum, non consurgant ".
DEUT|33|12|De Beniamin ait: Amantissimus Dominihabitabit confidenter in eo;Altissimus proteget eum tota dieet inter umeros illius requiescet ".
DEUT|33|13|De Ioseph quoque ait: Benedicta a Domino terra eius:donis caeli, roreatque abysso subiacente,
DEUT|33|14|fructibus soliset donis mensium,
DEUT|33|15|primitiis antiquorum montiumet donis collium aeternorum,
DEUT|33|16|frugibus terrae et plenitudine eius.Benedictio illius, qui apparuit in rubo,veniat super caput Iosephet super verticem nazaraei inter fratres suos;
DEUT|33|17|quasi primogeniti tauri pulchritudo eius,cornua unicornis cornua illius,in ipsis ventilabit gentesusque ad terminos terrae.Hae sunt multitudines Ephraim,et hae milia Manasse ".
DEUT|33|18|De Zabulon ait: Laetare, Zabulon, in exitu tuo,et Issachar, in tabernaculis tuis!
DEUT|33|19|Populos ad montem vocabunt,ibi immolabunt victimas iustitiae.Qui inundationem maris, quasi lac, sugentet thesauros absconditos arenarum ".
DEUT|33|20|De Gad ait: Benedictus, qui dilatat Gad!Quasi leo requiescitdilaceratque brachium et verticem.
DEUT|33|21|Et vidit primitias sibi,quia ibi pars ducis erat reposita;qui fuit cum principibus populiet fecit iustitiam Dominiet iudicia sua cum Israel ".
DEUT|33|22|De Dan quoque ait: Dan catulus leonisprosiliet largiter de Basan ".
DEUT|33|23|De Nephthali dixit: Nephthali satiabatur beneplacitoet plenus erit benedictione Domini:mare et meridiem possidebit ".
DEUT|33|24|De Aser quoque ait: Benedictus prae filiis Aser!Sit placens fratribus suiset tingat in oleo pedem suum.
DEUT|33|25|Ferrum et aes serae tuae,sicut dies tui robur tuum ".
DEUT|33|26|" Non est ut Deus Iesurun,qui ascendit super caelos ad auxilium tuumet in magnificentia sua super nubes.
DEUT|33|27|Habitaculum Deus antiquus,et subter brachia sempiterna.Eiciet a facie tua inimicumdicetque: "Conterere!".
DEUT|33|28|Habitabit Israel confidenter,et fons Iacob solus;stillabunt in terra frumenti et vini,caelique rorem.
DEUT|33|29|Beatus tu, Israel! Quis similis tui,popule, qui salvaris in Domino?Ipse est scutum auxilii tuiet gladius gloriae tuae.Blandientur tibi inimici tui,et tu eorum altitudines calcabis ".
DEUT|34|1|Ascendit ergo Moyses de campestribus Moab super montem Nabo in verticem Phasga contra Iericho; ostenditque ei Dominus omnem terram Galaad usque Dan
DEUT|34|2|et universum Nephthali terramque Ephraim et Manasse et omnem terram Iudae usque ad mare occidentale
DEUT|34|3|et Nageb et latitudinem campi Iericho civitatis palmarum usque Segor.
DEUT|34|4|Dixitque Dominus ad eum: " Haec est terra, pro qua iuravi Abraham, Isaac et Iacob, dicens: Semini tuo dabo eam. Vidisti eam oculis tuis et non transibis ad illam ".
DEUT|34|5|Mortuusque est ibi Moyses servus Domini in terra Moab, iubente Domino.
DEUT|34|6|Et sepelivit eum in valle in terra Moab contra Bethphegor; et non cognovit homo sepulcrum eius usque in praesentem diem.
DEUT|34|7|Moyses centum et viginti annorum erat, quando mortuus est; non caligavit oculus eius, nec robur illius defecit.
DEUT|34|8|Fleveruntque eum filii Israel in campestribus Moab triginta diebus; et completi sunt dies planctus lugentium Moysen.
DEUT|34|9|Iosue vero filius Nun repletus est spiritu sapientiae, quia Moyses posuit super eum manus suas; et oboedierunt ei filii Israel feceruntque, sicut praecepit Dominus Moysi.
DEUT|34|10|Et non surrexit ultra propheta in Israel sicut Moyses, quem nosset Dominus facie ad faciem,
DEUT|34|11|in omnibus signis atque portentis, quae misit per eum, ut faceret in terra Aegypti pharaoni et omnibus servis eius universaeque terrae illius,
DEUT|34|12|et in cuncta manu robusta magnisque mirabilibus, quae fecit Moyses coram universo Israel.
JOSH|1|1|Et factum est, ut post mortem Moysi servi Domini loqueretur Dominus ad Iosue filium Nun ministrum Moysi et diceret ei:
JOSH|1|2|" Moyses servus meus mortuus est; nunc igitur surge et transi Iordanem istum, tu et omnis populus iste, in terram, quam ego dabo filiis Israel.
JOSH|1|3|Omnem locum, quem calcaverit vestigium pedis vestri, vobis tradidi, sicut locutus sum Moysi.
JOSH|1|4|A deserto et Libano isto usque ad fluvium magnum Euphraten, omnis terra Hetthaeorum usque ad mare Magnum contra solis occasum erit terminus vester.
JOSH|1|5|Nullus tibi poterit resistere cunctis diebus vitae tuae: sicut fui cum Moyse, ero et tecum; non dimittam nec derelinquam te.
JOSH|1|6|Confortare et esto robustus; tu enim sorte divides populo huic terram, pro qua iuravi patribus suis, ut traderem eam illis.
JOSH|1|7|Confortare tantum et esto robustus valde, ut custodias et facias iuxta omnem legem, quam praecepit tibi Moyses servus meus. Ne declines ab ea ad dexteram vel ad sinistram, ut prospereris in omnibus, ad quaecumque perrexeris.
JOSH|1|8|Non recedat hoc volumen legis de ore tuo, sed meditaberis in eo diebus ac noctibus, ut custodias et facias iuxta omnia, quae scripta sunt in eo: tunc optime diriges viam tuam et tunc prosperaberis.
JOSH|1|9|Nonne praecepi tibi: Confortare et esto robustus, noli metuere et noli timere, quoniam tecum est Dominus Deus tuus in omnibus, ad quaecumque perrexeris?".
JOSH|1|10|Praecepitque Iosue praefectis populi dicens: " Transite per medium castrorum et imperate populo ac dicite:
JOSH|1|11|Praeparate vobis cibaria, quoniam post diem tertium transibitis Iordanem hunc et intrabitis ad possidendam terram, quam Dominus Deus vester daturus est vobis ".
JOSH|1|12|Rubenitis quoque et Gaditis et dimidiae tribui Manasse ait:
JOSH|1|13|" Mementote sermonis, quem praecepit vobis Moyses famulus Domini dicens: "Dominus Deus vester dedit vobis requiem et terram hanc".
JOSH|1|14|Uxores vestrae et filii ac iumenta manebunt in terra, quam tradidit vobis Moyses trans Iordanem; vos autem transibitis armati ante fratres vestros, omnes viri fortes, et adiuvabitis eos,
JOSH|1|15|donec det requiem Dominus fratribus vestris, sicut et vobis dedit, et possideant ipsi quoque terram, quam Dominus Deus vester daturus est eis. Et sic revertemini in terram possessionis vestrae et habitabitis in ea, quam vobis dedit Moyses famulus Domini trans Iordanem contra solis ortum.
JOSH|1|16|Responderuntque ad Iosue atque dixerunt: " Omnia, quae praecepisti nobis, faciemus et, quocumque miseris, ibimus.
JOSH|1|17|Sicut oboedivimus in cunctis Moysi, ita oboediemus et tibi; tantum sit Dominus Deus tuus tecum, sicut fuit cum Moyse.
JOSH|1|18|Quicumque contradixerit ori tuo et non oboedierit cunctis sermonibus, quos praeceperis ei, moriatur; tu tantum confortare et viriliter age ".
JOSH|2|1|Misit ergo Iosue filius Nun de Settim duos viros exploratores in abscondito et dixit eis; "Ite et considerate terram urbemque Iericho ". Qui pergentes ingressi sunt domum mulieris meretricis nomine Rahab et quieverunt ibi.
JOSH|2|2|Nuntiatumque est regi Iericho et dictum: " Ecce viri ingressi sunt huc per noctem de filiis Israel, ut explorarent terram ".
JOSH|2|3|Misitque rex Iericho ad Rahab dicens: " Educ viros, qui venerunt ad te et ingressi sunt domum tuam; exploratores quippe sunt et omnem terram considerare venerunt ".
JOSH|2|4|Tollensque mulier viros abscondit et ait: " Fateor, venerunt ad me, sed nesciebam unde essent;
JOSH|2|5|cumque porta clauderetur in tenebris, et illi pariter exierunt, nescio quo abierunt. Persequimini cito et comprehendetis eos ".
JOSH|2|6|Ipsa autem fecit ascendere viros in solarium domus suae operuitque eos lini stipula, quae ibi erat.
JOSH|2|7|Hi autem, qui missi fuerant, secuti sunt eos per viam, quae ducit ad vadum Iordanis; illisque egressis, statim porta clausa est.
JOSH|2|8|Necdum obdormierant qui latebant, et ecce mulier ascendit ad eos et ait:
JOSH|2|9|" Novi quod tradiderit Dominus vobis terram, et irruit in nos terror vester, et elanguerunt omnes habitatores terrae coram vobis.
JOSH|2|10|Audivimus enim quod siccaverit Dominus aquas maris Rubri ad vestrum introitum, quando egressi estis ex Aegypto, et quae feceritis duobus Amorraeorum regibus, qui erant trans Iordanem, Sehon et Og, quos interfecistis.
JOSH|2|11|Et haec audientes pertimuimus, et elanguit cor nostrum, nec remansit in nobis spiritus ad introitum vestrum; Dominus enim Deus vester ipse est Deus in caelo sursum et in terra deorsum.
JOSH|2|12|Nunc ergo iurate mihi per Dominum, ut, quomodo ego feci vobiscum misericordiam, ita et vos faciatis cum domo patris mei detisque mihi signum verum,
JOSH|2|13|ut salvetis patrem meum et matrem, fratres ac sorores meas et omnia, quae eorum sunt, et eruatis animas nostras de morte ".
JOSH|2|14|Qui responderunt ei: " Anima nostra sit pro vobis in mortem, si tamen non prodideris; cumque tradiderit nobis Dominus terram, faciemus in te misericordiam et veritatem ".
JOSH|2|15|Demisit ergo eos per funem de fenestra; domus enim eius haerebat muro, et in muro habitabat.
JOSH|2|16|Dixitque ad eos: " Ad montana pergite, ne forte occurrant vobis persecutores, ibique latete diebus tribus, donec redeant; et postea ibitis per viam vestram.
JOSH|2|17|Qui dixerunt ad eam: " Innoxii erimus a iuramento hoc, quo adiurasti nos,
JOSH|2|18|si, ingredientibus nobis terram, signum fuerit funiculus iste coccineus, et ligaveris eum in fenestra, per quam nos demisisti, et patrem tuum ac matrem fratresque et omnem cognationem tuam congregaveris in domum tuam.
JOSH|2|19|Qui ostium domus tuae egressus fuerit, sanguis ipsius erit in caput eius, et nos erimus innoxii; cunctorum autem sanguis, qui tecum fuerint in domo, redundabit in caput nostrum, si eos aliquis tetigerit.
JOSH|2|20|Quod si prodideris hoc verbum, erimus mundi ab hoc iuramento, quo adiurasti nos ".
JOSH|2|21|Et illa respondit: " Sicut locuti estis, ita fiat ". Dimittensque eos, ut pergerent, appendit funiculum coccineum in fenestra.
JOSH|2|22|Illi vero ambulantes pervenerunt ad montana et manserunt ibi tres dies, donec reverterentur, qui fuerant persecuti; quaerentes enim per omnem viam non reppererunt eos.
JOSH|2|23|Duo viri reversi sunt et descenderunt de monte et, transmisso Iordane, venerunt ad Iosue filium Nun narraveruntque ei omnia, quae acciderant sibi,
JOSH|2|24|atque dixerunt: " Tradidit Dominus in manus nostras omnem terram, et timore prostrati sunt cuncti habitatores eius in conspectu nostro ".
JOSH|3|1|Igitur Iosue de nocte consur gens movit castra. Egredientes que de Settim venerunt ad Iordanem, ipse et omnes filii Israel; et morati sunt ibi, antequam transirent.
JOSH|3|2|Tribus diebus evolutis, transierunt praefecti per castrorum medium
JOSH|3|3|et praeceperunt populo: " Quando videritis arcam foederis Domini Dei vestri et sacerdotes stirpis leviticae portantes eam, vos quoque consurgite et sequimini eam
JOSH|3|4|- sitque inter vos et arcam spatium cubitorum duum fere milium, et cavete, ne appropinquetis ad eam - ut sciatis per quam viam ingrediamini, quia prius non ambulastis per eam ".
JOSH|3|5|Dixitque Iosue ad populum: " Sanctificamini; cras enim faciet Dominus inter vos mirabilia ".
JOSH|3|6|Et ait ad sacerdotes: " Tollite arcam foederis et praecedite populum ". Qui tulerunt et ambulaverunt ante eos.
JOSH|3|7|Dixitque Dominus ad Iosue: " Hodie incipiam exaltare te coram omni Israel, ut sciant quod, sicut cum Moyse fui, ita et tecum sim.
JOSH|3|8|Tu autem praecipe sacerdotibus, qui portant arcam foederis, et dic eis: Cum veneritis ad oram aquae Iordanis, state in Iordane".
JOSH|3|9|Dixitque Iosue ad filios Israel: " Accedite huc et audite verba Domini Dei vestri ".
JOSH|3|10|Et rursum: " In hoc, inquit, scietis quod Deus vivens in medio vestri est et disperdet in conspectu vestro Chananaeum et Hetthaeum, Hevaeum et Pherezaeum, Gergesaeum quoque et Amorraeum et Iebusaeum.
JOSH|3|11|Ecce arca foederis Domini omnis terrae antecedet vos per Iordanem.
JOSH|3|12|Parate duodecim viros de tribubus Israel, singulos per singulas tribus;
JOSH|3|13|et cum posuerint vestigia pedum suorum sacerdotes, qui portant arcam Domini Dei universae terrae, in aquis Iordanis, aquae, quae inferiores sunt, decurrent, quae autem desuper veniunt, in una mole consistent ".
JOSH|3|14|Igitur egressus est populus de tabernaculis suis, ut transiret Iordanem; et sacerdotes, qui portabant arcam foederis, pergebant ante eum.
JOSH|3|15|Veneruntque usque ad Iordanem et, pedibus eorum in ora aquae tinctis - Iordanis autem omnes ripas alvei sui toto tempore messis impleverat -
JOSH|3|16|steterunt aquae desuper descendentes in loco uno instar molis procul valde apud urbem, quae vocatur Adam, ex latere Sarthan; quae autem inferiores erant, in mare Arabae, quod est mare Salsissimum, descenderunt, usquequo omnino deficerent.
JOSH|3|17|Populus autem incedebat contra Iericho, et sacerdotes, qui portabant arcam foederis Domini, stabant super siccam humum in medio Iordanis firmiter, donec omnis Israel compleret per arentem alveum transitum Iordanis.
JOSH|4|1|Quibus transgressis, dixit Dominus ad Iosue:
JOSH|4|2|" Sumite vobis de populo duodecim viros singulos per singulas tribus
JOSH|4|3|et praecipite eis, ut tollant de medio Iordanis alveo, ubi firmiter steterunt sacerdotum pedes, duodecim lapides; quos portabitis vobiscum et ponetis in loco castrorum, ubi fixeritis hac nocte tentoria ".
JOSH|4|4|Vocavitque Iosue duodecim viros, quos elegerat de filiis Israel, singulos de tribubus singulis,
JOSH|4|5|et ait ad eos: " Ite ante arcam Domini Dei vestri ad Iordanis medium et portate singuli singulos lapides in umeris vestris, iuxta numerum tribuum filiorum Israel,
JOSH|4|6|ut sit hoc signum inter vos. Quando interrogaverint vos filii vestri cras dicentes: "Quid sibi volunt isti lapides?",
JOSH|4|7|respondebitis eis: Defecerunt aquae Iordanis ante arcam foederis Domini, cum transiret eum; idcirco positi sunt lapides isti in monumentum filiis Israel usque in aeternum ".
JOSH|4|8|Fecerunt ergo filii Israel, sicut eis praecepit Iosue, portantes de medio Iordanis alveo duodecim lapides, ut ei Dominus imperarat, iuxta numerum tribuum filiorum Israel, usque ad locum, in quo castrametati sunt; ibique posuerunt eos.
JOSH|4|9|Alios quoque duodecim lapides posuit Iosue in medio Iordanis alveo, ubi steterunt sacerdotes, qui portabant arcam foederis; et sunt ibi usque in praesentem diem.
JOSH|4|10|Sacerdotes autem, qui portabant arcam, stabant in Iordanis medio, donec omnia complerentur, quae Iosue ut loqueretur ad populum praeceperat Dominus secundum omnia, quae dixerat ei Moyses. Festinavitque populus et transiit.
JOSH|4|11|Cumque transissent omnes, transivit et arca Domini; sacerdotesque pergebant ante populum.
JOSH|4|12|Filii quoque Ruben et Gad et dimidia tribus Manasse armati praecedebant filios Israel, sicut eis praeceperat Moyses;
JOSH|4|13|quadraginta fere milia expeditorum ad pugnam incedebant coram Domino in campestria Iericho.
JOSH|4|14|In illo die magnificavit Dominus Iosue coram omni Israel, ut timerent eum, sicut timuerant Moysen, omnibus diebus vitae suae.
JOSH|4|15|Dixitque ad eum:
JOSH|4|16|" Praecipe sacerdotibus, qui portant arcam testimonii, ut ascendant de Iordane ".
JOSH|4|17|Qui praecepit eis dicens: " Ascendite de Iordane ".
JOSH|4|18|Cumque ascendissent portantes arcam foederis Domini et siccam humum calcare coepissent, reversae sunt aquae in alveum suum et fluebant sicut ante super omnes ripas suas.
JOSH|4|19|Populus autem ascendit de Iordane decimo die mensis primi, et castrametati sunt in Galgalis, in termino orientali Iericho.
JOSH|4|20|Duodecim quoque lapides, quos de Iordanis alveo sumpserant, posuit Iosue in Galgalis.
JOSH|4|21|Et dixit ad filios Israel: " Quando interrogaverint filii vestri cras patres suos et dixerint eis: "Quid sibi volunt isti lapides?",
JOSH|4|22|docebitis eos atque dicetis: Per arentem alveum transivit Israel Iordanem istum,
JOSH|4|23|siccante Domino Deo vestro aquas eius in conspectu vestro, donec transiretis,
JOSH|4|24|sicut fecerat prius in mari Rubro, quod siccavit coram nobis, donec transiremus,
JOSH|4|25|ut cognoscant omnes terrarum populi fortissimam Domini manum, et ut vos timeatis Dominum Deum vestrum omni tempore ".
JOSH|5|1|Postquam ergo audierunt om nes reges Amorraeorum, qui ha bitabant trans Iordanem ad occidentalem plagam, et cuncti reges Chanaan, qui propinqua possidebant Magno mari loca, quod siccasset Dominus fluenta Iordanis coram filiis Israel, donec transirent, dissolutum est cor eorum, et non remansit in eis spiritus coram filiis Israel.
JOSH|5|2|Eo tempore ait Dominus ad Iosue: " Fac tibi cultros lapideos et circumcide iterum secundo filios Israel ".
JOSH|5|3|Fecit, quod iusserat Dominus, et circumcidit filios Israel in colle Praeputiorum.
JOSH|5|4|Haec autem causa est secundae circumcisionis: omnis populus, qui egressus est ex Aegypto, generis masculini, universi bellatores viri mortui sunt in deserto in via;
JOSH|5|5|qui omnes circumcisi erant. Populus autem, qui natus est in deserto, incircumcisus fuit.
JOSH|5|6|Per quadraginta enim annos ambulabant filii Israel, donec consumerentur omnes homines bellatores, qui non audierant vocem Domini, et quibus iuraverat, ut non ostenderet eis terram, super qua iuraverat patribus eorum, ut daret illis terram lacte et melle manantem.
JOSH|5|7|Horum filii in locum successerunt patrum et circumcisi sunt a Iosue, quia, sicut nati fuerant, in praeputio erant, nec eos in via aliquis circumciderat.
JOSH|5|8|Postquam autem omnes circumcisi sunt, manserunt in eodem castrorum loco, donec sanarentur.
JOSH|5|9|Dixitque Dominus ad Iosue: " Hodie abstuli opprobrium Aegypti a vobis ". Vocatumque est nomen loci illius Galgala usque in praesentem diem.
JOSH|5|10|Manseruntque filii Israel in Galgalis et fecerunt Pascha quarta decima die mensis ad vesperum in campestribus Iericho;
JOSH|5|11|et comederunt de frugibus terrae a die altero, azymos panes et polentam hoc ipso die.
JOSH|5|12|Defecitque manna a die sequenti, postquam comederunt de frugibus terrae, nec usi sunt ultra cibo illo filii Israel, sed comederunt de frugibus terrae Chanaan in anno illo.
JOSH|5|13|Cum autem esset Iosue in agro urbis Iericho, levavit oculos et vidit virum stantem contra se et evaginatum tenentem gladium; perrexitque ad eum et ait: " Noster es an adversariorum? ".
JOSH|5|14|Qui respondit: " Nequaquam, sed sum princeps exercitus Domini et nunc veni ".
JOSH|5|15|Cecidit Iosue pronus in terram et adorans ait: " Quid Dominus meus loquitur ad servum suum? ".
JOSH|5|16|Et dixit princeps exercitus Domini ad Iosue: " Solve calceamentum de pedibus tuis; locus enim, in quo stas, sanctus est ". Fecitque Iosue, ut sibi fuerat imperatum.
JOSH|6|1|Iericho autem erat munita et clausa coram filiis Israel, et nul lus egredi audebat aut ingredi.
JOSH|6|2|Dixitque Dominus ad Iosue: " Ecce dedi in manu tua Iericho et regem eius omnesque fortes viros.
JOSH|6|3|Circuite urbem cuncti bellatores semel per diem: sic facietis sex diebus.
JOSH|6|4|Septem sacerdotes portabunt septem bucinas, cornua arietum, ante arcam foederis. Die autem septimo septies circuibitis civitatem, et sacerdotes clangent bucinis.
JOSH|6|5|Cumque insonuerit vox tubae longior et in auribus vestris increpuerit, conclamabit omnis populus vociferatione maxima, et muri funditus corruent civitatis; ingredienturque singuli per locum, contra quem steterint ".
JOSH|6|6|Vocavit ergo Iosue filius Nun sacerdotes et dixit ad eos: " Tollite arcam foederis, et septem alii sacerdotes tollant septem bucinas et incedant ante arcam Domini ".
JOSH|6|7|Ad populum quoque ait: " Vadite et circuite civitatem, et viri armati praecedant arcam Domini ".
JOSH|6|8|Cumque Iosue verba finisset, septem sacerdotes septem bucinis clangebant ante arcam foederis Domini,
JOSH|6|9|omnisque armatus exercitus praecedebat sacerdotes clangentes, reliquum vulgus arcam sequebatur, ac bucinis omnia concrepabant.
JOSH|6|10|Praeceperat autem Iosue populo dicens: " Non clamabitis, nec audietur vox vestra, neque ullus sermo ex ore vestro egredietur, donec veniat dies, in quo dicam vobis: Clamate et vociferamini ".
JOSH|6|11|Circuivit ergo arca Domini civitatem per diem, et reversi in castra pernoctaverunt ibi.
JOSH|6|12|Igitur, Iosue de nocte consurgente, tulerunt sacerdotes arcam Domini,
JOSH|6|13|et septem ex eis septem bucinas, cornua arietum, praecedebantque arcam Domini ambulantes atque clangentes, et armatus populus ibat ante eos; vulgus autem reliquum sequebatur arcam, bucinis personantibus.
JOSH|6|14|Circuieruntque civitatem secundo die semel et reversi sunt in castra; sic fecerunt sex diebus.
JOSH|6|15|Die autem septimo, diluculo consurgentes circuierunt urbem eodem modo septies; in illo die tantum circuierunt urbem septies.
JOSH|6|16|Cumque septimo circuitu clangerent bucinis sacerdotes, dixit Iosue ad populum: " Vociferamini! Tradidit enim vobis Dominus civitatem.
JOSH|6|17|Sitque civitas anathema, ipsa et omnia, quae in ea sunt, Domino; sola Rahab meretrix vivat cum universis, qui cum ea in domo sunt: abscondit enim nuntios, quos direximus.
JOSH|6|18|Vos autem cavete, ne de anathemate quippiam auferatis et sitis praevaricationis rei, et omnia castra Israel anathema sint atque turbentur.
JOSH|6|19|Quidquid auri et argenti fuerit et vasorum aeneorum ac ferri, Domino consecretur repositum in thesauris eius ".
JOSH|6|20|Igitur, omni vociferante populo et clangentibus tubis, postquam in aures multitudinis vox sonitusque increpuit, muri ilico corruerunt; et ascendit unusquisque per locum, qui contra se erat, ceperuntque civitatem.
JOSH|6|21|Et interfecerunt omnia, quae erant in ea, a viro usque ad mulierem, ab infante usque ad senem; boves quoque et oves et asinos in ore gladii percusserunt.
JOSH|6|22|Duobus autem viris, qui exploratores missi fuerant, dixit Iosue: " Ingredimini domum mulieris meretricis et producite eam et omnia, quae illius sunt, sicut illi iuramento firmastis ".
JOSH|6|23|Ingressique iuvenes eduxerunt Rahab et parentes eius, fratres quoque et cunctam supellectilem ac cognationem illius et extra castra Israel manere fecerunt.
JOSH|6|24|Urbem autem et omnia, quae erant in ea, succenderunt, absque argento et auro et vasis aeneis ac ferro, quae in aerarium domus Domini consecrarunt.
JOSH|6|25|Rahab vero meretricem et domum patris eius et omnia, quae habebat, fecit Iosue vivere; et habitavit in medio Israel usque in praesentem diem, eo quod absconderit nuntios, quos miserat Iosue, ut explorarent Iericho.In tempore illo imprecatus est Iosue dicens:
JOSH|6|26|"Maledictus vir coram Domino, qui suscitaverit et aedificaverit civitatem Iericho; in primogenito suo fundamenta illius faciet et in novissimo liberorum ponet portas eius ".
JOSH|6|27|Fuit ergo Dominus cum Iosue, et nomen eius in omni terra vulgatum est.
JOSH|7|1|Filii autem Israel praevaricati sunt mandatum et usurpaverunt de anathemate: nam Achan filius Charmi filii Zabdi filii Zarae de tribu Iudae tulit aliquid de anathemate. Iratusque est Dominus contra filios Israel.
JOSH|7|2|Cumque mitteret Iosue de Iericho viros contra Hai, quae est iuxta Bethaven ad orientalem plagam oppidi Bethel, dixit eis: " Ascendite et explorate terram ". Qui praecepta complentes exploraverunt Hai
JOSH|7|3|et reversi dixerunt ei: " Non ascendat omnis populus, sed duo vel tria milia virorum pergant et deleant civitatem. Noli vexare omnem populum contra hostes paucissimos ".
JOSH|7|4|Ascenderunt ergo tria fere milia pugnatorum, qui statim terga verterunt coram viris urbis Hai,
JOSH|7|5|qui percusserunt ex eis circiter triginta et sex homines persecutique sunt eos de porta usque ad Sabarim et percusserunt eos in descensu; pertimuitque cor populi et instar aquae liquefactum est.
JOSH|7|6|Iosue vero scidit vestimenta sua et cecidit pronus in terram coram arca Domini usque ad vesperum, tam ipse quam omnes senes Israel; miseruntque pulverem super capita sua.
JOSH|7|7|Et dixit Iosue: " Heu, Domine Deus, quid voluisti traducere populum istum Iordanem fluvium, ut traderes nos in manus Amorraei et perderes? Utinam mansissemus trans Iordanem!
JOSH|7|8|Quaeso, Domine, quid dicam videns Israelem hostibus suis terga vertentem?
JOSH|7|9|Audient Chananaei et omnes habitatores terrae ac pariter conglobati circumdabunt nos atque delebunt nomen nostrum de terra. Et quid facies magno nomini tuo? ".
JOSH|7|10|Dixitque Dominus ad Iosue: " Surge! Cur iaces pronus in terra?
JOSH|7|11|Peccavit Israel et praevaricatus est pactum meum, quod mandaveram eis; tuleruntque de anathemate et furati sunt atque mentiti et absconderunt inter vasa sua.
JOSH|7|12|Nec poterunt filii Israel stare ante hostes suos eosque fugient, quia facti sunt anathema; non ero ultra vobiscum, donec conteratis anathema de medio vestri.
JOSH|7|13|Surge! Sanctifica populum et dic eis: Sanctificamini in crastinum. Haec enim dicit Dominus, Deus Israel: Anathema in medio tui est, Israel! Non poteris stare coram hostibus tuis, donec auferatis anathema de medio vestri.
JOSH|7|14|Accedetisque mane singuli per tribus vestras; et quamcumque tribum Dominus designaverit, accedet per cognationes suas et cognatio per domos domusque per viros:
JOSH|7|15|et quicumque ille in hoc facinore fuerit deprehensus, comburetur igni cum omnibus, quae ipsius sunt, quoniam praevaricatus est pactum Domini et fecit nefas in Israel ".
JOSH|7|16|Surgens itaque Iosue mane applicuit Israel per tribus suas, et inventa est tribus Iudae.
JOSH|7|17|Quae cum iuxta familias suas esset oblata, inventa est familia Zarae; illam quoque per domos offerens repperit Zabdi.
JOSH|7|18|Cuius domum in singulos dividens viros invenit Achan filium Charmi filii Zabdi filii Zarae de tribu Iudae.
JOSH|7|19|Et ait Iosue ad Achan: " Fili mi, da gloriam Domino, Deo Israel, et confitere atque indica mihi quid feceris; ne abscondas ".
JOSH|7|20|Responditque Achan Iosue et dixit ei: " Vere ego peccavi Domino, Deo Israel, et sic et sic feci:
JOSH|7|21|Vidi enim inter spolia pallium de Sennaar valde bonum et ducentos siclos argenti regulamque auream quinquaginta siclorum; et concupiscens abstuli et abscondi in terra contra medium tabernaculi mei argentumque subter ".
JOSH|7|22|Misit ergo Iosue ministros, qui currentes ad tabernaculum illius reppererunt cuncta abscondita in eodem loco et argentum simul;
JOSH|7|23|auferentesque de tentorio tulerunt ea ad Iosue et ad omnes filios Israel proieceruntque ante Dominum.
JOSH|7|24|Tollens itaque Iosue Achan filium Zarae argentumque et pallium et auream regulam filiosque eius et filias, boves et asinos et oves ipsumque tabernaculum et cunctam supellectilem - et omnis Israel cum eo - duxerunt eos ad vallem Achor,
JOSH|7|25|ubi dixit Iosue: " Quia turbasti nos, exturbet te Dominus in die hac ". Lapidavitque eum omnis Israel; et cuncta, quae illius erant, igne consumpta sunt.
JOSH|7|26|Congregaverunt quoque super eum acervum magnum lapidum, qui permanet usque in praesentem diem. Et aversus est furor Domini ab eis; vocatumque est nomen loci illius vallis Achor usque hodie.
JOSH|8|1|Dixit autem Dominus ad Iosue: " Ne timeas neque formides; tol le tecum omnem multitudinem pugnatorum et consurgens ascende in oppidum Hai: ecce tradidi in manu tua regem eius et populum urbemque et terram eius.
JOSH|8|2|Faciesque urbi Hai et regi eius, sicut fecisti Iericho et regi illius; praedam vero et omnia animantia diripietis vobis. Pone insidias urbi post eam ".
JOSH|8|3|Surrexitque Iosue et omnis exercitus bellatorum cum eo, ut ascenderent in Hai; et electa triginta milia virorum fortium misit nocte
JOSH|8|4|praecepitque eis dicens: "Collocamini in insidiis post civitatem nec longius recedatis ab illa; et eritis omnes parati.
JOSH|8|5|Ego autem et reliqua multitudo, quae mecum est, accedemus ex adverso contra urbem; cumque exierint contra nos sicut ante, fugiemus et terga vertemus,
JOSH|8|6|donec persequentes ab urbe longius protrahantur: putabunt enim nos fugere sicut prius.
JOSH|8|7|Nobis ergo fugientibus et illis sequentibus, consurgetis de insidiis et capietis civitatem; tradetque eam Dominus Deus vester in manus vestras.
JOSH|8|8|Cumque ceperitis, succendite eam; secundum verbum Domini facietis. Ecce mandavi vobis".
JOSH|8|9|Dimisitque eos, et perrexerunt ad insidiarum locum sederuntque inter Bethel et Hai ad occidentalem plagam urbis Hai. Iosue autem nocte illa in medio mansit populi.
JOSH|8|10|Surgensque diluculo recensuit populum et ascendit cum senioribus in fronte exercitus.
JOSH|8|11|Cumque omnes pugnatores cum eo ascendissent et appropinquassent civitati, steterunt ad septentrionalem urbis plagam, inter quam et eos vallis media erat.
JOSH|8|12|Et elegit fere quinque milia viros et posuit in insidiis inter Bethel et Hai ex occidentali parte eiusdem civitatis.
JOSH|8|13|Et posuit populus tota castra, quae erant in aquilone urbis, et agmen extremum ad occidentalem plagam urbis. Abiit ergo Iosue nocte illa et stetit in vallis medio.
JOSH|8|14|Quod cum vidisset rex Hai, festinavit mane et egressus est cum omni exercitu civitatis direxitque aciem contra Arabam ignorans quod post tergum laterent insidiae.
JOSH|8|15|Iosue vero et omnis Israel cesserunt loco simulantes metum et fugientes per solitudinis viam.
JOSH|8|16|Et convocatus est totus populus, qui erat in civitate, ad persequendum eos, et persecuti sunt eos. Cumque recessissent a civitate,
JOSH|8|17|et ne unus quidem in urbe Hai remansisset, qui non persequeretur Israel, et apertam urbem reliquissent,
JOSH|8|18|dixit Dominus ad Iosue: "Leva acinacem, quod in manu tua est, contra urbem Hai, quoniam tibi tradam eam ".
JOSH|8|19|Cumque elevasset acinacem ex adverso civitatis, insidiae, quae latebant, surrexerunt confestim et currentes ad civitatem ceperunt et cito succenderunt eam.
JOSH|8|20|Viri autem civitatis, qui persequebantur Iosue, respicientes et videntes fumum urbis ad caelum usque conscendere, non potuerunt ultra huc illucque diffugere, praesertim cum hi, qui simulaverant fugam et tendebant ad solitudinem, contra persequentes conversi essent.
JOSH|8|21|Vidensque Iosue et omnis Israel quod capta esset civitas, et fumus urbis ascenderet, reversi percusserunt viros Hai.
JOSH|8|22|Siquidem et illi, qui ceperant et succenderant civitatem, egressi sunt ex urbe in occursum eorum et hostes medios habuerunt. Cum ergo ex utraque parte adversarii caederentur, ita ut nullus de tanta multitudine salvaretur,
JOSH|8|23|regem quoque urbis Hai apprehenderunt viventem et obtulerunt Iosue.
JOSH|8|24|Igitur, omnibus habitatoribus Hai interfectis, qui Israelem ad deserta tendentem fuerant persecuti, et in eodem loco gladio corruentibus, reversi filii Israel percusserunt civitatem ore gladii.
JOSH|8|25|Erant autem, qui in eo die conciderant, a viro usque ad mulierem duodecim milia hominum omnes urbis Hai.
JOSH|8|26|Iosue vero non contraxit manum, quam in sublime porrexerat tenens acinacem, donec interficerentur omnes habitatores Hai.
JOSH|8|27|Iumenta tantum et praedam civitatis diviserunt sibi filii Israel, sicut praeceperat Dominus Iosue.
JOSH|8|28|Qui succendit urbem et fecit eam tumulum sempiternum, desolationem usque in praesentem diem.
JOSH|8|29|Regem quoque eius suspendit in ligno usque ad vesperum; et ad solis occasum praecepit Iosue, et deposuerunt cadaver eius de ligno proieceruntque in ipso introitu portae civitatis, congesto super eum magno acervo lapidum, qui permanet usque in praesentem diem.
JOSH|8|30|Tunc aedificavit Iosue altare Domino, Deo Israel, in monte Hebal,
JOSH|8|31|sicut praeceperat Moyses famulus Domini filiis Israel, et scriptum est in volumine legis Moysi, altare de lapidibus impolitis, quos ferrum non tetigit. Et obtulerunt super eo holocausta Domino immolaveruntque pacificas victimas.
JOSH|8|32|Et scripsit ibi super lapides exemplar legis Moysi, quod ille scripserat coram filiis Israel.
JOSH|8|33|Omnis autem populus et maiores natu praefectique ac iudices stabant ex utraque parte arcae in conspectu sacerdotum levitici generis, qui portabant arcam foederis Domini, ut advena ita et indigena. Media eorum pars iuxta montem Garizim et media iuxta montem Hebal, sicut praeceperat Moyses famulus Domini ad benedicendum populo Israel primum;
JOSH|8|34|post haec legit omnia verba legis, benedictionem et maledictionem, secundum cuncta, quae scripta erant in legis volumine.
JOSH|8|35|Nihil ex his, quae Moyses iusserat, omisit legere, sed universa replicavit coram omni congregatione Israel, mulieribus ac parvulis et advenis, qui inter eos morabantur.
JOSH|9|1|Quibus auditis, cuncti reges, qui trans Iordanem versabantur in montanis et in Sephela, in omni litore maris Magni, hi quoque, qui habitabant usque ad Libanum, Hetthaeus et Amorraeus, Chananaeus, Pherezaeus et Hevaeus et Iebusaeus
JOSH|9|2|congregati sunt pariter, ut pugnarent contra Iosue et Israel uno animo eademque sententia.
JOSH|9|3|At hi, qui habitabant in Gabaon, audientes cuncta, quae fecerat Iosue Iericho et Hai,
JOSH|9|4|et callide cogitantes tulerunt sibi cibaria, saccos veteres asinis imponentes et utres vinarios vetustos, scissos atque consutos,
JOSH|9|5|calceamentaque perantiqua, quae ad indicium vetustatis pittaciis consuta erant, induti veteribus vestimentis; panes quoque, quos portabant ob viaticum, duri erant et in frusta comminuti.
JOSH|9|6|Perrexeruntque ad Iosue, qui tunc morabatur in castris Galgalae, et dixerunt ei atque omni simul Israeli: " De terra longinqua venimus pactum vobiscum facere cupientes ". Responderuntque viri Israel ad Hevaeos atque dixerunt:
JOSH|9|7|" Ne forte in medio nostri habitetis, et non possimus foedus inire vobiscum ".
JOSH|9|8|At illi ad Iosue: " Servi, inquiunt, tui sumus ". Quibus Iosue ait: " Quinam estis et unde venistis? ".
JOSH|9|9|Responderunt: " De terra longinqua valde venerunt servi tui in nomine Domini Dei tui; audivimus enim famam potentiae eius, cuncta, quae fecit in Aegypto
JOSH|9|10|et duobus Amorraeorum regibus trans Iordanem, Sehon regi Hesebon et Og regi Basan, qui erat in Astharoth.
JOSH|9|11|Dixeruntque nobis seniores et omnes habitatores terrae nostrae: Tollite in manibus cibaria in viam et occurrite eis ac dicite: Servi vestri sumus; foedus inite nobiscum".
JOSH|9|12|En panes: quando egressi sumus de domibus nostris, ut veniremus ad vos, calidos sumpsimus; nunc sicci facti sunt et vetustate nimia comminuti.
JOSH|9|13|Utres vini novos implevimus, nunc rupti sunt et soluti; vestes et calceamenta, quibus induimur et quae habemus in pedibus, ob longitudinem largioris viae trita sunt et paene consumpta ".
JOSH|9|14|Susceperunt igitur viri de cibariis eorum et os Domini non interrogaverunt.
JOSH|9|15|Fecitque Iosue cum eis pacem et, inito foedere, pollicitus est quod viverent; principes quoque coetus iuraverunt eis.
JOSH|9|16|Post dies autem tres initi foederis, audierunt quod in vicino et inter eos habitarent.
JOSH|9|17|Moveruntque castra filii Israel et venerunt ad civitates eorum die tertio, quarum haec vocabula sunt: Gabaon et Cephira et Beroth et Cariathiarim;
JOSH|9|18|et non percusserunt eos filii Israel, eo quod iurassent eis principes coetus in nomine Domini, Dei Israel. Murmuravit itaque omnis coetus contra principes,
JOSH|9|19|qui responderunt eis: "Iuravimus illis in nomine Domini, Dei Israel, et idcirco non possumus eos contingere.
JOSH|9|20|Sed hoc faciemus eis: reserventur quidem, ut vivant, ne contra nos ira Domini concitetur, si peieraverimus;
JOSH|9|21|sed sic vivant, ut in usus universae multitudinis ligna caedant aquasque comportent ".Quibus haec loquentibus,
JOSH|9|22|vocavit Gabaonitas Iosue et dixit eis: " Cur nos decipere fraude voluistis, ut diceretis: "Procul valde habitamus a vobis", cum in medio nostri sitis?
JOSH|9|23|Itaque sub maledictione eritis, et non deficiet de stirpe vestra servus ligna caedens aquasque comportans in domum Dei mei".
JOSH|9|24|Qui responderunt: " Nuntiatum est nobis servis tuis, quod mandasset Dominus Deus tuus Moysi servo suo, ut traderet vobis omnem terram et disperderet cunctos habitatores eius; timuimus igitur valde pro animabus nostris, vestro terrore compulsi, et hoc consilium inivimus.
JOSH|9|25|Nunc autem in manu tua sumus: quod tibi bonum et rectum videtur, fac nobis ".
JOSH|9|26|Fecit ergo Iosue, ut dixerat, et liberavit eos de manu filiorum Israel, ut non occiderentur.
JOSH|9|27|Decrevitque in illo die esse eos in ministerium cuncti populi et altaris Domini caedentes ligna et aquas comportantes usque in praesens tempus pro loco, quem Dominus elegisset.
JOSH|10|1|Quae cum audisset Adonise dec rex Ierusalem, quod scili cet cepisset Iosue Hai et subvertisset eam - sicut enim fecerat Iericho et regi eius, sic fecit Hai et regi illius - et quod pacem fecissent Gabaonitae cum Israel et essent in medio eorum,
JOSH|10|2|timuerunt valde. Urbs enim magna erat Gabaon, sicut una regalium civitatum, et maior oppido Hai, omnesque viri eius bellatores fortissimi.
JOSH|10|3|Misit ergo Adonisedec rex Ierusalem ad Oham regem Hebron et ad Pharam regem Ierimoth, ad Iaphia quoque regem Lachis et ad Dabir regem Eglon dicens:
JOSH|10|4|" Ascendite ad me et ferte praesidium, ut expugnemus Gabaon, quia fecit pacem cum Iosue et filiis Israel ".
JOSH|10|5|Congregati igitur ascenderunt quinque reges Amorraeorum: rex Ierusalem, rex Hebron, rex Ierimoth, rex Lachis, rex Eglon simul cum exercitibus suis; et castrametati sunt circa Gabaon oppugnantes eam.
JOSH|10|6|Habitatores autem Gabaon miserunt ad Iosue, qui tunc morabatur in castris apud Galgalam, et dixerunt ei: " Ne retrahas manus tuas ab auxilio servorum tuorum! Ascende cito et libera nos ferque praesidium: convenerunt enim adversum nos omnes reges Amorraeorum, qui habitant in montanis ".
JOSH|10|7|Ascenditque Iosue de Galgalis, et omnis exercitus bellatorum cum eo, viri fortissimi.
JOSH|10|8|Dixitque Dominus ad Iosue: "Ne timeas eos! In manus enim tuas tradidi illos; nullus tibi ex eis resistere poterit ".
JOSH|10|9|Irruit itaque Iosue super eos repente tota ascendens nocte de Galgalis,
JOSH|10|10|et conturbavit eos Dominus a facie Israel; contrivitque plaga magna in Gabaon ac persecutus est per viam ascensus Bethoron et percussit usque Azeca et Maceda.
JOSH|10|11|Cumque fugerent filios Israel et essent in descensu Bethoron, Dominus misit super eos lapides magnos de caelo usque Azeca, et mortui sunt multo plures lapidibus grandinis, quam quos gladio percusserant filii Israel.
JOSH|10|12|Tunc locutus est Iosue Domino in die, qua tradidit Amorraeum in conspectu filiorum Israel, dixitque coram Israel: Sol, in Gabaon ne movearis,et luna, in valle Aialon ".
JOSH|10|13|Steteruntque sol et luna,donec ulcisceretur se gens de inimicis suis.Nonne scriptum est hoc in libro Iusti? Stetit itaque sol in medio caeli et non festinavit occumbere spatio unius fere diei.
JOSH|10|14|Non fuit antea et postea sicut dies illa, oboediente Domino voci hominis, quia Dominus pugnavit pro Israel.
JOSH|10|15|Reversusque est Iosue cum omni Israel in castra Galgalae.
JOSH|10|16|Fugerant autem quinque reges et se absconderant in spelunca urbis Maceda.
JOSH|10|17|Nuntiatumque est Iosue quod inventi essent quinque reges latentes in spelunca urbis Maceda.
JOSH|10|18|Qui praecepit: " Volvite saxa ingentia ad os speluncae et ponite viros, qui clausos custodiant.
JOSH|10|19|Vos autem nolite stare, sed persequimini hostes et extremos quoque fugientium caedite; ne dimittatis eos urbium suarum intrare praesidia, quia tradidit eos Dominus Deus vester in manus vestras ".
JOSH|10|20|Caesis igitur adversariis plaga maxima usque ad internecionem, ut reliquiae tantum ex eis effugere possent in civitates munitas,
JOSH|10|21|reversus est omnis exercitus ad Iosue in Maceda ad castra, sani et integri; nullusque contra filios Israel mutire ausus est.
JOSH|10|22|Praecepitque Iosue dicens: " Aperite os speluncae et producite ad me quinque reges, qui in ea latitant ".
JOSH|10|23|Feceruntque sic et eduxerunt ad eum quinque reges de spelunca: regem Ierusalem, regem Hebron, regem Ierimoth, regem Lachis, regem Eglon.
JOSH|10|24|Cumque educti essent ad eum, vocavit omnes viros Israel et ait ad principes exercitus, qui secum erant: "Accedite et ponite pedes super colla regum istorum". Qui cum accessissent et subiectorum colla pedibus calcarent,
JOSH|10|25|rursum ait ad eos: " Nolite timere nec paveatis; confortamini et estote robusti! Sic enim faciet Dominus cunctis hostibus vestris, adversum quos dimicatis ".
JOSH|10|26|Percussitque Iosue et interfecit eos atque suspendit super quinque ligna; fueruntque suspensi usque ad vesperum.
JOSH|10|27|Cumque occumberet sol, praecepit Iosue, ut deponerent eos de lignis; et depositos proiecerunt in speluncam, in qua latuerant, et posuerunt super os eius saxa ingentia, quae permanent usque in praesens.
JOSH|10|28|Eodem quoque die Macedam cepit Iosue et percussit eam in ore gladii regemque illius interfecit et omnes habitatores eius; non dimisit in ea ullas reliquias fecitque regi Maceda, sicut fecerat regi Iericho.
JOSH|10|29|Transivit cum omni Israel de Maceda in Lobna et pugnabat contra eam.
JOSH|10|30|Quam tradidit Dominus cum rege suo in manu Israel, percusseruntque urbem in ore gladii et omnes habitatores eius; non dimiserunt in ea ullas reliquias feceruntque regi Lobna, sicut fecerant regi Iericho.
JOSH|10|31|De Lobna transivit Iosue in Lachis cum omni Israel et, exercitu per gyrum disposito, oppugnabat eam.
JOSH|10|32|Tradiditque Dominus Lachis in manu Israel, qui cepit eam die altero; atque percussit in ore gladii omnemque animam, quae fuerat in ea, sicut fecerat Lobna.
JOSH|10|33|Eo tempore ascendit Horam rex Gazer, ut auxiliaretur Lachis; quem percussit Iosue cum omni populo eius usque ad internecionem.
JOSH|10|34|Transivitque de Lachis in Eglon cum omni Israel et circumdedit
JOSH|10|35|atque expugnavit eam eadem die percussitque in ore gladii omnes animas, quae erant in ea, iuxta omnia, quae fecerat Lachis.
JOSH|10|36|Ascendit quoque cum omni Israel de Eglon in Hebron et pugnavit contra eam.
JOSH|10|37|Cepitque eam et percussit in ore gladii, regem quoque eius et omnia oppida eius universasque animas, quae ibi fuerant commoratae; non reliquit ullas reliquias: sicut fecerat Eglon, sic fecit et Hebron, cuncta, quae in ea repperit, consumens gladio.
JOSH|10|38|Inde reversus cum omni Israel in Dabir oppugnavit
JOSH|10|39|et cepit eam; regem quoque eius et omnia oppida eius percussit in ore gladii; non dimisit in ea ullas reliquias: sicut fecerat Hebron et Lobna et regibus earum, sic fecit Dabir et regi illius.
JOSH|10|40|Percussit itaque Iosue omnem terram: montanam et Nageb atque Sephelam et declivia cum regibus suis; non dimisit in ea ullas reliquias, sed omne, quod spirare poterat, interfecit, sicut praeceperat Dominus, Deus Israel.
JOSH|10|41|Et percussit eos a Cadesbarne usque Gazam, omnem terram Gosen usque Gabaon,
JOSH|10|42|universosque reges et regiones eorum uno cepit impetu; Dominus enim, Deus Israel, pugnabat pro Israel.
JOSH|10|43|Reversusque est Iosue cum omni Israel ad locum castrorum in Galgala.
JOSH|11|1|Quae cum audisset Iabin rex Asor, misit ad Iobab regem Madon et ad regern Semeron atque ad regem Achsaph,
JOSH|11|2|ad reges quoque aquilonis, qui habitabant in montanis et in Araba contra meridiem Chenereth, in Sephela quoque et in regionibus Dor iuxta mare,
JOSH|11|3|Chananaeum in oriente et occidente, et Amorraeum atque Hetthaeum ac Pherezaeum et Iebusaeum in montanis, Hevaeum quoque, qui habitabat ad radices Hermon in terra Maspha.
JOSH|11|4|Egressique sunt omnes cum turmis suis, populus multus nimis sicut arena, quae est in litore maris, equi quoque et currus immensae multitudinis;
JOSH|11|5|conveneruntque omnes reges isti et castrametati sunt in unum ad aquas Merom, ut pugnarent contra Israel.
JOSH|11|6|Dixitque Dominus ad Iosue: "Ne timeas eos! Cras enim hac eadem hora ego tradam omnes istos occisos in conspectu Israel: equos eorum subnervabis et currus igne combures ".
JOSH|11|7|Venitque Iosue et omnis exercitus cum eo adversus illos ad aquas Merom subito, et irruerunt super eos.
JOSH|11|8|Tradiditque illos Dominus in manu Israel; qui percusserunt eos et persecuti sunt usque ad Sidonem magnam et Maserephoth in occidente campumque Maspha in oriente. Ita percussit omnes, ut nullas dimitteret ex eis reliquias;
JOSH|11|9|fecit sicut praeceperat ei Dominus: equos eorum subnervavit currusque combussit.
JOSH|11|10|Reversusque tempore illo cepit Asor et regem eius percussit gladio. Asor enim antiquitus inter omnia regna haec principatum tenebat.
JOSH|11|11|Percussitque omnes animas, quae ibidem morabantur; non dimisit in ea ullas reliquias, sed usque ad internecionem universa vastavit ipsamque urbem peremit incendio.
JOSH|11|12|Et omnes per circuitum civitates regesque earum cepit, percussit atque delevit, sicut praeceperat Moyses famulus Domini.
JOSH|11|13|Urbes tantum, quae erant in tumulis earum sitae, non succendit Israel; unam Asor solam Iosue flamma consumpsit.
JOSH|11|14|Omnemque praedam istarum urbium ac iumenta diviserunt sibi filii Israel, cunctis hominibus interfectis; nullum vivum reliquerunt.
JOSH|11|15|Sicut praeceperat Dominus Moysi servo suo, ita praecepit Moyses Iosue, et ille universa complevit; non praeteriit de universis mandatis ne unum quidem verbum, quod iusserat Dominus Moysi.
JOSH|11|16|Cepit itaque Iosue omnem terram hanc, montanam et Nageb terramque Gosen et Sephelam et Arabam montemque Israel et campestria eius,
JOSH|11|17|a monte Calvo, qui ascendit Seir, usque Baalgad in planitie Libani subter montem Hermon; omnes reges eorum cepit, percussit et occidit.
JOSH|11|18|Multo tempore pugnavit Iosue contra reges istos.
JOSH|11|19|Non fuit civitas, quae foedus iniret cum filiis Israel, praeter Hevaeum, qui habitabat in Gabaon: omnes bellando cepit.
JOSH|11|20|Domini enim sententia fuerat, ut indurarentur corda eorum, et pugnarent contra Israel et caderent et non mererentur ullam clementiam ac perirent, sicut praeceperat Dominus Moysi.
JOSH|11|21|In tempore illo venit Iosue et interfecit Enacim de montanis Hebron et Dabir et Anab et de omni monte Iudae et Israel urbesque eorum delevit.
JOSH|11|22|Non reliquit ullum de stirpe Enacim in terra filiorum Israel, absque civitatibus Gaza et Geth et Azoto, in quibus solis relicti sunt.
JOSH|11|23|Cepit ergo Iosue omnem terram, sicut locutus est Dominus ad Moysen, et tradidit eam in possessionem filiis Israel secundum partes et tribus suas; quievitque terra a proeliis.
JOSH|12|1|Hi sunt reges, quos percusserunt filii Israel et possederunt terram eorum trans Iordanem ad solis ortum, a torrente Arnon usque ad montem Hermon et omnem orientalem plagam Arabae.
JOSH|12|2|Sehon rex Amorraeorum, qui habitavit in Hesebon, dominatus est ab Aroer, quae sita est super ripam torrentis Arnon, et a media parte vallis et in dimidia parte Galaad usque ad torrentem Iaboc, qui est terminus filiorum Ammon;
JOSH|12|3|et in Araba usque ad mare Chenereth in oriente et usque ad mare Arabae, quod est mare Salsissimum, ad orientalem plagam in via, quae ducit Bethiesimoth, et in australi parte, quae iacet ad radices Phasga.
JOSH|12|4|Terminus Og regis Basan de reliquiis Raphaim, qui habitavit in Astharoth et in Edrai,
JOSH|12|5|et dominatus est in monte Hermon et in Salcha atque in universa Basan usque ad terminos Gesuri et Maachathi et in dimidia parte Galaad usque ad terminos Sehon regis Hesebon.
JOSH|12|6|Moyses famulus Domini et filii Israel percusserunt eos; tradiditque terram eorum Moyses in possessionem Rubenitis et Gaditis et dimidiae tribui Manasse.
JOSH|12|7|Hi sunt reges terrae, quos percussit Iosue et filii Israel trans Iordanem ad occidentalem plagam, a Baalgad in campo Libani usque ad montem Calvum, qui ascendit in Seir; tradiditque eam Iosue in possessionem tribubus Israel, singulis partes suas,
JOSH|12|8|tam in montanis quam in Sephela, in Araba et in declivibus et in solitudine ac in Nageb; Hetthaeus fuit et Amorraeus, Chananaeus et Pherezaeus, Hevaeus et Iebusaeus:
JOSH|12|9|rex Iericho unus, rex Hai, quae est ex latere Bethel, unus,
JOSH|12|10|rex Ierusalem unus, rex Hebron unus,
JOSH|12|11|rex Ierimoth unus, rex Lachis unus,
JOSH|12|12|rex Eglon unus, rex Gazer unus,
JOSH|12|13|rex Dabir unus, rex Gader unus,
JOSH|12|14|rex Horma unus, rex Arad unus,
JOSH|12|15|rex Lobna unus, rex Odollam unus,
JOSH|12|16|rex Maceda unus, rex Bethel unus,
JOSH|12|17|rex Thapphua unus, rex Opher unus,
JOSH|12|18|rex Aphec unus, rex Saron unus,
JOSH|12|19|rex Madon unus, rex Asor unus,
JOSH|12|20|rex Semeron unus, rex Achsaph unus,
JOSH|12|21|rex Thanach unus, rex Mageddo unus,
JOSH|12|22|rex Cedes unus, rex Iecnaam Carmeli unus,
JOSH|12|23|rex Dor et provinciae Dor unus, rex gentium Galgal unus,
JOSH|12|24|rex Thersa unus: omnes reges triginta unus.
JOSH|13|1|Iosue senex provectaeque aetatis erat, et dixit Dominus ad eum: " Senuisti et longaevus es; terraque latissima adhuc superest, quae necdum occupata est.
JOSH|13|2|Omnis videlicet Galilaea, regio Philisthim et universa Gesuri,
JOSH|13|3|a fluvio Sihor, qui est ad orientem Aegypti, usque ad terminos Accaron contra aquilonem, terra Chananaea, quae in quinque principes Philisthim dividitur, Gazaeos et Azotios, Ascalonitas, Getthaeos et Accaronitas ac Hevaei
JOSH|13|4|meridie; et omnis terra Chanaan de Ara Sidoniorum usque Apheca et terminos Amorraei;
JOSH|13|5|et terra Gibliorum et omnis Libanus in oriente a Baalgad sub monte Hermon usque ad introitum Emath,
JOSH|13|6|omnes, qui habitant in monte a Libano usque ad Maserephoth in occidente, universi Sidonii. Ego sum qui delebo eos a facie filiorum Israel. Sorte tantum distribue terram Israel in hereditatem, sicut praecepi tibi.
JOSH|13|7|Et nunc divide terram hanc in possessionem novem tribubus et dimidiae tribui Manasse ".
JOSH|13|8|Cum qua Ruben et Gad possederunt terram, quam tradidit eis Moyses famulus Domini trans fluenta Iordanis ad orientalem plagam:
JOSH|13|9|ab Aroer, quae sita est in ripa torrentis Arnon, et civitate in vallis medio, universaque campestria Medaba usque Dibon;
JOSH|13|10|et cunctas civitates Sehon regis Amorraei, qui regnavit in Hesebon, usque ad terminos filiorum Ammon;
JOSH|13|11|et Galaad ac terminos Gesuri et Maachathi omnemque montem Hermon et universam Basan usque Salcha,
JOSH|13|12|omne regnum Og in Basan, qui regnavit in Astharoth et Edrai - ipse fuit de reliquiis Raphaim C; percussitque eos Moyses atque delevit.
JOSH|13|13|Non autem disperdiderunt filii Israel Gesuri et Maachathi, et habitaverunt in medio Israel usque in praesentem diem.
JOSH|13|14|Tribui tantum Levi non dedit possessionem, sed sacrificia Domini, Dei Israel: ipsa est eius hereditas, sicut locutus est illi.
JOSH|13|15|Dedit ergo Moyses possessionem tribui filiorum Ruben iuxta cognationes suas.
JOSH|13|16|Fuitque terminus eorum ab Aroer, quae sita est in ripa torrentis Arnon, et a civitate in valle eiusdem torrentis media, et universa planities usque Medaba,
JOSH|13|17|Hesebon cunctaque oppida eius, quae sunt in campestribus: Dibon et Bamothbaal et Bethbaalmeon
JOSH|13|18|et Iasa et Cademoth et Mephaath,
JOSH|13|19|Cariathaim et Sabama et Serethsahar in monte convallis,
JOSH|13|20|Bethphegor et declivia Phasga et Bethiesimoth
JOSH|13|21|et omnes urbes campestres universumque regnum Sehon regis Amorraei, qui regnavit in Hesebon, quem percussit Moyses, ipsum et principes Madian, Evi et Recem et Sur et Hur et Rebe, duces Sehon habitatores terrae.
JOSH|13|22|Et Balaam filium Beor hariolum occiderunt filii Israel gladio cum ceteris interfectis.
JOSH|13|23|Factusque est terminus filiorum Ruben Iordanis fluvius. Haec est possessio Rubenitarum per cognationes suas, urbes et viculi earum.
JOSH|13|24|Deditque Moyses tribui Gad, filiis Gad, per cognationes suas possessionem, cuius hic est
JOSH|13|25|terminus: Iazer et omnes civitates Galaad dimidiaque pars terrae filiorum Ammon usque ad Aroer, quae est contra Rabba;
JOSH|13|26|et ab Hesebon usque Ramothmaspha et Betonim et a Mahanaim usque ad terminos Lodabar,
JOSH|13|27|in valle quoque Betharan et Bethnemra et Succoth et Saphon, reliqua pars regni Sehon regis Hesebon; Iordanis et terminus usque ad extremam partem maris Chenereth trans Iordanem ad orientalem plagam.
JOSH|13|28|Haec est possessio filiorum Gad per familias suas, civitates et villae earum.
JOSH|13|29|Dedit Moyses et dimidiae tribui filiorum Manasse, iuxta cognationes suas possessionem:
JOSH|13|30|Manasse, a Mahanaim universam Basan, cunctum regnum Og regis Basan omnesque vicos Iair, qui sunt in Basan, sexaginta oppida;
JOSH|13|31|et dimidiam partem Galaad et Astharoth et Edrai, urbes regni Og in Basan, filiis Machir filii Manasse, dimidiae parti filiorum Machir, iuxta cognationes suas.
JOSH|13|32|Hanc possessionem divisit Moyses in campestribus Moab trans Iordanem contra Iericho ad orientalem plagam.
JOSH|13|33|Tribui autem Levi non dedit possessionem, quoniam Dominus, Deus Israel, ipse est possessio eius, ut locutus est illi.
JOSH|14|1|Hoc est, quod hereditave runt filii Israel in terra Cha naan, quod dederunt eis Eleazar sacerdos et Iosue filius Nun et principes familiarum tribuum Israel,
JOSH|14|2|sorte omnia dividentes, sicut praeceperat Dominus in manu Moysi, novem tribubus et dimidiae tribui.
JOSH|14|3|Duabus enim tribubus et dimidiae dederat Moyses trans Iordanem possessionem, absque Levitis, quibus nihil dedit inter fratres suos;
JOSH|14|4|sed sunt filii Ioseph in duas divisi tribus, Manasse et Ephraim, nec acceperunt Levitae aliam in terra partem, nisi urbes ad habitandum et suburbana earum ad alenda iumenta et pecora sua.
JOSH|14|5|Sicut praeceperat Dominus Moysi, ita fecerunt filii Israel et diviserunt terram.
JOSH|14|6|Accesserunt itaque filii Iudae ad Iosue in Galgala, locutusque est ad eum Chaleb filius Iephonne Cenezaeus: " Nosti quid locutus sit Dominus ad Moysen hominem Dei de me et te in Cadesbarne.
JOSH|14|7|Quadraginta annorum eram, quando me misit Moyses famulus Domini de Cadesbarne, ut considerarem terram; nuntiavique ei quod mihi verum videbatur.
JOSH|14|8|Fratres autem mei, qui ascenderant mecum, dissolverunt cor populi, et nihilominus ego adimplevi, ut sequerer Dominum Deum meum.
JOSH|14|9|Iuravitque Moyses in die illo dicens: "Terra, quam calcavit pes tuus, erit possessio tua et filiorum tuorum in aeternum, quia adimplevisti, ut sequereris Dominum Deum meum".
JOSH|14|10|Concessit ergo Dominus vitam mihi, sicut pollicitus est, usque in praesentem diem. Quadraginta et quinque anni sunt ex quo locutus est Dominus verbum istud ad Moysen, quando ambulabat Israel per solitudinem; hodie octoginta quinque annorum sum,
JOSH|14|11|sic valens ut eo valebam tempore, quando ad explorandum missus sum; illius in me temporis fortitudo usque hodie perseverat tam ad bellandum quam ad gradiendum.
JOSH|14|12|Da ergo mihi montem istum, quem pollicitus est Dominus die illo, te quoque audiente quod Enacim ibi sunt et urbes magnae atque munitae; si forte sit Dominus mecum, et potuero delere eos, sicut promisit mihi ".
JOSH|14|13|Benedixitque ei Iosue et tradidit Hebron in possessionem;
JOSH|14|14|atque ex eo fuit Hebron Chaleb filio Iephonne Cenezaeo usque in praesentem diem, quia adimplevit, ut sequeretur Dominum, Deum Israel.
JOSH|14|15|Nomen Hebron antea vocabatur Cariatharbe (id est civitas Arbe), hominis maximi inter Enacim. Et terra cessavit a proeliis.
JOSH|15|1|Sors tribus filiorum Iudae per cognationes suas ista fuit: usque ad terminum Edom, ad desertum Sin contra Nageb, usque ad extremam partem australis plagae.
JOSH|15|2|Terminus eius meridionalis a summitate maris Salsissimi et a lingua eius, quae respicit meridiem.
JOSH|15|3|Egrediturque contra ascensum Acrabbim et pertransit in Sin ascenditque in meridie Cadesbarne et pervenit in Esron ascendens ad Addar et vertitur in Carca;
JOSH|15|4|atque inde pertransiens in Asemona pervenit ad torrentem Aegypti; eruntque exitus eius ad mare Magnum: hic erit vobis finis meridianae plagae.
JOSH|15|5|Ab oriente vero terminus erit mare Salsissimum usque ad extrema Iordanis. Terminus aquilonis a lingua maris et ab extremis Iordanis
JOSH|15|6|ascendit in Bethagla et transit ab aquilone Betharaba ascendens ad lapidem Boen filii Ruben
JOSH|15|7|et ascendens ad Dabir de valle Achor et contra aquilonem vergens ad Galiloth (hi sunt circuli), qui sunt ex adverso ascensionis Adommim, quae est ab australi parte torrentis, transit ad aquas, quae vocantur fons Solis, et erunt exitus eius ad fontem Rogel.
JOSH|15|8|Ascenditque per convallem Benennom ex latere Iebusaei ad meridiem - haec est Ierusalem - et inde se erigens ad verticem montis, qui est contra vallem Ennom ad occidentem in extrema parte vallis Raphaim contra aquilonem;
JOSH|15|9|pertransitque a vertice montis usque ad fontem aquae Nephtoa et pervenit usque ad vicos montis Ephron inclinaturque in Baala, quae est Cariathiarim.
JOSH|15|10|Et vergit de Baala contra occidentem usque ad montem Seir transitque iuxta latus montis Iarim ad aquilonem - id est Cheslon - et descendit in Bethsames transitque in Thamna
JOSH|15|11|et pervenit ad latus septentrionale Accaron inclinaturque in Sechron et transit montem Baala pervenitque in Iebneel et finitur mari. Terminus occidentalis est mare Magnum.
JOSH|15|12|Hi sunt termini filiorum Iudae per circuitum in cognationibus suis.
JOSH|15|13|Chaleb vero filio Iephonne dedit partem in medio filiorum Iudae, sicut praeceperat Dominus Iosue: Cariatharbe (id est civitas Arbe), patris Enac, ipsa est Hebron.
JOSH|15|14|Delevitque ex ea Chaleb tres filios Enac: Sesai et Ahiman et Tholmai de stirpe Enac.
JOSH|15|15|Atque inde conscendens venit ad habitatores Dabir, quae prius vocabatur Cariathsepher (id est civitas Litterarum).
JOSH|15|16|Dixitque Chaleb: " Qui percusserit Cariathsepher et ceperit eam, dabo illi Axam filiam meam uxorem ".
JOSH|15|17|Cepitque eam Othoniel filius Cenez frater Chaleb, deditque ei Axam filiam suam uxorem.
JOSH|15|18|Quae cum veniret, suasit viro suo, ut peteret a patre suo agrum; descenditque de asino. Cui Chaleb: " Quid habes? ", inquit.
JOSH|15|19|At illa respondit: " Da mihi benedictionem. Terram Nageb arentem dedisti mihi; iunge et irriguam ". Dedit itaque ei Chaleb irriguum superius et inferius.
JOSH|15|20|Haec est possessio tribus filiorum Iudae per cognationes suas.
JOSH|15|21|Erantque civitates ab extremis partibus filiorum Iudae iuxta terminos Edom in Nageb: Cabseel et Eder et Iagur
JOSH|15|22|et Cina et Dimona et Adada
JOSH|15|23|et Cades et Asor et Iethnan,
JOSH|15|24|Ziph et Telem et Baloth
JOSH|15|25|et Asorhadatta et Carioth, Esron - haec est Asor -
JOSH|15|26|Amam et Sama et Molada
JOSH|15|27|et Asargadda et Hasemon et Bethphelet
JOSH|15|28|et Asarsual et Bersabee et Baziothia,
JOSH|15|29|Baala et Iim et Esem
JOSH|15|30|et Eltholad et Cesil et Horma
JOSH|15|31|et Siceleg et Madmena et Sensenna
JOSH|15|32|et Lebaoth et Selim et Enremmon: omnes civitates viginti novem et villae earum.
JOSH|15|33|In campestribus vero: Esthaol et Saraa et Asena
JOSH|15|34|et Zanoa et Engannim, Thapphua et Enaim,
JOSH|15|35|Ierimoth et Odollam, Socho et Azeca
JOSH|15|36|et Saarim et Adithaim et Gedera et Gederothaim: urbes quattuordecim et villae earum.
JOSH|15|37|Sanan et Hadasa et Magdalgad
JOSH|15|38|et Delean et Maspha et Iecethel,
JOSH|15|39|Lachis et Bascath et Eglon
JOSH|15|40|et Chebbon et Lehemas et Cethlis
JOSH|15|41|et Gederoth, Bethdagon et Naama et Maceda: civitates sedecim et villae earum.
JOSH|15|42|Lobna et Ether et Asan
JOSH|15|43|et Iephtha et Esna et Nesib
JOSH|15|44|et Ceila et Achzib et Maresa: civitates novem et villae earum.
JOSH|15|45|Accaron cum filiabus et villulis suis;
JOSH|15|46|ab Accaron usque ad mare: omnia, quae sunt ad latus Azoti, et viculos eorum,
JOSH|15|47|Azotus cum filiabus et villulis suis, Gaza cum filiabus et villulis suis usque ad torrentem Aegypti, et mare Magnum terminus.
JOSH|15|48|Et in monte: Samir et Iether et Socho
JOSH|15|49|et Danna et Cariathsenna - haec est Dabir -
JOSH|15|50|et Anab et Esthemo et Anim
JOSH|15|51|et Gosen et Helon et Gilo: civitates undecim et villae earum.
JOSH|15|52|Arab et Duma et Esaan
JOSH|15|53|et Ianum et Beththapphua et Apheca
JOSH|15|54|et Ammatha et Cariatharbe - haec est Hebron - et Sior: civitates novem et villae earum.
JOSH|15|55|Maon et Carmel et Ziph et Iutta
JOSH|15|56|et Iezrahel et Iucadam et Zanoa,
JOSH|15|57|Accain, Gabaa et Thamna: civitates decem et villae earum.
JOSH|15|58|Halhul, Bethsur et Gedor
JOSH|15|59|et Mareth et Bethanoth et Eltecon: civitates sex et villae earum. Thecue et Ephratha - haec est Bethlehem - et Phegor et Etam et Culon et Tatam et Sores et Carem et Gallim et Bether et Manahath: civitates undecim et villae earum.
JOSH|15|60|Cariathbaal - haec est Cariathiarim (urbs Silvarum) - et Arebba: civitates duae et villae earum.
JOSH|15|61|In deserto: Betharaba, Meddin et Sachacha
JOSH|15|62|et Nebsan et civitas Salis et Engaddi: civitates sex et villae earum.
JOSH|15|63|Iebusaeum autem habitatorem Ierusalem non potuerunt filii Iudae delere; habitavitque Iebusaeus cum filiis Iudae in Ierusalem usque in praesentem diem.
JOSH|16|1|Cecidit quoque sors filiorum Ioseph ab Iordane contra Ie richo et aquas eius ab oriente, solitudo, quae ascendit de Iericho ad montem Bethel
JOSH|16|2|et egreditur de Bethel Luz transitque per terminum Arachitarum in Ataroth
JOSH|16|3|et descendit ad occidentem ad terminum Iephlethi usque ad terminos Bethoron inferioris et Gazer; finiunturque regiones eius mari Magno.
JOSH|16|4|Hereditaverunt illas filii Ioseph Manasses et Ephraim.
JOSH|16|5|Et factus est terminus filiorum Ephraim per cognationes suas et possessio eorum contra orientem Atarothaddar usque Bethoron superiorem;
JOSH|16|6|egrediunturque confinia in mare, Machmethath vero aquilonem respicit et vertitur terminus contra orientem in Thanathselo et pertransit ab oriente Ianoe.
JOSH|16|7|Descenditque de Ianoe in Ataroth et Naaratha et pervenit in Iericho et egreditur ad Iordanem.
JOSH|16|8|De Thapphua pertransit terminus ad occidentem ad torrentem Cana, suntque egressus eius in mare: haec est possessio tribus filiorum Ephraim per familias suas,
JOSH|16|9|urbesque separatae filiis Ephraim in medio possessionis filiorum Manasse, omnes urbes et villae earum.
JOSH|16|10|Et non interfecerunt filii Ephraim Chananaeum, qui habitabat in Gazer; habitavitque Chananaeus in medio Ephraim usque in diem hanc et factus est tributarius.
JOSH|17|1|Cecidit autem sors tribui Manasse - ipse est enim pri mogenitus Ioseph C; Machir primogenito Manasse patri Galaad, quia fuit vir pugnator, accepit in possessionem Galaad et Basan.
JOSH|17|2|Et reliqui filiorum Manasse acceperunt iuxta familias suas: filii Abiezer et filii Helec et filii Asriel et filii Sechem et filii Hepher et filii Semida: isti sunt filii Manasse filii Ioseph, mares per cognationes suas.
JOSH|17|3|Salphaad vero filio Hepher filii Galaad filii Machir filii Manasse non erant filii, sed solae filiae, quarum ista sunt nomina: Maala et Noa, Hegla et Melcha et Thersa.
JOSH|17|4|Veneruntque in conspectu Eleazari sacerdotis et Iosue filii Nun et principum dicentes: " Dominus praecepit per manum Moysi, ut daretur nobis possessio in medio fratrum nostrorum ". Deditque eis iuxta imperium Domini possessionem in medio fratrum patris earum.
JOSH|17|5|Et ceciderunt funiculi Manasse decem, absque terra Galaad et Basan trans Iordanem.
JOSH|17|6|Filiae enim Manasse acceperunt hereditatem in medio filiorum eius. Terra autem Galaad cecidit in sortem filiorum Manasse, qui reliqui erant.
JOSH|17|7|Fuitque terminus Manasse ab Aser: Machmethath, quae respicit Sichem et egreditur ad dextram in Iasib apud fontem Thapphuae.
JOSH|17|8|Etenim in sorte Manasse ceciderat terra Thapphuae; Thapphua autem ipsa, quae est iuxta terminos Manasse, fuit filiis Ephraim.
JOSH|17|9|Descenditque terminus ad torrentem Cana. In meridie torrentis civitates sunt Ephraim in medio urbium Manasse. Terminus Manasse est ab aquilone torrentis, et exitus eius pergit ad mare,
JOSH|17|10|ita ut ab austro sit possessio Ephraim et ab aquilone Manasse, et utramque claudat mare, et attingunt tribum Aser ab aquilone et tribum Issachar ab oriente.
JOSH|17|11|Fuitque hereditas Manasse in Issachar et in Aser: Bethsan et filiae eius et Ieblaam cum filiabus suis et habitatores Dor cum filiabus suis, habitatores quoque Endor cum filiabus suis; similiterque habitatores Thanach cum filiabus suis et habitatores Mageddo cum filiabus suis et tertia pars regionis Nopheth.
JOSH|17|12|Nec potuerunt filii Manasse has occupare civitates, sed Chananaeus permansit in terra ista.
JOSH|17|13|Postquam autem convaluerunt filii Israel, subiecerunt Chananaeos et fecerunt sibi tributarios nec expulerunt eos.
JOSH|17|14|Locutique sunt filii Ioseph ad Iosue atque dixerunt: " Quare dedisti mihi possessionem sortis et funiculi unius, cum sim tantae multitudinis et benedixerit mihi Dominus? ".
JOSH|17|15|Ad quos Iosue ait: " Si populus multus es, ascende in silvam et succide tibi spatia in terra Pherezaei et Raphaim, quia angusta est tibi possessio montis Ephraim ".
JOSH|17|16|Cui responderunt filii Ioseph: " Montana non sufficiunt nobis, et ferreis curribus utuntur omnes Chananaei, qui habitant in terra campestri, Bethsan cum filiabus suis et illi, qui sunt in planitie Iezrahel ".
JOSH|17|17|Dixitque Iosue ad domum Ioseph, Ephraim et Manasse: "Populus multus es et magnae fortitudinis; non habebis sortem unam,
JOSH|17|18|sed transibis ad montem et succides tibi atque purgabis ad habitandum spatia; et poteris ultra procedere cum subverteris Chananaeum, qui ferreos habet currus et est fortis ".
JOSH|18|1|Congregatique sunt omnes filii Israel in Silo ibique fixe runt tabernaculum conventus, et fuit eis terra subiecta.
JOSH|18|2|Remanserant autem filiorum Israel septem tribus, quae necdum acceperant possessiones suas.
JOSH|18|3|Ad quos Iosue ait: " Usquequo marcetis ignavia et non intratis ad possidendam terram, quam Dominus, Deus patrum vestrorum,dedit vobis?
JOSH|18|4|Eligite de singulis tribubus ternos viros, ut mittam eos, et surgant atque circumeant terram et describant eam iuxta numerum uniuscuiusque multitudinis referantque ad me, quod descripserint.
JOSH|18|5|Dividite vobis terram in septem partes: Iudas sit in terminis suis in australi plaga, et domus Ioseph in aquilone.
JOSH|18|6|Reliquam terram in septem partes describite; et huc afferetis ad me, ut coram Domino Deo nostro mittam vobis hic sortem,
JOSH|18|7|quia non est inter vos pars Levitarum, sed sacerdotium Domini est eorum hereditas. Gad autem et Ruben et dimidia tribus Manasse iam acceperant possessiones suas trans Iordanem ad orientalem plagam, quas dedit eis Moyses famulus Domini ".
JOSH|18|8|Cumque surrexissent viri, ut pergerent ad describendam terram, praecepit eis Iosue dicens: "Circuite terram et describite eam ac revertimini ad me, ut hic coram Domino in Silo mittam vobis sortem ".
JOSH|18|9|Itaque perrexerunt et lustrantes terram secundum urbes in septem partes diviserunt scribentes in volumine; reversique sunt ad Iosue in castra Silo.
JOSH|18|10|Qui misit eis sortes coram Domino in Silo divisitque ibi terram filiis Israel secundum partes eorum.
JOSH|18|11|Et ascendit sors prima filiorum Beniamin per familias suas, ut possiderent terram inter filios Iudae et filios Ioseph.
JOSH|18|12|Fuitque terminus eorum contra aquilonem a Iordane pergens iuxta latus Iericho septentrionalis plagae et inde contra occidentem ad montana conscendens et perveniens in solitudinem Bethaven;
JOSH|18|13|atque pertransiens iuxta Luzam ad meridiem - ipsa est Bethel - descendit in Atarothaddar in montem, qui est ad meridiem Bethoron inferioris,
JOSH|18|14|et inclinatur vergens contra mare ad meridiem a monte, qui respicit Bethoron contra meridiem; suntque exitus eius in Cariathbaal, quae vocatur et Cariathiarim, urbem filiorum Iudae. Haec est plaga ad occidentem.
JOSH|18|15|In plaga autem ad meridiem, ex parte Cariathiarim egreditur terminus in Gasim et pervenit usque ad fontem aquarum Nephtoa
JOSH|18|16|descenditque in extremam partem montis, qui respicit vallem Benennom et est contra septentrionalem plagam in extrema parte vallis Raphaim; descenditque in vallem Ennom, iuxta latus Iebusaei ad austrum, et pervenit ad fontem Rogel
JOSH|18|17|transiens ad aquilonem et egrediens ad Ensemes (id est fontem Solis). Et pertransit usque ad Galiloth (hi sunt circuli), qui sunt e regione ascensus Adommim, descenditque ad Abenboen (id est lapidem Boen) filii Ruben
JOSH|18|18|et pertransit ex latere aquilonis Betharaba descenditque in Arabam.
JOSH|18|19|Et praetergreditur contra aquilonem Bethagla; suntque exitus eius contra linguam maris Salsissimi ab aquilone in fine Iordanis. Haec est australis plaga.
JOSH|18|20|Iordanis autem est terminus ab oriente. Haec est possessio filiorum Beniamin per terminos suos in circuitu secundum familias suas.
JOSH|18|21|Fueruntque civitates eius: Iericho et Bethagla et Ameccasis
JOSH|18|22|et Betharaba et Semaraim et Bethel
JOSH|18|23|et Avim et Phara et Ophra,
JOSH|18|24|Capharemona et Ophni et Gabaa: civitates duodecim et villae earum.
JOSH|18|25|Gabaon et Rama et Beroth
JOSH|18|26|et Maspha et Cephira et Mosa
JOSH|18|27|et Recem, Iaraphel et Tharala
JOSH|18|28|et Sela, Eleph et Iebus, quae est Ierusalem, Gabaath et Cariath: civitates quattuordecim et villae earum. Haec est possessio filiorum Beniamin iuxta familias suas.
JOSH|19|1|Et egressa est sors secunda fi liorum Simeon per cognatio nes suas; fuitque hereditas
JOSH|19|2|eorum in medio possessionis filiorum Iudae. Bersabee et Sama et Molada
JOSH|19|3|et Asarsual et Bala et Esem
JOSH|19|4|et Eltholad et Bethul et Horma
JOSH|19|5|et Siceleg et Bethmarchaboth et Asarsusa
JOSH|19|6|et Bethlebaoth et Sarohen: civitates tredecim et villae earum.
JOSH|19|7|Ain et Remmon et Ethar et Asan: civitates quattuor et villae earum.
JOSH|19|8|Omnes viculi per circuitum urbium istarum usque ad Baalathbeer, Ramathnageb: haec est hereditas filiorum Simeon iuxta cognationes suas.
JOSH|19|9|Sumpta est de funiculo filiorum Iudae, quia maior erat; et idcirco possederunt filii Simeon in medio hereditatis eorum.
JOSH|19|10|Ceciditque sors tertia filiorum Zabulon per cognationes suas. Et factus est terminus possessionis eorum usque Sarid
JOSH|19|11|ascenditque contra occidentem et Merala et pervenit in Debbaseth usque ad torrentem, qui est contra Iecnaam,
JOSH|19|12|et revertitur de Sarid contra orientem in fines Ceseleththabor et egreditur ad Dabereth ascenditque contra Iaphia.
JOSH|19|13|Et inde pertransit usque ad orientalem plagam Gethhepher, Etthacasin et egreditur in Remmon et inclinatur in Noa;
JOSH|19|14|et vergit ad aquilonem ad Hanathon. Suntque egressus eius vallis Iephthael;
JOSH|19|15|et Cateth et Naalol et Semeron et Iedala et Bethlehem: civitates duodecim et villae earum.
JOSH|19|16|Haec est hereditas tribus filiorum Zabulon per cognationes suas, urbes et viculi earum.
JOSH|19|17|Issachar egressa est sors quarta per cognationes suas.
JOSH|19|18|Fuitque eius hereditas Iezrahel et Chasaloth et Sunam
JOSH|19|19|et Hapharaim et Seon et Anaharath
JOSH|19|20|et Rabbith et Cesion et Abes
JOSH|19|21|et Rameth et Engannim et Enhadda et Bethpheses.
JOSH|19|22|Et pervenit terminus eius usque Thabor et Sehesima et Bethsames; suntque exitus eius ad Iordanem; civitates sedecim et villae earum.
JOSH|19|23|Haec est possessio filiorum Issachar per cognationes suas, urbes et viculi earum.
JOSH|19|24|Ceciditque sors quinta tribui filiorum Aser per cognationes suas.
JOSH|19|25|Fuitque terminus eorum Helcath et Chali et Beten et Achsaph
JOSH|19|26|et Elmelech et Amaad et Masal et pervenit usque ad Carmelum in occidente et ad Sihorlabanath;
JOSH|19|27|ac revertitur contra orientem in Bethdagon et pertransit usque Zabulon et vallem Iephthael contra aquilonem in Bethemec et Neiel. Egrediturque ad laevam Chabul
JOSH|19|28|et Abran et Rohob et Hamon et Cana usque ad Sidonem magnam
JOSH|19|29|revertiturque in Rama usque ad civitatem munitissimam Tyrum et revertitur in Hosa; suntque exitus eius in mare; Mahaleb, Achazib
JOSH|19|30|et Amma et Aphec et Rohob: civitates viginti duae et villae earum.
JOSH|19|31|Haec est possessio filiorum Aser per cognationes suas, urbes et viculi earum.
JOSH|19|32|Filiorum Nephthali sexta sors cecidit per familias suas.
JOSH|19|33|Et coepit terminus de Heleph et de quercu in Saananim et Adamineceb et Iebnael usque Lecum et egressus eius usque ad Iordanem;
JOSH|19|34|revertiturque terminus contra occidentem in Aznotthabor atque inde egreditur in Hucoc et attingit Zabulon contra meridiem et Aser contra occidentem et Iordanem contra ortum solis;
JOSH|19|35|civitates munitissimae Assedim, Ser et Ammath, Reccath et Chenereth
JOSH|19|36|et Edema et Rama, Asor
JOSH|19|37|et Cedes et Edrai et Enasor,
JOSH|19|38|Ieron et Magdalel, Horem et Bethanath et Bethsames: civitates decem et novem et villae earum.
JOSH|19|39|Haec est possessio tribus filiorum Nephthali per cognationes suas, urbes et viculi earum.
JOSH|19|40|Tribui filiorum Dan per familias suas egressa est sors septima.
JOSH|19|41|Et fuit terminus possessionis eius Saraa et Esthaol et Hirsemes (id est civitas Solis)
JOSH|19|42|et Selebin et Aialon et Iethela
JOSH|19|43|et Elon et Thamna et Accaron
JOSH|19|44|et Elthece et Gebbethon et Baalath
JOSH|19|45|et Iud et Benebarach et Gethremmon
JOSH|19|46|et Meiarcon et Areccon cum termino, qui respicit Ioppen.
JOSH|19|47|Et terminus filiorum Dan effugit ab eis. Ascenderuntque filii Dan et pugnaverunt contra Lesem ceperuntque eam; et percusserunt in ore gladii ac possederunt et habitaverunt in ea, vocantes Lesemdan ex nomine Dan patris sui.
JOSH|19|48|Haec est possessio tribus filiorum Dan per cognationes suas, urbes et viculi earum.
JOSH|19|49|Cumque complessent terram sorte dividere singulis per tribus suas, dederunt filii Israel possessionem Iosue filio Nun in medio sui,
JOSH|19|50|iuxta praeceptum Domini, urbem quam postulavit: Thamnathsare in monte Ephraim. Et aedificavit civitatem habitavitque in ea.
JOSH|19|51|Hae sunt possessiones, quas sorte diviserunt Eleazar sacerdos et Iosue filius Nun et principes familiarum tribuum filiorum Israel in Silo coram Domino ad ostium tabernaculi conventus; compleveruntque partiri terram.
JOSH|20|1|Et locutus est Dominus ad Iosue dicens: " Loquere filiis Israel et dic eis:
JOSH|20|2|Separate vobis urbes fugitivorum, de quibus locutus sum ad vos per manum Moysi,
JOSH|20|3|ut confugiat ad eas, quicumque animam percusserit per errorem nescius, et possit evadere iram proximi, qui ultor est sanguinis.
JOSH|20|4|Cum ad unam harum confugerit civitatum, stabit ante portam civitatis et loquetur senioribus urbis illius ea, quae se comprobent innocentem; sicque suscipient eum et dabunt ei locum ad habitandum.
JOSH|20|5|Cumque ultor sanguinis eum fuerit persecutus, non tradent in manus eius, quia ignorans percussit proximum suum nec ante biduum triduumve eius probatur inimicus.
JOSH|20|6|Et habitabit in civitate illa, donec stet ante coetum ad iudicium, causam reddens facti sui, donec moriatur sacerdos magnus, qui fuerit in illo tempore. Tunc revertetur homicida et ingredietur civitatem suam et domum suam, de qua fugerat ".
JOSH|20|7|Decreveruntque Cedes in Galilaea montis Nephthali et Sichem in monte Ephraim et Cariatharbe - ipsa est Hebron - in monte Iudae;
JOSH|20|8|et trans Iordanem contra orientalem plagam Iericho statuerunt Bosor, quae sita est in campestri solitudine de tribu Ruben, et Ramoth in Galaad de tribu Gad et Golan in Basan de tribu Manasse.
JOSH|20|9|Hae civitates constitutae sunt cunctis filiis Israel et advenis, qui habitant inter eos, ut fugeret ad eas, qui animam nescius percussisset et non moreretur in manu proximi effusum sanguinem vindicare cupientis, donec staret ante populum expositurus causam suam.
JOSH|21|1|Accesseruntque principes familiarum Levi ad Eleazarum sacerdotem et Iosue filium Nun et ad duces cognationum per singulas tribus filiorum Israel
JOSH|21|2|locutique sunt ad eos in Silo terrae Chanaan atque dixerunt: " Dominus praecepit per manum Moysi, ut darentur nobis urbes ad habitandum et suburbana earum ad alenda iumenta ".
JOSH|21|3|Dederuntque filii Israel Levitis de possessionibus suis, iuxta imperium Domini, civitates illas et suburbana earum.
JOSH|21|4|Egressaque est sors in familias Caath: et acceperunt filii Aaron sacerdotis de tribubus Iudae et Simeon et Beniamin civitates tredecim.
JOSH|21|5|Et reliqui filiorum Caath, id est Levitae, acceperunt de tribubus Ephraim et Dan et dimidia tribu Manasse civitates decem.
JOSH|21|6|Porro filiis Gerson egressa est sors, ut acciperent de tribubus Issachar et Aser et Nephthali dimidiaque tribu Manasse in Basan civitates numero tredecim.
JOSH|21|7|Et filiis Merari per cognationes suas de tribubus Ruben et Gad et Zabulon urbes duodecim.
JOSH|21|8|Dederuntque filii Israel Levitis civitates illas et suburbana earum, sicut praecepit Dominus per manum Moysi, singulis sorte tribuentes.
JOSH|21|9|De tribubus filiorum Iudae et Simeon dederunt civitates, quarum ista sunt nomina,
JOSH|21|10|filiis Aaron ex familiis Caath levitici generis - prima enim sors illis egressa est C:
JOSH|21|11|Cariatharbe (id est civitas Arbe), patris Enac, quae vocatur Hebron, in monte Iudae et suburbana eius per circuitum.
JOSH|21|12|Agros vero et villas eius dederant Chaleb filio Iephonne ad possidendum.
JOSH|21|13|Dederunt ergo filiis Aaron sacerdotis Hebron confugii civitatem ac suburbana eius et Lobnam cum suburbanis suis
JOSH|21|14|et Iether et Esthemo
JOSH|21|15|et Helon et Dabir
JOSH|21|16|et Ain et Iutta et Bethsames cum suburbanis suis: civitates novem de tribubus illis duabus.
JOSH|21|17|De tribu autem Beniamin Gabaon et Gabaa
JOSH|21|18|et Anathoth et Almath cum suburbanis suis: civitates quattuor.
JOSH|21|19|Omnes simul civitates filiorum Aaron sacerdotis tredecim cum suburbanis suis.
JOSH|21|20|Reliquis vero ex familiis filiorum Caath Levitis haec est data possessio:
JOSH|21|21|de tribu Ephraim urbs confugii Sichem cum suburbanis suis in monte Ephraim et Gazer
JOSH|21|22|et Cibsaim et Bethoron cum suburbanis suis: civitates quattuor.
JOSH|21|23|De tribu quoque Dan Elthece et Gebbethon
JOSH|21|24|et Aialon et Gethremmon cum suburbanis suis: civitates quattuor.
JOSH|21|25|Porro de dimidia tribu Manasse Thanach et Gethremmon cum suburbanis suis: civitates duae.
JOSH|21|26|Omnes civitates decem et suburbana earum datae sunt filiis Caath inferioris gradus.
JOSH|21|27|Filiis quoque Gerson levitici generis dederunt de dimidia tribu Manasse confugii civitatem Golan in Basan et Astharoth cum suburbanis suis: civitates duas.
JOSH|21|28|Porro de tribu Issachar Cesion et Dabereth
JOSH|21|29|et Iaramoth et Engannim cum suburbanis suis: civitates quattuor.
JOSH|21|30|De tribu autem Aser Masal et Abdon
JOSH|21|31|et Helcath et Rohob cum suburbanis suis: civitates quattuor.
JOSH|21|32|De tribu quoque Nephthali civitas confugii Cedes in Galilaea et Ammothdor et Carthan cum suburbanis suis: civitates tres.
JOSH|21|33|Omnes urbes familiarum Gerson tredecim cum suburbanis suis.
JOSH|21|34|Filiis autem Merari Levitis inferioris gradus per familias suas data est de tribu Zabulon Iecnaam et Cartha
JOSH|21|35|et Remmon et Naalol: civitates quattuor cum suburbanis suis.
JOSH|21|36|De tribu Ruben ultra Iordanem contra Iericho civitas refugii Bosor in solitudine planitiei et Iasa
JOSH|21|37|et Cademoth et Mephaath: civitates quattuor cum suburbanis suis.
JOSH|21|38|Et de tribu Gad civitas confugii Ramoth in Galaad et Mahanaim
JOSH|21|39|et Hesebon et Iazer: civitates quattuor cum suburbanis suis.
JOSH|21|40|Omnes urbes filiorum Merari per familias reliquas de cognationibus Levitarum duodecim.
JOSH|21|41|Itaque universae civitates Levitarum in medio possessionis filiorum Israel fuerunt quadraginta octo
JOSH|21|42|cum suburbanis suis, singulae cum suburbanis suis in circuitu.
JOSH|21|43|Deditque Dominus Israeli omnem terram, quam traditurum se patribus eorum iuraverat, et possederunt illam atque habitaverunt in ea.
JOSH|21|44|Deditque Dominus eis requiem secundum omnia, quae iuraverat patribus eorum, nullusque eis hostium resistere ausus est, sed cunctos in eorum dicionem redegit.
JOSH|21|45|Ne unum quidem verbum bonum, quod locutus est ad domum Israel, irritum fuit, sed rebus expleta sunt omnia.
JOSH|22|1|Tunc vocavit Iosue Rubenitas et Gaditas et dimidiam tribum Manasse
JOSH|22|2|dixitque ad eos: "Fecistis omnia, quae vobis praecepit Moyses famulus Domini; mihi quoque in omnibus, quae praecepi vobis, oboedistis
JOSH|22|3|nec reliquistis fratres vestros hoc longo tempore usque in praesentem diem custodientes imperium Domini Dei vestri.
JOSH|22|4|Quia igitur dedit Dominus Deus vester fratribus vestris quietem ac pacem, sicut eis pollicitus est, revertimini nunc et ite in tabernacula vestra et in terram possessionis, quam tradidit vobis Moyses famulus Domini trans Iordanem;
JOSH|22|5|ita dumtaxat ut custodiatis attente et opere compleatis mandatum et legem, quam praecepit vobis Moyses servus Domini, ut diligatis Dominum Deum vestrum et ambuletis in omnibus viis eius et observetis mandata illius adhaereatisque ei ac serviatis in omni corde et in omni anima vestra ".
JOSH|22|6|Benedixitque eis Iosue et dimisit eos, qui reversi sunt in tabernacula sua.
JOSH|22|7|Dimidiae autem tribui Manasse possessionem Moyses dederat in Basan; et idcirco mediae, quae superfuit, dedit Iosue sortem inter ceteros fratres suos trans Iordanem ad occidentalem eius plagam. Cumque dimitteret eos in tabernacula sua et benedixisset illis,
JOSH|22|8|dixit ad eos: "Cum multis divitiis revertimini ad sedes vestras, cum argento et auro, aere ac ferro et veste multiplici; dividite praedam hostium cum fratribus vestris ".
JOSH|22|9|Reversique sunt et abierunt filii Ruben et filii Gad et dimidia tribus Manasse a filiis Israel de Silo, quae sita est in Chanaan, ut intrarent Galaad terram possessionis suae, quam obtinuerant iuxta imperium Domini in manu Moysi.
JOSH|22|10|Cumque venissent ad circulos Iordanis in terra Chanaan, aedificaverunt iuxta Iordanem altare ingens aspectu.
JOSH|22|11|Cum audissent filii Israel aedificasse filios Ruben et Gad et dimidiam tribum Manasse altare e regione terrae Chanaan ad Iordanis circulos ex adverso filiorum Israel,
JOSH|22|12|convenerunt omnes in Silo, ut ascenderent et dimicarent contra eos.
JOSH|22|13|Et interim miserunt ad illos in terram Galaad Phinees filium Eleazari sacerdotem
JOSH|22|14|et decem principes cum eo, singulos de tribubus, unusquisque erat caput familiae in cognationibus Israel.
JOSH|22|15|Qui venerunt ad filios Ruben et Gad et dimidiam tribum Manasse in terram Galaad dixeruntque ad eos:
JOSH|22|16|" Haec mandat omnis coetus Domini: Quae est ista transgressio? Cur reliquistis Dominum, Deum Israel, aedificantes vobis altare sacrilegum et a cultu illius recedentes?
JOSH|22|17|An parum vobis est peccatum Phegor, et usque in praesentem diem macula huius sceleris in nobis permanet, et facta est plaga in coetu Domini?
JOSH|22|18|Et vos hodie reliquistis Dominum, et factum est ut rebellaretis contra Dominum; et cras in universum coetum Israel eius ira desaeviet.
JOSH|22|19|Quod si putatis immundam esse terram possessionis vestrae, transite ad terram possessionis Domini, in qua habitaculum Domini est, et habitate inter nos; tantum ut contra Dominum non rebelletis nec nos rebellare faciatis aedificantes altare praeter altare Domini Dei nostri.
JOSH|22|20|Nonne Achan filius Zarae praeteriit mandatum Domini de anathemate, et super omnem coetum Israel ira Domini incubuit? Et ille erat unus homo; atque utinam solus perisset in scelere suo! ".
JOSH|22|21|Responderuntque filii Ruben et Gad et dimidia tribus Manasse principibus legationis Israel:
JOSH|22|22|" Fortissimus Deus Dominus, fortissimus Deus Dominus ipse novit, et Israel simul intelleget: si rebellionis, si praevaricationis animo contra Dominum hoc altare construximus, non salvet nos, sed puniat in praesenti;
JOSH|22|23|et si ea mente fecimus, ut recedamus a Domino et holocausta et oblationes et pacificas victimas super eo imponeremus, Dominus ipse quaerat et iudicet;
JOSH|22|24|et si non ea magis sollicitudine et cogitatione fecimus hoc dicentes: Cras dicent filii vestri filiis nostris: "Quid vobis et Domino, Deo Israel?
JOSH|22|25|Terminum posuit Dominus inter nos et vos, o filii Ruben et filii Gad, Iordanem fluvium, et idcirco partem non habetis in Domino"; et per hanc occasionem avertent filii vestri filios nostros a timore Domini. Putavimus itaque melius
JOSH|22|26|et diximus: Exstruamus nobis altare non in holocausta neque ad victimas offerendas,
JOSH|22|27|sed in testimonium inter nos et vos et sobolem nostram vestramque progeniem, ut serviamus Domino, et iuris nostri sit offerre holocausta et victimas et pacificas hostias, et nequaquam dicant cras filii vestri filiis nostris: "Non est vobis pars in Domino".
JOSH|22|28|Quod si voluerint dicere, respondebunt eis: "Ecce similitudo altaris Domini, quam fecerunt patres nostri non in holocausta neque in sacrificia, sed in testimonium inter nos et vos".
JOSH|22|29|Absit a nobis hoc scelus, ut recedamus a Domino et eius vestigia relinquamus, exstructo altari ad holocausta et oblationes et victimas offerendas, praeter altare Domini Dei nostri, quod est ante habitaculum eius ".
JOSH|22|30|Quibus auditis, Phinees sacerdos et principes legationis Israel, qui erant cum eo, placati sunt et verba filiorum Ruben et Gad et dimidiae tribus Manasse libentissime susceperunt;
JOSH|22|31|dixitque Phinees filius Eleazar sacerdos ad eos: " Nunc scimus quod nobiscum sit Dominus, quoniam alieni estis a praevaricatione hac et liberastis filios Israel de manu Domini ".
JOSH|22|32|Reversusque est cum principibus a filiis Ruben et Gad de terra Galaad in terram Chanaan ad filios Israel et rettulit eis.
JOSH|22|33|Placuitque sermo cunctis audientibus, et laudaverunt Deum filii Israel; et nequaquam ultra dixerunt, ut ascenderent contra eos in bellum et delerent terram, in qua habitabant filii Ruben et Gad.
JOSH|22|34|Vocaveruntque filii Ruben et filii Gad altare, quod exstruxerant, Testem; dixerunt enim: " Testis est inter nos quod Dominus ipse sit Deus.
JOSH|23|1|Evoluto autem multo tem pore, postquam pacem Do minus dederat Israeli ab omnibus in gyro nationibus et Iosue iam longaevo et persenilis aetatis,
JOSH|23|2|vocavit Iosue omnem Israelem maioresque natu et principes ac iudices et praefectos dixitque ad eos: " Ego senui et progressioris aetatis sum,
JOSH|23|3|vosque vidistis omnia, quae fecerit Dominus Deus vester cunctis nationibus istis, quomodo pro vobis ipse pugnaverit.
JOSH|23|4|Videte, sorte divisi vobis gentes, quae supersunt, in possessionem tribuum vestrarum, sicut omnes, quas delevi, a Iordane usque ad mare Magnum in occidente.
JOSH|23|5|Dominus Deus vester disperdet eas et auferet a facie vestra, et possidebitis terram eorum, sicut vobis pollicitus est.
JOSH|23|6|Tantum confortamini, ut custodiatis cuncta, quae scripta sunt in volumine legis Moysi, et non declinetis ab eis nec ad dexteram nec ad sinistram;
JOSH|23|7|ne conveniatis cum gentibus, quae inter vos residuae sunt, et iuretis in nomine deorum earum et serviatis eis et adoretis illos;
JOSH|23|8|sed adhaereatis Domino Deo vestro, quod fecistis usque in diem hanc.
JOSH|23|9|Et expulit Dominus in conspectu vestro gentes magnas et robustissimas, et nullus vobis resistere potuit:
JOSH|23|10|unus e vobis persequitur hostium mille viros, quia Dominus Deus vester pro vobis ipse pugnat, sicut pollicitus est;
JOSH|23|11|hoc tantum diligentissime praecavete, ut diligatis Dominum Deum vestrum.
JOSH|23|12|Quod si volueritis gentium harum, quae inter vos residuae sunt, erroribus adhaerere et cum eis miscere conubia atque amicitias copulare,
JOSH|23|13|iam nunc scitote quod Dominus Deus vester non eas deleat ante faciem vestram; sed sint vobis in rete, foveam ac laqueum et flagellum ex latere vestro, et spinae in oculis vestris, donec vos disperdat de terra hac optima, quam tradidit vobis.
JOSH|23|14|En ego hodie ingredior viam universae terrae; et toto animo cognoscetis quod de omnibus verbis bonis, quae Dominus Deus vester locutus est vobis, non praeterierit ne unum quidem incassum.
JOSH|23|15|Sicut ergo implevit opere, quod promisit, et prospera cuncta venerunt, sic adducet super vos quidquid malorum comminatus est, donec vos disperdat de terra hac optima, quam tradidit vobis.
JOSH|23|16|Si praeterieritis pactum Domini Dei vestri, quod mandavit vobis, et servieritis diis alienis et adoraveritis eos, consurget in vos furor Domini, et cito peribitis ab hac terra optima, quam tradidit vobis ".
JOSH|24|1|Congregavitque Iosue omnes tribus Israel in Sichem et vocavit maiores natu ac principes et iudices et praefectos, steteruntque in conspectu Dei;
JOSH|24|2|et ad totum populum sic locutus est: " Haec dicit Dominus, Deus Israel: Trans fluvium habitaverunt patres vestri ab initio, Thare pater Abraham et Nachor, servieruntque diis alienis.
JOSH|24|3|Tuli ergo patrem vestrum Abraham de Mesopotamiae finibus et adduxi eum per totam terram Chanaan multiplicavique semen eius.
JOSH|24|4|Et dedi ei Isaac illique rursum dedi Iacob et Esau; e quibus Esau dedi montem Seir ad possidendum, Iacob vero et filii eius descenderunt in Aegyptum.
JOSH|24|5|Misique Moysen et Aaron et percussi Aegyptum signis, quae feci in medio eius, et postea eduxi vos.
JOSH|24|6|Eduxique patres vestros de Aegypto, et venistis ad mare. Persecutique sunt Aegyptii patres vestros cum curribus et equitatu usque ad mare Rubrum.
JOSH|24|7|Clamaverunt autem ad Dominum, qui posuit tenebras inter vos et Aegyptios et adduxit super eos mare et operuit illos. Viderunt oculi vestri, quae in Aegypto fecerim; et habitastis in solitudine multo tempore.
JOSH|24|8|Et introduxi vos ad terram Amorraei, qui habitabat trans Iordanem; cumque pugnarent contra vos, tradidi eos in manus vestras, et occupastis terram eorum atque interfecistis illos.
JOSH|24|9|Surrexit autem Balac filius Sephor rex Moab et pugnavit contra Israelem; misitque et vocavit Balaam filium Beor, ut malediceret vobis.
JOSH|24|10|Et ego nolui audire eum, sed e contrario benedixit vobis, et liberavi vos de manu eius.
JOSH|24|11|Transistisque Iordanem et venistis ad Iericho; pugnaveruntque contra vos viri civitatis illius, Amorraeus et Pherezaeus et Chananaeus et Hetthaeus et Gergesaeus et Hevaeus et Iebusaeus; et tradidi illos in manus vestras.
JOSH|24|12|Misique ante vos crabrones, et eiecerunt eos coram vobis - duos reges Amorraeorum - non in gladio nec in arcu tuo.
JOSH|24|13|Dedique vobis terram, de qua non laborastis, et urbes, quas non aedificastis, et habitatis in eis, vineas et oliveta, quae non plantastis, et manducatis ex eis.
JOSH|24|14|Nunc ergo timete Dominum et servite ei perfecto corde atque verissimo; et auferte deos, quibus servierunt patres vestri in Mesopotamia et in Aegypto, ac servite Domino.
JOSH|24|15|Sin autem malum vobis videtur, ut Domino serviatis, eligite vobis hodie, cui servire vultis, utrum diis, quibus servierunt patres vestri in Mesopotamia, an diis Amorraeorum, in quorum terra habitatis. Ego autem et domus mea serviemus Domino ".
JOSH|24|16|Responditque populus et ait: " Absit a nobis, ut relinquamus Dominum et serviamus diis alienis.
JOSH|24|17|Dominus Deus noster ipse eduxit nos et patres nostros de terra Aegypti, de domo servitutis; fecitque videntibus nobis signa ingentia et custodivit nos in omni via, per quam ambulavimus, et in cunctis populis, per quos transivimus;
JOSH|24|18|et eiecit universas gentes, Amorraeum habitatorem terrae, quam nos intravimus. Serviemus igitur etiam nos Domino, quia ipse est Deus noster.
JOSH|24|19|Dixitque Iosue ad populum: " Non poteritis servire Domino. Deus enim sanctus et Deus aemulator est nec ignoscet sceleribus vestris atque peccatis.
JOSH|24|20|Si dimiseritis Dominum et servieritis diis alienis, convertet se et affliget vos atque subvertet, postquam vobis praestiterit bona ".
JOSH|24|21|Dixitque populus ad Iosue: " Nequaquam, sed Domino serviemus ".
JOSH|24|22|Et Iosue ad populum: " Testes, inquit, vos estis contra vos quia ipsi elegeritis vobis Dominum, ut serviatis ei ". Responderuntque: " Testes ".
JOSH|24|23|" Nunc ergo, ait, auferte deos alienos de medio vestri et inclinate corda vestra ad Dominum, Deum Israel".
JOSH|24|24|Dixitque populus ad Iosue: "Domino Deo nostro serviemus; oboedientes erimus praeceptis eius ".
JOSH|24|25|Percussit igitur Iosue in die illo foedus populo et proposuit ei praecepta atque iudicia in Sichem.
JOSH|24|26|Scripsitque verba haec in volumine legis Dei; et tulit lapidem pergrandem posuitque eum ibi subter quercum, quae erat in sanctuario Domini,
JOSH|24|27|et dixit ad omnem populum: " En lapis iste erit adversus vos in testimonium quia audivit omnia verba Domini, quae locutus est inter nos, ne forte postea negare velitis et mentiri Domino Deo vestro ".
JOSH|24|28|Dimisitque populum, singulos in possessionem suam.
JOSH|24|29|Et post haec mortuus est Iosue filius Nun, servus Domini, centum decem annorum.
JOSH|24|30|Sepelieruntque eum in finibus possessionis suae in Thamnathsare, quae sita est in monte Ephraim a septentrionali parte montis Gaas.
JOSH|24|31|Servivitque Israel Domino cunctis diebus Iosue et seniorum, qui longo vixerunt tempore post Iosue et qui noverunt omnia opera Domini, quae fecerat Israel.
JOSH|24|32|Ossa quoque Ioseph, quae tulerant filii Israel de Aegypto, sepelierunt in Sichem, in parte agri, quem emerat Iacob a filiis Hemmor patris Sichem centum argenteis, et fuit in possessionem filiorum Ioseph.
JOSH|24|33|Eleazar quoque filius Aaron mortuus est; et sepelierunt eum in Gabaa Phinees filii eius, quae data est ei in monte Ephraim.
JUDG|1|1|Post mortem Iosue consulue runt filii Israel Dominum dicen tes: " Quis nostrum primus ascendet ad Chananaeum ad pugnandum contra eum? ".
JUDG|1|2|Dixitque Dominus: " Iudas ascendet: ecce tradidi terram in manus eius ".
JUDG|1|3|Et ait Iudas Simeoni fratri suo: " Ascende mecum in sorte mea, et pugnemus contra Chananaeum, et ego pergam tecum in sorte tua ". Et abiit cum eo Simeon.
JUDG|1|4|Ascenditque Iudas, et tradidit Dominus Chananaeum ac Pherezaeum in manus eorum, et percusserunt in Bezec decem milia virorum.
JUDG|1|5|Inveneruntque Adonibezec in Bezec et pugnaverunt contra eum ac percusserunt Chananaeum et Pherezaeum.
JUDG|1|6|Fugit autem Adonibezec, quem persecuti comprehenderunt, caesis pollicibus manuum eius ac pedum.
JUDG|1|7|Dixitque Adonibezec: " Septuaginta reges, amputatis manuum ac pedum pollicibus, colligebant sub mensa mea ciborum reliquias. Sicut feci, ita reddidit mihi Deus ". Adduxeruntque eum in Ierusalem, et ibi mortuus est.
JUDG|1|8|Oppugnantes ergo filii Iudae Ierusalem ceperunt eam; et percusserunt in ore gladii tradentes incendio civitatem.
JUDG|1|9|Et postea descendentes pugnaverunt contra Chananaeum, qui habitabat in montanis et in Nageb et in Sephela.
JUDG|1|10|Pergensque Iuda contra Chananaeum, qui habitabat in Hebron, cui nomen fuit antiquitus Cariatharbe, percussit Sesai et Ahiman et Tholmai.
JUDG|1|11|Atque inde profectus abiit ad habitatores Dabir, cuius nomen vetus erat Cariathsepher (id est civitas Litterarum).
JUDG|1|12|Dixitque Chaleb: " Qui percusserit Cariathsepher et ceperit eam, dabo ei Axam filiam meam uxorem ".
JUDG|1|13|Cumque cepisset eam Othoniel filius Cenez frater Chaleb minor, dedit ei Axam filiam suam coniugem.
JUDG|1|14|Quae cum veniret, incitavit eum, ut peteret a patre suo agrum. Demisit ergo se de asino, et dixit ei Chaleb: " Quid habes? ".
JUDG|1|15|At illa respondit: " Da mihi benedictionem; quia terram arentem dedisti mihi, da et irriguam aquis ". Dedit ergo ei Chaleb irriguum superius et irriguum inferius.
JUDG|1|16|Filii autem Hobab Cinaei cognati Moysi ascenderunt de civitate Palmarum cum filiis Iudae in desertum Iudae, quod est ad meridiem Arad, et habitaverunt cum Amalecitis.
JUDG|1|17|Abiit autem Iudas cum Simeone fratre suo et percusserunt simul Chananaeum, qui habitabat in Sephath, et percusserunt urbem anathemate. Vocatumque est nomen eius Horma (id est Anathema).
JUDG|1|18|Cepitque Iudas Gazam cum finibus suis et Ascalonem atque Accaron cum terminis suis.
JUDG|1|19|Fuitque Dominus cum Iuda, et montana possedit; nec potuit expellere habitatores vallis, quia falcatis curribus abundabant.
JUDG|1|20|Dederuntque Chaleb Hebron, sicut dixerat Moyses, qui expulit ex ea tres filios Enac.
JUDG|1|21|Iebusaeum autem habitatorem Ierusalem non expulerunt filii Beniamin, habitavitque Iebusaeus cum filiis Beniamin in Ierusalem usque in praesentem diem.
JUDG|1|22|Domus quoque Ioseph ascendit Bethel, fuitque Dominus cum eis.
JUDG|1|23|Nam, cum explorarent urbem, quae prius Luza vocabatur,
JUDG|1|24|viderunt custodes hominem egredientem de civitate dixeruntque ad eum: " Ostende nobis introitum civitatis, et faciemus tecum misericordiam ".
JUDG|1|25|Qui cum ostendisset eis, percusserunt urbem in ore gladii; hominem autem illum et omnem cognationem eius dimiserunt.
JUDG|1|26|Qui dimissus abiit in terram Hetthim et aedificavit ibi civitatem vocavitque eam Luzam, quae ita appellatur usque in praesentem diem.
JUDG|1|27|Manasses quoque non occupavit Bethsan et Thanach cum viculis suis nec expulit habitatores Dor et Ieblaam et Mageddo cum viculis suis; mansitque Chananaeus in terra hac.
JUDG|1|28|Postquam autem confortatus est Israel, fecit eos tributarios et expellere noluit.
JUDG|1|29|Ephraim etiam non expulit Chananaeum, qui habitabat in Gazer, sed habitavit Chananaeus in medio eius in Gazer.
JUDG|1|30|Zabulon non expulit habitatores Cetron et Naalol, sed habitavit Chananaeus in medio eius factusque est ei tributarius.
JUDG|1|31|Aser quoque non expulit habitatores Achcho et Sidonis, Ahalab et Achazib et Helba et Aphec et Rohob;
JUDG|1|32|habitavitque Aser in medio Chananaei habitatoris illius terrae, quia non expulit eum.
JUDG|1|33|Nephthali non expulit habitatores Bethsames et Bethanath et habitavit inter Chananaeum habitatorem terrae, fueruntque ei Bethsamitae et Bethanitae tributarii.
JUDG|1|34|Artavitque Amorraeus filios Dan in montem nec dedit eis locum, ut ad planiora descenderent.
JUDG|1|35|Habitavitque Amorraeus in Hathares, in Aialon et Salebim; et aggravata est manus domus Ioseph, factusque est ei tributarius.
JUDG|1|36|Fuit autem terminus Amorraei ab ascensu Acrabbim ad Petram et superiora loca.
JUDG|2|1|Ascenditque angelus Domini de Galgalis in Bochim et ait: " Eduxi vos de Aegypto et introduxi in terram, pro qua iuravi patribus vestris et pollicitus sum, ut non facerem irritum pactum meum vobiscum in sempiternum,
JUDG|2|2|ita dumtaxat ut non feriretis foedus cum habitatoribus terrae huius, sed aras eorum subverteretis. Et noluistis audire vocem meam. Cur hoc fecistis?
JUDG|2|3|Quam ob rem nolui expellere eos a facie vestra, ut sint vobis in laqueum, et dii eorum in ruinam ".
JUDG|2|4|Cumque loqueretur angelus Domini verba haec ad omnes filios Israel, elevaverunt vocem suam et fleverunt.
JUDG|2|5|Et vocatum est nomen loci illius Bochim (id est locus Flentium); immolaveruntque ibi hostias Domino.
JUDG|2|6|Dimisit ergo Iosue populum, et abierunt filii Israel unusquisque in possessionem suam, ut obtinerent terram.
JUDG|2|7|Servieruntque Domino cunctis diebus Iosue et seniorum, qui longo post eum vixerunt tempore et viderant universum opus magnum Domini, quod fecerat cum Israel.
JUDG|2|8|Mortuus est autem Iosue filius Nun famulus Domini centum et decem annorum;
JUDG|2|9|et sepelierunt eum in finibus possessionis suae in Thamnathsare in monte Ephraim a septentrionali plaga montis Gaas.
JUDG|2|10|Omnisque illa generatio congregata est ad patres suos, et surrexerunt alii post illam, qui non noverant Dominum et opus, quod fecerat cum Israel.
JUDG|2|11|Feceruntque filii Israel malum in conspectu Domini et servierunt Baalim
JUDG|2|12|ac dimiserunt Dominum, Deum patrum suorum, qui eduxerat eos de terra Aegypti, et secuti sunt deos alienos, de diis populorum, qui habitabant in circuitu eorum, et adoraverunt eos et ad iracundiam concitaverunt Dominum
JUDG|2|13|dimittentes eum et servientes Baal et Astharoth.
JUDG|2|14|Iratusque Dominus contra Israel tradidit eos in manibus diripientium, qui diripuerunt eos, et vendidit eos hostibus, qui habitabant per gyrum, nec potuerunt resistere adversariis suis;
JUDG|2|15|sed, quocumque pergere voluissent, manus Domini erat super eos ad malum, sicut locutus est et iuravit eis, et vehementer afflicti sunt.
JUDG|2|16|Suscitavitque Dominus iudices, qui liberarent eos de vastantium manibus;
JUDG|2|17|sed nec illos audire voluerunt fornicantes cum diis alienis et adorantes eos. Cito deseruerunt viam, per quam ingressi fuerant patres eorum audientes mandata Domini, et omnia fecere contraria.
JUDG|2|18|Cumque Dominus iudices suscitaret eis, erat Dominus cum iudice et liberabat eos de manu hostium eorum toto tempore iudicis, quia flectebatur misericordia et audiebat gemitus afflictorum.
JUDG|2|19|Postquam autem mortuus esset iudex, revertebantur et multo faciebant peiora quam fecerant patres sui, sequentes deos alienos, servientes eis et adorantes illos: non dimiserunt opera sua et viam durissimam, per quam ambulare consueverant.
JUDG|2|20|Iratusque est furor Domini in Israel et ait: " Quia irritum fecit gens ista pactum meum, quod pepigeram cum patribus eorum, et vocem meam audire contempsit,
JUDG|2|21|et ego non expellam gentes, quas dimisit Iosue et mortuus est;
JUDG|2|22|ut in ipsis experiar Israel, utrum custodiant viam Domini et ambulent in ea, sicut custodierunt patres eorum, an non ".
JUDG|2|23|Dimisit ergo Dominus has nationes et cito expellere noluit nec tradidit in manibus Iosue.
JUDG|3|1|Hae sunt gentes, quas Dominus dereliquit, ut erudiret in eis Is raelem, omnes, qui non noverant bella Chananaeorum,
JUDG|3|2|ut discerent certare cum hostibus generationes filiorum Israel, quae non habebant consuetudinem proeliandi:
JUDG|3|3|quinque satrapae Philisthinorum omnisque Chananaeus et Sidonius atque Hevaeus, qui habitabat in monte Libano de monte Baalhermon usque ad introitum Emath.
JUDG|3|4|Dimisitque eos, ut in ipsis experiretur Israelem, utrum audiret mandata Domini, quae praeceperat patribus eorum per manum Moysi, an non.
JUDG|3|5|Itaque filii Israel habitaverunt in medio Chananaei et Hetthaei et Amorraei et Pherezaei et Hevaei et Iebusaei
JUDG|3|6|et duxerunt uxores filias eorum, ipsique filias suas eorum filiis tradiderunt, et servierunt diis eorum.
JUDG|3|7|Feceruntque filii Israel malum in conspectu Domini et obliti sunt Domini Dei sui servientes Baalim et Astharoth.
JUDG|3|8|Iratusque Dominus contra Israel tradidit eos in manus Chusanrasathaim regis Mesopotamiae, servieruntque ei octo annis.
JUDG|3|9|Et clamaverunt ad Dominum, qui suscitavit eis salvatorem et liberavit eos, Othoniel videlicet filium Cenez fratrem Chaleb minorem.
JUDG|3|10|Fuitque in eo spiritus Domini, et iudicavit Israelem egressusque est ad pugnam; et tradidit Dominus in manu eius Chusanrasathaim regem Mesopotamiae, et praevaluit adversus eum.
JUDG|3|11|Quievitque terra quadraginta annis, et mortuus est Othoniel filius Cenez.
JUDG|3|12|Addiderunt autem filii Israel facere malum in conspectu Domini, qui confortavit adversum eos Eglon regem Moab, quia fecerunt malum in conspectu Domini.
JUDG|3|13|Et copulavit sibi Eglon filios Ammon et Amalec abiitque et percussit Israel atque possedit urbem Palmarum.
JUDG|3|14|Servieruntque filii Israel Eglon regi Moab decem et octo annis.
JUDG|3|15|Et clamaverunt filii Israel ad Dominum, qui suscitavit eis salvatorem Aod filium Gera de Beniamin, qui sinistra manu utebatur pro dextera. Miseruntque filii Israel per illum munera Eglon regi Moab.
JUDG|3|16|Fecitque Aod sibi gladium ancipitem longitudinis palmae manus et accinctus est eo subter vestem in dextro femore
JUDG|3|17|obtulitque munera Eglon regi Moab. Erat autem Eglon crassus nimis.
JUDG|3|18|Cumque obtulisset ei munera, dimisit socios, qui illa portaverant;
JUDG|3|19|et reversus de Galgalis, ubi erant idola, dixit ad regem: " Verbum secretum habeo ad te, o rex ". Et ille imperavit silentium; egressique sunt omnes, qui circa eum erant.
JUDG|3|20|Aod autem ingressus erat ad eum, cum sederet in aestivo cenaculo, quod ipsi soli erat, dixitque: " Verbum Dei habeo ad te ". Qui statim surrexit de throno.
JUDG|3|21|Extenditque Aod manum sinistram et tulit sicam de dextro femore suo infixitque eam in ventre eius
JUDG|3|22|tam valide, ut capulus ferrum sequeretur in vulnere ac pinguissimo adipe stringeretur. Nec eduxit gladium, sed ita, ut percusserat, reliquit in corpore; statimque per secreta naturae alvi stercora proruperunt.
JUDG|3|23|Aod autem egressus in atrium clausit ostium cenaculi post se et obfirmavit sera.
JUDG|3|24|Egresso illo, servi regis venerunt et, cum viderent clausas fores cenaculi, dixerunt: " Certe purgat alvum in aestivo cubiculo ".
JUDG|3|25|Exspectantesque diu, donec erubescerent, et videntes quod nullus aperiret, tulerunt clavem et aperientes invenerunt dominum suum iacentem in terra mortuum.
JUDG|3|26|Aod autem, dum illi cunctarentur, effugerat et pertransiit locum idolorum, unde reversus fuerat, venitque in Seira.
JUDG|3|27|Et statim insonuit bucina in monte Ephraim; descenderuntque cum eo filii Israel, ipso in fronte gradiente.
JUDG|3|28|Qui dixit ad eos: " Sequimini me; tradidit enim Dominus inimicos vestros Moabitas in manus vestras ". Descenderuntque post eum et occupaverunt vada Iordanis, quae transmittunt in Moab, et non dimiserunt transire quemquam,
JUDG|3|29|sed percusserunt Moabitas in tempore illo circiter decem milia, omnes robustos et fortes viros. Nullus eorum evadere potuit.
JUDG|3|30|Humiliatusque est Moab die illo sub manu Israel; et quievit terra octoginta annis.
JUDG|3|31|Post hunc fuit Samgar filius Anath, qui percussit de Philisthim sescentos viros stimulo boum; et ipse quoque salvum fecit Israel.
JUDG|4|1|Addideruntque filii Israel facere malum in conspectu Domini post mortem Aod,
JUDG|4|2|et tradidit illos Dominus in manu Iabin regis Chanaan, qui regnavit in Asor. Habuitque ducem exercitus sui nomine Sisaram: ipse autem habitabat in Haroseth gentium.
JUDG|4|3|Clamaveruntque filii Israel ad Dominum; nongentos enim habebat falcatos currus et per viginti annos vehementer oppresserat eos.
JUDG|4|4|Erat autem Debora prophetis, uxor Lapidoth, quae iudicabat Israel in illo tempore.
JUDG|4|5|Et sedebat sub palma Deborae inter Rama et Bethel in monte Ephraim; ascendebantque ad eam filii Israel in iudicium.
JUDG|4|6|Quae misit et vocavit Barac filium Abinoem de Cedes Nephthali dixitque ad eum: " Praecepit tibi Dominus, Deus Israel: Vade et duc exercitum in montem Thabor tollesque tecum decem milia pugnatorum de filiis Nephthali et de filiis Zabulon.
JUDG|4|7|Ego autem ducam ad te in loco torrentis Cison Sisaram principem exercitus Iabin et currus eius atque omnem multitudinem et tradam eum in manu tua ".
JUDG|4|8|Dixitque ad eam Barac: " Si venis mecum, vadam; si nolueris venire mecum, non pergam ".
JUDG|4|9|Quae dixit ad eum: " Ibo quidem tecum; sed in hac via non erit tibi gloria, quia in manu mulieris tradet Dominus Sisaram ".Surrexit itaque Debora et perrexit cum Barac in Cedes.
JUDG|4|10|Qui, accitis Zabulon et Nephthali in Cedes, ascendit cum decem milibus pugnatorum habens Deboram in comitatu suo.
JUDG|4|11|Haber autem Cinaeus recesserat a ceteris Cinaeis fratribus suis filiis Hobab cognati Moysi et tetendit tabernaculum usque ad quercum in Saananim iuxta Cedes.
JUDG|4|12|Nuntiatumque est Sisarae quod ascendisset Barac filius Abinoem in montem Thabor,
JUDG|4|13|et congregavit omnes nongentos falcatos currus omnemque exercitum, qui cum eo erat, de Haroseth gentium ad torrentem Cison.
JUDG|4|14|Dixitque Debora ad Barac: " Surge: haec est enim dies, in qua tradidit Dominus Sisaram in manus tuas. En ipse ductor est tuus ". Descendit itaque Barac de monte Thabor, et decem milia pugnatorum cum eo.
JUDG|4|15|Perterruitque Dominus Sisaram et omnes currus eius universamque multitudinem in ore gladii ad conspectum Barac, in tantum ut Sisara de curru desiliens pedibus fugeret,
JUDG|4|16|et Barac persequeretur fugientes currus et exercitum usque ad Haroseth gentium, et omnis hostium multitudo usque ad internecionem caderet.
JUDG|4|17|Sisara autem fugiens pervenit ad tentorium Iahel uxoris Haber Cinaei; erat enim pax inter Iabin regem Asor et domum Haber Cinaei.
JUDG|4|18|Egressa igitur Iahel in occursum Sisarae dixit ad eum: " Intra ad me, domine mi; intra, ne timeas ". Qui ingressus tabernaculum eius et opertus ab ea panno,
JUDG|4|19|dixit ad eam: " Da mihi, obsecro, paululum aquae, quia sitio ". Quae aperuit utrem lactis et dedit ei bibere et operuit illum.
JUDG|4|20|Dixitque Sisara ad eam: " Sta ante ostium tabernaculi et, cum venerit aliquis interrogans te et dicens: "Numquid hic est aliquis?", respondebis: Nullus est" ".
JUDG|4|21|Tulit porro Iahel uxor Haber clavum tabernaculi assumens pariter malleum; et ingressa abscondite et cum silentio, posuit supra tempus capitis eius clavum, percussumque malleo defixit in cerebrum usque ad terram; qui soporem morti socians defecit et mortuus est.
JUDG|4|22|Et ecce Barac sequens Sisaram veniebat; egressaque Iahel in occursum eius dixit ei: " Veni, et ostendam tibi virum, quem quaeris ". Qui cum intrasset ad eam, vidit Sisaram iacentem mortuum et clavum infixum in tempore eius.
JUDG|4|23|Humiliavit ergo Deus in die illo Iabin regem Chanaan coram filiis Israel,
JUDG|4|24|qui crescebant cotidie et forti manu opprimebant Iabin regem Chanaan, donec delerent eum.
JUDG|5|1|Cecineruntque Debora et Barac filius Abinoem in die illo dicen tes:
JUDG|5|2|" Quia comae excussae sunt in Israel,cum sponte se obtulit populus,benedicite Domino!
JUDG|5|3|Audite, reges, percipite auribus, principes;ego sum, ego sum, quae Domino canam,psallam Domino, Deo Israel!
JUDG|5|4|Domine, cum exires de Seir,incederes de regione Edom,terra mota est, caelique stillaverunt, ac nubes stillaverunt aquis;
JUDG|5|5|montes fluxerunt a facie Domini Sinai,a facie Domini, Dei Israel.
JUDG|5|6|In diebus Samgar filii Anath,in diebus Iahel quieverunt semitae; et, qui ingrediebantur per eas,ambulaverunt per calles devios.
JUDG|5|7|Cessaverunt fortes in Israel et quieverunt,donec surgeres, Debora,surgeres mater in Israel.
JUDG|5|8|Elegerunt deos novos;tunc erat pugna in portis.Clipeus et hasta non apparueruntin quadraginta milibus Israel.
JUDG|5|9|Cor meum diligit principes Israel.Qui sponte obtulistis vos in populo, benedicite Domino!
JUDG|5|10|Qui ascenditis super nitentes asinaset sedetis super tapetiaet ambulatis in via, loquimini.
JUDG|5|11|Ad vocem eorum,qui distribuunt aquas ad canales,ibi narrant iustitias Domini,iustitias fortitudinis eius in Israel:tunc descendit populus Domini ad portas.
JUDG|5|12|Surge, surge, Debora;surge, surge et loquere canticum!Surge, Barac, et apprehende captivos tuos,fili Abinoem!
JUDG|5|13|Tunc descenderunt reliquiae ad inclitos,populus Domini descendit pro eo in fortibus.
JUDG|5|14|Ex Ephraim venerunt principes in vallempost te, Beniamin, in populis tuis.De Machir principes descenderunt, et de Zabulon, qui tenent sceptrum, praefecti.
JUDG|5|15|Duces Issachar fuere cum Debora;sic Barac in vallem missus cum peditibus suis.In pagis Ruben magna consilia cordis.
JUDG|5|16|Quare sedebas inter caulas,ut audires sibilos tibiae apud greges?Pagis Ruben magnae investigationes cordis.
JUDG|5|17|Galaad trans Iordanem quiescebat;et Dan cur peregrinus vacabat navibus?Aser habitabat in litore mariset in portibus morabatur.
JUDG|5|18|Zabulon vero obtulit animam suam morti,et Nephthali super excelsa regionis.
JUDG|5|19|Venerunt reges et pugnaverunt,pugnaverunt reges Chanaanin Thanach iuxta aquas Mageddo, praedam argenti non tulere!
JUDG|5|20|De caelo dimicaverunt stellae,cursu suo adversus Sisaram pugnaverunt.
JUDG|5|21|Torrens Cison traxit cadavera eorum,torrens proeliorum, torrens Cison; incede, anima mea, fortiter.
JUDG|5|22|Tunc calcaverunt ungulae equorumin cursu praecipiti fortium suorum.
JUDG|5|23|Maledicite, Meroz, dixit angelus Domini,maledicite habitatoribus eius,quia non venerunt ad auxilium Domini,in adiutorium Domini in fortibus.
JUDG|5|24|Benedicta prae mulieribus Iahel uxor Haber Cinaei,prae mulieribus tabernaculi benedicatur!
JUDG|5|25|Aquam petenti lac deditet in phiala principum obtulit butyrum.
JUDG|5|26|Sinistram manum misit ad clavumet dextram ad fabrorum malleum:percussitque Sisaram quaerens in capite vulneri locumet tempus valide perforans.
JUDG|5|27|Inter pedes eius ruit, cecidit, iacebat;inter pedes eius ruit, cecidit;ubi ruit, ibi iacebat exanimis.
JUDG|5|28|Per fenestram prospiciens eiulabatmater Sisarae per cancellos:Cur moratur regredi currus eius? Quare tardant rotae quadrigarum illius?".
JUDG|5|29|Una sapientior ceteris uxoribus respondit ei,et ipsa sibi repetit verba illius:
JUDG|5|30|"Certo nunc dividunt inventa spolia, unam, duas feminas singulis viris;duas vestes diversorum colorumSisarae in praedam;unam, duas texturas discolorescollo meo in praedam".
JUDG|5|31|Sic pereant omnes inimici tui, Domine!Qui autem diligunt eum, rutilent,sicut sol in ortu suo splendet ".
JUDG|5|32|Quievitque terra per quadraginta annos.
JUDG|6|1|Fecerunt autem filii Israel malum in conspectu Domini, qui tradidit eos in manu Madian septem annis.
JUDG|6|2|Et oppressi sunt valde ab eis. Feceruntque sibi antra et speluncas in montibus et tutissima loca.
JUDG|6|3|Cumque sevisset Israel, ascendebat Madian et Amalec ceterique orientalium nationum
JUDG|6|4|et apud eos figentes tentoria, sicut erant in herbis, cuncta vastabant usque ad introitum Gazae nihilque omnino ad vitam pertinens relinquebant in Israel, non oves, non boves, non asinos.
JUDG|6|5|Ipsi enim et universi greges eorum veniebant cum tabernaculis suis et, instar locustarum, universa complebant, innumera multitudo hominum et camelorum, quidquid tetigerant devastantes.
JUDG|6|6|Humiliatusque est Israel valde in conspectu Madian.
JUDG|6|7|Et clamavit ad Dominum postulans auxilium contra Madianitas.
JUDG|6|8|Qui misit ad eos virum prophetam, et locutus est: " Haec dicit Dominus, Deus Israel: Ego vos feci conscendere de Aegypto et eduxi vos de domo servitutis
JUDG|6|9|et liberavi de manu Aegyptiorum et omnium inimicorum, qui affligebant vos, eiecique eos ad introitum vestrum et tradidi vobis terram eorum.
JUDG|6|10|Et dixi: Ego Dominus Deus vester, ne timeatis deos Amorraeorum, in quorum terra habitatis. Et noluistis audire vocem meam ".
JUDG|6|11|Venit autem angelus Domini et sedit sub quercu, quae erat in Ephra et pertinebat ad Ioas de familia Abiezer. Cumque Gedeon filius eius excuteret atque purgaret frumenta in torculari, ut absconderet a Madian,
JUDG|6|12|apparuit ei angelus Domini et ait: " Dominus tecum, vir fortis! ".
JUDG|6|13|Dixitque ei Gedeon: " Obsecro, domine mi, si Dominus nobiscum est, cur apprehenderunt nos haec omnia? Ubi sunt omnia mirabilia eius, quae narraverunt patres nostri atque dixerunt: "De Aegypto eduxit nos Dominus"? Nunc autem dereliquit nos Dominus et tradidit in manu Madian ".
JUDG|6|14|Respexitque ad eum Dominus et ait: " Vade in hac fortitudine tua et liberabis Israel de manu Madian; scito quod miserim te ".
JUDG|6|15|Qui respondens ait: " Obsecro, Domine, in quo liberabo Israel? Ecce familia mea infima est in Manasse, et ego minimus in domo patris mei ".
JUDG|6|16|Dixitque ei Dominus: " Ego ero tecum, et percuties Madian quasi unum virum ".
JUDG|6|17|Et ille: " Si inveni, inquit, gratiam coram te, da mihi signum quod tu sis, qui loquaris ad me;
JUDG|6|18|ne recedas hinc, donec revertar ad te portans oblationem et offerens tibi ". Qui respondit: " Ego praestolabor adventum tuum ".
JUDG|6|19|Ingressus est itaque Gedeon et coxit haedum et de farinae ephi azymos panes; carnesque ponens in canistro et ius carnium mittens in ollam tulit omnia sub quercum et obtulit ei.
JUDG|6|20|Cui dixit angelus Dei: " Tolle carnes et panes azymos et pone super petram illam et ius desuper funde ". Cumque fecisset ita,
JUDG|6|21|extendit angelus Domini summitatem virgae, quam tenebat in manu, et tetigit carnes et azymos panes, ascenditque ignis de petra et carnes azymosque panes consumpsit. Angelus autem Domini evanuit ex oculis eius.
JUDG|6|22|Vidensque Gedeon quod esset angelus Domini ait: "Heu mihi, Domine Deus, quia vidi angelum Domini facie ad faciem! ".
JUDG|6|23|Dixitque ei Dominus: " Pax tecum, ne timeas, non morieris! ".
JUDG|6|24|Aedificavit ergo ibi Gedeon altare Domino vocavitque illud: " Dominus pax "; usque in praesentem diem adhuc est in Ephra filiorum Abiezer.
JUDG|6|25|Nocte illa dixit Dominus ad eum: " Tolle taurum patris tui, alterum taurum scilicet annorum septem, destruesque aram Baal, quae est patris tui, et palum, qui iuxta aram est, succide;
JUDG|6|26|et aedificabis altare Domino Deo tuo in summitate petrae huius secundum ordinem; tollesque taurum secundum et offeres holocaustum super struem lignorum pali, quem succideris ".
JUDG|6|27|Assumptis igitur Gedeon decem viris de servis suis, fecit, sicut praeceperat Dominus; timens autem domum patris sui et homines illius civitatis per diem facere noluit, sed omnia nocte complevit.
JUDG|6|28|Cumque surrexissent viri oppidi eius mane, viderunt destructam aram Baal palumque succisum et taurum alterum impositum super altare, quod tunc aedificatum erat.
JUDG|6|29|Dixeruntque ad invicem: " Quis hoc fecit? ". Cumque perquirerent auctorem facti, dictum est: " Gedeon filius Ioas fecit haec omnia ".
JUDG|6|30|Et dixerunt ad Ioas: " Produc filium tuum, ut moriatur, quia destruxit aram Baal et succidit palum ".
JUDG|6|31|Respondit Ioas omnibus, qui circumdabant eum: " Numquid certare vultis pro Baal et salvare eum? Qui certabit pro Baal, morietur usque mane. Si Deus est, certet pro seipso contra eum, qui destruxit aram eius ".
JUDG|6|32|Ex illo die vocatus est Gedeon Ierobbaal, eo quod dicebatur: " Certet contra eum Baal, quia destruxit altare eius ".
JUDG|6|33|Igitur omnis Madian et Amalec et orientales populi congregati sunt simul et transeuntes Iordanem castrametati sunt in valle Iezrahel.
JUDG|6|34|Spiritus autem Domini induit Gedeon, qui clangens bucina convocavit domum Abiezer, ut sequeretur.
JUDG|6|35|Misitque nuntios in universum Manassen, qui et ipse secutus est eum; et alios nuntios in Aser et Zabulon et Nephthali, qui occurrerunt ei.
JUDG|6|36|Dixitque Gedeon ad Deum: " Si salvum facis per manum meam Israel, sicut locutus es,
JUDG|6|37|ponam vellus lanae in area: si ros in solo vellere fuerit, et in omni terra siccitas, sciam quod per manum meam, sicut locutus es, liberabis Israel ".
JUDG|6|38|Factumque est ita. Et de nocte consurgens, expresso vellere concham rore complevit.
JUDG|6|39|Dixitque rursus ad Deum: " Ne irascatur furor tuus contra me, si adhuc semel tentavero signum quaerens in vellere. Oro, ut solum vellus siccum sit, et omnis terra rore madens ".
JUDG|6|40|Fecitque Deus nocte illa, ut postulaverat; et fuit siccitas in solo vellere, et ros in omni terra.
JUDG|7|1|Igitur Ierobbaal, qui et Gedeon, de nocte consurgens et omnis populus cum eo castrame tati sunt ad fontem, qui vocatur Harad. Erant autem castra Madian in valle ad septentrionalem plagam collis Moreh.
JUDG|7|2|Dixitque Dominus ad Gedeon: " Maior tecum est populus, quam ut tradatur Madian in manus eius, ne glorietur contra me Israel et dicat: "Meis viribus liberatus sum".
JUDG|7|3|Loquere ad populum et, cunctis audientibus, praedica: "Qui formidolosus et timidus est, revertatur et recedat de monte Gelboe" ". Et reversa sunt ex populo viginti duo milia virorum; et tantum decem milia remanserunt.
JUDG|7|4|Dixitque Dominus ad Gedeon: " Adhuc populus multus est; duc eos ad aquas, et ibi probabo illos, et, de quo dixero tibi ut tecum vadat, ipse pergat; quem ire prohibuero, revertatur ".
JUDG|7|5|Cumque deduxisset populum ad aquas, dixit Dominus ad Gedeon: " Qui lingua lambuerint aquas, sicut solent canes lambere, separabis eos seorsum; qui autem curvatis genibus biberint, in altera parte erunt ".
JUDG|7|6|Fuit itaque numerus eorum, qui manu ad os proiciente aquas lambuerant, trecenti viri; omnis autem reliqua multitudo flexo poplite biberat.
JUDG|7|7|Et ait Dominus ad Gedeon: " In trecentis viris, qui lambuerunt aquas, liberabo vos et tradam Madian in manu tua; omnis autem reliqua multitudo revertatur in locum suum ".
JUDG|7|8|Sumptis itaque pro numero cibariis et tubis, omnem reliquam multitudinem abire praecepit ad tabernacula sua et ipse trecentos viros tenuit. Castra autem Madian erant subter eum in valle.
JUDG|7|9|Eadem nocte dixit Dominus ad eum: " Surge et descende in castra, quia tradidi ea in manu tua.
JUDG|7|10|Sin autem ire formidas, descendat tecum Phara puer tuus.
JUDG|7|11|Et, cum audieris quid loquantur, tunc confortabuntur manus tuae, et securior ad hostium castra descendes ". Descendit ergo ipse et Phara puer eius in partem castrorum, ubi erant armatorum vigiliae.
JUDG|7|12|Madian autem et Amalec et omnes orientales populi fusi iacebant in valle ut locustarum multitudo; cameli quoque innumerabiles erant sicut arena, quae iacet in litoribus maris.
JUDG|7|13|Cumque venisset Gedeon, narrabat aliquis somnium proximo suo et dicebat: " Ecce vidi somnium, et videbatur mihi quasi subcinericius panis ex hordeo volvi et in Madian castra descendere; cumque pervenisset ad tabernaculum, percussit illud atque subvertit et terrae funditus coaequavit ".
JUDG|7|14|Respondit is, cui loquebatur: "Non est hoc aliud nisi gladius Gedeonis filii Ioas viri Israelitae; tradidit Deus in manu eius Madian et omnia castra eius ".
JUDG|7|15|Cumque audisset Gedeon somnium et interpretationem eius, adoravit et reversus ad castra Israel ait: " Surgite, tradidit enim Dominus in manus vestras castra Madian ".
JUDG|7|16|Divisitque trecentos viros in tres partes et dedit tubas in manibus eorum lagoenasque vacuas ac lampades in medio lagoenarum
JUDG|7|17|et dixit ad eos: " Quod me facere videritis, hoc facite; ingrediar extremam partem castrorum, et, quod fecero, sectamini.
JUDG|7|18|Quando personaverit tuba in manu mea et omnium eorum, qui mecum sunt, vos quoque per castrorum circuitum clangite et conclamate: "Domino et Gedeoni!" ".
JUDG|7|19|Ingressusque est Gedeon et trecenti viri, qui erant cum eo, extremam partem castrorum, incipientibus vigiliis noctis mediae, cum eo ipso tempore custodes mutati essent, et coeperunt bucinis clangere et conterere lagoenas.
JUDG|7|20|Cumque in tribus personarent turmis et hydrias confregissent, tenuerunt sinistris manibus lampades et dextris sonantes tubas clamaveruntque: " Gladius Domino et Gedeoni! ",
JUDG|7|21|stantes singuli in loco suo per circuitum castrorum hostilium. Omnia itaque castra turbata sunt, et vociferantes ululantesque fugerunt.
JUDG|7|22|Et insistebant trecenti viri bucinis personantes. Immisitque Dominus gladium in omnibus castris, et mutua se caede truncabant fugientes usque Bethsetta, Sareda et crepidinem Abelmehula in Tebbath.
JUDG|7|23|Convocati autem viri Israel de Nephthali et Aser et omni Manasse persequebantur Madian.
JUDG|7|24|Misitque Gedeon nuntios in omnem montem Ephraim dicens: " Descendite in occursum Madian et occupate aquas usque Bethbera atque Iordanem ". Omnis Ephraim praeoccupavit aquas usque Bethbera atque Iordanem.
JUDG|7|25|Apprehensosque duos principes Madian Oreb et Zeb interfecit Oreb in Petra Oreb, Zeb vero in Torculari Zeb; et persecuti sunt Madian capita Oreb et Zeb portantes ad Gedeon trans fluenta Iordanis.
JUDG|8|1|Dixeruntque ad eum viri Ephraim: " Quid est hoc quod nobis facere voluisti, ut non nos vocares, cum ad pugnam pergeres contra Madian? ", iurgantes fortiter et prope vim inferentes.
JUDG|8|2|Quibus ille respondit: " Quid enim tale facere potui, quale vos fecistis? Nonne melior est racemus Ephraim vindemiis Abiezer?
JUDG|8|3|In manus vestras Deus tradidit principes Madian Oreb et Zeb. Quid tale facere potui, quale vos fecistis? ". Quod cum locutus esset, requievit spiritus eorum, quo tumebant contra eum.
JUDG|8|4|Cumque venisset Gedeon ad Iordanem, transivit eum cum trecentis viris, qui secum erant et prae lassitudine fugientes persequi vix poterant.
JUDG|8|5|Dixitque ad viros Succoth: "Date, obsecro, panes populo, qui mecum est, quia valde defecerunt, et ego persequor Zebee et Salmana reges Madian ".
JUDG|8|6|Responderunt principes Succoth: " Forsitan palmae manuum Zebee et Salmana in manu tua sunt, ut demus exercitui tuo panes? ".
JUDG|8|7|Quibus ille ait: " Cum ergo tradiderit Dominus Zebee et Salmana in manus meas, triturabo carnes vestras cum spinis deserti et tribulis ".
JUDG|8|8|Et inde conscendens venit in Phanuel locutusque est ad viros eius loci similia. Cui et illi responderunt, sicut responderant viri Succoth.
JUDG|8|9|Dixit itaque et eis: "Cum reversus fuero in pace, destruam turrim hanc".
JUDG|8|10|Zebee autem et Salmana requiescebant in Carcar cum omni exercitu suo, quasi quindecim milia viri, qui remanserant ex omnibus turmis orientalium populorum, caesis centum viginti milibus bellatorum educentium gladium.
JUDG|8|11|Ascendensque Gedeon per viam eorum, qui in tabernaculis morabantur ad orientalem partem Nobe et Iegbaa, percussit castra hostium, qui securi erant et nihil adversi suspicabantur.
JUDG|8|12|Fugeruntque Zebee et Salmana. Persequens Gedeon comprehendit duos reges Madian Zebee et Salmana, turbato omni exercitu eorum.
JUDG|8|13|Revertensque Gedeon filius Ioas de bello per ascensum Hares,
JUDG|8|14|apprehendit puerum de viris Succoth interrogavitque eum nomina principum et seniorum Succoth, qui scripsit ei septuaginta septem viros.
JUDG|8|15|Venitque ad viros Succoth et dixit eis: "En Zebee et Salmana, super quibus exprobrastis mihi dicentes: "Forsitan manus Zebee et Salmana in manibus tuis sunt, ut demus viris tuis, qui lassi sunt, panes?" ".
JUDG|8|16|Tulit ergo seniores civitatis et spinas deserti ac tribulos; et trituravit cum eis viros Succoth.
JUDG|8|17|Turrim quoque Phanuel subvertit, occisis habitatoribus civitatis.
JUDG|8|18|Dixitque ad Zebee et Salmana: " Quales fuerunt viri, quos occidistis in Thabor? ". Qui responderunt: " Similes tui, et unusquisque ex eis quasi filius regis ".
JUDG|8|19|Quibus ille ait: " Fratres mei fuerunt, filii matris meae. Vivit Dominus, si servassetis eos, non vos occiderem! ".
JUDG|8|20|Dixitque Iether primogenito suo: " Surge et interfice eos! ". Qui non eduxit gladium; timebat enim, quia adhuc puer erat.
JUDG|8|21|Dixeruntque Zebee et Salmana: " Tu surge et irrue in nos, quia iuxta aetatem robur est hominis ". Surrexit Gedeon et interfecit Zebee et Salmana et tulit lunulas, quibus colla camelorum eorum decorata erant.
JUDG|8|22|Dixeruntque viri Israel ad Gedeon: " Dominare nostri, tu et filius tuus et filius filii tui, quia liberasti nos de manu Madian ".
JUDG|8|23|Quibus ille ait: " Non dominabor vestri, nec dominabitur in vos filius meus, sed dominabitur Dominus ".
JUDG|8|24|Dixitque ad eos: " Unam petitionem postulo a vobis: date mihi unusquisque anulum ex praeda sua ". Anulos enim aureos Ismaelitae habere consuerant.
JUDG|8|25|Qui responderunt: " Libentissime dabimus ". Expandentesque super terram pallium proiecerunt in eo unusquisque anulum de praeda sua.
JUDG|8|26|Et fuit pondus postulatorum anulorum mille septingenti auri sicli absque lunulis et inauribus et vestibus purpureis, quibus Madian reges uti soliti erant, et praeter torques camelorum.
JUDG|8|27|Fecitque ex eo Gedeon ephod et posuit illud in civitate sua Ephra. Fornicatusque est omnis Israel in eo, et factum est Gedeoni et omni domui eius in ruinam.
JUDG|8|28|Humiliatus est autem Madian coram filiis Israel, nec potuerunt ultra elevare cervices, sed quievit terra per quadraginta annos, quibus Gedeon vivebat.
JUDG|8|29|Abiit itaque Ierobbaal filius Ioas et habitavit in domo sua;
JUDG|8|30|habuitque Gedeon septuaginta filios, qui egressi sunt de femore eius, eo quod multas haberet uxores.
JUDG|8|31|Concubina quoque illius, quam habebat in Sichem, genuit ei filium, cui ipse nomen imposuit Abimelech.
JUDG|8|32|Mortuusque est Gedeon filius Ioas in senectute bona et sepultus est in sepulcro Ioas patris sui in Ephra filiorum Abiezer.
JUDG|8|33|Postquam autem mortuus est Gedeon, aversi sunt filii Israel et fornicati cum Baalim posuerunt sibi Baalberith in deum.
JUDG|8|34|Nec recordati sunt Domini Dei sui, qui eruit eos de manu omnium inimicorum suorum per circuitum,
JUDG|8|35|nec fecerunt misericordiam cum domo Ierobbaal Gedeon iuxta omnia bona, quae fecerat Israeli.
JUDG|9|1|Abiit autem Abimelech filius Ierobbaal in Sichem ad fratres matris suae et locutus est ad eos et ad omnem cognationem familiae matris suae dicens:
JUDG|9|2|" Loquimini ad omnes viros Sichem: "Quid vobis est melius, ut dominentur vestri septuaginta viri, omnes filii Ierobbaal, an ut dominetur vobis unus vir? Simulque considerate quod os vestrum et caro vestra sum" ".
JUDG|9|3|Locutique sunt fratres matris eius de eo ad omnes viros Sichem universos sermones istos et inclinaverunt cor eorum post Abimelech dicentes: " Frater noster est ".
JUDG|9|4|Dederuntque illi septuaginta pondo argenti de fano Baalberith; qui conduxit sibi ex eo viros inopes et vagos, secutique sunt eum.
JUDG|9|5|Et venit in domum patris sui Ephra et occidit fratres suos filios Ierobbaal septuaginta viros super lapidem unum. Remansitque Ioatham filius Ierobbaal minimus, quia absconditus erat.
JUDG|9|6|Congregati sunt autem omnes viri Sichem et universae domus Mello abieruntque et constituerunt regem Abimelech iuxta quercum, quae stabat in Sichem.
JUDG|9|7|Quod cum nuntiatum esset Ioatham, ivit et stetit in vertice montis Garizim elevataque voce clamavit et dixit: " Audite me, viri Sichem, ut audiat vos Deus.
JUDG|9|8|Ierunt ligna, ut ungerent super se regem, dixeruntque olivae: "Impera nobis".
JUDG|9|9|Quae respondit: "Numquid possum deserere pinguedinem meam, qua et dii honorantur et homines, et venire, ut super ligna movear?".
JUDG|9|10|Dixeruntque ligna ad arborem ficum: "Veni et super nos regnum accipe".
JUDG|9|11|Quae respondit eis: "Numquid possum deserere dulcedinem meam fructusque suavissimos et ire, ut super cetera ligna movear?".
JUDG|9|12|Locuta quoque sunt ligna ad vitem: "Veni et impera nobis".
JUDG|9|13|Quae respondit: "Numquid possum deserere vinum meum, quod laetificat deos et homines, et super ligna cetera commoveri?".
JUDG|9|14|Dixeruntque omnia ligna ad rhamnum: "Veni et impera super nos".
JUDG|9|15|Quae respondit eis: "Si vere me regem vobis constituitis, venite et sub mea umbra requiescite; sin autem non vultis, egrediatur ignis de rhamno et devoret cedros Libani!".
JUDG|9|16|Nunc igitur, si recte et absque peccato constituistis super vos regem Abimelech et bene egistis cum Ierobbaal et cum domo eius et reddidistis vicem beneficiis eius,
JUDG|9|17|qui pugnavit pro vobis et animam suam dedit periculis, ut erueret vos de manu Madian,
JUDG|9|18|qui nunc surrexistis contra domum patris mei et interfecistis filios eius septuaginta viros super unum lapidem et constituistis regem Abimelech filium ancillae eius super habitatores Sichem, eo quod frater vester sit;
JUDG|9|19|si ergo recte et absque vitio egistis cum Ierobbaal et domo eius hodie, laetamini in Abimelech, et ille laetetur in vobis.
JUDG|9|20|Sin autem perverse, egrediatur ignis ex Abimelech et consumat habitatores Sichem et domum Mello, egrediaturque ignis de viris Sichem et de domo Mello et devoret Abimelech! ".
JUDG|9|21|Quae cum Ioatham dixisset, fugit et abiit in Bera habitavitque ibi metu Abimelech fratris sui.
JUDG|9|22|Regnavit itaque Abimelech super Israel tribus annis.
JUDG|9|23|Misitque Deus spiritum pessimum inter Abimelech et habitatores Sichem, qui rebellaverunt contra eum,
JUDG|9|24|ut scelus interfectionis septuaginta filiorum Ierobbaal et effusio sanguinis eorum veniret super Abimelech fratrem suum et in viros Sichimorum, qui eum adiuverant.
JUDG|9|25|Posueruntque insidias adversus eum in montium summitate et exercebant latrocinia agentes praedas de omnibus praetereuntibus. Nuntiatumque est Abimelech.
JUDG|9|26|Venit autem Gaal filius Ebed cum fratribus suis et transivit in Sichimam, et confisi sunt habitatores Sichem in eo.
JUDG|9|27|Egressi in agros vindemiaverunt vineas uvasque calcaverunt et, factis cantantium choris, ingressi sunt fanum dei sui et inter epulas et pocula maledicebant Abimelech,
JUDG|9|28|clamante Gaal filio Ebed: " Quis est Abimelech, et quae est Sichem, ut serviamus ei? Numquid non est filius Ierobbaal et Zebul praefectus eius? Servite viris Hemmor patris Sichem! Cur serviemus ei?
JUDG|9|29|Utinam daret aliquis populum istum sub manu mea, ut auferrem de medio Abimelech et dicerem ei: Congrega exercitus multitudinem et veni ".
JUDG|9|30|Zebul princeps civitatis, auditis sermonibus Gaal filii Ebed, iratus est valde
JUDG|9|31|et misit clam ad Abimelech nuntios dicens: " Ecce Gaal filius Ebed venit in Sichimam cum fratribus suis et excitant adversum te civitatem.
JUDG|9|32|Surge itaque nocte cum populo, qui tecum est, et latita in agro.
JUDG|9|33|Et primo mane, oriente sole, irrue super civitatem; illo autem egrediente adversum te cum populo suo, fac ei, quod potueris ".
JUDG|9|34|Surrexit itaque Abimelech cum omni exercitu suo nocte et tetendit insidias iuxta Sichimam in quattuor locis.
JUDG|9|35|Egressusque est Gaal filius Ebed et stetit in introitu portae civitatis; surrexit autem Abimelech et omnis exercitus cum eo de insidiarum loco.
JUDG|9|36|Cumque vidisset populum Gaal, dixit ad Zebul: " Ecce de montibus multitudo descendit ". Cui ille respondit: " Umbras montium vides quasi homines ".
JUDG|9|37|Rursumque Gaal ait: " Ecce populus de Umbilico terrae descendit, et unus cuneus venit per viam Quercus Augurum ".
JUDG|9|38|Cui dixit Zebul: " Ubi est nunc os tuum, quo loquebaris: "Quis est Abimelech, ut serviamus ei?". Nonne iste est populus, quem despiciebas? Egredere et pugna contra eum ".
JUDG|9|39|Abiit ergo Gaal, spectante Sichimorum populo, et pugnavit contra Abimelech.
JUDG|9|40|Qui persecutus est eum fugientem, cecideruntque ex parte eius plurimi usque ad portam civitatis.
JUDG|9|41|Et Abimelech sedit in Aruma; Zebul autem Gaal et fratres eius expulit de urbe nec in ea passus est commorari.
JUDG|9|42|Sequenti ergo die egressus est populus in campum. Quod cum nuntiatum esset Abimelech,
JUDG|9|43|tulit exercitum suum et divisit in tres turmas tendens insidias in agris. Vidensque quod egrederetur populus de civitate, surrexit et percussit eos.
JUDG|9|44|Irruensque cum cuneo suo obsedit ingressum portae civitatis; duae autem turmae palantes per campum adversarios percusserunt.
JUDG|9|45|Porro Abimelech omni illo die oppugnabat urbem, quam cepit, interfectis habitatoribus eius ipsaque destructa, ita ut sal in ea dispergeret.
JUDG|9|46|Quod cum audissent, qui habitabant in turre Sichimorum, ingressi sunt cryptam fani Elberith (id est dei Foederis).
JUDG|9|47|Abimelech quoque audiens omnes viros turris Sichimorum pariter conglobatos,
JUDG|9|48|ascendit in montem Selmon cum omni populo suo et, arrepta securi, praecidit arboris ramum impositumque ferens umero dixit ad socios: " Quod me viditis facere, cito facite ".
JUDG|9|49|Igitur certatim ramos de arboribus praecidentes sequebantur ducem, quos circumdantes cryptae succenderunt; atque ita factum est, ut fumo et igne omnes homines necarentur, circiter mille viri pariter ac mulieres, habitatores turris Sichem.
JUDG|9|50|Abimelech autem inde proficiscens venit ad oppidum Thebes, quod obsidebat et cepit.
JUDG|9|51|Erat autem turris fortis in media civitate, ad quam confugerant viri simul ac mulieres et omnes cives civitatis, clausa firmissime ianua, et super turris tectum stantes per propugnacula.
JUDG|9|52|Accedensque Abimelech iuxta turrim pugnabat fortiter et appropinquans ostio ignem supponere nitebatur.
JUDG|9|53|Et ecce una mulier superiorem molam desuper iaciens illisit capiti Abimelech et confregit cerebrum eius.
JUDG|9|54|Qui vocavit cito armigerum suum et ait ad eum: " Evagina gladium tuum et percute me, ne forte dicatur quod a femina interfectus sim ". Qui transfodit eum.
JUDG|9|55|Illoque mortuo, omnes viri Israel hoc videntes reversi sunt in sedes suas.
JUDG|9|56|Et reddidit Deus malum, quod fecerat Abimelech contra patrem suum, interfectis septuaginta fratribus suis.
JUDG|9|57|Sichimitis quoque, quod operati erant, retributum est, et venit super eos maledictio Ioatham filii Ierobbaal.
JUDG|10|1|Post Abimelech surrexit dux ad salvandum Israel Thola fi lius Phua filii Dodo, vir de Issachar, qui habitavit in Samir montis Ephraim.
JUDG|10|2|Et iudicavit Israel viginti et tribus annis mortuusque ac sepultus est in Samir.
JUDG|10|3|Huic successit Iair Galaadites, qui iudicavit Israel per viginti et duos annos
JUDG|10|4|habens triginta filios sedentes super triginta pullos asinarum, et ipsis erant triginta civitates, quae appellatae sunt Havoth Iair (id est villae Iair) usque in praesentem diem, in terra Galaad.
JUDG|10|5|Mortuusque est Iair ac sepultus in Camon.
JUDG|10|6|Filii autem Israel peccatis veteribus iungentes nova fecerunt malum in conspectu Domini et servierunt Baalim et Astharoth et diis Syriae ac Sidonis et Moab et filiorum Ammon et Philisthim; dimiseruntque Dominum et non colebant eum.
JUDG|10|7|Contra quos iratus tradidit eos in manu Philisthim et filiorum Ammon.
JUDG|10|8|Afflictique sunt et vehementer oppressi per annos decem et octo omnes filii Israel, qui habitabant trans Iordanem in terra Amorraei in Galaad;
JUDG|10|9|in tantum ut filii Ammon Iordanem transirent ad pugnandum etiam contra Iudam et Beniamin et domum Ephraim; afflictusque est Israel nimis.
JUDG|10|10|Et clamantes filii Israel ad Dominum dixerunt: " Peccavimus tibi, quia dereliquimus Deum nostrum et servivimus Baalim ".
JUDG|10|11|Quibus locutus est Dominus: " Numquid non Aegyptii et Amorraei filiique Ammon et Philisthim,
JUDG|10|12|Sidonii quoque et Amalec et Madian oppresserunt vos, et clamastis ad me, et erui vos de manu eorum?
JUDG|10|13|Et tamen reliquistis me et coluistis deos alienos; idcirco non addam ut ultra vos liberem.
JUDG|10|14|Ite et invocate deos, quos elegistis: ipsi vos liberent in tempore angustiae! ".
JUDG|10|15|Dixeruntque filii Israel ad Dominum: "Peccavimus; redde tu nobis, quidquid tibi placet, tantum nunc libera nos ".
JUDG|10|16|Quae dicentes omnia de finibus suis alienorum deorum idola proiecerunt et servierunt Domino, qui doluit super miseriis Israel.
JUDG|10|17|Itaque filii Ammon convocati in Galaad fixere tentoria; contra quos congregati filii Israel in Maspha castrametati sunt.
JUDG|10|18|Dixeruntque populus, principes Galaad, singuli ad proximos suos: " Qui primus contra filios Ammon coeperit dimicare, erit dux omnium habitatorum Galaad ".
JUDG|11|1|Fuit Iephte Galaadites vir fortissimus, filius meretricis mulieris, quem genuit Galaad.
JUDG|11|2|Habuit autem Galaad uxorem, de qua suscepit filios, qui, postquam creverant, eiecerunt Iephte dicentes: " Heres in domo patris nostri esse non poteris, quia de altera matre generatus es ".
JUDG|11|3|Quos ille fugiens atque devitans habitavit in terra Tob; congregatique sunt ad eum viri inopes et exierunt cum eo.
JUDG|11|4|In illis diebus pugnabant filii Ammon contra Israel.
JUDG|11|5|Quibus acriter instantibus, perrexerunt maiores natu de Galaad, ut tollerent in auxilium sui Iephte de terra Tob.
JUDG|11|6|Dixeruntque ad eum: " Veni et esto princeps noster, et pugnemus contra filios Ammon ".
JUDG|11|7|Quibus ille respondit: " Nonne vos estis, qui odistis me et eiecistis de domo patris mei? Et nunc venistis ad me necessitate compulsi ".
JUDG|11|8|Dixeruntque principes Galaad ad Iephte: " Ob hanc igitur causam nunc ad te venimus, ut proficiscaris nobiscum et pugnes contra filios Ammon sisque dux omnium, qui habitant in Galaad ".
JUDG|11|9|Iephte quoque dixit eis: " Si revocatis me, ut pugnem pro vobis contra filios Ammon, tradideritque eos Dominus in manus meas, ego ero princeps vester ".
JUDG|11|10|Qui responderunt ei: " Dominus, qui haec audit, ipse mediator ac testis est quod secundum verbum tuum faciemus ".
JUDG|11|11|Abiit itaque Iephte cum principibus Galaad, fecitque eum omnis populus principem sui. Locutusque est Iephte omnes sermones suos coram Domino in Maspha.
JUDG|11|12|Et misit Iephte nuntios ad regem filiorum Ammon, qui ex persona sua dicerent: " Quid mihi et tibi est, quia venisti contra me, ut invaderes terram meam? ".
JUDG|11|13|Quibus ille respondit: " Quia tulit Israel terram meam, quando ascendit de Aegypto, a finibus Arnon usque Iaboc atque Iordanem; nunc igitur cum pace redde mihi eam ".
JUDG|11|14|Rursumque Iephte nuntios misit et imperavit eis, ut dicerent regi Ammon:
JUDG|11|15|" Haec dicit Iephte: Non tulit Israel terram Moab nec terram filiorum Ammon.
JUDG|11|16|Sed, quando de Aegypto conscenderunt, ambulavit Israel per solitudinem usque ad mare Rubrum et venit in Cades;
JUDG|11|17|misitque nuntios ad regem Edom dicens: "Dimitte, ut transeam per terram tuam". Qui noluit acquiescere precibus eius. Misit quoque et ad regem Moab, qui et ipse transitum praebere contempsit. Mansit itaque Israel in Cades
JUDG|11|18|et pertransiens desertum circuivit ex latere terram Edom et terram Moab venitque contra orientalem plagam terrae Moab et castrametatus est trans Arnon nec voluit intrare terminos Moab; Arnon quippe confinium est terrae Moab.
JUDG|11|19|Misit itaque Israel nuntios ad Sehon regem Amorraeorum, regem Hesebon, et dixit ei: "Dimitte, ut transeam per terram tuam usque ad locum meum".
JUDG|11|20|Qui et ipse Israel verbis diffidens non dimisit eum transire per terminos suos, sed, omni populo suo congregato, egressus est contra eum in Iasa et fortiter resistebat.
JUDG|11|21|Tradiditque eum Dominus in manu Israel cum omni exercitu suo, qui percussit eum et possedit omnem terram Amorraei habitatoris regionis illius,
JUDG|11|22|universos fines eius de Arnon usque Iaboc et de solitudine usque ad Iordanem.
JUDG|11|23|Dominus ergo, Deus Israel, subvertit Amorraeum coram populo suo Israel; et tu nunc vis possidere terram eius?
JUDG|11|24|Nonne ea, quae tibi Chamos deus tuus in possessionem dat, tibi iure debentur? Quae autem Dominus Deus noster victor obtinuit, in nostram cedunt possessionem.
JUDG|11|25|Num quid melior es Balac filio Sephor rege Moab? Numquid iurgatus est contra Israel et pugnavit contra eum?
JUDG|11|26|Quando habitabat in Hesebon et viculis eius et in Aroer et villis illius et in cunctis civitatibus iuxta Arnon per trecentos annos, quare tanto tempore nihil super hac repetitione tentastis?
JUDG|11|27|Igitur non ego pecco in te, sed tu contra me male agis indicens mihi bella non iusta. Iudicet Dominus arbiter huius diei inter filios Israel et inter filios Ammon ".
JUDG|11|28|Noluitque acquiescere rex filiorum Ammon verbis Iephte, quae per nuntios mandaverat.
JUDG|11|29|Factus est ergo super Iephte spiritus Domini, et pertransiens Galaad et Manasse venit in Maspha Galaad et inde ad filios Ammon.
JUDG|11|30|Votum autem vovit Domino dicens: " Si tradideris filios Ammon in manus meas,
JUDG|11|31|quicumque primus fuerit egressus de foribus domus meae mihique occurrerit revertenti cum pace a filiis Ammon, eum holocaustum offeram Domino ".
JUDG|11|32|Transivitque Iephte ad filios Ammon, ut pugnaret contra eos; quos tradidit Dominus in manus eius.
JUDG|11|33|Percussitque eos ab Aroer usque dum venias in Mennith viginti civitates et usque ad Abelcharmim plaga magna nimis; humiliatique sunt filii Ammon a filiis Israel.
JUDG|11|34|Revertenti autem Iephte in Maspha domum suam occurrit unigenita filia cum tympanis et choris: non enim habebat alios liberos.
JUDG|11|35|Qua visa, scidit vestimenta sua et ait: " Heu, filia mi, incurvans incurvasti me! Et tu es in eis, qui me perturbant! Aperui enim os meum ad Dominum et aliud facere non potero ".
JUDG|11|36|Cui illa respondit: " Pater mi, si aperuisti os tuum ad Dominum, fac mihi, quodcumque pollicitus es, concessa tibi a Domino ultione atque victoria de hostibus tuis filiis Ammon ".
JUDG|11|37|Dixitque ad patrem: " Hoc solum mihi praesta, quod deprecor: Dimitte me, ut duobus mensibus circumeam montes et plangam virginitatem meam cum sodalibus meis ".
JUDG|11|38|Cui ille respondit: " Vade! ". Et dimisit eam duobus mensibus. Cumque abisset cum sodalibus suis, flebat virginitatem suam in montibus.
JUDG|11|39|Expletisque duobus mensibus, reversa est ad patrem suum; et fecit ei, sicut voverat, quae non cognoverat virum. Exinde mos increbuit in Israel, et consuetudo servata est,
JUDG|11|40|ut post anni circulum conveniant in unum filiae Israel et plangant filiam Iephte Galaaditae diebus quattuor.
JUDG|12|1|Ecce autem convocatus vir Ephraim transiit contra aqui lonem, et dixerunt ad Iephte: " Quare vadens ad pugnam contra filios Ammon vocare nos noluisti, ut pergeremus tecum? Igitur incendemus domum tuam super te.
JUDG|12|2|Quibus ille respondit: " Disceptatio erat mihi et populo meo contra filios Ammon vehemens, vocavique vos, ut mihi praeberetis auxilium, et facere noluistis.
JUDG|12|3|Quod cernens posui in manibus meis animam meam transivique ad filios Ammon, et tradidit eos Dominus in manus meas. Quid commerui, ut hodie adversum me consurgatis in proelium? ".
JUDG|12|4|Vocatis itaque ad se cunctis viris Galaad, pugnabat contra Ephraim. Percusseruntque viri Galaad Ephraim, quia dixerat: " Fugitivi de Ephraim estis; Galaad habitat in medio Ephraim et Manasse ".
JUDG|12|5|Occupaveruntque Galaaditae vada Iordanis, per quae Ephraim reversurus erat. Cumque venisset ad ea de Ephraim numero fugiens atque dixisset: " Obsecro, ut me transire permittatis ", dicebant ei Galaaditae: " Numquid Ephrathaeus es? ". Quo dicente: " Non sum ",
JUDG|12|6|interrogabant eum: " Dic ergo: Scibboleth " (quod interpretatur Spica). Qui respondebat: " Sibboleth ", illud recte exprimere non valens. Statimque apprehensum iugulabant in ipso Iordanis transitu. Et ceciderunt in illo tempore de Ephraim quadraginta duo milia.
JUDG|12|7|Iudicavitque Iephte Galaadites Israel sex annis et mortuus est ac sepultus in civitate sua in Galaad.
JUDG|12|8|Post hunc iudicavit Israel Abesan de Bethlehem.
JUDG|12|9|Qui habuit triginta filios et totidem filias emittens foras maritis dedit; et eiusdem numeri filiis suis accepit uxores forinsecus. Qui septem annis iudicavit Israel;
JUDG|12|10|mortuusque est ac sepultus in Bethlehem.
JUDG|12|11|Cui successit Ahialon Zabulonites et iudicavit Israel decem annis;
JUDG|12|12|mortuusque est ac sepultus in Ahialon terrae Zabulon.
JUDG|12|13|Post hunc iudicavit Israel Abdon filius Illel Pharathonites.
JUDG|12|14|Qui habuit quadraginta filios et triginta ex eis nepotes ascendentes super septuaginta pullos asinarum. Et iudicavit Israel octo annis;
JUDG|12|15|mortuusque est ac sepultus in Pharathon terrae Ephraim in monte Amalecite.
JUDG|13|1|Rursumque filii Israel fece runt malum in conspectu Do mini, qui tradidit eos in manus Philisthinorum quadraginta annis.
JUDG|13|2|Erat autem vir quidam de Saraa et de stirpe Dan nomine Manue habens uxorem sterilem.
JUDG|13|3|Cui apparuit angelus Domini et dixit ad eam: " Ecce sterilis es et absque liberis, sed concipies et paries filium.
JUDG|13|4|Cave ergo, ne vinum bibas ac siceram nec immundum quidquam comedas,
JUDG|13|5|quia ecce concipies et paries filium, cuius non tanget caput novacula: erit enim puer nazaraeus Dei ex matris utero et ipse incipiet liberare Israel de manu Philisthinorum ".
JUDG|13|6|Quae cum venisset ad maritum, dixit ei: " Vir Dei venit ad me habens aspectum sicut angelus Domini, terribilis nimis. Non interrogavi eum, unde esset, nec ipse nomen suum mihi indicavit.
JUDG|13|7|Et dixit mihi: "Ecce concipies et paries filium; cave, ne vinum bibas et siceram et ne aliquo vescaris immundo: erit enim puer nazaraeus Dei ex utero matris usque ad diem mortis suae" ".
JUDG|13|8|Oravit itaque Manue Dominum et ait: " Obsecro, Domine, ut vir Dei, quem misisti, veniat iterum et doceat nos, quid debeamus facere de puero, qui nasciturus est ".
JUDG|13|9|Exaudivitque Deus precantem Manue, et venit rursum angelus Dei ad mulierem sedentem in agro. Manue autem maritus eius non erat cum ea.
JUDG|13|10|Festinavit ergo et cucurrit ad virum suum nuntiavitque ei dicens: " Ecce apparuit mihi vir, qui illo die venerat ad me ".
JUDG|13|11|Qui surrexit et secutus est uxorem suam veniensque ad virum dixit ei: " Tu es, qui locutus es mulieri? ". Et ille respondit: " Ego sum ".
JUDG|13|12|Cui Manue: " Quando, inquit, sermo tuus fuerit expletus, quid circa puerum observare et facere debemus? ".
JUDG|13|13|Dixitque angelus Domini ad Manue: " Ab omnibus, quae locutus sum uxori tuae, abstineat se;
JUDG|13|14|et, quidquid ex vinea nascitur, non comedat, vinum et siceram non bibat, nullo vescatur immundo et, quod ei praecepi, custodiat ".
JUDG|13|15|Dixitque Manue ad angelum Domini: " Obsecro, ut retineamus te et faciamus tibi haedum de capris ".
JUDG|13|16|Cui respondit angelus Domini: " Si me retines, non comedam panes tuos; sin autem vis holocaustum facere, offer illud Domino ". Et nesciebat Manue quod angelus Domini esset.
JUDG|13|17|Dixitque ad eum: " Quod est tibi nomen, ut, si sermo tuus fuerit expletus, honoremus te? ".
JUDG|13|18|Cui ille respondit: " Cur quaeris nomen meum, quod est mirabile? ".
JUDG|13|19|Tulit itaque Manue haedum de capris et oblationem similae et posuit super petram offerens Domino, qui facit mirabilia; ipse autem et uxor eius intuebantur.
JUDG|13|20|Cumque ascenderet flamma de altari in caelum, angelus Domini in flamma pariter ascendit. Quod cum vidisset Manue et uxor eius, proni ceciderunt in terram;
JUDG|13|21|et ultra non eis apparuit angelus Domini. Statimque intellexit Manue angelum esse Domini
JUDG|13|22|et dixit ad uxorem suam: " Morte moriemur, quia vidimus Deum ".
JUDG|13|23|Cui respondit mulier: " Si Dominus nos vellet occidere, de manibus nostris holocaustum et oblationem non suscepisset nec ostendisset nobis haec omnia neque talia dixisset ".
JUDG|13|24|Peperit itaque filium et vocavit nomen eius Samson. Crevitque puer, et benedixit ei Dominus.
JUDG|13|25|Coepitque spiritus Domini impellere eum in Castris Dan inter Saraa et Esthaol.
JUDG|14|1|Descendit igitur Samson in Thamna vidensque ibi mulie rem de filiabus Philisthim
JUDG|14|2|ascendit et nuntiavit patri suo et matri dicens: " Vidi mulierem in Thamna de filiabus Philisthinorum, quam quaeso ut mihi accipiatis uxorem.
JUDG|14|3|Cui dixerunt pater et mater sua: " Numquid non est mulier in filiabus fratrum tuorum et in omni populo meo, quia vis accipere uxorem de Philisthim, qui incircumcisi sunt? ". Dixitque Samson ad patrem suum: " Hanc mihi accipe, quia placuit oculis meis ".
JUDG|14|4|Parentes autem eius nesciebant quod res a Domino fieret, et quaereret occasionem contra Philisthim. Eo enim tempore Philisthim dominabantur Israeli.
JUDG|14|5|Descendit itaque Samson cum patre suo et matre in Thamna. Cumque venissent ad vineas oppidi, apparuit catulus leonis rugiens et occurrit ei.
JUDG|14|6|Irruit autem spiritus Domini in Samson, et dilaceravit leonem, quasi haedum in frusta concerperet, nihil omnino habens in manu; et hoc patri et matri noluit indicare.
JUDG|14|7|Descenditque et locutus est mulieri, quae placuerat oculis eius.
JUDG|14|8|Et post aliquot dies revertens, ut acciperet eam, declinavit, ut videret cadaver leonis; et ecce examen apum in corpore leonis erat ac favus mellis.
JUDG|14|9|Quem, cum sumpsisset in manibus, comedebat in via; veniensque ad patrem suum et matrem dedit eis partem, qui et ipsi comederunt. Nec tamen eis voluit indicare quod mel de corpore leonis assumpserat.
JUDG|14|10|Descendit itaque pater eius ad mulierem, et fecit ibi Samson convivium; sic enim iuvenes facere consuerant.
JUDG|14|11|Cum ergo cives loci illius vidissent eum, dederunt ei sodales triginta, qui essent cum eo.
JUDG|14|12|Quibus locutus est Samson: " Proponam vobis problema, quod si solveritis mihi intra septem dies convivii, dabo vobis triginta tunicas et totidem vestes mutatorias;
JUDG|14|13|sin autem non potueritis solvere, vos dabitis mihi triginta tunicas et eiusdem numeri vestes mutatorias ". Qui responderunt ei: " Propone problema, ut audiamus ".
JUDG|14|14|Dixitque eis: De comedente exivit cibus,et de forti est egressa dulcedo ".Nec potuerunt per tres dies propositionem solvere.
JUDG|14|15|Cumque adesset dies quartus, dixerunt ad uxorem Samson: " Blandire viro tuo et suade ei, ut indicet tibi quid significet problema. Quod si facere nolueris, incendemus et te et domum patris tui. An idcirco nos vocastis ad nuptias, ut spoliaretis? ".
JUDG|14|16|Quae fundebat apud Samson lacrimas et querebatur dicens: " Odisti me et non diligis; idcirco problema, quod proposuisti filiis populi mei, non vis mihi exponere ". At ille respondit: " Patri meo et matri nolui dicere et tibi indicare potero? ".
JUDG|14|17|Septem igitur diebus convivii flebat apud eum; tandemque die septimo, cum ei molesta esset, exposuit. Quae statim indicavit civibus suis,
JUDG|14|18|et illi dixerunt ei die septimo ante solis occubitum: Quid dulcius melle,et quid leone fortius? ".Qui ait ad eos: Si non arassetis in vitula mea,non invenissetis propositionem meam ".
JUDG|14|19|Irruit itaque in eo spiritus Domini, descenditque Ascalonem et percussit ibi triginta viros, quorum ablatas vestes dedit iis, qui problema solverant; iratusque nimis ascendit in domum patris sui.
JUDG|14|20|Uxor autem eius accepit maritum unum de amicis eius, qui erat pronubus.
JUDG|15|1|Post aliquantum autem tem poris, cum dies triticeae mes sis instarent, venit Samson invisere volens uxorem suam et attulit ei haedum de capris. Cumque ad eam vellet intrare, prohibuit eum pater illius
JUDG|15|2|dicens: " Putavi quod odisses eam et ideo tradidi illam amico tuo; sed habet sororem iuniorem, quae pulchrior illa est; sit tibi pro ea uxor ".
JUDG|15|3|Dixitque eis Samson: " Hac vice non erit culpa in me contra Philisthaeos, cum faciam eis mala ".
JUDG|15|4|Perrexitque et cepit trecentas vulpes caudasque earum iunxit ad caudas sumensque faces ligavit singulas in medio binarum caudarum;
JUDG|15|5|facibusque igne succensis, dimisit vulpes in segetes Philisthinorum. Et comportatae iam fruges et adhuc stantes in stipula concrematae sunt in tantum, ut vineas quoque et oliveta flamma consumeret.
JUDG|15|6|Dixeruntque Philisthim: " Quis fecit hanc rem? ". Quibus dictum est: " Samson gener Thamnathaei, quia tulit uxorem eius et alteri tradidit, haec operatus est ". Ascenderuntque Philisthim et combusserunt tam mulierem quam patrem eius.
JUDG|15|7|Quibus ait Samson: " Si talia facitis, utique ex vobis expetam ultionem et tunc quiescam ".
JUDG|15|8|Percussitque eos ingenti plaga, suram ad femur. Et descendens habitavit in spelunca petrae Etam.
JUDG|15|9|Igitur ascendentes Philisthim in terra Iudae castrametati sunt, et in Lehi (id est Maxilla) eorum est fusus exercitus.
JUDG|15|10|Dixeruntque ad eos viri de tribu Iudae: " Cur ascendistis adversum nos?. Qui responderunt: " Ut ligemus Samson venimus et reddamus ei, quae in nos operatus est ".
JUDG|15|11|Descenderunt ergo tria milia virorum de Iuda ad specum petrae Etam dixeruntque ad Samson: " Nescis quod Philisthim imperent nobis? Quare hoc nobis facere voluisti? ". Quibus ille ait: " Sicut fecerunt mihi, feci eis.
JUDG|15|12|" Ligare, inquiunt, te venimus et tradere in manus Philisthinorum ". " Iurate, respondit, mihi quod non me occidatis ".
JUDG|15|13|Dixerunt: " Non te occidemus, sed vinctum trademus ". Ligaveruntque eum duobus novis funibus et tulerunt de petra Etam.
JUDG|15|14|Qui cum venisset in Lehi, et Philisthim vociferantes occurrissent ei, irruit spiritus Domini in eum, et, sicut solent ad odorem ignis lina consumi, ita vincula, quibus brachia eius ligata erant, dissipata sunt et soluta.
JUDG|15|15|Inventamque maxillam asini recentem arripiens percussit in ea mille viros
JUDG|15|16|et ait: In maxilla asiniacervum feci ex eis!In mandibula asinipercussi mille viros! ".
JUDG|15|17|Cumque haec canens verba complesset, proiecit mandibulam de manu et vocavit nomen loci illius Ramathlehi (quod interpretatur Elevatio maxillae).
JUDG|15|18|Sitiensque valde clamavit ad Dominum et ait: " Tu dedisti in manu servi tui salutem hanc maximam atque victoriam; et en siti morior incidamque in manus incircumcisorum ".
JUDG|15|19|Aperuit itaque Deus fossam in Lehi, et egressae sunt inde aquae; quibus haustis, refocillavit spiritum et vires recepit. Idcirco appellatum est nomen fontis illius fons Invocantis, qui est in Lehi usque in praesentem diem.
JUDG|15|20|Iudicavitque Israel in diebus Philisthim viginti annis.
JUDG|16|1|Abiit Samson in Gazam et vidit ibi meretricem mulie rem ingressusque est ad eam.
JUDG|16|2|Cum nuntiatum esset Gazaeis intrasse urbem Samson, circuierunt et insidiabantur ei in porta civitatis; tota autem nocte quieverunt praestolantes, ut, facto mane, exeuntem occiderent.
JUDG|16|3|Dormivit autem Samson usque ad noctis medium et inde consurgens apprehendit ambas portae fores cum postibus suis et evellit eas cum sera, impositasque umeris portavit ad verticem montis, qui respicit Hebron.
JUDG|16|4|Post haec amavit mulierem, quae habitabat in valle Sorec et vocabatur Dalila.
JUDG|16|5|Veneruntque ad eam principes Philisthinorum atque dixerunt: " Decipe eum et disce ab illo in quo tantam habeat fortitudinem, et quomodo eum superare valeamus et vinctum humiliare; quod si feceris, dabimus tibi singuli mille centum argenteos ".
JUDG|16|6|Locuta est ergo Dalila ad Samson: " Dic mihi, obsecro, in quo sit tua maxima fortitudo, et quid sit, quo ligatus humilieris ".
JUDG|16|7|Cui respondit Samson: " Si septem nerviceis funibus necdum siccis et adhuc humentibus ligatus fuero, deficiam eroque ut ceteri homines ".
JUDG|16|8|Attuleruntque ad eam satrapae Philisthinorum septem funes, ut dixerat; quibus vinxit eum,
JUDG|16|9|latentibus apud se insidiis in cubiculo. Clamavitque ad eum: " Philisthim super te, Samson! ". Qui rupit vincula, quomodo si rumpat quis filum de stuppa tortum, cum odorem ignis acceperit; et non est cognitum in quo esset fortitudo eius.
JUDG|16|10|Dixitque ad eum Dalila: " Ecce illusisti mihi et falsum locutus es; saltem nunc indica mihi quo ligari debeas ".
JUDG|16|11|Cui ille respondit: " Si ligatus fuero novis funibus, qui numquam fuerunt in opere, infirmus ero et aliorum hominum similis ".
JUDG|16|12|Quibus rursum Dalila vinxit eum et clamavit: " Philisthim super te, Samson! ", in cubiculo insidiis praeparatis. Qui ita rupit vincula brachiorum quasi fila telarum.
JUDG|16|13|Dixitque Dalila rursum ad eum: " Usquequo decipis me et falsum loqueris? Ostende quo vinciri debeas ". Cui respondit Samson: " Si septem crines nexos capitis mei cum licio plexueris et paxillo fixeris, deficiam eroque ut ceteri homines ".
JUDG|16|14|Quae cum dormire eum fecisset et septem crines nexos capitis eius cum licio plexisset et paxillo fixisset, dixit ad eum: " Philisthim super te, Samson! ". Qui consurgens de somno extraxit paxillum cum navicula et licio.
JUDG|16|15|Dixitque ad eum Dalila: " Quomodo dicis quod ames me, cum animus tuus non sit mecum? Per tres vices mentitus es mihi et noluisti dicere in quo sit tua maxima fortitudo ".
JUDG|16|16|Cumque molesta ei esset et per multos dies iugiter eum urgeret, defecit anima eius et ad mortem usque lassata est.
JUDG|16|17|Tunc aperiens ei totum cor suum dixit ad eam: " Novacula numquam ascendit super caput meum, quia nazaraeus consecratus Deo sum de utero matris meae; si rasum fuerit caput meum, recedet a me fortitudo mea, et deficiam eroque ut ceteri homines ".
JUDG|16|18|Videns illa quod confessus ei esset omnem animum suum, misit ad principes Philisthinorum atque mandavit: " Ascendite adhuc semel, quia nunc mihi aperuit totum cor suum ". Qui ascenderunt, assumpta pecunia, quam promiserant.
JUDG|16|19|At illa dormire eum fecit super genua sua vocavitque tonsorem et fecit radere septem crines eius et coepit humiliare eum; statim enim ab eo fortitudo discessit.
JUDG|16|20|Dixitque: " Philisthim super te, Samson! ". Qui de somno consurgens dixit in animo suo: " Egrediar, sicut ante feci, et me excutiam ", nesciens quod Dominus recessisset ab eo.
JUDG|16|21|Quem cum apprehendissent Philisthim, statim eruerunt oculos eius et duxerunt Gazam vinctum duabus catenis aeneis et clausum in carcere molere fecerunt.
JUDG|16|22|Iamque capilli eius renasci coeperant, postquam rasi sunt.
JUDG|16|23|Principes autem Philisthinorum convenerunt in unum, ut immolarent hostias magnificas Dagon deo suo et epularentur dicentes: Tradidit deus nosterin manus nostrasinimicum nostrum Samson ".
JUDG|16|24|Quem etiam populus videns laudabat deum suum eademque dicebat: Tradidit deus noster in manus nostrasadversarium nostrum,qui vastavit terram nostramet occidit plurimos nostrum ".
JUDG|16|25|Cum enim iam hilariores essent, postulaverunt, ut vocaretur Samson et ante eos luderet. Qui adductus de carcere ludebat ante eos; feceruntque eum stare inter duas columnas.
JUDG|16|26|Qui dixit puero tenenti manum suam: " Dimitte me, ut tangam columnas, quibus imminet domus, et recliner super eas et paululum requiescam ".
JUDG|16|27|Domus autem plena erat virorum ac mulierum; et erant ibi omnes principes Philisthinorum, ac de tecto circiter tria milia utriusque sexus spectabant ludentem Samson.
JUDG|16|28|At ille invocavit Dominum dicens: " Domine Deus, memento mei! Et redde mihi tantum hac vice fortitudinem pristinam, Deus, ut ulciscar me de Philisthim saltem pro uno duorum luminum meorum! ".
JUDG|16|29|Et tangens ambas columnas medias, quibus innitebatur domus, obnixusque contra alteram earum dextera et contra alteram laeva
JUDG|16|30|ait: " Moriatur anima mea cum Philisthim! ". Concussisque fortiter columnis, cecidit domus super omnes principes et ceteram multitudinem, quae ibi erat; multoque plures interfecit moriens, quam ante vivus occiderat.
JUDG|16|31|Descendentes autem fratres eius et universa cognatio tulerunt corpus eius et sepelierunt inter Saraa et Esthaol in sepulcro patris sui Manue; iudicavitque Israel viginti annis.
JUDG|17|1|Fuit vir quidam de monte Ephraim nomine Michas,
JUDG|17|2|qui dixit matri suae: " Mille centum argenteos, qui ablati sunt a te et super quibus, me audiente, maledicens iuraveras, ecce ego habeo; ego abstuli ". Cui illa respondit: " Benedictus filius meus Domino! ".
JUDG|17|3|Reddidit ergo eos matri suae, quae dixit ei: " Consecravi et vovi argentum hoc Domino: de manu mea suscipiat pro filio meo, ut faciat sculptile atque conflatile. Et nunc trado illud tibi ".
JUDG|17|4|Reddiditque eos matri suae, quae tulit ducentos argenteos et dedit eos argentario, ut faceret ex eis sculptile atque conflatile, quod fuit in domo Michae,
JUDG|17|5|qui aediculam Dei habens fecit ephod ac theraphim implevitque unius filiorum suorum manum, et factus est ei sacerdos.
JUDG|17|6|In diebus illis non erat rex in Israel, sed unusquisque, quod sibi rectum videbatur, hoc faciebat.
JUDG|17|7|Fuit quoque adulescens de Bethlehem Iudae ex cognatione Iudae; eratque ipse Levites et habitabat ibi ut advena.
JUDG|17|8|Egressusque de civitate Bethlehem peregrinari voluit ubicumque sibi commodum repperisset. Cumque iter faciens venisset in monte Ephraim usque ad domum Michae,
JUDG|17|9|interrogatus est ab eo unde venisset. Qui respondit: " Levita sum de Bethlehem Iudae et vado, ut habitem, ubi potuero et utile mihi esse perspexero ".
JUDG|17|10|Dixitque Michas: " Mane apud me et esto mihi parens ac sacerdos; daboque tibi per annos singulos decem argenteos ac vestium apparatum et quae ad victum sunt necessaria ".
JUDG|17|11|Acquievit et mansit apud hominem fuitque illi quasi unus de filiis.
JUDG|17|12|Implevitque Michas manum eius et habuit puerum sacerdotem apud se,
JUDG|17|13|" nunc scio, dicens, quod benefaciet mihi Dominus habenti levitici generis sacerdotem ".
JUDG|18|1|In diebus illis non erat rex in Israel, et tribus Dan quaere bat possessionem sibi, ut habitaret in ea; usque ad illum enim diem inter ceteras tribus sortem non acceperat.
JUDG|18|2|Miserunt igitur filii Dan stirpis et familiae suae quinque viros fortissimos de Saraa et Esthaol, ut explorarent terram et diligenter inspicerent, dixeruntque eis: " Ite et considerate terram ". Qui cum venissent in montem Ephraim usque ad domum Michae, pernoctaverunt ibi.
JUDG|18|3|Cum essent prope domum Michae, agnoscentes vocem adulescentis Levitae declinaverant illuc dicentes ad eum: " Quis te huc adduxit? Quid hic agis? Quam ob causam huc venire voluisti? ".
JUDG|18|4|Qui respondit eis: " Haec et haec praestitit mihi Michas et me mercede conduxit, ut sim ei sacerdos ".
JUDG|18|5|Rogaveruntque eum, ut consuleret Deum, ut scire possent an prospero itinere pergerent, et res haberet effectum.
JUDG|18|6|Qui respondit eis: " Ite cum pace; Dominus respicit viam vestram et iter, quo pergitis ".
JUDG|18|7|Euntes itaque quinque viri venerunt Lais videruntque populum habitantem in ea absque ullo timore iuxta Sidoniorum consuetudinem, securum et quietum, nullo eis penitus resistente, magnarumque opum et procul a Sidoniis neque in societate cum Syria.
JUDG|18|8|Reversique ad fratres suos in Saraa et Esthaol et quid egissent sciscitantibus, responderunt:
JUDG|18|9|" Surgite, et ascendamus adversus eos. Vidimus enim terram valde opulentam et uberem, et vos neglegetis? Nolite cessare; eamus et possideamus eam.
JUDG|18|10|Intrabimus ad securos in regionem latissimam; tradetque nobis Deus locum, in quo nullius rei est penuria eorum, quae sunt in terra ".
JUDG|18|11|Profecti igitur sunt de cognatione Dan, de Saraa et Esthaol, sescenti viri accincti armis bellicis.
JUDG|18|12|Ascendentesque castrametati sunt in Cariathiarim Iudae, qui locus ex eo tempore Castrorum Dan nomen accepit et est post tergum Cariathiarim.
JUDG|18|13|Inde transierunt in montem Ephraim.Cumque venissent usque ad domum Michae,
JUDG|18|14|dixerunt quinque viri, qui prius missi fuerant ad considerandam terram Lais, fratribus suis: " Nostis quod in domibus istis sit ephod et theraphim et sculptile atque conflatile? Videte quid vobis placeat, ut faciatis ".
JUDG|18|15|Et, cum paululum declinassent, ingressi sunt domum adulescentis Levitae, domum Michae, salutaveruntque eum verbis pacificis.
JUDG|18|16|Sescenti autem viri, ita ut erant armati, stabant ante ostium.
JUDG|18|17|At illi, qui ingressi fuerant domum iuvenis, sculptile et ephod et theraphim atque conflatile tulerunt; et sacerdos stabat ante ostium et sescenti viri armati.
JUDG|18|18|Tulerunt igitur, qui intraverant domum, sculptile, ephod et theraphim atque conflatile. Quibus dixit sacerdos: " Quid facitis? ".
JUDG|18|19|Cui responderunt: " Tace et pone digitum super os tuum venique nobiscum, ut habeamus te patrem et sacerdotem. Quid tibi melius est, ut sis sacerdos in domo unius viri, an in una tribu et familia in Israel? ".
JUDG|18|20|Et gavisus est sacerdos tulitque ephod et theraphim ac sculptile et profectus est in medio populi.
JUDG|18|21|Qui cum pergerent et ante se ire fecissent parvulos et iumenta et omne, quod erat pretiosum,
JUDG|18|22|iamque a domo Michae essent procul, viri, qui habitabant in aedibus prope domum Michae, convocati secuti sunt filios Dan
JUDG|18|23|et post tergum clamare coeperunt. Qui cum respexissent, dixerunt ad Micham: " Quid tibi vis? Cur concurritis? ".
JUDG|18|24|Qui respondit: " Deos meos, quos mihi feci, tulistis, et sacerdotem et omnia, quae habeo, et dicitis: "Quid tibi est?" ".
JUDG|18|25|Dixeruntque ei filii Dan: " Cave, ne ultra loquaris ad nos, et irruant in te viri animo concitati, et ipse cum omni domo tua pereas ".
JUDG|18|26|Et sic, coepto itinere, perrexerunt. Videns autem Michas quod fortiores se essent, reversus est in domum suam.
JUDG|18|27|Sescenti autem viri tulerunt, quod Michas fecerat, et sacerdotem eius veneruntque in Lais ad populum quiescentem atque securum et percusserunt eos in ore gladii urbemque incendio tradiderunt,
JUDG|18|28|nullo penitus ferente praesidium, eo quod procul habitarent a Sidone neque cum Syria haberent quidquam societatis ac negotii.Erat autem civitas sita in regione Rohob; quam rursum exstruentes habitaverunt in ea,
JUDG|18|29|vocato nomine civitatis Dan iuxta vocabulum patris sui, quem genuerat Israel, quae prius Lais dicebatur.
JUDG|18|30|Posueruntque sibi sculptile; et Ionathan filius Gersam filii Moysi ac filii eius sacerdotes erant in tribu Dan usque ad diem captivitatis terrae;
JUDG|18|31|mansitque apud eos idolum Michae omni tempore, quo fuit domus Dei in Silo.
JUDG|18|32|In diebus illis non erat rex in Israel.
JUDG|19|1|Fuit quidam vir Levi tes habitans ut advena in extrema parte montis Ephraim, qui accepit concubinam de Bethlehem Iudae.
JUDG|19|2|Quae irritata reversa est in domum patris sui in Bethlehem mansitque apud eum quattuor mensibus.
JUDG|19|3|Secutusque est eam vir suus volens loqui ad cor eius et secum reducere habens in comitatu puerum et duos asinos. Quae suscepit eum et introduxit in domum patris sui. Quem cum socer eius vidisset, occurrit ei laetus
JUDG|19|4|et retinuit hominem. Mansitque gener in domo soceri tribus diebus comedens cum eo et bibens familiariter.
JUDG|19|5|Die autem quarto, cum de nocte consurrexissent, et ille proficisci vellet, socer ait ad eum: " Gusta prius pauxillum panis et conforta cor tuum et sic proficisceris ".
JUDG|19|6|Sederuntque ambo simul et comederunt ac biberunt. Dixitque pater puellae ad generum suum: " Quaeso te, ut hodie hic maneas, pariterque laetemur ".
JUDG|19|7|At ille consurgens coepit velle proficisci. Et nihilominus obnixe eum socer tenuit et apud se fecit manere.
JUDG|19|8|Mane autem facto, quinta die parabat Levites iter; cui socer rursum: " Oro te, inquit, ut confortes cor tuum". Et tardabant, donec declinaret dies; et ambo comederunt simul.
JUDG|19|9|Surrexitque adulescens, ut pergeret cum uxore sua et puero. Cui rursum locutus est socer eius pater puellae: " Considera quod dies ad occasum declivior sit et propinquet ad vesperum; manete apud me etiam hodie, pernocta hic et esto laeto animo, et cras mane proficiscemini, ut vadas in domum tuam ".
JUDG|19|10|Noluit gener acquiescere sermonibus eius, sed statim perrexit et venit contra Iebus, id est Ierusalem, ducens secum duos asinos onustos et concubinam.
JUDG|19|11|Iamque aderant iuxta Iebus, et dies mutabatur in noctem; dixitque puer ad dominum suum: " Veni, obsecro, declinemus ad urbem Iebusaeorum et maneamus in ea ".
JUDG|19|12|Cui respondit dominus: " Non ingrediamur oppidum gentis alienae, quae non est de filiis Israel, sed transibimus usque Gabaa ".
JUDG|19|13|Dixitque puero suo: "Veni, accedamus ad unum de locis et manebimus in Gabaa aut Rama ".
JUDG|19|14|Transierunt igitur Iebus et coeptum carpebant iter; occubuitque eis sol iuxta Gabaa, quae est in tribu Beniamin.
JUDG|19|15|Diverteruntque ad eam, ut manerent ibi; quo cum intrassent, sedebant in platea civitatis, et nullus eos recipere volebat hospitio.
JUDG|19|16|Et ecce apparuit homo senex revertens de agro et de opere suo vespere, qui et ipse erat de monte Ephraim et peregrinus habitabat in Gabaa; homines autem loci illius erant de tribu Beniamin.
JUDG|19|17|Elevatisque oculis, vidit senex sedentem hominem viatorem in platea civitatis et dixit ad eum: " Unde venis et quo vadis? ".
JUDG|19|18|Qui respondit ei: " Profecti sumus de Bethlehem Iudae et pergimus ad locum meum, qui est in extrema parte montis Ephraim, unde profectus sum in Bethlehem. Et nunc vado ad domum meam, nullusque sub tectum suum me vult recipere
JUDG|19|19|habentem paleas et pabulum pro asinis nostris et panem ac vinum in meos et ancillae tuae usus et pueri, qui cum servo tuo sunt; nulla re indigemus nisi hospitio ".
JUDG|19|20|Cui respondit senex: " Pax tecum sit! Ego praebebo omnia, quae necessaria sunt; tantum, quaeso, ne in platea maneas ".
JUDG|19|21|Introduxitque eum in domum suam et commixtum migma asinis praebuit; ac, postquam laverunt pedes suos, recepit eos in convivium.
JUDG|19|22|Illis laeto corde epulantibus, venerunt viri civitatis illius filii Belial et circumdantes domum senis fores pulsare coeperunt clamantes ad dominum domus atque dicentes: " Educ virum, qui ingressus est domum tuam, ut abutamur eo ".
JUDG|19|23|Egressusque est ad eos senex et ait: " Nolite, fratres, nolite facere malum hoc, quia ingressus est homo hospitium meum, et cessate ab hac stultitia.
JUDG|19|24|Habeo filiam virginem, et hic homo habet concubinam; educam eas ad vos, ut humilietis eas et faciatis eis, quod vobis placuerit; tantum, obsecro, ne scelus hoc operemini in virum ".
JUDG|19|25|Nolebant acquiescere sermonibus eius; quod cernens homo apprehendit et eduxit ad eos concubinam suam. Qua cum abusi essent et tota nocte ei illusissent, dimiserunt eam mane.
JUDG|19|26|At mulier, recedentibus tenebris, venit ad ostium domus, ubi manebat dominus suus, et ibi corruit.
JUDG|19|27|Mane facto surrexit homo et aperuit ostium, ut coeptam expleret viam; et ecce concubina eius iacebat ante ostium, sparsis in limine manibus.
JUDG|19|28|Cui ille loquebatur: " Surge, ut ambulemus ". Qua nihil respondente, intellegens quod erat mortua, tulit eam et imposuit asino; reversusque est in domum suam.
JUDG|19|29|Quam cum esset ingressus, arripuit gladium et cadaver uxoris secundum ossa sua in duodecim partes ac frusta concidens misit in omnes terminos Israel.
JUDG|19|30|Quod cum vidissent singuli, conclamabant: " Numquam res talis facta et visa est in Israel ex eo die, quo ascenderunt patres nostri de Aegypto, usque in praesens tempus! ". Praeceperat enim viris, quos miserat, dicens: Haec dicite omni viro Israel: Si factum est quidquam tale ex die, quo ascenderunt filii Israel de terra Aegypti, usque ad praesentem diem? Attendite ad hoc, consiliamini et decernite quid facto opus sit!".
JUDG|20|1|Egressi sunt itaque omnes fi lii Israel et pariter congrega ti, quasi vir unus, de Dan usque Bersabee et terra Galaad ad Dominum in Maspha.
JUDG|20|2|Omnisque populi anguli et cunctae tribus Israel in ecclesiam populi Dei convenerunt: quadringenta milia peditum pugnatorum.
JUDG|20|3|Nec latuit filios Beniamin, quod ascendissent filii Israel in Maspha. Interrogatusque Levita maritus mulieris interfectae quo modo tantum scelus perpetratum esset,
JUDG|20|4|respondit: " Veni in Gabaa Beniamin cum uxore mea illucque diverti.
JUDG|20|5|Et ecce homines civitatis illius circumdederunt nocte domum, in qua manebam, volentes me occidere et uxorem meam incredibili libidinis furore vexantes; denique mortua est.
JUDG|20|6|Quam arreptam in frusta concidi misique partes in omnes terminos possessionis Israel, quia fecerunt nefas et piaculum in Israel.
JUDG|20|7|Adestis omnes, filii Israel: decernite quid facere debeatis ".
JUDG|20|8|Stansque omnis populus quasi unius hominis sermone respondit: " Non recedemus in tabernacula nostra, nec suam quisquam intrabit domum,
JUDG|20|9|sed hoc contra Gabaa in commune faciemus secundum sortem:
JUDG|20|10|decem viri eligantur e centum ex omnibus tribubus Israel et centum de mille et mille de decem milibus, ut comportent exercitui cibaria illis, qui venerunt, ut reddant Gabaa Beniamin pro scelere, quod meretur ".
JUDG|20|11|Convenitque universus Israel ad civitatem quasi unus homo, eadem mente unoque consilio,
JUDG|20|12|et miserunt nuntios ad omnem tribum Beniamin, qui dicerent: " Quale nefas in vobis repertum est!
JUDG|20|13|Tradite homines filios Belial in Gabaa, qui hoc flagitium perpetrarunt, ut moriantur, et auferatur malum de Israel ".Qui noluerunt fratrum suorum filiorum Israel audire mandatum,
JUDG|20|14|sed ex cunctis urbibus, quae suae sortis erant, convenerunt in Gabaa, ut illis ferrent auxilium et contra universum Israel populum dimicarent.
JUDG|20|15|Recensitique sunt in die illa viginti sex milia de civitatibus Beniamin educentium gladium, praeter habitatores Gabaa, qui septingenti erant viri fortissimi.
JUDG|20|16|In universo hoc populo erant septingenti viri electi, qui sinistra pro dextra utebantur et sic fundis lapides ad certum iaciebant, ut capillum quoque possent percutere, et nequaquam in alteram partem ictus lapidis deferretur.
JUDG|20|17|Virorum quoque Israel, absque filiis Beniamin, recensita sunt quadringenta milia educentium gladios et paratorum ad pugnam.
JUDG|20|18|Qui surgentes venerunt in Bethel consulueruntque Deum atque dixerunt: " Quis erit in exercitu nostro princeps certaminis contra filios Beniamin?. Quibus respondit Dominus: " Iuda ascendet primus ".
JUDG|20|19|Statimque filii Israel surgentes mane castrametati sunt contra Gabaa;
JUDG|20|20|et inde procedentes ad pugnam contra Beniamin, contra urbem aciem direxerunt.
JUDG|20|21|Egressique filii Beniamin de Gabaa occiderunt de filiis Israel die illo viginti duo milia viros.
JUDG|20|22|Rursum filii Israel confortati in eodem loco, in quo prius certaverant, aciem direxerunt,
JUDG|20|23|ita tamen ut prius ascenderent et flerent coram Domino usque ad noctem consulerentque eum et dicerent: " Debeo ultra procedere ad dimicandum contra filios Beniamin fratres meos, an non? ". Quibus ille respondit: " Ascendite ad eos ".
JUDG|20|24|Cumque filii Israel altero die contra filios Beniamin ad proelium processissent,
JUDG|20|25|eruperunt filii Beniamin de Gabaa et occurrentes eis iterum decem et octo milia virorum educentium gladium prostraverunt.
JUDG|20|26|Quam ob rem omnes filii Israel, universus populus, venerunt in Bethel et sedentes flebant coram Domino ieiunaveruntque die illo usque ad vesperam et obtulerunt ei holocausta et pacificas victimas
JUDG|20|27|et super statu suo interrogaverunt. Eo tempore ibi erat arca foederis Dei,
JUDG|20|28|et Phinees filius Eleazari filii Aaron stabat coram eo. Consuluerunt igitur Dominum atque dixerunt: " Exire ultra debemus ad pugnam contra filios Beniamin fratres nostros, an quiescere? ". Quibus ait Dominus: " Ascendite, cras enim tradam eos in manus vestras ".
JUDG|20|29|Posueruntque filii Israel insidias per circuitum urbis Gabaa
JUDG|20|30|et tertia vice sicut semel et bis contra Beniamin et Gabaa exercitum produxerunt.
JUDG|20|31|Sed et filii Beniamin eruperunt in occursum populi et abstracti de civitate coeperunt caedere ex eis sicut primo et secundo die, per duas semitas terga vertentes, quarum una ferebat in Bethel, altera in Gabaa, atque prosternere in campo triginta circiter viros.
JUDG|20|32|Putaverunt enim solito eos more percussos cedere; qui fugam simulaverunt, ut abstraherent eos de civitate et quasi fugientes ad supradictas semitas perducerent.
JUDG|20|33|Omnes itaque viri Israel surgentes de sedibus suis tetenderunt aciem in loco, qui vocatur Baalthamar. Insidiae quoque eruperunt de loco suo, de regione in occidente Gabaa.
JUDG|20|34|Venerunt ergo adversus Gabaa decem milia virorum electorum de universo Israel. Ingravatumque est bellum contra filios Beniamin, et non intellexerunt quod ex omni parte illis instaret interitus.
JUDG|20|35|Percussitque eos Dominus in conspectu filiorum Israel, et interfecerunt ex eis in illo die viginti quinque milia et centum viros, omnes bellatores et educentes gladium.
JUDG|20|36|Filii autem Beniamin, cum se inferiores esse vidissent, coeperunt fugere. Quod cernentes filii Israel, dederunt eis ad fugiendum locum, quia confidebant in insidiis, quas iuxta urbem posuerant.
JUDG|20|37|Qui cum repente de latibulis surrexissent, irruerunt super Gabaa et ingressi celeriter percusserunt totam civitatem in ore gladii.
JUDG|20|38|Signum autem dederant filii Israel his, quos in insidiis collocaverant, ut ignem accenderent et, ascendente in altum fumo, captam urbem demonstrarent.
JUDG|20|39|Verterant ergo terga filii Israel in ipso certamine positi, et filii Beniamin putantes quod percussissent eos sicut in priore pugna, coeperant de exercitu eorum caedere triginta fere viros.
JUDG|20|40|Cum autem columna fumi de civitate conscendere coepisset, et Beniamin quoque retro aspiciens cerneret de civitate flammas in sublime ferri,
JUDG|20|41|cumque vir Israel versa facie aggrederetur, vir Beniamin conturbatus est, quia vidit se apprehensum a malo.
JUDG|20|42|Et ad viam deserti ire coeperunt, illuc quoque eos adversariis persequentibus. Sed et hi, qui urbem succenderant, occurrerunt eis,
JUDG|20|43|atque ita factum est ut ex utraque parte ab hostibus caederentur, nec erat eis ulla requies. Prostrati sunt usque ad orientalem plagam urbis Gabaa.
JUDG|20|44|Fuerunt autem, qui interfecti sunt de Beniamin, decem et octo milia virorum omnes robustissimi pugnatores.
JUDG|20|45|Qui remanserant, fugerunt in solitudinem et pergebant ad petram, cuius vocabulum est Remmon. Quasi racemos colligentes occiderunt in viis quinque milia viros. Et cum instantius eos persequerentur usque Gadaam, interfecerunt etiam alios duo milia.
JUDG|20|46|Et sic factum est ut omnes, qui ceciderant de Beniamin in die illa, essent viginti quinque milia pugnatores ad bella promptissimi.
JUDG|20|47|Remanserunt itaque, qui evadere potuerant et fugere in solitudinem, sescenti viri; sederuntque in petra Remmon mensibus quattuor.
JUDG|20|48|Regressi autem filii Israel ex civitatibus a viris usque ad iumenta, usque ad omne, quod inveniri poterat, gladio percusserunt, cunctasque urbes et viculos Beniamin vorax flamma consumpsit.
JUDG|21|1|Iuraverunt autem filii Israel in Maspha et dixerunt: " Nullus nostrum dabit filiis Beniamin de filiabus suis uxorem ".
JUDG|21|2|Venitque populus in Bethel, et in conspectu Dei sedentes usque ad vesperam levaverunt vocem et magno ululatu coeperunt flere dicentes:
JUDG|21|3|" Quare, Domine, Deus Israel, factum est hoc in populo tuo, ut hodie una tribus auferretur de Israel? ".
JUDG|21|4|Altera autem die diluculo consurgentes exstruxerunt altare obtuleruntque ibi holocausta et pacificas victimas
JUDG|21|5|et dixerunt: " Quis non ascendit in congregationem ad Dominum de universis tribubus Israel? ". Grandi enim se iuramento constrinxerant interfici eos, qui non ascendissent ad Dominum in Maspha.
JUDG|21|6|Ductique paenitentia filii Israel super fratre suo Beniamin coeperunt dicere: " Ablata est hodie una tribus de Israel.
JUDG|21|7|Quid faciemus, ut, qui remanserunt, uxores accipiant? Omnes enim in commune iuravimus per Dominum non daturos nos his filias nostras ".
JUDG|21|8|Idcirco dixerunt: " Quis est de universis tribubus Israel, qui non ascendit ad Dominum in Maspha? ". Et ecce nemo de Iabes Galaad in castra venerat ad congregationem,
JUDG|21|9|et, cum populus recenseretur, nullus ex eis repertus est.
JUDG|21|10|Misit itaque coetus decem milia viros robustissimos et praeceperunt eis: " Ite et percutite habitatores Iabes Galaad in ore gladii tam uxores quam parvulos eorum.
JUDG|21|11|Et hoc erit, quod observare debetis: Omne generis masculini et mulieres, quae cognoverunt viros, interficite; virgines autem reservate ".
JUDG|21|12|Inventaeque sunt de Iabes Galaad quadringentae virgines, quae nescierunt viri torum, et adduxerunt eas in castra in Silo in terra Chanaan.
JUDG|21|13|Misitque coetus nuntios ad filios Beniamin, qui erant in petra Remmon, et dederunt eis pacem.
JUDG|21|14|Veneruntque filii Beniamin in illo tempore, et datae sunt eis uxores de filiabus Iabes Galaad; alias autem non reppererunt, quas simili modo traderent.
JUDG|21|15|Populusque valde doluit de Beniamin, quia fecerat Dominus confractionem in tribubus Israel.
JUDG|21|16|Dixeruntque seniores coetus: " Quid faciemus reliquis, qui non acceperunt uxores? Omnes in Beniamin feminae conciderunt ".
JUDG|21|17|Et dixerunt: " Possessio eorum, qui effugerunt, erit Beniamin, ne una tribus deleatur ex Israel.
JUDG|21|18|Filias autem nostras eis dare non possumus, constricti hoc iuramento: Maledictus, qui dederit de filiabus suis uxorem Beniamin!" ".
JUDG|21|19|Ceperuntque consilium atque dixerunt: " Ecce sollemnitas Domini est in Silo anniversaria, quae sita est ad septentrionem urbis Bethel et ad orientalem plagam viae, quae de Bethel tendit ad Sichimam et ad meridiem oppidi Lebona ".
JUDG|21|20|Praeceperuntque filiis Beniamin atque dixerunt: "Ite et latitate in vineis;
JUDG|21|21|cumque videritis filias Silo ad ducendos choros ex more procedere, exite repente de vineis et rapite ex eis singuli uxores singulas et pergite in terram Beniamin ".
JUDG|21|22|Cumque venerint patres earum ac fratres et apud nos queri coeperint, dicemus eis: " Miseremini nostri et eorum; non enim acceperunt unusquisque uxorem in bello, et vos, si dedissetis eis, deliquissetis ".
JUDG|21|23|Feceruntque filii Beniamin, ut sibi fuerat imperatum, et iuxta numerum suum rapuerunt sibi de his, quae ducebant choros, uxores singulas; abieruntque in possessionem suam aedificantes urbes et habitantes in eis.
JUDG|21|24|Filii quoque Israel reversi sunt inde illo tempore unusquisque ad tribum et familiam suam in possessionem suam.
JUDG|21|25|In diebus illis non erat rex in Israel, sed unusquisque, quod sibi rectum videbatur, hoc faciebat.
RUTH|1|1|In diebus, quando iudices praeerant, facta est fames in ter ra. Abiitque homo de Bethlehem Iudae, ut peregrinaretur in regione Moabitide cum uxore sua ac duobus liberis.
RUTH|1|2|Ipse vocabatur Elimelech et uxor eius Noemi et duo filii alter Mahalon et alter Chelion Ephrathaei de Bethlehem Iudae. Ingressique regionem Moabitidem morabantur ibi.
RUTH|1|3|Et mortuus est Elimelech maritus Noemi, remansitque ipsa cum filiis,
RUTH|1|4|qui acceperunt uxores Moabitidas, quarum una vocabatur Orpha, altera Ruth; manseruntque ibi decem fere annis.
RUTH|1|5|Et ambo mortui sunt, Mahalon videlicet et Chelion; remansitque mulier orbata duobus liberis ac marito.
RUTH|1|6|Et surrexit, ut in patriam pergeret cum utraque nuru sua de regione Moabitide; audierat enim quod respexisset Dominus populum suum et dedisset eis escas.
RUTH|1|7|Egressa est itaque de loco peregrinationis suae cum utraque nuru et, iam in via posita revertendi in terram Iudae,
RUTH|1|8|dixit ad eas: " Ite in domum matris vestrae; faciat Dominus vobiscum misericordiam, sicut fecistis cum mortuis et mecum:
RUTH|1|9|det vobis invenire requiem in domibus virorum, quos sortiturae estis ". Et osculata est eas. Quae elevata voce flere coeperunt
RUTH|1|10|et dicere: " Tecum pergemus ad populum tuum ".
RUTH|1|11|Quibus illa respondit: " Revertimini, filiae meae; cur venitis mecum? Num ultra habeo filios in utero meo, ut viros ex me sperare possitis?
RUTH|1|12|Revertimini, filiae meae, abite; iam enim senectute confecta sum nec apta vinculo coniugali; etiamsi possem hac nocte concipere et parere filios,
RUTH|1|13|numquid exspectare velitis et abstinere vos a matrimonio, donec crescant et annos impleant pubertatis? Nolite, quaeso, filiae meae; quia amaritudo est mihi magis quam vobis, et egressa est manus Domini contra me.
RUTH|1|14|Elevata igitur voce, rursum flere coeperunt. Orpha osculata socrum est ac reversa; Ruth autem adhaesit socrui suae.
RUTH|1|15|Cui dixit Noemi: " En reversa est cognata tua ad populum suum et ad deos suos; vade cum ea".
RUTH|1|16|Quae respondit: "Noli instare mihi, ut relinquam te et abeam; quocumque perrexeris, pergam; ubi morata fueris, et ego pariter morabor: populus tuus populus meus et Deus tuus Deus meus.
RUTH|1|17|Quae te morientem terra susceperit, in ea moriar ibique locum accipiam sepulturae. Haec mihi faciat Dominus et haec addat, si non sola mors me et te separaverit ".
RUTH|1|18|Videns ergo Noemi quod obstinato Ruth animo decrevisset secum pergere, adversari noluit nec ultra ad suos reditum persuadere.
RUTH|1|19|Profectaeque sunt simul et venerunt in Bethlehem. Quibus urbem ingressis, tota urbs commota est super eas; dicebantque mulieres: "Haec est illa Noemi!".
RUTH|1|20|Quibus ait: "Ne vocetis me Noemi (id est Pulchram), sed vocate me Mara hoc est Amaram), quia valde me amaritudine replevit Omnipotens.
RUTH|1|21|Egressa sum plena, et vacuam reduxit me Dominus; cur igitur vocatis me Noemi, quam humiliavit Dominus, et afflixit Omnipotens? ".
RUTH|1|22|Venit ergo Noemi cum Ruth Moabitide nuru sua de terra peregrinationis suae ac reversa est in Bethlehem, quando hordea metere incipiebant.
RUTH|2|1|Erat autem Noemi consangui neus viri sui homo potens et for tis nomine Booz.
RUTH|2|2|Dixitque Ruth Moabitis ad socrum suam: " Si permittis, vadam in agrum et colligam spicas, quae fugerint manus metentium, ubicumque clementis in me patris familias repperero gratiam". Cui illa respondit: " Vade, filia mea.
RUTH|2|3|Abiit itaque et colligebat spicas post terga metentium. Accidit autem ut ager ille haberet dominum nomine Booz, qui erat de cognatione Elimelech.
RUTH|2|4|Et ecce ipse veniebat de Bethlehem dixitque messoribus: "Dominus vobiscum". Qui responderunt ei: " Benedicat tibi Dominus ".
RUTH|2|5|Dixitque Booz iuveni, qui messoribus praeerat: " Cuius est haec puella?.
RUTH|2|6|Qui respondit: " Haec est Moabitis, quae venit cum Noemi de regione Moabitide
RUTH|2|7|et rogavit, ut spicas colligeret remanentes sequens messorum vestigia; et de mane usque nunc stat in agro et nunc tantum ad momentum requievit ".
RUTH|2|8|Et ait Booz ad Ruth: " Audi, filia: ne vadas ad colligendum in alterum agrum nec recedas ab hoc loco, sed iungere puellis meis.
RUTH|2|9|Vide et, ubi messuerint, sequere eas; mandavi enim pueris, ut nemo tibi molestus sit; sed, si sitieris, vade ad sarcinulas et bibe de aqua, quam pueri hauserint ".
RUTH|2|10|Quae cadens in faciem suam et adorans super terram dixit ad eum: " Unde mihi hoc, ut invenirem gratiam ante oculos tuos, et nosse me dignareris peregrinam mulierem? ".
RUTH|2|11|Cui ille respondit: " Nuntiata sunt mihi omnia, quae feceris socrui tuae post mortem viri tui et quod dereliqueris parentes tuos et terram, in qua nata es, et veneris ad populum, quem ante nesciebas.
RUTH|2|12|Reddat tibi Dominus pro opere tuo, et plenam mercedem recipias a Domino, Deo Israel, ad quem venisti et sub cuius confugisti alas ".
RUTH|2|13|Quae ait: " Inveniam gratiam ante oculos tuos, domine mi, qui consolatus es me et locutus es ad cor ancillae tuae, quae non sum similis unius puellarum tuarum ".
RUTH|2|14|Dixitque ad eam Booz hora vescendi: "Veni huc et comede panem et intinge buccellam tuam in aceto ". Sedit itaque ad messorum latus, et porrexit ei polentam, comeditque et saturata est et tulit reliquias.
RUTH|2|15|Atque inde surrexit, ut spicas ex more colligeret. Praecepit autem Booz pueris suis dicens: "Etiam inter manipulos colligat, ne prohibeatis eam;
RUTH|2|16|quin et de fasciculis spicas proicite et remanere permittite, ut colligat, et colligentem nemo corripiat ".
RUTH|2|17|Collegit ergo in agro usque ad vesperam; et, quae collegerat virga excutiens, invenit hordei quasi ephi mensuram (id est tres modios).
RUTH|2|18|Quos portans reversa est in civitatem et ostendit socrui suae, quae collegerat; insuper protulit et dedit ei de reliquiis cibi sui, quo saturata fuerat.
RUTH|2|19|Dixitque ei socrus: " Ubi hodie collegisti et ubi fecisti opus? Sit benedictus, qui misertus est tui! ". Indicavitque ei apud quem esset operata et dixit: " Nomen viri est Booz ".
RUTH|2|20|Cui respondit Noemi: " Benedictus sit a Domino, quia non subtraxit gratiam suam nec vivis nec mortuis! ". Rursumque ait: " Propinquus noster est homo ex eis, qui pro nobis ius redemptionis habent ".
RUTH|2|21|Et Ruth: " Hoc quoque, inquit, praecepit mihi, ut tamdiu messoribus eius iungerer, donec omnes segetes meterentur ".
RUTH|2|22|Cui dixit socrus: " Melius est, filia mea, ut cum puellis eius exeas ad metendum, ne in alieno agro quispiam tibi molestus sit ".
RUTH|2|23|Iuncta est itaque puellis Booz usque ad finem messis hordei et tritici; et mansit cum socru sua.
RUTH|3|1|Et dixit ad eam Noemi socrus sua: " Filia mea, quaeram tibi requiem et providebo, ut bene sit tibi.
RUTH|3|2|Booz propinquus noster, cuius puellis in agro iuncta eras, ecce ipse hac nocte aream hordei ventilat.
RUTH|3|3|Lavare igitur, ungere et induere pallio tuo ac descende in aream; non te videat homo, donec esum potumque finierit.
RUTH|3|4|Quando autem ierit ad dormiendum, nota locum, in quo dormiat; veniesque et discooperies pallium, quo operitur a parte pedum, et ibi iacebis. Ipse autem dicet tibi quid agere debeas ".
RUTH|3|5|Quae respondit: " Quidquid praeceperis, faciam ".
RUTH|3|6|Descenditque in aream et fecit omnia, quae sibi imperaverat socrus.
RUTH|3|7|Cumque comedisset Booz et bibisset et factus esset hilarior issetque ad dormiendum in extrema parte acervi manipulorum, venit abscondite et, discooperto a pedibus eius pallio, se proiecit.
RUTH|3|8|Et ecce, nocte iam media, expavit homo et erexit se viditque mulierem iacentem ad pedes suos.
RUTH|3|9|Et ait illi: " Quae es? ". Illaque respondit: " Ego sum Ruth ancilla tua. Expande pallium tuum super famulam tuam, quia tibi est ius redemptionis ".
RUTH|3|10|Et ille: " Benedicta, inquit, es a Domino, filia; et priorem pietatem posteriore superasti, quia non es secuta iuvenes pauperes sive divites.
RUTH|3|11|Noli ergo metuere, sed, quidquid dixeris mihi, faciam tibi; scit enim omnis populus, qui habitat intra portas urbis meae, mulierem te esse fortem.
RUTH|3|12|Nec abnuo me propinquum, sed est alius me propinquior.
RUTH|3|13|Quiesce hac nocte et, facto mane, si te voluerit propinquitatis iure suscipere, bene, suscipiat; sin autem ille noluerit, vivit Dominus, ego te absque ulla dubitatione suscipiam! Dormi usque mane ".
RUTH|3|14|Dormivit itaque ad pedes eius usque ad noctis abscessum. Surrexitque, antequam homines se cognoscerent mutuo, et dixit Booz: " Cave, ne quis noverit quod huc veneris ".
RUTH|3|15|Et rursum: " Expande, inquit, palliolum tuum, quo operiris, et tene utraque manu ". Qua extendente et tenente, mensus est sex modios hordei et posuit super eam; quae portans ingressa est civitatem
RUTH|3|16|et venit ad socrum suam. Quae dixit ei: " Quid egisti, filia? ". Narravitque ei omnia, quae sibi fecisset homo,
RUTH|3|17|et ait: " Ecce sex modios hordei dedit mihi et ait: " Nolo vacuam te reverti ad socrum tuam ".
RUTH|3|18|Dixitque Noemi: " Exspecta, filia, donec videamus quem res exitum habeat; neque enim cessabit homo, nisi compleverit hodie, quod locutus est.
RUTH|4|1|Ascendit ergo Booz ad portam et sedit ibi. Cumque vidisset propinquum praeterire, de quo locutus erat, dixit ad eum: " Declina paulisper et sede hic ", vocans eum nomine suo. Qui divertit et sedit.
RUTH|4|2|Tollens autem Booz decem viros de senioribus civitatis dixit ad eos: " Sedete hic ".
RUTH|4|3|Quibus sedentibus, locutus est ad propinquum: " Partem agri fratris nostri Elimelech vendit Noemi, quae reversa est de regione Moabitide.
RUTH|4|4|Quod audire te volui et tibi dicere: Coram cunctis sedentibus et maioribus natu de populo meo, si vis possidere iure propinquitatis, eme et posside; sin autem tibi displicet, hoc ipsum indica mihi, ut sciam quid facere debeam. Nullus est enim propinquus, excepto te, qui prior es, et me, qui secundus sum ". At ille respondit: " Ego agrum emam ".
RUTH|4|5|Cui dixit Booz: " Quando emeris agrum de manu Noemi, Ruth quoque Moabitidem, quae uxor defuncti fuit, debes accipere, ut suscites nomen defuncti propinqui tui in hereditate sua ".
RUTH|4|6|Qui respondit: " Cedo iure propinquitatis; neque enim possessionem familiae meae delere debeo. Tu meo utere privilegio, quo me libenter carere profiteor ".
RUTH|4|7|Hic autem erat mos antiquitus in Israel pro redemptione et commutatione: ut esset firma concessio, solvebat homo calceamentum suum et dabat proximo suo. Hoc erat testimonium cessionis in Israel.
RUTH|4|8|Dixit ergo propinquus ad Booz: " Eme tibi ". Et solvit calceamentum suum de pede suo.
RUTH|4|9|Et Booz maioribus natu et universo populo: " Testes, inquit, vos estis hodie quod acquisierim omnia, quae fuerunt Elimelech et Chelion et Mahalon, tradente Noemi,
RUTH|4|10|et etiam Ruth Moabitidem uxorem Mahalon in coniugium sumpserim, ut suscitem nomen defuncti in hereditate sua, ne vocabulum eius de fratribus suis et de porta loci sui deleatur. Vos, inquam, huius rei hodie testes estis ".
RUTH|4|11|Respondit omnis populus, qui erat in porta, et maiores natu: " Nos testes sumus; faciat Dominus hanc mulierem, quae ingreditur domum tuam, sicut Rachel et Liam, quae aedificaverunt ambae domum Israel.Fortiter age in Ephrathaet fac tibi celebre nomen in Bethlehem!
RUTH|4|12|Fiatque domus tua sicut domus Phares, quem Thamar peperit Iudae, de semine, quod dederit Dominus tibi ex hac puella! ".
RUTH|4|13|Tulit itaque Booz Ruth et accepit uxorem; ingressusque est ad eam, et dedit illi Dominus, ut conciperet et pareret filium.
RUTH|4|14|Dixeruntque mulieres ad Noemi: " Benedictus Dominus, qui non est passus, ut deficeret tibi hodie, qui redimit familiam tuam, et vocetur nomen eius in Israel
RUTH|4|15|et consoletur animam tuam et enutriat senectutem; de nuru enim tua natus est, quae te diligit et multo tibi est melior quam septem filii ".
RUTH|4|16|Susceptumque Noemi puerum posuit in sinu suo et gerulae officio fungebatur.
RUTH|4|17|Vicinae autem mulieres congratulantes ei et dicentes: " Natus est filius Noemi! ", vocaverunt nomen eius Obed. Hic est pater Isai patris David.
RUTH|4|18|Hae sunt generationes Phares: Phares genuit Esrom,
RUTH|4|19|Esrom genuit Aram, Aram genuit Aminadab,
RUTH|4|20|Aminadab genuit Naasson, Naasson genuit Salmon,
RUTH|4|21|Salmon genuit Booz, Booz genuit Obed,
RUTH|4|22|Obed genuit Iesse, Iesse genuit David.
1SAM|1|1|Fuit vir unus de Ramathaim Suphita de monte Ephraim, et nomen eius Elcana filius Ieroham filii Eliu filii Thohu filii Suph, Ephrathaeus.
1SAM|1|2|Et habuit duas uxores: nomen uni Anna et nomen secundae Phenenna. Fueruntque Phenennae filii, Annae autem non erant liberi.
1SAM|1|3|Et ascendebat vir ille de civitate sua singulis annis, ut adoraret et sacrificaret Domino exercituum in Silo. Erant autem ibi duo filii Heli, Ophni et Phinees, sacerdotes Domini.
1SAM|1|4|Venit ergo dies, et immolavit Elcana dabatque Phenennae uxori suae et cunctis filiis eius et filiabus partes;
1SAM|1|5|Annae autem dabat unam partem electam, quia Annam diligebat; Dominus autem concluserat vulvam eius.
1SAM|1|6|Affligebat quoque eam aemula eius et vehementer angebat, ut conturbaret eam, quod conclusisset Dominus vulvam eius.
1SAM|1|7|Sicque faciebat per singulos annos, cum, redeunte tempore, ascenderent templum Domini, et sic provocabat eam. Porro illa flebat et non capiebat cibum.
1SAM|1|8|Dixit ergo ei Elcana vir suus: " Anna, cur fles et quare non comedis? Et quam ob rem affligitur cor tuum? Numquid non ego melior sum tibi quam decem filii? ".
1SAM|1|9|Surrexit autem Anna, postquam comederant et biberant in Silo, et Heli sacerdote sedente super sellam ante postes templi Domini.
1SAM|1|10|Cum esset Anna amaro animo, oravit Dominum flens largiter
1SAM|1|11|et votum vovit dicens: " Domine exercituum, si respiciens videris afflictionem famulae tuae et recordatus mei fueris nec oblitus ancillae tuae dederisque servae tuae sexum virilem, dabo eum Domino omnes dies vitae eius, et novacula non ascendet super caput eius ".
1SAM|1|12|Factum est ergo, cum illa multiplicaret preces coram Domino, ut Heli observaret os eius.
1SAM|1|13|Porro Anna loquebatur in corde suo; tantumque labia illius movebantur, et vox penitus non audiebatur. Aestimavit igitur eam Heli temulentam
1SAM|1|14|dixitque ei: " Usquequo ebria eris? Digere paulisper vinum, quo mades!.
1SAM|1|15|Respondens Anna: " Nequaquam, inquit, domine mi; nam mulier infelix nimis ego sum: vinumque et omne, quod inebriare potest, non bibi, sed effudi animam meam in conspectu Domini.
1SAM|1|16|Ne reputes ancillam tuam quasi unam de filiabus Belial, quia ex multitudine doloris et maeroris mei locuta sum usque in praesens ".
1SAM|1|17|Tunc Heli ait ei: " Vade in pace, et Deus Israel det tibi petitionem, quam rogasti eum ".
1SAM|1|18|Et illa dixit: " Utinam inveniat ancilla tua gratiam in oculis tuis ". Et abiit mulier in viam suam et comedit; vultusque illius non fuerunt amplius sicut prius.
1SAM|1|19|Et surrexerunt mane et adoraverunt coram Domino.Reversique sunt et venerunt in domum suam in Rama. Cognovit autem Elcana Annam uxorem suam, et recordatus est eius Dominus.
1SAM|1|20|Et factum est post circulum dierum concepit Anna et peperit filium vocavitque nomen eius Samuel, eo quod a Domino postulasset eum.
1SAM|1|21|Ascendit autem vir Elcana et omnis domus eius, ut immolaret Domino hostiam annuam et votum suum.
1SAM|1|22|Et Anna non ascendit; dixit enim viro suo: " Non vadam, donec ablactetur infans, et ducam eum, et appareat ante conspectum Domini et maneat ibi iugiter ".
1SAM|1|23|Et ait ei Elcana vir suus: " Fac, quod bonum tibi videtur, et mane, donec ablactes eum; precorque, ut impleat Dominus verbum suum ". Mansit ergo mulier et lactavit filium suum, donec amoveret eum a lacte.
1SAM|1|24|Et adduxit eum secum, postquam ablactaverat, cum vitulo trium annorum et tribus modiis farinae et utre vini; et adduxit eum ad domum Domini in Silo. Puer autem erat adhuc infantulus.
1SAM|1|25|Et immolaverunt vitulum et obtulerunt puerum Heli,
1SAM|1|26|et ait Anna: " Obsecro, mi domine; vivit anima tua, domine, ego sum illa mulier, quae steti coram te hic orans Dominum.
1SAM|1|27|Pro puero isto oravi, et dedit mihi Dominus petitionem meam, quam postulavi eum.
1SAM|1|28|Idcirco et ego commodavi eum Domino; cunctis diebus, quibus vivet, postulatus erit pro Domino ".Et adoraverunt ibi Dominum.
1SAM|2|1|Et oravit Anna et ait: Exsultavit cor meum in Do mino,exaltatum est cornu meum in Deo meo;dilatatum est os meum super inimicos meos,quoniam laetata sum in salutari tuo.
1SAM|2|2|Non est sanctus ut est Dominus;neque enim est alius extra te,et non est fortis sicut Deus noster.
1SAM|2|3|Nolite multiplicare loqui sublimia gloriantes.Recedant superba de ore vestro,quia Deus scientiarum Dominus est, et ab eo ponderantur actiones.
1SAM|2|4|Arcus fortium confractus est,et infirmi accincti sunt robore.
1SAM|2|5|Saturati prius pro pane se locaverunt,et famelici non eguerunt amplius.Sterilis peperit plurimos,et, quae multos habebat filios, emarcuit.
1SAM|2|6|Dominus mortificat et vivificat,deducit ad infernum et reducit.
1SAM|2|7|Dominus pauperem facit et ditat,humiliat et sublevat;
1SAM|2|8|suscitat de pulvere egenumet de stercore elevat pauperem,ut sedeat cum principibuset solium gloriae teneat.Domini enim sunt cardines terrae, et posuit super eos orbem.
1SAM|2|9|Pedes sanctorum suorum servabit,et impii in tenebris conticescent,quia non in fortitudine sua roborabitur vir.
1SAM|2|10|Dominus conteret adversarios suos;super ipsos in caelis tonabit.Dominus iudicabit fines terraeet dabit imperium regi suoet sublimabit cornu christi sui ".
1SAM|2|11|Et abiit Elcana in Rama in domum suam. Puer autem erat minister in conspectu Domini ante faciem Heli sacerdotis.
1SAM|2|12|Porro filii Heli filii Belial nescientes Dominum
1SAM|2|13|neque officium sacerdotum ad populum, sed, quicumque immolasset victimam, veniebat puer sacerdotis, dum coquerentur carnes, et habebat fuscinulam tridentem in manu sua
1SAM|2|14|et mittebat eam in lebetem vel in caldariam aut in ollam sive in cacabum et omne, quod levabat fuscinula, tollebat sacerdos sibi. Sic faciebant universo Israeli venienti in Silo.
1SAM|2|15|Etiam, antequam adolerent adipem, veniebat puer sacerdotis et dicebat immolanti: " Da mihi carnem, ut coquam sacerdoti; non enim accipiet a te carnem coctam sed crudam ".
1SAM|2|16|Dicebatque illi immolans: " Incendatur primum iuxta morem hodie adeps, et tolle tibi, quantumcumque desiderat anima tua ". Qui respondens aiebat ei: " Nequaquam; nunc enim dabis, alioquin tollam vi ".
1SAM|2|17|Erat ergo peccatum puerorum grande nimis coram Domino, quia detrahebant sacrificio Domini.
1SAM|2|18|Samuel autem ministrabat ante faciem Domini, puer accinctus ephod lineo.
1SAM|2|19|Et tunicam parvam faciebat ei mater sua, quam afferebat ei singulis annis ascendens cum viro suo, ut immolaret hostiam annuam.
1SAM|2|20|Et benedicebat Heli Elcanae et uxori eius dicebatque: " Reddat tibi Dominus semen de muliere hac pro petitione, quae postulata est pro Domino. Et abierunt in locum suum.
1SAM|2|21|Visitavit ergo Dominus Annam, et concepit et peperit tres filios et duas filias. Et crevit puer Samuel apud Dominum.
1SAM|2|22|Heli autem erat senex valde et audivit omnia, quae faciebant filii sui universo Israeli et quomodo dormiebant cum mulieribus, quae ministrabant ad ostium tabernaculi,
1SAM|2|23|et dixit eis: " Quare facitis res huiuscemodi, quas ego audio, res pessimas, ab omni populo?
1SAM|2|24|Nolite, filii mei; non enim est bona fama, quam ego audio, ut transgredi faciatis populum Domini.
1SAM|2|25|Si peccaverit vir in virum,arbiter ei potest esse Deus;si autem in Dominum peccaverit vir,quis intercedet pro eo? ".Et non audierunt vocem patris sui, quia voluit Dominus occidere eos.
1SAM|2|26|Puer autem Samuel proficiebat atque crescebat et placebat tam Domino quam hominibus.
1SAM|2|27|Venit autem vir Dei ad Heli et ait ad eum: " Haec dicit Dominus: Numquid non aperte revelatus sum domui patris tui, cum esset in Aegypto in domo pharaonis?
1SAM|2|28|Et elegi eum ex omnibus tribubus Israel mihi in sacerdotem, ut ascenderet ad altare meum et adoleret mihi incensum et portaret ephod coram me; et dedi domui patris tui omnia de sacrificiis filiorum Israel.
1SAM|2|29|Quare calce abicitis victimam meam et munera mea, quae praecepi, ut offerrentur in templo, et magis honorasti filios tuos quam me, ut impinguaremini primitiis omnis sacrificii Israel populi mei?
1SAM|2|30|Propterea ait Dominus, Deus Israel: Loquens locutus sum, ut domus tua et domus patris tui ministraret in conspectu meo usque in sempiternum. Nunc autem, dicit Dominus, absit hoc a me. Sed quicumque glorificaverit me, glorificabo eum; qui autem contemnunt me, erunt ignobiles.
1SAM|2|31|Ecce dies veniunt, et praecidam brachium tuum et brachium domus patris tui, ut non sit senex in domo tua.
1SAM|2|32|Et videbis aemulum tuum in templo in universis prosperis Israel; et non erit senex in domo tua omnibus diebus.
1SAM|2|33|Verumtamen non auferam penitus virum ex te ab altari meo; sed ut deficiant oculi tui, et tabescat anima tua, et pars magna domus tuae morietur, cum ad virilem aetatem venerit.
1SAM|2|34|Hoc autem erit tibi signum, quod venturum est duobus filiis tuis Ophni et Phinees: in die uno morientur ambo.
1SAM|2|35|Et suscitabo mihi sacerdotem fidelem, qui iuxta cor meum et animam meam faciat; et aedificabo ei domum fidelem, et ambulabit coram christo meo cunctis diebus.
1SAM|2|36|Futurum est autem ut quicumque remanserit in domo tua, veniat, ut procidat ante illum pro nummo argenteo et torta panis dicatque: "Dimitte me, obsecro, ad unam partem sacerdotalem, ut comedam buccellam panis" ".
1SAM|3|1|Puer autem Samuel ministrabat Domino coram Heli. Et sermo Domini erat pretiosus in diebus illis: non erat visio frequens.
1SAM|3|2|Factum est ergo in die quadam, Heli iacebat in loco suo, et oculi eius caligaverant, nec poterat videre.
1SAM|3|3|Lucerna Dei nondum exstincta erat, et Samuel dormiebat in templo Domini, ubi erat arca Dei.
1SAM|3|4|Et vocavit Dominus Samuel, qui respondens ait: " Ecce ego ".
1SAM|3|5|Et cucurrit ad Heli et dixit: " Ecce ego; vocasti enim me ". Qui dixit: Non vocavi. Revertere; dormi! ". Et abiit et dormivit.
1SAM|3|6|Et Dominus rursum vocavit Samuel. Consurgensque Samuel abiit ad Heli et dixit: " Ecce ego, quia vocasti me ". Qui respondit: " Non vocavi te, fili mi. Revertere et dormi! ".
1SAM|3|7|Porro Samuel necdum sciebat Dominum, neque revelatus fuerat ei sermo Domini.
1SAM|3|8|Et Dominus rursum vocavit Samuel tertio, qui consurgens abiit ad Heli
1SAM|3|9|et ait: " Ecce ego, quia vocasti me ". Intellexit igitur Heli quia Dominus vocaret puerum, et ait ad Samuel: " Vade et dormi; et, si deinceps vocaverit te, dices: " Loquere, Domine, quia audit servus tuus" ". Abiit ergo Samuel et dormivit in loco suo.
1SAM|3|10|Et venit Dominus et stetit et vocavit, sicut vocaverat prius: " Samuel, Samuel ". Et ait Samuel: " Loquere, quia audit servus tuus ".
1SAM|3|11|Et dixit Dominus ad Samuel: " Ecce ego facio verbum in Israel, quod quicumque audierit, tinnient ambae aures eius.
1SAM|3|12|In die illo suscitabo adversum Heli omnia, quae locutus sum super domum eius: incipiam et complebo.
1SAM|3|13|Praedixi enim ei quod iudicaturus essem domum eius in aeternum propter iniquitatem, eo quod noverat filios suos contemnere Deum et non corripuit eos.
1SAM|3|14|Idcirco iuravi domui Heli quod non expietur iniquitas domus eius victimis et muneribus usque in aeternum ".
1SAM|3|15|Dormivit autem Samuel usque mane aperuitque ostia domus Domini. Et Samuel timebat indicare visionem Heli.
1SAM|3|16|Vocavit ergo Heli Samuelem et dixit: " Samuel, fili mi ". Qui respondens ait: " Praesto sum ".
1SAM|3|17|Et interrogavit eum: " Quis est sermo, quem locutus est ad te? Oro te, ne celaveris me. Haec faciat tibi Deus et haec addat, si absconderis a me sermonem ex omnibus verbis, quae dicta sunt tibi ".
1SAM|3|18|Indicavit itaque ei Samuel universos sermones et non abscondit ab eo. Et ille respondit: " Dominus est! Quod bonum est in oculis suis, faciat ".
1SAM|3|19|Crevit autem Samuel, et Dominus erat cum eo, et non cecidit ex omnibus verbis eius in terram.
1SAM|3|20|Et cognovit universus Israel a Dan usque Bersabee quod constitutus esset Samuel propheta Domini.
1SAM|3|21|Et addidit Dominus ut appareret in Silo, quoniam revelatus fuerat Dominus Samueli in Silo iuxta verbum Domini. Et evenit sermo Samuelis universo Israeli.
1SAM|4|1|Et factum est in diebus illis, convenerunt Philisthim in pu gnam; et egressus est Israel obviam Philisthim in proelium et castrametatus est iuxta Abenezer. Porro Philisthim venerunt in Aphec
1SAM|4|2|et instruxerunt aciem contra Israel. Crescente autem certamine, terga vertit Israel Philisthaeis; et caesi sunt in illo certamine passim per agros quasi quattuor milia virorum.
1SAM|4|3|Et reversus est populus ad castra, dixeruntque maiores natu de Israel: " Quare percussit nos Dominus hodie coram Philisthim? Afferamus ad nos de Silo arcam foederis Domini, et veniat in medium nostri, ut salvet nos de manu inimicorum nostrorum ".
1SAM|4|4|Misit ergo populus in Silo, et tulerunt inde arcam foederis Domini exercituum sedentis super cherubim; erantque duo filii Heli cum arca foederis Dei, Ophni et Phinees.
1SAM|4|5|Cumque venisset arca foederis Domini in castra, vociferatus est omnis Israel clamore grandi, et personuit terra.
1SAM|4|6|Et audierunt Philisthim vocem clamoris dixeruntque: " Quaenam est haec vox clamoris magni in castris Hebraeorum? ". Et cognoverunt quod arca Domini venisset in castra.
1SAM|4|7|Timueruntque Philisthim dicentes: " Venit Deus in castra! ". Et ingemuerunt dicentes:
1SAM|4|8|" Vae nobis! Non enim fuit tanta exsultatio heri et nudiustertius. Vae nobis! Quis nos servabit de manu deorum sublimium istorum? Hi sunt dii, qui percusserunt Aegyptum omni plaga in deserto.
1SAM|4|9|Confortamini et estote viri, Philisthim, ne serviatis Hebraeis, sicut illi servierunt vobis. Estote viri et bellate! ".
1SAM|4|10|Pugnaverunt ergo Philisthim, et caesus est Israel, et fugit unusquisque in tabernaculum suum; et facta est plaga magna nimis, et ceciderunt de Israel triginta milia peditum.
1SAM|4|11|Et arca Dei capta est; duoque filii Heli mortui sunt, Ophni et Phinees.
1SAM|4|12|Currens autem vir de Beniamin ex acie venit in Silo in die illo scissa veste et conspersus pulvere caput.
1SAM|4|13|Cumque ille venisset, Heli sedebat super sellam iuxta portam aspectans viam; erat enim cor eius pavens pro arca Dei. Vir autem ille, postquam ingressus est, nuntiavit urbi; et ululavit omnis civitas.
1SAM|4|14|Et audivit Heli sonitum clamoris dixitque: " Quis est hic sonitus tumultus huius? ". At ille festinavit et venit et nuntiavit Heli.
1SAM|4|15|Heli autem erat nonaginta et octo annorum, et oculi eius caligaverant, et videre non poterat.
1SAM|4|16|Et dixit ad Heli: " Ego sum qui veni de proelio et ego qui de acie fugi hodie ". Cui ille ait: " Quid actum est, fili mi? ".
1SAM|4|17|Respondens autem, qui nuntiabat: " Fugit, inquit, Israel coram Philisthim, et ruina magna facta est in populo; insuper et duo filii tui mortui sunt, Ophni et Phinees, et arca Dei capta est ".
1SAM|4|18|Cumque ille nominasset arcam Dei, cecidit de sella retrorsum iuxta ostium et, fractis cervicibus, mortuus est; senex enim erat vir et gravis. Et ipse iudicavit Israel quadraginta annis.
1SAM|4|19|Nurus autem eius, uxor Phinees, praegnans erat vicinaque partui. Et, audito nuntio quod capta esset arca Dei et mortuus socer suus et vir suus, incurvavit se et peperit; irruerant enim in eam dolores subiti.
1SAM|4|20|In ipso autem momento mortis eius dixerunt ei, quae stabant circa eam: Ne timeas, quia filium peperisti ". Quae non respondit eis neque animadvertit.
1SAM|4|21|Et vocavit puerum Ichabod dicens: " Translata est gloria de Israel! ", quia capta est arca Dei et pro socero suo et pro viro suo.
1SAM|4|22|Et ait: " Translata est gloria ab Israel, eo quod capta est arca Dei!.
1SAM|5|1|Philisthim autem tulerunt arcam Dei et asportaverunt eam a Abenezer in Azotum.
1SAM|5|2|Tulerunt Philisthim arcam Dei et intulerunt eam in templum Dagon et statuerunt eam iuxta Dagon.
1SAM|5|3|Cumque surrexissent Azotii altera die, ecce Dagon iacebat pronus in terram ante arcam Domini; et tulerunt Dagon et restituerunt eum in loco suo.
1SAM|5|4|Rursumque mane die altera consurgentes invenerunt Dagon iacentem super faciem suam in terram coram arca Domini; caput autem Dagon et duae palmae manuum eius abscisae erant super limen:
1SAM|5|5|porro Dagon truncus solus remanserat in loco suo. Propter hanc causam non calcant sacerdotes Dagon et omnes, qui ingrediuntur templum eius, super limen Dagon in Azoto usque in hodiernum diem.
1SAM|5|6|Aggravata est autem manus Domini super Azotios, et demolitus est eos et percussit eos tumoribus, Azotum et fines eius.
1SAM|5|7|Videntes autem viri Azotii huiuscemodi plagam dixerunt: " Non maneat arca Dei Israel apud nos, quoniam dura est manus eius super nos et super Dagon deum nostrum ".
1SAM|5|8|Et mittentes congregaverunt omnes principes Philisthinorum ad se et dixerunt: " Quid faciemus de arca Dei Israel? ". Responderuntque: " In Geth circumducatur arca Dei Israel ". Et circumduxerunt arcam Dei Israel.
1SAM|5|9|Postquam autem circumduxerunt eam, facta est manus Domini super civitatem, pavor magnus nimis; et percussit viros urbis a parvo usque ad maiorem, et eruperunt eis tumores.
1SAM|5|10|Miserunt ergo arcam Dei in Accaron.Cumque venisset arca Dei in Accaron, exclamaverunt Accaronitae dicentes: " Adduxerunt ad nos arcam Dei Israel, ut interficiat nos et populum nostrum!.
1SAM|5|11|Miserunt itaque et congregaverunt omnes principes Philisthinorum et dixerunt: " Dimittite arcam Dei Israel, et revertatur in locum suum et non interficiat nos cum populo nostro ".
1SAM|5|12|Fiebat enim pavor mortis in tota civitate, et gravissima valde manus Dei. Viri quoque, qui mortui non fuerant, percutiebantur tumoribus, et ascendebat ululatus civitatis in caelum.
1SAM|6|1|Fuit ergo arca Domini in regio ne Philisthinorum septem mensi bus;
1SAM|6|2|et vocaverunt Philisthim sacerdotes et divinos dicentes: " Quid faciemus de arca Domini? Indicate nobis quomodo remittemus eam in locum suum ".Qui dixerunt:
1SAM|6|3|" Si remittitis arcam Dei Israel, nolite dimittere eam vacuam, sed, quod debetis, reddite ei pro peccato, et tunc curabimini; scietis quare non recedat manus eius a vobis ".
1SAM|6|4|Qui dixerunt: " Quid est quod pro delicto reddere debeamus ei? ". Responderuntque illi:
1SAM|6|5|" Iuxta numerum principum Philisthinorum quinque tumores aureos facietis et quinque mures aureos, quia plaga una fuit omnibus vobis et principibus vestris. Facietisque similitudines tumorum vestrorum et similitudines murium, qui demoliti sunt terram, et dabitis Deo Israel gloriam, si forte relevet manum suam a vobis et a diis vestris et a terra vestra.
1SAM|6|6|Quare gravatis corda vestra, sicut aggravavit Aegyptus et pharao cor suum? Nonne, postquam percussit eos, tunc dimiserunt eos, et abierunt?
1SAM|6|7|Nunc ergo arripite et facite plaustrum novum unum et duas vaccas fetas, quibus non est impositum iugum, iungite in plaustro; et recludite vitulos earum domi.
1SAM|6|8|Tolletisque arcam Domini et ponetis in plaustro; et similitudines aureas, quas exsolvistis ei pro delicto, ponetis in capsella ad latus eius et dimittite eam, ut vadat,
1SAM|6|9|et aspicietis. Et siquidem per viam finium suorum ascenderit contra Bethsames, ipse fecit nobis hoc malum grande; sin autem minime, sciemus quia nequaquam manus eius tetigit nos, sed casu accidit ".
1SAM|6|10|Fecerunt ergo illi hoc modo et tollentes duas vaccas, quae lactabant vitulos, iunxerunt ad plaustrum vitulosque earum concluserunt domi;
1SAM|6|11|et posuerunt arcam Dei super plaustrum et capsellam, quae habebat mures aureos et similitudines tumorum.
1SAM|6|12|Ibant autem in directum vaccae per viam, quae ducit Bethsames, et itinere uno gradiebantur pergentes et mugientes et non declinabant neque ad dextram neque ad sinistram. Sed et principes Philisthim sequebantur usque ad terminos Bethsames.
1SAM|6|13|Porro Bethsamitae metebant triticum in valle; et elevantes oculos viderunt arcam et gavisi sunt, cum vidissent.
1SAM|6|14|Et plaustrum venit in agrum Iosue Bethsamitae et stetit ibi. Erat autem ibi lapis magnus; et conciderunt ligna plaustri vaccasque imposuerunt super ea holocaustum Domino.
1SAM|6|15|Levitae autem deposuerunt arcam Dei et capsellam, quae erat iuxta eam, in qua erant similitudines aureae; et posuerunt super lapidem grandem. Viri autem Bethsamitae obtulerunt holocausta et immolaverunt victimas in die illa Domino.
1SAM|6|16|Et quinque principes Philisthinorum viderunt et reversi sunt in Accaron in die illa.
1SAM|6|17|Hi sunt autem tumores aurei, quos reddiderunt Philisthim pro delicto Domino: Azotus unum, Gaza unum, Ascalon unum, Geth unum, Accaron unum;
1SAM|6|18|et mures aureos secundum numerum urbium Philisthim quinque principum, ab urbe murata usque ad villam, quae erat absque muro; et lapis ille magnus, super quem posuerunt arcam Domini, testis est usque in hunc diem in agro Iosue Bethsamitis.
1SAM|6|19|Filii autem Iechoniae non sunt gavisi super viros Bethsamites quia viderant arcam Domini; et percussit Dominus de populo septuaginta viros. Luxitque populus eo quod Dominus percussisset plebem plaga magna;
1SAM|6|20|et dixerunt viri Bethsamitae: " Quis poterit stare in conspectu Domini, Dei sancti huius? Et ad quem ascendet a nobis? ".
1SAM|6|21|Miseruntque nuntios ad habitatores Cariathiarim dicentes: " Reduxerunt Philisthim arcam Domini. Descendite et ducite eam sursum ad vos ".
1SAM|7|1|Venerunt ergo viri Cariathiarim et duxerunt arcam Domini sursum et intulerunt eam in domum Abinadab in colle; Eleazarum autem filium eius sanctificaverunt, ut custodiret arcam Domini.
1SAM|7|2|Et factum est, ex qua die mansit arca Domini in Cariathiarim, multiplicati sunt dies; erat quippe iam annus vicesimus, et ingemuit omnis domus Israel post Dominum.
1SAM|7|3|Ait autem Samuel ad universam domum Israel dicens: " Si in toto corde vestro revertimini ad Dominum, auferte deos alienos de medio vestri et Astharoth et praeparate corda vestra Domino et servite ei soli, et eruet vos de manu Philisthim ".
1SAM|7|4|Abstulerunt ergo filii Israel Baalim et Astharoth et servierunt Domino soli.
1SAM|7|5|Dixit autem Samuel: " Congregate universum Israel in Maspha, ut orem pro vobis Dominum ".
1SAM|7|6|Et convenerunt in Maspha hauseruntque aquam et effuderunt in conspectu Domini et ieiunaverunt in die illa et dixerunt ibi: " Peccavimus Domino ". Iudicavitque Samuel filios Israel in Maspha.
1SAM|7|7|Et audierunt Philisthim quod congregati essent filii Israel in Maspha, et ascenderunt principes Philisthinorum ad Israel. Quod cum audissent filii Israel, timuerunt a facie Philisthinorum
1SAM|7|8|dixeruntque ad Samuel: " Ne cesses pro nobis clamare ad Dominum Deum nostrum, ut salvet nos de manu Philisthinorum ".
1SAM|7|9|Tulit ergo Samuel agnum lactantem unum et obtulit illum holocaustum integrum Domino; et clamavit Samuel ad Dominum pro Israel, et exaudivit eum Dominus.
1SAM|7|10|Factum est autem cum Samuel offerret holocaustum, Philisthim iniere proelium contra Israel. Intonuit autem Dominus fragore magno in die illa super Philisthim et exterruit eos, et caesi sunt a facie Israel.
1SAM|7|11|Egressique viri Israel de Maspha persecuti sunt Philisthaeos et percusserunt eos usque ad locum, qui erat subter Bethchar.
1SAM|7|12|Tulit autem Samuel lapidem unum et posuit eum inter Maspha et inter Sen et vocavit nomen loci illius Abenezer (id est Lapis adiutorii) dixitque: " Hucusque auxiliatus est nobis Dominus ".
1SAM|7|13|Et humiliati sunt Philisthim nec apposuerunt ultra ut venirent in terminos Israel. Facta est itaque manus Domini super Philisthaeos cunctis diebus Samuel.
1SAM|7|14|Et redditae sunt urbes, quas tulerant Philisthim ab Israel, Israeli ab Accaron usque Geth; et terminos earum liberavit Israel de manu Philisthinorum. Eratque pax inter Israel et Amorraeum.
1SAM|7|15|Iudicabat quoque Samuel Israel cunctis diebus vitae suae
1SAM|7|16|et ibat per singulos annos circumiens Bethel et Galgala et Maspha et iudicabat Israelem in supradictis locis. Revertebaturque in Rama; ibi enim erat domus eius, et ibi iudicabat Israelem. Aedificavit etiam ibi altare Domino.
1SAM|8|1|Factum est autem cum senuis set, Samuel posuit filios suos iu dices Israel.
1SAM|8|2|Fuitque nomen filii eius primogeniti Ioel et nomen secundi Abia; iudicabant in Bersabee.
1SAM|8|3|Et non ambulaverunt filii illius in viis eius, sed declinaverunt post avaritiam acceperuntque munera et perverterunt iudicium.
1SAM|8|4|Congregati ergo universi maiores natu Israel venerunt ad Samuel in Rama
1SAM|8|5|dixeruntque ei: " Ecce tu senuisti, et filii tui non ambulant in viis tuis; nunc ergo constitue nobis regem, ut iudicet nos, sicut universae habent nationes ".
1SAM|8|6|Displicuitque sermo in oculis Samuelis, eo quod dixissent: " Da nobis regem, ut iudicet nos ". Et oravit Samuel ad Dominum.
1SAM|8|7|Dixit autem Dominus ad Samuel: " Audi vocem populi in omnibus, quae loquuntur tibi; non enim te abiecerunt, sed me abiecerunt, ne regnem super eos.
1SAM|8|8|Iuxta omnia opera sua, quae fecerunt a die, qua eduxi eos de Aegypto, usque ad diem hanc, sicut dereliquerunt me et servierunt diis alienis, sic faciunt etiam tibi.
1SAM|8|9|Nunc ergo audi vocem eorum; verumtamen contestare eos et praedic eis ius regis, qui regnaturus est super eos ".
1SAM|8|10|Dixit itaque Samuel omnia verba Domini ad populum, qui petierat a se regem,
1SAM|8|11|et ait: " Hoc erit ius regis, qui imperaturus est vobis: Filios vestros tollet et ponet in curribus suis facietque sibi equites, et current ante quadrigas eius;
1SAM|8|12|et constituet sibi tribunos et centuriones et aratores agrorum suorum et messores segetum et fabros armorum et curruum suorum.
1SAM|8|13|Filias quoque vestras faciet sibi unguentarias et focarias et panificas.
1SAM|8|14|Agros quoque vestros et vineas et oliveta optima tollet et dabit servis suis.
1SAM|8|15|Sed et segetes vestras et vinearum reditus addecimabit, ut det eunuchis et famulis suis.
1SAM|8|16|Servos etiam vestros et ancillas et boves vestros optimos et asinos auferet et ponet in opere suo.
1SAM|8|17|Greges vestros addecimabit, vosque eritis ei servi.
1SAM|8|18|Et clamabitis in die illa a facie regis vestri, quem elegistis vobis, et non exaudiet vos Dominus in die illa ".
1SAM|8|19|Noluit autem populus audire vocem Samuel, sed dixerunt: " Nequaquam: rex enim erit super nos,
1SAM|8|20|et erimus nos quoque sicut omnes gentes; et iudicabit nos rex noster et egredietur ante nos et pugnabit bella nostra pro nobis ".
1SAM|8|21|Et audivit Samuel omnia verba populi et locutus est ea in auribus Domini.
1SAM|8|22|Dixit autem Dominus ad Samuel: " Audi vocem eorum et constitue super eos regem ". Et ait Samuel ad viros Israel: " Vadat unusquisque in civitatem suam ".
1SAM|9|1|Et erat vir de Beniamin nomine Cis filius Abiel filii Seror filii Be chorath filii Aphia, Beniaminita vir potens.
1SAM|9|2|Et erat ei filius vocabulo Saul electus et bonus, et non erat vir de filiis Israel melior illo; ab umero et sursum eminebat super omnem populum.
1SAM|9|3|Perierant autem asinae Cis patris Saul, et dixit Cis ad Saul filium suum: " Tolle tecum unum de pueris et consurgens vade et quaere asinas ". Qui cum transissent per montem Ephraim
1SAM|9|4|et per terram Salisa et non invenissent, transierunt etiam per terram Salim, et non erant, sed et per terram Iemini et minime reppererunt.
1SAM|9|5|Cum autem venissent in terram Suph, dixit Saul ad puerum suum, qui erat cum eo: " Veni, et revertamur, ne forte dimiserit pater meus asinas et sollicitus sit pro nobis ".
1SAM|9|6|Qui ait ei: " Ecce est vir Dei in civitate hac, vir nobilis. Omne quod loquitur, absque ambiguitate venit. Nunc ergo eamus illuc, si forte indicet nobis de via nostra, propter quam venimus ".
1SAM|9|7|Dixitque Saul ad puerum suum: " Ecce ibimus; quid feremus ad virum? Panis defecit in sitarciis nostris, et sportulam non habemus, ut demus homini Dei. Quid habemus? ".
1SAM|9|8|Rursum puer respondit Sauli et ait: " Ecce inventa est in manu mea quarta pars sicli argenti; demus homini Dei, ut indicet nobis viam nostram. -
1SAM|9|9|Olim in Israel sic loquebatur unusquisque vadens consulere Deum: " Venite, et eamus ad videntem "; qui enim propheta dicitur hodie, vocabatur olim videns. -
1SAM|9|10|Et dixit Saul ad puerum suum: " Optimus sermo tuus; veni, eamus ". Et ierunt in civitatem, in qua erat vir Dei.
1SAM|9|11|Cumque ascenderent clivum civitatis, invenerunt puellas egredientes ad hauriendam aquam et dixerunt eis: " Num hic est videns? ".
1SAM|9|12|Quae respondentes dixerunt illis: " Hic est: ecce ante te, festina nunc; hodie enim venit in civitatem, quia sacrificium est hodie populo in excelso.
1SAM|9|13|Ingredientes urbem statim invenietis eum, antequam ascendat excelsum ad vescendum; neque enim comesurus est populus, donec ille veniat, quia ipse benedicit hostiae, et deinceps comedunt, qui vocati sunt. Nunc ergo conscendite, quia statim reperietis eum ".
1SAM|9|14|Et ascenderunt in civitatem. Cumque illi intrarent in urbem, apparuit Samuel egrediens obviam eis, ut ascenderet in excelsum.
1SAM|9|15|Dominus autem revelaverat Samuel, ante unam diem quam veniret Saul, dicens:
1SAM|9|16|" Hac ipsa, quae nunc est hora, cras mittam ad te virum de terra Beniamin, et unges eum ducem super populum meum Israel, et salvabit populum meum de manu Philisthinorum, quia respexi populum meum; venit enim clamor eorum ad me ".
1SAM|9|17|Cumque aspexisset Samuel Saulem, Dominus ait ei: " Ecce vir, quem dixeram tibi; iste dominabitur populo meo ".
1SAM|9|18|Accessit autem Saul ad Samuelem in medio portae et ait: " Indica, oro, mihi: Ubi est domus videntis? ".
1SAM|9|19|Et respondit Samuel Sauli dicens: " Ego sum videns. Ascende ante me in excelsum, ut comedatis mecum hodie. Et dimittam te mane et omnia, quae sunt in corde tuo, indicabo tibi;
1SAM|9|20|et de asinis, quas perdidisti nudiustertius, ne sollicitus sis, quia inventae sunt. Et cuius erunt optima quaeque Israel? Nonne tibi et omni domui patris tui? ".
1SAM|9|21|Respondens autem Saul ait: "Numquid non Beniaminita ego sum de minima tribu Israel, et cognatio mea novissima inter omnes familias de tribu Beniamin? Quare ergo locutus es mihi sermonem istum? ".
1SAM|9|22|Assumens itaque Samuel Saulem et puerum eius introduxit eos in triclinium et dedit eis locum in capite eorum, qui fuerant invitati: erant enim quasi triginta viri.
1SAM|9|23|Dixitque Samuel coco: " Da partem, quam dedi tibi et praecepi, ut reponeres seorsum apud te ".
1SAM|9|24|Levavit autem cocus armum et caudam et posuit ante Saul. Dixitque Samuel: " Ecce quod remansit; pone ante te et comede, quia de industria servatum est tibi, quando populum vocavi ". Et comedit Saul cum Samuel in die illa.
1SAM|9|25|Et descenderunt de excelso in oppidum. Et straverunt pro Saul in solario, et dormivit.
1SAM|9|26|Cumque mane surrexissent, et iam elucesceret, vocavit Samuel Saul in solario dicens: " Surge, ut dimittam te ". Et surrexit Saul. Egressique sunt ambo, ipse videlicet et Samuel.
1SAM|9|27|Cumque descenderent in extrema parte civitatis, Samuel dixit ad Saul: " Dic puero, ut antecedat nos - et ille antecessit C; tu autem subsiste paulisper, ut indicem tibi verbum Domini ".
1SAM|10|1|Tulit autem Samuel lenticulam olei et effudit super caput eius et deosculatus eum ait: " Ecce unxit te Dominus in principem super populum suum, super Israel. Et tu dominaberis populo Domini et tu liberabis eum de manu inimicorum eius, qui in circuitu eius sunt. Et hoc tibi signum quia unxit te Deus in principem super hereditatem suam:
1SAM|10|2|cum abieris hodie a me, invenies duos viros iuxta sepulcrum Rachel in finibus Beniamin, dicentque tibi: "Inventae sunt asinae, ad quas ieras perquirendas; et intermissis pater tuus asinis sollicitus est pro vobis et dicit: Quid faciam de filio meo?".
1SAM|10|3|Cumque abieris inde et ultra transieris et veneris ad quercum Thabor, invenient te ibi tres viri ascendentes ad Deum in Bethel: unus portans tres haedos et alius tres tortas panis et alius portans utrem vini.
1SAM|10|4|Cumque te salutaverint, dabunt tibi duos panes, et accipies de manu eorum.
1SAM|10|5|Post haec venies in Gabaa Dei, ubi est statio Philisthinorum; et, cum ingressus fueris ibi urbem, obviam habebis gregem prophetarum descendentium de excelso et ante eos psalterium et tympanum et tibiam et citharam ipsosque prophetantes.
1SAM|10|6|Et insiliet in te spiritus Domini, et prophetabis cum eis et mutaberis in virum alium.
1SAM|10|7|Quando ergo evenerint signa haec omnia tibi, fac, quaecumque invenerit manus tua, quia Dominus tecum est.
1SAM|10|8|Et descendes ante me in Galgala. Ego quippe descendam ad te, ut offeram oblationem et immolem victimas pacificas. Septem diebus exspectabis, donec veniam ad te et ostendam tibi, quae facias ".
1SAM|10|9|Itaque, cum avertisset umerum suum, ut abiret a Samuele, immutavit ei Deus cor aliud, et venerunt omnia signa haec in die illa.
1SAM|10|10|Veneruntque inde in Gabaa, et ecce grex prophetarum obvius ei; et insiluit super eum spiritus Dei, et prophetavit in medio eorum.
1SAM|10|11|Videntes autem omnes, qui noverant eum heri et nudiustertius, quod esset cum prophetis et prophetaret, dixerunt ad invicem: " Quaenam res accidit filio Cis? Num et Saul inter prophetas? ".
1SAM|10|12|Responditque vir loci illius dicens: " Et quis pater eorum? ". Propterea versum est in proverbium: " Num et Saul inter prophetas? ".
1SAM|10|13|Cessavit autem prophetare et venit in Gabaa;
1SAM|10|14|dixitque patruus Saul ad eum et ad puerum eius: " Quo abistis? ". Qui respondit: " Quaerere asinas; quas cum non repperissemus, venimus ad Samuelem".
1SAM|10|15|Et dixit ei patruus suus: "Indica mihi quid dixerit tibi Samuel".
1SAM|10|16|Et ait Saul ad patruum suum: " Indicavit nobis quia inventae essent asinae ". De sermone autem regni non indicavit ei, quem locutus illi fuerat Samuel.
1SAM|10|17|Et convocavit Samuel populum ad Dominum in Maspha
1SAM|10|18|et ait ad filios Israel: " Haec dicit Dominus, Deus Israel: Ego eduxi Israel de Aegypto et erui vos de manu Aegyptiorum et de manu omnium regnorum, quae affligebant vos.
1SAM|10|19|Vos autem hodie proiecistis Deum vestrum, qui solus salvavit vos de universis malis et tribulationibus vestris, et dixistis: "Nequaquam, sed regem constitue super nos!". Nunc ergo state coram Domino per tribus vestras et per familias ".
1SAM|10|20|Et applicuit Samuel omnes tribus Israel; et cecidit sors in tribum Beniamin.
1SAM|10|21|Et applicuit tribum Beniamin et cognationes eius; et cecidit in cognationem Metri et pervenit usque ad Saul filium Cis. Quaesierunt ergo eum, et non est inventus.
1SAM|10|22|Et consuluerunt post haec Dominum, utrumnam venisset illuc vir. Responditque Dominus: " Ecce absconditus est inter sarcinas ".
1SAM|10|23|Cucurrerunt itaque et tulerunt eum inde; stetitque in medio populi et altior fuit universo populo ab umero et sursum.
1SAM|10|24|Et ait Samuel ad omnem populum: Certe videtis, quem elegit Dominus, quoniam non sit similis ei in omni populo ". Et clamavit cunctus populus et ait: " Vivat rex! ".
1SAM|10|25|Locutus est autem Samuel ad populum legem regni et scripsit in libro et reposuit coram Domino; et dimisit Samuel omnem populum, singulos in domum suam.
1SAM|10|26|Sed et Saul abiit in domum suam in Gabaa; et abierunt cum eo viri fortes, quorum tetigerat Deus corda.
1SAM|10|27|Filii vero Belial dixerunt: " Num salvare nos poterit iste? ". Et despexerunt eum et non attulerunt ei munera; ille vero dissimulabat se audire.
1SAM|11|1|Ascendit autem Naas Am monites et pugnare coepit ad versum Iabes Galaad. Dixeruntque omnes viri Iabes ad Naas: " Habeto nos foederatos, et serviemus tibi ".
1SAM|11|2|Et respondit ad eos Naas Ammonites: " In hoc feriam vobiscum foedus, ut eruam omnium vestrum oculos dextros ponamque vos opprobrium in universo Israel ".
1SAM|11|3|Et dixerunt ad eum seniores Iabes: " Concede nobis septem dies, ut mittamus nuntios in universos terminos Israel; et, si non fuerit qui defendat nos, egrediemur ad te ".
1SAM|11|4|Venerunt ergo nuntii in Gabaa Saulis et locuti sunt verba audiente populo; et levavit omnis populus vocem suam et flevit.
1SAM|11|5|Et ecce Saul veniebat sequens boves de agro et ait: " Quid habet populus quod plorat? ". Et narraverunt ei verba virorum Iabes.
1SAM|11|6|Et insilivit spiritus Domini in Saul, cum audisset verba haec; et iratus est furor eius nimis.
1SAM|11|7|Et assumens par boum concidit in frusta misitque in omnes terminos Israel per manum nuntiorum dicens: " Quicumque non exierit secutusque fuerit Saul et Samuel, sic fiet bobus eius ". Invasit ergo timor Domini populum, et egressi sunt quasi vir unus.
1SAM|11|8|Et recensuit eos in Bezec: fueruntque filiorum Israel trecenta milia; virorum autem Iudae triginta milia.
1SAM|11|9|Et dixit nuntiis, qui venerant: " Sic dicetis viris, qui sunt in Iabes Galaad: Cras erit vobis salus, cum incaluerit sol ". Venerunt ergo nuntii et annuntiaverunt viris Iabes, qui laetati sunt
1SAM|11|10|et dixerunt: "Mane exibimus ad vos, et facietis nobis omne, quod placuerit vobis ".
1SAM|11|11|Et factum est, cum venisset dies crastinus, constituit Saul populum in tres partes; et ingressi sunt media castra in vigilia matutina et percusserunt Ammon, usque dum incalesceret dies. Reliqui autem dispersi sunt, ita ut non relinquerentur in eis duo pariter.
1SAM|11|12|Et ait populus ad Samuel: " Quis est iste qui dixit: "Saul num regnabit super nos?". Date viros, et interficiemus eos ".
1SAM|11|13|Et ait Saul: " Non occidetur quisquam in die hac, quia hodie fecit Dominus salutem in Israel".
1SAM|11|14|Dixit autem Samuel ad populum: " Venite, et eamus in Galgala et innovemus ibi regnum ".
1SAM|11|15|Et perrexit omnis populus in Galgala, et fecerunt ibi regem Saul coram Domino in Galgala; et immolaverunt ibi victimas pacificas coram Domino. Et laetatus est ibi Saul et cuncti viri Israel nimis.
1SAM|12|1|Dixit autem Samuel ad universum Israel: " Ecce audivi vocem vestram iuxta omnia, quae locuti estis ad me, et constitui super vos regem;
1SAM|12|2|et nunc rex graditur ante vos. Ego autem senui et incanui; porro filii mei vobiscum sunt. Itaque conversatus coram vobis ab adulescentia mea usque ad hanc diem;
1SAM|12|3|ecce praesto sum. Loquimini contra me coram Domino et coram christo eius, utrum bovem cuiusquam tulerim an asinum, si quempiam calumniatus sum, si oppressi aliquem, si de manu cuiusquam munus accepi, ut oculos meos clauderem in eius causa. Restituam vobis ".
1SAM|12|4|Et dixerunt: " Non es calumniatus nos neque oppressisti neque tulisti de manu alicuius quippiam ".
1SAM|12|5|Dixitque ad eos: " Testis Dominus adversum vos, et testis christus eius in die hac, quia non inveneritis in manu mea quippiam ". Et dixerunt: " Testis ".
1SAM|12|6|Et ait Samuel ad populum: " Testis est Dominus, qui fecit Moysen et Aaron et eduxit patres nostros de terra Aegypti.
1SAM|12|7|Nunc ergo state, ut iudicio contendam adversum vos coram Domino de omnibus misericordiis Domini, quas fecit vobiscum et cum patribus vestris:
1SAM|12|8|quomodo ingressus est Iacob in Aegyptum, et oppresserunt eos Aegyptii; et clamaverunt patres vestri ad Dominum, et misit Dominus Moysen et Aaron et eduxit patres vestros ex Aegypto et collocavit eos in loco hoc;
1SAM|12|9|qui obliti sunt Domini Dei sui, et tradidit eos in manu Sisarae magistri militiae Asor et in manu Philisthinorum et in manu regis Moab, et pugnaverunt adversum eos.
1SAM|12|10|Postea autem clamaverunt ad Dominum et dixerunt: "Peccavimus, quia dereliquimus Dominum et servivimus Baalim et Astharoth; nunc ergo erue nos de manu inimicorum nostrorum, et serviemus tibi".
1SAM|12|11|Et misit Dominus Ierobbaal et Barac et Iephte et Samuel et eruit vos de manu inimicorum vestrorum per circuitum; et habitastis confidenter.
1SAM|12|12|Videntes autem quod Naas rex filiorum Ammon venisset adversum vos, dixistis mihi: "Nequaquam, sed rex imperabit nobis!", cum Dominus Deus vester regnaret in vobis.
1SAM|12|13|Nunc ergo praesto est rex vester, quem elegistis et petistis; ecce dedit vobis Dominus regem.
1SAM|12|14|Si timueritis Dominum et servieritis ei et audieritis vocem eius et non contempseritis sermonem Domini, eritis et vos et rex, qui imperat vobis, sequentes Dominum Deum vestrum.
1SAM|12|15|Si autem non audieritis vocem Domini, sed contempseritis sermonem Domini, erit manus Domini super vos et super regem vestrum, ut disperdat vos.
1SAM|12|16|Sed et nunc state et videte rem istam grandem, quam facturus est Dominus in conspectu vestro.
1SAM|12|17|Numquid non messis tritici est hodie? Invocabo Dominum, et dabit tonitrua et pluvias; et scietis et videbitis quia grande malum feceritis vobis in conspectu Domini petentes super vos regem ".
1SAM|12|18|Et clamavit Samuel ad Dominum, et dedit Dominus tonitrua et pluviam in die illa.
1SAM|12|19|Et timuit omnis populus nimis Dominum et Samuel; dixitque universus populus ad Samuel: " Ora pro servis tuis ad Dominum Deum tuum, ut non moriamur: addidimus enim universis peccatis nostris malum, ut peteremus nobis regem ".
1SAM|12|20|Dixit autem Samuel ad populum: " Nolite timere. Vos fecistis universum malum hoc; verumtamen nolite recedere a tergo Domini et servite Domino in omni corde vestro;
1SAM|12|21|et nolite declinare post vana, quae non proderunt vobis neque eruent vos, quia vana sunt;
1SAM|12|22|profecto non derelinquet Dominus populum suum propter nomen suum magnum, quia dignatus est Dominus facere vos sibi populum.
1SAM|12|23|Absit autem a me hoc peccatum in Dominum, ut cessem orare pro vobis et docere vos viam bonam et rectam.
1SAM|12|24|Igitur timete Dominum et servite ei in veritate et ex toto corde vestro; vidistis enim magnifica, quae in vobis gesserit.
1SAM|12|25|Quod si perseveraveritis in malitia, et vos et rex vester pariter peribitis ".
1SAM|13|1|Filius annorum Saul, cum regnare coepisset; duobus au tem annis regnavit super Israel.
1SAM|13|2|Et elegit sibi Saul tria milia de Israel: et erant cum Saul duo milia in Machmas et in monte Bethel, mille autem cum Ionathan in Gabaa Beniamin. Porro ceterum populum remisit unumquemque in tabernacula sua.
1SAM|13|3|Et percussit Ionathan stationem Philisthinorum, quae erat in Gabaa. Quod audierunt Philisthim; Saul autem cecinit bucina in omni terra dicens: " Audiant Hebraei! ".
1SAM|13|4|Et universus Israel audivit huiuscemodi famam: " Percussit Saul stationem Philisthinorum; et factus est Israel odiosus Philisthim ". Ergo populus congregatus est post Saul in Galgala.
1SAM|13|5|Et Philisthim congregati sunt ad proeliandum contra Israel: tria milia curruum et sex milia equitum et reliquum vulgus plurimum sicut arena, quae est in litore maris. Et ascendentes castrametati sunt in Machmas ad orientem Bethaven.
1SAM|13|6|Quod cum vidissent viri Israel se in arto sitos - afflictus est enim populus - absconderunt se in speluncis et in abditis, in petris quoque et in antris et in cisternis.
1SAM|13|7|Hebraei autem transierunt Iordanem in terram Gad et Galaad.Cumque adhuc esset Saul in Galgalis, universus populus perterritus est, qui sequebatur eum.
1SAM|13|8|Et exspectavit septem diebus iuxta placitum Samuel, et non venit Samuel in Galgala; dilapsusque est populus ab eo.
1SAM|13|9|Ait ergo Saul: " Afferte mihi holocaustum et pacifica ". Et obtulit holocaustum.
1SAM|13|10|Cumque complesset offerens holocaustum, ecce Samuel veniebat; et egressus est Saul obviam ei, ut salutaret eum.
1SAM|13|11|Locutusque est ad eum Samuel: " Quid fecisti? ". Respondit Saul: " Quia vidi quod dilaberetur populus a me, et tu non veneras iuxta placitos dies, porro Philisthim congregati fuerant in Machmas,
1SAM|13|12|dixi: Nunc descendent Philisthim ad me in Galgala, et faciem Domini non placavi. Necessitate compulsus obtuli holocaustum ".
1SAM|13|13|Dixitque Samuel ad Saul: " Stulte egisti. Utinam custodisses mandata Domini Dei tui, quae praecepit tibi! Profecto nunc confirmasset Dominus regnum tuum super Israel in sempiternum;
1SAM|13|14|sed nequaquam regnum tuum ultra consurget. Quaesivit sibi Dominus virum iuxta cor suum; et constituit eum Dominus ducem super populum suum, eo quod non servaveris, quae praecepit Dominus ".
1SAM|13|15|Surrexit autem Samuel et ascendit de Galgalis et abiit per viam suam. Et reliquus populus ascendit post Saul obviam exercitui bellatorum. Et venerunt de Galgalis in Gabaa Beniamin. Et recensuit Saul populum, qui inventi fuerant cum eo, quasi sescentos viros.
1SAM|13|16|Et Saul et Ionathan filius eius populusque, qui erat cum eis, erat in Gabaa Beniamin; porro Philisthim consederant in Machmas.
1SAM|13|17|Et egressi sunt ad praedandum de castris Philisthinorum tres cunei: unus cuneus pergebat contra viam Ophra ad terram Sual,
1SAM|13|18|porro alius ingrediebatur per viam Bethoron, tertius autem verterat se ad iter termini imminentis valli Seboim contra desertum.
1SAM|13|19|Porro faber ferrarius non inveniebatur in omni terra Israel; caverant enim Philisthim, ne forte facerent Hebraei gladium aut lanceam.
1SAM|13|20|Descendebat ergo omnis Israel ad Philisthim, ut exacueret unusquisque vomerem suum et ligonem et securim et falcem.
1SAM|13|21|Pretium autem exacutionis erat: pro vomeribus et ligonibus duae partes sicli, et tertia pars sicli ad acuendas secures et ad stimulum corrigendum.
1SAM|13|22|Cumque venisset dies proelii Machmas, non est inventus ensis et lancea in manu totius populi, qui erat cum Saul et cum Ionathan, excepto Saul et Ionathan filio eius.
1SAM|13|23|Egressa est autem statio Philisthim ad fauces Machmas.
1SAM|14|1|Et accidit quadam die, ut diceret Ionathan filius Saul ad adulescentem armigerum suum: " Veni, et transeamus ad stationem Philisthim, quae est ibi ex adverso ". Patri autem suo hoc ipsum non indicavit.
1SAM|14|2|Porro Saul morabatur in extrema parte Gabaa sub malogranato, quae erat in Magron; et erat populus cum eo quasi sescentorum virorum.
1SAM|14|3|Et Ahias filius Achitob fratris Ichabod filii Phinees, qui ortus fuerat ex Heli sacerdote Domini in Silo, portabat ephod. Sed et populus ignorabat quod isset Ionathan.
1SAM|14|4|Erant autem inter ascensus, per quos nitebatur Ionathan transire ad stationem Philisthinorum, dens rupis hinc ex una parte et dens rupis illinc ex altera parte: nomen uni Boses et nomen alteri Sene;
1SAM|14|5|unus scopulus prominens ad aquilonem ex adverso Machmas et alter a meridie contra Gabaa.
1SAM|14|6|Dixit autem Ionathan ad adulescentem armigerum suum: " Veni, transeamus ad stationem incircumcisorum horum, si forte faciat Dominus pro nobis; quia non est Domino difficile salvare vel in multitudine vel in paucis ".
1SAM|14|7|Dixitque ei armiger suus: " Fac omnia, quae placent animo tuo. Perge quo cupis; ego ero tecum ubicumque volueris ".
1SAM|14|8|Et ait Ionathan: " Ecce nos transimus ad viros istos. Cumque apparuerimus eis,
1SAM|14|9|si taliter locuti fuerint ad nos: "Manete, donec veniamus ad vos", stemus in loco nostro nec ascendamus ad eos.
1SAM|14|10|Si autem dixerint: "Ascendite ad nos", ascendamus, quia tradidit eos Dominus in manibus nostris; hoc erit nobis signum ".
1SAM|14|11|Apparuit igitur uterque stationi Philisthinorum. Dixeruntque Philisthim: " En Hebraei egrediuntur de cavernis, in quibus absconditi fuerant ".
1SAM|14|12|Et locuti sunt viri de statione ad Ionathan et ad armigerum eius dixeruntque: " Ascendite ad nos, et ostendimus vobis rem ". Et ait Ionathan ad armigerum suum: " Ascendamus; sequere me, tradidit enim eos Dominus in manu Israel ".
1SAM|14|13|Ascendit autem Ionathan reptans manibus et pedibus et armiger eius post eum; Philisthim cadebant ante Ionathan, et eos armiger eius interficiebat sequens eum.
1SAM|14|14|Et facta est plaga prima, qua percussit Ionathan et armiger eius quasi viginti viros in media fere parte iugeri.
1SAM|14|15|Et factus est terror in castris per agros; sed et omnis populus stationis eorum et, qui ierant ad praedandum, obstupuerunt; et conturbata est terra, et factus est terror a Deo.
1SAM|14|16|Et respexerunt speculatores Saul, qui erant in Gabaa Beniamin; et ecce multitudo fluctuabat huc illucque diffugiens.
1SAM|14|17|Et ait Saul populo, qui erat cum eo: " Requirite et videte quis abierit ex nobis ". Cumque requisissent, repertum est non adesse Ionathan et armigerum eius.
1SAM|14|18|Et ait Saul ad Ahiam: " Applica ephod ". Ipse enim portabat ephod in die illa in conspectu filiorum Israel.
1SAM|14|19|Cumque loqueretur Saul ad sacerdotem, tumultus maior fiebat in castris Philisthinorum, crescebatque paulatim et clarius reboabat. Et ait Saul ad sacerdotem: " Contrahe manum tuam ".
1SAM|14|20|Congregati ergo sunt Saul et omnis populus, qui erat cum eo, et venerunt usque ad locum certaminis. Et ecce versus fuerat gladius uniuscuiusque ad proximum suum: perturbatio magna nimis.
1SAM|14|21|Sed et Hebraei, qui fuerant cum Philisthim heri et nudiustertius ascenderantque cum eis in castris, reversi sunt et ipsi, ut essent cum Israel, qui erant cum Saul et Ionathan.
1SAM|14|22|Omnes quoque Israelitae, qui se absconderant in monte Ephraim, audientes quod fugissent Philisthim, sociaverunt se et ipsi cum suis in proelio.
1SAM|14|23|Et salvavit Dominus in die illa Israel; pugna autem pervenit ultra Bethaven.
1SAM|14|24|Et viri Israel comprimebant se in die illa. Adiuravit autem Saul populum dicens: " Maledictus vir, qui comederit panem usque ad vesperam, donec ulciscar de inimicis meis! ". Et non manducavit universus populus panem.
1SAM|14|25|Omneque terrae vulgus venit in saltum, in quo erat mel super faciem agri.
1SAM|14|26|Ingressus est itaque populus saltum, et apparuit fluens mel. Nullusque applicuit manum ad os suum; timebat enim populus iuramentum.
1SAM|14|27|Porro Ionathan non audierat, cum adiuraret pater eius populum; extenditque summitatem virgae, quam habebat in manu, et intinxit in favo mellis et convertit manum suam ad os suum, et illuminati sunt oculi eius.
1SAM|14|28|Respondensque unus de populo ait: " Iureiurando constrinxit pater tuus populum dicens: "Maledictus, qui comederit panem hodie!". Defecit autem populus ".
1SAM|14|29|Dixitque Ionathan: " Turbavit pater meus terram! Videte quia illuminati sunt oculi mei, eo quod gustaverim paululum de melle isto;
1SAM|14|30|quanto magis si comedisset hodie populus de praeda inimicorum suorum, quam repperit? Nonne nunc maior facta fuisset plaga in Philisthim? ".
1SAM|14|31|Percusserunt ergo in die illa Philisthaeos a Machmis usque in Aialon; defatigatus est autem populus nimis.
1SAM|14|32|Et versus ad praedam tulit oves et boves et vitulos; et mactaverunt in terra, comeditque populus cum sanguine.
1SAM|14|33|Nuntiaverunt autem Saul dicentes: " Ecce populus peccat Domino comedens cum sanguine ". Qui ait: " Praevaricati estis! Volvite ad me huc saxum grande ".
1SAM|14|34|Et dixit Saul: " Dispergimini in vulgus et dicite eis, ut adducat ad me unusquisque bovem suum et arietem, et occidite super istud et vescimini; et non peccabitis Domino comedentes cum sanguine ". Adduxit itaque omnis populus, unusquisque quod erat in manu sua illa nocte, et occiderunt ibi.
1SAM|14|35|Aedificavit autem Saul altare Domino. Tuncque primum coepit aedificare altare Domino.
1SAM|14|36|Et dixit Saul: " Irruamus super Philisthim nocte et vastemus eos, usquedum illucescat mane; nec relinquamus de eis virum ". Dixitque populus: " Omne, quod bonum videtur in oculis tuis, fac ". Et ait sacerdos: " Accedamus huc ad Deum ".
1SAM|14|37|Et consuluit Saul Deum: " Num persequar Philisthim? Numquid trades eos in manu Israel? ". Et non respondit ei in die illa.
1SAM|14|38|Dixitque Saul: " Accedite huc, universi duces populi, et scitote et videte per quem acciderit peccatum hoc hodie.
1SAM|14|39|Vivit Dominus, salvator Israel, quia si per Ionathan filium meum factum est, absque retractatione morietur ". Ad quod nullus contradixit ei de omni populo.
1SAM|14|40|Et ait ad universum Israel: " Separamini vos in partem unam, et ego cum Ionathan filio meo ero in parte altera ". Respondit populus ad Saul: " Quod bonum videtur in oculis tuis, fac ".
1SAM|14|41|Et dixit Saul ad Dominum, Deum Israel: " Quid est quod non responderis servo tuo hodie? Si est in me aut in Ionathan filio meo iniquitas ista, Domine, Deus Israel, da Urim; sed, si est haec iniquitas in populo tuo Israel, da Tummim ". Et deprehensus est Ionathan et Saul; populus autem salvus evasit.
1SAM|14|42|Et ait Saul: " Mittite sortem inter me et inter Ionathan filium meum ". Et captus est Ionathan.
1SAM|14|43|Dixit autem Saul ad Ionathan: " Indica mihi quid feceris ". Et indicavit ei Ionathan et ait: " Gustans gustavi in summitate virgae, quae erat in manu mea, paululum mellis et ecce ego morior ".
1SAM|14|44|Et ait Saul: " Haec faciat mihi Deus et haec addat, nisi morte morieris, Ionathan ".
1SAM|14|45|Dixitque populus ad Saul: " Ergone Ionathan morietur, qui fecit salutem hanc magnam in Israel? Hoc nefas est; vivit Dominus, quia non cadet capillus de capite eius in terram, quia cum Deo operatus est hodie ". Liberavit ergo populus Ionathan, ut non moreretur.
1SAM|14|46|Recessitque Saul nec persecutus est Philisthim; porro Philisthim abierunt in loca sua.
1SAM|14|47|At Saul, confirmato regno super Israel, pugnabat per circuitum adversum omnes inimicos eius: contra Moab et filios Ammon et Edom et reges Soba et Philisthaeos; et, quocumque se verterat, superabat.
1SAM|14|48|Fortiter egit et percussit Amalec et eruit Israel de manu vastatorum eius.
1SAM|14|49|Fuerunt autem filii Saul Ionathan et Isui et Melchisua. Nomina duarum filiarum eius: nomen primogenitae Merob et nomen minoris Michol.
1SAM|14|50|Et nomen uxoris Saul Achinoam filia Achimaas, et nomen principis militiae eius Abner filius Ner patrui Saul.
1SAM|14|51|Porro Cis pater Saul et Ner pater Abner fuerunt filii Abiel.
1SAM|14|52|Erat autem bellum potens adversum Philisthaeos omnibus diebus Saul; nam, quemcumque viderat Saul virum fortem et aptum ad proelium, sociabat eum sibi.
1SAM|15|1|Et dixit Samuel ad Saul: " Me misit Dominus, ut unge rem te in regem super populum eius Israel. Nunc ergo audi vocem Domini.
1SAM|15|2|Haec dicit Dominus exercituum: "Recensui, quaecumque fecit Amalec Israeli, quomodo restitit ei in via, cum ascenderet de Aegypto.
1SAM|15|3|Nunc igitur vade et demolire Amalec et percute anathemate universa eius; non parcas ei, sed interfice a viro usque ad mulierem et parvulum atque lactantem, bovem et ovem, camelum et asinum" ".
1SAM|15|4|Convocavit itaque Saul populum et recensuit eos in Telem: ducenta milia peditum et decem milia virorum Iudae.
1SAM|15|5|Cumque venisset Saul usque ad civitatem Amalec, tetendit insidias in torrente
1SAM|15|6|dixitque Saul Cinaeo: " Abite, recedite atque descendite ab Amalec, ne forte perdam te cum eo; tu enim fecisti misericordiam cum omnibus filiis Israel, cum ascenderent de Aegypto ". Et recessit Cinaeus de medio Amalec.
1SAM|15|7|Percussitque Saul Amalec ab Hevila usque ad Sur, quae est e regione Aegypti.
1SAM|15|8|Et apprehendit Agag regem Amalec vivum; omne autem vulgus interfecit in ore gladii.
1SAM|15|9|Et pepercit Saul et populus Agag et optimis gregibus ovium et armentorum, pinguibus scilicet pecoribus et agnis et universis, quae pulchra erant, nec voluerunt disperdere ea; quidquid vero vile fuit et reprobum, hoc demoliti sunt.
1SAM|15|10|Factum est autem verbum Domini ad Samuel dicens:
1SAM|15|11|" Paenitet me quod constituerim Saul regem, quia dereliquit me et verba mea opere non implevit ". Contristatusque est Samuel et clamavit ad Dominum tota nocte.
1SAM|15|12|Cumque de nocte surrexisset Samuel, ut iret ad Saul mane, nuntiatum est Samueli quod venisset Saul in Carmel et erexisset sibi trophaeum et reversus transisset descendissetque in Galgala.
1SAM|15|13|Et cum venisset Samuel ad Saul, dixit ei Saul: " Benedictus tu Domino; implevi verbum Domini ".
1SAM|15|14|Dixitque Samuel: " Et quae est haec vox gregum, quae resonat in auribus meis, et armentorum, quam ego audio? ".
1SAM|15|15|Et ait Saul: " De Amalec adduxerunt ea; pepercit enim populus melioribus ovibus et armentis, ut immolarentur Domino Deo tuo; reliqua vero occidimus ".
1SAM|15|16|Dixit autem Samuel ad Saul: " Sine me, et indicabo tibi, quae locutus sit Dominus ad me nocte ". Dixitque ei: " Loquere ".
1SAM|15|17|Et ait Samuel: " Nonne, cum parvulus esses in oculis tuis, caput in tribubus Israel factus es? Unxitque te Dominus regem super Israel
1SAM|15|18|et misit te Dominus in viam et ait: " Vade et interfice peccatores Amalec et pugnabis contra eos usque ad internecionem eorum ".
1SAM|15|19|Quare ergo non audisti vocem Domini, sed versus ad praedam es et fecisti malum in oculis Domini? ".
1SAM|15|20|Et ait Saul ad Samuelem: " Immo audivi vocem Domini et ambulavi in via, per quam misit me Dominus; et adduxi Agag regem Amalec et Amalec interfeci.
1SAM|15|21|Tulit autem populus de praeda oves et boves, primitias eorum, quae caesa sunt, ut immolet Domino Deo tuo in Galgalis ".
1SAM|15|22|Et ait Samuel: " Numquid vult Dominus holocausta aut victimas et non potius ut oboediatur voci Domini? Melior est enim oboedientia quam victimae, et auscultare magis quam offerre adipem arietum.
1SAM|15|23|Vere peccatum hariolandi est repugnare, et scelus idololatriae nolle acquiescere: pro eo ergo quod abiecisti sermonem Domini, abiecit te, ne sis rex ".
1SAM|15|24|Dixitque Saul ad Samuelem: " Peccavi, quia praevaricatus sum sermonem Domini et verba tua timens populum et oboediens voci eorum;
1SAM|15|25|sed nunc tolle, quaeso, peccatum meum et revertere mecum, ut adorem Dominum ".
1SAM|15|26|Et ait Samuel ad Saul: " Non revertar tecum, quia proiecisti sermonem Domini; et proiecit te Dominus, ne sis rex super Israel ".
1SAM|15|27|Et conversus est Samuel, ut abiret; ille autem apprehendit summitatem pallii eius, quae et scissa est.
1SAM|15|28|Et ait ad eum Samuel: " Scidit Dominus regnum Israel a te hodie et tradidit illud proximo tuo meliori te.
1SAM|15|29|Porro Gloria Israel non mentitur et paenitudine non flectitur; neque enim homo est, ut agat paenitentiam ".
1SAM|15|30|At ille ait: " Peccavi, sed nunc honora me coram senibus populi mei et coram Israel; et revertere mecum, ut adorem Dominum Deum tuum ".
1SAM|15|31|Reversus ergo Samuel secutus est Saulem et adoravit Saul Dominum.
1SAM|15|32|Dixitque Samuel: " Adducite ad me Agag regem Amalec ". Et oblatus est ei Agag tremens. Et dixit Agag: " Certe secessit amaritudo mortis! ".
1SAM|15|33|Et ait Samuel: " Sicut fecit absque liberis mulieres gladius tuus, sic absque liberis erit inter mulieres mater tua ". Et in frusta concidit Samuel Agag coram Domino in Galgalis.
1SAM|15|34|Abiit autem Samuel in Rama; Saul vero ascendit in domum suam in Gabaa Saulis.
1SAM|15|35|Et non vidit Samuel ultra Saul usque ad diem mortis suae; verumtamen lugebat Samuel Saul, quoniam Dominum paenitebat quod constituisset Saul regem super Israel.
1SAM|16|1|Dixitque Dominus ad Samuelem: " Usquequo tu luges Saul, cum ego proiecerim eum, ne regnet super Israel? Imple cornu tuum oleo et veni, ut mittam te ad Isai Bethlehemitem; providi enim in filiis eius mihi regem ".
1SAM|16|2|Et ait Samuel: " Quomodo vadam? Audiet enim Saul et interficiet me ". Et ait Dominus: " Vitulam de armento tolles in manu tua et dices: "Ad immolandum Domino veni".
1SAM|16|3|Et vocabis Isai ad victimam; et ego ostendam tibi quid facias, et unges quemcumque monstravero tibi ".
1SAM|16|4|Fecit ergo Samuel, sicut locutus est ei Dominus, venitque in Bethlehem. Et expaverunt seniores civitatis occurrentes ei dixeruntque: " Pacificusne ingressus tuus? ".
1SAM|16|5|Et ait: " Pacificus; ad immolandum Domino veni. Sanctificamini et venite mecum, ut immolem ". Sanctificavit ergo Isai et filios eius et vocavit eos ad sacrificium.
1SAM|16|6|Cumque ingressi essent, vidit Eliab et ait: " Absque dubio coram Domino est christus eius! ".
1SAM|16|7|Et dixit Dominus ad Samuelem: " Ne respicias vultum eius neque altitudinem staturae eius, quoniam abieci eum; nec iuxta intuitum hominis iudico: homo enim videt ea, quae parent, Dominus autem intuetur cor ".
1SAM|16|8|Et vocavit Isai Abinadab et adduxit eum coram Samuele, qui dixit: " Nec hunc elegit Dominus ".
1SAM|16|9|Adduxit autem Isai Samma, de quo ait: " Etiam hunc non elegit Dominus ".
1SAM|16|10|Adduxit itaque Isai septem filios suos coram Samuele, et ait Samuel ad Isai: " Non elegit Dominus ex istis ".
1SAM|16|11|Dixitque Samuel ad Isai: " Numquid iam completi sunt filii? ". Qui respondit: " Adhuc reliquus est minimus et pascit oves ". Et ait Samuel ad Isai: " Mitte et adduc eum; nec enim discumbemus prius quam huc ille venerit ".
1SAM|16|12|Misit ergo et adduxit eum; erat autem rufus et pulcher aspectu decoraque facie. Et ait Dominus: " Surge, unge eum; ipse est enim ".
1SAM|16|13|Tulit igitur Samuel cornu olei et unxit eum in medio fratrum eius; et directus est spiritus Domini in David a die illa et in reliquum. Surgensque Samuel abiit in Rama.
1SAM|16|14|Spiritus autem Domini recessit a Saul, et exagitabat eum spiritus nequam a Domino.
1SAM|16|15|Dixeruntque servi Saul ad eum: " Ecce spiritus Dei malus exagitat te.
1SAM|16|16|Iubeat dominus noster, et servi tui, qui coram te sunt, quaerant hominem scientem psallere cithara, ut, quando arripuerit te spiritus Dei malus, psallat manu sua, et levius feras ".
1SAM|16|17|Et ait Saul ad servos suos: " Providete mihi aliquem bene psallentem et adducite eum ad me ".
1SAM|16|18|Et respondens unus de pueris ait: " Ecce vidi filium Isai Bethlehemitae scientem psallere et fortissimum robore et virum bellicosum et prudentem in verbis et virum pulchrum; et Dominus est cum eo ".
1SAM|16|19|Misit ergo Saul nuntios ad Isai dicens: " Mitte ad me David filium tuum, qui est in pascuis ".
1SAM|16|20|Tulitque Isai asinum cum pane et utre vini et haedo de capris uno et misit per manum David filii sui Sauli.
1SAM|16|21|Et venit David ad Saul et stetit coram eo; at ille dilexit eum nimis, et factus est eius armiger.
1SAM|16|22|Misitque Saul ad Isai dicens: " Stet David in conspectu meo; invenit enim gratiam in oculis meis ".
1SAM|16|23|Igitur, quandocumque spiritus Dei arripiebat Saul, David tollebat citharam et percutiebat manu sua; et refocillabatur Saul et levius habebat: recedebat enim ab eo spiritus malus.
1SAM|17|1|Congregantes vero Phili sthim agmina sua in proe lium, convenerunt in Socho Iudae et castrametati sunt inter Socho et Azeca in Aphesdommim.
1SAM|17|2|Porro Saul et viri Israel congregati venerunt in vallem Terebinthi et instruxerunt aciem ad pugnandum contra Philisthim.
1SAM|17|3|Et Philisthim stabant super montem ex hac parte, et Israel stabat super montem ex altera parte; vallisque erat inter eos.
1SAM|17|4|Et egressus est vir propugnator de castris Philisthinorum nomine Goliath de Geth altitudinis sex cubitorum et palmi.
1SAM|17|5|Et cassis aerea super caput eius, et lorica squamata induebatur; porro pondus loricae eius quinque milia siclorum aeris.
1SAM|17|6|Et ocreas aereas habebat in cruribus, et acinaces aereus erat inter umeros eius.
1SAM|17|7|Hastile autem hastae eius erat quasi liciatorium texentium, ipsum autem ferrum hastae eius sescentos siclos habebat ferri; et armiger eius antecedebat eum.
1SAM|17|8|Stansque clamabat adversum agmina Israel et dicebat eis: " Quare venitis parati ad proelium? Numquid ego non sum Philisthaeus, et vos servi Saul? Eligite ex vobis virum, et descendat ad singulare certamen!
1SAM|17|9|Si quiverit pugnare mecum et percusserit me, erimus vobis servi; si autem ego praevaluero et percussero eum, vos servi eritis et servietis nobis ".
1SAM|17|10|Et aiebat Philisthaeus: " Ego exprobravi agminibus Israel hodie: Date mihi virum, et ineat mecum singulare certamen! ".
1SAM|17|11|Audiens autem Saul et omnes Israelitae sermones Philisthaei huiuscemodi stupebant et metuebant nimis.
1SAM|17|12|David autem erat filius viri Ephrathaei, de quo supra dictum est, de Bethlehem Iudae, cui erat nomen Isai; qui habebat octo filios et erat vir in diebus Saul senex et grandaevus inter viros.
1SAM|17|13|Abierunt autem tres filii eius maiores post Saul in proelium; et nomina trium filiorum eius, qui perrexerant ad bellum: Eliab primogenitus et secundus Abinadab tertiusque Samma.
1SAM|17|14|David autem erat minimus; tribus ergo maioribus secutis Saulem,
1SAM|17|15|ibat David et revertebatur a Saul, ut pasceret gregem patris sui in Bethlehem.
1SAM|17|16|Procedebat vero Philisthaeus mane et vespere et stabat quadraginta diebus.
1SAM|17|17|Dixit autem Isai ad David filium suum: " Accipe fratribus tuis ephi frumenti tosti et decem panes istos et curre in castra ad fratres tuos.
1SAM|17|18|Et decem formellas casei has deferes ad tribunum, et fratres tuos visitabis, si recte agant; et pignus ab eis referes ".
1SAM|17|19|Saul autem et illi et omnes filii Israel in valle Terebinthi pugnabant adversum Philisthim.
1SAM|17|20|Surrexit itaque David mane et commendavit gregem custodi et onustus abiit, sicut praeceperat ei Isai. Et venit ad carraginem, dum exercitus egrediebatur ad pugnam et vociferabatur in certamine.
1SAM|17|21|Direxerunt ergo Israel et Philisthim aciem adversus aciem.
1SAM|17|22|Derelinquens autem David vasa, quae attulerat, sub manu custodis ad sarcinas, cucurrit ad locum certaminis et interrogabat, si omnia recte agerentur erga fratres suos.
1SAM|17|23|Cumque adhuc ille loqueretur eis, apparuit vir ille propugnator ascendens, Goliath nomine, Philisthaeus de Geth, ex castris Philisthinorum; et loquente eo haec eadem verba, audivit David.
1SAM|17|24|Omnes autem Israelitae, cum vidissent virum, fugerunt a facie eius timentes eum valde.
1SAM|17|25|Et dixit unus quispiam de Israel: " Num vidistis virum hunc, qui ascendit? Ad exprobrandum enim Israeli ascendit. Virum ergo, qui percusserit eum, ditabit rex divitiis magnis et filiam suam dabit ei; et domum patris eius faciet absque tributo in Israel ".
1SAM|17|26|Et ait David ad viros, qui stabant secum, dicens: " Quid dabitur viro, qui percusserit Philisthaeum hunc et tulerit opprobrium de Israel? Quis est enim hic Philisthaeus incircumcisus, qui exprobravit acies Dei viventis? ".
1SAM|17|27|Referebat autem ei populus eundem sermonem dicens: " Haec dabuntur viro, qui percusserit eum ".
1SAM|17|28|Quod cum audisset Eliab frater eius maior, loquente eo cum aliis, iratus est contra David et ait: " Quare venisti et cui dereliquisti pauculas oves illas in deserto? Ego novi superbiam tuam et nequitiam cordis tui, quia ut videres proelium descendisti ".
1SAM|17|29|Et dixit David: " Quid feci? Numquid non verbum est? ".
1SAM|17|30|Et declinavit paululum ab eo ad alium dixitque eundem sermonem; et respondit ei populus verbum sicut prius.
1SAM|17|31|Audita sunt autem verba, quae locutus est David, et annuntiata in conspectu Saul.
1SAM|17|32|Ad quem cum fuisset adductus, locutus est ei: " Non concidat cor cuiusquam in eo; ego servus tuus vadam et pugnabo adversus Philisthaeum istum ".
1SAM|17|33|Et ait Saul ad David: " Non vales resistere Philisthaeo isti nec pugnare adversus eum, quia puer es; hic autem vir bellator ab adulescentia sua ".
1SAM|17|34|Dixitque David ad Saul: " Pascebat servus tuus patris sui gregem, et veniebat leo vel ursus tollebatque arietem de medio gregis.
1SAM|17|35|Et sequebar eos et percutiebam eruebamque de ore eorum; et illi consurgebant adversum me, et apprehendebam mentum eorum et percutiebam interficiebamque eos.
1SAM|17|36|Nam et leonem et ursum interfecit servus tuus; erit igitur et Philisthaeus hic incircumcisus quasi unus ex eis, quia ausus est maledicere exercitum Dei viventis ".
1SAM|17|37|Et ait David: " Dominus, qui eruit me de manu leonis et de manu ursi, ipse liberabit me de manu Philisthaei huius ". Dixit autem Saul ad David: Vade, et Dominus tecum sit ".
1SAM|17|38|Et induit Saul David vestimentis suis et imposuit galeam aeream super caput eius et vestivit eum lorica.
1SAM|17|39|Accinctus ergo David gladio eius super vestem suam coepit tentare, si armatus posset incedere; non enim habebat consuetudinem. Dixitque David ad Saul: " Non possum sic incedere, quia nec usum habeo ". Et deposuit ea
1SAM|17|40|et tulit baculum suum in manu sua; et elegit sibi quinque levissimos lapides de torrente et misit eos in peram pastoralem, qua ut sacculo lapidum utebatur, et fundam manu tulit et processit adversum Philisthaeum.
1SAM|17|41|Ibat autem Philisthaeus incedens et appropinquans adversum David, et armiger eius ante eum.
1SAM|17|42|Cumque inspexisset Philisthaeus et vidisset David, despexit eum; erat enim adulescens rufus et pulcher aspectu.
1SAM|17|43|Et dixit Philisthaeus ad David: " Numquid ego canis sum, quod tu venis ad me cum baculo? ". Et maledixit Philisthaeus David in diis suis;
1SAM|17|44|dixitque ad David: " Veni ad me, et dabo carnes tuas volatilibus caeli et bestiis terrae ".
1SAM|17|45|Dixit autem David ad Philisthaeum: " Tu venis ad me cum gladio et hasta et acinace; ego autem venio ad te in nomine Domini exercituum, Dei agminum Israel, quibus exprobrasti.
1SAM|17|46|Hodie dabit te Dominus in manu mea, et percutiam te et auferam caput tuum a te; et dabo cadaver tuum et cadavera castrorum Philisthim hodie volatilibus caeli et bestiis terrae, ut sciat omnis terra quia est Deus in Israel,
1SAM|17|47|et noverit universa ecclesia haec quia non in gladio nec in hasta salvat Dominus: ipsius enim est bellum, et tradet vos in manus nostras ".
1SAM|17|48|Cum ergo surrexisset Philisthaeus et veniret et appropinquaret contra David, festinavit David et cucurrit ad pugnam adversum Philisthaeum.
1SAM|17|49|Et misit manum suam in peram tulitque unum lapidem et funda iecit; et percussit Philisthaeum in fronte, et infixus est lapis in fronte eius, et cecidit in faciem suam super terram.
1SAM|17|50|Praevaluitque David adversum Philisthaeum in funda et in lapide; percussumque Philisthaeum interfecit. Cumque gladium non haberet in manu, David
1SAM|17|51|cucurrit et stetit super Philisthaeum; et tulit gladium eius et eduxit eum de vagina sua et interfecit eum praeciditque caput eius.Videntes autem Philisthim quod mortuus esset fortissimus eorum fugerunt.
1SAM|17|52|Et consurgentes viri Israel et Iudae vociferati sunt et persecuti Philisthaeos usque dum venirent ad Geth et usque ad portas Accaron. Cecideruntque vulnerati de Philisthim in via a Saarim usque ad Geth et usque ad Accaron.
1SAM|17|53|Et revertentes filii Israel, postquam persecuti fuerant Philisthaeos, praedati sunt castra eorum.
1SAM|17|54|Assumens autem David caput Philisthaei attulit illud in Ierusalem; arma vero eius posuit in tabernaculo.
1SAM|17|55|Eo autem tempore, quo viderat Saul David egredientem contra Philisthaeum, ait ad Abner principem militiae: " De qua stirpe descendit hic adulescens, Abner? ". Dixitque Abner: " Vivit anima tua, rex, quia non novi ".
1SAM|17|56|Et ait rex: " Interroga tu, cuius filius sit iste puer ".
1SAM|17|57|Cumque regressus esset David, percusso Philisthaeo, tulit eum Abner et introduxit coram Saul caput Philisthaei habentem in manu.
1SAM|17|58|Et ait ad eum Saul: " De qua progenie es, o adulescens? ". Dixitque David: " Filius servi tui Isai Bethlehemitae ego sum ".
1SAM|18|1|Et factum est cum complesset loqui ad Saul, anima Ionathan colligata est animae David, et dilexit eum Ionathan quasi animam suam.
1SAM|18|2|Tulitque eum Saul in die illa et non concessit ei, ut reverteretur in domum patris sui.
1SAM|18|3|Inierunt autem Ionathan et David foedus; diligebat enim eum quasi animam suam.
1SAM|18|4|Et exspoliavit se Ionathan tunicam, qua erat vestitus, et dedit eam David et reliqua vestimenta sua usque ad gladium et arcum suum et usque ad balteum.
1SAM|18|5|Egrediebatur quoque David ad omnia, quaecumque misisset eum Saul, et prospere agebat; posuitque eum Saul super viros belli, et acceptus erat in oculis universi populi, etiam in conspectu famulorum Saul.
1SAM|18|6|Porro cum reverterentur, cum rediret David, percusso Philisthaeo, egressae sunt mulieres de universis urbibus Israel cantantes chorosque ducentes in occursum Saul regis in tympanis et in canticis laetitiae et in sistris.
1SAM|18|7|Et praecinebant mulieres ludentes atque dicentes: Percussit Saul milia sua,et David decem milia sua ".
1SAM|18|8|Iratus est autem Saul nimis, et displicuit in oculis eius iste sermo, dixitque: " Dederunt David decem milia et mihi dederunt milia; quid ei superest nisi solum regnum? ".
1SAM|18|9|Non rectis ergo oculis Saul aspiciebat David ex die illa et deinceps.
1SAM|18|10|Post diem autem alteram invasit spiritus Dei malus Saul, et vaticinabatur in medio domus suae; David autem psallebat manu sua sicut per singulos dies, tenebatque Saul lanceam.
1SAM|18|11|Et sustulit eam putans quod configere posset David cum pariete; et declinavit David a facie eius secundo.
1SAM|18|12|Et timuit Saul David, eo quod esset Dominus cum eo et a se recessisset.
1SAM|18|13|Amovit ergo eum Saul a se et fecit eum tribunum super mille viros; et egrediebatur et intrabat in conspectu populi.
1SAM|18|14|In omnibus quoque viis suis David prospere agebat, et Dominus erat cum eo.
1SAM|18|15|Vidit itaque Saul quod prospere ageret nimis et coepit pavere eum;
1SAM|18|16|omnis autem Israel et Iuda diligebat David; ipse enim egrediebatur et ingrediebatur ante eos.
1SAM|18|17|Dixit autem Saul ad David: " Ecce filia mea maior Merob, ipsam dabo tibi uxorem; tantummodo esto mihi vir fortis et proeliare bella Domini ". Saul autem reputabat dicens: " Non sit manus mea in eo, sed sit super illum manus Philisthinorum ".
1SAM|18|18|Ait autem David ad Saul: " Quis ego sum, aut quae est vita mea aut cognatio patris mei in Israel, ut fiam gener regis? ".
1SAM|18|19|Factum est autem tempus, cum deberet dari Merob filia Saul David, data est Hadriel Molathitae uxor.
1SAM|18|20|Dilexit autem Michol filia Saul altera David, et nuntiatum est Saul, et placuit ei;
1SAM|18|21|dixitque Saul: " Dabo eam illi, ut fiat ei in scandalum, et sit super eum manus Philisthinorum ". Dixit ergo Saul ad David altera vice: " Gener meus eris hodie ".
1SAM|18|22|Et mandavit Saul servis suis: " Loquimini ad David secreto dicentes: Ecce places regi, et omnes servi eius diligunt te; nunc ergo esto gener regis" ".
1SAM|18|23|Et locuti sunt servi Saul in auribus David omnia verba haec, et ait David: " Num parum vobis videtur generum esse regis? Ego autem sum vir pauper et tenuis ".
1SAM|18|24|Et renuntiaverunt servi Saul dicentes: " Huiuscemodi verba locutus est David ".
1SAM|18|25|Dixit autem Saul: " Sic loquimini ad David: "Non habet necesse rex sponsalia, nisi tantum centum praeputia Philisthinorum, ut fiat ultio de inimicis regis" ". Porro Saul cogitabat tradere David in manibus Philisthinorum.
1SAM|18|26|Cumque renuntiassent servi eius David verba, quae dixerat Saul, placuit sermo in oculis David, ut fieret gener regis.
1SAM|18|27|Et nondum erant dies impleti, cum David surgens abiit cum viris, qui sub eo erant, et percussit ex Philisthim ducentos viros; et attulit praeputia eorum, et annumeraverunt ea regi, ut esset gener eius.Dedit itaque ei Saul Michol filiam suam uxorem.
1SAM|18|28|Et vidit Saul et intellexit quia Dominus esset cum David; Michol autem filia Saul diligebat eum.
1SAM|18|29|Et Saul magis coepit timere David; factusque est Saul inimicus David cunctis diebus.
1SAM|18|30|Et egressi sunt principes Philisthinorum; et, quotiescumque egrediebantur, prospere agebat David magis quam omnes servi Saul, et celebre factum est nomen eius nimis.
1SAM|19|1|Locutus est autem Saul ad Ionathan filium suum et ad omnes servos suos de occisione David; porro Ionathan filius Saul diligebat David valde.
1SAM|19|2|Et indicavit Ionathan David dicens: " Quaerit Saul pater meus occidere te; quapropter observa te, quaeso, mane; et manebis clam et absconderis.
1SAM|19|3|Ego autem egrediens stabo iuxta patrem meum in agro, ubicumque fueris; et ego loquar de te ad patrem meum et, quodcumque videro, nuntiabo tibi ".
1SAM|19|4|Locutus est ergo Ionathan de David bona ad Saul patrem suum dixitque ad eum: " Ne peccet rex in servum suum David, quia non peccavit tibi, et opera eius bona sunt tibi valde.
1SAM|19|5|Et posuit animam suam in manu sua et percussit Philisthaeum, et fecit Dominus victoriam magnam universo Israeli; vidisti et laetatus es. Quare ergo peccas in sanguine innoxio interficiens David, qui est absque culpa?.
1SAM|19|6|Quod cum audisset Saul, placatus voce Ionathan iuravit: " Vivit Dominus quia non occidetur ".
1SAM|19|7|Vocavit itaque Ionathan David et indicavit ei omnia verba haec; et introduxit lonathan David ad Saul, et fuit ante eum, sicut fuerat heri et nudiustertius.
1SAM|19|8|Motum est autem rursum bellum, et egressus David pugnavit adversum Philisthim percussitque eos plaga magna; et fugerunt a facie eius.
1SAM|19|9|Et factus est spiritus Domini malus in Saul; sedebat autem in domo sua et tenebat lanceam, porro David psallebat in manu sua.
1SAM|19|10|Nisusque est Saul configere lancea David in pariete; et declinavit David a facie Saul, lancea autem, casso vulnere, perlata est in parietem. Et David fugit et salvatus est nocte illa.
1SAM|19|11|Misit ergo Saul satellites suos in domum David, ut custodirent eum, et interficeretur mane.Quod cum annuntiasset David Michol uxor sua dicens: " Nisi salvaveris te nocte hac, cras morieris ",
1SAM|19|12|deposuit eum per fenestram. Porro ille abiit et aufugit atque salvatus est.
1SAM|19|13|Tulit autem Michol theraphim et posuit eum super lectum; et pellem pilosam caprarum posuit ad caput eius et operuit eum vestimentis.
1SAM|19|14|Misit autem Saul nuntios, qui raperent David, et responsum est quod aegrotaret.
1SAM|19|15|Rursumque misit Saul nuntios, ut viderent David, dicens: " Afferte eum ad me in lecto, ut occidatur ".
1SAM|19|16|Cumque venissent nuntii, inventus est theraphim super lectum, et pellis caprarum ad caput eius.
1SAM|19|17|Dixitque Saul ad Michol: " Quare sic illusisti mihi et dimisisti inimicum meum, ut fugeret? ". Et respondit Michol ad Saul: " Quia ipse locutus est mihi: "Dimitte me, alioquin interficiam te" ".
1SAM|19|18|David autem fugiens salvatus est et venit ad Samuel in Rama et nuntiavit ei omnia, quae fecerat sibi Saul. Et abierunt ipse et Samuel et morati sunt in Naioth.
1SAM|19|19|Nuntiatum est autem Sauli a dicentibus: " Ecce David in Naioth in Rama.
1SAM|19|20|Misit ergo Saul nuntios, ut raperent David. Qui cum vidissent cuneum prophetarum vaticinantium et Samuel stantem super eos, factus est in illis spiritus Dei, et vaticinari coeperunt etiam ipsi.
1SAM|19|21|Quod cum nuntiatum esset Sauli, misit alios nuntios; vaticinati sunt autem et illi. Et rursum Saul misit tertios nuntios, qui et ipsi vaticinati sunt.
1SAM|19|22|Abiit autem etiam ipse in Rama et venit usque ad cisternam magnam, quae est in Socho; et interrogavit et dixit: " In quo loco sunt Samuel et David? ". Dictumque est ei: " Ecce in Naioth sunt in Rama ".
1SAM|19|23|Et abiit inde in Naioth in Rama; et factus est etiam super eum spiritus Dei, et ambulabat ingrediens et vaticinans, usquedum veniret in Naioth in Rama.
1SAM|19|24|Et exspoliavit se etiam ipse vestimentis suis et vaticinatus est cum ceteris coram Samuel; et cecidit nudus tota die illa et nocte, unde et exivit proverbium: " Num et Saul inter prophetas? ".
1SAM|20|1|Fugit autem David de Naioth, quae est in Rama, veniensque locutus est coram Ionathan: " Quid feci? Quae est iniquitas mea et quod peccatum meum in patrem tuum, quia quaerit animam meam? ".
1SAM|20|2|Qui dixit ei: " Absit, non morieris; neque enim faciet pater meus quidquam grande vel parvum, nisi prius indicaverit mihi; hoc ergo celavit me pater meus tantummodo? Nequaquam erit istud ".
1SAM|20|3|Et rursum respondit David et ait: " Scit profecto pater tuus quia inveni gratiam in oculis tuis et dixit: "Nesciat hoc Ionathan, ne forte tristetur". Quinimmo vivit Dominus, et vivit anima tua, quia uno tantum gradu ego morsque dividimur ".
1SAM|20|4|Et ait Ionathan ad David: " Quid desiderat anima tua, ut faciam tibi? ".
1SAM|20|5|Dixit autem David ad Ionathan: " Ecce neomenia est crastino, et ego ex more sedere soleo iuxta regem ad vescendum; dimitte ergo me, ut abscondar in agro usque ad vesperam diei tertiae.
1SAM|20|6|Si requisierit me pater tuus, respondebis ei: "Rogavit me David, ut iret celeriter in Bethlehem civitatem suam, quia victimae annuae ibi sunt universis contribulibus eius".
1SAM|20|7|Si dixerit: "Bene", pax erit servo tuo; si autem fuerit iratus, scito quia malum decretum est ab eo.
1SAM|20|8|Fac ergo misericordiam in servum tuum, quia foedus Domini me famulum tuum tecum inire fecisti; si autem est in me aliqua iniquitas, tu me interfice et ad patrem tuum ne introducas me ".
1SAM|20|9|Et ait Ionathan: " Absit hoc a te; neque enim fieri potest ut, si certo cognovero malum decretum esse a patre meo contra te, non annuntiem tibi ".
1SAM|20|10|Responditque David ad Ionathan: " Quis nuntiabit mihi, si quid forte responderit tibi pater tuus dure? ".
1SAM|20|11|Et ait Ionathan ad David: " Veni, egrediamur foras in agrum ". Cumque exissent ambo in agrum,
1SAM|20|12|ait Ionathan ad David: " Vivit Dominus, Deus Israel, investigabo sententiam patris mei hoc fere tempore cras vel perendie; et si aliquid boni fuerit super David, et non statim miserim ad te et notum tibi fecerim,
1SAM|20|13|haec faciat Dominus in Ionathan et haec augeat! Si autem perseveraverit patris mei malitia adversum te, hoc quoque notum faciam tibi et dimittam te, ut vadas in pace. Et sit Dominus tecum, sicut fuit cum patre meo.
1SAM|20|14|Et, si vixero, facies mihi misericordiam Domini; si vero mortuus fuero,
1SAM|20|15|non auferas misericordiam tuam a domo mea usque in sempiternum, quando eradicaverit Dominus inimicos David unumquemque de terra ".
1SAM|20|16|Pepigit ergo foedus Ionathan cum domo David dicens: " Requirat Dominus de manu inimicorum David! ".
1SAM|20|17|Et addidit Ionathan ut faceret David iurare per dilectionem suam erga illum; sicut animam enim suam, ita diligebat eum.
1SAM|20|18|Dixitque ad eum Ionathan: " Cras neomenia est, et requireris;
1SAM|20|19|vacua erit enim sessio tua. Perendie descendes festinus et venies in locum, ubi abscondisti te in die facti illius; et sedebis iuxta acervum illum.
1SAM|20|20|Et ego tres sagittas mittam iuxta eum et iaciam quasi exercens me ad signum.
1SAM|20|21|Mittam quoque et puerum dicens ei: "Vade et affer mihi sagittas".
1SAM|20|22|Si dixero puero: "Ecce sagittae intra te sunt, tolle eas", tu veni ad me, quia pax tibi est, et nihil est mali, vivit Dominus. Si autem sic locutus fuero puero: "Ecce sagittae ultra te sunt", vade, quia dimisit te Dominus.
1SAM|20|23|De verbo autem, quod locuti fuimus, ego et tu, sit Dominus inter me et te usque in sempiternum ".
1SAM|20|24|Absconditus est ergo David in agro; et venit neomenia, et sedit rex ad mensam ad comedendum.
1SAM|20|25|Cumque sedisset rex super cathedram suam secundum consuetudinem, quae erat iuxta parietem, sedit Ionathan ex adverso, et sedit Abner ex latere Saul; vacuusque apparuit locus David.
1SAM|20|26|Et non est locutus Saul quidquam in die illa; cogitabat enim quod forte evenisset ei, ut non esset mundus nec purificatus.
1SAM|20|27|Cumque illuxisset dies secunda post neomeniam, rursum vacuus apparuit locus David; dixitque Saul ad Ionathan filium suum: " Cur non venit filius Isai nec heri nec hodie ad vescendum? ".
1SAM|20|28|Et respondit Ionathan Sauli: " Rogavit me obnixe, ut iret in Bethlehem,
1SAM|20|29|et ait: "Dimitte me, quoniam sacrificium familiae est in civitate, et frater meus ipse accersivit me; nunc ergo, si inveni gratiam in oculis tuis, vadam cito et videbo fratres meos". Ob hanc causam non venit ad mensam regis ".
1SAM|20|30|Iratus autem Saul adversum Ionathan dixit ei: " Fili mulieris perversae, numquid ignoro quia diligis filium Isai in confusionem tuam et in confusionem nuditatis matris tuae?
1SAM|20|31|Omnibus enim diebus, quibus filius Isai vixerit super terram, non stabilieris tu neque regnum tuum; itaque iam nunc mitte et adduc eum ad me, quia filius mortis est ".
1SAM|20|32|Respondens autem Ionathan Sauli patri suo ait: " Quare morietur? Quid fecit? ".
1SAM|20|33|Et arripuit Saul lanceam, ut percuteret eum; et intellexit Ionathan quod definitum esset patri suo, ut interficeret David.
1SAM|20|34|Surrexit ergo Ionathan a mensa in ira furoris et non comedit in die neomeniae secunda panem; contristatus est enim super David, eo quod confudisset eum pater suus.
1SAM|20|35|Cumque illuxisset mane, venit Ionathan in agrum ad locum constitutum a David et puer parvulus cum eo;
1SAM|20|36|et ait ad puerum suum: " Vade et affer mihi sagittas, quas ego iacio ". Cumque puer cucurrisset, iecit sagittam trans puerum.
1SAM|20|37|Venit itaque puer ad locum sagittae, quam miserat Ionathan, et clamavit Ionathan post tergum pueri et ait: " Ecce ibi est sagitta porro ultra te.
1SAM|20|38|Clamavitque Ionathan post tergum pueri: " Festina velociter, ne steteris ". Sustulit autem puer Ionathae sagittam et attulit ad dominum suum
1SAM|20|39|et quid ageretur penitus ignorabat, tantummodo enim Ionathan et David rem noverant.
1SAM|20|40|Dedit igitur Ionathan arma sua puero et dixit ei: " Vade, defer in civitatem ".
1SAM|20|41|Cumque abisset puer, surrexit David de latere acervi et cadens pronus in terram adoravit tertio; et osculantes alterutrum fleverunt pariter, David autem amplius.
1SAM|20|42|Dixit ergo Ionathan ad David: " Vade in pace; iuravimus enim ambo in nomine Domini dicentes: Dominus erit inter me et te et inter semen meum et semen tuum usque in sempiternum ".
1SAM|21|1|Et surrexit David et abiit; sed et Ionathan ingressus est civitatem.
1SAM|21|2|Venit autem David in Nob ad Achimelech sacerdotem, et obstupuit Achimelech eo quod venisset David, et dixit ei: " Quare tu solus et nullus est tecum? ".
1SAM|21|3|Et ait David ad Achimelech sacerdotem: " Rex praecepit mihi negotium et dixit: "Nemo sciat rem, propter quam a me missus es, et cuiusmodi tibi praecepta dederim"; pueris vero condixi in illum et illum locum.
1SAM|21|4|Nunc igitur, si habes ad manum quinque panes, da mihi, aut quidquid inveneris ".
1SAM|21|5|Et respondens sacerdos David ait ei: " Non habeo panes laicos ad manum, sed tantum panem sanctum; si mundi sunt pueri maxime a mulieribus? ".
1SAM|21|6|Et respondit David sacerdoti et dixit ei: " Equidem, si de mulieribus agitur, continuimus nos ab heri et nudiustertius. Quando egrediebar, fuerunt corpora puerorum sancta, quamvis iter esset profanum. Quanto magis hodie sunt sancti quoad corpora ".
1SAM|21|7|Dedit ergo ei sacerdos sanctificatum panem; neque enim erat ibi panis, nisi tantum panes propositionis, qui sublati fuerant a facie Domini, ut ponerentur panes calidi.
1SAM|21|8|Erat autem ibi vir de servis Saul in die illa retentus ante Dominum; et nomen eius Doeg Idumaeus, potentissimus pastorum Saul.
1SAM|21|9|Dixit autem David ad Achimelech: " Si habes hic ad manum hastam aut gladium? Quia gladium meum et arma mea non tuli mecum; negotium enim regis urgebat ".
1SAM|21|10|Et dixit sacerdos: " Ecce hic gladius Goliath Philisthaei, quem percussisti in valle Terebinthi; est involutus pallio post ephod. Si istum vis tollere, tolle, neque enim est alius hic absque eo ". Et ait David: " Non est huic alter similis; da mihi eum ".
1SAM|21|11|Surrexit itaque David et fugit in die illa a facie Saul et venit ad Achis regem Geth.
1SAM|21|12|Dixeruntque ei servi Achis: " Numquid non iste est David rex terrae? Nonne huic cantabant per choros dicentes: "Percussit Saul milia sua, et David decem milia sua"? ".
1SAM|21|13|Posuit autem David sermones istos in corde suo et extimuit valde a facie Achis regis Geth.
1SAM|21|14|Et immutavit os suum coram eis; et insaniebat inter manus eorum et impingebat in ostia portae, defluebantque salivae in barbam.
1SAM|21|15|Et ait Achis ad servos suos: " Vidistis hominem insanum. Quare adduxistis eum ad me?
1SAM|21|16|An desunt nobis furiosi, quod introduxistis istum, ut fureret, me praesente? Hicine ingredietur domum meam? ".
1SAM|22|1|Abiit ergo inde David et fugit in speluncam Odollam; quod cum audissent fratres eius et omnis domus patris eius, descenderunt ad eum illuc.
1SAM|22|2|Et convenerunt ad eum omnes, qui erant in angustia constituti et oppressi aere alieno et amaro animo; et factus est eorum princeps, fueruntque cum eo quasi quadringenti viri.
1SAM|22|3|Et profectus est David inde in Maspha, quae est Moab, et dixit ad regem Moab: " Maneat, oro, pater meus et mater mea vobiscum, donec sciam quid faciat mihi Deus ".
1SAM|22|4|Et reliquit eos ante faciem regis Moab; manseruntque apud eum cunctis diebus, quibus David fuit in praesidio.
1SAM|22|5|Dixitquc Gad propheta ad David: " Noli manere in praesidio. Proficiscere et vade in terram Iudae ". Et profectus David venit in saltum Haret.
1SAM|22|6|Et audivit Saul quod detectus fuisset David et viri, qui erant cum eo. Saul autem, cum maneret in Gabaa et esset sub myrice, quae est in excelso, hastam manu tenens, cunctique servi eius circumstarent eum,
1SAM|22|7|ait ad servos suos, qui assistebant ei: " Audite, Beniaminitae. Etiam omnibus vobis dabit filius Isai agros et vineas et universos vos faciet tribunos et centuriones,
1SAM|22|8|quoniam coniurastis omnes adversum me. Et non est qui mihi renuntiet quod filius meus foedus iunxerit cum filio Isai; non est qui vicem meam doleat ex vobis, nec qui annuntiet mihi quod suscitaverit filius meus servum meum adversum me insidiantem mihi sicut hodie ".
1SAM|22|9|Respondens autem Doeg Idumaeus, qui assistebat cum servis Saul: " Vidi, inquit, filium Isai in Nob apud Achimelech filium Achitob;
1SAM|22|10|qui consuluit pro eo Dominum et cibaria dedit ei, sed et gladium Goliath Philisthaei dedit illi ".
1SAM|22|11|Misit ergo rex ad accersendum Achimelech sacerdotem filium Achitob et omnem domum patris eius, sacerdotum, qui erant in Nob; qui venerunt universi ad regem.
1SAM|22|12|Et ait Saul: " Audi, fili Achitob ". Qui respondit: " Praesto sum, domine ".
1SAM|22|13|Dixitque ad eum Saul: " Quare coniurastis adversum me, tu et filius Isai, et dedisti ei panes et gladium et consuluisti pro eo Deum, ut consurgeret adversum me insidiator, sicut est hodie? ".
1SAM|22|14|Respondensque Achimelech regi ait: " Et quis in omnibus servis tuis sicut David fidelis et gener regis et dux satellitum tuorum et gloriosus in domo tua?
1SAM|22|15|Num hodie coepi consulere pro eo Deum? Absit hoc a me, ne suspicetur rex adversus servum suum rem huiuscemodi, adversus universam domum patris mei; non enim scivit servus tuus quidquam super hoc negotio, vel modicum vel grande ".
1SAM|22|16|Dixitque rex: " Morte morieris, Achimelech, tu et omnis domus patris tui ".
1SAM|22|17|Et ait rex emissariis, qui circumstabant eum: " Convertimini et interficite sacerdotes Domini, nam manus eorum cum David est; scientes quod fugisset, non indicaverunt mihi ". Noluerunt autem servi regis extendere manum suam in sacerdotes Domini.
1SAM|22|18|Et ait rex ad Doeg: " Convertere tu et irrue in sacerdotes ". Conversusque Doeg Idumaeus irruit in sacerdotes; et trucidavit in die illa octoginta quinque viros vestitos ephod lineo.
1SAM|22|19|Nob autem civitatem sacerdotum percussit in ore gladii, viros et mulieres, parvulos et lactantes, bovem et asinum et ovem in ore gladii.
1SAM|22|20|Evadens autem unus filius Achimelech filii Achitob, cuius nomen erat Abiathar, fugit ad David
1SAM|22|21|et annuntiavit ei quod occidisset Saul sacerdotes Domini.
1SAM|22|22|Et ait David ad Abiathar: " Sciebam in die illa quod, cum ibi esset Doeg Idumaeus, procul dubio annuntiaret Saul; ego sum reus omnium animarum domus patris tui.
1SAM|22|23|Mane mecum, ne timeas; qui enim quaerit animam meam, quaerit et animam tuam, mecumque servaberis ".
1SAM|23|1|Et nuntiaverunt David di centes: " Ecce Philisthim op pugnant Ceila et diripiunt areas ".
1SAM|23|2|Consuluit igitur David Dominum dicens: " Num vadam et percutiam Philisthaeos istos? ". Et ait Dominus ad David: " Vade et percuties Philisthaeos et salvabis Ceila ".
1SAM|23|3|Et dixerunt viri, qui erant cum David, ad eum: " Ecce nos hic in Iuda consistentes timemus; quanto magis si ierimus in Ceila adversum agmina Philisthinorum? ".
1SAM|23|4|Rursum ergo David consuluit Dominum, qui respondens ei ait: " Surge et vade in Ceila; ego enim tradam Philisthaeos in manu tua ".
1SAM|23|5|Abiit ergo David et viri eius in Ceila et pugnavit adversum Philisthaeos et abegit iumenta eorum et percussit eos plaga magna: et salvavit David habitatores Ceilae.
1SAM|23|6|Porro cum fugisset Abiathar filius Achimelcch ad David, et ipse cum David in Ceila ephod secum habens descenderat.
1SAM|23|7|Nuntiatum est autem Saul quod venisset David in Ceila, et ait Saul: " Tradidit eum Deus in manus meas; conclususque est introgressus urbem, in qua portae et serae sunt ".
1SAM|23|8|Et convocavit Saul omnem populum, ut ad pugnam descenderet in Ceila et obsideret David et viros eius.
1SAM|23|9|Quod cum rescisset David quia praepararet ei Saul clam malum, dixit ad Abiathar sacerdotem: " Applica ephod ".
1SAM|23|10|Et ait David: " Domine, Deus Israel, audivit famam servus tuus quod disponat Saul venire ad Ceila, ut evertat urbem propter me.
1SAM|23|11|Si tradent me viri Ceilae in manus eius? Et si descendet Saul, sicut audivit servus tuus? Domine, Deus Israel, indica servo tuo ". Et ait Dominus: " Descendet ".
1SAM|23|12|Dixitque David: " Si tradent viri Ceilae me et viros, qui sunt mecum, in manu Saul? ". Et dixit Dominus: " Tradent ".
1SAM|23|13|Surrexit ergo David et viri eius quasi sescenti et egressi de Ceila huc atque illuc vagabantur incerti. Nuntiatumque est Saul quod fugisset David de Ceila, quam ob rem destitit exire.
1SAM|23|14|Morabatur autem David in deserto in locis firmissimis mansitque in monte, in deserto Ziph; et quaerebat eum Saul cunctis diebus, sed non tradidit eum Deus in manus eius.
1SAM|23|15|Et cognovit David quod egressus esset Saul, ut quaereret animam eius; porro David erat in deserto Ziph in Horesa.
1SAM|23|16|Et surrexit Ionathan filius Saul et abiit ad David in Horesa; et confortavit manus eius in Deo dixitque ei:
1SAM|23|17|" Ne timeas, neque enim inveniet te manus Saul patris mei; et tu regnabis super Israel, et ego ero tibi secundus; sed et Saul pater meus scit hoc ".
1SAM|23|18|Percussit igitur uterque foedus coram Domino; mansitque David in Horesa, Ionathan autem reversus est in domum suam.
1SAM|23|19|Ascenderunt autem Ziphaei ad Saul in Gabaa dicentes: " Nonne David latitat apud nos in locis tutissimis in Horesa, in colle Hachila, quae est ad meridiem deserti?
1SAM|23|20|Nunc ergo, si desideravit anima tua, rex, ut descenderes, descende; nostrum autem erit ut tradamus eum in manus regis ".
1SAM|23|21|Dixitque Saul: " Benedicti vos a Domino, quia doluistis vicem meam.
1SAM|23|22|Abite, oro, et diligentius praeparate et curiosius agite; et considerate locum, ubi sit pes eius, vel quis viderit eum ibi; dictum est enim ad me quod callidus sit valde.
1SAM|23|23|Considerate et videte omnia latibula eius, in quibus absconditur, et revertimini ad me ad certum locum, ut vadam vobiscum; quodsi fuerit in regione, perscrutabor eum in cunctis regionibus Iudae ".
1SAM|23|24|At illi surgentes abierunt in Ziph ante Saul.David autem et viri eius erant in deserto Maon, in Araba ad meridiem deserti.
1SAM|23|25|Ivit ergo Saul et socii eius ad quaerendum eum, et nuntiatum est David; descenditque ad petram et versabatur in deserto Maon. Quod cum audisset Saul, persecutus est David in deserto Maon.
1SAM|23|26|Et ibat Saul ad latus montis ex parte una, David autem et viri eius erant in latere montis ex parte altera; porro David praeceps fugiebat a facie Saul. Itaque Saul et viri eius in modum coronae cingebant David et viros eius, ut caperent eos.
1SAM|23|27|Et nuntius venit ad Saul dicens: " Festina et veni, quoniam infuderunt se Philisthim super terram ".
1SAM|23|28|Reversus est ergo Saul desistens persequi David; et perrexit in occursum Philisthinorum. Propter hoc vocaverunt locum illum: " Petram dividentem ".
1SAM|24|1|Ascendit ergo David inde et habitavit in locis tutissimis Engaddi.
1SAM|24|2|Cumque reversus esset Saul, postquam persecutus est Philisthaeos, nuntiaverunt ei dicentes: " Ecce David in deserto est Engaddi ".
1SAM|24|3|Assumens ergo Saul tria milia electorum virorum ex omni Israel perrexit ad investigandum David et viros eius ad rupes ibicum.
1SAM|24|4|Et venit ad caulas ovium, quae se offerebant vianti.Eratque ibi spelunca, quam ingressus est Saul, ut purgaret ventrem; porro David et viri eius in interiore parte speluncae latebant.
1SAM|24|5|Et dixerunt viri David ad eum: " Ecce dies, de qua locutus est Dominus ad te: "Ego trado tibi inimicum tuum, ut facias ei sicut placuerit in oculis tuis" ". Surrexit ergo David et praecidit oram chlamydis Saul silenter.
1SAM|24|6|Post haec cor David percussit eum, eo quod abscidisset oram chlamydis Saul,
1SAM|24|7|dixitque ad viros suos: " Propitius mihi sit Dominus, ne faciam hanc rem domino meo, christo Domini, ut mittam manum meam in eum, quoniam christus Domini est ".
1SAM|24|8|Et cohibuit David viros suos sermonibus et non permisit eos, ut consurgerent in Saul.Porro Saul exsurgens de spelunca pergebat coepto itinere.
1SAM|24|9|Surrexit autem et David post eum et egressus de spelunca clamavit post tergum Saul dicens: " Domine mi rex! ". Et respexit Saul post se, et inclinans se David pronus in terram adoravit
1SAM|24|10|dixitque ad Saul: " Quare audis verba hominum loquentium: "David quaerit malum adversum te?".
1SAM|24|11|Ecce hodie viderunt oculi tui quod tradiderit te Dominus hodie in manu mea in spelunca; et dictum est mihi, ut occiderem te, sed pepercit tibi oculus meus. Dixi enim: Non extendam manum meam in dominum meum, quia christus Domini est
1SAM|24|12|et pater meus. Quin potius vide et cognosce oram chlamydis tuae in manu mea, quoniam, cum praeciderem summitatem chlamydis tuae, nolui occidere te. Animadverte et vide quoniam non est in manu mea malum neque iniquitas, neque peccavi in te; tu autem insidiaris animae meae, ut auferas eam.
1SAM|24|13|Iudicet Dominus inter me et te et ulciscatur me Dominus ex te; manus autem mea non sit in te.
1SAM|24|14|Sicut et in proverbio antiquo dicitur: "Ab impiis egredietur impietas", manus ergo mea non sit in te.
1SAM|24|15|Quem sequitur rex Israel? Quem persequeris? Canem mortuum et pulicem unum.
1SAM|24|16|Sit Dominus iudex et iudicet inter me et te et videat et diiudicet causam meam et eruat me de manu tua ".
1SAM|24|17|Cum autem complesset David loquens sermones huiuscemodi ad Saul, dixit Saul: " Numquid vox haec tua est, fili mi David? ". Et levavit Saul vocem suam et flevit.
1SAM|24|18|Dixitque ad David: " Iustior tu es quam ego; tu enim tribuisti mihi bona, ego autem reddidi tibi mala.
1SAM|24|19|Et tu indicasti hodie, quae feceris mihi bona, quomodo tradiderit me Dominus in manu tua, et non occideris me.
1SAM|24|20|Quis enim, cum invenerit inimicum suum, dimittet eum in via bona? Sed Dominus reddat tibi vicissitudinem hanc, pro eo quod hodie operatus es in me.
1SAM|24|21|Et nunc, quia scio quod certissime regnaturus sis et habiturus in manu tua regnum Israel,
1SAM|24|22|iura mihi in Domino, ne deleas semen meum post me neque auferas nomen meum de domo patris mei ".
1SAM|24|23|Et iuravit David Sauli. Abiit ergo Saul in domum suam, et David et viri eius ascenderunt ad praesidium.
1SAM|25|1|Mortuus est autem Samuel; et congregatus est universus Israel, et planxerunt eum et sepelierunt eum in domo sua in Rama.Consurgensque David descendit in desertum Maon.
1SAM|25|2|Erat autem vir quispiam in solitudine Maon, et possessio eius in Carmel; et homo ille magnus nimis; erantque ei oves tria milia et mille caprae. Et accidit ut tonderet gregem suum in Carmel.
1SAM|25|3|Nomen autem viri illius erat Nabal et nomen uxoris eius Abigail. Eratque mulier illa prudentissima et speciosa; porro vir eius durus et moribus malis; erat autem de genere Chaleb.
1SAM|25|4|Cum ergo audisset David in deserto quod tonderet Nabal gregem suum,
1SAM|25|5|misit decem iuvenes et dixit eis: " Ascendite in Carmel et venietis ad Nabal et salutabitis eum ex nomine meo pacifice
1SAM|25|6|et dicetis fratri meo: "Et tibi pax et domui tuae pax et omnibus, quaecumque habes, sit pax!
1SAM|25|7|Et nunc audivi quod tonsores essent apud te. Pastores autem tui erant nobiscum in deserto; numquam eis molesti fuimus, nec aliquando defuit eis quidquam de grege omni tempore, quo fuerunt nobiscum in Carmel.
1SAM|25|8|Interroga pueros tuos, et indicabunt tibi. Nunc ergo inveniant pueri isti gratiam in oculis tuis, in die enim bona venimus; quodcumque invenerit manus tua, da servis tuis et filio tuo David" ".
1SAM|25|9|Cumque venissent pueri David, locuti sunt ad Nabal omnia verba haec ex nomine David et siluerunt.
1SAM|25|10|Respondens autem Nabal pueris David ait: " Quis est David, et quis est filius Isai? Hodie increverunt servi, qui fugiunt dominos suos.
1SAM|25|11|Tollam ergo panes meos et aquas meas et carnes pecorum, quae occidi, tonsoribus meis et dabo viris, quos nescio unde sint? ".
1SAM|25|12|Regressi sunt itaque pueri David per viam suam et reversi venerunt et nuntiaverunt ei omnia verba haec.
1SAM|25|13|Tunc David ait viris suis: " Accingatur unusquisque gladio suo! ". Et accincti sunt singuli gladio suo, accinctusque est et David ense suo, et secuti sunt David quasi quadringenti viri; porro ducenti remanserunt ad sarcinas.
1SAM|25|14|Abigail autem uxori Nabal nuntiavit unus de pueris suis dicens: " Ecce misit David nuntios de deserto, ut benedicerent domino nostro, sed aversatus est eos.
1SAM|25|15|Homines isti boni satis fuerunt nobis et non molesti; nec quidquam aliquando periit omni tempore, quo sumus conversati cum eis in deserto.
1SAM|25|16|Pro muro erant nobis tam in nocte quam in die omnibus diebus, quibus pavimus apud eos greges.
1SAM|25|17|Quam ob rem considera et recogita quid facias, quoniam malum decretum est adversus dominum nostrum et adversus domum eius universam. Et ipse filius Belial est, ita ut nemo ei possit loqui ".
1SAM|25|18|Festinavit igitur Abigail et tulit ducentos panes et duos utres vini et quinque arietes coctos et quinque sata frumenti tosti et centum ligaturas uvae passae et ducentas massas caricarum et imposuit super asinos.
1SAM|25|19|Dixitque pueris suis: " Praecedite me, ecce ego post tergum sequar vos. Viro autem suo Nabal non indicavit.
1SAM|25|20|Cum ergo ascendisset asinum et descenderet in tegmine montis, David et viri eius descendebant in occursum eius; quibus et illa occurrit.
1SAM|25|21|Et aiebat David: " Vere frustra servavi omnia, quae huius erant in deserto, et non periit quidquam de cunctis, quae ad eum pertinebant; et reddidit mihi malum pro bono.
1SAM|25|22|Haec faciat Deus inimicis David et haec addat, si reliquero de omnibus, quae ad eum pertinent, usque mane quidquid masculini sexus ".
1SAM|25|23|Cum autem vidisset Abigail David, festinavit et descendit de asino et procidit coram David super faciem suam et adoravit super terram.
1SAM|25|24|Et cecidit ad pedes eius et dixit: " In me sit, domine mi, haec iniquitas; loquatur, obsecro, ancilla tua in auribus tuis, et audi verba famulae tuae.
1SAM|25|25|Ne ponat, oro, dominus meus cor suum super virum istum iniquum Nabal, quia secundum nomen suum stultus est, et est stultitia cum eo; ego autem ancilla tua non vidi pueros domini mei, quos misisti.
1SAM|25|26|Nunc ergo, domine mi, vivit Dominus, et vivit anima tua, quia Dominus prohibuit te, ne venires in sanguine et salvares te manu tua; et nunc fiant sicut Nabal inimici tui et qui quaerunt domino meo malum.
1SAM|25|27|Quapropter suscipe benedictionem hanc, quam attulit ancilla tua domino meo, et da pueris, qui sequuntur dominum meum.
1SAM|25|28|Aufer iniquitatem famulae tuae. Faciens enim faciet Dominus domino meo domum fidelem, quia proelia Domini dominus meus proeliatur; malitia ergo non inveniatur in te omnibus diebus vitae tuae.
1SAM|25|29|Si enim surrexerit aliquando homo persequens te et quaerens animam tuam, erit anima domini mei custodita in fasciculo vitae apud Dominum Deum tuum; sed inimicorum tuorum animam ipse iaciat in impetu et circulo fundae.
1SAM|25|30|Cum ergo fecerit Dominus domino meo omnia, quae locutus est, bona de te et constituerit te ducem super Israel,
1SAM|25|31|non erit tibi hoc in singultum et in scrupulum cordis domino meo, quod effuderis sanguinem innoxium et ipse te ultus fueris; et cum benefecerit Dominus domino meo, recordaberis ancillae tuae ".
1SAM|25|32|Et ait David ad Abigail: " Benedictus Dominus, Deus Israel, qui misit te hodie in occursum meum. Et benedicta prudentia tua,
1SAM|25|33|et benedicta tu, quae prohibuisti me hodie, ne irem ad sanguinem et ulciscerer me manu mea.
1SAM|25|34|Alioquin, vivit Dominus, Deus Israel, qui prohibuit me malum facere tibi, nisi cito venisses in occursum mihi, non remansisset Nabal usque ad lucem matutinam quidquid masculini sexus ".
1SAM|25|35|Suscepit ergo David de manu eius omnia, quae attulerat ei, dixitque ei: Vade pacifice in domum tuam. Ecce audivi vocem tuam et honoravi faciem tuam ".
1SAM|25|36|Venit autem Abigail ad Nabal; et ecce erat ei convivium in domo eius quasi convivium regis, et cor Nabal iucundum; erat enim ebrius nimis. Et non indicavit ei verbum pusillum aut grande usque in mane.
1SAM|25|37|Diluculo autem, cum digessisset vinum Nabal, haec indicavit ei uxor sua; et emortuum est cor eius intrinsecus, et factus est quasi lapis.
1SAM|25|38|Cumque pertransissent decem dies, percussit Dominus Nabal, et mortuus est.
1SAM|25|39|Quod cum audisset David mortuum Nabal, ait: " Benedictus Dominus, qui iudicavit causam opprobrii mei de manu Nabal et servum suum custodivit a malo et malitiam Nabal reddidit Dominus in caput eius ".Misit ergo David et locutus est ad Abigail, ut sumeret eam sibi in uxorem.
1SAM|25|40|Et venerunt pueri David ad Abigail in Carmel et locuti sunt ad eam dicentes: " David misit nos ad te, ut accipiat te sibi in uxorem ".
1SAM|25|41|Quae consurgens adoravit prona in terram et ait: " Ecce famula tua sit in ancillam, ut lavet pedes servorum domini mei ".
1SAM|25|42|Et festinavit et surrexit Abigail et ascendit super asinum, et quinque puellae ierunt cum ea pedisequae eius; et secuta est nuntios David et facta est illi uxor.
1SAM|25|43|Sed et Achinoam accepit David de Iezrahel, et fuit utraque uxor eius.
1SAM|25|44|Saul autem dedit Michol filiam suam uxorem David Phalti filio Lais, qui erat de Gallim.
1SAM|26|1|Et venerunt Ziphaei ad Saul in Gabaa dicentes: " Ecce David absconditus est in colle Hachila, quae est ex adverso solitudinis ".
1SAM|26|2|Et surrexit Saul et descendit in desertum Ziph, et cum eo tria milia virorum de electis Israel, ut quaereret David in deserto Ziph.
1SAM|26|3|Et castrametatus est Saul in colle Hachila, quae erat ex adverso solitudinis in via. David autem habitabat in deserto; videns autem quod venisset Saul post se in desertum,
1SAM|26|4|misit exploratores et didicit quod illuc venisset certissime.
1SAM|26|5|Et surrexit David et venit ad locum, ubi erat Saul. Cumque vidisset locum, in quo dormiebat Saul et Abner filius Ner princeps militiae eius, Saulem dormientem in carragine et reliquum vulgus per circuitum eius,
1SAM|26|6|ait David ad Achimelech Hetthaeum et Abisai filium Sarviae fratrem Ioab dicens: " Quis descendet mecum ad Saul in castra? ". Dixitque Abisai: " Ego descendam tecum ".
1SAM|26|7|Venerunt ergo David et Abisai ad populum nocte et invenerunt Saul iacentem et dormientem in carragine et hastam fixam in terra ad caput eius, Abner autem et populum dormientes in circuitu eius.
1SAM|26|8|Dixitque Abisai ad David: " Conclusit Deus hodie inimicum tuum in manus tuas; nunc ergo perfodiam eum lancea in terra semel, et secundo opus non erit ".
1SAM|26|9|Et dixit David ad Abisai: " Ne interficias eum; quis enim extendit manum suam in christum Domini et innocens erit? ".
1SAM|26|10|Et dixit David: " Vivit Dominus quia Dominus percutiet eum, aut dies eius veniet, ut moriatur, aut in proelium descendens peribit.
1SAM|26|11|Propitius mihi sit Dominus, ne extendam manum meam in christum Domini. Nunc igitur tolle hastam, quae est ad caput eius, et scyphum aquae, et abeamus ".
1SAM|26|12|Tulit ergo David hastam et scyphum aquae, qui erat ad caput Saul, et abierunt; et non erat quisquam, qui videret et intellegeret et vigilaret, sed omnes dormiebant, quia sopor Domini irruerat super eos.
1SAM|26|13|Cumque transisset David ex adverso et stetisset in vertice montis de longe, et esset grande intervallum inter eos,
1SAM|26|14|clamavit David ad populum et ad Abner filium Ner dicens: " Nonne respondebis, Abner? ". Et respondens Abner ait: " Quis es tu? Clamasti ad regem! ".
1SAM|26|15|Et ait David ad Abner: " Numquid non vir tu es? Et quis alius similis tui in Israel? Quare ergo non custodisti dominum tuum regem? Ingressus est enim unus de turba, ut interficeret regem dominum tuum.
1SAM|26|16|Non est bonum hoc, quod fecisti. Vivit Dominus quoniam filii mortis estis vos, qui non custodistis dominum vestrum, christum Domini. Nunc ergo vide, ubi sit hasta regis et ubi scyphus aquae, qui erat ad caput eius ".
1SAM|26|17|Cognovit autem Saul vocem David et dixit: " Num vox tua haec est, fili mi David? ". Et ait David: " Vox mea, domine mi rex ".
1SAM|26|18|Et ait: " Quam ob causam dominus meus persequitur servum suum? Quid feci? Aut quod est in manu mea malum?
1SAM|26|19|Nunc ergo audiat, oro, dominus meus rex verba servi sui: Si Dominus incitat te adversum me, odoretur sacrificium; si autem filii hominum, maledicti sint in conspectu Domini, quia eiecerunt me hodie, ut non habitem in hereditate Domini dicentes: "Vade, servi diis alienis".
1SAM|26|20|Et nunc non effundatur sanguis meus in terra longe a facie Domini; quia egressus est rex Israel, ut quaerat pulicem unum, sicut persequitur quis perdicem in montibus ".
1SAM|26|21|Et ait Saul: " Peccavi. Revertere, fili mi David; nequaquam enim ultra malefaciam tibi, eo quod pretiosa fuerit anima mea in oculis tuis hodie; apparet quod stulte egerim et erraverim multum nimis ".
1SAM|26|22|Et respondens David ait: " Ecce hasta regis; transeat unus de pueris et tollat eam.
1SAM|26|23|Dominus autem retribuet unicuique secundum iustitiam suam et fidem; tradidit enim te Dominus hodie in manu mea, et nolui extendere manum meam in christum Domini.
1SAM|26|24|Et sicut magnificata est anima tua hodie in oculis meis, sic magnificetur anima mea in oculis Domini, et liberet me de omni angustia ".
1SAM|26|25|Ait ergo Saul ad David: " Benedictus tu, fili mi David; et quidem faciens facies et potens poteris ". Abiit autem David in viam suam, et Saul reversus est in locum suum.
1SAM|27|1|Et ait David in corde suo: " Aliquando incidam in uno die in manu Saul; nonne melius est ut fugiam et salver in terra Philisthinorum, ut desperet Saul cessetque me quaerere in cunctis finibus Israel? Fugiam ergo manus eius ".
1SAM|27|2|Et surrexit David et abiit ipse et sescenti viri cum eo ad Achis filium Maoch regem Geth.
1SAM|27|3|Et habitavit David cum Achis in Geth ipse et viri eius unusquisque cum domo sua; David et duae uxores eius, Achinoam Iezrahelites et Abigail uxor Nabal de Carmel.
1SAM|27|4|Et nuntiatum est Saul quod fugisset David in Geth, et non addidit ultra ut quaereret eum.
1SAM|27|5|Dixit autem David ad Achis: " Si inveni gratiam in oculis tuis, detur mihi locus in una urbium regionis huius, ut habitem ibi. Cur enim manet servus tuus in civitate regis tecum? ".
1SAM|27|6|Dedit itaque ei Achis in die illa Siceleg; propter quam causam facta est Siceleg regum Iudae usque in diem hanc.
1SAM|27|7|Fuit autem numerus dierum, quibus habitavit David in regione Philisthinorum, annus et quattuor menses.
1SAM|27|8|Et ascendit David et viri eius et agebant praedas de Gesuri et de Gerzi et de Amalecitis; hae enim gentes habitabant terram, quae est a Telem in via Sur et usque ad terram Aegypti.
1SAM|27|9|Et percutiebat David omnem terram nec relinquebat viventem virum et mulierem; tollensque oves et boves et asinos et camelos et vestes revertebatur et veniebat ad Achis.
1SAM|27|10|Dicebat autem ei Achis: " In quem irruistis hodie? ". Respondebatque David: " Contra Nageb Iudae vel contra Nageb Ierameel vel contra Nageb Ceni ".
1SAM|27|11|Viro et mulieri non parcebat David nec adducebat in Geth dicens: " Ne forte loquantur adversum nos: "Haec fecit David" ". Et hoc erat decretum illi omnibus diebus, quibus habitavit in regione Philisthinorum.
1SAM|27|12|Credidit ergo Achis David dicens: " Valde odiosum se fecit populo suo Israel; eritigitur mihi servus sempiternus ".
1SAM|28|1|Factum est autem in diebus illis, congregaverunt Phili sthim agmina sua, ut praepararentur ad bellum contra Israel. Dixitque Achis ad David: " Sciens nunc scito quoniam mecum egredieris in castris tu et viri tui ".
1SAM|28|2|Dixitque David ad Achis: " Ideo tu quoque scies, quae facturus est servus tuus ". Et ait Achis ad David: " Ideo custodem capitis mei ponam te cunctis diebus ".
1SAM|28|3|Samuel autem mortuus erat; planxeratque eum omnis Israel, et sepelierant eum in Rama urbe sua. Et Saul abstulerat magos et hariolos de terra.
1SAM|28|4|Congregatique sunt Philisthim et venerunt et castrametati sunt in Sunam. Congregavit autem et Saul universum Israel, et castrametati sunt in Gelboe.
1SAM|28|5|Et vidit Saul castra Philisthim et timuit, et expavit cor eius nimis.
1SAM|28|6|Consuluitque Dominum, et non respondit ei neque per somnia neque per Urim neque per prophetas.
1SAM|28|7|Dixitque Saul servis suis: " Quaerite mihi mulierem habentem pythonem, et vadam ad eam et sciscitabor per illam ". Et dixerunt servi eius ad eum: Est mulier habens pythonem in Endor ".
1SAM|28|8|Mutavit ergo habitum suum vestitusque est aliis vestimentis et abiit ipse et duo viri cum eo; veneruntque ad mulierem nocte, et ait: " Divina mihi in pythone et suscita mihi, quem dixero tibi ".
1SAM|28|9|Et ait mulier ad eum: " Ecce tu nosti, quanta fecerit Saul et quomodo eraserit magos et hariolos de terra; quare ergo insidiaris animae meae, ut occidar? ".
1SAM|28|10|Et iuravit ei Saul in Domino dicens: " Vivit Dominus quia non veniet tibi quidquam mali propter hanc rem ".
1SAM|28|11|Dixitque ei mulier: " Quem suscitabo tibi? ". Qui ait: " Samuelem suscita mihi ".
1SAM|28|12|Cum autem vidisset mulier Samuelem, exclamavit voce magna et dixit ad Saul: " Quare imposuisti mihi? Tu es enim Saul! ".
1SAM|28|13|Dixitque ei rex: " Noli timere. Quid vidisti? ". Et ait mulier ad Saul: Hominem divinum vidi ascendentem de terra ".
1SAM|28|14|Dixitque ei: " Qualis est forma eius? ". Quae ait: " Vir senex ascendit et ipse amictus est pallio ". Intellexit Saul quod Samuel esset et inclinavit se super faciem suam in terra et adoravit.
1SAM|28|15|Dixit autem Samuel ad Saul: " Quare inquietasti me, ut suscitarer? ". Et ait Saul: " Coartor nimis. Siquidem Philisthim pugnant adversum me, et Deus recessit a me et exaudire me noluit neque in manu prophetarum neque per somnia; vocavi ergo te, ut ostenderes mihi quid faciam ".
1SAM|28|16|Et ait Samuel: " Quid interrogas me, cum Dominus recesserit a te et factus est adversarius tuus?
1SAM|28|17|Fecit enim Dominus, sicut locutus est in manu mea, et scidit regnum de manu tua et dedit illud proximo tuo David,
1SAM|28|18|quia non oboedisti voci Domini neque fecisti iram furoris eius in Amalec. Idcirco quod pateris, fecit tibi Dominus hodie.
1SAM|28|19|Et dabit Dominus etiam Israel tecum in manu Philisthim; cras autem tu et filii tui mecum eritis, sed et castra Israel tradet Dominus in manu Philisthim ".
1SAM|28|20|Statimque Saul cecidit porrectus in terram; extimuerat enim verba Samuel, et robur non erat in eo, quia non comederat panem tota die illa et tota nocte illa.
1SAM|28|21|Accessit itaque mulier ad Saul et vidit quod conturbatus esset valde; dixitque ad eum: " Ecce audivit ancilla tua vocem tuam, et posui animam meam in manu mea et oboedivi sermonibus tuis, quos locutus es ad me.
1SAM|28|22|Nunc igitur audi et tu vocem ancillae tuae, ut ponam coram te buccellam panis, et comedens convalescas, ut possis iter facere ".
1SAM|28|23|Qui renuit et ait: " Non comedam ". Coegerunt autem eum servi sui et mulier; et tandem, audita voce eorum, surrexit de terra et sedit super lectum.
1SAM|28|24|Mulier autem illa habebat vitulum pascualem in domo; et festinavit et occidit eum, tollensque farinam miscuit eam et coxit azyma.
1SAM|28|25|Et posuit ante Saul et ante servos eius. Qui cum comedissent, surrexerunt et abierunt hac eadem nocte.
1SAM|29|1|Congregata sunt ergo Philisthim universa agmina in Aphec; sed et Israel castrametatus est super fontem, qui erat in Iezrahel.
1SAM|29|2|Et principes quidem Philisthim incedebant in centuriis et milibus; David autem et viri eius incedebant in novissimo agmine cum Achis.
1SAM|29|3|Dixeruntque principes Philisthim: " Quid sibi volunt Hebraei isti? ". Et ait Achis ad principes Philisthim: " Nonne iste est David, qui fuit servus Saul regis Israel et est apud me multis diebus vel annis, et non inveni in eo quidquam ex die, qua transfugit ad me, usque ad diem hanc? ".
1SAM|29|4|Irati sunt autem adversus eum principes Philisthim et dixerunt ei: " Revertatur vir iste et sedeat in loco suo, in quo constituisti eum, et non descendat nobiscum in proelium, ne fiat nobis adversarius, cum proeliari coeperimus. Quomodo enim aliter placare poterit dominum suum nisi in capitibus horum virorum?
1SAM|29|5|Nonne iste est David, cui cantabant in choris dicentes: "Percussit Saul milia sua, et David decem milia sua"? ".
1SAM|29|6|Vocavit ergo Achis David et ait ei: " Vivit Dominus quia rectus es tu, et bonus est in conspectu meo exitus tuus et introitus tuus mecum in castris, et non inveni in te quidquam mali ex die, qua venisti ad me, usque ad diem hanc. Sed principibus non places.
1SAM|29|7|Revertere ergo et vade in pace et non offendes oculos principum Philisthim ".
1SAM|29|8|Dixitque David ad Achis: " Quid enim feci, et quid invenisti in me servo tuo a die, qua fui in conspectu tuo, usque in diem hanc, ut non veniam et pugnem contra inimicos domini mei regis? ".
1SAM|29|9|Respondens autem Achis locutus est ad David: " Scio quia bonus es tu in oculis meis sicut angelus Dei; sed principes Philisthim dixerunt: "Non ascendet nobiscum in proelium".
1SAM|29|10|Igitur consurge mane, tu et servi domini tui, qui venerunt tecum, et, cum de nocte surrexeritis et coeperit dilucescere, pergite ".
1SAM|29|11|Surrexit itaque de nocte David ipse et viri eius, ut proficiscerentur mane et reverterentur ad terram Philisthim. Philisthim autem ascenderunt in Iezrahel.
1SAM|30|1|Cumque venissent David et viri eius in Siceleg die tertia, Amalecitae impetum fecerant contra Nageb et contra Siceleg et percusserant Siceleg et succenderant eam igni;
1SAM|30|2|et captivas duxerant mulieres et omnes in ea a minimo usque ad magnum et non interfecerant quemquam, sed secum duxerant et pergebant in itinere suo.
1SAM|30|3|Cum ergo venisset David et viri eius ad civitatem et invenissent eam succensam igni et uxores suas et filios suos et filias ductas esse captivas,
1SAM|30|4|levaverunt David et populus, qui erat cum eo, voces suas et planxerunt, donec deficerent in eis lacrimae.
1SAM|30|5|Siquidem et duae uxores David captivae ductae fuerant, Achinoam Iezrahelites et Abigail uxor Nabal de Carmel.
1SAM|30|6|Et angustiatus est David valde; volebat enim eum populus lapidare, quia amara erat anima uniuscuiusque viri super filiis suis et filiabus. Confortatus est autem David in Domino Deo suo
1SAM|30|7|et ait ad Abiathar sacerdotem filium Achimelech: " Applica ad me ephod. Et applicuit Abiathar ephod ad David.
1SAM|30|8|Et consuluit David Dominum dicens: " Persequar latrunculos hos et comprehendam eos an non? ". Dixitque ei: " Persequere; absque dubio enim comprehendes eos et excuties praedam ".
1SAM|30|9|Abiit ergo David ipse et sescenti viri, qui erant cum eo, et venerunt usque ad torrentem Besor, et lassi quidam substiterunt.
1SAM|30|10|Persecutus est autem David ipse et quadringenti viri; et reliqui substiterunt: ducenti, qui lassi transire non poterant torrentem Besor.
1SAM|30|11|Et invenerunt virum Aegyptium in agro et adduxerunt eum ad David; dederuntque ei panem, et comedit, et dederunt ei aquam bibere,
1SAM|30|12|sed et dederunt ei fragmen massae caricarum et duas ligaturas uvae passae. Quae cum comedisset, reversus est spiritus eius; non enim comederat panem neque biberat aquam tribus diebus et tribus noctibus.
1SAM|30|13|Dixit itaque ei David: " Cuius es tu vel unde? ". Qui ait ei: " Puer Aegyptius ego sum servus viri Amalecitae; dereliquit autem me dominus meus, quia aegrotare coepi nudiustertius.
1SAM|30|14|Siquidem nos erupimus contra Nageb Cherethi et contra Nageb Iudae et Nageb Chaleb et Siceleg succendimus igni ".
1SAM|30|15|Dixitque ei David: " Potes me ducere ad istum cuneum? ". Qui ait: " Iura mihi per Deum quod non occidas me et non tradas me in manu domini mei, et ducam te ad cuneum istum ". Et iuravit ei David.
1SAM|30|16|Qui cum duxisset eum, ecce illi discumbebant super faciem universae terrae comedentes et bibentes et festum celebrantes pro cuncta praeda et spoliis, quae ceperant de terra Philisthim et de terra Iudae.
1SAM|30|17|Et percussit eos David die altera a diluculo usque ad vesperam, et non evasit ex eis quisquam, nisi quadringenti viri adulescentes, qui ascenderant camelos et fugerant.
1SAM|30|18|Eruit ergo David omnia, quae ceperant Amalecitae, et duas uxores suas eruit.
1SAM|30|19|Nec defuit quidquam a parvo usque ad magnum tam de filiis quam de filiabus et de spoliis, et, quaecumque rapuerant, omnia reduxit David.
1SAM|30|20|Cepit ergo David universos greges et armenta, et minaverunt ante faciem eius possessionem hanc dixeruntque: " Haec est praeda David ".
1SAM|30|21|Venit autem David ad ducentos viros, qui lassi substiterant nec sequi potuerant David, et residere eos iusserat in torrente Besor. Qui egressi sunt obviam David et populo, qui erat cum eo. Accedens autem David ad populum salutavit eos pacifice.
1SAM|30|22|Respondensque omnis vir pessimus et iniquus de viris, qui ierant cum David, dixit: " Quia non venerunt nobiscum, non dabimus eis quidquam de praeda, quam eruimus; sed sufficiat unicuique uxor sua et filii; quos cum acceperint, recedant ".
1SAM|30|23|Dixit autem David: " Non sic facietis, fratres mei, de his, quae tradidit Dominus nobis, et custodivit nos et dedit latrunculos, qui eruperant adversum nos, in manu nostra;
1SAM|30|24|nec audiet vos quisquam super sermone hoc; aequa enim pars erit descendentis ad proelium et remanentis ad sarcinas, et similiter divident.
1SAM|30|25|Et factum est hoc ex die illa et deinceps constitutum ut praeceptum et quasi lex in Israel usque ad diem hanc.
1SAM|30|26|Venit ergo David in Siceleg et misit dona de praeda senioribus Iudae proximis suis dicens: " Accipite benedictionem de praeda hostium Domini ";
1SAM|30|27|his, qui erant in Bethul et qui in Ramathnageb et qui in Iether
1SAM|30|28|et qui in Aroer et qui in Sephamoth et qui in Esthemo
1SAM|30|29|et qui in Carmel et qui in urbibus Ierameeli et qui in urbibus Ceni
1SAM|30|30|et qui in Horma et qui in Borasan et qui in Athach
1SAM|30|31|et qui in Hebron et reliquis locis, in quibus commoratus fuerat David ipse et viri eius.
1SAM|31|1|Philisthim autem pugnabant adversum Israel; et fugerunt viri Israel ante faciem Philisthim et ceciderunt interfecti in monte Gelboe.
1SAM|31|2|Irrueruntque Philisthim in Saul et filios eius et percusserunt Ionathan et Abinadab et Melchisua filios Saul.
1SAM|31|3|Totumque pondus proelii versum est in Saul; et consecuti sunt eum viri arcu, et vulneratus est vehementer a sagittariis.
1SAM|31|4|Dixitque Saul ad armigerum suum: " Evagina gladium tuum et percute me, ne forte veniant incircumcisi isti et confodiant me et illudant mihi ". Et noluit armiger eius; erat enim nimio timore perterritus. Arripuit itaque Saul gladium et irruit super eum.
1SAM|31|5|Quod cum vidisset armiger eius, videlicet quod mortuus esset Saul, irruit etiam ipse super gladium suum et mortuus est cum eo.
1SAM|31|6|Mortuus est ergo Saul et tres filii eius et armiger illius et universi viri eius in die illa pariter.
1SAM|31|7|Videntes autem viri Israel, qui erant trans vallem et trans Iordanem, quod fugissent viri Israelitae et quod mortuus esset Saul et filii eius, reliquerunt civitates suas et fugerunt. Veneruntque Philisthim et habitaverunt ibi.
1SAM|31|8|Facta autem die altera, venerunt Philisthim, ut spoliarent interfectos, et invenerunt Saul et tres filios eius iacentes in monte Gelboe.
1SAM|31|9|Et praeciderunt caput Saul et exspoliaverunt eum armis, quae miserunt in terram Philisthinorum per circuitum, ut annuntiaretur in templis idolorum suorum et populo.
1SAM|31|10|Et posuerunt arma eius in templo Astharoth, corpus vero eius suspenderunt in muro Bethsan.
1SAM|31|11|Quod cum audissent habitatores Iabes Galaad, quaecumque fecerant Philisthim Saul,
1SAM|31|12|surrexerunt omnes viri fortissimi et ambulaverunt tota nocte et tulerunt cadaver Saul et cadavera filiorum eius de muro Bethsan; veneruntque Iabes et combusserunt ea ibi.
1SAM|31|13|Et tulerunt ossa eorum et sepelierunt sub myrice in Iabes et ieiunaverunt septem diebus.
2SAM|1|1|Factum est autem, postquam mortuus est Saul, ut David re verteretur a caede Amalec et maneret in Siceleg dies duos.
2SAM|1|2|In die autem tertia apparuit homo veniens de castris Saul veste conscissa et pulvere aspersus caput; et, ut venit ad David, cecidit super faciem suam et adoravit.
2SAM|1|3|Dixitque ad eum David: " Unde venis? ". Qui ait ad eum: " De castris Israel fugi ".
2SAM|1|4|Et dixit ad eum David: " Quid enim factum est? Indica mihi ". Qui ait: " Fugit populus ex proelio, et multi corruentes e populo mortui sunt; sed et Saul et Ionathan filius eius interierunt ".
2SAM|1|5|Dixitque David ad adulescentem, qui nuntiabat ei: " Unde scis quia mortuus est Saul et Ionathan filius eius? ".
2SAM|1|6|Et ait adulescens, qui narrabat ei: " Casu veni in montem Gelboe, et Saul incumbebat super hastam suam. Porro currus et equites appropinquabant ei,
2SAM|1|7|et conversus post tergum suum vidensque me vocavit. Cui cum respondissem: Adsum,
2SAM|1|8|dixit mihi: "Quisnam es tu?". Et dixi ad eum: Amalecites ego sum.
2SAM|1|9|Et locutus est mihi: "Sta super me et interfice me, quoniam tenent me angustiae, et adhuc tota anima mea in me est".
2SAM|1|10|Stansque super eum occidi illum; sciebam enim quod vivere non poterat post ruinam. Et tuli diadema, quod erat in capite eius, et armillam de brachio illius et attuli ad te dominum meum huc ".
2SAM|1|11|Apprehendens autem David vestimenta sua scidit omnesque viri, qui erant cum eo;
2SAM|1|12|et planxerunt et fleverunt et ieiunaverunt usque ad vesperam super Saul et super Ionathan filium eius et super populum Domini et super domum Israel, quod corruissent gladio.
2SAM|1|13|Dixitque David ad iuvenem, qui nuntiaverat ei: " Unde es? ". Qui respondit: " Filius hominis advenae Amalecitae ego sum ".
2SAM|1|14|Et ait ad eum David: " Quare non timuisti mittere manum tuam, ut occideres christum Domini? ".
2SAM|1|15|Vocansque David unum de pueris ait: " Accedens irrue in eum ". Qui percussit illum, et mortuus est.
2SAM|1|16|Et ait ad eum David: " Sanguis tuus super caput tuum; os enim tuum locutum est adversum te dicens: "Ego interfeci christum Domini" ".
2SAM|1|17|Planxit autem David planctum huiuscemodi super Saul et super Ionathan filium eius;
2SAM|1|18|et praecepit, ut docerent filios Iudae canticum Arcus, sicut scriptum est in libro Iusti, et ait:
2SAM|1|19|" Incliti, o Israel, super montes tuos interfecti,quomodo ceciderunt fortes!
2SAM|1|20|Nolite annuntiare in Gethneque annuntietis in compitis Ascalonis,ne forte laetentur filiae Philisthim,ne exsultent filiae incircumcisorum.
2SAM|1|21|Montes Gelboe, nec ros nec pluviae veniant super vos,neque sint agri oblationum!Quia ibi abiectus est clipeus fortium,clipeus Saul, quasi non esset unctus oleo.
2SAM|1|22|A sanguine interfectorum, ab adipe fortiumarcus Ionathan numquam rediit retrorsum,et gladius Saul non est reversus inanis.
2SAM|1|23|Saul et Ionathan amabiles et decori in vita sua,in morte quoque non sunt divisi,aquilis velociores, leonibus fortiores.
2SAM|1|24|Filiae Israel, super Saul flete,qui vestiebat vos coccino in deliciis, qui praebebat ornamenta aurea cultui vestro.
2SAM|1|25|Quomodo ceciderunt fortes in proelio!Ionathan in excelsis tuis occisus est.
2SAM|1|26|Doleo super te, frater mi Ionathan,suavis nimis mihi;mirabilis amor tuus mihisuper amorem mulierum.
2SAM|1|27|Quomodo ceciderunt fortes,et perierunt arma bellica! ".
2SAM|2|1|Igitur post haec consuluit David Dominum dicens: " Num ascendam in unam de civitatibus Iudae? ". Et ait Dominus ad eum: " Ascende ". Dixitque David: " Quo ascendam? ". Et respondit ei: " In Hebron ".
2SAM|2|2|Ascendit ergo David et duae uxores eius, Achinoam Iezrahelites et Abigail uxor Nabal de Carmel;
2SAM|2|3|sed et viros, qui erant cum eo, duxit David singulos cum domo sua, et manserunt in oppidis Hebron.
2SAM|2|4|Veneruntque viri Iudae et unxerunt ibi David, ut regnaret super domum Iudae.Et nuntiatum est David quod viri Iabes Galaad sepelissent Saul.
2SAM|2|5|Misit ergo David nuntios ad viros Iabes Galaad dixitque ad eos: " Benedicti vos Domino, qui fecistis misericordiam hanc cum domino vestro Saul et sepelistis eum.
2SAM|2|6|Et nunc faciat quidem vobis Dominus misericordiam et veritatem; sed et ego reddam vobis similiter bonum, eo quod feceritis istud.
2SAM|2|7|Nunc autem confortentur manus vestrae, et estote fortes; licet enim mortuus sit dominus vester Saul, tamen me unxit domus Iudae in regem sibi.
2SAM|2|8|Abner autem filius Ner princeps exercitus Saul tulit Isbaal filium Saul et duxit eum in Mahanaim
2SAM|2|9|regemque constituit super Galaad et super Aser et super Iezrahel et super Ephraim et super Beniamin et super Israel universum.
2SAM|2|10|Quadraginta annorum erat Isbaal filius Saul, cum regnare coepisset super Israel, et duobus annis regnavit; sola autem domus Iudae sequebatur David.
2SAM|2|11|Et fuit numerus dierum, quos commoratus est David imperans in Hebron super domum Iudae, septem annorum et sex mensium.
2SAM|2|12|Egressusque est Abner filius Ner et pueri Isbaal filii Saul de Mahanaim in Gabaon.
2SAM|2|13|Porro Ioab filius Sarviae et pueri David egressi sunt et occurrerunt eis iuxta piscinam Gabaon; et, cum in unum convenissent e regione, constiterunt hi ex una parte piscinae et illi ex altera.
2SAM|2|14|Dixitque Abner ad Ioab: " Surgant pueri et ludant coram nobis ". Et respondit Ioab: " Surgant ".
2SAM|2|15|Surrexerunt ergo et transierunt numero duodecim de Beniamin ex parte Isbaal filii Saul, et duodecim de pueris David.
2SAM|2|16|Apprehensoque unusquisque capite comparis sui, defixit gladium in latus contrarii, et ceciderunt simul; vocatumque est nomen loci illius ager Laterum in Gabaon.
2SAM|2|17|Et ortum est bellum durum valde in die illa, fugatusque est Abner et viri Israel a pueris David.
2SAM|2|18|Erant autem ibi tres filii Sarviae: Ioab et Abisai et Asael. Porro Asael cursor velocissimus fuit quasi unus ex capreis, quae morantur in campis.
2SAM|2|19|Persequebatur autem Asael Abner et non declinavit ad dextram sive ad sinistram omittens persequi Abner.
2SAM|2|20|Respexit itaque Abner post tergum suum et ait: " Tune es Asael? ". Qui respondit: " Ego sum ".
2SAM|2|21|Dixitque ei Abner: " Vade ad dextram sive ad sinistram et apprehende unum de adulescentibus et tolle tibi spolia eius ". Noluit autem Asael omittere quin urgeret eum.
2SAM|2|22|Rursumque locutus est Abner ad Asael: " Recede, noli me sequi, ne compellar confodere te in terram et levare non potero faciem meam ad Ioab fratrem tuum ".
2SAM|2|23|Qui audire contempsit et noluit declinare. Percussit ergo eum Abner, aversa hasta in inguine, et exiit hasta retrorsum, et mortuus est ibi. Omnesque qui transibant per locum, in quo ceciderat Asael et mortuus erat, subsistebant.
2SAM|2|24|Persequentibus autem Ioab et Abisai fugientem Abner, sol occubuit; et venerunt usque ad collem Amma, qui est ex adverso Gaiah in via deserti in Gabaon.
2SAM|2|25|Congregatique sunt filii Beniamin ad Abner et conglobati in unum cuneum steterunt in summitate tumuli unius.
2SAM|2|26|Et exclamavit Abner ad Ioab et ait: " Num usque ad internecionem tuus mucro desaeviet? An ignoras quod periculosa sit desperatio? Usquequo non dicis populo, ut omittat persequi fratres suos? ".
2SAM|2|27|Et ait Ioab: " Vivit Deus, nisi locutus fuisses, usque mane non recessisset populus persequens unusquisque fratrem suum ".
2SAM|2|28|Insonuit ergo Ioab bucina, et stetit omnis exercitus; nec persecuti sunt ultra Israel neque certaverunt amplius.
2SAM|2|29|Abner autem et viri eius abierunt per Arabam tota nocte illa et transierunt Iordanem et, lustrato toto saltu Bethron, venerunt Mahanaim.
2SAM|2|30|Porro Ioab reversus, omisso Abner, congregavit omnem populum; et defuerunt de pueris David decem et novem viri, excepto Asaele;
2SAM|2|31|servi autem David percusserunt de Beniamin et ex viris, qui erant cum Abner, trecentos sexaginta, qui et mortui sunt.
2SAM|2|32|Tuleruntque Asael et sepelierunt eum in sepulcro patris sui in Bethlehem. Et ambulaverunt tota nocte Ioab et viri, qui erant cum eo, et in ipso crepusculo pervenerunt in Hebron.
2SAM|3|1|Facta est ergo longa concertatio inter domum Saul et inter do mum David: David semper invalescens, domus autem Saul decrescens cotidie.
2SAM|3|2|Nati quoque sunt filii David in Hebron. Fuitque primogenitus eius Amnon de Achinoam Iezrahelitide,
2SAM|3|3|et post eum Cheleab de Abigail uxore Nabal de Carmel, porro tertius Absalom filius Maacha filiae Tholmai regis Gesur,
2SAM|3|4|quartus autem Adonias filius Haggith et quintus Saphatia filius Abital,
2SAM|3|5|sextus quoque Iethraam de Egla uxore David. Hi nati sunt David in Hebron.
2SAM|3|6|Cum ergo esset proelium inter domum Saul et domum David, Abner filius Ner regebat domum Saul.
2SAM|3|7|Fuerat autem Sauli concubina nomine Respha filia Aia. Dixitque Isbaal ad Abner:
2SAM|3|8|" Quare ingressus es ad concubinam patris mei? ". Qui iratus nimis propter verba Isbaal ait: " Numquid caput canis ego sum de Iuda? Hodie facio misericordiam super domum Saul patris tui et super fratres et proximos eius et non tradidi te in manu David. Et tu requisisti in me quod argueres pro muliere hodie.
2SAM|3|9|Haec faciat Deus Abner et haec addat ei, nisi, quomodo iuravit Dominus David, sic faciam cum eo,
2SAM|3|10|ut transferatur regnum de domo Saul, et confirmetur thronus David super Israel et super Iudam a Dan usque Bersabee ".
2SAM|3|11|Et non potuit respondere ei quidquam, quia metuebat illum.
2SAM|3|12|Misit ergo Abner nuntios ad David pro se dicentes: " Cuius est terra?, et ut loquerentur: " Fac mecum amicitias, et erit manus mea tecum, et reducam ad te universum Israel ".
2SAM|3|13|Qui ait: " Optime, ego faciam tecum amicitias, sed unam rem peto a te dicens: Non videbis faciem meam, nisi prius adduxeris Michol filiam Saul; et sic venies et videbis me ".
2SAM|3|14|Misit autem David nuntios ad Isbaal filium Saul dicens: "Redde uxorem meam Michol, quam despondi mihi centum praeputiis Philisthim ".
2SAM|3|15|Misit ergo Isbaal et tulit eam a viro suo Phaltiel filio Lais.
2SAM|3|16|Sequebaturque eam vir suus plorans usque Bahurim; et dixit ad eum Abner: " Vade, revertere ". Qui reversus est.
2SAM|3|17|Sermonem quoque intulit Abner ad seniores Israel dicens: " Tam heri quam nudiustertius quaerebatis David, ut regnaret super vos;
2SAM|3|18|nunc ergo facite, quoniam Dominus locutus est ad David dicens: "In manu servi mei David salvabo populum meum Israel de manu Philisthim et omnium inimicorum eius" ".
2SAM|3|19|Locutus est autem Abner etiam ad Beniamin; et abiit, ut loqueretur ad David in Hebron omnia, quae placuerant Israel et universo Beniamin.
2SAM|3|20|Venitque ad David in Hebron cum viginti viris, et fecit David Abner et viris eius, qui venerant cum eo, convivium.
2SAM|3|21|Et dixit Abner ad David: " Surgam, ut congregem ad te dominum meum regem omnem Israel, et ineant tecum foedus, et imperes omnibus, sicut desiderat anima tua ".Cum ergo deduxisset David Abner, et ille isset in pace,
2SAM|3|22|pueri David et Ioab venerunt ab expeditione cum praeda magna. Abner autem non erat cum David in Hebron, quia iam dimiserat eum, et profectus fuerat in pace,
2SAM|3|23|et Ioab et omnis exercitus, qui erat cum eo, postea venerant. Nuntiatum est itaque Ioab a narrantibus: " Venit Abner filius Ner ad regem, et dimisit eum, et abiit in pace ".
2SAM|3|24|Et ingressus est Ioab ad regem et ait: " Quid fecisti? Ecce venit Abner ad te; quare dimisisti eum, et abiit et recessit?
2SAM|3|25|Ignoras Abner filium Ner? Certe ad hoc venit, ut deciperet te et sciret exitum tuum et introitum tuum et nosset omnia quae agis ".
2SAM|3|26|Egressus itaque Ioab a David misit nuntios post Abner, et reduxerunt eum a cisterna Sira, ignorante David.
2SAM|3|27|Cumque redisset Abner in Hebron, seorsum abduxit eum Ioab ad medium portae, ut loqueretur ei quiete, et percussit illum ibi in inguine, et mortuus est in ultionem sanguinis Asael fratris eius.
2SAM|3|28|Quod cum audisset David rem iam gestam, ait: " Mundus ego sum et regnum meum apud Dominum usque in sempiternum a sanguine Abner filii Ner;
2SAM|3|29|et veniat super caput Ioab et super omnem domum patris eius, nec deficiat de domo Ioab fluxum morbidum sustinens, leprosus et tenens fusum et cadens gladio et indigens pane ".
2SAM|3|30|Igitur Ioab et Abisai frater eius interfecerunt Abner, eo quod occidisset Asael fratrem eorum in Gabaon in proelio.
2SAM|3|31|Dixit autem David ad Ioab et ad omnem populum, qui erat cum eo: " Scindite vestimenta vestra et accingimini saccis et plangite ante exequias Abner ". Porro rex David sequebatur feretrum.
2SAM|3|32|Cumque sepelissent Abner in Hebron, levavit rex David vocem suam et flevit super tumulum Abner; flevit autem et omnis populus.
2SAM|3|33|Plangensque rex et lugens Abner ait: Numquid, ut mori solent insensati,mori debuit Abner?
2SAM|3|34|Manus tuae ligatae non erant,et pedes tui non erant compedibus aggravati;sed, sicut solent cadere coram filiis iniquitatis, corruisti ".Congeminansque omnis populus flevit super eum.
2SAM|3|35|Cumque venisset universa multitudo reficere David pane clara adhuc die, iuravit David dicens: " Haec faciat mihi Deus et haec addat, si ante occasum solis gustavero panem vel aliud quidquam ".
2SAM|3|36|Omnisque populus audivit; et placuit eis, sicut cuncta, quae fecit rex, bona erant in conspectu totius populi.
2SAM|3|37|Et cognovit omne vulgus et universus Israel in die illa quoniam non actum fuisset a rege, ut occideretur Abner filius Ner.
2SAM|3|38|Dixit quoque rex ad servos suos: " Num ignoratis quoniam princeps et maximus cecidit hodie in Israel?
2SAM|3|39|Ego vero adhuc debilis sum, quamvis sim unctus rex; viri autem isti filii Sarviae duriores sunt quam ego. Retribuat Dominus facienti malum iuxta malitiam suam ".
2SAM|4|1|Audivit autem Isbaal filius Saul quod cecidisset Abner in He bron, et dissolutae sunt manus eius, omnisque Israel perturbatus est.
2SAM|4|2|Duo autem viri duces turmarum erant filio Saul, nomen uni Baana et nomen alteri Rechab filii Remmon Berothitae de filiis Beniamin; siquidem et Beroth reputata est in Beniamin.
2SAM|4|3|Fugerant enim Berothitae in Getthaim, factique sunt ibi advenae usque in tempus hoc.
2SAM|4|4|Erat autem Ionathan filio Saul filius debilis pedibus. Quinquennis enim fuit, quando venit nuntius de Saul et Ionathan ex Iezrahel. Tollens itaque eum nutrix sua fugit; cumque festinaret, ut fugeret, cecidit et claudus effectus est habuitque vocabulum Meribbaal.
2SAM|4|5|Venientes igitur filii Remmon Berothitae, Rechab et Baana, ingressi sunt, fervente die, domum Isbaal, qui dormiebat super stratum suum meridie; et ostiaria domus purgans triticum obdormivit.
2SAM|4|6|Ingressi sunt ergo usque interiora domus et percusserunt eum in inguine Rechab et Baana frater eius et fugerunt.
2SAM|4|7|Cum autem ingressi fuissent domum, ille dormiebat super lectum suum in conclavi, et percutientes interfecerunt eum; sublatoque capite eius, abierunt per viam Arabae tota nocte.
2SAM|4|8|Et attulerunt caput Isbaal ad David in Hebron dixeruntque ad regem: " Ecce caput Isbaal filii Saul inimici tui, qui quaerebat animam tuam; et dedit Dominus domino meo regi ultiones hodie de Saul et de semine eius ".
2SAM|4|9|Respondens autem David Rechab et Baana fratri eius filiis Remmon Berothitae dixit ad eos: " Vivit Dominus, qui eruit animam meam de omni angustia,
2SAM|4|10|quoniam eum, qui annuntiaverat mihi et dixerat: "Mortuus est Saul", qui putabat se prospera nuntiare, tenui et occidi in Siceleg, cui oportebat me dare mercedem pro nuntio;
2SAM|4|11|quanto magis nunc, cum homines impii interfecerunt virum innoxium in domo sua super lectum suum, non quaeram sanguinem eius de manu vestra et auferam vos de terra? ".
2SAM|4|12|Praecepit itaque David pueris, et interfecerunt eos; praecidentesque manus et pedes eorum suspenderunt eos super piscinam in Hebron. Caput autem Isbaal tulerunt et sepelierunt in sepulcro Abner in Hebron.
2SAM|5|1|Et venerunt universae tribus Is rael ad David in Hebron dicen tes: " Ecce nos os tuum et caro tua sumus.
2SAM|5|2|Sed et heri et nudiustertius, cum esset Saul rex super nos, tu eras educens et reducens Israel. Dixit autem Dominus ad te: "Tu pasces populum meum Israel et tu eris dux super Israel" ".
2SAM|5|3|Venerunt quoque omnes senes Israel ad regem in Hebron, et percussit cum eis rex David foedus in Hebron coram Domino; unxeruntque David in regem super Israel.
2SAM|5|4|Triginta annorum erat David, cum regnare coepisset, et quadraginta annis regnavit:
2SAM|5|5|in Hebron regnavit super Iudam septem annis et sex mensibus; in Ierusalem autem regnavit triginta tribus annis super omnem Israel et Iudam.
2SAM|5|6|Et abiit rex et omnes viri, qui erant cum eo, in Ierusalem ad Iebusaeum habitatorem terrae. Qui dixit ad David: "Non ingredieris huc, sed depellent te caeci et claudi ", significantes: " Non ingredietur David huc.
2SAM|5|7|Cepit autem David arcem Sion: haec est civitas David.
2SAM|5|8|Dixerat enim David in die illa: " Omnis, qui percutiet Iebusaeum, attingat per cuniculum fontis claudos et caecos exosos animae David ". Idcirco dicitur in proverbio: " Caecus et claudus non intrabunt in domum.
2SAM|5|9|Habitavit autem David in arce et vocavit eam Civitatem David; et aedificavit per gyrum a Mello et intrinsecus.
2SAM|5|10|Et ibat proficiens atque succrescens, et Dominus, Deus exercituum, erat cum eo.
2SAM|5|11|Misit quoque Hiram rex Tyri nuntios ad David et ligna cedrina et artifices lignorum artificesque lapidum pro parietibus; et aedificaverunt domum David.
2SAM|5|12|Et cognovit David quoniam confirmasset eum Dominus regem super Israel et quoniam exaltasset regnum eius super populum suum Israel.
2SAM|5|13|Accepitque David adhuc concubinas et uxores de Ierusalem, postquam venerat de Hebron; natique sunt David et alii filii et filiae.
2SAM|5|14|Et haec nomina eorum, qui nati sunt ei in Ierusalem: Samua et Sobab et Nathan et Salomon
2SAM|5|15|et Iebahar et Elisua et Napheg
2SAM|5|16|et Iaphia et Elisama et Eliada et Eliphalet.
2SAM|5|17|Audierunt vero Philisthim quod unxissent David regem super Israel et ascenderunt universi, ut quaererent David. Quod cum audisset David, descendit in praesidium;
2SAM|5|18|Philisthim autem venientes diffusi sunt in valle Raphaim.
2SAM|5|19|Et consuluit David Dominum dicens: " Si ascendam ad Philisthim? Et si dabis eos in manu mea? ". Et dixit Dominus ad David: "Ascende, quia tradens dabo Philisthim in manu tua ".
2SAM|5|20|Venit ergo David in Baalpharasim (id est Dominus diruptionum); et percussit eos ibi et dixit: "Divisit Dominus inimicos meos coram me, sicut dividuntur aquae ". Propterea vocatum est nomen loci illius Baalpharasim.
2SAM|5|21|Et reliquerunt ibi sculptilia sua, quae tulit David et viri eius.
2SAM|5|22|Et addiderunt adhuc Philisthim ut ascenderent et diffusi sunt in valle Raphaim.
2SAM|5|23|Consuluit autem David Dominum, qui respondit: " Non ascendas, sed gyra post tergum eorum et venies ad eos ex adverso arborum celthium
2SAM|5|24|et, cum audieris sonitum gradientis in cacumine arborum celthium, tunc inibis proelium, quia tunc egredietur Dominus ante faciem tuam, ut percutiat castra Philisthim ".
2SAM|5|25|Fecit itaque David, sicut praeceperat ei Dominus; et percussit Philisthim de Gabaon usque dum venias Gazer.
2SAM|6|1|Congregavit autem rursum Da vid omnes electos ex Israel tri ginta milia.
2SAM|6|2|Surrexitque David et abiit, et universus populus, qui erat cum eo, in Baala Iudae, ut adducerent inde arcam Dei, super quam invocatum est nomen Domini exercituum sedentis in cherubim super eam.
2SAM|6|3|Et imposuerunt arcam Dei super plaustrum novum tuleruntque eam de domo Abinadab, qui erat in colle. Oza autem et Ahio filii Abinadab minabant plaustrum:
2SAM|6|4|Oza ambulabat iuxta arcam, et Ahio praecedebat eam.
2SAM|6|5|David autem et omnis Israel ludebant coram Domino omni virtute in canticis et citharis et lyris et tympanis et sistris et cymbalis.
2SAM|6|6|Postquam autem venerunt ad aream Nachon, extendit manum Oza ad arcam Dei et tenuit eam, quoniam boves lascivientes proruperunt.
2SAM|6|7|Iratusque est indignatione Dominus contra Ozam et percussit eum super temeritate; qui mortuus est ibi iuxta arcam Dei.
2SAM|6|8|Contristatus autem est David, eo quod diruptionem dirupisset Dominus in Ozam; et vocatum est nomen loci illius Pharesoza (id est Diruptio Ozae) usque in diem hanc.
2SAM|6|9|Et extimuit David Dominum in die illa dicens: " Quomodo ingredietur ad me arca Domini? ".
2SAM|6|10|Et noluit divertere ad se arcam Domini in civitate David, sed divertit eam in domum Obededom Getthaei.
2SAM|6|11|Et habitavit arca Domini in domo Obededom Getthaei tribus mensibus, et benedixit Dominus Obededom et omnem domum eius.
2SAM|6|12|Nuntiatumque est regi David: " Benedixit Dominus Obededom et omnia eius propter arcam Dei ". Abiit ergo David et adduxit arcam Dei de domo Obededom in civitatem David cum gaudio.
2SAM|6|13|Cumque progressi essent, qui portabant arcam Domini, sex passus, immolavit bovem et vitulum saginatum,
2SAM|6|14|et David saltabat totis viribus ante Dominum. Porro David erat accinctus ephod lineo.
2SAM|6|15|Et David et omnis domus Israel ducebant arcam Domini in iubilo et in clangore bucinae.
2SAM|6|16|Cumque intrasset arca Domini in civitatem David, Michol filia Saul prospiciens per fenestram vidit regem David subsilientem atque saltantem coram Domino et despexit eum in corde suo.
2SAM|6|17|Et introduxerunt arcam Domini et posuerunt eam in loco suo in medio tabernaculi, quod tetenderat ei David; et obtulit David coram Domino holocausta et pacifica.
2SAM|6|18|Cumque complesset offerens holocaustum et pacifica, benedixit populo in nomine Domini exercituum.
2SAM|6|19|Et partitus est multitudini universae Israel tam viro quam mulieri singulis collyridam panis unam et laganum palmarum unum et palatham unam. Et abiit omnis populus unusquisque in domum suam.
2SAM|6|20|Reversusque est et David, ut benediceret domui suae, et egressa Michol filia Saul in occursum David ait: " Quam gloriosus fuit hodie rex Israel discooperiens se ante ancillas servorum suorum, quasi si nudetur unus de scurris! ".
2SAM|6|21|Dixitque David ad Michol: " Ante Dominum salto. Benedictus Dominus, qui elegit me potius quam patrem tuum et quam omnem domum eius, ut constitueret me ducem super populum Domini, super Israel!
2SAM|6|22|Ludam in conspectu Domini et vilior fiam plus quam factus sum et ero deiectus in oculis meis, sed apud ancillas, de quibus locuta es, gloriosior apparebo ".
2SAM|6|23|Igitur Michol filiae Saul non est natus filius usque ad diem mortis suae.
2SAM|7|1|Factum est autem cum sedisset rex in domo sua, et Dominus de disset ei requiem undique ab universis inimicis suis,
2SAM|7|2|dixit ad Nathan prophetam: " Videsne quod ego habitem in domo cedrina, et arca Dei posita sit in medio pellium? ".
2SAM|7|3|Dixitque Nathan ad regem: " Omne, quod est in corde tuo, vade, fac, quia Dominus tecum est ".
2SAM|7|4|Factum est autem in nocte illa, et ecce sermo Domini ad Nathan dicens:
2SAM|7|5|" Vade et loquere ad servum meum David: Haec dicit Dominus: Numquid tu aedificabis mihi domum ad habitandum?
2SAM|7|6|Numquam enim habitavi in domo ex die, qua eduxi filios Israel de terra Aegypti, usque in diem hanc, sed ambulabam in tabernaculo et in tentorio.
2SAM|7|7|Per cuncta loca, quae transivi cum omnibus filiis Israel, numquid loquens locutus sum ad unum de iudicibus Israel, cui praecepi, ut pasceret populum meum Israel, dicens: Quare non aedificastis mihi domum cedrinam?
2SAM|7|8|Et nunc haec dices servo meo David: Haec dicit Dominus exercituum: Ego tuli te de pascuis sequentem greges, ut esses dux super populum meum Israel,
2SAM|7|9|et fui tecum in omnibus, ubicumque ambulasti, et interfeci universos inimicos tuos a facie tua; fecique tibi nomen grande iuxta nomen magnorum, qui sunt in terra.
2SAM|7|10|Et ponam locum populo meo Israel et plantabo eum, et habitabit in eo et non turbabitur amplius; nec addent filii iniquitatis ut affligant eum sicut prius
2SAM|7|11|et ex die, qua constitui iudices super populum meum Israel, et requiem dabo tibi ab omnibus inimicis tuis. Praedicitque tibi Dominus quod domum faciat tibi Dominus.
2SAM|7|12|Cumque completi fuerint dies tui, et dormieris cum patribus tuis, suscitabo semen tuum post te, quod egredietur de visceribus tuis; et firmabo regnum eius.
2SAM|7|13|Ipse aedificabit domum nomini meo, et stabiliam thronum regni eius usque in sempiternum.
2SAM|7|14|Ego ero ei in patrem, et ipse erit mihi in filium; qui si inique aliquid gesserit, arguam eum in virga virorum et in plagis filiorum hominum.
2SAM|7|15|Misericordiam autem meam non auferam ab eo, sicut abstuli a Saul, quem amovi a facie tua;
2SAM|7|16|et stabilis erit domus tua et regnum tuum usque in aeternum ante faciem meam, et thronus tuus erit firmus iugiter ".
2SAM|7|17|Secundum omnia verba haec et iuxta universam visionem istam sic locutus est Nathan ad David.
2SAM|7|18|Ingressus est autem rex David et sedit coram Domino et dixit: " Quis ego sum, Domine Deus, et quae domus mea, quia adduxisti me hucusque?
2SAM|7|19|Sed et hoc parum visum est in conspectu tuo, Domine Deus, et locutus es etiam de domo servi tui in longinquum, et ista est lex hominis, Domine Deus!
2SAM|7|20|Quid ergo addere poterit adhuc David, ut loquatur ad te? Tu enim scis servum tuum, Domine Deus.
2SAM|7|21|Propter verbum tuum et secundum cor tuum fecisti omnia magnalia haec, ita ut nota faceres servo tuo.
2SAM|7|22|Idcirco magnus es, Domine Deus, quia non est similis tui; neque est Deus extra te, iuxta omnia, quae audivimus auribus nostris.
2SAM|7|23|Quae est autem ut populus tuus Israel una gens in terra, propter quam ivit Deus, ut redimeret eam sibi in populum et poneret sibi nomen faceretque eis magnalia et horribilia, ut eiceres a facie populi tui, quem redemisti tibi ex Aegypto, gentes et deos eorum?
2SAM|7|24|Et firmasti tibi populum tuum Israel in populum sempiternum; et tu, Domine, factus es eis in Deum.
2SAM|7|25|Nunc ergo, Domine Deus, verbum, quod locutus es super servum tuum et super domum eius, confirma in sempiternum et fac, sicut locutus es!
2SAM|7|26|Et magnificetur nomen tuum usque in sempiternum, atque dicatur: Dominus exercituum est Deus super Israel". Et domus servi tui David erit stabilita coram te,
2SAM|7|27|quia tu, Domine exercituum, Deus Israel, revelasti aurem servi tui dicens: "Domum aedificabo tibi". Propterea invenit servus tuus cor suum, ut oraret te oratione hac.
2SAM|7|28|Nunc ergo, Domine Deus, tu es Deus, et verba tua erunt vera; cum ergo locutus sis ad servum tuum bona haec,
2SAM|7|29|dignare igitur benedicere domui servi tui, ut sit in sempiternum coram te, quia tu, Domine Deus, locutus es, et benedictione tua benedicetur domus servi tui in sempiternum ".
2SAM|8|1|Factum est autem post haec, percussit David Philisthim et humiliavit eos; et tulit David Geth et urbes eius de manu Philisthim.
2SAM|8|2|Et percussit Moab et mensus est eos funiculo sternens eos in terra; mensus est autem duos funiculos ad occidendum et unum funiculum plenum ad vivificandum; factusque est Moab David serviens sub tributo.
2SAM|8|3|Et percussit David Adadezer filium Rohob regem Soba, quando profectus est, ut dominaretur super flumen Euphraten.
2SAM|8|4|Et captis David ex parte eius mille septingentis equitibus et viginti milibus peditum, subnervavit omnes iugales curruum; dereliquit autem ex eis centum currus.
2SAM|8|5|Venit quoque Syria Damasci, ut praesidium ferret Adadezer regi Soba, et percussit David de Syria viginti duo milia virorum;
2SAM|8|6|et posuit David praesidium in Syria Damasci; factaque est Syria David serviens sub tributo. Et auxiliatus est Dominus David in omnibus, ad quaecumque profectus est.
2SAM|8|7|Et tulit David arma aurea, quae habebant servi Adadezer, et detulit ea in Ierusalem;
2SAM|8|8|et de Tebah et de Berothai civitatibus Adadezer tulit rex David aes multum nimis.
2SAM|8|9|Audivit autem Thou rex Emath quod percussisset David omne robur Adadezer
2SAM|8|10|et misit Thou Adoram filium suum ad regem David, ut salutaret eum congratulans et gratias ageret eo quod pugnasset cum Adadezer et percussisset eum; hostis quippe erat Thou Adadezer. Attulit autem Adoram et vasa argentea et vasa aurea et vasa aerea,
2SAM|8|11|quae et ipsa sanctificavit rex David Domino cum argento et auro, quae sanctificaverat de universis gentibus, quas subegerat:
2SAM|8|12|de Syria et Moab et filiis Ammon et Philisthim et Amalec et de manibus Adadezer filii Rohob regis Soba.
2SAM|8|13|Fecit quoque sibi David nomen cum reverteretur, percussa Idumaea in valle Salis, caesis decem et octo milibus.
2SAM|8|14|Et posuit in Idumaea praesidia; et facta est universa Idumaea serviens David. Et auxiliatus est Dominus David in omnibus, ad quaecumque profectus est.
2SAM|8|15|Et regnavit David super omnem Israel; faciebat quoque David iudicium et iustitiam omni populo suo.
2SAM|8|16|Ioab autem filius Sarviae erat super exercitum; porro Iosaphat filius Ahilud erat a commentariis,
2SAM|8|17|et Sadoc filius Achitob et Abiathar filius Achimelech sacerdotes, et Saraias scriba.
2SAM|8|18|Banaias autem filius Ioiadae super Cherethi et Phelethi; filii autem David sacerdotes erant.
2SAM|9|1|Et dixit David: " Putasne est aliquis, qui remanserit adhuc de domo Saul, ut faciam cum eo misericordiam propter Ionathan? ".
2SAM|9|2|Erat autem de domo Saul servus nomine Siba; quem cum vocasset rex ad se, dixit ei: " Tune es Siba? ". Et ille respondit: " Ego sum, servus tuus ".
2SAM|9|3|Et ait rex: " Num superest aliquis de domo Saul, ut faciam cum eo misericordiam Dei? ". Dixitque Siba regi: " Superest filius Ionathan, debilis pedibus ".
2SAM|9|4|" Ubi, inquit, est? ". Et Siba ad regem: " Ecce, ait, in domo est Machir filii Ammiel in Lodabar ".
2SAM|9|5|Misit ergo rex David et tulit eum de domo Machir filii Ammiel de Lodabar.
2SAM|9|6|Cum autem venisset Meribbaal filius Ionathan filii Saul ad David, corruit in faciem suam et adoravit. Dixitque David: " Meribbaal ". Qui respondit: " Adsum servus tuus ".
2SAM|9|7|Et ait ei David: "Ne timeas, quia faciens faciam in te misericordiam propter Ionathan patrem tuum; et restituam tibi omnes agros Saul patris tui, et tu comedes panem in mensa mea semper ".
2SAM|9|8|Qui adorans eum dixit: " Quis ego sum servus tuus, quoniam respexisti super canem mortuum similem mei? ".
2SAM|9|9|Vocavit itaque rex Sibam puerum Saul et dixit ei: " Omnia, quaecumque fuerunt Saul et universae domui eius, do filio domini tui.
2SAM|9|10|Operare igitur ei terram, tu et filii tui et servi tui, et, quod inferes, sit cibus domui domini tui, quo alantur; Meribbaal autem filius domini tui comedet semper panem super mensam meam ". Erant autem Sibae quindecim filii et viginti servi.
2SAM|9|11|Dixitque Siba ad regem: " Sicut iussisti, domine mi rex, servo tuo, sic faciet servus tuus ". Meribbaal autem comedebat super mensam eius quasi unus de filiis regis.
2SAM|9|12|Habebat autem Meribbaal filium parvulum nomine Micha; omnes vero, qui habitabant in domo Sibae, serviebant Meribbaal.
2SAM|9|13|Porro Meribbaal habitabat in Ierusalem, quia de mensa regis iugiter vescebatur; et erat claudus utroque pede.
2SAM|10|1|Factum est autem post haec, ut moreretur rex filiorum Ammon, et regnaret Hanon filius eius pro eo.
2SAM|10|2|Dixitque David: " Faciam misericordiam cum Hanon filio Naas, sicut fecit pater eius mecum misericordiam ". Misit ergo David consolans eum per servos suos super patris interitu. Cum autem venissent servi David in terram filiorum Ammon,
2SAM|10|3|dixerunt principes filiorum Ammon ad Hanon dominum suum: " Putas quod propter honorem patris tui David miserit ad te consolatores; et non ideo, ut investigaret et exploraret civitatem et everteret eam, misit David servos suos ad te? ".
2SAM|10|4|Tulit itaque Hanon servos David rasitque dimidiam partem barbae eorum et praecidit vestes eorum medias usque ad nates et dimisit eos.
2SAM|10|5|Quod cum nuntiatum esset David, misit in occursum eorum - erant enim viri confusi turpiter valde - et mandavit eis David: " Manete Iericho, donec crescat barba vestra, et tunc revertimini ".
2SAM|10|6|Videntes autem filii Ammon quod exosos se fecissent David, miserunt et conduxerunt mercede a Syria Bethrohob et a Syria Soba viginti milia peditum et a rege Maacha mille viros et a viris Tob duodecim milia virorum.
2SAM|10|7|Quod cum audisset David, misit Ioab et omnem exercitum, viros fortissimos.
2SAM|10|8|Egressi sunt ergo filii Ammon et direxerunt aciem ante ipsum introitum portae; Syri autem Soba et Rohob et viri Tob et Maacha seorsum erant in campo.
2SAM|10|9|Videns igitur Ioab quod praeparatum esset adversum se proelium et ex adverso et post tergum, elegit ex omnibus electis Israel et instruxit aciem contra Syros;
2SAM|10|10|reliquam autem partem populi tradidit Abisai fratri suo, qui direxit aciem adversus filios Ammon.
2SAM|10|11|Et ait Ioab: " Si praevaluerint adversum me Syri, eris mihi in adiutorium; si autem filii Ammon praevaluerint adversum te, auxiliabor tibi.
2SAM|10|12|Esto vir fortis, et fortiter agamus pro populo nostro et civitatibus Dei nostri; Dominus autem faciet, quod bonum est in conspectu suo ".
2SAM|10|13|Iniit itaque Ioab et populus, qui erat cum eo, certamen contra Syros, qui fugerunt a facie eius.
2SAM|10|14|Filii autem Ammon videntes quod fugissent Syri, fugerunt et ipsi a facie Abisai et ingressi sunt civitatem. Reversusque est Ioab a filiis Ammon et venit Ierusalem.
2SAM|10|15|Videntes igitur Syri quoniam corruissent coram Israel, congregati sunt pariter.
2SAM|10|16|Misitque Adadezer et eduxit Syros, qui erant trans fluvium, et venerunt in Elam; Sobach autem magister militiae Adadezer erat princeps eorum.
2SAM|10|17|Quod cum nuntiatum esset David, contraxit omnem Israelem et transivit Iordanem venitque in Elam. Et direxerunt aciem Syri ex adverso David et pugnaverunt contra eum.
2SAM|10|18|Fugeruntque Syri a facie Israel; et occidit David de Syris septingentos currus et quadraginta milia peditum et Sobach principem militiae percussit, qui ibi mortuus est.
2SAM|10|19|Videntes autem universi reges, qui erant in praesidio Adadezer, se victos esse ab Israel, fecerunt pacem cum Israel et servierunt eis. Timueruntque Syri auxilium praebere ultra filiis Ammon.
2SAM|11|1|Factum est autem vertente anno, eo tempore quo solent reges ad bella procedere, misit David Ioab et servos suos cum eo et universum Israel, et vastaverunt filios Ammon et obsederunt Rabba; David autem remansit in Ierusalem.
2SAM|11|2|Et factum est vespere, ut surgeret David de strato suo et deambularet in solario domus regiae. Viditque de solario mulierem se lavantem; erat autem mulier pulchra valde.
2SAM|11|3|Misit ergo rex et requisivit quae esset mulier; nuntiatumque ei est quod ipsa esset Bethsabee filia Eliam uxor Uriae Hetthaei.
2SAM|11|4|Missis itaque David nuntiis, tulit eam; quae cum ingressa esset ad illum, dormivit cum ea, quae se sanctificaverat ab immunditia sua.
2SAM|11|5|Et reversa est domum suam; cum autem concepisset, mittens nuntiavit David et ait: " Concepi ".
2SAM|11|6|Misit autem David ad Ioab dicens: " Mitte ad me Uriam Hetthaeum ". Misitque Ioab Uriam ad David,
2SAM|11|7|et venit Urias ad David. Quaesivitque David quam recte ageret Ioab et populus, et quomodo administraretur bellum;
2SAM|11|8|et dixit David ad Uriam: " Descende in domum tuam et lava pedes tuos ". Et egressus est Urias de domo regis; secutusque est eum cibus regius.
2SAM|11|9|Dormivit autem Urias ante portam domus regiae cum aliis servis domini sui et non descendit ad domum suam.
2SAM|11|10|Nuntiatumque est David a dicentibus: " Non ivit Urias ad domum suam ". Et ait David ad Uriam: " Numquid non de via venisti? Quare non descendisti ad domum tuam? ".
2SAM|11|11|Et ait Urias ad David: " Arca et Israel et Iuda habitant in papilionibus, et dominus meus Ioab et servi domini mei super faciem terrae manent; et ego ingrediar domum meam, ut comedam et bibam et dormiam cum uxore mea? Per salutem tuam et per salutem animae tuae, non faciam rem hanc! ".
2SAM|11|12|Ait ergo David ad Uriam: " Mane hic etiam hodie, et cras dimittam te ". Mansit Urias in Ierusalem die illa et altera.
2SAM|11|13|Vocavit enim eum David, ut comederet coram se et biberet, et inebriavit eum. Qui egressus vespere dormivit in strato suo cum servis domini sui et in domum suam non descendit.
2SAM|11|14|Factum est ergo mane, et scripsit David epistulam ad Ioab misitque per manum Uriae
2SAM|11|15|scribens in epistula: " Ponite Uriam in prima acie, ubi fortissimum est proelium, et recedite ab eo, ut percussus intereat ".
2SAM|11|16|Igitur cum Ioab obsideret urbem, posuit Uriam in loco, quo sciebat viros esse fortissimos.
2SAM|11|17|Egressique viri de civitate bellabant adversum Ioab; et ceciderunt de populo, de servis David, et mortuus est etiam Urias Hetthaeus.
2SAM|11|18|Misit itaque Ioab et nuntiavit David omnia de proelio;
2SAM|11|19|praecepitque nuntio dicens: " Cum compleveris universos sermones proelii ad regem,
2SAM|11|20|si eum videris indignari et dixerit: "Quare accessistis ad urbem, ut proeliaremini? An ignorabatis quod desuper ex muro tela mittantur?
2SAM|11|21|Quis percussit Abimelech filium Ierobbaal? Nonne mulier misit super eum molam versatilem de muro, et mortuus est in Thebes? Quare iuxta murum accessistis?", dices: Etiam servus tuus Urias Hetthaeus occubuit ".
2SAM|11|22|Abiit ergo nuntius et venit et narravit David omnia, quae ei praeceperat Ioab.
2SAM|11|23|Et dixit nuntius ad David: " Quia praevaluerunt adversum nos viri et egressi sunt ad nos in agrum, nos, facto impetu, persecuti eos sumus usque ad portam civitatis.
2SAM|11|24|Et direxerunt iacula sagittarii ad servos tuos ex muro desuper; mortuique sunt de servis regis, quin etiam servus tuus Urias Hetthaeus mortuus est ".
2SAM|11|25|Et dixit David ad nuntium: " Haec dices Ioab: Non te affligat ista res; varius enim eventus est belli, et nunc hunc, nunc illum consumit gladius; corrobora proelium tuum adversus urbem, ut destruas eam. Et tu conforta eum ".
2SAM|11|26|Audivit autem uxor Uriae quod mortuus esset Urias vir suus et planxit eum.
2SAM|11|27|Transactoque luctu, misit David et introduxit eam domum suam, et facta est ei uxor peperitque ei filium. Et displicuit, quod fecerat David, coram Domino.
2SAM|12|1|Misit ergo Dominus Nathan ad David. Qui cum venisset ad eum, dixit ei: " Duo viri erant in civitate una, unus dives et alter pauper.
2SAM|12|2|Dives habebat oves et boves plurimos valde.
2SAM|12|3|Pauper autem nihil habebat omnino praeter ovem unam parvulam, quam emerat et nutrierat, et quae creverat apud eum cum filiis eius simul de pane illius comedens et de calice eius bibens et in sinu illius dormiens; eratque illi sicut filia.
2SAM|12|4|Cum autem peregrinus quidam venisset ad divitem, parcens ille sumere de ovibus et de bobus suis, ut exhiberet convivium peregrino illi, qui venerat ad se, tulit ovem viri pauperis et praeparavit cibos homini, qui venerat ad se ".
2SAM|12|5|Iratus autem indignatione David adversus hominem illum nimis dixit ad Nathan: " Vivit Dominus, quoniam filius mortis est vir, qui fecit hoc;
2SAM|12|6|ovem reddet in quadruplum, eo quod fecerit istud et non pepercerit ".
2SAM|12|7|Dixit autem Nathan ad David: " Tu es ille vir! Haec dicit Dominus, Deus Israel: Ego unxi te in regem super Israel et ego erui te de manu Saul;
2SAM|12|8|et dedi tibi domum domini tui et uxores domini tui in sinu tuo dedique tibi domum Israel et Iudae et, si parva sunt ista, adiciam tibi multo maiora.
2SAM|12|9|Quare ergo contempsisti verbum Domini, ut faceres malum in conspectu eius? Uriam Hetthaeum percussisti gladio et uxorem illius accepisti uxorem tibi et interfecisti eum gladio filiorum Ammon.
2SAM|12|10|Quam ob rem non recedet gladius de domo tua usque in sempiternum, eo quod despexeris me et tuleris uxorem Uriae Hetthaei, ut esset uxor tua.
2SAM|12|11|Itaque haec dicit Dominus: Ecce ego suscitabo super te malum de domo tua et tollam uxores tuas in oculis tuis et dabo proximo tuo, et dormiet cum uxoribus tuis in oculis solis huius.
2SAM|12|12|Tu enim fecisti abscondite; ego vero faciam istud in conspectu omnis Israel et in conspectu solis ".
2SAM|12|13|Et dixit David ad Nathan: " Peccavi Domino ". Dixitque Nathan ad David: Dominus quoque transtulit peccatum tuum; non morieris.
2SAM|12|14|Verumtamen quoniam blasphemare fecisti inimicos Domini propter hoc, filius, qui natus est tibi, morte morietur ".
2SAM|12|15|Et reversus est Nathan domum suam.Percussitque Dominus parvulum, quem peperat uxor Uriae David, et graviter aegrotavit;
2SAM|12|16|deprecatusque est David Dominum pro parvulo et ieiunavit David ieiunio et ingressus domum pernoctabat iacens super terram.
2SAM|12|17|Steterunt autem seniores domus eius iuxta eum cogentes eum, ut surgeret de terra; qui noluit neque comedit cum eis cibum.
2SAM|12|18|Accidit autem die septima, ut moreretur infans. Timueruntque servi David nuntiare ei quod mortuus esset parvulus; dixerunt enim: " Ecce, cum parvulus adhuc viveret, loquebamur ad eum, et non audiebat vocem nostram. Nunc quomodo dicemus: "Mortuus est puer"? Peius patrabit! ".
2SAM|12|19|Cum ergo vidisset David servos suos mussitantes, intellexit quod mortuus esset infantulus dixitque ad servos suos: " Num mortuus est puer?. Qui responderunt ei: " Mortuus est ".
2SAM|12|20|Surrexit igitur David de terra et lotus unctusque est; cumque mutasset vestem, ingressus est domum Domini et adoravit et venit in domum suam petivitque, ut ponerent ei panem, et comedit.
2SAM|12|21|Dixerunt autem ei servi sui: " Quid est quod fecisti? Propter infantem, cum adhuc viveret, ieiunasti et flebas; mortuo autem puero, surrexisti et comedisti panem ".
2SAM|12|22|Qui ait: " Propter infantem, dum adhuc viveret, ieiunavi et flevi. Dicebam enim: Quis scit, si forte miserebitur mei Dominus, et vivet infans?
2SAM|12|23|Nunc autem, quia mortuus est, quare ieiuno? Numquid potero revocare eum amplius? Ego vadam magis ad eum, ille vero non revertetur ad me ".
2SAM|12|24|Et consolatus est David Bethsabee uxorem suam ingressusque ad eam dormivit cum ea, quae genuit filium; et vocavit nomen eius Salomon. Et Dominus dilexit eum
2SAM|12|25|misitque in manu Nathan prophetae et vocavit nomen eius Iedidia (id est Amabilis Domino) propter Dominum.
2SAM|12|26|Igitur pugnavit Ioab contra Rabba filiorum Ammon et expugnavit urbem regiam.
2SAM|12|27|Misitque Ioab nuntios ad David dicens: " Dimicavi adversum Rabba et cepi urbem aquarum;
2SAM|12|28|nunc igitur congrega reliquam partem populi et obside civitatem et cape eam, ne, cum a me capta fuerit urbs, nomine meo vocetur ".
2SAM|12|29|Congregavit itaque David omnem populum et profectus est adversum Rabba; cumque dimicasset, cepit eam.
2SAM|12|30|Et tulit diadema Melchom de capite eius, pondo auri talentum, habens gemmam pretiosissimam, quod venit super caput David. Sed et praedam civitatis asportavit multam valde,
2SAM|12|31|populum quoque eius educens condemnavit ad operam lapicidinarum et ad secures et dolabras ferreas et transtulit eos ad opus laterum; sic fecit universis civitatibus filiorum Ammon. Et reversus est David et omnis exercitus Ierusalem.
2SAM|13|1|Factum est autem post haec, ut Absalom filii David soro rem speciosissimam, vocabulo Thamar, adamaret Amnon filius David.
2SAM|13|2|Et angustiatus est Amnon, ita ut aegrotaret propter amorem Thamar sororis suae, quia, cum esset virgo, difficile ei videbatur ut quippiam inhoneste ageret cum ea.
2SAM|13|3|Erat autem Amnonis amicus nomine Ionadab filius Samma fratris David, vir callidus valde.
2SAM|13|4|Qui dixit ad eum: " Quare sic attenuaris macie, fili regis, per singulos dies? Cur non indicas mihi? ". Dixitque ei Amnon: " Thamar sororem Absalom fratris mei amo ".
2SAM|13|5|Cui respondit Ionadab: " Cuba super lectulum tuum et languorem simula. Cumque venerit pater tuus, ut visitet te, dic ei: "Veniat, oro, Thamar soror mea, ut det mihi cibum et faciat in oculis meis pulmentum, ut videam et comedam de manu eius" ".
2SAM|13|6|Accubuit itaque Amnon et simulavit languorem. Cumque venisset rex ad visitandum eum, ait Amnon ad regem: " Veniat, obsecro, Thamar soror mea, ut faciat in oculis meis duas sorbitiunculas, et cibum capiam de manu eius.
2SAM|13|7|Misit ergo David ad Thamar domum dicens: " Veni in domum Amnon fratris tui et fac ei pulmentum ".
2SAM|13|8|Venitque Thamar in domum Amnon fratris sui; ille autem iacebat. Quae tollens farinam commiscuit et conficiens in oculis eius coxit sorbitiunculas.
2SAM|13|9|Tollensque sartaginem effudit, quod coxerat, et posuit coram eo. Noluit comedere; dixitque Amnon: " Eicite universos a me ". Cumque exissent omnes,
2SAM|13|10|dixit Amnon ad Thamar: " Infer cibum in conclave, ut vescar de manu tua. Tulit ergo Thamar sorbitiunculas, quas fecerat, et intulit ad Amnon fratrem suum in conclave.
2SAM|13|11|Cumque obtulisset ei cibum, apprehendit eam et ait: " Veni, cuba mecum, soror mea ".
2SAM|13|12|Quae respondit ei: " Noli, frater mi, noli opprimere me! Neque enim hoc fas est in Israel; noli facere stultitiam hanc.
2SAM|13|13|Et ego quo ibo in opprobrio meo? Et tu eris quasi unus de insipientibus in Israel; quin potius loquere ad regem, et non negabit me tibi ".
2SAM|13|14|Noluit autem acquiescere precibus eius, sed praevalens viribus oppressit eam et cubavit cum illa.
2SAM|13|15|Et exosam eam habuit Amnon magno odio nimis, ita ut maius esset odium, quo oderat eam, amore, quo ante dilexerat. Dixitque ei Amnon: " Surge, vade! ".
2SAM|13|16|Quae respondit ei: " Ne fiat, frater mi, quia maius est hoc malum, quod nunc agis adversum me expellens me, quam quod ante fecisti ". Et noluit audire eam;
2SAM|13|17|sed vocato puero, qui ministrabat ei, dixit: " Eice hanc a me foras et claude ostium post eam ".
2SAM|13|18|Quae induta erat talari tunica; huiusmodi enim filiae regis virgines palliis vestibus utebantur. Eiecit itaque eam minister illius foras clausitque fores post eam.
2SAM|13|19|Quae aspergens pulverem capiti suo, scissa talari tunica impositisque manibus super caput suum, ibat ingrediens et clamans.
2SAM|13|20|Dixit autem ei Absalom frater suus: " Num Amnon frater tuus fuit tecum? Sed nunc, soror, tace: frater tuus est; neque affligas cor tuum pro re hac. Mansit itaque Thamar desolata in domo Absalom fratris sui.
2SAM|13|21|Cum autem audisset rex David omnia haec, iratus est valde; et noluit contristare spiritum Amnon filii sui, quoniam diligebat eum, quia primogenitus erat ei.
2SAM|13|22|Porro non est locutus Absalom ad Amnon nec malum nec bonum; oderat enim Absalom Amnon, eo quod violasset Thamar sororem suam.
2SAM|13|23|Factum est autem post tempus biennii, ut tonderentur oves Absalom in Baalhasor, quae est iuxta Ephraim; et vocavit Absalom omnes filios regis.
2SAM|13|24|Venitque ad regem et ait ad eum: " Ecce tondentur oves servi tui; veniat, oro, rex cum servis suis ad servum tuum ".
2SAM|13|25|Dixitque rex ad Absalom: " Noli, fili mi, noli rogare, ut veniamus omnes et gravemus te ". Cum autem cogeret eum, et noluisset ire, benedixit ei.
2SAM|13|26|Et ait Absalom: " Si non vis venire, veniat, obsecro, nobiscum saltem Amnon frater meus ". Dixitque ad eum rex: " Cur vadet tecum? ".
2SAM|13|27|Coegit itaque eum Absalom, et dimisit cum eo Amnon et universos filios regis.Fecitque Absalom convivium quasi convivium regis.
2SAM|13|28|Praecepit autem Absalom pueris suis dicens: " Observate. Cum hilarior fuerit Amnon vino, et dixero vobis: Percutite Amnon et interficite eum!, nolite timere; ego enim sum, qui praecepi vobis. Roboramini et estote viri fortes ".
2SAM|13|29|Fecerunt ergo pueri Absalom adversum Amnon, sicut praeceperat eis Absalom; surgentesque omnes filii regis ascenderunt singuli mulos suos et fugerunt.
2SAM|13|30|Cumque adhuc pergerent in itinere, fama praevenit ad David dicens: " Percussit Absalom omnes filios regis, et non remansit ex eis saltem unus.
2SAM|13|31|Surrexit itaque rex et scidit vestimenta sua et prostravit se super terram; et omnes servi ipsius, qui assistebant ei, sciderunt vestimenta sua.
2SAM|13|32|Respondens autem Ionadab filius Samma fratris David dixit: " Ne aestimet dominus meus quod omnes pueri filii regis occisi sint; Amnon solus mortuus est, quoniam in ore Absalom hoc erat positum ex die, qua oppressit Thamar sororem eius.
2SAM|13|33|Nunc ergo ne ponat dominus meus rex super cor suum verbum istud dicens: Omnes filii regis occisi sunt", quoniam Amnon solus mortuus est ".
2SAM|13|34|Fugit autem Absalom.Et levavit puer speculator oculos suos et aspexit, et ecce populus multus veniebat per viam Oronaim ex latere montis in descensu; et venit speculator et nuntiavit regi dicens: " Video homines per viam Oronaim ".
2SAM|13|35|Dixit autem Ionadab ad regem: " Ecce filii regis adsunt! Iuxta verbum servi tui sic factum est ".
2SAM|13|36|Cumque cessasset loqui, apparuerunt et filii regis et intrantes levaverunt vocem suam et fleverunt; sed et rex et omnes servi eius fleverunt ploratu magno nimis.
2SAM|13|37|Porro Absalom fugiens abiit ad Tholmai filium Ammiud regem Gesur. Luxit ergo David filium suum cunctis diebus.
2SAM|13|38|Absalom autem, cum fugisset et venisset in Gesur, fuit ibi tribus annis.
2SAM|13|39|Cessavitque spiritus regis adversari Absalom, eo quod consolatus esset super Amnon interitu.
2SAM|14|1|Intellegens autem Ioab filius Sarviae quod cor regis ver sum esset ad Absalom,
2SAM|14|2|misit Thecuam et tulit inde mulierem sapientem dixitque ad eam: " Lugere te simula et induere veste lugubri et ne ungaris oleo, ut sis quasi mulier plurimo iam tempore lugens mortuum.
2SAM|14|3|Et ingredieris ad regem et loqueris ad eum sermones huiuscemodi ". Posuit autem Ioab verba in ore eius.
2SAM|14|4|Itaque, cum ingressa fuisset mulier Thecuites ad regem, cecidit coram eo super terram et adoravit et dixit: " Serva me, rex ".
2SAM|14|5|Et ait ad eam rex: " Quid causae habes? ". Quae respondit: " Heu, mulier vidua ego sum: mortuus est vir meus.
2SAM|14|6|Et ancillae tuae erant duo filii, qui rixati sunt adversum se in agro, nullusque erat, qui eos interveniens prohibere posset; et percussit alter alterum et interfecit eum.
2SAM|14|7|Et ecce consurgens universa cognatio adversum ancillam tuam dicit: Trade eum, qui percussit fratrem suum, ut occidamus eum pro anima fratris sui, quem interfecit, et deleamus heredem". Et quaerunt exstinguere scintillam meam, quae relicta est, ut non supersit viro meo nomen et reliquiae super terram ".
2SAM|14|8|Et ait rex ad mulierem: " Vade in domum tuam, et ego iubebo de te ".
2SAM|14|9|Dixitque mulier Thecuites ad regem: " In me, domine mi rex, iniquitas et in domum patris mei; rex autem et thronus eius sit innocens ".
2SAM|14|10|Et ait rex: " Qui contradixerit tibi, adduc eum ad me, et ultra non addet ut tangat te ".
2SAM|14|11|Quae ait: " Recordetur rex Domini Dei sui, ut non augeat ultor sanguinis perniciem, et nequaquam interficiant filium meum ". Qui ait: " Vivit Dominus, quia non cadet de capillis filii tui super terram ".
2SAM|14|12|Dixit ergo mulier: " Loquatur ancilla tua ad dominum meum regem verbum. Et ait: " Loquere ".
2SAM|14|13|Dixitque mulier: " Quare cogitasti istiusmodi rem contra populum Dei? Eo enim quod rex locutus est verbum istud, hoc est quasi delictum, quia rex noluit reducere eiectum suum.
2SAM|14|14|Omnes morimur et quasi aquae sumus, quae delabuntur in terram, quae non colliguntur; nec tamen vult perire Deus animam, sed retractat cogitans, ne penitus pereat, qui abiectus est.
2SAM|14|15|Nunc igitur veni, ut loquar ad regem dominum meum verbum hoc, quia populus terruit me. Et dixit ancilla tua: Loquar ad regem, si quo modo faciat rex verbum ancillae suae.
2SAM|14|16|Nam audiet rex, ut liberet ancillam suam de manu illius, qui vult delere me et filium meum simul de hereditate Dei.
2SAM|14|17|Dixit ergo ancilla tua: Fiat verbum domini mei regis mihi in quietem. Sicut enim angelus Dei, sic est dominus meus rex, ut audiat et discernat bonum et malum. Et Dominus Deus tuus sit tecum! ".
2SAM|14|18|Et respondens rex dixit ad mulierem: " Ne abscondas a me verbum, quod te interrogo ". Dixitque mulier: " Loquatur dominus meus rex ".
2SAM|14|19|Et ait rex: " Numquid manus Ioab tecum est in omnibus istis? ". Respondit mulier et ait: " Per salutem animae tuae, domine mi rex, nec ad dextram nec ad sinistram potest deviari ab omnibus his, quae locutus est dominus meus rex; servus enim tuus Ioab ipse praecepit mihi et ipse posuit in os ancillae tuae omnia verba haec;
2SAM|14|20|ut verterem figuram rei huius, servus tuus Ioab fecit istud. Tu autem, domine mi, sapiens es, sicut habet sapientiam angelus Dei, ut intellegas omnia, quae fiunt super terram ".
2SAM|14|21|Et ait rex ad Ioab: " Ecce hoc facio; vade igitur et revoca puerum Absalom ".
2SAM|14|22|Cadensque Ioab super faciem suam in terram adoravit et benedixit regi. Et dixit Ioab: " Hodie intellexit servus tuus quia inveni gratiam in oculis tuis, domine mi rex; fecisti enim sermonem servi tui ".
2SAM|14|23|Surrexit ergo Ioab et abiit in Gesur et adduxit Absalom in Ierusalem.
2SAM|14|24|Dixit autem rex: " Revertatur in domum suam et faciem meam non videat. Reversus est itaque Absalom in domum suam et faciem regis non vidit.
2SAM|14|25|Porro sicut Absalom vir non erat pulcher in omni Israel, qui valde laudaretur, a vestigio pedis usque ad verticem non erat in eo ulla macula.
2SAM|14|26|Et quando tondebatur capillus - semel autem in anno tondebatur, quia gravabat eum caesaries - ponderabat capillos capitis sui ducentis siclis pondere regio.
2SAM|14|27|Nati sunt autem Absalom filii tres et filia una, nomine Thamar, eleganti forma.
2SAM|14|28|Mansitque Absalom Ierusalem duobus annis et faciem regis non vidit.
2SAM|14|29|Misit itaque ad Ioab, ut mitteret eum ad regem; qui noluit venire ad eum. Cumque secundo misisset, et ille noluisset venire,
2SAM|14|30|dixit servis suis: " Videte agrum Ioab iuxta agrum meum habentem messem hordei; ite igitur et succendite eum igni ". Succenderunt ergo servi Absalom segetem igni. Et venientes servi Ioab, scissis vestibus suis, dixerunt: " Succenderunt servi Absalom agrum igni! ".
2SAM|14|31|Surrexitque Ioab et venit ad Absalom in domum eius et dixit: " Quare succenderunt servi tui segetem meam igni? ".
2SAM|14|32|Et respondit Absalom ad Ioab: " Misi ad te obsecrans, ut venires ad me, et mitterem te ad regem, ut diceres ei: "Quare veni de Gesur? Melius mihi erat adhuc ibi esse". Obsecro ergo, ut videam faciem regis; quod si est in me iniquitas, interficiat me ".
2SAM|14|33|Ingressus Ioab ad regem nuntiavit ei. Vocatusque Absalom intravit ad regem et adoravit super faciem in terra coram eo; osculatusque est rex Absalom.
2SAM|15|1|Post haec fecit sibi Absalom currus et equos et quinqua ginta viros, qui praecederent eum.
2SAM|15|2|Et mane consurgens Absalom stabat iuxta viam portae; et omnem virum, qui habebat negotium, ut veniret ad regis iudicium, vocabat Absalom ad se et dicebat: " De qua civitate es tu? ". Qui respondens aiebat: " Ex una tribu Israel ego sum servus tuus ".
2SAM|15|3|Respondebatque ei Absalom: " Vide, sermones tui sunt boni et iusti, sed non est qui te audiat constitutus a rege ". Dicebatque Absalom:
2SAM|15|4|" Quis me constituat iudicem in terra, ut ad me veniant omnes, qui habent negotium iudicandum, et iustificem eos? ".
2SAM|15|5|Sed et cum accederet ad eum homo, ut se prostraret coram illo, extendebat manum suam et apprehendens osculabatur eum.
2SAM|15|6|Faciebatque hoc omni Israel, qui veniebat ad iudicium, ut audiretur a rege, et sollicitabat corda virorum Israel.
2SAM|15|7|Post quattuor autem annos dixit Absalom ad regem: " Vadam, quaeso, et reddam in Hebron vota mea, quae vovi Domino.
2SAM|15|8|Votum enim vovit servus tuus, cum esset in Gesur Syriae, dicens: Si reduxerit me Dominus in Ierusalem, sacrificabo Domino ".
2SAM|15|9|Dixitque ei rex. " Vade in pace ". Et surrexit et abiit in Hebron.
2SAM|15|10|Misit autem Absalom exploratores in universas tribus Israel dicens: " Statim ut audieritis clangorem bucinae, dicite: "Factus est rex Absalom in Hebron" ".
2SAM|15|11|Porro cum Absalom ierunt ducenti viri de Ierusalem vocati, euntes simplici corde et causam penitus ignorantes.
2SAM|15|12|Accersivit quoque Absalom, cum immolaret victimas, Achitophel Gilonitem consiliarium David de civitate sua Gilo. Et facta est coniuratio valida; populusque concurrens augebatur cum Absalom.
2SAM|15|13|Venit igitur nuntius ad David dicens: " Toto corde universus Israel sequitur Absalom ".
2SAM|15|14|Et ait David servis suis, qui erant cum eo in Ierusalem: " Surgite, fugiamus; neque enim erit nobis effugium a facie Absalom. Festinate egredi, ne festinans occupet nos et impellat super nos ruinam et percutiat civitatem in ore gladii ".
2SAM|15|15|Dixeruntque servi regis ad eum: " In omnibus, quaecumque elegerit dominus noster rex, ecce servi tui sumus ".
2SAM|15|16|Egressus est ergo rex et universa domus eius post eum et dereliquit rex decem mulieres concubinas ad custodiendam domum.
2SAM|15|17|Egressusque rex et omnis populus post eum steterunt ad ultimam domum.
2SAM|15|18|Et universi servi eius transierunt iuxta eum; et omnes Cherethi et Phelethi et omnes Getthaei, sescenti viri, qui secuti eum fuerant de Geth, transierunt coram rege.
2SAM|15|19|Dixit autem rex ad Ethai Getthaeum: " Cur venis etiam tu nobiscum? Revertere et habita cum rege, quia alienigena es, immo et exsul de loco tuo.
2SAM|15|20|Heri venisti, et hodie compellam te vagari nobiscum, cum ego vadam, quo iturus sum? Revertere et reduc tecum fratres tuos, et Dominus faciat tecum misericordiam et veritatem ".
2SAM|15|21|Et respondit Ethai regi dicens: " Vivit Dominus et vivit dominus meus rex, in quocumque loco fuerit dominus meus rex, sive ad mortem sive ad vitam, ibi erit servus tuus ".
2SAM|15|22|Et ait David Ethai: " Veni et transi ". Et transivit Ethai Getthaeus et omnes viri eius et omnes parvuli, qui cum eo erant.
2SAM|15|23|Omnisque terra flebat voce magna, et universus populus transibat. Rex quoque transgrediebatur torrentem Cedron, et cunctus populus incedebat contra viam deserti.
2SAM|15|24|Venit autem et Sadoc et universi Levitae cum eo portantes arcam foederis Dei; et deposuerunt arcam Dei. Et sacrificavit Abiathar, donec omnis populus egressus fuerat de civitate.
2SAM|15|25|Et dixit rex ad Sadoc: " Reporta arcam Dei in urbem. Si invenero gratiam in oculis Domini, reducet me et ostendet mihi eam et habitationem suam.
2SAM|15|26|Si autem dixerit: "Non places mihi", praesto sum: faciat, quod bonum est coram se ".
2SAM|15|27|Et dixit rex ad Sadoc sacerdotem: " Videsne? Revertere in civitatem in pace; et Achimaas filius tuus et Ionathan filius Abiathar, duo filii vestri sint vobiscum.
2SAM|15|28|Ecce ego morabor ad vada deserti, donec veniat sermo a vobis indicans mihi ".
2SAM|15|29|Reportaverunt igitur Sadoc et Abiathar arcam Dei Ierusalem et manserunt ibi.
2SAM|15|30|Porro David ascendebat clivum Olivarum scandens et flens, operto capite et nudis pedibus incedens; sed et omnis populus, qui erat cum eo, operto capite ascendebat plorans.
2SAM|15|31|Nuntiatum est autem David quod et Achitophel esset in coniuratione cum Absalom; dixitque David: " Infatua, quaeso, Domine, consilium Achitophel.
2SAM|15|32|Cumque ascendisset David summitatem montis, in quo adorabatur Deus, ecce occurrit ei Chusai Arachites, scissa veste et terra pleno capite.
2SAM|15|33|Et dixit ei David: " Si veneris mecum, eris mihi oneri;
2SAM|15|34|Si autem in civitatem revertaris et dixeris Absalom: "Servus tuus ego, rex, ero; servus patris tui ego fui prius, nunc autem ego sum servus tuus", dissipabis mihi consilium Achitophel.
2SAM|15|35|Habes autem tecum Sadoc et Abiathar sacerdotes; et omne verbum, quodcumque audieris de domo regis, indicabis Sadoc et Abiathar sacerdotibus.
2SAM|15|36|Sunt autem cum eis duo filii eorum: Achimaas Sadoc et Ionathan Abiathar; et mittetis per eos ad me omne verbum, quod audieritis ".
2SAM|15|37|Veniente ergo Chusai amico David in civitatem, Absalom quoque ingressus est Ierusalem.
2SAM|16|1|Cumque David transisset paululum montis verticem, apparuit Siba puer Meribbaal in occursum eius cum duobus asinis stratis, qui onerati erant ducentis panibus et centum alligaturis uvae passae et centum fasciculis fructuum aestivorum et utre vini.
2SAM|16|2|Et dixit rex Sibae: " Quid sibi volunt haec? ". Responditque Siba: " Asini domesticis regis ad sedendum; et panes et fructus aestivi ad vescendum pueris tuis; vinum autem, ut bibat, si quis defecerit in deserto.
2SAM|16|3|Et ait rex: " Ubi est filius domini tui? ". Responditque Siba regi: " Remansit in Ierusalem dicens: "Hodie restituet mihi domus Israel regnum patris mei" ".
2SAM|16|4|Et ait rex Sibae: " Ecce, tua sint omnia, quae fuerunt Meribbaal ". Dixitque Siba: " Adoro; inveniam gratiam coram te, domine mi rex ".
2SAM|16|5|Venit ergo rex David usque Bahurim, et ecce egrediebatur inde vir de cognatione domus Saul nomine Semei filius Gera; procedebat egrediens et maledicens
2SAM|16|6|mittebatque lapides contra David et contra universos servos regis David. Omnis autem populus et universi viri fortissimi a dextro et sinistro latere regis incedebant.
2SAM|16|7|Ita autem loquebatur Semei, cum malediceret regi: " Egredere, egredere, vir sanguinum et vir Belial!
2SAM|16|8|Reddidit tibi Dominus universum sanguinem domus Saul, quoniam invasisti regnum eius; et dedit Dominus regnum in manu Absalom filii tui; et ecce premunt te mala tua, quoniam vir sanguinum es ".
2SAM|16|9|Dixit autem Abisai filius Sarviae regi: " Quare maledicit canis hic mortuus domino meo regi? Vadam et amputabo caput eius ".
2SAM|16|10|Et ait rex: "Quid mihi et vobis filii Sarviae? Si maledicit, et si Dominus praecepit ei, ut malediceret David, quis est qui audeat dicere: Quare sic fecisti?" ".
2SAM|16|11|Et ait rex Abisai et universis servis suis: " Ecce filius meus, qui egressus est de visceribus meis, quaerit animam meam; quanto magis nunc iste filius Beniaminita. Dimittite eum, ut maledicat iuxta praeceptum Domini.
2SAM|16|12|Fortasse respiciet Dominus afflictionem meam et reddet mihi bonum pro maledictione hac hodierna ".
2SAM|16|13|Ambulabat itaque David et socii eius per viam; Semei autem per iugum montis ex latere gradiebatur maledicens et mittens lapides adversum eum terramque spargens.
2SAM|16|14|Venit itaque rex et universus populus cum eo lassus usque ad aquas, et refocillati sunt ibi.
2SAM|16|15|Absalom autem et omnis populus eius, viri Israel, ingressi sunt Ierusalem, sed et Achitophel cum eo.
2SAM|16|16|Cum autem venisset Chusai Arachites amicus David ad Absalom, locutus est ad eum: " Vivat rex! Vivat rex! ".
2SAM|16|17|Ad quem Absalom: "Haec est, inquit, gratia tua ad amicum tuum? Quare non isti cum amico tuo? ".
2SAM|16|18|Responditque Chusai ad Absalom: " Nequaquam; quia, quem elegit Dominus, et hic populus et omnis Israel, illius ero et cum eo manebo.
2SAM|16|19|Sed, ut et hoc inferam, cui ego serviturus sum? Nonne filio regis? Sicut parui patri tuo, sic parebo et tibi ".
2SAM|16|20|Dixit autem Absalom ad Achitophel: " Inite consilium quid agere debeamus ".
2SAM|16|21|Et ait Achitophel ad Absalom: " Ingredere ad concubinas patris tui, quas dimisit ad custodiendam domum; ut, cum audierit omnis Israel quod foedaveris patrem tuum, roborentur manus omnium, qui tecum sunt ".
2SAM|16|22|Tetenderunt igitur Absalom tabernaculum in solario; ingressusque est ad concubinas patris sui coram universo Israel.
2SAM|16|23|Consilium autem Achitophel, quod dabat in diebus illis, quasi si quis consuleret Deum; sic erat omne consilium Achitophel, et cum esset cum David et cum esset cum Absalom.
2SAM|17|1|Dixitque Achitophel ad Ab salom: " Eligam mihi duode cim milia virorum et consurgens persequar David hac nocte
2SAM|17|2|et irruens super eum, quippe qui lassus est et solutis manibus, terrebo eum. Cumque fugerit omnis populus, qui cum eo est, percutiam regem desolatum
2SAM|17|3|et reducam universum populum ad te, sicut revertitur sponsa ad virum suum; unius solummodo viri animam quaeris, et omnis populus erit in pace.
2SAM|17|4|Placuitque sermo eius Absalom et cunctis maioribus natu Israel.
2SAM|17|5|Ait autem Absalom: " Vocate et Chusai Arachiten, et audiamus quid etiam ipse dicat ".
2SAM|17|6|Cumque venisset Chusai ad Absalom, ait Absalom ad eum: " Huiuscemodi sermonem locutus est Achitophel; verbum eius facere debemus an non? Tu loquere ".
2SAM|17|7|Et dixit Chusai ad Absalom: " Non bonum consilium, quod dedit Achitophel hac vice ".
2SAM|17|8|Et rursum intulit Chusai: " Tu nosti patrem tuum et viros, qui cum eo sunt, esse fortissimos et amaro animo, veluti ursa in saltu catulis orbata; sed et pater tuus vir bellator est nec morabitur cum populo:
2SAM|17|9|ecce nunc latitat in aliqua fovea aut in aliquo alio loco. Et, cum ceciderit unus quilibet in principio, certo audient et dicent: "Facta est plaga in populo, qui sequitur Absalom".
2SAM|17|10|Et fortissimus quoque, cuius cor est quasi leonis, pavore solvetur; scit enim omnis Israel fortem esse patrem tuum et robustos omnes, qui cum eo sunt.
2SAM|17|11|Sed hoc mihi videtur rectum esse consilium: congregetur ad te universus Israel a Dan usque Bersabee, quasi arena maris innumerabilis, et tu ipse gradieris in proelium;
2SAM|17|12|et irruemus super eum, in quocumque loco fuerit inventus, et operiemus eum sicut cadere solet ros super terram; et non remanebit de eo et de omnibus viris, qui cum eo sunt, ne unus quidem.
2SAM|17|13|Quod si urbem aliquam fuerit ingressus, applicabit omnis Israel civitati illi funes, et trahemus eam in torrentem, ut non reperiatur nec calculus quidem ex ea ".
2SAM|17|14|Dixitque Absalom et omnis vir Israel: " Melius consilium Chusai Arachitae consilio Achitophel ". Dominus enim statuerat dissipare consilium Achitophel utile, ut induceret Dominus super Absalom malum.
2SAM|17|15|Et ait Chusai Sadoc et Abiathar sacerdotibus: " Hoc et hoc modo consilium dedit Achitophel Absalom et senibus Israel, et ego tale et tale dedi consilium;
2SAM|17|16|nunc ergo mittite cito et nuntiate David dicentes: "Ne moreris nocte hac ad vada deserti, sed absque dilatione transgredere, ne absorbeatur rex et omnis populus, qui cum eo est" ".
2SAM|17|17|Ionathan autem et Achimaas stabant iuxta fontem Rogel; abiit ancilla et nuntiavit eis, et illi profecti sunt, ut referrent ad regem David nuntium; non enim poterant introire civitatem, ne viderentur.
2SAM|17|18|Vidit autem eos quidam iuvenis et indicavit Absalom; illi vero concito gradu profecti ingressi sunt domum cuiusdam viri in Bahurim, qui habebat puteum in vestibulo suo, et descenderunt in eum.
2SAM|17|19|Tulit autem mulier et expandit velamen super os putei et sparsit super illud ptisanas, et sic res latuit.
2SAM|17|20|Cumque venissent servi Absalom ad mulierem in domum, dixerunt: " Ubi est Achimaas et Ionathan? ". Et respondit eis mulier: " Transierunt hinc ad aquas ". At hi, qui quaerebant, cum non repperissent, reversi sunt Ierusalem.
2SAM|17|21|Cumque abissent, ascenderunt illi de puteo et pergentes nuntiaverunt regi David atque dixerunt: " Surgite et transite cito fluvium, quoniam huiuscemodi dedit consilium contra vos Achitophel ".
2SAM|17|22|Surrexit ergo David et omnis populus, qui erat cum eo, et transierunt Iordanem, donec dilucesceret; et ne unus quidem residuus fuit, qui non transisset fluvium.
2SAM|17|23|Porro Achitophel videns quod non fuisset factum consilium suum, stravit asinum suum et surrexit et abiit in domum suam in civitatem suam et, disposita domo sua, laqueo se suspendit et interiit; et sepultus est in sepulcro patris sui.
2SAM|17|24|David autem venit in Mahanaim, et Absalom transivit Iordanem, ipse et omnis vir Israel cum eo.
2SAM|17|25|Amasam vero constituerat Absalom pro Ioab super exercitum; Amasa autem erat filius viri, qui vocabatur Iether Ismaelites, qui ingressus est ad Abigail filiam Isai sororem Sarviae, quae fuit mater Ioab.
2SAM|17|26|Et castrametatus est Israel cum Absalom in terra Galaad.
2SAM|17|27|Cumque venisset David in Mahanaim, Sobi filius Naas de Rabba filiorum Ammon et Machir filius Ammiel de Lodabar et Berzellai Galaadites de Rogelim
2SAM|17|28|obtulerunt ei stratoria et tapetia et pelves et vasa fictilia, frumentum et hordeum et farinam, frixum cicer et fabam et lentem
2SAM|17|29|et mel et butyrum, oves et pingues vitulos; dederuntque David et populo, qui cum eo erat, ad vescendum; suspicati enim sunt populum fame et siti fuisse fatigatum in deserto.
2SAM|18|1|Igitur, recensito David populo suo, constituit super eum tribunos et centuriones.
2SAM|18|2|Et divisit David populum in tres partes: tertiam partem sub manu Ioab et tertiam sub manu Abisai filii Sarviae fratris Ioab et tertiam in manu Ethai, qui erat de Geth. Dixitque rex ad populum: " Egrediar et ego vobiscum ".
2SAM|18|3|Et respondit populus: " Non exibis. Sive enim fugerimus, non magnopere ad eos de nobis pertinebit; et si media pars ceciderit e nobis, non satis curabunt, sed tu unus pro decem milibus computaris. Melius est igitur, ut sis nobis ex urbe praesidio ".
2SAM|18|4|Ad quos rex ait: " Quod vobis rectum videtur, hoc faciam ". Stetit ergo rex iuxta portam; egrediebaturque populus per turmas suas centeni et milleni.
2SAM|18|5|Et praecepit rex Ioab et Abisai et Ethai dicens: " Leniter mihi agite cum puero Absalom ". Et omnis populus audiebat praecipientem regem cunctis principibus pro Absalom.
2SAM|18|6|Itaque egressus est populus in campum contra Israel, et factum est proelium in saltu Ephraim.
2SAM|18|7|Et caesus est ibi populus Israel ab exercitu David; factaque est ibi plaga magna in die illa viginti milium hominum.
2SAM|18|8|Fuit autem ibi proelium dispersum super faciem omnis terrae; et multo plures erant, quos saltus consumpserat de populo, quam hi, quos voraverat gladius in die illa.
2SAM|18|9|Accidit autem, ut occurreret Absalom servis David sedens mulo; cumque ingressus fuisset mulus subter condensam quercum et magnam, adhaesit caput eius quercui, et mansit suspensus inter caelum et terram; mulus, cui insederat, pertransivit.
2SAM|18|10|Vidit autem hoc quispiam et nuntiavit Ioab dicens: " Vidi Absalom pendere de quercu ".
2SAM|18|11|Et ait Ioab viro, qui nuntiaverat ei: " Si vidisti, quare non confodisti eum in terra? Ego vero dedissem tibi decem argenti siclos et unum balteum ".
2SAM|18|12|Qui dixit ad Ioab: " Et si appenderes in manibus meis mille argenteos, nequaquam mitterem manum meam in filium regis. Audientibus enim nobis, praecepit rex tibi et Abisai et Ethai dicens: "Custodite, quisquis sit, puerum Absalom!".
2SAM|18|13|Sed et si fecissem contra animam meam infideliter, nequaquam hoc regem latere potuisset, et tu stares ex adverso ".
2SAM|18|14|Et ait Ioab: " Non ita praestolabor coram te ". Tulit ergo tres lanceas in manu sua et infixit eas in corde Absalom, cum adhuc palpitaret haerens in quercu;
2SAM|18|15|et cucurrerunt decem iuvenes armigeri Ioab et percutientes interfecerunt eum.
2SAM|18|16|Cecinit autem Ioab bucina, et destitit populus persequi fugientem Israel, quia Ioab retinuit populum.
2SAM|18|17|Et tulerunt Absalom et proiecerunt eum in saltu in foveam grandem et erexerunt super eum acervum lapidum magnum nimis; omnis autem Israel fugit in tabernacula sua.
2SAM|18|18|Porro Absalom erexerat sibi, cum adhuc viveret, lapidem, qui est in valle Regis; dixerat enim: " Non habeo filium, qui memoriam servabit nominis mei ". Vocavitque titulum nomine suo, et appellatur Manus Absalom usque ad hanc diem.
2SAM|18|19|Achimaas autem filius Sadoc ait: " Curram et nuntiabo regi, quia iudicium fecerit ei Dominus de manu inimicorum eius ".
2SAM|18|20|Ad quem Ioab dixit: " Non es vir boni nuntii in hac die, sed nuntiabis in alia; hodie enim non nuntiabis bona, eo quod filius regis est mortuus.
2SAM|18|21|Et ait Ioab Aethiopi: " Vade et nuntia regi, quae vidisti ". Adoravit Aethiops Ioab et cucurrit.
2SAM|18|22|Rursus autem Achimaas filius Sadoc dixit ad Ioab: " Quidquid evenerit, etiam ego curram post Aethiopem! ". Dixitque Ioab: " Quid vis currere, fili mi? Non erit tibi merces pro bono nuntio ".
2SAM|18|23|Qui respondit: " Quidquid evenerit, curram ". Et ait ei: " Curre! ". Currens ergo Achimaas per viam regionis transivit Aethiopem.
2SAM|18|24|David autem sedebat inter duas portas; speculator vero, qui ierat in solarium portae super murum, elevans oculos vidit hominem currentem solum
2SAM|18|25|et exclamans indicavit regi. Dixitque rex: " Si solus est, bonus est nuntius in ore eius ". Properante autem illo et accedente propius,
2SAM|18|26|vidit speculator hominem alterum currentem, et clamavit speculator ad ianitorem: " Apparet mihi homo currens solus ". Dixitque rex: " Et iste bonus est nuntius ".
2SAM|18|27|Speculator autem: " Contemplor, ait, cursum prioris quasi cursum Achimaas filii Sadoc ". Et ait rex: " Vir bonus est et nuntium portans bonum venit ".
2SAM|18|28|Clamans autem Achimaas dixit ad regem: " Pax! ". Et adorans regem pronus in terram ait: " Benedictus Dominus Deus tuus, qui conclusit homines, qui levaverunt manus suas contra dominum meum regem! ".
2SAM|18|29|Et ait rex: " Estne pax puero Absalom? ". Dixitque Achimaas: " Vidi tumultum magnum, cum mitteret Ioab servum regis et me servum tuum, sed nescio quid fuerit ".
2SAM|18|30|Ad quem rex: " Recede, ait, et sta illic ". Cumque ille recessisset et staret,
2SAM|18|31|apparuit Aethiops et veniens ait: " Bonum apporto nuntium, domine mi rex; iudicavit enim pro te Dominus hodie salvans te de manu omnium, qui surrexerunt contra te ".
2SAM|18|32|Dixit autem rex ad Aethiopem: " Estne pax puero Absalom? ". Cui respondens Aethiops: " Fiant, inquit, sicut puer inimici domini mei regis et universi, qui consurrexerunt adversus eum in malum! ".
2SAM|19|1|Contremuit itaque rex et ascendit cenaculum portae et flevit. Et sic loquebatur vadens: " Fili mi Absalom, fili mi, fili mi Absalom! Quis mihi tribuat, ut ego moriar pro te? Absalom fili mi, fili mi! ".
2SAM|19|2|Nuntiatum est autem Ioab quod rex fleret et lugeret filium suum.
2SAM|19|3|Et versa est victoria in die illa in luctum omni populo; audivit enim populus in die illa dici: " Dolet rex super filio suo ".
2SAM|19|4|Et furtim ingressus est populus in die illa civitatem, quomodo reverti solet populus confusus, cum fugit de proelio.
2SAM|19|5|Porro rex operuit vultum suum et clamabat voce magna: " Fili mi Absalom, Absalom fili mi, fili mi! ".
2SAM|19|6|Ingressus ergo Ioab ad regem in domo dixit: " Confudisti hodie vultus omnium servorum tuorum, qui salvam fecerunt animam tuam hodie et animam filiorum tuorum et filiarum tuarum et animam uxorum tuarum et animam concubinarum tuarum.
2SAM|19|7|Diligis odientes te et odio habes diligentes te. Ostendisti hodie quia non curas de ducibus tuis et de servis tuis; et vere cognovi modo quia, si Absalom viveret, et nos omnes occubuissemus, tunc placeret tibi.
2SAM|19|8|Nunc igitur surge et procede et loquere ad cor servorum tuorum; iuro enim tibi per Dominum quod si non exieris, ne unus quidem remansurus sit tecum nocte hac, et peius erit hoc tibi quam omnia mala, quae venerunt super te ab adulescentia tua usque in praesens ".
2SAM|19|9|Surrexit ergo rex et sedit in porta, et omni populo nuntiatum est quod rex sederet in porta; venitque universa multitudo coram rege.Israel autem fugerat in tabernacula sua.
2SAM|19|10|Omnis quoque populus certabat in cunctis tribubus Israel dicens: " Rex liberavit nos de manu inimicorum nostrorum, ipse salvavit nos de manu Philisthinorum; et nunc fugit de terra ab Absalom.
2SAM|19|11|Absalom autem, quem unximus super nos, mortuus est in bello. Quare nunc siletis et non reducitis regem? ".
2SAM|19|12|Sermo autem omnis Israel pervenerat ad regem in domo eius. Tunc rex David misit ad Sadoc et Abiathar sacerdotes dicens: " Loquimini ad maiores natu Iudae dicentes: Cur estis novissimi ad reducendum regem in domum suam?
2SAM|19|13|Fratres mei vos, os meum et caro mea vos; quare novissimi reducitis regem?
2SAM|19|14|Et Amasae dicite: Nonne os meum es et caro mea? Haec faciat mihi Deus et haec addat, si non magister militiae fueris coram me omni tempore pro Ioab! ".
2SAM|19|15|Et inclinavit cor omnium virorum Iudae quasi viri unius; miseruntque ad regem dicentes: " Revertere tu et omnes servi tui ".
2SAM|19|16|Et reversus est rex et venit usque ad Iordanem; et Iuda venit in Galgala, ut occurreret regi et traduceret eum Iordanem.
2SAM|19|17|Festinavit autem Semei filius Gera Beniaminita de Bahurim et descendit cum viris Iudae in occursum regis David;
2SAM|19|18|mille viri de Beniamin et Siba puer de domo Saul et quindecim filii eius ac viginti servi erant cum eo. Irruperant autem Iordanem iam ante regem
2SAM|19|19|et transierant vada, ut traducerent domum regis et facerent iuxta placitum eius. Semei autem filius Gera prostratus coram rege, cum transiturus esset Iordanem,
2SAM|19|20|dixit ad eum: " Ne reputes mihi, domine mi, iniquitatem neque memineris iniuriam servi tui in die, qua egressus es, domine mi rex, de Ierusalem; neque ponas, rex, in corde tuo.
2SAM|19|21|Agnosco enim servus tuus peccatum meum et idcirco hodie primus veni de omni domo Ioseph descendique in occursum domini mei regis ".
2SAM|19|22|Respondens vero Abisai filius Sarviae dixit: " Numquid non occidetur Semei, pro hoc quia maledixit christo Domini? ".
2SAM|19|23|Et ait David: " Quid mihi et vobis, filii Sarviae, quia efficimini mihi hodie in satan? Ergone hodie interficietur vir in Israel? An ignoro hodie me factum regem super Israel? ".
2SAM|19|24|Et ait rex Semei: " Non morieris! ". Iuravitque ei.
2SAM|19|25|Meribbaal quoque filius Saul descendit in occursum regis; non laverat pedes nec circumcidit ungues nec totonderat barbam vestesque suas non laverat a die, qua egressus fuerat rex, usque ad diem reversionis eius in pace.
2SAM|19|26|Cumque de Ierusalem occurrisset regi, dixit ei rex: " Quare non venisti mecum, Meribbaal? ".
2SAM|19|27|Qui respondens ait: " Domine mi rex, servus meus decepit me! Nam dixeram ei ego famulus tuus: Sternere faciam mihi asinum et ascendens abibo cum rege; claudus enim sum servus tuus.
2SAM|19|28|Insuper et fraudulenter accusavit me servum tuum ad te dominum meum regem. Tu autem, domine mi rex, sicut angelus Dei es; fac, quod placitum est tibi.
2SAM|19|29|Neque enim fuit domus patris mei nisi morti obnoxia domino meo regi; tu autem posuisti me servum tuum inter convivas mensae tuae. Quid ultra igitur habeo iustitiae, ut vociferer ad regem? ".
2SAM|19|30|Ait ergo ei rex: " Quid ultra loqueris? Dixi: Tu et Siba dividite possessiones ".
2SAM|19|31|Responditque Meribbaal regi: " Etiam cuncta accipiat, postquam reversus est dominus meus rex pacifice in domum suam! ".
2SAM|19|32|Berzellai quoque Galaadites descenderat de Rogelim et traduxit regem Iordanem, ut dimitteret eum ad Iordanem.
2SAM|19|33|Erat autem Berzellai Galaadites senex valde, id est octogenarius; et ipse praebuerat alimenta regi, cum moraretur in Mahanaim; erat quippe vir dives nimis.
2SAM|19|34|Dixit itaque rex ad Berzellai: " Veni mecum et praebebo tibi alimenta apud me in Ierusalem ".
2SAM|19|35|Et ait Berzellai ad regem: " Quot sunt dies annorum vitae meae, ut ascendam cum rege Ierusalem?
2SAM|19|36|Octogenarius sum hodie; numquid vigent sensus mei ad discernendum suave aut amarum? Aut delectare potest servum tuum cibus et potus? Vel audire ultra possum vocem cantorum atque cantricum? Quare servus tuus esset ultra oneri domino meo regi?
2SAM|19|37|Paululum procedam famulus tuus ab Iordane tecum. Et cur dabit rex mihi hanc vicissitudinem?
2SAM|19|38|Sed obsecro, ut revertar servus tuus et moriar in civitate mea iuxta sepulcrum patris mei et matris meae. Sed ecce servus tuus Chamaam; ipse vadat tecum, domine mi rex, et fac ei, quod tibi bonum videtur ".
2SAM|19|39|Dixitque rex: " Mecum transeat Chamaam, et ego faciam ei, quidquid tibi placuerit; et omne, quod petieris a me, impetrabis ".
2SAM|19|40|Cumque transisset universus populus et rex Iordanem, osculatus est rex Berzellai et benedixit ei; et ille reversus est in locum suum.
2SAM|19|41|Transivit ergo rex in Galgala, et Chamaam cum eo. Omnis autem populus Iudae traduxerat regem, et etiam media pars populi Israel.
2SAM|19|42|Et ecce omnes viri Israel concurrentes ad regem dixerunt ei: " Quare te furati sunt fratres nostri viri Iudae et traduxerunt regem et domum eius Iordanem omnesque viros David cum eo? ".
2SAM|19|43|Et respondit omnis vir Iudae ad virum Israel: " Quia propior mihi est rex. Cur irasceris super hac re? Numquid comedimus aliquid ex rege, aut munera nobis data sunt? ".
2SAM|19|44|Et respondit vir Israel ad virum Iudae et ait: " Decem partes mihi sunt in rege et ideo etiam in David. Ego sum potior te; cur contempsisti me? Et non ego prior locutus sum, ut reducerem regem meum? ". Durius autem responderunt viri Iudae viris Israel.
2SAM|20|1|Accidit quoque, ut ibi esset vir Belial nomine Seba filius Bochri Beniaminita; et cecinit bucina et ait: Non est nobis pars in David,neque hereditas in filio Isai!Vir Israel, in tabernacula tua! ".
2SAM|20|2|Et separatus est omnis vir Israel a David secutusque est Seba filium Bochri; viri autem Iudae adhaeserunt regi suo a Iordane usque Ierusalem.
2SAM|20|3|Cumque venisset rex in domum suam Ierusalem, tulit decem mulieres concubinas, quas dereliquerat ad custodiendam domum, et tradidit eas in custodiam alimenta eis praebens. Et non est ingressus ad eas, sed erant clausae usque ad diem mortis suae in viduitate viventes.
2SAM|20|4|Dixit autem rex Amasae: " Convoca mihi omnes viros Iudae in diem tertium et tu adesto praesens ".
2SAM|20|5|Abiit ergo Amasa, ut convocaret Iudam; et moratus est ultra tempus, quod ei constituerat.
2SAM|20|6|Ait autem David ad Abisai: " Nunc magis afflicturus est nos Seba filius Bochri quam Absalom; tolle igitur servos domini tui et persequere eum, ne inveniat civitates munitas et effugiat nos ".
2SAM|20|7|Egressi sunt ergo cum eo viri Ioab, Cherethi quoque et Phelethi et omnes fortissimi; exierunt de Ierusalem ad persequendum Seba filium Bochri.
2SAM|20|8|Cumque illi essent iuxta lapidem grandem, qui est in Gabaon, Amasa venerat ante eos. Porro Ioab accinctus erat habitu suo, et in cingulo super lumbos gladius absconditus erat, qui levi motu ex vagina in manum suam cecidit.
2SAM|20|9|Dixitque Ioab ad Amasam: " Estne pax tibi, mi frater? ". Et tenuit manu dextera mentum Amasae, ut oscularetur eum.
2SAM|20|10|Porro Amasa non observavit gladium in manu Ioab, qui percussit eum in inguine et effudit intestina eius in terram, nec secundum vulnus apposuit; et mortuus est. Ioab autem et Abisai frater eius persecuti sunt Seba filium Bochri.
2SAM|20|11|Interea quidam de pueris Ioab stetit iuxta cadaver Amasae et dixit: " Qui esse vult cum Ioab et pro David, sequatur Ioab! ".
2SAM|20|12|Amasa autem conspersus sanguine iacebat in media via. Vidit hoc vir quod subsisteret omnis populus ad videndum eum; et amovit Amasam de via in agrum operuitque eum vestimento, cum videret quod omnes transeuntes propter eum subsisterent.
2SAM|20|13|Amoto igitur illo de via, transibat omnis vir sequens Ioab ad persequendum Seba filium Bochri.
2SAM|20|14|Porro ille transierat per omnes tribus Israel usque in Abelbethmaacha; omnesque Bochritae congregati sunt et ingressi sunt etiam post eum.
2SAM|20|15|Venerunt itaque et oppugnabant eum in Abelbethmaacha et fuderunt contra civitatem aggerem, qui stetit contra antemurale; et omnis populus, qui erat cum Ioab, moliebatur destruere muros.
2SAM|20|16|Et exclamavit mulier sapiens de civitate: " Audite, audite! Dicite Ioab: "Appropinqua huc, et loquar tecum" ".
2SAM|20|17|Qui cum accessisset ad eam, ait illi: " Tu es Ioab? ". Et ille respondit: " Ego ". Ad quem sic locuta est: " Audi sermones ancillae tuae. Qui respondit: " Audio ".
2SAM|20|18|Rursumque illa: " Sermo, inquit, dicebatur in vetere proverbio: Interrogent in Abel, et sic perficient rem".
2SAM|20|19|Ego pacifica fidelium Israel, et tu quaeris subruere civitatem et evertere matrem in Israel. Quare praecipitas hereditatem Domini? ".
2SAM|20|20|Respondensque Ioab ait: " Absit, absit hoc a me; non praecipito neque demolior.
2SAM|20|21|Non se sic habet res, sed homo de monte Ephraim, Seba filius Bochri cognomine, levavit manum suam contra regem David; tradite illum solum, et recedam a civitate". Et ait mulier ad Ioab: " Ecce, caput eius mittetur ad te per murum ".
2SAM|20|22|Ingressa est ergo ad omnem populum et locuta est eis sapienter. Qui abscissum caput Seba filii Bochri proiecerunt ad Ioab. Et ille cecinit tuba, et recesserunt ab urbe unusquisque in tabernacula sua. Ioab autem reversus est Ierusalem ad regem.
2SAM|20|23|Erat ergo Ioab super omnem exercitum Israel; Banaias autem filius Ioiadae super Cherethaeos et Phelethaeos;
2SAM|20|24|Adoniram vero super onera; porro Iosaphat filius Ahilud a commentariis.
2SAM|20|25|Siva autem scriba, Sadoc vero et Abiathar sacerdotes;
2SAM|20|26|Hira quoque Iairites erat sacerdos David.
2SAM|21|1|Facta est fames in diebus David tribus annis iugiter. Et consuluit David oraculum Domini, dixitque Dominus: " Super Saul et super domum eius est sanguis, quia occidit Gabaonitas ".
2SAM|21|2|Vocatis ergo Gabaonitis, rex dixit ad eos - porro Gabaonitae non sunt de filiis Israel, sed reliquiae Amorraeorum; filii quippe Israel iuraverant eis, sed voluit Saul percutere eos zelo suo pro filiis Israel et Iudae -;
2SAM|21|3|dixit ergo David ad Gabaonitas: " Quid faciam vobis? Et quod erit vestri piaculum, ut benedicatis hereditati Domini? ".
2SAM|21|4|Dixeruntque ei Gabaonitae: " Non est nobis super argento et auro quaestio contra Saul et contra domum eius; neque nobis licet interficere hominem de Israel ". Ad quos ait: " Quod ergo dixeritis, faciam vobis ".
2SAM|21|5|Qui dixerunt regi: " De filiis viri, qui attrivit nos et cogitavit delere nos ita ut ne unus quidem nostrum residuus esset in cunctis finibus Israel,
2SAM|21|6|dentur nobis septem viri, et suspendamus eos in patibulis Domino in Gabaon in monte Domini ". Et ait rex: " Ego dabo ".
2SAM|21|7|Pepercitque rex Meribbaal filio Ionathan filii Saul propter iusiurandum Domini, quod fuerat inter David et inter Ionathan filium Saul.
2SAM|21|8|Tulit itaque rex duos filios Respha filiae Aia, quos peperit Saul, Armoni et Meribbaal, et quinque filios Merob filiae Saul, quos genuerat Hadrieli filio Berzellai, qui fuit de Molathi,
2SAM|21|9|et dedit eos in manu Gabaonitarum, qui suspenderunt illos in monte coram Domino. Et ceciderunt hi septem simul, occisi in diebus messis primis, incipiente messione hordei.
2SAM|21|10|Tollens autem Respha filia Aia cilicium substravit sibi super petram ab initio messis, donec stillaret aqua super eos de caelo, et non dimisit aves caeli considere super eos per diem neque bestias campi per noctem.
2SAM|21|11|Et nuntiata sunt David, quae fecerat Respha filia Aia concubina Saul.
2SAM|21|12|Et abiit David et tulit ossa Saul et ossa Ionathan filii eius a civibus Iabes Galaad, qui furati fuerant ea de platea Bethsan, in qua suspenderant eos Philisthim, cum interfecissent Saul in Gelboe,
2SAM|21|13|et asportavit inde ossa Saul et ossa Ionathan filii eius; et colligentes ossa eorum, qui suspensi fuerant,
2SAM|21|14|sepelierunt ea cum ossibus Saul et Ionathan filii eius in terra Beniamin in Sela, in sepulcro Cis patris eius. Feceruntque omnia, quae praeceperat rex; et repropitiatus est Deus terrae post haec.
2SAM|21|15|Factum est autem rursum proelium Philisthinorum adversum Israel, et descendit David et servi eius cum eo, et pugnabant contra Philisthim, et fatigatus est David.
2SAM|21|16|Iesbibenob, qui fuit de genere Rapha - ferrum hastae trecentos siclos appendebat - et accinctus erat ense novo, nisus est percutere David;
2SAM|21|17|praesidioque ei fuit Abisai filius Sarviae et percussum Philisthaeum interfecit. Tunc iuraverunt viri David dicentes: " Iam non egredieris nobiscum in bellum, ne exstinguas lucernam Israel ".
2SAM|21|18|Fuitque rursum bellum in Gob contra Philisthaeos; tunc percussit Sobbochai de Husa Saph de stirpe Rapha.
2SAM|21|19|Et fuit iterum bellum in Gob contra Philisthaeos, in quo percussit Elchanan filius Iair Bethlehemites Goliath Getthaeum, cuius hastile hastae erat quasi liciatorium texentium.
2SAM|21|20|Et adhuc fuit bellum in Geth, in quo vir excelsus, qui senos in manibus pedibusque habebat digitos, id est viginti et quattuor, et is quoque erat de origine Rapha,
2SAM|21|21|exprobravit Israel; percussit autem eum Ionathan filius Samma fratris David.
2SAM|21|22|Hi quattuor erant de genere Rapha ex Geth et ceciderunt per manum David et servorum eius.
2SAM|22|1|Locutus est autem David Domino verba carminis huius in die, qua liberavit eum Dominus de manu omnium inimicorum suorum et de manu Saul,
2SAM|22|2|et ait: Dominus petra mea et arx mea et salvator meus;
2SAM|22|3|Deus meus, rupes mea, in quam confugiam,scutum meum et cornu salutis meae!Munimentum meum et refugium meum.Salvator meus, de violentia liberabis me.
2SAM|22|4|Laudabilem invocabo Dominumet ab inimicis meis salvus ero.
2SAM|22|5|Quia circumdederunt me fluctus mortis,torrentes Belial terruerunt me;
2SAM|22|6|praeoccupaverunt me laquei mortis.
2SAM|22|7|In tribulatione mea invocavi Dominumet ad Deum meum clamavi;et exaudivit de templo suo vocem meam,et clamor meus venit ad aures eius.
2SAM|22|8|Commota est et contremuit terra;fundamenta caelorum concussa suntet conquassata, quoniam iratus est.
2SAM|22|9|Ascendit fumus de naribus eius,et ignis de ore eius vorabat;carbones incensi sunt ab eo.
2SAM|22|10|Et inclinavit caelos et descendit,et caligo sub pedibus eius.
2SAM|22|11|Et ascendit super cherub et volavitet devolavit super pennas venti.
2SAM|22|12|Posuit tenebras in circuitu suo tabernaculum suum,tenebrosas aquas, nubes densissimas.
2SAM|22|13|Prae fulgore in conspectu eiusincensi sunt carbones ignis.
2SAM|22|14|Intonuit de caelo Dominus,et Excelsus dedit vocem suam.
2SAM|22|15|Misit sagittas et dissipavit eos,fulguravit fulmina et conturbavit eos.
2SAM|22|16|Et apparuerunt effusiones maris,et revelata sunt fundamenta orbisab increpatione Domini,ab inspiratione spiritus furoris eius.
2SAM|22|17|Misit de excelso et assumpsit me,traxit me de aquis multis;
2SAM|22|18|liberavit me ab inimico meo potentissimo,ab his, qui oderant me, qui robustiores me erant.
2SAM|22|19|Praevenerunt me in die afflictionis meae,et factus est Dominus firmamentum meum;
2SAM|22|20|et eduxit me in latitudinem,liberavit me, quia complacui ei.
2SAM|22|21|Retribuit mihi Dominus secundum iustitiam meamet secundum munditiam manuum mearum reddit mihi,
2SAM|22|22|quia custodivi vias Dominiet non egi impie a Deo meo.
2SAM|22|23|Omnia enim iudicia eius in conspectu meo,et a praeceptis eius non recessi;
2SAM|22|24|et fui immaculatus cum eoet custodivi me ab iniquitate mea.
2SAM|22|25|Et retribuet mihi Dominus secundum iustitiam meamet secundum munditiam meam in conspectu oculorum suorum.
2SAM|22|26|Cum sancto sanctus eriset cum viro innocente innocens eris;
2SAM|22|27|cum electo electus eriset cum perverso callidus eris.
2SAM|22|28|Et populum pauperem salvum facieset oculos superborum humiliabis,
2SAM|22|29|quia tu lucerna mea, Domine,et Deus meus illuminat tenebras meas.
2SAM|22|30|In te enim aggrediar hostium turmas,in Deo meo transiliam murum.
2SAM|22|31|Deus, immaculata via eius,eloquium Domini igne examinatum;scutum est omnium sperantium in se.
2SAM|22|32|Quoniam quis est Deus praeter Dominum?Et quae rupes praeter Deum nostrum?
2SAM|22|33|Deus, qui accinxit me fortitudineet complanavit perfectam viam meam,
2SAM|22|34|coaequans pedes meos cerviset super excelsa statuens me;
2SAM|22|35|docens manus meas ad proelium,et tendunt arcum aereum brachia mea.
2SAM|22|36|Dedisti mihi clipeum salutis tuae,et exauditio tua magnificavit me.
2SAM|22|37|Dilatasti gressus meos subtus me,et non sunt infirmati tali mei.
2SAM|22|38|Persequebar inimicos meos et conterebamet non convertebar, donec consumerem eos.
2SAM|22|39|Consumpsi eos et confregi, ut non consurgerent:ceciderunt sub pedibus meis.
2SAM|22|40|Accinxisti me fortitudine ad proelium,incurvasti insurgentes in me subtus me.
2SAM|22|41|Inimicos meos dedisti mihi dorsum,odientes me, et disperdidi eos.
2SAM|22|42|Clamaverunt, et non erat qui salvaret,ad Dominum, et non exaudivit eos.
2SAM|22|43|Contrivi eos ut pulverem terrae,quasi lutum platearum comminui eos.
2SAM|22|44|Salvasti me a contradictionibus populi mei,constituisti me in caput gentium.Populus, quem ignorabam, servit mihi,
2SAM|22|45|filii alieni blandiuntur mihi,auditu auris oboediunt mihi.
2SAM|22|46|Filii alieni defluuntet contremiscunt ex arcibus suis.
2SAM|22|47|Vivit Dominus, et benedicta petra mea,et exaltetur Deus, petra salutis meae.
2SAM|22|48|Deus, qui das vindictas mihiet deicis populos sub me.
2SAM|22|49|Qui educis me ab inimicis meiset ab insurgentibus in me elevas me;a viro iniquo liberas me.
2SAM|22|50|Propterea confitebor tibi, Domine, in gentibus,et nomini tuo cantabo:
2SAM|22|51|Magnificat salutes regis suiet facit misericordiam christo suo Davidet semini eius in sempiternum ".
2SAM|23|1|Haec autem sunt verba David novissima: Dixit David filius Isai,dixit vir constitutus in alto,christus Dei Iacob,suavis psalta Israel.
2SAM|23|2|Spiritus Domini locutus est per me, et sermo eius super linguam meam.
2SAM|23|3|Locutus est Deus Israel,mihi dixit Petra Israel:Dominator hominum iustus,dominator in timore Dei
2SAM|23|4|est sicut lux aurorae, oriente sole,mane absque nubibus;de splendore post pluviamherba oritur de terra".
2SAM|23|5|Nonne sic est domus mea cum Deo?Quia pactum aeternum statuit mihi,dispositum in omnibus atque munitum.Cunctam enim salutem meam et omne desiderabilenonne faciet germinare?
2SAM|23|6|Praevaricatores autemquasi spinae abiectae universi,quae non tolluntur manibus;
2SAM|23|7|et si quis tangere voluerit eas,armabitur ferro et ligno lanceato,igneque succensae comburentur ".
2SAM|23|8|Haec nomina fortium David:Iesbaal Hachamonites, princeps inter tres, ipse levavit hastam suam super octingentos, quos interfecit impetu uno.
2SAM|23|9|Post hunc Eleazar filius Dodo Ahohites, inter tres fortes. Qui erat cum David in Aphesdommim, quando Philisthim congregati sunt illuc in proelium.
2SAM|23|10|Cumque ascendissent viri Israel, ipse stetit et percussit Philisthaeos, donec deficeret manus eius et obrigesceret cum gladio; fecitque Dominus salutem magnam in die illa, et populus reversus est tantum ad spolia detrahenda.
2SAM|23|11|Et post hunc Samma filius Age Ararites. Et congregati sunt Philisthim in Lehi; erat quippe ibi ager lente plenus. Cumque fugisset populus a facie Philisthim,
2SAM|23|12|stetit ille in medio agri et tuitus est eum percussitque Philisthaeos, et fecit Dominus salutem magnam.
2SAM|23|13|Et descenderunt tres de triginta et venerunt tempore messis ad David in speluncam Odollam; castra autem Philisthinorum erant posita in valle Raphaim.
2SAM|23|14|Et David erat tunc in praesidio; porro statio Philisthinorum tunc erat in Bethlehem.
2SAM|23|15|Desideravit igitur David et ait: " O si quis mihi daret potum aquae de cisterna, quae est in Bethlehem iuxta portam! ".
2SAM|23|16|Irruperunt ergo tres fortes castra Philisthinorum et hauserunt aquam de cisterna Bethlehem, quae erat iuxta portam, et attulerunt ad David. At ille noluit bibere, sed libavit illam Domino
2SAM|23|17|dicens: " Propitius mihi sit Dominus, ne faciam hoc. Num sanguinem hominum istorum, qui profecti sunt in animarum periculo, bibam? ". Noluit ergo bibere. Haec fecerunt tres robustissimi.
2SAM|23|18|Abisai autem frater Ioab filius Sarviae princeps erat de triginta. Ipse est qui elevavit hastam suam contra trecentos, quos interfecit. Nominatus in triginta
2SAM|23|19|et inter triginta nobilior eratque eorum princeps; sed usque ad tres primos non pervenerat.
2SAM|23|20|Et Banaias filius Ioiadae vir fortissimus magnorum operum de Cabseel. Ipse percussit duos filios Ariel de Moab, et ipse descendit et percussit leonem in media cisterna in diebus nivis.
2SAM|23|21|Ipse quoque interfecit virum Aegyptium, virum procerae staturae habentem in manu hastam; itaque cum descendisset ad eum cum baculo, vi extorsit hastam de manu Aegyptii et interfecit eum hasta sua.
2SAM|23|22|Haec fecit Banaias filius Ioiadae, et ipse nominatus inter triginta fortissimos.
2SAM|23|23|Erat autem nobilior inter triginta; verumtamen usque ad tres non pervenerat. Fecitque eum David sibi caput satellitum suorum.
2SAM|23|24|Asael frater Ioab erat inter triginta. Elchanan filius Dodo de Bethlehem,
2SAM|23|25|Samma de Harod, Elica de Harod,
2SAM|23|26|Heles de Phalti, Hira filius Acces de Thecua,
2SAM|23|27|Abiezer de Anathoth, Sobbochai de Husa,
2SAM|23|28|Selmon Ahohites, Maharai Netophathites,
2SAM|23|29|Heled filius Baana Netophathites, Ithai filius Ribai de Gabaa filiorum Beniamin,
2SAM|23|30|Banaia Pharathonites, Heddai de torrentibus Gaas,
2SAM|23|31|Abibaal Arbathites, Azmaveth de Bahurim,
2SAM|23|32|Eliaba de Saalbon, Iasen de Gun,
2SAM|23|33|Ionathan filius Samma de Arar, Ahiam filius Sarar Ararites.
2SAM|23|34|Eliphalet filius Aasbai Maachathitae, Eliam filius Achitophel Gilonites,
2SAM|23|35|Hesro de Carmel, Pharai de Arab,
2SAM|23|36|Igal filius Nathan de Soba, Bani de Gad,
2SAM|23|37|Selec de Ammon, Naharai Berothites armiger Ioab filii Sarviae,
2SAM|23|38|Hira Iethrites, Gareb et ipse Iethrites,
2SAM|23|39|Urias Hetthaeus.Omnes triginta septem.
2SAM|24|1|Et addidit furor Domini ira sci contra Israel; commovit que David contra eos dicens: " Vade, numera Israel et Iudam ".
2SAM|24|2|Dixitque rex ad Ioab et ad principes exercitus sui, qui erant cum eo: " Perambula omnes tribus Israel a Dan usque Bersabee, et numerate populum, ut sciam numerum eius ".
2SAM|24|3|Dixitque Ioab regi: " Adaugeat Dominus Deus tuus ad populum, quantus nunc est, centuplum in conspectu domini mei regis! Sed quid sibi dominus meus rex vult in re huiuscemodi? ".
2SAM|24|4|Praevaluit autem sermo regis contra Ioab et principes exercitus; egressusque est Ioab et principes militum a facie regis, ut numerarent populum Israel.
2SAM|24|5|Cumque pertransissent Iordanem, inceperunt ab Aroer et ab urbe, quae est in media valle, transeuntes ad Gaditas et ad Iazer.
2SAM|24|6|Et pervenerunt in Galaad et in terram Hetthaeorum in Cades et venerunt in Dan. Et a Dan converterunt se ad Sidonem
2SAM|24|7|et pervenerunt ad arcem Tyri et omnes urbes Hevaei et Chananaei exieruntque ad Nageb Iudae in Bersabee.
2SAM|24|8|Et, lustrata universa terra, affuerunt post novem menses et viginti dies in Ierusalem.
2SAM|24|9|Dedit ergo Ioab numerum descriptionis populi regi; et inventa sunt de Israel octingenta milia virorum fortium, qui educerent gladium, et de Iuda quingenta milia pugnatorum.
2SAM|24|10|Percussit autem cor David eum, postquam numeratus est populus, et dixit David ad Dominum: " Peccavi valde in hoc facto; nunc vero precor, Domine, ut transferas iniquitatem servi tui, quia stulte egi nimis ".
2SAM|24|11|Surrexit itaque David mane, et sermo Domini factus est ad Gad propheten, videntem David, dicens:
2SAM|24|12|" Vade et loquere ad David: Haec dicit Dominus: Trium tibi datur optio; elige unum, quod volueris ex his, ut faciam tibi ".
2SAM|24|13|Cumque venisset Gad ad David, nuntiavit ei dicens: " Aut tribus annis veniet tibi fames in terra tua, aut tribus mensibus fugies adversarios tuos, et illi te persequentur, aut certe tribus diebus erit pestilentia in terra tua. Nunc ergo delibera et vide quem respondeam ei, qui me misit, sermonem ".
2SAM|24|14|Dixit autem David ad Gad: " Artor nimis; sed melius est, ut incidamus in manu Domini - multae enim misericordiae eius sunt - quam in manu hominum! ".
2SAM|24|15|Et elegit sibi David pestilentiam; et erant dies messis tritici. Immisitque Dominus pestilentiam in Israel de mane usque ad tempus constitutum, et mortui sunt ex populo a Dan usque Bersabee septuaginta milia virorum.
2SAM|24|16|Cumque extendisset manum suam angelus super Ierusalem, ut disperderet eam, misertus est Dominus super afflictione et ait angelo percutienti populum: " Sufficit; nunc contine manum tuam! ".Erat autem angelus Domini iuxta aream Areuna Iebusaei.
2SAM|24|17|Dixitque David ad Dominum, cum vidisset angelum caedentem populum: " Ego sum qui peccavi, ego inique egi; isti, qui oves sunt, quid fecerunt? Vertatur, obsecro, manus tua contra me et contra domum patris mei ".
2SAM|24|18|Venit autem Gad ad David in die illa et dixit ei: " Ascende, constitue Domino altare in area Areuna Iebusaei ".
2SAM|24|19|Et ascendit David iuxta sermonem Gad, quem praeceperat ei Dominus.
2SAM|24|20|Conspiciensque Areuna animadvertit regem et servos eius transire ad se
2SAM|24|21|et egressus adoravit regem prono vultu in terra et ait: " Quid causae est, ut veniat dominus meus rex ad servum suum? ". Cui David ait: " Ut emam a te aream et aedificem altare Domino, et cesset interfectio, quae grassatur in populo ".
2SAM|24|22|Et ait Areuna ad David: " Accipiat et offerat dominus meus rex, sicut ei placet. Ecce boves in holocaustum et plaustrum et iuga boum in usum lignorum.
2SAM|24|23|Omnia dat Areuna, o rex, regi ". Dixitque Areuna ad regem: " Dominus Deus tuus suscipiat votum tuum! ".
2SAM|24|24|Cui respondens rex ait: " Nequaquam; sed emam pretio a te et non offeram Domino Deo meo holocausta gratuita ". Emit ergo David aream et boves argenti siclis quinquaginta.
2SAM|24|25|Et aedificavit ibi David altare Domino et obtulit holocausta et pacifica.Et repropitiatus est Dominus terrae, et cohibita est plaga ab Israel.
1KGS|1|1|Et rex David senuerat habebat que aetatis plurimos dies; cum que operiretur vestibus, non calefiebat.
1KGS|1|2|Dixerunt ergo ei servi sui: " Quaeratur domino nostro regi adulescentula virgo et stet coram rege et curam eius agat dormiatque in sinu tuo et calefaciat dominum nostrum regem ".
1KGS|1|3|Quaesierunt igitur adulescentulam speciosam in omnibus finibus Israel et invenerunt Abisag Sunamitin et adduxerunt eam ad regem.
1KGS|1|4|Erat autem puella pulchra nimis et curam agebat regis et ministrabat ei; rex vero non cognovit eam.
1KGS|1|5|Adonias autem filius Haggith elevabatur dicens: " Ego regnabo! ". Fecitque sibi currum et equites et quinquaginta viros, qui ante eum currerent.
1KGS|1|6|Nec corripuit eum pater suus aliquando dicens: " Quare hoc fecisti? ". Erat autem et ipse pulcher valde, secundus natu post Absalom.
1KGS|1|7|Et sermo ei cum Ioab filio Sarviae et cum Abiathar sacerdote, qui adiuvabant partes Adoniae.
1KGS|1|8|Sadoc vero sacerdos et Banaias filius Ioiadae et Nathan propheta et Semei et Rei et robur exercitus David non erat cum Adonia.
1KGS|1|9|Immolatis ergo Adonias ovibus et vitulis et pinguibus iuxta lapidem Zoheleth, qui erat vicinus fonti Rogel, vocavit universos fratres suos filios regis et omnes viros Iudae servos regis;
1KGS|1|10|Nathan autem prophetam et Banaiam et robustos quosque et Salomonem fratrem suum non vocavit.
1KGS|1|11|Dixit itaque Nathan ad Bethsabee matrem Salomonis: " Num audisti quod regnaverit Adonias filius Haggith, et dominus noster David hoc ignorat?
1KGS|1|12|Nunc ergo veni, accipe a me consilium et salva animam tuam filiique tui Salomonis.
1KGS|1|13|Vade et ingredere ad regem David et dic ei: Nonne tu, domine mi rex, iurasti mihi ancillae tuae dicens: "Salomon filius tuus regnabit post me et ipse sedebit in solio meo"? Quare ergo regnat Adonias?
1KGS|1|14|Et, adhuc ibi te loquente cum rege, ego veniam post te et complebo sermones tuos ".
1KGS|1|15|Ingressa est itaque Bethsabee ad regem in cubiculo; rex autem senuerat nimis, et Abisag Sunamitis ministrabat ei.
1KGS|1|16|Inclinavit se Bethsabee et adoravit regem; ad quam rex: " Quid tibi, inquit, vis? ".
1KGS|1|17|Quae respondens ait: " Domine mi, tu iurasti per Dominum Deum tuum ancillae tuae: "Salomon filius tuus regnabit post me, et ipse sedebit in solio meo";
1KGS|1|18|et ecce nunc Adonias regnat, te, domine mi rex, ignorante.
1KGS|1|19|Mactavit boves et pinguia quaeque et oves plurimas et vocavit omnes filios regis, Abiathar quoque sacerdotem et Ioab principem militiae; Salomonem autem servum tuum non vocavit.
1KGS|1|20|Verumtamen, domine mi rex, in te oculi respiciunt totius Israel, ut indices eis quis sedere debeat in solio tuo, domine mi rex, post te.
1KGS|1|21|Eritque, cum dormierit dominus meus rex cum patribus suis, erimus ego et filius meus Salomon peccatores ".
1KGS|1|22|Adhuc illa loquente cum rege, Nathan propheta venit;
1KGS|1|23|et nuntiaverunt regi dicentes: " Adest Nathan propheta ". Cumque introisset ante conspectum regis et adorasset eum pronus in terram,
1KGS|1|24|dixit Nathan: " Domine mi rex, tu ergo dixisti: "Adonias regnet post me, et ipse sedeat super thronum meum"?
1KGS|1|25|Quia descendit hodie et immolavit boves et pinguia et arietes plurimos et vocavit universos filios regis et principes exercitus, Abiathar quoque sacerdotem; illique vescentes et bibentes coram eo dixerunt: "Vivat rex Adonias!".
1KGS|1|26|Me autem servum tuum et Sadoc sacerdotem et Banaiam filium Ioiadae et Salomonem famulum tuum non vocavit.
1KGS|1|27|Numquid a domino meo rege exivit hoc verbum, et mihi non indicasti servo tuo quis sessurus esset super thronum domini mei regis post eum? ".
1KGS|1|28|Et respondit rex David dicens: " Vocate ad me Bethsabee ". Quae cum fuisset ingressa coram rege et stetisset ante eum,
1KGS|1|29|iuravit rex et ait: " Vivit Dominus, qui eruit animam meam de omni angustia,
1KGS|1|30|quia, sicut iuravi tibi per Dominum, Deum Israel, dicens: Salomon filius tuus regnabit post me et ipse sedebit super solium meum pro me, sic faciam hodie ".
1KGS|1|31|Summissoque Bethsabee in terram vultu, adoravit regem dicens: " Vivat dominus meus rex David in aeternum! ".
1KGS|1|32|Dixit quoque rex David: " Vocate mihi Sadoc sacerdotem et Nathan prophetam et Banaiam filium Ioiadae ". Qui cum ingressi fuissent coram rege,
1KGS|1|33|dixit ad eos: " Tollite vobiscum servos domini vestri et imponite Salomonem filium meum, super mulam meam et ducite eum in Gihon,
1KGS|1|34|et ungat eum ibi Sadoc sacerdos et Nathan propheta in regem super Israel, et canetis bucina atque dicetis: "Vivat rex Salomon!".
1KGS|1|35|Et ascendetis post eum, et veniet et sedebit super solium meum, et ipse regnabit pro me; illique praecipiam, ut sit dux super Israel et super Iudam ".
1KGS|1|36|Et respondit Banaias filius Ioiadae regi dicens: " Amen, sic loquatur Dominus Deus domini mei regis.
1KGS|1|37|Quomodo fuit Dominus cum domino meo rege, sic sit cum Salomone et sublimius faciat solium eius a solio domini mei regis David ".
1KGS|1|38|Descendit ergo Sadoc sacerdos et Nathan propheta et Banaias filius Ioiadae et Cherethi et Phelethi, et imposuerunt Salomonem super mulam regis David et adduxerunt eum in Gihon.
1KGS|1|39|Sumpsitque Sadoc sacerdos cornu olei de tabernaculo et unxit Salomonem; et cecinerunt bucina, et dixit omnis populus: " Vivat rex Salomon! ".
1KGS|1|40|Et ascendit universa multitudo post eum, et populus canebat tibiis et laetabatur gaudio magno, et insonuit terra ad clamorem eorum.
1KGS|1|41|Audivit autem Adonias et omnes, qui invitati fuerant ab eo; iamque convivium finitum erat. Sed et Ioab, audita voce tubae, ait: " Quid sibi vult clamor civitatis tumultuantis? ".
1KGS|1|42|Adhuc illo loquente, Ionathan filius Abiathar sacerdotis venit; cui dixit Adonias: " Ingredere, quia vir strenuus es et bona nuntians ".
1KGS|1|43|Responditque Ionathan Adoniae: " Nequaquam! Dominus enim noster, rex David, regem constituit Salomonem
1KGS|1|44|misitque cum eo Sadoc sacerdotem et Nathan prophetam et Banaiam filium Ioiadae et Cherethi et Phelethi, et imposuerunt eum super mulam regis;
1KGS|1|45|unxeruntque eum Sadoc sacerdos et Nathan propheta regem in Gihon. Et ascenderunt inde laetantes, et insonuit civitas; haec est vox, quam audistis.
1KGS|1|46|Sed et Salomon sedit super solio regni,
1KGS|1|47|et ingressi servi regis benedixerunt domino nostro regi David dicentes: Amplificet Deus nomen Salomonis super nomen tuum et magnificet thronum eius super thronum tuum". Et adoravit rex in lectulo suo.
1KGS|1|48|Insuper et haec locutus est: "Benedictus Dominus, Deus Israel, qui dedit hodie sedentem in solio meo, videntibus oculis meis" ".
1KGS|1|49|Territi sunt ergo et surrexerunt omnes, qui invitati fuerant ab Adonia, et ivit unusquisque in viam suam.
1KGS|1|50|Adonias autem timens Salomonem surrexit et abiit tenuitque cornua altaris.
1KGS|1|51|Et nuntiaverunt Salomoni dicentes: " Ecce Adonias timens regem Salomonem tenuit cornua altaris dicens: "Iuret mihi hodie rex Salomon quod non interficiat servum suum gladio"".
1KGS|1|52|Dixitque Salomon: " Si fuerit vir bonus, non cadet ne unus quidem capillus eius in terram; sin autem malum inventum fuerit in eo, morietur.
1KGS|1|53|Misit ergo rex Salomon et eduxit eum ab altari, et ingressus adoravit regem Salomonem; dixitque ei Salomon: " Vade in domum tuam ".
1KGS|2|1|Appropinquaverant autem dies David ut moreretur, praecepit que Salomoni filio suo dicens:
1KGS|2|2|" Ego ingredior viam universae terrae; confortare et esto vir
1KGS|2|3|et observa decreta Domini Dei tui, ut ambules in viis eius et custodias statuta eius et praecepta eius et iudicia et testimonia, sicut scriptum est in lege Moysi, ut prospere agas in universis, quae facis et quocumque te verteris;
1KGS|2|4|ut confirmet Dominus sermonem suum, quem locutus est de me dicens: "Si custodierint filii tui viam suam et ambulaverint coram me in veritate, in omni corde suo et in omni anima sua, non auferetur tibi vir de solio Israel".
1KGS|2|5|Tu quoque nosti, quae fecerit mihi Ioab filius Sarviae, quae fecerit duobus principibus exercitus Israel, Abner filio Ner et Amasae filio Iether, quos occidit; et effudit sanguinem belli in pace et posuit cruorem proelii in balteo suo, qui erat circa lumbos eius, et in calceamento suo, quod erat in pedibus eius.
1KGS|2|6|Facies ergo iuxta sapientiam tuam et non deduces canitiem eius pacifice ad inferos.
1KGS|2|7|Sed filiis Berzellai Galaaditis reddes gratiam, eruntque comedentes in mensa tua; occurrerunt enim mihi, quando fugiebam a facie Absalom fratris tui.
1KGS|2|8|Habes quoque apud te Semei filium Gera de Beniamin de Bahurim, qui maledixit mihi maledictione pessima, quando ibam ad Mahanaim; sed quia descendit mihi in occursum ad Iordanem, et iuravi ei per Dominum dicens: Non te interficiam gladio.
1KGS|2|9|Tu noli pati esse eum innoxium; vir autem sapiens es et scies, quae facias ei deducesque canos eius cum sanguine ad infernum ".
1KGS|2|10|Dormivit igitur David cum patribus suis et sepultus est in civitate David.
1KGS|2|11|Dies autem, quibus regnavit David super Israel, quadraginta anni sunt: in Hebron regnavit septem annis, in Ierusalem triginta tribus.
1KGS|2|12|Salomon autem sedit super thronum David patris sui, et firmatum est regnum eius nimis.
1KGS|2|13|Et ingressus est Adonias filius Haggith ad Bethsabee matrem Salomonis, quae dixit ei: " Pacificusne ingressus tuus? ". Qui respondit: " Pacificus.
1KGS|2|14|Addiditque: " Sermo mihi est ad te ". Cui ait: " Loquere ". Et ille:
1KGS|2|15|" Tu, inquit, nosti quia meum erat regnum, et me proposuerat omnis Israel sibi in regem, sed translatum est regnum et factum est fratris mei; a Domino enim constitutum est ei.
1KGS|2|16|Nunc ergo petitionem unam deprecor a te; ne confundas faciem meam ". Quae dixit ad eum: " Loquere ".
1KGS|2|17|Et ille ait: " Precor, ut dicas Salomoni regi - neque enim negare tibi quidquam potest - ut det mihi Abisag Sunamitin uxorem ".
1KGS|2|18|Et ait Bethsabee: " Bene, ego loquar pro te regi ".
1KGS|2|19|Venit ergo Bethsabee ad regem Salomonem, ut loqueretur ei pro Adonia. Et surrexit rex in occursum eius adoravitque eam et sedit super thronum suum; positus quoque est thronus matri regis, quae sedit ad dexteram eius.
1KGS|2|20|Dixitque ei: " Petitionem unam parvulam ego deprecor a te; ne confundas faciem meam". Dixit ei rex: " Pete, mater mi, neque enim fas est, ut avertam faciem tuam ".
1KGS|2|21|Quae ait: " Detur Abisag Sunamitis Adoniae fratri tuo uxor ".
1KGS|2|22|Responditque rex Salomon et dixit matri suae: " Quare postulas Abisag Sunamitin Adoniae? Postula ei et regnum! Ipse est enim frater meus maior me et habet Abiathar sacerdotem et Ioab filium Sarviae ".
1KGS|2|23|Iuravit itaque rex Salomon per Dominum dicens: " Haec faciat mihi Deus et haec addat, certe contra animam suam locutus est Adonias verbum hoc.
1KGS|2|24|Et nunc, vivit Dominus, qui firmavit me et collocavit me super solium David patris mei et qui fecit mihi domum, sicut locutus est, certe hodie occidetur Adonias ".
1KGS|2|25|Misitque rex Salomon per manum Banaiae filii Ioiadae, qui interfecit eum, et mortuus est.
1KGS|2|26|Abiathar quoque sacerdoti dixit rex: " Vade in Anathoth ad agrum tuum; es quidem vir mortis, sed hodie te non interficiam, quia portasti arcam Domini Dei coram David patre meo et sustinuisti laborem in omnibus, in quibus laboravit pater meus ".
1KGS|2|27|Eiecit ergo Salomon Abiathar, ut non esset sacerdos Domini, ut impleretur sermo Domini, quem locutus est super domum Heli in Silo.
1KGS|2|28|Venit autem nuntius ad Ioab. Ioab autem declinaverat post Adoniam, cum post Absalom non declinasset; fugit ergo Ioab in tabernaculum Domini et apprehendit cornua altaris.
1KGS|2|29|Nuntiatumque est regi Salomoni, quod fugisset Ioab in tabernaculum Domini et esset iuxta altare; misitque Salomon Banaiam filium Ioiadae dicens: " Vade, interfice eum! ".
1KGS|2|30|Venit Banaias ad tabernaculum Domini et dixit ei: " Haec dicit rex: Egredere!". Qui ait: " Non egrediar, sed hic moriar ". Renuntiavit Banaias regi sermonem dicens: " Haec locutus est Ioab et haec respondit mihi ".
1KGS|2|31|Dixitque ei rex: " Fac, sicut locutus est, et interfice eum et sepeli; et amovebis sanguinem innocentem, qui effusus est a Ioab, a me et a domo patris mei.
1KGS|2|32|Et reddet Dominus sanguinem eius super caput eius, quia interfecit duos viros iustos melioresque se et occidit eos gladio, patre meo David ignorante: Abner filium Ner principem militiae Israel et Amasam filium Iether principem exercitus Iudae.
1KGS|2|33|Et revertetur sanguis illorum in caput Ioab et in caput seminis eius in sempiternum; David autem et semini eius et domui et throno illius sit pax usque in aeternum a Domino ".
1KGS|2|34|Ascendit itaque Banaias filius Ioiadae et aggressus eum interfecit; sepultusque est in domo sua in deserto.
1KGS|2|35|Et constituit rex Banaiam filium Ioiadae pro eo super exercitum et Sadoc sacerdotem posuit pro Abiathar.
1KGS|2|36|Misit quoque rex et vocavit Semei dixitque ei: " Aedifica tibi domum in Ierusalem et habita ibi et non egredieris inde huc atque illuc;
1KGS|2|37|quacumque autem die egressus fueris et transieris torrentem Cedron, scito te interficiendum; sanguis tuus erit super caput tuum ".
1KGS|2|38|Dixitque Semei regi: " Bonus sermo; sicut locutus est dominus meus rex, sic faciet servus tuus ". Habitavit itaque Semei in Ierusalem diebus multis.
1KGS|2|39|Factum est autem post annos tres, ut fugerent duo servi Semei ad Achis filium Maacha regem Geth; nuntiatumque est Semei quod servi eius essent in Geth.
1KGS|2|40|Et surrexit Semei et stravit asinum suum ivitque in Geth ad Achis ad requirendos servos suos et adduxit eos de Geth.
1KGS|2|41|Nuntiatum est autem Salomoni quod isset Semei in Geth de Ierusalem et redisset.
1KGS|2|42|Et mittens vocavit eum dixitque illi: " Nonne testificatus sum tibi per Dominum et praedixi tibi: Quacumque die egressus ieris huc et illuc, scito te esse moriturum? Et respondisti mihi "Bonus sermo; audivi".
1KGS|2|43|Quare ergo non custodisti iusiurandum Domini et praeceptum, quod praeceperam tibi? ".
1KGS|2|44|Dixitque rex ad Semei: " Tu nosti omne malum, cuius tibi conscium est cor tuum, quod fecisti David patri meo; reddit Dominus malitiam tuam in caput tuum.
1KGS|2|45|Et rex Salomon benedictus, et thronus David erit stabilis coram Domino usque in sempiternum ".
1KGS|2|46|Iussit itaque rex Banaiae filio Ioiadae, qui egressus percussit eum, et mortuus est. Confirmatum est igitur regnum in manu Salomonis.
1KGS|3|1|Et affinitate coniunctus est pharaoni regi Aegypti. Accepit namque filiam eius et adduxit in civitatem David, donec compleret aedificans domum suam et domum Domini et murum Ierusalem per circuitum.
1KGS|3|2|Attamen populus immolabat in excelsis; non enim aedificatum erat templum nomini Domini usque in diem illum.
1KGS|3|3|Dilexit autem Salomon Dominum ambulans in praeceptis David patris sui, excepto quod in excelsis immolabat et accendebat thymiama.
1KGS|3|4|Abiit itaque in Gabaon, ut immolaret ibi; illud quippe erat excelsum maximum. Mille hostias in holocaustum obtulit Salomon super altare illud.
1KGS|3|5|In Gabaon apparuit Dominus Salomoni per somnium nocte dicens: " Postula quod vis, ut dem tibi ".
1KGS|3|6|Et ait Salomon: " Tu fecisti cum servo tuo David patre meo misericordiam magnam, sicut ambulavit in conspectu tuo in veritate et iustitia et recto corde tecum; custodisti ei misericordiam tuam grandem et dedisti ei filium sedentem super thronum eius, sicut est hodie.
1KGS|3|7|Et nunc, Domine Deus meus, tu regnare fecisti servum tuum pro David patre meo. Ego autem sum puer parvus et ignorans egressum et introitum meum;
1KGS|3|8|et servus tuus in medio est populi, quem elegisti, populi infiniti, qui numerari et supputari non potest prae multitudine.
1KGS|3|9|Da ergo servo tuo cor docile, ut iudicare possit populum tuum et discernere inter bonum et malum. Quis enim potest iudicare populum tuum hunc multum? ".
1KGS|3|10|Placuit ergo sermo coram Domino quod Salomon rem huiuscemodi postulasset,
1KGS|3|11|et dixit Deus Salomoni: " Quia postulasti verbum hoc et non petisti tibi dies multos nec divitias aut animam inimicorum tuorum, sed postulasti tibi sapientiam ad discernendum iudicium,
1KGS|3|12|ecce feci tibi secundum sermones tuos et dedi tibi cor sapiens et intellegens, in tantum ut nullus ante te similis tui fuerit nec post te surrecturus sit;
1KGS|3|13|sed et haec, quae non postulasti, dedi tibi, divitias scilicet et gloriam, ut nemo fuerit similis tui in regibus cunctis diebus tuis.
1KGS|3|14|Si autem ambulaveris in viis meis et custodieris praecepta mea et mandata mea, sicut ambulavit David pater tuus, longos faciam dies tuos ".
1KGS|3|15|Igitur evigilavit Salomon et intellexit quod esset somnium. Cumque venisset Ierusalem, stetit coram arca foederis Domini et obtulit holocausta et fecit victimas pacificas et convivium universis famulis suis.
1KGS|3|16|Tunc venerunt duae mulieres meretrices ad regem steteruntque coram eo.
1KGS|3|17|Quarum una ait: " Obsecro, mi domine; ego et mulier haec habitabamus in domo una, et peperi apud eam in domo;
1KGS|3|18|tertia vero die, postquam ego peperi, peperit et haec; et eramus simul, nullusque alius nobiscum in domo, exceptis nobis duabus.
1KGS|3|19|Mortuus est autem filius mulieris huius nocte; dormiens quippe oppressit eum.
1KGS|3|20|Et consurgens intempesta nocte, silentio tulit filium meum de latere meo ancillae tuae dormientis et collocavit in sinu suo; suum autem filium, qui erat mortuus, posuit in sinu meo.
1KGS|3|21|Cumque surrexissem mane, ut darem lac filio meo, apparuit mortuus; quem diligentius intuens clara luce, deprehendi non esse meum, quem genueram ".
1KGS|3|22|Responditque altera mulier: " Non est ita, sed filius meus vivit, tuus autem mortuus est ". E contrario illa dicebat: " Mentiris. Filius quippe tuus mortuus est, meus autem vivit ". Atque in hunc modum contendebant coram rege.
1KGS|3|23|Tunc rex ait: " Haec dicit: "Filius meus vivit, et filius tuus mortuus est"; et ista respondit: "Non, sed filius tuus mortuus est, et filius meus vivit" ".
1KGS|3|24|Dixit ergo rex: " Afferte mihi gladium! ". Cumque attulissent gladium coram rege:
1KGS|3|25|" Dividite, inquit, infantem vivum in duas partes, et date dimidiam partem uni et dimidiam partem alteri ".
1KGS|3|26|Dixit autem mulier, cuius filius erat vivus, ad regem - commota sunt quippe viscera eius super filio suo -: " Obsecro, domine, date illi infantem vivum et nolite interficere eum ". E contrario illa dicebat: " Nec mihi nec tibi sit; dividatur ".
1KGS|3|27|Respondens rex ait: " Date huic infantem vivum, et non occidatur; haec est mater eius ".
1KGS|3|28|Audivit itaque omnis Israel iudicium, quod iudicasset rex; et timuerunt regem videntes sapientiam Dei esse in eo ad faciendum iudicium.
1KGS|4|1|Erat autem rex Salomon regnans super omnem Israel.
1KGS|4|2|Et hi principes quos habebat: Azarias filius Sadoc sacerdos;
1KGS|4|3|Elihoreph et Ahia filii Sisa scribae; Iosaphat filius Ahilud cancellarius;
1KGS|4|4|Banaias filius Ioiadae super exercitum; Sadoc autem et Abiathar sacerdotes;
1KGS|4|5|Azarias filius Nathan super praefectos; Zabud filius Nathan sacerdos amicus regis;
1KGS|4|6|et Ahisar praepositus domus et Adoniram filius Abda super tributa.
1KGS|4|7|Habebat autem Salomon duodecim praefectos super omnem Israel, qui praebebant annonam regi et domui eius; per singulos enim menses in anno singuli necessaria ministrabant.
1KGS|4|8|Et haec nomina eorum: Benhur in monte Ephraim;
1KGS|4|9|Bendecar in Maces et in Salebim et in Bethsames et in Elon et in Bethanan;
1KGS|4|10|Benhesed in Aruboth, ipsius erat Socho et omnis terra Epher;
1KGS|4|11|Benabinadab, cuius omnis regio Dor, Tapheth filiam Salomonis habebat uxorem;
1KGS|4|12|Baana filius Ahilud regebat Thanach et Mageddo et universam Bethsan, quae est iuxta Sarthan subter Iezrahel, a Bethsan usque Abelmehula et usque ultra Iecmaam;
1KGS|4|13|Bengaber in Ramoth Galaad habebat villas Iair filii Manasse in Galaad: ipse praeerat in omni regione Argob, quae est in Basan, sexaginta civitatibus magnis atque muratis, quae habebant seras aereas;
1KGS|4|14|Ahinadab filius Addo praeerat in Mahanaim;
1KGS|4|15|Achimaas in Nephthali, sed et ipse habebat Basemath filiam Salomonis in coniugio;
1KGS|4|16|Baana filius Chusai in Aser et in Baloth;
1KGS|4|17|Iosaphat filius Pharue in Issachar;
1KGS|4|18|Semei filius Ela in Beniamin;
1KGS|4|19|Gaber filius Uri in terra Galaad, in terra Sehon regis Amorraei et Og regis Basan, ut praefectus unus, qui erat in terra.
1KGS|4|20|Iuda et Israel innumerabiles, sicut arena maris in multitudine, comedentes et bibentes atque laetantes.
1KGS|5|1|Salomon autem erat in dicione sua habens omnia regna a Flu mine usque ad terram Philisthim et ad terminum Aegypti offerentium sibi munera et servientium ei cunctis diebus vitae eius.
1KGS|5|2|Erat autem cibus Salomonis per dies singulos triginta chori similae et sexaginta chori farinae,
1KGS|5|3|decem boves pingues et viginti boves pascuales et centum oves, excepta venatione cervorum, caprearum atque bubalorum et avium altilium.
1KGS|5|4|Ipse enim obtinebat omnem regionem, quae erat trans Flumen, a Thaphsa usque Gazam, et cunctos reges illarum regionum; et habebat pacem ex omni parte in circuitu.
1KGS|5|5|Habitabatque Iuda et Israel absque timore ullo, unusquisque sub vite sua et sub ficu sua a Dan usque Bersabee cunctis diebus Salomonis.
1KGS|5|6|Et habebat Salomon quattuor milia praesepia equorum currulium et duodecim milia equestres.
1KGS|5|7|Et praebebant supradicti praefecti necessaria mensae regis Salomonis et convivarum eius cum ingenti cura, unusquisque in suo mense.
1KGS|5|8|Hordeum quoque et paleas equorum et iumentorum deferebant in locum, ubi erat unicuique constitutum.
1KGS|5|9|Dedit quoque Deus sapientiam Salomoni et prudentiam multam nimis et latitudinem cordis quasi arenam, quae est in litore maris.
1KGS|5|10|Et praecedebat sapientia Salomonis sapientiam omnium Orientalium et Aegyptiorum;
1KGS|5|11|et erat sapientior cunctis hominibus, sapientior Ethan Ezrahita et Heman et Chalchol et Darda filiis Mahol et erat nominatus in universis gentibus per circuitum.
1KGS|5|12|Locutus est quoque Salomon tria milia parabolas, et fuerunt carmina eius quinque et mille.
1KGS|5|13|Et disputavit super lignis, a cedro, quae est in Libano, usque ad hyssopum, quae egreditur de pariete; et disseruit de iumentis et volucribus et reptilibus et piscibus.
1KGS|5|14|Et veniebant de cunctis populis ad audiendam sapientiam Salomonis, ab universis regibus terrae, qui audiebant sapientiam eius.
1KGS|5|15|Misit quoque Hiram rex Tyri servos suos ad Salomonem; audivit enim quod ipsum unxissent regem pro patre eius, quia amicus fuerat Hiram David omni tempore.
1KGS|5|16|Misit autem et Salomon ad Hiram dicens:
1KGS|5|17|" Tu scis voluntatem David patris mei et quia non potuerit aedificare domum nomini Domini Dei sui propter bella imminentia per circuitum, donec daret Dominus eos sub vestigio pedum eius.
1KGS|5|18|Nunc autem requiem dedit Dominus Deus meus mihi per circuitum; non est adversarius neque occursus malus.
1KGS|5|19|Quam ob rem cogito aedificare templum nomini Domini Dei mei, sicut locutus est Dominus David patri meo dicens: "Filius tuus, quem dabo pro te super solium tuum, ipse aedificabit domum nomini meo".
1KGS|5|20|Praecipe igitur, ut praecidant mihi cedros de Libano, et servi mei sint cum servis tuis; mercedem autem servorum tuorum dabo tibi quamcumque praeceperis; scis enim quoniam non est in populo meo vir, qui noverit ligna caedere sicut Sidonii ".
1KGS|5|21|Cum ergo audisset Hiram verba Salomonis, laetatus est valde et ait: " Benedictus Dominus hodie, qui dedit David filium sapientissimum super populum hunc plurimum ".
1KGS|5|22|Et misit Hiram ad Salomonem dicens: " Audivi, quaecumque mandasti mihi; ego faciam omnem voluntatem tuam in lignis cedrinis et abiegnis.
1KGS|5|23|Servi mei deponent ea de Libano ad mare, et ego componam ea in ratibus in mari usque ad locum, quem significaveris mihi, et applicabo ea ibi, et tu tolles ea; praebebisque necessaria mihi, ut detur cibus domui meae ".
1KGS|5|24|Itaque Hiram dabat Salomoni ligna cedrina et ligna abiegna iuxta omnem voluntatem eius.
1KGS|5|25|Salomon autem praebebat Hiram viginti milia chororum tritici in cibum domui eius et viginti choros purissimi olei; haec tribuebat Salomon Hiram per annos singulos.
1KGS|5|26|Dedit quoque Dominus sapientiam Salomoni, sicut locutus est ei; et erat pax inter Hiram et Salomonem, et percusserunt foedus ambo.
1KGS|5|27|Elegitque rex Salomon operas de omni Israel, et erat indictio triginta milia virorum.
1KGS|5|28|Mittebatque eos in Libanum decem milia per menses singulos vicissim, ita ut duobus mensibus essent in domibus suis; et Adoniram erat super huiuscemodi indictione.
1KGS|5|29|Fueruntque Salomoni septuaginta milia eorum, qui onera portabant, et octoginta milia latomorum in monte,
1KGS|5|30|absque praepositis, qui praeerant singulis operibus numero trium milium et trecentorum praecipientium populo, his, qui faciebant opus.
1KGS|5|31|Praecepitque rex, ut tollerent lapides grandes, lapides pretiosos in fundamentum templi, lapides quadratos;
1KGS|5|32|dolaverunt ergo caementarii Salomonis, caementarii Hiram et Giblii ligna et lapides et praeparaverunt ad aedificandam domum.
1KGS|6|1|Factum est igitur quadringente simo et octogesimo anno egres sionis filiorum Israel de terra Aegypti, in anno quarto, mense Ziv - ipse est mensis secundus - regni Salomonis super Israel, aedificare coepit domum Domino.
1KGS|6|2|Domus autem, quam aedificabat rex Salomon Domino, habebat sexaginta cubitos in longitudine et viginti cubitos in latitudine et triginta cubitos in altitudine.
1KGS|6|3|Et porticus erat ante templum viginti cubitorum longitudinis iuxta mensuram latitudinis templi et habebat decem cubitos latitudinis ante faciem templi.
1KGS|6|4|Fecitque in templo fenestras cum marginibus et cancellis.
1KGS|6|5|Et aedificavit contra parietem templi tabulata per gyrum in parietibus domus per circuitum templi et Dabir et fecit latera in circuitu.
1KGS|6|6|Tabulatum, quod subter erat, quinque cubitos habebat latitudinis et medium tabulatum sex cubitorum latitudinis et tertium tabulatum septem habens cubitos latitudinis; gradus enim posuit in domo per circuitum forinsecus, ut non ingrederentur trabes in muros templi.
1KGS|6|7|Domus autem cum aedificaretur, lapidibus dedolatis atque perfectis aedificata est; et malleus et securis et omne ferramentum non sunt audita in domo, cum aedificaretur.
1KGS|6|8|Ostium lateris inferioris in parte erat domus dextrae, et per cochleam ascendebant in medium latus et a medio in tertium.
1KGS|6|9|Et aedificavit domum et consummavit eam; texit quoque domum laquearibus cedrinis.
1KGS|6|10|Aedificavit ergo stratum contra omnem domum quinque cubitis altitudinis et iunxit domui lignis cedrinis.
1KGS|6|11|Et factus est sermo Domini ad Salomonem dicens:
1KGS|6|12|" Domus haec, quam aedificas, si ambulaveris in praeceptis meis et iudicia mea feceris et custodieris omnia mandata mea gradiens per ea, firmabo sermonem meum tibi, quem locutus sum ad David patrem tuum;
1KGS|6|13|et habitabo in medio filiorum Israel et non derelinquam populum meum Israel ".
1KGS|6|14|Igitur aedificavit Salomon domum et consummavit eam.
1KGS|6|15|Et aedificavit parietes domus intrinsecus tabulis cedrinis; a pavimento domus usque ad summitatem parietum et usque ad laquearia operuit lignis intrinsecus et texit pavimentum domus tabulis abiegnis.
1KGS|6|16|Aedificavitque viginti cubitorum a posteriore parte templi tabulis cedrinis a pavimento usque ad superiora; et fecit ei intrinsecus Dabir, id est sancta sanctorum.
1KGS|6|17|Porro quadraginta cubitorum erat ipsum templum ante illud.
1KGS|6|18|Et cedrus in domo intrinsecus sculptas habebat colocynthidas et calices apertos florum. Omnia cedrinis tabulis vestiebantur, nec omnino lapis apparere poterat in pariete.
1KGS|6|19|Dabir autem in medio domus in interiori parte fecerat, ut poneret ibi arcam foederis Domini.
1KGS|6|20|Habebat viginti cubitos longitudinis et viginti cubitos latitudinis et viginti cubitos altitudinis; et vestivit illud auro purissimo et fecit altare cedrinum ante Dabir.
1KGS|6|21|Domum quoque operuit Salomon intrinsecus auro purissimo et posuit catenas aureas ante Dabir.
1KGS|6|22|Nihilque erat in templo, quod non auro tegeretur; sed et totum altare Dabir texit auro.
1KGS|6|23|Et fecit in Dabir duos cherubim de lignis oleastri decem cubitorum altitudinis.
1KGS|6|24|Quinque cubitorum ala cherub una et quinque cubitorum ala cherub altera, id est decem cubitos habentes a summitate alae unius usque ad alae alterius summitatem.
1KGS|6|25|Decem quoque cubitorum erat cherub secundus, mensura par et effigies una erat duobus cherubim;
1KGS|6|26|altitudinem habebat unus cherub decem cubitorum et similiter cherub secundus.
1KGS|6|27|Posuitque cherubim in medio templi interioris; extendebant autem alas suas cherubim, et tangebat ala una parietem et ala cherub secundi tangebat parietem alterum; alae autem alterae in media parte templi se invicem contingebant.
1KGS|6|28|Texit quoque cherubim auro.
1KGS|6|29|Et omnes parietes templi per circuitum scalpsit variis caelaturis; et fecit in eis cherubim et palmas et calices apertos florum intrinsecus et foras.
1KGS|6|30|Sed et pavimentum domus texit auro intrinsecus et extrinsecus.
1KGS|6|31|Et pro ingressu Dabir fecit valvas de lignis oleastri postesque cum marginibus quinque.
1KGS|6|32|Et in duabus valvis de lignis oleastri scalpsit cherubim et palmas et calices apertos florum et vestivit ea auro operiens tam cherubim quam palmas et cetera auro.
1KGS|6|33|Fecitque eodem modo pro introitu templi postes cum quattuor marginibus de lignis oleastri
1KGS|6|34|et duas valvas de lignis abiegnis; et utraque valva duplex erat et versatilis.
1KGS|6|35|Et scalpsit cherubim et palmas et calices apertos florum operuitque omnia laminis aureis.
1KGS|6|36|Et aedificavit atrium interius tribus ordinibus lapidum politorum et uno ordine lignorum cedri.
1KGS|6|37|Anno quarto fundata est domus Domini in mense Ziv;
1KGS|6|38|et in anno undecimo, mense Bul - ipse est mensis octavus - perfecta est domus in omni opere suo et in universis utensilibus; aedificavitque eam annis septem.
1KGS|7|1|Domum autem suam aedificavit Salomon tredecim annis et ad perfectum usque perduxit.
1KGS|7|2|Aedificavit quoque domum Saltus Libani centum cubitorum longitudinis et quinquaginta cubitorum latitudinis et triginta cubitorum altitudinis super quattuor ordines columnarum cedrinarum, et ligna cedrina super columnas.
1KGS|7|3|Et erat tectum cedrinum in alto super tabulas quadraginta quinque, quae erant super columnas, quindecim in uno ordine,
1KGS|7|4|et marginum tres ordines, fenestra iuxta fenestram tribus vicibus.
1KGS|7|5|Ostia, id est postes, habebant quadruplicem marginem.
1KGS|7|6|Et porticum columnarum fecit quinquaginta cubitorum longitudinis et triginta cubitorum latitudinis, et alteram porticum in facie maioris porticus et columnas et cancellos ante eas.
1KGS|7|7|Porticum quoque solii, in qua tribunal erat, fecit et texit lignis cedrinis a pavimento usque ad pavimentum.
1KGS|7|8|Et domus, in qua habitabat, erat in altero atrio intro a porticu et simili opere. Domum quoque fecit filiae pharaonis, quam uxorem duxerat Salomon, tali opere quali et hanc porticum.
1KGS|7|9|Omnia lapidibus pretiosis, qui ad normam quandam atque mensuram tam intrinsecus quam extrinsecus serrati erant, a fundamento usque ad summitatem parietum, et extrinsecus usque ad atrium maius.
1KGS|7|10|Fundamenta autem de lapidibus pretiosis, lapidibus magnis decem sive octo cubitorum.
1KGS|7|11|Et desuper lapides pretiosi secundum mensuram secti et ligna cedrina.
1KGS|7|12|Et atrium maius in circuitu habebat tres ordines de lapidibus sectis et unum ordinem de dolata cedro; necnon et atrium domus Domini interius et porticus domus.
1KGS|7|13|Misit quoque rex Salomon et tulit Hiram de Tyro,
1KGS|7|14|filium mulieris viduae de tribu Nephthali, patre Tyrio, artificem aerarium et plenum sapientia et intellegentia et doctrina ad faciendum omne opus ex aere. Qui, cum venisset ad regem Salomonem, fecit omne opus eius.
1KGS|7|15|Et finxit duas columnas aereas, decem et octo cubitorum altitudinis columnam unam, et linea duodecim cubitorum ambiebat columnam, et grossitudo eius quattuor digitorum, et intrinsecus cava erat; sic et columna altera.
1KGS|7|16|Duo quoque capitella fecit, quae ponerentur super capita columnarum, fusili aere; quinque cubitorum altitudinis capitellum unum et quinque cubitorum altitudinis capitellum alterum,
1KGS|7|17|et serta quasi in modum texturae, fimbriae in modum catenarum sibi invicem miro opere contextarum in capitellis, quae erant super caput columnarum, septem in capitello uno et septem in capitello altero.
1KGS|7|18|Et fecit malogranatorum duos ordines per circuitum super sertum unum, ut tegerent capitella, quae erant super summitatem columnarum; eodem modo fecit et capitello secundo.
1KGS|7|19|Capitella autem, quae erant super capita columnarum, quasi opere lilii fabricata erant in porticu, quattuor cubitorum.
1KGS|7|20|Et rursum alia capitella in summitate duarum columnarum etiam desuper, iuxta alvum, quae erat super sertum. Malogranatorum autem ducentorum duo ordines erant in circuitu capitelli primi et eodem modo in circuitu capitelli secundi.
1KGS|7|21|Et statuit duas columnas in porticum templi; cumque statuisset columnam dexteram, vocavit eam nomine Iachin, similiter erexit columnam sinistram et vocavit nomen eius Booz.
1KGS|7|22|Et super capita columnarum opus in modum lilii posuit; per fectumque est opus columnarum.
1KGS|7|23|Fecit quoque mare fusile decem cubitorum a labio usque ad labium, rotundum in circuitu, quinque cubitorum altitudo eius; et resticula triginta cubitorum cingebat illud per circuitum.
1KGS|7|24|Et scalptura colocynthidum subter labium circuibat illud, duo ordines scalpturarum fusilium in una fusione cum mari.
1KGS|7|25|Et stabat super duodecim boves, e quibus tres respiciebant ad aquilonem et tres ad occidentem et tres ad meridiem et tres ad orientem, et mare super eos desuper erat; quorum posteriora universa intrinsecus latitabant.
1KGS|7|26|Grossitudo autem luteris habebat mensuram palmi, labiumque eius erat quasi labium calicis et folium repandi lilii; duo milia batos capiebat.
1KGS|7|27|Et fecit bases decem aereas, quattuor cubitorum longitudinis bases singulas et quattuor cubitorum latitudinis et trium cubitorum altitudinis.
1KGS|7|28|Hoc autem erat opus basium: limbos habebant, insuper et limbos inter columellas.
1KGS|7|29|Super limbos inter columellas erant leones et boves et cherubim, et super columellas similiter; supra et infra leones et boves erant coronae, opus malleatum.
1KGS|7|30|Et quattuor rotae per bases singulas et axes aerei, et quattuor pedes et quasi umeruli subter luterem fusiles, contra singulos coronae.
1KGS|7|31|Et os eius erat rotundum, opus basis, unius cubiti et dimidii; etiam in ore eius variae caelaturae erant, limbi autem eius erant quadrati, non rotundi.
1KGS|7|32|Quattuor quoque rotae subter limbis erant, et fulcra rotarum cohaerebant basi; una rota habebat altitudinis cubitum et semis.
1KGS|7|33|Tales autem rotae erant, quales solent in curru fieri, et fulcra earum et canthi et radii et modioli, omnia fusilia.
1KGS|7|34|Nam et umeruli illi quattuor per singulos angulos basis unius ex ipsa basi fusiles et coniuncti erant.
1KGS|7|35|In summitate autem basis erat quaedam rotunditas dimidii cubiti, et in summitate basis fulcra eius et limbi eius ex semetipsa.
1KGS|7|36|Scalpsit quoque in tabulatis illis, fulcris eius et super limbos eius cherubim et leones et palmas secundum vacuum singulorum, et coronas per circuitum.
1KGS|7|37|In hunc modum fecit decem bases, fusura una, et mensura scalpturaque consimili.
1KGS|7|38|Fecit quoque decem luteres aereos; quadraginta batos capiebat luter unus, eratque quattuor cubitorum; singulosque luteres per singulas, id est decem bases posuit.
1KGS|7|39|Et constituit decem bases, quinque ad dexteram partem templi et quinque ad sinistram; mare autem posuit ad dexteram partem templi contra orientem ad meridiem.
1KGS|7|40|Fecit quoque Hiram lebetes et vatilla et phialas et perfecit omne opus regi Salomoni in templo Domini;
1KGS|7|41|columnas duas et globos capitellorum super capita columnarum duos et serta duo, ut operirent duos globos, qui erant super capita columnarum;
1KGS|7|42|et malogranata quadringenta in duobus sertis, duos versus malogranatorum in sertis singulis, ad operiendos globos capitellorum, qui erant super faciem columnarum;
1KGS|7|43|et bases decem et luteres decem super bases
1KGS|7|44|et mare unum et boves duodecim subter mare;
1KGS|7|45|et lebetes et vatilla et phialas. Omnia vasa, quae fecit Hiram regi Salomoni in domo Domini, de aere polito erant.
1KGS|7|46|In campestri regione Iordanis fudit ea rex in argillosa terra inter Succoth et Sarthan.
1KGS|7|47|Et posuit Salomon omnia vasa; propter multitudinem autem nimiam ignorabatur pondus aeris.
1KGS|7|48|Fecitque Salomon omnia vasa in domo Domini: altare aureum et mensam, super quam ponerentur panes propositionis, auream;
1KGS|7|49|et candelabra, quinque ad dexteram et quinque ad sinistram contra Dabir, ex auro puro, et florem et lucernas desuper aureas; et forcipes aureos
1KGS|7|50|et pateras et cultros et phialas et sartagines et turibula de auro purissimo; et cardines ostiorum domus interioris Sancti sanctorum et ostiorum domus templi ex auro.
1KGS|7|51|Et perfecit omne opus, quod faciebat Salomon in domo Domini, et intulit Salomon, quae sanctificaverat David pater suus, argentum et aurum et vasa, reposuitque in thesauris domus Domini.
1KGS|8|1|Tunc congregavit Salomon om nes maiores natu Israel - om nes principes tribuum, duces familiarum filiorum Israel ad regem Salomonem - in Ierusalem, ut deferrent arcam foederis Domini de civitate David, id est de Sion.
1KGS|8|2|Convenitque ad regem Salomonem universus Israel in mense Ethanim in sollemnitate, ipse est mensis septimus.
1KGS|8|3|Veneruntque cuncti senes Israel, et tulerunt sacerdotes arcam
1KGS|8|4|et portaverunt arcam Domini et tabernaculum conventus et omnia vasa sanctuarii, quae erant in tabernaculo; et ferebant ea sacerdotes et Levitae.
1KGS|8|5|Rex autem Salomon et universus coetus Israel, qui convenerat ad eum, cum illo ante arcam immolabant oves et boves absque aestimatione et numero.
1KGS|8|6|Et intulerunt sacerdotes arcam foederis Domini in locum suum in Dabir templi, in sanctum sanctorum, subter alas cherubim;
1KGS|8|7|siquidem cherubim expandebant alas super locum arcae et protegebant arcam et vectes eius desuper.
1KGS|8|8|Cumque eminerent vectes et apparerent summitates eorum foris in sanctuario ante Dabir, non apparebant ultra extrinsecus; qui et fuerunt ibi usque in praesentem diem.
1KGS|8|9|In arca autem non erat aliud nisi duae tabulae lapideae, quas posuerat in ea Moyses in Horeb, quando pepigit Dominus foedus cum filiis Israel, cum egrederentur de terra Aegypti.
1KGS|8|10|Factum est autem cum exissent sacerdotes de sanctuario, nebula implevit domum Domini,
1KGS|8|11|et non poterant sacerdotes stare et ministrare propter nebulam; impleverat enim gloria Domini domum Domini.
1KGS|8|12|Tunc ait Salomon: Dominus dixit ut habitaret in nebula.
1KGS|8|13|Aedificans aedificavi domum in habitaculum tuum,firmissimum solium tuum in sempiternum ".
1KGS|8|14|Convertitque rex faciem suam et benedixit omni ecclesiae Israel; omnis enim ecclesia Israel stabat.
1KGS|8|15|Et ait: " Benedictus Dominus, Deus Israel, qui locutus est ore suo ad David patrem meum et in manibus suis perfecit dicens:
1KGS|8|16|"A die qua eduxi populum meum Israel de Aegypto, non elegi civitatem de universis tribubus Israel, ut aedificaretur domus, et esset nomen meum ibi; sed elegi David, ut esset super populum meum Israel".
1KGS|8|17|Voluitque David pater meus aedificare domum nomini Domini, Dei Israel,
1KGS|8|18|et ait Dominus ad David patrem meum: "Quod cogitasti in corde tuo aedificare domum nomini meo, bene fecisti hoc ipsum mente tractans;
1KGS|8|19|verumtamen tu non aedificabis domum sed filius tuus, qui egredietur de lumbis tuis, ipse aedificabit domum nomini meo".
1KGS|8|20|Confirmavit Dominus sermonem suum, quem locutus est; stetique pro David patre meo et sedi super thronum Israel, sicut locutus est Dominus, et aedificavi domum nomini Domini, Dei Israel.
1KGS|8|21|Et constitui ibi locum arcae, in qua foedus est Domini, quod percussit cum patribus nostris, quando eduxit eos de terra Aegypti ".
1KGS|8|22|Stetit autem Salomon ante altare Domini in conspectu omnis ecclesiae Israel et expandit manus suas in caelum
1KGS|8|23|et ait: " Domine, Deus Israel, non est similis tui Deus in caelo desuper et super terra deorsum, qui custodis pactum et misericordiam servis tuis, qui ambulant coram te in toto corde suo;
1KGS|8|24|qui custodisti servo tuo David patri meo, quae locutus es ei; ore locutus es et manibus perfecisti, ut et haec dies probat.
1KGS|8|25|Nunc igitur, Domine, Deus Israel, conserva famulo tuo David patri meo, quae locutus es ei dicens: "Non auferetur de te vir coram me, qui sedeat super thronum Israel, ita tamen, si custodierint filii tui viam suam, ut ambulent coram me, sicut tu ambulasti in conspectu meo".
1KGS|8|26|Et nunc, Domine, Deus Israel, firmentur verba tua, quae locutus es servo tuo David patri meo.
1KGS|8|27|Ergone putandum est quod vere Deus habitet super terram? Si enim caelum et caeli caelorum te capere non possunt, quanto magis domus haec, quam aedificavi!
1KGS|8|28|Sed respice ad orationem servi tui et ad preces eius, Domine Deus meus; audi clamorem et orationem, quam servus tuus orat coram te hodie,
1KGS|8|29|ut sint oculi tui aperti super domum hanc nocte ac die, super locum, de quo dixisti: "Erit nomen meum ibi", ut exaudias orationem, qua orat te servus tuus in loco isto,
1KGS|8|30|ut exaudias deprecationem servi tui et populi tui Israel, quodcumque oraverint in loco isto, et exaudies in loco habitaculi tui in caelo et, cum exaudieris, propitius eris.
1KGS|8|31|Si peccaverit homo in proximum suum et habuerit aliquod iuramentum, quo teneatur astrictus, et venerit propter iuramentum coram altari tuo in domum istam,
1KGS|8|32|tu exaudies in caelo et facies et iudicabis servos tuos condemnans impium et reddens viam suam super caput eius iustificansque iustum et retribuens ei secundum iustitiam suam.
1KGS|8|33|Si superatus fuerit populus tuus Israel ab inimicis suis, quia peccaturus est tibi, et agentes paenitentiam et confitentes nomini tuo venerint et oraverint et deprecati te fuerint in domo hac,
1KGS|8|34|exaudi in caelo et dimitte peccatum populi tui Israel et reduces eos in terram, quam dedisti patribus eorum.
1KGS|8|35|Si clausum fuerit caelum et non pluerit propter peccata eorum, et oraverint in loco isto confessi nomini tuo et a peccatis suis conversi propter afflictionem suam,
1KGS|8|36|exaudi eos in caelo et dimitte peccata servorum tuorum et populi tui Israel et ostende eis viam bonam, per quam ambulent, et da pluviam super terram tuam, quam dedisti populo tuo in possessionem.
1KGS|8|37|Fames si oborta fuerit in terra aut pestilentia aut uredo aut aurugo aut locusta vel bruchus, et afflixerit eum inimicus eius portas obsidens, omnis plaga, universa infirmitas,
1KGS|8|38|cuncta oratio et deprecatio, quae acciderit omni homini de populo tuo Israel; si quis cognoverit plagam cordis sui et expanderit manus suas in domo hac,
1KGS|8|39|tu audies in caelo in loco habitationis tuae et repropitiaberis et facies, ut des unicuique secundum omnes vias suas, sicut videris cor eius, quia tu nosti solus cor omnium filiorum hominum,
1KGS|8|40|ut timeant te cunctis diebus, quibus vivunt super faciem terrae, quam dedisti patribus nostris.
1KGS|8|41|Insuper et alienigena, qui non est de populo tuo Israel, cum venerit de terra longinqua propter nomen tuum
1KGS|8|42|- audietur enim nomen tuum magnum et manus tua fortis et brachium tuum extentum ubique - cum venerit ergo et oraverit in hoc loco,
1KGS|8|43|tu exaudies in caelo in loco habitationis tuae et facies omnia, pro quibus invocaverit te alienigena, ut sciant universi populi terrarum nomen tuum et timeant te, sicut populus tuus Israel, et probent quia nomen tuum invocatum est super domum hanc, quam aedificavi.
1KGS|8|44|Si egressus fuerit populus tuus ad bellum contra inimicos suos per viam, quocumque miseris eos, et oraverint te contra viam civitatis, quam elegisti, et contra domum, quam aedificavi nomini tuo,
1KGS|8|45|exaudies in caelo orationes eorum et preces eorum et facies iudicium eorum.
1KGS|8|46|Quod si peccaverint tibi - non est enim homo qui non peccet - et iratus tradideris eos inimicis suis, et captivi ducti fuerint in terram inimicorum longe vel prope
1KGS|8|47|et egerint paenitentiam in corde suo in loco captivitatis et conversi deprecati te fuerint in captivitate sua dicentes: "Peccavimus, inique egimus, impie gessimus";
1KGS|8|48|et reversi fuerint ad te in universo corde suo et tota anima sua in terra inimicorum suorum, ad quam captivi ducti sunt, et oraverint te contra viam terrae suae, quam dedisti patribus eorum, et civitatis, quam elegisti, et templi, quod aedificavi nomini tuo,
1KGS|8|49|exaudies in caelo in firmamento solii tui orationes eorum et preces eorum et facies iudicium eorum;
1KGS|8|50|et propitiaberis populo tuo, qui peccavit tibi, et omnibus iniquitatibus eorum, quibus praevaricati sunt in te, et dabis misericordiam coram eis, qui eos captivos habuerint, ut misereantur eis
1KGS|8|51|- populus enim tuus est et hereditas tua, quos eduxisti de terra Aegypti de medio fornacis ferreae -
1KGS|8|52|ut sint oculi tui aperti ad deprecationem servi tui et populi tui Israel, et exaudias eos in universis, pro quibus invocaverint te.
1KGS|8|53|Tu enim separasti eos tibi in hereditatem de universis populis terrae, sicut locutus es per Moysen servum tuum, quando eduxisti patres nostros de Aegypto, Domine Deus ".
1KGS|8|54|Factum est autem cum complesset Salomon orans Dominum omnem orationem et deprecationem hanc, surrexit de conspectu altaris Domini; utrumque enim genu in terram fixerat et manus expanderat in caelum.
1KGS|8|55|Stetit ergo et benedixit omni ecclesiae Israel voce magna dicens:
1KGS|8|56|" Benedictus Dominus, qui dedit requiem populo suo Israel iuxta omnia, quae locutus est; non cecidit ne unus quidem sermo ex omnibus bonis, quae locutus est per Moysen servum suum.
1KGS|8|57|Sit Dominus Deus noster nobiscum, sicut fuit cum patribus nostris, non derelinquens nos neque proiciens,
1KGS|8|58|sed inclinet corda nostra ad se, ut ambulemus in universis viis eius et custodiamus mandata eius et decreta et iudicia, quaecumque mandavit patribus nostris.
1KGS|8|59|Et sint sermones mei isti, quibus deprecatus sum coram Domino, appropinquantes Domino Deo nostro die ac nocte, ut faciat iudicium servo suo et populo suo Israel per singulos dies,
1KGS|8|60|ut sciant omnes populi terrae quia Dominus ipse est Deus, et non est ultra absque eo.
1KGS|8|61|Sit quoque cor vestrum perfectum cum Domino Deo nostro, ut ambuletis in decretis eius et custodiatis mandata eius sicut et hodie ".
1KGS|8|62|Igitur rex et omnis Israel cum eo immolabant victimas coram Domino.
1KGS|8|63|Mactavitque Salomon hostias pacificas, quas immolavit Domino, boum viginti duo milia et ovium centum viginti milia. Et dedicaverunt templum Domini rex et omnes filii Israel.
1KGS|8|64|In die illa sanctificavit rex medium atrii, quod erat ante domum Domini; fecit quippe holocaustum ibi et oblationem et adipem pacificorum, quoniam altare aereum, quod erat coram Domino, minus erat et capere non poterat holocaustum et oblationem et adipem pacificorum.
1KGS|8|65|Fecit ergo Salomon in tempore illo festivitatem celebrem, et omnis Israel cum eo, ecclesia magna ab introitu Emath usque ad rivum Aegypti, coram Domino Deo nostro septem diebus.
1KGS|8|66|Et in die octava dimisit populos; qui benedicentes regi profecti sunt in tabernacula sua laetantes et alacri corde super omnibus bonis, quae fecerat Dominus David servo suo et Israel populo suo.
1KGS|9|1|Factum est autem cum perfecisset Salomon aedificium domus Domini et aedificium regis et omne, quod optaverat et voluerat facere,
1KGS|9|2|apparuit ei Dominus secundo, sicut apparuerat ei in Gabaon.
1KGS|9|3|Dixitque Dominus ad eum: " Exaudivi orationem tuam et deprecationem tuam, quam deprecatus es coram me; sanctificavi domum hanc, quam aedificasti, ut ponerem nomen meum ibi in sempiternum; et erunt oculi mei et cor meum ibi cunctis diebus.
1KGS|9|4|Tu quoque, si ambulaveris coram me, sicut ambulavit David pater tuus in simplicitate cordis et in aequitate, et feceris omnia, quae praecepi tibi, et legitima mea et iudicia mea servaveris,
1KGS|9|5|ponam thronum regni tui super Israel in sempiternum, sicut locutus sum David patri tuo dicens: Non auferetur de genere tuo vir de solio Israel.
1KGS|9|6|Si autem aversione aversi fueritis vos et filii vestri non sequentes me nec custodientes mandata mea et decreta mea, quae proposui vobis, sed abieritis et colueritis deos alienos et adoraveritis eos,
1KGS|9|7|auferam Israel de superficie terrae, quam dedi eis, et templum, quod sanctificavi nomini meo, proiciam a conspectu meo; eritque Israel in proverbium et in fabulam cunctis populis,
1KGS|9|8|et domus haec erit in ruinas. Omnis, qui transierit per eam, stupebit et sibilabit et dicet: "Quare fecit Dominus sic terrae huic et domui huic?".
1KGS|9|9|Et respondebunt: "Quia dereliquerunt Dominum Deum suum, qui eduxit patres eorum de terra Aegypti, et secuti sunt deos alienos et adoraverunt eos et coluerunt eos; idcirco induxit Dominus super eos omne malum hoc" ".
1KGS|9|10|Expletis autem annis viginti, postquam aedificaverat Salomon duas domos, id est domum Domini et domum regis
1KGS|9|11|- Hiram rege Tyri praebente Salomoni ligna cedrina et abiegna et aurum iuxta omne quod opus habuerat - tunc dedit Salomon Hiram viginti oppida in terra Galilaeae.
1KGS|9|12|Et egressus est Hiram de Tyro, ut videret oppida, quae dederat ei Salomon, et non placuerunt ei;
1KGS|9|13|et ait: " Haeccine sunt civitates, quas dedisti mihi, frater? ". Et appellavit eas terram Chabul usque in diem hanc.
1KGS|9|14|Misit quoque Hiram ad regem centum viginti talenta auri.
1KGS|9|15|Haec est summa indictionis, quam constituit rex Salomon ad aedificandam domum Domini et domum suam et Mello et murum Ierusalem et Asor et Mageddo et Gazer.
1KGS|9|16|Pharao rex Aegypti ascendit et cepit Gazer succenditque eam igni et Chananaeum, qui habitabat in civitate, interfecit; et dedit eam in dotem filiae suae uxori Salomonis.
1KGS|9|17|Aedificavit ergo Salomon Gazer et Bethoron inferiorem
1KGS|9|18|et Baalath et Thamar in terra solitudinis
1KGS|9|19|et omnes civitates horreorum, quae ad se pertinebant, et civitates curruum et civitates equorum et quodcumque ei placuit, ut aedificaret in Ierusalem et in Libano et in omni terra potestatis suae.
1KGS|9|20|Universum populum, qui remanserat de Amorraeis et Hetthaeis et Pherezaeis et Hevaeis et Iebusaeis, qui non erant de filiis Israel,
1KGS|9|21|horum filios, qui remanserant post eos in terra, quos scilicet non potuerant filii Israel exterminare, fecit Salomon tributarios usque in diem hanc.
1KGS|9|22|De filiis autem Israel non constituit Salomon servire quemquam, sed erant viri bellatores et ministri eius et principes et pugnatores eius et praefecti curruum et equitum.
1KGS|9|23|Erant autem principes eorum, qui super omnia opera Salomonis praepositi erant, quingenti quinquaginta; qui habebant subiectum populum et statutis operibus imperabant.
1KGS|9|24|Filia autem pharaonis ascendit de civitate David in domum suam, quam aedificaverat ei; tunc aedificavit Mello.
1KGS|9|25|Offerebat quoque Salomon tribus vicibus per annos singulos holocausta et pacificas victimas super altare, quod aedificaverat Domino, et adolebat coram Domino; perfectumque est templum.
1KGS|9|26|Classem quoque fecit rex Salomon in Asiongaber, quae est iuxta Ailath in litore maris Rubri in terra Idumaea.
1KGS|9|27|Misitque Hiram in classe illa servos suos viros nauticos gnaros maris cum servis Salomonis.
1KGS|9|28|Qui, cum venissent in Ophir, sumptum inde aurum quadringentorum viginti talentorum detulerunt ad regem Salomonem.
1KGS|10|1|Sed et regina Saba, audita fama Salomonis - in hono rem nominis Domini - venit tentare eum in aenigmatibus.
1KGS|10|2|Et ingressa Ierusalem multo cum comitatu et divitiis, camelis portantibus aromata et aurum infinitum nimis et gemmas pretiosas, venit ad Salomonem et locuta est ei universa, quae habebat in corde suo.
1KGS|10|3|Et docuit eam Salomon omnia verba, quae proposuerat: non fuit sermo, qui regem posset latere, et non responderet ei.
1KGS|10|4|Videns autem regina Saba omnem sapientiam Salomonis et domum, quam aedificaverat,
1KGS|10|5|et cibos mensae eius et sessionem servorum et ordinem ministrantium vestesque eorum et pincernas et holocausta, quae offerebat in domo Domini, non habebat ultra spiritum
1KGS|10|6|dixitque ad regem: " Verus est sermo, quem audivi in terra mea super rebus tuis et super sapientia tua!
1KGS|10|7|Et non credebam narrantibus mihi, donec ipsa veni et vidi oculis meis et probavi quod media pars mihi nuntiata non fuerit; maior est sapientia et bona tua quam rumor, quem audivi.
1KGS|10|8|Beati viri tui et beati servi tui hi, qui stant coram te semper et audiunt sapientiam tuam!
1KGS|10|9|Sit Dominus Deus tuus benedictus, cui placuisti, et posuit te super thronum Israel, eo quod dilexerit Dominus Israel in sempiternum et constituit te regem, ut faceres iudicium et iustitiam ".
1KGS|10|10|Dedit ergo regi centum viginti talenta auri et aromata multa nimis et gemmas pretiosas; non sunt allata ultra aromata tam multa quam ea, quae dedit regina Saba regi Salomoni.
1KGS|10|11|Sed et classis Hiram, quae portabat aurum de Ophir, attulit ex Ophir ligna thyina multa nimis et gemmas pretiosas.
1KGS|10|12|Fecitque rex de lignis thyinis fulcra domus Domini et domus regiae et citharas lyrasque cantoribus. Non sunt allata huiuscemodi ligna thyina neque visa usque in praesentem diem.
1KGS|10|13|Rex autem Salomon dedit reginae Saba omnia, quae voluit et petivit ab eo, praeter ea, quae ultro obtulerat ei munere regio. Quae reversa est et abiit in terram suam cum servis suis.
1KGS|10|14|Erat autem pondus auri, quod afferebatur Salomoni per annos singulos, sescentorum sexaginta sex talentorum auri,
1KGS|10|15|praeter id, quod proveniebat ex tributis subiectorum et commercio negotiatorum et omnium regum Arabiae et ducum terrae.
1KGS|10|16|Fecit quoque rex Salomon ducenta scuta de auro puro, sescentos auri siclos dedit in laminas scuti unius;
1KGS|10|17|et trecentas peltas ex auro probato, tres minae auri unam peltam vestiebant; posuitque ea rex in domo Saltus Libani.
1KGS|10|18|Fecit etiam rex Salomon thronum de ebore grandem et vestivit eum auro fulvo nimis.
1KGS|10|19|Qui habebat sex gradus, et summitas throni rotunda erat in parte posteriori, et duae manus hinc atque inde tenentes sedile, et duo leones stabant iuxta manus;
1KGS|10|20|et duodecim leunculi stantes super sex gradus hinc atque inde. Non est factum tale opus in universis regnis.
1KGS|10|21|Sed et omnia vasa, quibus potabat rex Salomon, erant aurea, et universa supellex domus Saltus Libani de auro purissimo; non erat argentum nec alicuius pretii putabatur in diebus Salomonis,
1KGS|10|22|quia classis Tharsis, quae regi erat, per mare cum classe Hiram semel per tres annos redibat deferens aurum et argentum et ebur et simias et pavos.
1KGS|10|23|Magnificatus est ergo rex Salomon super omnes reges terrae divitiis et sapientia.
1KGS|10|24|Et universa terra desiderabat vultum Salomonis, ut audiret sapientiam eius, quam dederat Deus in corde eius.
1KGS|10|25|Et singuli deferebant ei munera, vasa argentea et aurea, vestes et arma bellica, aromata quoque et equos et mulos per annos singulos.
1KGS|10|26|Congregavitque Salomon currus et equites, et facti sunt ei mille quadringenti currus et duodecim milia equitum; et disposuit eos per civitates quadrigarum et cum rege in Ierusalem.
1KGS|10|27|Fecitque ut tanta esset abundantia argenti in Ierusalem quanta et lapidum; et cedrorum praebuit multitudinem quasi sycomoros, quae nascuntur in Sephela.
1KGS|10|28|Et educebantur equi Salomoni de Aegypto et de Coa; negotiatores enim regis emebant de Coa statuto pretio.
1KGS|10|29|Constabat autem et egrediebatur quadriga ex Aegypto sescentis siclis argenti, et equus centum quinquaginta; atque in hunc modum cunctis regibus Hetthaeorum et Syriae per manus suas venundabant.
1KGS|11|1|Rex autem Salomon amavit mulieres alienigenas multas, filiam quoque pharaonis et Moabitidas et Ammonitidas, Idumaeas et Sidonias et Hetthaeas,
1KGS|11|2|de gentibus, super quibus dixit Dominus filiis Israel: " Non ingrediemini ad eas, neque de illis ingredientur ad vestras; certissime enim avertent corda vestra, ut sequamini deos earum ". His itaque copulatus est Salomon amore;
1KGS|11|3|fueruntque ei uxores quasi reginae septingentae et concubinae trecentae, et averterunt mulieres cor eius.
1KGS|11|4|Cumque iam esset senex, depravatum est cor eius per mulieres, ut sequeretur deos alienos; nec erat cor eius perfectum cum Domino Deo suo sicut cor David patris eius,
1KGS|11|5|sed colebat Salomon Astharthen, deam Sidoniorum, et Melchom idolum Ammonitarum.
1KGS|11|6|Fecitque Salomon quod non placuerat coram Domino et non adimplevit ut sequeretur Dominum sicut David pater eius.
1KGS|11|7|Tunc aedificavit Salomon fanum Chamos idolo Moab in monte, qui est contra Ierusalem, et Melchom idolo filiorum Ammon;
1KGS|11|8|atque in hunc modum fecit universis uxoribus suis alienigenis, quae adolebant et immolabant diis suis.
1KGS|11|9|Igitur iratus est Dominus Salomoni, quod aversa esset mens eius a Domino, Deo Israel, qui apparuerat ei bis
1KGS|11|10|et praeceperat de verbo hoc, ne sequeretur deos alienos; et non custodivit, quae mandavit ei Dominus.
1KGS|11|11|Dixit itaque Dominus Salomoni: " Quia habuisti hoc apud te et non custodisti pactum meum et praecepta mea, quae mandavi tibi, disrumpens scindam regnum tuum a te et dabo illud servo tuo.
1KGS|11|12|Verumtamen in diebus tuis non faciam propter David patrem tuum; de manu filii tui scindam illud.
1KGS|11|13|Nec totum regnum auferam, sed tribum unam dabo filio tuo propter David servum meum et Ierusalem, quam elegi ".
1KGS|11|14|Suscitavit autem Dominus adversarium Salomoni Adad Idumaeum, qui erat de semine regio, in Edom.
1KGS|11|15|Cum enim vicisset David Idumaeam, et ascendisset Ioab princeps militiae ad sepeliendum eos, qui fuerant interfecti, et occidisset omne masculinum in Idumaea
1KGS|11|16|- sex enim mensibus ibi moratus est Ioab et omnis Israel, donec interimerent omne masculinum in Idumaea -
1KGS|11|17|fugit Adad ipse et viri Idumaei de servis patris eius cum eo, ut ingrederetur Aegyptum; erat autem Adad puer parvulus.
1KGS|11|18|Cumque surrexissent de Madian, venerunt in Pharan tuleruntque secum viros de Pharan et introierunt Aegyptum ad pharaonem regem Aegypti, qui dedit ei domum et cibos constituit et terram delegavit.
1KGS|11|19|Et invenit Adad gratiam coram pharao valde, in tantum ut daret ei uxorem sororem uxoris suae germanam Taphnes reginae.
1KGS|11|20|Genuitque ei soror Taphnes Genubath filium et ablactavit eum Taphnes in domo pharaonis, eratque Genubath habitans apud pharaonem cum filiis eius.
1KGS|11|21|Cumque audisset Adad in Aegypto dormisse David cum patribus suis et mortuum esse Ioab principem militiae, dixit pharaoni: " Dimitte me, ut vadam in terram meam ".
1KGS|11|22|Dixitque ei pharao: " Qua enim re apud me indiges, ut quaeras ire ad terram tuam? ". At ille respondit: " Nulla; sed obsecro, ut dimittas me ".
1KGS|11|23|Suscitavit quoque Deus Salomoni adversarium Razon filium Eliada, qui fugerat ab Adadezer rege Soba domino suo.
1KGS|11|24|Et congregavit ad se viros et factus est princeps turmae, cum interficeret eos David; abieruntque Damascum et habitaverunt ibi et regnaverunt in Damasco.
1KGS|11|25|Eratque adversarius Israeli cunctis diebus Salomonis; et hoc cum malo, quod erat Adad. Et detestatus est Israel regnavitque in Syria.
1KGS|11|26|Ieroboam quoque filius Nabat, Ephrathaeus de Sareda, servus Salomonis, cuius mater erat nomine Sarva mulier vidua, levavit manum contra regem.
1KGS|11|27|Et haec causa rebellionis adversus eum: Salomon aedificavit Mello et coaequavit voraginem civitatis David patris sui.
1KGS|11|28|Erat autem Ieroboam vir fortis et strenuus; vidensque Salomon adulescentem industrium constituerat eum praefectum super labores universae domus Ioseph.
1KGS|11|29|Factum est igitur in tempore illo, ut Ieroboam egrederetur de Ierusalem, et inveniret eum Ahias Silonites propheta in via opertus pallio novo; erant autem duo tantum in agro.
1KGS|11|30|Apprehendensque Ahias pallium suum novum, quo coopertus erat, scidit in duodecim partes
1KGS|11|31|et ait ad Ieroboam: " Tolle tibi decem scissuras; haec enim dicit Dominus, Deus Israel: Ecce ego scindam regnum de manu Salomonis et dabo tibi decem tribus.
1KGS|11|32|Porro una tribus remanebit ei propter servum meum David et Ierusalem civitatem, quam elegi ex omnibus tribubus Israel;
1KGS|11|33|eo quod dereliquerint me et adoraverint Astharthen deam Sidoniorum et Chamos deum Moab et Melchom deum filiorum Ammon et non ambulaverint in viis meis, ut facerent iustitiam coram me et praecepta mea et iudicia sicut David pater eius.
1KGS|11|34|Nec auferam omne regnum de manu eius, sed ducem ponam eum cunctis diebus vitae suae propter David servum meum, quem elegi, qui custodivit mandata mea et praecepta mea.
1KGS|11|35|Auferam autem regnum de manu filii eius et dabo tibi decem tribus;
1KGS|11|36|filio autem eius dabo tribum unam, ut remaneat lucerna David servo meo cunctis diebus coram me in Ierusalem civitate, quam elegi, ut esset nomen meum ibi.
1KGS|11|37|Te autem assumam, et regnabis super omnia, quae desiderat anima tua, erisque rex super Israel.
1KGS|11|38|Si igitur audieris omnia, quae praecepero tibi, et ambulaveris in viis meis et feceris, quod rectum est coram me custodiens mandata mea et praecepta mea, sicut fecit David servus meus, ero tecum et aedificabo tibi domum stabilem, quomodo aedificavi David, et tradam tibi Israel
1KGS|11|39|et affligam semen David super hoc, verumtamen non cunctis diebus ".
1KGS|11|40|Voluit ergo Salomon interficere Ieroboam, qui surrexit et aufugit in Aegyptum ad Sesac regem Aegypti et fuit in Aegypto usque ad mortem Salomonis.
1KGS|11|41|Reliqua autem gestorum Salomonis, omnia, quae fecit, et sapientia eius, ecce universa scripta sunt in libro gestorum Salomonis;
1KGS|11|42|dies autem, quos regnavit Salomon in Ierusalem super omnem Israel, quadraginta anni sunt.
1KGS|11|43|Dormivitque Salomon cum patribus suis et sepultus est in civitate David patris sui; regnavitque Roboam filius eius pro eo.
1KGS|12|1|Venit autem Roboam in Sichem; illuc enim congregatus erat omnis Israel ad constituendum eum regem.
1KGS|12|2|At Ieroboam filius Nabat, cum adhuc esset in Aegypto profugus a facie regis Salomonis, audito hoc nuntio, reversus est de Aegypto.
1KGS|12|3|Miseruntque et vocaverunt eum. Venit ergo Ieroboam et omnis multitudo Israel, et locuti sunt ad Roboam dicentes:
1KGS|12|4|" Pater tuus durissimum iugum imposuit nobis; tu itaque nunc imminue paululum de imperio patris tui durissimo et de iugo gravissimo, quod imposuit nobis, et serviemus tibi ".
1KGS|12|5|Qui ait eis: " Ite usque ad tertium diem et revertimini ad me ".Cumque abisset populus,
1KGS|12|6|iniit consilium rex Roboam cum senioribus, qui assistebant coram Salomone patre eius, cum adhuc viveret, et ait: " Quod mihi datis consilium, ut respondeam populo huic? ".
1KGS|12|7|Qui dixerunt ei: " Si hodie oboedieris populo huic et servieris et petitioni eorum cesseris locutusque fueris ad eos verba lenia, erunt tibi servi cunctis diebus ".
1KGS|12|8|Qui dereliquit consilium senum, quod dederant ei, et adhibuit adulescentes, qui nutriti fuerant cum eo et assistebant illi,
1KGS|12|9|dixitque ad eos: " Quod mihi datis consilium, ut respondeam populo huic, qui dixerunt mihi: "Levius fac iugum, quod imposuit pater tuus super nos"?.
1KGS|12|10|Et dixerunt ei iuvenes, qui nutriti fuerant cum eo: " Sic loquere populo huic, qui locuti sunt ad te dicentes: "Pater tuus aggravavit iugum nostrum, tu releva nos"; sic loqueris ad eos: Minimus digitus meus grossior est lumbis patris mei.
1KGS|12|11|Et nunc, pater meus posuit super vos iugum grave, ego autem addam super iugum vestrum; pater meus cecidit vos flagellis, ego autem caedam scorpionibus ".
1KGS|12|12|Venit ergo Ieroboam et omnis populus ad Roboam die tertia, sicut locutus fuerat rex dicens: " Revertimini ad me die tertia ".
1KGS|12|13|Responditque rex populo dura, derelicto consilio seniorum, quod ei dederant,
1KGS|12|14|et locutus est eis secundum consilium iuvenum dicens: Pater meus aggravavit iugum vestrum,ego autem addam iugo vestro;pater meus cecidit vos flagellis,ego autem caedam vos scorpionibus ".
1KGS|12|15|Ergo non acquievit rex populo, quoniam dispositum erat a Domino, ut suscitaret verbum suum, quod locutus fuerat in manu Ahiae Silonitae ad Ieroboam filium Nabat.
1KGS|12|16|Videns itaque omnis Israel quod noluisset eos audire rex, respondit ei dicens: Quae nobis pars in David,vel quae hereditas in filio Isai?Vade in tabernacula tua, Israel!Nunc vide domum tuam, David! ". Et abiit Israel in tabernacula sua.
1KGS|12|17|Super filios autem Israel, quicumque habitabant in civitatibus Iudae, regnavit Roboam.
1KGS|12|18|Misit rex Roboam Adoniram, qui erat super servitutem; et lapidavit eum omnis Israel, et mortuus est. Porro rex Roboam festinus ascendit currum et fugit in Ierusalem.
1KGS|12|19|Recessitque Israel a domo David usque in praesentem diem.
1KGS|12|20|Factum est autem cum audisset omnis Israel quod reversus esset Ieroboam, miserunt et vocaverunt eum, congregato coetu, et constituerunt eum regem super omnem Israel; nec secutus est quisquam domum David praeter tribum Iudae solam.
1KGS|12|21|Venit autem Roboam Ierusalem et congrcgavit universam domum Iudae et tribum Beniamin, centum octoginta milia electorum virorum bellatorum, ut pugnaret contra domum Israel et reduceret regnum Roboam filio Salomonis.
1KGS|12|22|Factus est vero sermo Domini ad Semeiam virum Dei dicens:
1KGS|12|23|" Loquere ad Roboam filium Salomonis regem Iudae et ad omnem domum Iudae et Beniamin et reliquos de populo dicens:
1KGS|12|24|Haec dicit Dominus: Non ascendetis neque bellabitis contra fratres vestros, filios Israel; revertatur vir in domum suam; a me enim factum est hoc ". Audierunt sermonem Domini et reversi sunt de itinere, sicut eis praeceperat Dominus.
1KGS|12|25|Aedificavit autem Ieroboam Sichem in monte Ephraim et habitavit ibi; et egressus inde aedificavit Phanuel.
1KGS|12|26|Dixitque Ieroboam in corde suo: " Nunc revertetur regnum ad domum David,
1KGS|12|27|si ascenderit populus iste, ut faciat sacrificia in domo Domini in Ierusalem, et convertetur cor populi huius ad dominum suum Roboam regem Iudae, interficientque me et revertentur ad Roboam regem Iudae ".
1KGS|12|28|Et excogitato consilio, fecit rex duos vitulos aureos et dixit ad populum: " Nolite ultra ascendere in Ierusalem! Ecce dii tui, Israel, qui te eduxerunt de terra Aegypti ".
1KGS|12|29|Posuitque unum in Bethel et alterum donavit in Dan;
1KGS|12|30|et factum est hoc in peccatum: ibat enim populus coram uno usque in Dan.
1KGS|12|31|Et fecit fana in excelsis et sacerdotes de extremis populi, qui non erant de filiis Levi.
1KGS|12|32|Constituitque diem sollemnem in mense octavo, quinta decima die mensis, in similitudinem sollemnitatis, quae celebratur in Iuda. Et ascendit altare; sic fecit in Bethel, ut immolaret vitulis, quos fabricatus erat; constituitque in Bethel sacerdotes excelsorum, quae fecerat.
1KGS|12|33|Et ascendit super altare, quod exstruxerat in Bethel, quinta decima die mensis octavi, quem finxerat de corde suo; et fecit sollemnitatem filiis Israel et ascendit super altare, ut adoleret.
1KGS|13|1|Et ecce vir Dei venit de Iuda in sermone Domini in Bethel, Ieroboam stante super altare ad adolendum;
1KGS|13|2|et exclamavit contra altare in sermone Domini et ait: " Altare, altare, haec dicit Dominus: Ecce filius nascetur domui David, Iosias nomine, et immolabit super te sacerdotes excelsorum, qui nunc in te immolant, et ossa hominum super te incendent ".
1KGS|13|3|Deditque in illa die signum dicens: " Hoc erit signum, quod locutus est Dominus: ecce altare scindetur, et effundetur cinis, qui in eo est ".
1KGS|13|4|Cumque audisset rex sermonem hominis Dei, quem inclamaverat contra altare in Bethel, extendit manum suam de altari dicens: " Apprehendite eum! ". Et exaruit manus eius, quam extenderat contra eum, nec valuit retrahere eam ad se.
1KGS|13|5|Altare quoque scissum est, et effusus est cinis de altari iuxta signum, quod praedixerat vir Dei in sermone Domini.
1KGS|13|6|Et ait rex ad virum Dei: " Deprecare faciem Domini Dei tui et ora pro me, ut restituatur manus mea mihi ". Oravit vir Dei faciem Domini, et reversa est manus regis ad eum et facta est sicut prius fuerat.
1KGS|13|7|Locutus est autem rex ad virum Dei: " Veni mecum domum, ut prandeas, et dabo tibi munera ".
1KGS|13|8|Responditque vir Dei ad regem: " Si dederis mihi mediam partem domus tuae, non veniam tecum nec comedam panem neque bibam aquam in loco isto;
1KGS|13|9|sic enim mandatum est mihi in sermone Domini praecipientis: "Non comedes panem neque bibes aquam nec reverteris per viam, qua venisti" ".
1KGS|13|10|Abiit ergo per aliam viam et non est reversus per iter, quo venerat in Bethel.
1KGS|13|11|Prophetes autem quidam senex habitabat in Bethel; ad quem venerunt filii sui et narraverunt ei omnia opera, quae fecerat vir Dei illa die in Bethel, et verba, quae locutus fuerat ad regem, narraverunt quoque patri suo.
1KGS|13|12|Et dixit eis pater eorum: " Per quam viam abiit? ". Ostenderunt ei filii sui viam, per quam abierat vir Dei, qui venerat de Iuda.
1KGS|13|13|Et ait filiis suis: " Sternite mihi asinum ". Qui cum stravissent, ascendit
1KGS|13|14|et abiit post virum Dei et invenit eum sedentem subtus terebinthum et ait illi: " Tune es vir Dei, qui venisti de Iuda?". Respondit ille: " Ego sum ".
1KGS|13|15|Dixit ad eum: " Veni mecum domum, ut comedas panem ".
1KGS|13|16|Qui ait: " Non possum reverti neque venire tecum nec comedam panem neque bibam aquam in loco isto;
1KGS|13|17|sic enim dictum est mihi in sermone Domini: "Non comedes panem et non bibes ibi aquam nec reverteris per viam, qua ieris" ".
1KGS|13|18|Qui ait illi: " Et ego propheta sum similis tui; et angelus locutus est mihi in sermone Domini dicens: "Reduc eum tecum in domum tuam, et comedat panem et bibat aquam" ". Fefellit eum
1KGS|13|19|et reduxit secum; comedit ergo panem in domo eius et bibit aquam.
1KGS|13|20|Cumque sederent ad mensam, factus est sermo Domini ad prophetam, qui reduxerat eum,
1KGS|13|21|et exclamavit ad virum Dei, qui venerat de Iuda, dicens: " Haec dicit Dominus: Quia non oboediens fuisti ori Domini et non custodisti mandatum, quod praecepit tibi Dominus Deus tuus,
1KGS|13|22|et reversus es et comedisti panem et bibisti aquam in loco, in quo praecepit tibi, ne comederes panem neque biberes aquam, non inferetur cadaver tuum in sepulcrum patrum tuorum ".
1KGS|13|23|Cumque comedisset panem et bibisset, stravit sibi asinum prophetae, qui reduxerat eum;
1KGS|13|24|et, cum abisset, invenit eum leo in via et occidit, et erat cadaver eius proiectum in itinere; asinus autem stabat iuxta illum, et leo stabat iuxta cadaver.
1KGS|13|25|Et ecce viri transeuntes viderunt cadaver proiectum in via et leonem stantem iuxta cadaver; et venerunt et divulgaverunt in civitate, in qua prophetes ille senex habitabat.
1KGS|13|26|Quod cum audisset propheta ille, qui reduxerat eum de via, ait: " Vir Dei est, qui inoboediens fuit ori Domini, et tradidit eum Dominus leoni; et confregit eum et occidit iuxta verbum Domini, quod locutus est ei ".
1KGS|13|27|Dixitque ad filios suos: " Sternite mihi asinum! ". Qui cum stravissent,
1KGS|13|28|et ille abisset, invenit cadaver eius proiectum in via et asinum et leonem stantes iuxta cadaver; non comedit leo de cadavere nec laesit asinum.
1KGS|13|29|Tulit ergo prophetes cadaver viri Dei et posuit illud super asinum et reversus intulit in civitatem prophetae senis, ut plangerent eum et sepelirent.
1KGS|13|30|Et posuit cadaver eius in sepulcro suo, et planxerunt eum: " Heu, heu, mi frater! ".
1KGS|13|31|Cumque sepelissent eum, dixit ad filios suos: " Cum mortuus fuero, sepelite me in sepulcro, in quo vir Dei sepultus est; iuxta ossa eius ponite ossa mea.
1KGS|13|32|Profecto enim veniet sermo, quem praedixit in sermone Domini contra altare, quod est in Bethel, et contra omnia fana excelsorum, quae sunt in urbibus Samariae ".
1KGS|13|33|Post haec non est reversus Ieroboam de via sua pessima, sed iterum faciebat de novissimis populi sacerdotes excelsorum; quicumque volebat, implebat eius manum, ut fieret sacerdos excelsorum.
1KGS|13|34|Et propter hanc causam peccavit domus Ieroboam, et eversa est et deleta de superficie terrae.
1KGS|14|1|In tempore illo aegrotavit Abia filius Ieroboam,
1KGS|14|2|dixitque Ieroboam uxori suae: " Surge et commuta habitum, ne cognoscaris quod sis uxor Ieroboam, et vade in Silo, ubi est Ahias propheta, qui locutus est mihi quod regnaturus essem super populum hunc.
1KGS|14|3|Tolle quoque in manu tua decem panes et crustula et vas mellis et vade ad illum: ipse indicabit tibi quid eventurum sit puero ".
1KGS|14|4|Fecit, ut dixerat, uxor Ieroboam et consurgens abiit in Silo et venit in domum Ahiae; at ille non poterat videre, quia caligaverant oculi eius prae senectute.
1KGS|14|5|Dixerat autem Dominus ad Ahiam: " Ecce uxor Ieroboam ingredietur, ut consulat te super filio suo, qui aegrotat; haec et haec loqueris ei. Cum intret, simulabit se peregrinam esse ".
1KGS|14|6|Cum ergo audiret Ahias sonitum pedum eius introeuntis per ostium, ait: " Ingredere, uxor Ieroboam. Quare aliam te esse simulas? Ego autem missus sum ad te durus nuntius.
1KGS|14|7|Vade et dic Ieroboam: "Haec dicit Dominus, Deus Israel: Quia exaltavi te de medio populi et dedi te ducem super populum meum Israel
1KGS|14|8|et scidi regnum a domo David et dedi illud tibi, et non fuisti sicut servus meus David, qui custodivit mandata mea et secutus est me in toto corde suo faciens quod placitum esset in conspectu meo,
1KGS|14|9|sed operatus es mala super omnes, qui fuerunt ante te, et fecisti tibi deos alienos et conflatiles, ut me ad iracundiam provocares, me autem proiecisti post tergum tuum:
1KGS|14|10|idcirco ecce ego inducam mala super domum Ieroboam et percutiam de Ieroboam quidquid masculini sexus, impuberem et puberem in Israel; et mundabo reliquias domus Ieroboam, sicut mundari solet fimus usque ad purum.
1KGS|14|11|Qui mortui fuerint de Ieroboam in civitate, comedent eos canes; qui autem mortui fuerint in agro, vorabunt eos aves caeli, quia Dominus locutus est.
1KGS|14|12|Tu igitur surge et vade in domum tuam, et in ipso introitu pedum tuorum in urbem morietur puer,
1KGS|14|13|et planget eum omnis Israel et sepeliet; iste enim solus inferetur de Ieroboam in sepulcrum, quia inventum est in eo, quod bonum erat Domino, Deo Israel, in domo Ieroboam.
1KGS|14|14|Constituet autem sibi Dominus regem super Israel, qui percutiat domum Ieroboam.
1KGS|14|15|Et percutiet Dominus Israel, ut moveatur sicut arundo in aqua, et evellet Israel de terra bona hac, quam dedit patribus eorum; et ventilabit eos trans Flumen, quia fecerunt sibi palos, ut irritarent Dominum.
1KGS|14|16|Et tradet Dominus Israel propter peccata Ieroboam, qui peccavit et peccare fecit Israel" ".
1KGS|14|17|Surrexit itaque uxor Ieroboam et abiit et venit in Thersa; cumque illa ingrederetur limen domus, puer mortuus est.
1KGS|14|18|Et sepelierunt eum, et planxit illum omnis Israel iuxta sermonem Domini, quem locutus est in manu servi sui Ahiae prophetae.
1KGS|14|19|Reliqua autem gestorum Ieroboam, quomodo pugnaverit et quomodo regnaverit, ecce scripta sunt in libro annalium regum Israel.
1KGS|14|20|Dies autem, quibus regnavit Ieroboam, viginti duo anni sunt; et dormivit cum patribus suis. Regnavitque Nadab filius eius pro eo.
1KGS|14|21|Porro Roboam filius Salomonis regnavit in Iuda. Quadraginta et unius anni erat Roboam, cum regnare coepisset, et decem et septem annos regnavit in Ierusalem civitate, quam elegit Dominus, ut poneret nomen suum ibi ex omnibus tribubus Israel. Nomen autem matris eius Naama Ammanites.
1KGS|14|22|Et fecit Iuda malum coram Domino, et irritaverunt eum super omnibus, quae fecerant patres eorum in peccatis suis, quae peccaverant;
1KGS|14|23|aedificaverunt enim et ipsi sibi excelsa et lapides et palos super omnem collem excelsum et subter omnem arborem frondosam.
1KGS|14|24|Sed et prostibula fuerunt in terra; feceruntque omnes abominationes gentium, quas attrivit Dominus ante faciem filiorum Israel.
1KGS|14|25|In quinto autem anno regni Roboam ascendit Sesac rex Aegypti in Ierusalem
1KGS|14|26|et tulit thesauros domus Domini et thesauros regios et universa diripuit, scuta quoque aurea omnia, quae fecerat Salomon.
1KGS|14|27|Pro quibus fecit rex Roboam scuta aerea et tradidit ea in manu ducum cursorum, qui excubabant ante ostium domus regis.
1KGS|14|28|Cumque ingrederetur rex in domum Domini, portabant ea cursores et postea reportabant ad armamentarium cursorum.
1KGS|14|29|Reliqua autem gestorum Roboam et omnia, quae fecit, ecce scripta sunt in libro annalium regum Iudae.
1KGS|14|30|Fuitque bellum inter Roboam et Ieroboam cunctis diebus.
1KGS|14|31|Dormivit itaque Roboam cum patribus suis et sepultus est cum eis in civitate David; nomen autem matris eius Naama Ammanites. Et regnavit Abiam filius eius pro eo.
1KGS|15|1|Igitur in octavo decimo anno regni Ieroboam filii Nabat regnavit Abiam super Iudam.
1KGS|15|2|Tribus annis regnavit in Ierusalem; nomen matris eius Maacha filia Abessalom.
1KGS|15|3|Ambulavitque in omnibus peccatis patris sui, quae fecerat ante eum; nec erat cor eius perfectum cum Domino Deo suo sicut cor David patris eius.
1KGS|15|4|Sed propter David dedit ei Dominus Deus suus lucernam in Ierusalem, ut suscitaret filium eius post eum et statueret Ierusalem;
1KGS|15|5|eo quod fecisset David rectum in oculis Domini et non declinasset ab omnibus, quae praeceperat ei, cunctis diebus vitae suae, excepta re Uriae Hetthaei. (6)
1KGS|15|6|attamen bellum fuit inter Roboam et inter Hieroboam omni tempore vitae eius
1KGS|15|7|Reliqua autem gestorum Abiam et omnia, quae fecit, nonne haec scripta sunt in libro annalium regum Iudae? Fuitque bellum inter Abiam et inter Ieroboam.
1KGS|15|8|Et dormivit Abiam cum patribus suis, et sepelierunt eum in civitate David; regnavitque Asa filius eius pro eo.
1KGS|15|9|In anno ergo vicesimo Ieroboam regis Israel regnavit Asa rex Iudae
1KGS|15|10|et quadraginta et uno anno regnavit in Ierusalem. Nomen matris eius Maacha filia Abessalom.
1KGS|15|11|Et fecit Asa rectum ante conspectum Domini sicut David pater eius.
1KGS|15|12|Et abstulit prostibula de terra purgavitque universas sordes idolorum, quae fecerant patres eius.
1KGS|15|13|Insuper et Maacham matrem suam amovit, ne esset domina, eo quod fecisset abominationem Aserae; confregitque Asa simulacrum turpissimum et combussit in torrente Cedron.
1KGS|15|14|Excelsa autem non abstulit; verumtamen cor Asa perfectum erat coram Domino cunctis diebus suis.
1KGS|15|15|Et intulit ea, quae sanctificaverat pater suus et quae ipse voverat, in domum Domini, argentum et aurum et vasa.
1KGS|15|16|Bellum autem erat inter Asa et Baasa regem lsrael cunctis diebus eorum.
1KGS|15|17|Ascendit quoque Baasa rex Israel in Iudam et aedificavit Rama, ut non posset quispiam egredi vel ingredi de parte Asa regis Iudae.
1KGS|15|18|Tollens itaque Asa omne argentum et aurum, quod remanserat in thesauris domus Domini et in thesauris domus regiae, dedit illud in manu servorum suorum et misit ad Benadad filium Tabremmon filii Hezion regem Syriae, qui habitabat in Damasco, dicens:
1KGS|15|19|" Foedus est inter me et te et inter patrem meum et patrem tuum; ideo misi tibi munera, argentum et aurum, et peto, ut irritum facias foedus, quod habes cum Baasa rege Israel, et recedat a me ".
1KGS|15|20|Acquiescens Benadad regi Asa misit principes exercituum suorum in civitates Israel, et percusserunt Ahion et Dan et Abelbethmaacha et universam Chenereth cum omni terra Nephthali.
1KGS|15|21|Quod cum audisset Baasa, cessavit aedificare Rama et reversus est in Thersa.
1KGS|15|22|Rex autem Asa convocavit omnem Iudam, nullo excusato; et tulerunt lapides Rama et ligna eius, quibus aedificaverat Baasa, et exstruxit de eis rex Asa Gabaa Beniamin et Maspha.
1KGS|15|23|Reliqua autem omnium gestorum Asa et universa fortitudo eius et cuncta, quae fecit, et civitates, quas exstruxit, nonne haec scripta sunt in libro annalium regum Iudae? Verumtamen in tempore senectutis suae doluit pedes;
1KGS|15|24|et dormivit cum patribus suis et sepultus est cum eis in civitate David patris sui. Regnavitque Iosaphat filius eius pro eo.
1KGS|15|25|Nadab vero filius Ieroboam regnavit super Israel anno secundo Asa regis Iudae; regnavitque super Israel duobus annis.
1KGS|15|26|Et fecit, quod malum est in conspectu Domini, et ambulavit in viis patris sui et in peccato eius, quo peccare fecit Israel.
1KGS|15|27|Insidiatus est autem ei Baasa filius Ahiae de domo Issachar et percussit eum in Gebbethon, quae est urbs Philisthinorum; siquidem Nadab et omnis Israel obsidebant Gebbethon.
1KGS|15|28|Interfecit igitur illum Baasa in anno tertio Asa regis Iudae et regnavit pro eo.
1KGS|15|29|Cumque regnasset, percussit omnem domum Ieroboam; non dimisit ne unam quidem animam de semine eius, donec deleret eam iuxta verbum Domini, quod locutus fuerat in manu servi sui Ahiae Silonitis
1KGS|15|30|propter peccata Ieroboam, quae peccaverat et quibus peccare fecerat Israel, et propter delictum, quo irritaverat Dominum, Deum Israel.
1KGS|15|31|Reliqua autem gestorum Nadab et omnia, quae fortiter operatus est, nonne haec scripta sunt in libro annalium regum Israel?
1KGS|15|32|Fuitque bellum inter Asa et Baasa regem Israel cunctis diebus eorum.
1KGS|15|33|Anno tertio Asa regis Iudae regnavit Baasa filius Ahiae super omnem Israel in Thersa viginti quattuor annis;
1KGS|15|34|et fecit malum coram Domino ambulavitque in via Ieroboam et in peccato eius, quo peccare fecit Israel.
1KGS|16|1|Factus est autem sermo Domini ad Iehu filium Hanani contra Baasa dicens:
1KGS|16|2|" Pro eo quod exaltavi te de pulvere et posui te ducem super populum meum Israel, tu autem ambulasti in via Ieroboam et peccare fecisti populum meum Israel, ut me irritares in peccatis eorum,
1KGS|16|3|ecce ego demetam posteriora Baasa et posteriora domus eius et faciam domum tuam sicut domum Ieroboam filii Nabat.
1KGS|16|4|Qui mortuus fuerit de Baasa in civitate, comedent eum canes; et, qui mortuus fuerit ex eo in agro, comedent eum volucres caeli".
1KGS|16|5|Reliqua autem gestorum Baasa et quaecumque fecit et fortitudo eius, nonne haec scripta sunt in libro annalium regum Israel?
1KGS|16|6|Dormivit ergo Baasa cum patribus suis sepultusque est in Thersa; et regnavit Ela filius eius pro eo.
1KGS|16|7|Sed et in manu Iehu filii Hanani prophetae verbum Domini factum est ad Baasa et ad domum eius propter omne malum, quod fecerat coram Domino ad irritandum eum in operibus manuum suarum, ut fieret sicut domus Ieroboam, eo quod percussisset eam.
1KGS|16|8|Anno vicesimo sexto Asa regis Iudae regnavit Ela filius Baasa super Israel in Thersa duobus annis.
1KGS|16|9|Et rebellavit contra eum servus suus Zamri dux mediae partis curruum. Erat autem Ela in Thersa bibens et temulentus in domo Arsa praefecti domus in Thersa;
1KGS|16|10|irruens ergo Zamri percussit et occidit eum anno vicesimo septimo Asa regis Iudae et regnavit pro eo.
1KGS|16|11|Cumque regnasset et sedisset super solium eius, percussit omnem domum Baasa et non dereliquit ex eo quidquid masculini sexus et propinquos et amicos eius.
1KGS|16|12|Delevitque Zamri omnem domum Baasa iuxta verbum Domini, quod locutus fuerat ad Baasa in manu Iehu prophetae,
1KGS|16|13|propter universa peccata Baasa et peccata Ela filii eius, qui peccaverunt et peccare fecerunt Israel provocantes Dominum, Deum Israel, in vanitatibus suis.
1KGS|16|14|Reliqua autem gestorum Ela et omnia, quae fecit, nonne haec scripta sunt in libro annalium regum Israel?
1KGS|16|15|Anno vicesimo septimo Asa regis Iudae regnavit Zamri septem diebus in Thersa. Porro exercitus obsidebat Gebbethon urbem Philisthinorum.
1KGS|16|16|Cumque audisset rebellasse Zamri et occidisse regem, fecit sibi regem omnis Israel Amri, qui erat princeps militiae super Israel in die illa in castris.
1KGS|16|17|Ascendit ergo Amri et omnis Israel cum eo de Gebbethon, et obsidebant Thersa;
1KGS|16|18|videns autem Zamri quod expugnanda esset civitas, ingressus est palatium et succendit super se domum regiam et mortuus est igne
1KGS|16|19|in peccatis suis, quae peccaverat faciens malum coram Domino et ambulans in via Ieroboam et in peccato eius, quo fecit peccare Israel.
1KGS|16|20|Reliqua autem gestorum Zamri et rebellio, quam fecit, nonne haec scripta sunt in libro annalium regum Israel?
1KGS|16|21|Tunc divisus est populus Israel in duas partes: media pars populi sequebatur Thebni filium Gineth, ut constitueret eum regem, et media pars Amri.
1KGS|16|22|Praevaluit autem populus, qui erat cum Amri, populo, qui sequebatur Thebni filium Gineth; mortuusque est Thebni, et regnavit Amri.
1KGS|16|23|Anno tricesimo primo Asa regis Iudae regnavit Amri super Israel duodecim annis; in Thersa regnavit sex annis.
1KGS|16|24|Emitque montem Samariae a Somer duobus talentis argenti et aedificavit eum et vocavit nomen civitatis, quam exstruxerat, nomine Somer domini montis Samariae.
1KGS|16|25|Fecit autem Amri malum in conspectu Domini et operatus est nequiter super omnes, qui fuerunt ante eum;
1KGS|16|26|ambulavitque in omni via Ieroboam filii Nabat et in peccato eius, quo peccare fecerat Israel, ut irritaret Dominum, Deum Israel, in vanitatibus suis.
1KGS|16|27|Reliqua autem gestorum Amri et proelia eius, quae fortiter gessit, nonne haec scripta sunt in libro annalium regum Israel?
1KGS|16|28|Et dormivit Amri cum patribus suis et sepultus est in Samaria; regnavitque Achab filius eius pro eo.
1KGS|16|29|Achab vero filius Amri regnavit super Israel anno tricesimo octavo Asa regis Iudae; et regnavit Achab filius Amri super Israel in Samaria viginti et duobus annis.
1KGS|16|30|Et fecit Achab filius Amri malum in conspectu Domini super omnes, qui fuerunt ante eum.
1KGS|16|31|Nec suffecit ei, ut ambularet in peccatis Ieroboam filii Nabat; insuper duxit uxorem Iezabel filiam Ethbaal regis Sidoniorum et abiit et servivit Baal et adoravit eum.
1KGS|16|32|Et posuit aram Baal in templo Baal, quod aedificaverat in Samaria,
1KGS|16|33|et fecit Achab palum. Et addidit Achab in opere suo irritans Dominum, Deum Israel, super omnes reges Israel, qui fuerant ante eum.
1KGS|16|34|In diebus eius aedificavit Hiel de Bethel Iericho; in Abiram primitivo suo fundavit eam et in Segub novissimo suo posuit portas eius, iuxta verbum Domini, quod locutus fuerat in manu Iosue filii Nun.
1KGS|17|1|Et dixit Elias Thesbites de Thesbi in Galaad ad Achab: " Vivit Dominus, Deus Israel, in cuius conspectu sto. Non erit annis his ros et pluvia, nisi iuxta oris mei verba! ".
1KGS|17|2|Et factum est verbum Domini ad eum dicens:
1KGS|17|3|" Recede hinc et vade contra orientem et abscondere in torrente Charith, qui est contra Iordanem,
1KGS|17|4|et ibi de torrente bibes; corvisque praecepi, ut pascant te ibi ".
1KGS|17|5|Abiit ergo et fecit iuxta verbum Domini; cumque abisset, sedit in torrente Charith, qui est contra Iordanem.
1KGS|17|6|Corvi quoque deferebant ei panem et carnes mane, similiter panem et carnes vesperi; et bibebat de torrente.
1KGS|17|7|Post dies autem siccatus est torrens; non enim pluerat super terram.
1KGS|17|8|Factus est igitur sermo Domini ad eum dicens:
1KGS|17|9|" Surge et vade in Sarepta Sidoniorum et manebis ibi; praecepi enim ibi mulieri viduae, ut pascat te ".
1KGS|17|10|Surrexit et abiit Sareptam. Cumque venisset ad portam civitatis, apparuit ei mulier vidua colligens ligna; et vocavit eam dixitque: " Da mihi paululum aquae in vase, ut bibam ".
1KGS|17|11|Cumque illa pergeret, ut afferret, clamavit post tergum eius dicens: " Affer mihi, obsecro, et buccellam panis in manu tua ".
1KGS|17|12|Quae respondit: " Vivit Dominus Deus tuus, non habeo panem, nisi quantum pugillus capere potest farinae in hydria et paululum olei in lecytho. En colligo duo ligna, ut ingrediar et faciam illud mihi et filio meo, ut comedamus et moriamur ".
1KGS|17|13|Ad quam Elias ait: " Noli timere, sed vade et fac, sicut dixisti; verumtamen mihi primum fac de ipsa farinula subcinericium panem parvulum et affer ad me; tibi autem et filio tuo facies postea.
1KGS|17|14|Haec autem dicit Dominus, Deus Israel: "Hydria farinae non deficiet, nec lecythus olei minuetur usque ad diem, in qua daturus est Dominus pluviam super faciem terrae" ".
1KGS|17|15|Quae abiit et fecit iuxta verbum Eliae et comedit illa et ipse et domus eius per dies.
1KGS|17|16|Hydria farinae non defecit, et lecythus olei non est imminutus iuxta verbum Domini, quod locutus fuerat in manu Eliae.
1KGS|17|17|Factum est autem post haec, aegrotavit filius mulieris matris familiae; et erat languor fortis nimis, ita ut non remaneret in eo halitus.
1KGS|17|18|Dixit ergo ad Eliam: " Quid mihi et tibi, vir Dei? Ingressus es ad me, ut rememorarentur iniquitates meae, et interficeres filium meum? ".
1KGS|17|19|Et ait ad eam: " Da mihi filium tuum ". Tulitque eum de sinu illius et portavit in cenaculum, ubi ipse manebat, et posuit super lectulum suum;
1KGS|17|20|clamavitque ad Dominum et dixit: " Domine Deus meus, etiamne viduam, apud quam ego ut hospes habito, afflixisti, ut interficeres filium eius?.
1KGS|17|21|Et expandit se atque mensus est super puerum tribus vicibus et clamavit ad Dominum et ait: " Domine Deus meus, revertatur, oro, anima pueri huius in viscera eius ".
1KGS|17|22|Et exaudivit Dominus vocem Eliae, et reversa est anima pueri intra eum, et revixit.
1KGS|17|23|Tulitque Elias puerum et deposuit eum de cenaculo in inferiorem domum et tradidit matri suae et ait illi: " En vivit filius tuus ".
1KGS|17|24|Dixitque mulier ad Eliam: " Nunc in isto cognovi quoniam vir Dei es tu, et verbum Domini in ore tuo verum est ".
1KGS|18|1|Post dies multos factum est verbum Domini ad Eliam in anno tertio dicens: " Vade et ostende te Achab, ut dem pluviam super faciem terrae ".
1KGS|18|2|Ivit ergo Elias, ut ostenderet se Achab.Erat autem fames vehemens in Samaria.
1KGS|18|3|Vocavitque Achab Abdiam dispensatorem domus suae. Abdias autem timebat Dominum valde;
1KGS|18|4|nam, cum interficeret Iezabel prophetas Domini, tulit ille centum prophetas et abscondit eos quinquagenos et quinquagenos in speluncis et pavit eos pane et aqua.
1KGS|18|5|Dixit ergo Achab ad Abdiam: " Vade in terra ad universos fontes aquarum et in cunctas valles, si forte invenire possimus herbam, ut salvemus equos et mulos et nullum de iumentis interficere debeamus ".
1KGS|18|6|Diviseruntque sibi regiones, ut circuirent eas: Achab ibat per viam unam, et Abdias per viam alteram seorsum.
1KGS|18|7|Cumque esset Abdias in via, Elias occurrit ei; qui cum cognovisset eum, cecidit super faciem suam et ait: " Num tu es, domine mi, Elias? ".
1KGS|18|8|Cui ille respondit: " Ego. Vade, dic domino tuo: "Adest Elias" ".
1KGS|18|9|Et ille: " Quid peccavi, inquit, quoniam trades me servum tuum in manu Achab, ut interficiat me?
1KGS|18|10|Vivit Dominus Deus tuus, non est gens aut regnum, quo non miserit dominus meus te requirens et, respondentibus cunctis: "Non est hic", adiuravit regna singula et gentes, eo quod minime reperireris.
1KGS|18|11|Et nunc dicis mihi: "Vade et dic domino tuo: Adest Elias".
1KGS|18|12|Cumque recessero a te, spiritus Domini asportabit te in locum, quem ego ignoro; et ingressus nuntiabo Achab, et non inveniet te et interficiet me. Servus autem tuus timet Dominum ab infantia sua.
1KGS|18|13|Numquid non indicatum est domino meo quid fecerim, cum interficeret Iezabel prophetas Domini: quod absconderim de prophetis Domini centum viros, quinquagenos et quinquagenos in speluncis et paverim eos pane et aqua?
1KGS|18|14|Et nunc tu dicis: "Vade et dic domino tuo: Adest Elias", ut interficiat me ".
1KGS|18|15|Dixit Elias: " Vivit Dominus exercituum ante cuius vultum sto: hodie apparebo ei ".
1KGS|18|16|Abiit ergo Abdias in occursum Achab et indicavit ei.Venitque Achab in occursum Eliae
1KGS|18|17|et, cum vidisset eum, ait: " Tune es, qui conturbas Israel? ".
1KGS|18|18|Et ille ait: " Non turbavi Israel, sed tu et domus patris tui, qui dereliquistis mandata Domini, et secutus es Baalim.
1KGS|18|19|Verumtamen nunc mitte et congrega ad me universum Israel in monte Carmeli et prophetas Baal quadringentos quinquaginta prophetasque Aserae quadringentos, qui comedunt de mensa Iezabel ".
1KGS|18|20|Misit Achab ad omnes filios Israel et congregavit prophetas in monte Carmeli.
1KGS|18|21|Accedens autem Elias ad omnem populum ait: " Usquequo claudicatis in duas partes? Si Dominus est Deus, sequimini eum; si autem Baal, sequimini illum ". Et non respondit ei populus verbum.
1KGS|18|22|Et ait rursus Elias ad populum: " Ego remansi propheta Domini solus; prophetae autem Baal quadringenti et quinquaginta viri sunt.
1KGS|18|23|Dentur nobis duo boves, et illi eligant sibi bovem unum et in frusta caedentes ponant super ligna; ignem autem non supponant. Et ego faciam bovem alterum et imponam super ligna; ignemque non supponam.
1KGS|18|24|Invocate nomen dei vestri, et ego invocabo nomen Domini; et Deus, qui exaudierit per ignem, ipse est Deus! ". Respondens omnis populus ait: " Optima propositio ".
1KGS|18|25|Dixit ergo Elias prophetis Baal: " Eligite vobis bovem unum et facite primi, quia vos plures estis; et invocate nomen dei vestri ignemque non supponatis ".
1KGS|18|26|Qui cum tulissent bovem, quem dederat eis, fecerunt et invocabant nomen Baal de mane usque ad meridiem dicentes: " Baal, exaudi nos! ". Et non erat vox, nec qui responderet. Saliebantque in circuitu altaris, quod fecerant.
1KGS|18|27|Cumque esset iam meridies, illudebat eis Elias dicens: " Clamate voce maiore; deus enim est et forsitan occupatus est aut secessit aut in itinere aut certe dormit, ut excitetur ".
1KGS|18|28|Clamabant ergo voce magna et incidebant se iuxta ritum suum cultris et lanceolis, donec perfunderentur sanguine.
1KGS|18|29|Postquam autem transiit meridies, et, illis prophetantibus, venerat tempus, quo sacrificium offerri solet, nec audiebatur vox, neque aliquis respondebat nec attendebat orantes,
1KGS|18|30|dixit Elias omni populo: " Venite ad me ". Et, accedente ad se populo, curavit altare Domini, quod destructum fuerat;
1KGS|18|31|et tulit duodecim lapides iuxta numerum tribuum filiorum Iacob, ad quem factus est sermo Domini dicens: " Israel erit nomen tuum ".
1KGS|18|32|Et aedificavit lapidibus altare in nomine Domini fecitque aquaeductum quasi pro duobus satis in circuitu altaris
1KGS|18|33|et composuit ligna divisitque per membra bovem et posuit super ligna
1KGS|18|34|et ait: " Implete quattuor hydrias aqua et fundite super holocaustum et super ligna ". Rursumque dixit: " Etiam secundo hoc facite ". Qui cum fecissent et secundo, ait: " Etiam tertio idipsum facite ". Feceruntque et tertio,
1KGS|18|35|et currebant aquae circum altare, et fossa aquaeductus repleta est.
1KGS|18|36|Cumque iam tempus esset, ut offerretur sacrificium, accedens Elias propheta ait: " Domine, Deus Abraham, Isaac et Israel, hodie ostende quia tu es Deus in Israel, et ego servus tuus et iuxta praeceptum tuum feci omnia haec.
1KGS|18|37|Exaudi me, Domine, exaudi me, ut discat populus iste quia tu, Domine, es Deus et tu convertisti cor eorum iterum! ".
1KGS|18|38|Cecidit autem ignis Domini et voravit holocaustum et ligna et lapides, pulverem quoque et aquam, quae erat in aquaeductu lambens.
1KGS|18|39|Quod cum vidisset omnis populus, cecidit in faciem suam et ait: " Dominus ipse est Deus, Dominus ipse est Deus! ".
1KGS|18|40|Dixitque Elias ad eos: " Apprehendite prophetas Baal, et ne unus quidem effugiat ex eis! ". Quos cum comprehendissent, duxit eos Elias ad torrentem Cison et interfecit eos ibi.
1KGS|18|41|Et ait Elias ad Achab: " Ascende, comede et bibe, quia sonus multae pluviae est ".
1KGS|18|42|Ascendit Achab, ut comederet et biberet. Elias autem ascendit in verticem Carmeli et pronus in terram posuit faciem inter genua sua
1KGS|18|43|et dixit ad puerum suum: " Ascende et prospice contra mare ". Qui, cum ascen disset et contemplatus esset, ait: " Non est quidquam ". Et rursum ait illi: " Revertere septem vicibus ".
1KGS|18|44|In septima autem vice dixit: " Ecce nubecula parva quasi manus hominis ascendit de mari ". Et ait: " Ascende et dic Achab: Iunge et descende, ne occupet te pluvia! ".
1KGS|18|45|Et factum est interea: ecce caeli contenebrati sunt, et nubes et ventus, et facta est pluvia grandis. Ascendens itaque Achab abiit in Iezrahel.
1KGS|18|46|Et manus Domini facta est super Eliam; accinctisque lumbis, currebat ante Achab, donec veniret in Iezrahel.
1KGS|19|1|Nuntiavit autem Achab Iezabel omnia, quae fecerat Elias, et quomodo occidisset universos prophetas gladio.
1KGS|19|2|Misitque Iezabel nuntium ad Eliam dicens: " Haec mihi faciant dii et haec addant, nisi hac hora cras posuero animam tuam sicut animam unius ex illis ".
1KGS|19|3|Timuit ergo Elias et surgens abiit, ut animam suam salvaret, venitque in Bersabee Iudae et dimisit ibi puerum suum.
1KGS|19|4|Et perrexit in desertum via unius diei; cumque venisset et sederet subter unam iuniperum, petivit animae suae, ut moreretur, et ait: " Sufficit mihi, Domine! Tolle animam meam; neque enim melior sum quam patres mei ".
1KGS|19|5|Proiecitque se et obdormivit in umbra iuniperi; et ecce angelus tetigit eum et dixit illi: " Surge, comede! ".
1KGS|19|6|Respexit, et ecce ad caput suum subcinericius panis et vas aquae; comedit ergo et bibit et rursum obdormivit.
1KGS|19|7|Reversusque est angelus Domini secundo et tetigit eum dixitque illi: " Surge, comede! Grandis enim tibi restat via ".
1KGS|19|8|Qui, cum surrexisset, comedit et bibit et ambulavit in fortitudine cibi illius quadraginta diebus et quadraginta noctibus usque ad montem Dei Horeb.
1KGS|19|9|Cumque venisset illuc, mansit in spelunca. Et ecce sermo Domini ad eum dixitque illi: " Quid hic agis, Elia? ".
1KGS|19|10|At ille respondit: " Zelo zelatus sum pro Domino, Deo exercituum, quia dereliquerunt pactum tuum filii Israel, altaria tua destruxerunt et prophetas tuos occiderunt gladio; et derelictus sum ego solus, et quaerunt animam meam, ut auferant eam ".
1KGS|19|11|Et ait ei: " Egredere et sta in monte coram Domino ". Et ecce Dominus transit, et ventus grandis et fortis subvertens montes et conterens petras ante Dominum; non in vento Dominus. Et post ventum, commotio; non in commotione Dominus.
1KGS|19|12|Et post commotionem, ignis; non in igne Dominus. Et post ignem, sibilus aurae tenuis.
1KGS|19|13|Quod cum audisset Elias, operuit vultum suum pallio et egressus stetit in ostio speluncae; et ecce vox ad eum dicens: " Quid agis hic, Elia? ".
1KGS|19|14|Et ille respondit: " Zelo zelatus sum pro Domino, Deo exercituum, quia dereliquerunt pactum tuum filii Israel, altaria tua destruxerunt et prophetas tuos occiderunt gladio; et derelictus sum ego solus, et quaerunt animam meam, ut auferant eam ".
1KGS|19|15|Et ait Dominus ad eum: " Vade et revertere in viam tuam per desertum in Damascum. Cumque perveneris, unges Hazael regem super Syriam;
1KGS|19|16|et Iehu filium Namsi unges regem super Israel; Eliseum autem filium Saphat, qui est de Abelmehula, unges prophetam pro te.
1KGS|19|17|Et erit: quicumque fugerit gladium Hazael, occidet eum Iehu; et, qui fugerit gladium Iehu, interficiet eum Eliseus.
1KGS|19|18|Et relinquam mihi in Israel septem milia: universorum genua, quae non sunt incurvata ante Baal, et omne os, quod non osculatum est eum ".
1KGS|19|19|Profectus ergo inde repperit Eliseum filium Saphat arantem duodecim iugis boum; et ipse cum duodecimo erat. Cumque venisset Elias ad eum, misit pallium suum super illum,
1KGS|19|20|qui statim, relictis bobus, cucurrit post Eliam et ait: " Osculer, oro, patrem meum et matrem meam, et sic sequar te ". Dixitque ei: " Vade et revertere; quid enim feci tibi? ".
1KGS|19|21|Reversus autem ab eo tulit par boum et mactavit illud et in iugo boum coxit carnes et dedit populo, et comederunt. Consurgensque abiit et secutus est Eliam et ministrabat ei.
1KGS|20|1|Porro Benadad rex Syriae congregavit omnem exerci tum suum et triginta duos reges secum et equos et currus et ascendens pugnabat contra Samariam et obsidebat eam.
1KGS|20|2|Mittensque nuntios ad Achab regem Israel in civitatem
1KGS|20|3|ait: " Haec dicit Benadad: Argentum tuum et aurum tuum meum est, et uxores tuae et filii tui optimi mei sunt ".
1KGS|20|4|Responditque rex Israel: " Iuxta verbum tuum, domine mi rex; tuus sum ego et omnia mea ".
1KGS|20|5|Revertentesque nuntii dixerunt: " Haec dicit Benadad: Quia misi ad te dicens: "Argentum tuum et aurum tuum et uxores tuas et filios tuos dabis mihi",
1KGS|20|6|profecto cras hac eadem hora mittam servos meos ad te, et scrutabuntur domum tuam et domum servorum tuorum; et omne, quod oculis tuis pretiosum est, ponent in manibus suis et auferent ".
1KGS|20|7|Vocavit autem rex Israel omnes seniores terrae et ait: " Animadvertite et videte quoniam insidietur nobis; misit enim ad me pro uxoribus meis et filiis et pro argento et auro, et non abnui ".
1KGS|20|8|Dixeruntque omnes maiores natu et universus populus ad eum: " Non audias neque acquiescas illi ".
1KGS|20|9|Respondit itaque nuntiis Benadad: " Dicite domino meo regi: Omnia, propter quae misisti ad me servum tuum initio, faciam; hanc autem rem facere non possum ". Reversique nuntii rettulerunt ei.
1KGS|20|10|Qui remisit et ait: " Haec faciant mihi dii et haec addant, si suffecerit pulvis Samariae pugillis omnis populi, qui sequitur me ".
1KGS|20|11|Et respondens rex Israel ait: " Dicite ei: Ne glorietur accinctus aeque ut discinctus ".
1KGS|20|12|Factum est autem, cum audisset verbum istud, bibebat ipse et reges in umbraculis et ait servis suis: " Circumdate civitatem! ". Et circumdederunt eam.
1KGS|20|13|Et ecce propheta unus accedens ad Achab regem Israel ait: " Haec dicit Dominus: Certe vidisti omnem multitudinem hanc nimiam. Ecce ego tradam eam in manu tua hodie, ut scias quia ego sum Dominus ".
1KGS|20|14|Et ait Achab: " Per quem? ". Dixitque ei: " Haec dicit Dominus: Per pedisequos principum provinciarum ". Et ait: " Quis incipiet proeliari? ". Et ille dixit: " Tu ".
1KGS|20|15|Recensuit ergo pueros principum provinciarum et repperit numerum ducentorum triginta duorum; et post eos recensuit populum, omnes filios Israel, septem milia.
1KGS|20|16|Et egressi sunt meridie. Benadad autem bibebat temulentus in umbraculis ipse et reges triginta duo cum eo, qui ad auxilium eius venerant.
1KGS|20|17|Egressi sunt autem pueri principum provinciarum in prima fronte. Misit itaque Benadad, qui nuntiaverunt ei dicentes: " Viri egressi sunt de Samaria ".
1KGS|20|18|At ille ait: " Sive pro pace veniunt, apprehendite eos vivos; sive ut proelientur, vivos eos capite ".
1KGS|20|19|Egressi erant ergo ex urbe pueri principum provinciarum, ac reliquus exercitus sequebatur,
1KGS|20|20|et percussit unusquisque virum, qui contra se venerat; fugeruntque Syri, et persecutus est eos Israel. Fugit quoque Benadad rex Syriae in equo cum equitibus.
1KGS|20|21|Necnon egressus rex Israel percussit equos et currus et percussit Syriam plaga magna.
1KGS|20|22|Accedens autem propheta ad regem Israel dixit ei: " Vade et confortare et scito et vide quid facias; vertente enim anno rex Syriae ascendet contra te ".
1KGS|20|23|Servi vero regis Syriae dixerunt ei: " Deus montium est Deus eorum, ideo superaverunt nos; sed pugnemus contra eos in campestribus et obtinebimus eos.
1KGS|20|24|Fac ergo hoc: Amove reges singulos a loco suo et pone principes pro eis;
1KGS|20|25|et instaura numerum militum, qui ceciderunt de tuis, et equos secundum equos pristinos et currus secundum currus, quos ante habuisti, et pugnabimus contra eos in campestribus: et videbis quod obtinebimus eos ". Credidit consilio eorum et fecit ita.
1KGS|20|26|Igitur vertente anno recensuit Benadad Syros et ascendit in Aphec, ut pugnaret contra Israel.
1KGS|20|27|Porro filii Israel recensiti sunt et, acceptis cibariis, profecti ex adverso castraque metati sunt contra eos, quasi duo parvi greges caprarum; Syri autem repleverunt terram.
1KGS|20|28|Et accedens vir Dei dixit ad regem Israel: " Haec dicit Dominus: Quia dixerunt Syri: "Deus montium est Dominus et non est Deus vallium", dabo omnem multitudinem hanc grandem in manu tua, et scietis quia ego Dominus.
1KGS|20|29|Dirigebant septem diebus ex adverso hi atque illi acies, septima autem die commissum est bellum; percusseruntque filii Israel de Syris centum milia peditum in die una.
1KGS|20|30|Fugerunt autem, qui remanserant in Aphec, in civitatem, et cecidit murus super viginti septem milia hominum, qui remanserant.Porro Benadad fugiens ingressus est civitatem in cubiculum, quod erat intra cubiculum.
1KGS|20|31|Dixeruntque ei servi sui: " Ecce audivimus quod reges domus Israel clementes sint; ponamus itaque saccos in lumbis nostris et funiculos in capitibus nostris et egrediamur ad regem Israel; forsitan salvabit animam tuam ".
1KGS|20|32|Accinxerunt saccis lumbos suos et posuerunt funes in capitibus suis veneruntque ad regem Israel et dixerunt: " Servus tuus Benadad dicit: Vivat, oro te, anima mea" ". Et ille ait: " Si adhuc vivit, frater meus est ".
1KGS|20|33|Quod acceperunt viri pro omine et festinantes rapuerunt verbum ex ore eius atque dixerunt: " Frater tuus Benadad ". Et dixit eis: " Ite et adducite eum ". Egressus est ergo ad eum Benadad, et levavit eum in currum suum.
1KGS|20|34|Qui dixit ei: " Civitates, quas tulit pater meus a patre tuo, reddam; et plateas fac tibi in Damasco, sicut fecit pater meus in Samaria ". Achab: " Ego autem, inquit, foederatum te dimittam ". Et pepigit ei foedus et dimisit eum.
1KGS|20|35|Tunc vir quidam de filiis prophetarum dixit ad socium suum in sermone Domini: " Percute me! ". At ille noluit percutere.
1KGS|20|36|Cui ait: " Quia noluisti audire vocem Domini, ecce recedes a me, et percutiet te leo ". Cumque paululum recessisset ab eo, invenit eum leo atque percussit.
1KGS|20|37|Sed et alterum inveniens virum dixit ad eum: " Percute me! ". Qui percussit eum et vulneravit.
1KGS|20|38|Abiit ergo propheta et occurrit regi in via et mutavit aspectum ponens fasciam super oculos suos.
1KGS|20|39|Cumque rex transiret, clamavit ad regem et ait: " Servus tuus egressus est ad proeliandum comminus; cumque fugisset vir unus, adduxit eum quidam ad me et ait: "Custodi virum istum! Qui si lapsus fuerit, erit anima tua pro anima eius, aut talentum argenti appendes".
1KGS|20|40|Dum autem ego turbatus huc illucque me verterem, subito non comparuit. Et ait rex Israel ad eum: " Hoc est iudicium tuum, quod ipse decrevisti.
1KGS|20|41|At ille statim abstulit fasciam de oculis suis, et cognovit eum rex Israel quod esset de prophetis.
1KGS|20|42|Qui ait ad eum: " Haec dicit Dominus: Quia dimisisti de manu tua virum, quem morti devoveram, erit anima tua pro anima eius, et populus tuus pro populo eius ".
1KGS|20|43|Reversus est igitur rex Israel in domum suam tristis et indignans venitque in Samariam.
1KGS|21|1|Postea autem factum est hoc. Vinea erat Naboth Iez rahelitae, quae erat in Iezrahel iuxta palatium Achab regis Samariae.
1KGS|21|2|Locutus est ergo Achab ad Naboth dicens: " Da mihi vineam tuam, ut faciam mihi hortum holerum, quia vicina est et prope domum meam. Daboque tibi pro ea vineam meliorem aut, si tibi commodius putas, argenti pretium quanto digna est ".
1KGS|21|3|Cui respondit Naboth: " Propitius mihi sit Dominus, ne dem hereditatem patrum meorum tibi ".
1KGS|21|4|Venit ergo Achab in domum suam tristis et indignans super verbo, quod locutus fuerat ad eum Naboth Iezrahelites dicens: " Non dabo tibi hereditatem patrum meorum ". Et proiciens se in lectulum suum avertit faciem ad parietem et non comedit panem.
1KGS|21|5|Ingressa est autem ad eum Iezabel uxor sua dixitque ei: " Quid est hoc, unde anima tua contristata est? Et quare non comedis panem? ".
1KGS|21|6|Qui respondit ei: " Quia locutus sum Naboth Iezrahelitae et dixi ei: Da mihi vineam tuam, accepta pecunia; aut, si tibi placet, dabo tibi vineam pro ea. Et ille ait: "Non dabo tibi vineam meam" ".
1KGS|21|7|Dixit ergo ad eum Iezabel uxor eius: " Grandis auctoritatis es et bene regis regnum Israel! Surge et comede panem et aequo esto animo; ego dabo tibi vineam Naboth Iezrahelitae ".
1KGS|21|8|Scripsit itaque litteras ex nomine Achab et signavit eas anulo eius et misit ad maiores natu et ad optimates, qui erant in civitate eius et habitabant cum Naboth.
1KGS|21|9|Litterarum autem haec erat sententia: " Praedicate ieiunium et sedere facite Naboth in capite populi
1KGS|21|10|et submittite duos viros filios Belial contra eum, et testimonium dicant: "Maledixisti Deum et regem"; et educite eum et lapidate, sicque moriatur ".
1KGS|21|11|Fecerunt ergo cives eius maiores natu et optimates, qui habitabant cum eo in urbe, sicut praeceperat eis Iezabel et sicut scriptum erat in litteris, quas miserat ad eos.
1KGS|21|12|Praedicaverunt ieiunium et sedere fecerunt Naboth in capite populi;
1KGS|21|13|et ingressi duo viri filii Belial sederunt contra eum et illi, ut viri diabolici, dixerunt contra eum testimonium coram multitudine: " Maledixit Naboth Deum et regem ". Quam ob rem eduxerunt eum extra civitatem et lapidibus interfecerunt;
1KGS|21|14|miseruntque ad Iezabel dicentes: " Lapidatus est Naboth et mortuus est.
1KGS|21|15|Factum est autem cum audisset Iezabel lapidatum Naboth et mortuum, locuta est ad Achab: " Surge, posside vineam Naboth Iezrahelitae, qui noluit tibi acquiescere et dare eam, accepta pecunia; non enim vivit Naboth, sed mortuus est ".
1KGS|21|16|Quod cum audisset Achab, mortuum videlicet Naboth, surrexit et descendebat in vineam Naboth Iezrahelitae, ut possideret eam.
1KGS|21|17|Factus est igitur sermo Domini ad Eliam Thesbiten dicens:
1KGS|21|18|" Surge et descende in occursum Achab regis Israel, qui est in Samaria; ecce est in vinea Naboth, ad quam descendit, ut possideat eam.
1KGS|21|19|Et loqueris ad eum dicens: Haec dicit Dominus: Occidisti, insuper et possedisti! Et post haec addes: Haec dicit Dominus: In loco, in quo linxerunt canes sanguinem Naboth, lambent tuum quoque sanguinem ".
1KGS|21|20|Et ait Achab ad Eliam: " Num invenisti me, inimice mi? ". Qui dixit: " Inveni, eo quod venumdatus sis, ut faceres malum in conspectu Domini.
1KGS|21|21|Ecce ego inducam super te malum et demetam posteriora tua et interficiam de Achab quidquid masculini sexus sive impuberem sive puberem in Israel.
1KGS|21|22|Et dabo domum tuam sicut domum Ieroboam filii Nabat et sicut domum Baasa filii Ahia, quia egisti, ut me ad iracundiam provocares, et peccare fecisti Israel.
1KGS|21|23|Sed et de Iezabel locutus est Dominus dicens: Canes comedent Iezabel in agro Iezrahel.
1KGS|21|24|Qui de Achab mortuus fuerit in civitate, comedent eum canes; qui autem mortuus fuerit in agro, comedent eum volucres caeli ".
1KGS|21|25|Igitur non fuit alter talis sicut Achab, qui venumdatus est, ut faceret malum in conspectu Domini; concitavit enim eum Iezabel uxor sua,
1KGS|21|26|et abominabilis effectus est, in tantum ut sequeretur idola secundum omnia, quae fecerant Amorraei, quos consumpsit Dominus a facie filiorum Israel.
1KGS|21|27|Itaque cum audisset Achab sermones istos, scidit vestem suam et operuit cilicio carnem suam ieiunavitque et dormivit in sacco et ambulabat demisso capite.
1KGS|21|28|Factus est autem sermo Domini ad Eliam Thesbiten dicens:
1KGS|21|29|Nonne vidisti humiliatum Achab coram me? Quia igitur humiliatus est mei causa, non inducam malum in diebus eius, sed in diebus filii sui inferam malum domui eius ".
1KGS|22|1|Transierunt igitur tres anni absque bello inter Syriam et Israel.
1KGS|22|2|In anno autem tertio descendit Iosaphat rex ludae ad regem Israel,
1KGS|22|3|dixitque rex Israel ad servos suos: " Ignoratis quod nostra sit Ramoth Galaad et neglegimus tollere eam de manu regis Syriae? ".
1KGS|22|4|Et ait ad Iosaphat: " Veniesne mecum ad proeliandum in Ramoth Galaad? ".
1KGS|22|5|Dixitque Iosaphat ad regem Israel: " Sicut ego sum, ita et tu; populus meus et populus tuus unum sunt, et equites mei et equites tui ". Dixitque Iosaphat ad regem Israel: " Quaere, oro te, hodie sermonem Domini ".
1KGS|22|6|Congregavit ergo rex Israel prophetas quadringentos circiter viros et ait ad eos: " Ire debeo in Ramoth Galaad ad bellandum, an quiescere? ". Qui responderunt: " Ascende, et dabit Dominus in manu regis ".
1KGS|22|7|Dixit autem Iosaphat: " Non est hic et alius propheta Domini, ut interrogemus per eum? ".
1KGS|22|8|Et ait rex Israel ad Iosaphat: " Remansit vir unus, per quem possimus interrogare Dominum; sed ego odi eum, quia non prophetat mihi bonum sed malum: Michaeas filius Iemla ". Cui Iosaphat ait: " Ne loquaris ita, rex.
1KGS|22|9|Vocavit ergo rex Israel eunuchum quendam et dixit ei: " Festina adducere Michaeam filium Iemla ".
1KGS|22|10|Rex autem Israel et Iosaphat rex Iudae sedebat unusquisque in solio suo vestiti cultu regio in area iuxta ostium portae Samariae; et universi prophetae prophetabant in conspectu eorum.
1KGS|22|11|Fecit quoque sibi Sedecias filius Chanaana cornua ferrea et ait: " Haec dicit Dominus: His ventilabis Syriam, donec deleas eam ".
1KGS|22|12|Omnesque prophetae similiter prophetabant dicentes: " Ascende in Ramoth Galaad et vade prospere, et tradet Dominus in manu regis ".
1KGS|22|13|Nuntius vero, qui ierat ut vocaret Michaeam, locutus est ad eum dicens: Ecce sermones prophetarum ore uno regi bona praedicant; sit ergo sermo tuus similis eorum, et loquere bona ".
1KGS|22|14|Cui Michaeas ait: " Vivit Dominus quia, quodcumque dixerit mihi Dominus, hoc loquar! ".
1KGS|22|15|Venit itaque ad regem, et ait illi rex: " Michaea, ire debemus in Ramoth Galaad ad proeliandum, an cessare? ". Cui ille respondit: " Ascende et vade prospere, et tradet Dominus in manu regis ".
1KGS|22|16|Dixit autem rex ad eum: " Iterum atque iterum adiuro te, ut non loquaris mihi, nisi quod verum est in nomine Domini ".
1KGS|22|17|Et ille ait: Vidi cunctum Israeldispersum in montibusquasi oves non habentes pastorem. Et ait Dominus: "Non habent isti dominum; revertatur unusquisque in domum suam in pace" ".
1KGS|22|18|Dixit ergo rex Israel ad Iosaphat: " Numquid non dixi tibi quia non prophetat mihi bonum sed semper malum? ".
1KGS|22|19|Ille vero addens ait: " Propterea audi sermonem Domini: Vidi Dominum sedentem super solium suum et omnem exercitum caeli assistentem ei a dextris et a sinistris.
1KGS|22|20|Et ait Dominus: "Quis decipiet Achab, ut ascendat et cadat in Ramoth Galaad?". Et dixit unus verba huiuscemodi et alius aliter.
1KGS|22|21|Egressus est autem spiritus et stetit coram Domino et ait: "Ego decipiam illum". Cui locutus est Dominus: "In quo?".
1KGS|22|22|Et ille ait: "Egrediar et ero spiritus mendax in ore omnium prophetarum eius". Et dixit Dominus: "Decipies et praevalebis; egredere et fac ita".
1KGS|22|23|Nunc igitur ecce dedit Dominus spiritum mendacii in ore omnium prophetarum tuorum, qui hic sunt, et Dominus locutus est contra te malum.
1KGS|22|24|Accessit autem Sedecias filius Chanaana et percussit Michaeam in maxillam et dixit: " Quomodo transivit spiritus Domini a me, ut loqueretur tibi? ".
1KGS|22|25|Et ait Michaeas: " Visurus es in die illa, quando ingredieris cubiculum intra cubiculum, ut abscondaris ".
1KGS|22|26|Et ait rex Israel: " Tolle Michaeam, et maneat apud Amon principem civitatis et apud Ioas filium regis,
1KGS|22|27|et dic eis: "Haec dicit rex: Mittite virum istum in carcerem et sustentate eum pane tribulationis et aqua angustiae, donec revertar in pace" ".
1KGS|22|28|Dixitque Michaeas: " Si reversus fueris in pace, non est locutus Dominus in me ". Et ait: " Audite, populi omnes! ".
1KGS|22|29|Ascendit itaque rex Israel et Iosaphat rex Iudae in Ramoth Galaad.
1KGS|22|30|Dixitque rex Israel ad Iosaphat: " Mutato aspectu ineundum est proelium; tu autem induere vestibus tuis ". Porro rex Israel mutavit aspectum et ingressus est bellum.
1KGS|22|31|Rex autem Syriae praeceperat principibus curruum triginta duobus dicens: " Non pugnabitis contra minorem et maiorem quempiam, nisi contra regem Israel solum ".
1KGS|22|32|Cum ergo vidissent principes curruum Iosaphat, suspicati sunt quod ipse esset rex Israel et impetu facto pugnabant contra eum. Et exclamavit Iosaphat;
1KGS|22|33|intellexeruntque principes curruum quod non esset rex Israel et cessaverunt ab eo.
1KGS|22|34|Vir autem quidam tetendit arcum in incertum sagittam dirigens et percussit regem Israel inter iuncturas et loricam. At ille dixit aurigae suo: " Verte manum tuam et eice me de exercitu, quia graviter vulneratus sum ".
1KGS|22|35|Aggravatum est ergo proelium in die illa; et rex Israel stabat in curru suo contra Syros et mortuus est vespere: fluebat autem sanguis plagae in sinum currus.
1KGS|22|36|Et clamor insonuit in universo exercitu ad solis occasum: " Unusquisque revertatur in civitatem et in terram suam! ".
1KGS|22|37|Mortuus est igitur rex et perlatus est Samariam; sepelieruntque regem in Samaria.
1KGS|22|38|Et laverunt currum eius in piscina Samariae; et linxerunt canes sanguinem eius, et scorta laverunt se iuxta verbum Domini, quod locutus fuerat.
1KGS|22|39|Reliqua vero gestorum Achab et universa, quae fecit, et domus eburnea, quam aedificavit, cunctaeque urbes, quas exstruxit, nonne haec scripta sunt in libro annalium regum Israel?
1KGS|22|40|Dormivit ergo Achab cum patribus suis; et regnavit Ochozias filius eius pro eo.
1KGS|22|41|Iosaphat vero filius Asa regnare coeperat super Iudam anno quarto Achab regis Israel;
1KGS|22|42|triginta quinque annorum erat, cum regnare coepisset, et viginti quinque annos regnavit in Ierusalem. Nomen matris eius Azuba filia Selachi.
1KGS|22|43|Et ambulavit in omni via Asa patris sui et non declinavit ex ea; fecitque, quod rectum erat in conspectu Domini.
1KGS|22|44|Verumtamen excelsa non abstulit; adhuc enim populus sacrificabat et adolebat in excelsis.
1KGS|22|45|Pacemque fecit Iosaphat cum rege Israel.
1KGS|22|46|Reliqua autem gestorum Iosaphat et opera eius, quae fortiter gessit, et proelia, nonne haec scripta sunt in libro annalium regum Iudae?
1KGS|22|47|Sed et reliquias prostibulorum, qui remanserant in diebus Asa patris eius, abstulit de terra.
1KGS|22|48|Nec erat tunc rex in Edom sed praefectus regius.
1KGS|22|49|Rex vero Iosaphat fecerat naves Tharsis, quae navigarent in Ophir propter aurum; et ire non potuerunt, quia confractae sunt in Asiongaber.
1KGS|22|50|Tunc ait Ochozias filius Achab ad Iosaphat: " Vadant servi mei cum servis tuis in navibus ". Et noluit Iosaphat.
1KGS|22|51|Dormivitque Iosaphat cum patribus suis et sepultus est cum eis in civitate David patris sui; regnavitque Ioram filius eius pro eo.
1KGS|22|52|Ochozias autem filius Achab regnare coeperat super Israel in Samaria anno septimo decimo Iosaphat regis Iudae regnavitque super Israel duobus annis.
1KGS|22|53|Et fecit malum in conspectu Domini et ambulavit in via patris sui et matris suae et in via Ieroboam filii Nabat, qui peccare fecit Israel;
1KGS|22|54|servivit quoque Baal et adoravit eum et irritavit Dominum, Deum Israel, iuxta omnia, quae fecerat pater eius.
2KGS|1|1|Praevaricatus est autem Moab in Israel, postquam mortuus est Achab.
2KGS|1|2|Ceciditque Ochozias per cancellos cenaculi sui, quod habebat in Samaria, et aegrotavit; misitque nuntios dicens ad eos: " Ite, consulite Beelzebub deum Accaron, utrum vivere queam de infirmitate mea hac ".
2KGS|1|3|Angelus autem Domini locutus est ad Eliam Thesbiten: " Surge, ascende in occursum nuntiorum regis Samariae et dices ad eos: Numquid non est Deus in Israel, ut eatis ad consulendum Beelzebub deum Accaron?
2KGS|1|4|Quam ob rem haec dicit Dominus: De lectulo, super quem ascendisti, non descendes, sed morte morieris ". Et abiit Elias.
2KGS|1|5|Reversique sunt nuntii ad Ochoziam, qui dixit eis: " Quare reversi estis? ".
2KGS|1|6|At illi responderunt ei: " Vir occurrit nobis et dixit ad nos: "Ite, revertimini ad regem, qui misit vos, et dicetis ei: Haec dicit Dominus: Numquid, quia non est Deus in Israel, mittis, ut consulatur Beelzebub deus Accaron? Idcirco de lectulo, super quem ascendisti, non descendes, sed morte morieris" ".
2KGS|1|7|Qui dixit eis: " Cuius figurae et habitus vir erat, qui occurrit vobis et locutus est verba haec? ".
2KGS|1|8|At illi dixerunt: " Vir in veste pilosa et zona pellicea accinctis renibus ". Qui ait: " Elias Thesbites est ".
2KGS|1|9|Misitque ad eum quinquagenarium principem et quinquaginta, qui erant sub eo; qui ascendit ad eum sedentique in vertice montis ait: " Homo Dei, rex praecepit, ut descendas ".
2KGS|1|10|Respondensque Elias dixit quinquagenario: " Si homo Dei sum, descendat ignis e caelo et devoret te et quinquaginta tuos ". Descendit itaque ignis e caelo et devoravit eum et quinquaginta, qui erant cum eo.
2KGS|1|11|Rursum misit ad eum principem quinquagenarium alterum et quinquaginta cum eo; qui locutus est illi: " Homo Dei, haec dicit rex: "Festina, descende!" ".
2KGS|1|12|Respondens Elias ait illis: " Si homo Dei ego sum, descendat ignis e caelo et devoret te et quinquaginta tuos ". Descendit ergo ignis Dei e caelo et devoravit illum et quinquaginta eius.
2KGS|1|13|Iterum misit principem quinquagenarium tertium et quinquaginta, qui erant cum eo; qui cum venisset, curvavit genua contra Eliam et precatus est eum et ait: " Homo Dei, noli despicere animam meam et animam servorum tuorum, qui mecum sunt.
2KGS|1|14|Ecce descendit ignis de caelo et devoravit duos principes quinquagenarios primos et quinquagenos, qui cum eis erant; sed nunc obsecro, ut miserearis animae meae ".
2KGS|1|15|Locutus est autem angelus Domini ad Eliam dicens: " Descende cum eo, ne timeas ". Surrexit igitur et descendit cum eo ad regem
2KGS|1|16|et locutus est ei: " Haec dicit Dominus: Quia misisti nuntios ad consulendum Beelzebub deum Accaron, quasi non esset Deus in Israel, a quo posses interrogare sermonem, ideo de lectulo, super quem ascendisti, non descendes, sed morte morieris ".
2KGS|1|17|Mortuus est ergo iuxta sermonem Domini, quem locutus est Elias. Et regnavit Ioram frater eius pro eo anno secundo Ioram filii Iosaphat regis Iudae; non enim habebat filium.
2KGS|1|18|Reliqua autem gestorum Ochoziae, quae operatus est, nonne haec scripta sunt in libro annalium regum Israel?
2KGS|2|1|Factum est autem cum levare vellet Dominus Eliam per turbi nem in caelum, ibant Elias et Eliseus de Galgalis;
2KGS|2|2|dixitque Elias ad Eliseum: " Sede hic, quia Dominus misit me usque Bethel ". Cui ait Eliseus: " Vivit Dominus, et vivit anima tua, quia non derelinquam te ". Cumque descendissent Bethel,
2KGS|2|3|egressi sunt filii prophetarum, qui erant in Bethel, ad Eliseum et dixerunt ei: "Numquid nosti quia hodie Dominus tollat dominum tuum desuper capite tuo? ". Qui respondit: " Et ego novi, silete ".
2KGS|2|4|Dixit autem ei Elias: " Elisee, sede hic, quia Dominus misit me in Iericho ". Et ille ait: " Vivit Dominus, et vivit anima tua, quia non derelinquam te ". Cumque venissent Ierichum,
2KGS|2|5|accesserunt filii prophetarum, qui erant in Iericho, ad Eliseum et dixerunt ei: " Numquid nosti quia hodie Dominus tollet dominum tuum desuper capite tuo? ". Et ait: " Et ego novi, silete ".
2KGS|2|6|Dixit autem ei Elias: " Sede hic, quia Dominus misit me ad Iordanem ". Qui ait: " Vivit Dominus, et vivit anima tua, quia non derelinquam te ". Ierunt igitur ambo pariter,
2KGS|2|7|et quinquaginta viri de filiis prophetarum secuti sunt, qui et steterunt e contra longe. Illi autem ambo stabant super Iordanem.
2KGS|2|8|Tulitque Elias pallium suum et involvit illud et percussit aquas, quae divisae sunt in utramque partem, et transierunt ambo per siccum.
2KGS|2|9|Cumque transissent, Elias dixit ad Eliseum: " Postula, quod vis, ut faciam tibi, antequam tollar a te ". Dixitque Eliseus: " Obsecro, ut fiant duae partes spiritus tui in me ".
2KGS|2|10|Qui respondit: " Rem difficilem postulasti. Attamen si videris me, quando tollor a te, erit tibi, quod petisti; si autem non videris, non erit ".
2KGS|2|11|Cumque pergerent et incedentes sermocinarentur, ecce currus igneus et equi ignei diviserunt utrumque; et ascendit Elias per turbinem in caelum.
2KGS|2|12|Eliseus autem videbat et clamabat: " Pater mi, pater mi, currus Israel et auriga eius! ". Et non vidit eum amplius; apprehenditque vestimenta sua et scidit illa in duas partes.
2KGS|2|13|Et levavit pallium Eliae, quod ceciderat ei, reversusque stetit super ripam Iordanis.
2KGS|2|14|Et pallio Eliae, quod ceciderat ei, percussit aquas et dixit: " Ubi est Deus Eliae etiam nunc? ". Percussitque aquas, et divisae sunt huc atque illuc, et transiit Eliseus.
2KGS|2|15|Videntes autem filii prophetarum, qui erant in Iericho de contra, dixerunt: " Requievit spiritus Eliae super Eliseum ". Et venientes in occursum eius adoraverunt eum proni in terram
2KGS|2|16|dixeruntque illi: " Ecce cum servis tuis sunt quinquaginta viri fortes, qui possunt ire et quaerere dominum tuum, ne forte tulerit eum spiritus Domini et proiecerit in uno montium aut in una vallium ". Qui ait: " Nolite mittere! ".
2KGS|2|17|Coegeruntque eum, donec acquiesceret et diceret: " Mittite ". Et miserunt quinquaginta viros. Qui cum quaesissent tribus diebus, non invenerunt
2KGS|2|18|et reversi sunt ad eum. At ille habitabat in Iericho dixitque eis: " Numquid non dixi vobis: Nolite ire?".
2KGS|2|19|Dixerunt quoque viri civitatis ad Eliseum: " Ecce habitatio civitatis huius optima est, sicut tu ipse, domine, perspicis; sed aquae pessimae sunt, et terra faciens abortium ".
2KGS|2|20|At ille ait: "Afferte mihi vas novum et mittite in illud sal ". Qui cum attulissent,
2KGS|2|21|egressus ad fontem aquarum misit in eum sal et ait: " Haec dicit Dominus: Sanavi aquas has, et non erit ultra in eis mors neque abortium ".
2KGS|2|22|Sanatae sunt ergo aquae usque ad diem hanc iuxta verbum Elisei, quod locutus est.
2KGS|2|23|Ascendit autem inde Bethel. Cumque ascenderet per viam, pueri parvi egressi sunt de civitate et illudebant ei dicentes: "Ascende, calve; ascende, calve! ".
2KGS|2|24|Qui cum respexisset, vidit eos et maledixit eis in nomine Domini; egressique sunt duo ursi de saltu et laceraverunt ex eis quadraginta duos pueros.
2KGS|2|25|Abiit autem inde in montem Carmeli et inde reversus est Samariam.
2KGS|3|1|Ioram vero filius Achab regnavit super Israel in Samaria anno decimo octavo Iosaphat regis Iudae regnavitque duodecim annis.
2KGS|3|2|Et fecit malum coram Domino, sed non sicut pater suus et mater; tulit enim lapidem Baal, quem fecerat pater eius.
2KGS|3|3|Verumtamen in peccatis Ieroboam filii Nabat, qui peccare fecit Israel, adhaesit nec recessit ab eis.
2KGS|3|4|Porro Mesa rex Moab nutriebat pecora multa et solvebat regi Israel centum milia agnorum et lanam centum milium arietum.
2KGS|3|5|Cumque mortuus fuisset Achab, praevaricatus est foedus, quod habebat cum rege Israel.
2KGS|3|6|Egressus est igitur rex Ioram in die illa de Samaria et recensuit universum Israel;
2KGS|3|7|profectusque misit ad Iosaphat regem Iudae dicens: " Rex Moab recessit a me. Vis venire mecum contra Moab ad proelium? ". Qui respondit: " Ascendam. Qui meus est tuus est, populus meus populus tuus, equi mei equi tui ".
2KGS|3|8|Dixitque: " Per quam viam ascendemus? ". At ille respondit: " Per desertum Idumaeae ".
2KGS|3|9|Perrexerunt igitur rex Israel et rex Iudae et rex Edom et circuierunt per viam septem dierum; nec erat aqua exercitui et iumentis, quae sequebantur eos.
2KGS|3|10|Dixitque rex Israel: " Heu! Congregavit nos Dominus tres reges, ut traderet in manu Moab ".
2KGS|3|11|Et ait Iosaphat: " Estne hic propheta Domini, ut interrogemus Dominum per eum? ". Et respondit unus de servis regis Israel: " Est hic Eliseus filius Saphat, qui fundebat aquam super manus Eliae ".
2KGS|3|12|Et ait Iosaphat: " Est apud eum sermo Domini ". Descenditque ad eum rex Israel et Iosaphat et rex Edom.
2KGS|3|13|Dixit autem Eliseus ad regem Israel: " Quid mihi et tibi est? Vade ad prophetas patris tui et ad prophetas matris tuae ". Et ait illi rex Israel: "Non, congregavit enim Dominus tres reges hos, ut traderet eos in manu Moab? ".
2KGS|3|14|Dixit autem Eliseus: " Vivit Dominus exercituum, in cuius conspectu sto, quod si non vultum Iosaphat regis Iudae revererer, ne attendissem quidem te nec respexissem;
2KGS|3|15|nunc autem adducite mihi psaltem ". Cumque caneret psaltes, facta est super eum manus Domini,
2KGS|3|16|et ait: " Haec dicit Dominus: Facite in torrente hoc fossas et fossas.
2KGS|3|17|Haec enim dicit Dominus: Non videbitis ventum neque pluviam, et torrens replebitur aquis; et bibetis vos et pecora et iumenta vestra.
2KGS|3|18|Parumque hoc est in conspectu Domini; insuper tradet etiam Moab in manu vestra,
2KGS|3|19|et percutietis omnem civitatem munitam et omnem urbem electam et universum lignum fructiferum succidetis cunctosque fontes aquarum obturabitis et omnem agrum egregium operietis lapidibus ".
2KGS|3|20|Factum est igitur mane, quando sacrificium offerri solet, et ecce aquae veniebant per viam Edom. Et repleta est terra aquis.
2KGS|3|21|Universi autem Moabitae audientes quod ascendissent reges, ut pugnarent adversum eos, convocaverunt omnes, qui accingi poterant balteo et desuper, et steterunt in terminis.
2KGS|3|22|Primoque mane surgentes et, orto iam sole super aquis, viderunt Moabitae e contra aquas rubras quasi sanguinem
2KGS|3|23|dixeruntque: "Sanguis est gladii! Pugnaverunt reges contra se et caesi sunt mutuo. Nunc perge ad praedam, Moab! ".
2KGS|3|24|Perrexeruntque in castra Israel. Porro consurgens Israel percussit Moab, at illi fugerunt coram eis. Venerunt igitur subsequentes et percutientes Moab.
2KGS|3|25|Et civitates destruxerunt et omnem agrum optimum mittentes singuli lapides repleverunt; et universos fontes aquarum obturaverunt et omnia ligna fructifera succiderunt, ita ut muri tantum Cirhareseth remanerent; et circumdederunt civitatem fundibularii et aggressi sunt.
2KGS|3|26|Quod cum vidisset rex Moab, praevaluisse scilicet hostes, tulit secum septingentos viros educentes gladium, ut irrumperet ad regem Edom; et non potuerunt.
2KGS|3|27|Arripiensque filium suum primogenitum, qui regnaturus erat pro eo, obtulit holocaustum super murum. Et facta est indignatio magna super Israel; statimque recesserunt ab eo et reversi sunt in terram suam.
2KGS|4|1|Mulier autem quaedam de uxoribus filiorum prophetarum clamabat ad Eliseum dicens: " Servus tuus vir meus mortuus est, et tu nosti quia servus tuus fuit timens Dominum; et ecce creditor venit, ut tollat duos filios meos ad serviendum sibi ".
2KGS|4|2|Cui dixit Eliseus: " Quid vis, ut faciam tibi? Dic mihi: Quid habes in domo tua? ". At illa respondit: " Non habeo ancilla tua quidquam in domo mea, nisi vasculum olei ".
2KGS|4|3|Cui ait: " Vade, pete mutuo ab omnibus vicinis tuis vasa vacua non pauca;
2KGS|4|4|et ingredere et claude ostium, cum intrinsecus fueris tu et filii tui, et mitte inde in omnia vasa haec et, cum plena fuerint, tolles ".
2KGS|4|5|Ivit itaque mulier et clausit ostium super se et super filios suos; illi offerebant vasa, et illa infundebat.
2KGS|4|6|Cumque plena fuissent vasa, dixit ad filium suum: " Affer mihi adhuc vas. Et ille respondit: " Non habeo ". Stetitque oleum.
2KGS|4|7|Venit autem illa et indicavit homini Dei. Et ille: " Vade, inquit, vende oleum et redde creditori tuo; tu autem et filii tui vivite de reliquo ".
2KGS|4|8|Facta est autem quaedam dies, et transibat Eliseus per Sunam. Erat autem ibi mulier magna, quae tenuit eum, ut comederet panem. Quotiescumque inde transibat, divertebat ad eam, ut comederet panem.
2KGS|4|9|Quae dixit ad virum suum: " Animadverto quod vir Dei sanctus est iste, qui transit per nos frequenter.
2KGS|4|10|Faciamus ergo cenaculum muratum parvum et ponamus ei in eo lectulum et mensam et sellam et candelabrum, ut, cum venerit ad nos, maneat ibi ".
2KGS|4|11|Facta est ergo dies quaedam, et veniens divertit in cenaculum et requievit ibi.
2KGS|4|12|Dixitque ad Giezi puerum suum: " Voca Sunamitin istam ". Qui cum vocasset eam, et illa stetisset coram eo,
2KGS|4|13|dixit ad puerum: " Loquere ad eam: Ecce sedule in omnibus ministrasti nobis; quid vis, ut faciam tibi? Numquid habes negotium et vis, ut loquar regi sive principi militiae? ". Quae respondit: " In medio populi mei habito ".
2KGS|4|14|Et ait: " Quid ergo vult, ut faciam ei? ". Dixitque Giezi: "Ne quaeras; filium enim non habet, et vir eius senex est ".
2KGS|4|15|Praecepit itaque, ut vocaret eam; quae cum vocata fuisset et stetisset ad ostium,
2KGS|4|16|dixit ad eam: " In tempore isto, in anno altero, amplexaberis filium ". At illa respondit: " Noli, quaeso, domine mi, vir Dei, noli mentiri ancillae tuae ".
2KGS|4|17|Et concepit mulier et peperit filium in tempore isto anni alterius, quo dixerat Eliseus.
2KGS|4|18|Crevit autem puer et, cum esset quaedam dies, et egressus isset ad patrem suum, ad messores,
2KGS|4|19|ait patri suo: " Caput meum, caput meum! ". At ille dixit servo: " Tolle et duc eum ad matrem suam ".
2KGS|4|20|Qui cum tulisset et adduxisset eum ad matrem suam, posuit eum illa super genua sua usque ad meridiem, et mortuus est.
2KGS|4|21|Ascendit autem et collocavit eum super lectulum hominis Dei et clausit ostium; et egressa
2KGS|4|22|vocavit virum suum et ait: "Mitte mecum, obsecro, unum de pueris et asinam, ut excurram usque ad hominem Dei et revertar ".
2KGS|4|23|Qui ait illi: " Quam ob causam vadis ad eum hodie? Non sunt calendae neque sabbatum ". Quae respondit: " Vale ".
2KGS|4|24|Stravitque asinam et praecepit puero: " Mina et propera, ne mihi moram facias in eundo, nisi praecepero tibi ".
2KGS|4|25|Profecta est igitur et venit ad virum Dei in montem Carmeli. Cumque vidisset eam vir Dei de contra, ait ad Giezi puerum suum: " Ecce Sunamitis illa.
2KGS|4|26|Vade cito in occursum eius et dic ei: Rectene agitur circa te et circa virum tuum et circa filium tuum? ". Quae respondit: " Recte ".
2KGS|4|27|Cumque venisset ad virum Dei in monte, apprehendit pedes eius; et accessit Giezi, ut amoveret eam, et ait homo Dei: " Dimitte illam; anima enim eius in amaritudine est, et Dominus celavit me et non indicavit mihi.
2KGS|4|28|Quae dixit illi: " Numquid petivi filium a domino meo? Numquid non dixi tibi: Ne illudas me? ".
2KGS|4|29|Et ille ait ad Giezi: " Accinge lumbos tuos et tolle baculum meum in manu tua et vade. Si occurrerit tibi homo, non salutes eum et, si salutaverit te quispiam, non respondeas illi. Et pones baculum meum super faciem pueri ".
2KGS|4|30|Porro mater pueri ait: " Vivit Dominus, et vivit anima tua, non dimittam te ". Surrexit ergo et secutus est eam.
2KGS|4|31|Giezi autem praecesserat eos et posuerat baculum super faciem pueri, et non erat vox neque sensus reversusque est in occursum eius et nuntiavit ei dicens: " Non evigilavit puer ".
2KGS|4|32|Ingressus est ergo Eliseus domum, et ecce puer mortuus iacebat in lectulo eius;
2KGS|4|33|ingressusque clausit ostium super se et puerum et oravit ad Dominum.
2KGS|4|34|Et ascendit et incubuit super puerum posuitque os suum super os eius et oculos suos super oculos eius et manus suas super manus eius et incurvavit se super eum, et calefacta est caro pueri.
2KGS|4|35|At ille reversus deambulavit in domo semel huc et illuc et ascendit et incubuit super eum, et sternutavit puer septies aperuitque oculos.
2KGS|4|36|Et ille vocavit Giezi et dixit ei: " Voca Sunamitin hanc ". Quae vocata ingressa est ad eum. Qui ait: " Tolle filium tuum ".
2KGS|4|37|Venit illa et corruit ad pedes eius et adoravit super terram; tulitque filium suum et egressa est.
2KGS|4|38|Et Eliseus reversus est in Galgala. Erat autem fames in terra, et filii prophetarum habitabant coram eo. Dixitque puero suo: " Pone ollam grandem et coque pulmentum filiis prophetarum ".
2KGS|4|39|Et egressus est unus in agrum, ut colligeret herbas agrestes; invenitque quasi vitem silvestrem et collegit ex ea colocynthidas agri. Et implevit pallium suum et reversus concidit in ollam pulmenti; nesciebat enim quid esset.
2KGS|4|40|Infuderunt ergo sociis, ut comederent. Cumque gustassent de coctione, exclamaverunt dicentes: " Mors in olla, vir Dei! ". Et non potuerunt comedere.
2KGS|4|41|At ille: " Afferte, inquit, farinam ". Cumque tulissent, misit in ollam et ait: " Infunde turbae, et comedat ". Et non fuit amplius quidquam amaritudinis in olla.
2KGS|4|42|Vir autem quidam venit de Baalsalisa deferens viro Dei panes primitiarum, viginti panes hordeaceos et frumentum novum in pera sua. At ille dixit: " Da populo, ut comedat ".
2KGS|4|43|Responditque ei minister eius: " Quantum est hoc, ut apponam coram centum viris? ". Rursum ille dixit: " Da populo, ut comedat. Haec enim dicit Dominus: "Comedent, et supererit" ".
2KGS|4|44|Posuit itaque coram eis, qui comederunt, et superfuit iuxta verbum Domini.
2KGS|5|1|Naaman princeps militiae regis Syriae erat vir magnus apud dominum suum et honoratus; per illum enim dedit Dominus salutem Syriae. Erat autem vir fortis leprosus.
2KGS|5|2|Porro de Syria egressa fuerat turma et captivam duxerat de terra Israel puellam parvulam, quae erat in obsequio uxoris Naaman.
2KGS|5|3|Quae ait ad dominam suam: " Utinam esset dominus meus ad prophetam, qui est in Samaria! Profecto curaret eum a lepra, quam habet ".
2KGS|5|4|Ingressus est itaque Naaman ad dominum suum et nuntiavit ei dicens: " Sic et sic locuta est puella de terra Israel ".
2KGS|5|5|Dixitque ei rex Syriae: " Vade, et mittam litteras ad regem Israel ". Qui cum profectus esset et tulisset secum decem talenta argenti et sex milia siclorum auri et decem mutatoria vestimentorum,
2KGS|5|6|detulit litteras ad regem Israel in haec verba: " Cum acceperis epistulam hanc, scito quod miserim ad te Naaman servum meum, ut cures eum a lepra sua ".
2KGS|5|7|Cumque legisset rex Israel litteras, scidit vestimenta sua et ait: " Numquid Deus sum, ut occidere possim et vivificare, quia iste mittit ad me, ut curem hominem a lepra sua? Animadvertite et videte quod occasiones quaerat adversum me ".
2KGS|5|8|Quod cum audisset Eliseus vir Dei, scidisse videlicet regem Israel vestimenta sua, misit ad eum dicens: " Quare scidisti vestimenta tua? Veniat ad me et sciat esse prophetam in Israel ".
2KGS|5|9|Venit ergo Naaman cum equis et curribus et stetit ad ostium domus Elisei.
2KGS|5|10|Misitque ad eum Eliseus nuntium dicens: " Vade et lavare septies in Iordane; et recipiet sanitatem caro tua, atque mundaberis ".
2KGS|5|11|Iratus Naaman recedebat dicens: " Putabam quod egrederetur ad me et stans invocaret nomen Domini Dei sui et tangeret manu sua locum leprae et curaret me.
2KGS|5|12|Numquid non meliores sunt Abana et Pharphar, fluvii Damasci, omnibus aquis Israel, ut laver in eis et munder? ". Cum ergo vertisset se et abiret indignans,
2KGS|5|13|accesserunt ad eum servi sui et locuti sunt ei: " Si rem grandem dixisset tibi propheta, certe faceres; quanto magis quia nunc dixit tibi: Lavare et mundaberis!" ".
2KGS|5|14|Descendit et intinxit se in Iordane septies iuxta sermonem viri Dei, et restituta est caro eius sicut caro pueri parvuli, et mundatus est.
2KGS|5|15|Reversusque ad virum Dei cum universo comitatu suo venit et stetit coram eo et ait: " Vere scio quod non sit Deus in universa terra, nisi tantum in Israel! Obsecro itaque, ut accipias benedictionem a servo tuo ".
2KGS|5|16|At ille respondit: " Vivit Dominus, ante quem sto, non accipiam ". Cumque vim faceret, penitus non acquievit.
2KGS|5|17|Dixitque Naaman: " Ut vis. Sed, obsecro, concedatur mihi servo tuo tantum terrae quantum onus duorum burdonum; non enim faciet ultra servus tuus holocaustum aut victimam diis alienis, nisi Domino.
2KGS|5|18|Hoc autem solum ignoscat Dominus servo tuo, quando ingreditur dominus meus templum Remmon, ut adoret ibi, et illo innitente super manum meam, si adoravero in templo Remmon, adorante eo in eodem loco, ut ignoscat mihi Dominus servo tuo pro hac re ".
2KGS|5|19|Qui dixit ei: " Vade in pace ". Abiit ergo ab eo viam modicam.
2KGS|5|20|Dixitque Giezi puer viri Dei: " Pepercit dominus meus Naaman Syro isti, ut non acciperet ab eo, quae attulit; vivit Dominus, curram post eum et accipiam ab eo aliquid ".
2KGS|5|21|Et secutus est Giezi post tergum Naaman. Quem cum vidisset ille currentem ad se, desiluit de curru in occursum eius et ait: " Rectene sunt omnia? ".
2KGS|5|22|Et ille ait: " Recte. Dominus meus misit me dicens: "Modo venerunt ad me duo adulescentes de monte Ephraim ex filiis prophetarum. Da eis talentum argenti et vestes mutatorias duplices" ".
2KGS|5|23|Dixitque Naaman: " Melius est, ut accipias duo talenta ". Et coegit eum ligavitque duo talenta argenti in duobus saccis et duplicia vestimenta et imposuit duobus pueris suis, qui et portaverunt coram eo.
2KGS|5|24|Cumque venisset ad collem, tulit de manu eorum et reposuit in domo; dimisitque viros et abierunt.
2KGS|5|25|Ipse autem ingressus stetit coram domino suo. Et dixit Eliseus: " Unde venis, Giezi? ". Qui respondit: " Non ivit servus tuus quoquam ".
2KGS|5|26|At ille: " Nonne, ait, cor meum in praesenti erat, quando reversus est homo de curru suo in occursum tui? Estne tempus accipere argentum et accipere vestes et oliveta et vineta et oves et boves et servos et ancillas?
2KGS|5|27|Sed et lepra Naaman adhaerebit tibi et semini tuo in sempiternum ". Et egressus est ab eo leprosus quasi nix.
2KGS|6|1|Dixerunt autem filii prophetarum ad Eliseum: " Ecce locus, in quo habitamus coram te, angustus est nobis.
2KGS|6|2|Eamus usque ad Iordanem, et tollant singuli de silva materias singulas, ut aedificemus nobis ibi locum ad habitandum ". Qui dixit: " Ite ".
2KGS|6|3|Et ait unus ex illis: " Veni ergo et tu cum servis tuis ". Respondit: " Ego veniam ".
2KGS|6|4|Et abiit cum eis. Cumque venissent ad Iordanem, caedebant ligna.
2KGS|6|5|Accidit autem, ut, cum unus materiam succidisset, caderet ferrum securis in aquam; exclamavitque ille et ait: " Heu, domine mi! Et hoc ipsum mutuo acceperam! ".
2KGS|6|6|Dixit autem homo Dei: " Ubi cecidit? ". At ille monstravit ei locum. Praecidit ergo lignum et misit illuc, natavitque ferrum.
2KGS|6|7|Et ait: " Tolle!". Qui extendit manum et tulit illud.
2KGS|6|8|Rex autem Syriae pugnabat contra Israel; consiliumque iniit cum servis suis dicens: " In loco illo et illo ponamus insidias ".
2KGS|6|9|Misit itaque vir Dei ad regem Israel dicens: " Cave, ne transeas in loco illo, quia ibi Syri in insidiis sunt ".
2KGS|6|10|Misit rex Israel ad locum, quem dixerat ei vir Dei et de quo praemonuerat eum, et observavit se ibi non semel neque bis.
2KGS|6|11|Conturbatumque est cor regis Syriae pro hac re et, convocatis servis suis, ait: " Quare non indicatis mihi quis proditor mei sit apud regem Israel? ".
2KGS|6|12|Dixitque unus servorum eius: " Nequaquam, domine mi rex. Sed Eliseus propheta, qui est in Israel, indicat regi Israel omnia verba, quaecumque locutus fueris in conclavi tuo ".
2KGS|6|13|Dixit eis: " Ite et videte ubi sit, ut mittam et capiam eum ". Annuntiaveruntque ei dicentes: " Ecce in Dothain ".
2KGS|6|14|Misit ergo illuc equos et currus et robur exercitus; qui cum venissent nocte, circumdederunt civitatem.
2KGS|6|15|Consurgens autem diluculo minister viri Dei egressus est viditque exercitum in circuitu civitatis et equos et currus nuntiavitque ei dicens: Heu, domine mi, quid faciemus? ".
2KGS|6|16|At ille respondit: "Noli timere; plures enim nobiscum sunt quam cum illis".
2KGS|6|17|Oravitque Eliseus dicens: " Domine, aperi oculos huius, ut videat ". Et aperuit Dominus oculos pueri, et vidit, et ecce mons plenus equorum et curruum igneorum in circuitu Elisei.
2KGS|6|18|Hostes vero descenderunt ad eum. Porro Eliseus oravit Dominum dicens: " Percute, obsecro, gentem hanc caecitate! ". Percussitque eos Dominus, ne viderent iuxta verbum Elisei.
2KGS|6|19|Dixit autem ad eos Eliseus: " Non est haec via, nec ista est civitas; sequimini me, et ostendam vobis virum, quem quaeritis ". Duxit ergo eos in Samariam.
2KGS|6|20|Cumque ingressi fuissent in Samaria, dixit Eliseus: " Domine, aperi oculos istorum, ut videant ". Aperuitque Dominus oculos eorum, et viderunt esse se in medio Samariae.
2KGS|6|21|Dixitque rex Israel ad Eliseum, cum vidisset eos: " Numquid percutiam eos, pater mi? ".
2KGS|6|22|At ille ait: " Non percuties; neque enim, quos cepisti gladio et arcu tuo, percutis. Pone panem et aquam coram eis, ut comedant et bibant et vadant ad dominum suum ".
2KGS|6|23|Appositaque est eis ciborum magna praeparatio, et comederunt et biberunt, et dimisit eos; abieruntque ad dominum suum, et ultra non venerunt turmae Syriae in terram Israel.
2KGS|6|24|Factum est autem post haec, congregavit Benadad rex Syriae universum exercitum suum et ascendit et obsidebat Samariam.
2KGS|6|25|Factaque est fames magna in Samaria et tamdiu obsessa est, donec venumdaretur caput asini octoginta argenteis et quarta pars cabi stercoris columbarum quinque argenteis.
2KGS|6|26|Cumque rex Israel transiret per murum, mulier exclamavit ad eum dicens: Salva me, domine mi rex! ".
2KGS|6|27|Qui ait: " Non, salvet te te Dominus. Unde salvare te possum? De area an de torculari? ". Dixitque ad eam rex: " Quid tibi vis? ". Quae respondit:
2KGS|6|28|" Mulier ista dixit mihi: "Da filium tuum, ut comedamus eum hodie, et filium meum comedemus cras".
2KGS|6|29|Coximus ergo filium meum et comedimus. Dixique ei die altera: Da filium tuum, ut comedamus eum; quae abscondit filium suum ".
2KGS|6|30|Quod cum audisset rex, scidit vestimenta sua. Et transibat super murum, viditque omnis populus cilicium, quo vestitus erat ad carnem intrinsecus.
2KGS|6|31|Et ait: " Haec mihi faciat Deus et haec addat, si steterit caput Elisei filii Saphat super eum hodie ".
2KGS|6|32|Eliseus autem sedebat in domo sua, et senes sedebant cum eo. Praemisit itaque rex virum. Sed antequam veniret nuntius, Eliseus dixit ad senes: " Numquid scitis quod miserit filius homicidae hic, ut praecidatur caput meum? Videte ergo, cum venerit nuntius, claudite ostium et non sinatis eum introire; ecce enim sonitus pedum domini eius post eum est ".
2KGS|6|33|Et adhuc illo loquente eis, apparuit rex, qui veniebat ad eum, et ait: Ecce, tantum malum a Domino est; quid amplius exspectabo a Domino? ".
2KGS|7|1|Dixit autem Eliseus: " Audite verbum Domini. Haec dicit Dominus: In tempore hoc cras modius similae uno statere erit, et duo modii hordei statere uno in porta Samariae ".
2KGS|7|2|Respondens dux, super cuius manum rex incumbebat, homini Dei ait: " Si Dominus fecerit etiam cataractas in caelo, numquid poterit esse, quod loqueris? ". Qui ait: " Videbis oculis tuis et inde non comedes ".
2KGS|7|3|Quattuor ergo viri erant leprosi iuxta introitum portae; qui dixerunt ad invicem: " Quid hic esse volumus, donec moriamur?
2KGS|7|4|Sive ingredi voluerimus civitatem, fame moriemur; sive manserimus hic, moriendum nobis est. Venite igitur, et transfugiamus ad castra Syriae. Si pepercerint nobis, vivemus; si autem occidere voluerint, nihilominus moriemur ".
2KGS|7|5|Surrexerunt igitur vesperi, ut venirent ad castra Syriae. Cumque venissent ad principium castrorum Syriae, nullum ibidem reppererunt.
2KGS|7|6|Siquidem Dominus sonitum audiri fecerat in castris Syriae curruum et equorum et exercitus plurimi; dixeruntque ad invicem: " Ecce mercede conduxit adversum nos rex Israel reges Hetthaeorum et Aegyptiorum, ut venirent contra nos ".
2KGS|7|7|Surrexerunt ergo et fugerunt in tenebris et dereliquerunt tentoria sua et equos et asinos, castra, sicut erant; fugeruntque animas tantum suas salvare cupientes.
2KGS|7|8|Igitur cum venissent leprosi illi ad principium castrorum, ingressi sunt unum tabernaculum et comederunt et biberunt; tuleruntque inde argentum et aurum et vestes et abierunt et absconderunt. Et rursum reversi sunt ad aliud tabernaculum, et inde similiter auferentes absconderunt.
2KGS|7|9|Dixeruntque ad invicem: " Non recte facimus; haec enim dies boni nuntii est, et nos tacemus. Si noluerimus nuntiare usque mane, sceleris arguemur; venite, eamus et nuntiemus in aula regis ".
2KGS|7|10|Cumque venissent, vocaverunt portarios civitatis et narraverunt eis dicentes: " Ivimus ad castra Syriae et nullum ibidem repperimus hominum nisi equos et asinos alligatos et tentoria, sicut erant ".
2KGS|7|11|Clamaverunt ergo portarii et nuntiaverunt in palatio regis intrinsecus.
2KGS|7|12|Qui surrexit nocte et ait ad servos suos: " Dico vobis quid fecerint nobis Syri. Sciunt quia fame laboramus, et idcirco egressi sunt de castris et latitant in agris dicentes: "Cum egressi fuerint de civitate, capiemus eos viventes, et tunc civitatem ingredi poterimus" ".
2KGS|7|13|Respondit autem unus servorum eius: " Tollamus quinque equos, qui remanserunt in urbe; fiant sicut universa multitudo Israel, quae consumpta est; mittamus ergo et videamus ".
2KGS|7|14|Adduxerunt ergo duos currus cum equis, misitque rex post exercitum Syrorum dicens: " Ite et videte ".
2KGS|7|15|Qui abierunt post eos usque ad Iordanem; ecce autem omnis via plena erat vestibus et vasis, quae proiecerant Syri, cum turbarentur. Reversique nuntii indicaverunt regi.
2KGS|7|16|Et egressus populus diripuit castra Syriae; factusque est modius similae statere uno, et duo modii hordei statere uno iuxta verbum Domini.
2KGS|7|17|Porro rex ducem illum, in cuius manu incumbebat, constituit ad portam; quem conculcavit turba in introitu, et mortuus est iuxta quod locutus fuerat vir Dei, quando descenderat rex ad eum.
2KGS|7|18|Factumque est secundum sermonem viri Dei, quem dixerat regi, quando ait: " Duo modii hordei statere uno erunt, et modius similae statere uno hoc eodem tempore cras in porta Samariae ";
2KGS|7|19|quando responderat dux ille viro Dei et dixerat: " Etiamsi Dominus fecerit cataractas in caelo, numquid fieri poterit, quod loqueris? ", et dixerat ei: " Videbis oculis tuis et inde non comedes ".
2KGS|7|20|Evenit ergo ei, sicut praedictum erat, et conculcavit eum populus in porta, et mortuus est.
2KGS|8|1|Eliseus autem locutus est ad mulierem, cuius vivere fecerat fi lium, dicens: " Surge, vade tu et domus tua et peregrinare ubicumque reppereris; vocavit enim Dominus famem, et veniet super terram septem annis ".
2KGS|8|2|Quae surrexit et fecit iuxta verbum hominis Dei et vadens cum domo sua peregrinata est in terra Philisthim septem annis.
2KGS|8|3|Cumque finiti essent anni septem, reversa est mulier de terra Philisthim; et egressa est, ut interpellaret regem pro domo sua et agris suis.
2KGS|8|4|Rex autem loquebatur cum Giezi puero viri Dei dicens: " Narra mihi omnia magnalia, quae fecit Eliseus ".
2KGS|8|5|Cumque ille narraret regi quomodo mortuum suscitasset, apparuit mulier, cuius vivificaverat filium, clamans ad regem pro domo sua et pro agris suis. Dixitque Giezi: " Domine mi rex, haec est mulier, et hic filius eius, quem suscitavit Eliseus ".
2KGS|8|6|Et interrogavit rex mulierem, quae narravit ei. Deditque ei rex eunuchum unum dicens: " Restitue ei omnia, quae sua sunt, et universos reditus agrorum a die, qua reliquit terram usque ad praesens ".
2KGS|8|7|Venit quoque Eliseus Damascum, et Benadad rex Syriae aegrotabat. Nuntiaveruntque ei dicentes: " Venit vir Dei huc ".
2KGS|8|8|Et ait rex ad Hazael: " Tolle tecum munera et vade in occursum viri Dei et consule Dominum per eum dicens: Si evadere potero de infirmitate mea hac? ".
2KGS|8|9|Ivit igitur Hazael in occursum eius habens secum munera et omnia bona Damasci, onera quadraginta camelorum. Cumque stetisset coram eo, ait: " Filius tuus Benadad rex Syriae misit me ad te dicens: "Si sanari potero de infirmitate mea hac?" ".
2KGS|8|10|Dixitque ei Eliseus: " Vade, dic ei: Sanaberis. Porro ostendit mihi Dominus quia morte morietur ".
2KGS|8|11|Stetitque facies eius, et conturbatus est usque ad suffusionem vultus flevitque vir Dei.
2KGS|8|12|Cui Hazael ait: " Quare dominus meus flet? ". At ille respondit: " Quia scio, quae facturus sis filiis Israel mala: civitates eorum munitas igne succendes et iuvenes eorum interficies gladio et parvulos eorum elides et praegnantes discindes ".
2KGS|8|13|Dixitque Hazael: " Quid enim sum servus tuus canis, ut faciam rem istam magnam? ". Et ait Eliseus: " Ostendit mihi Dominus te regem Syriae fore ".
2KGS|8|14|Qui cum recessisset ab Eliseo, venit ad dominum suum. Qui ait ei: " Quid tibi dixit Eliseus? ". At ille respondit: " Dixit mihi: Recipies sanitatem ".
2KGS|8|15|Cumque venisset dies altera, tulit stragulum et intinxit aqua et expandit super faciem eius, et mortuus est; regnavitque Hazael pro eo.
2KGS|8|16|Anno quinto Ioram filii Achab regis Israel - Iosaphat autem erat rex Iudae - regnavit Ioram filius Iosaphat regis Iudae.
2KGS|8|17|Triginta duorum erat annorum, cum regnare coepisset, et octo annis regnavit in Ierusalem.
2KGS|8|18|Ambulavitque in viis regum Israel, sicut ambulaverat domus Achab; filia enim Achab erat uxor eius. Et fecit, quod malum est coram Domino.
2KGS|8|19|Noluit autem Dominus disperdere Iudam propter David servum suum, sicut promiserat ei, ut daret illi lucernam et filiis eius cunctis diebus.
2KGS|8|20|In diebus eius recessit Edom, ne esset sub Iuda, et constituit sibi regem.
2KGS|8|21|Venitque Ioram Seira et omnis currus cum eo; et surrexit nocte percussitque Idumaeos, qui eum circumdederant, et principes curruum; et populus fugit in tabernacula sua.
2KGS|8|22|Recessit ergo Edom, ne esset sub Iuda, usque ad diem hanc. Tunc recessit et Lobna in tempore illo.
2KGS|8|23|Reliqua autem gestorum Ioram et universa, quae fecit, nonne haec scripta sunt in libro annalium regum Iudae?
2KGS|8|24|Et dormivit Ioram cum patribus suis sepultusque est cum eis in civitate David; et regnavit Ochozias filius eius pro eo.
2KGS|8|25|Anno duodecimo Ioram filii Achab regis Israel regnavit Ochozias filius Ioram regis Iudae.
2KGS|8|26|Viginti duorum annorum erat Ochozias, cum regnare coepisset, et uno anno regnavit in Ierusalem. Nomen matris eius Athalia filia Amri regis Israel.
2KGS|8|27|Et ambulavit in viis domus Achab et fecit, quod malum est coram Domino, sicut domus Achab; gener enim domus Achab fuit.
2KGS|8|28|Abiit quoque cum Ioram filio Achab ad proeliandum contra Hazael regem Syriae in Ramoth Galaad; et vulneraverunt Syri Ioram.
2KGS|8|29|Qui reversus est, ut curaretur in Iezrahel de vulneribus, quibus vulneraverant eum Syri in Rama proeliantem contra Hazael regem Syriae. Porro Ochozias filius Ioram rex Iudae descendit invisere Ioram filium Achab in Iezrahel, quia aegrotabat.
2KGS|9|1|Eliseus autem prophetes vocavit unum de filiis prophetarum et ait illi: Accinge lumbos tuos et tolle lenticulam olei hanc in manu tua et vade in Ramoth Galaad.
2KGS|9|2|Cumque veneris illuc, videbis Iehu filium Iosaphat filii Namsi et ingressus suscitabis eum de medio fratrum suorum et introduces interius cubiculum.
2KGS|9|3|Tenensque lenticulam olei fundes super caput eius et dices: " Haec dicit Dominus: Unxi te regem super Israel ". Aperiesque ostium et fugies et non ibi subsistes ".
2KGS|9|4|Abiit ergo adulescens puer prophetae Ramoth Galaad
2KGS|9|5|et ingressus est. Ecce autem principes exercitus sedebant, et ait: " Verbum mihi ad te, princeps ". Dixitque Iehu: " Ad quem ex omnibus nobis?. At ille dixit: " Ad te, o princeps ".
2KGS|9|6|Et surrexit et ingressus est cubiculum. At ille fudit oleum super caput eius et ait: " Haec dicit Dominus, Deus Israel: Unxi te regem super populum Domini, super Israel.
2KGS|9|7|Percuties domum Achab domini tui, ut ulciscar sanguinem servorum meorum prophetarum et sanguinem omnium servorum Domini de manu Iezabel.
2KGS|9|8|Perdamque omnem domum Achab et interficiam de Achab quidquid masculini sexus et impuberem et puberem in Israel.
2KGS|9|9|Et dabo domum Achab sicut domum Ieroboam filii Nabat et sicut domum Baasa filii Ahiae.
2KGS|9|10|Iezabel quoque comedent canes in agro Iezrahel, nec erit qui sepeliat eam ". Aperuitque ostium et fugit.
2KGS|9|11|Iehu autem egressus est ad servos domini sui, qui dixerunt ei: " Rectene sunt omnia? Quid venit insanus iste ad te? ". Qui ait eis: " Nostis hominem et loquelam eius ".
2KGS|9|12|At illi responderunt: " Mendacium! Narra nobis! ". Qui ait eis: " Haec et haec locutus est mihi dicens: "Haec dicit Dominus: Unxi te regem super Israel" ".
2KGS|9|13|Festinaverunt itaque et unusquisque tollens pallium suum posuerunt sub pedibus eius super structuram graduum et cecinerunt tuba atque dixerunt: " Regnavit Iehu! ".
2KGS|9|14|Coniuravit ergo Iehu filius Iosaphat filii Namsi contra Ioram. Porro Ioram defenderat Ramoth Galaad ipse et omnis Israel contra Hazael regem Syriae
2KGS|9|15|et reversus fuerat, ut curaretur in Iezrahel propter vulnera, quia percusserant eum Syri proeliantem contra Hazael regem Syriae. Dixitque Iehu: " Si placet vobis, nemo egrediatur profugus de civitate, ne vadat et nuntiet in Iezrahel ".
2KGS|9|16|Et ascendit et profectus est in Iezrahel; Ioram enim aegrotabat ibi, et Ochozias rex Iudae descenderat ad visitandum Ioram.
2KGS|9|17|Igitur speculator, qui stabat super turrim Iezrahel, vidit globum Iehu venientis et ait: " Video ego globum ". Dixitque Ioram: " Tolle equitem et mitte in occursum eorum, et dicat vadens: "Rectene sunt omnia?" ".
2KGS|9|18|Abiit igitur, qui ascenderat equum in occursum eius, et ait: " Haec dicit rex: Pacatane sunt omnia? ". Dixitque ei Iehu: " Quid tibi et paci? Transi et sequere me ". Nuntiavit quoque speculator dicens: " Venit nuntius ad eos et non revertitur ".
2KGS|9|19|Misit etiam equitem secundum; venitque ad eos et ait: " Haec dicit rex: Num pax est? ". Et ait Iehu: " Quid tibi et paci? Transi et sequere me ".
2KGS|9|20|Nuntiavit autem speculator dicens: " Venit usque ad eos et non revertitur. Est autem incessus quasi incessus Iehu filii Namsi; praeceps enim graditur ".
2KGS|9|21|Et ait Ioram: " Iunge currum! ". Iunxeruntque currum eius, et egressus est Ioram rex Israel et Ochozias rex Iudae singuli in curribus suis. Egressique sunt in occursum Iehu et invenerunt eum in agro Naboth Iezrahelitis.
2KGS|9|22|Cumque vidisset Ioram Iehu, dixit: " Estne pax, Iehu? ". At ille respondit: " Quae pax? Adhuc fornicationes Iezabel matris tuae et veneficia eius multa vigent! ".
2KGS|9|23|Convertit autem Ioram manum suam et fugiens ait ad Ochoziam: " Insidiae, Ochozia! ".
2KGS|9|24|Porro Iehu tetendit arcum manu et percussit Ioram inter scapulas. Et egressa est sagitta per cor eius; statimque corruit in curru suo.
2KGS|9|25|Dixitque Iehu ad Badacer ducem: " Tolle, proice eum in agro Naboth Iezrahelitae! Memento enim: ego et tu eramus cum his, qui vectabantur gemini post Achab patrem huius, quando Dominus onus hoc levavit super eum dicens:
2KGS|9|26|"Pro sanguine Naboth et pro sanguine filiorum eius, quem vidi heri, ait Dominus, reddam tibi in agro isto, dicit Dominus". Nunc igitur tolle, proice eum in agro iuxta verbum Domini ".
2KGS|9|27|Ochozias autem rex Iudae videns hoc fugit per viam Bethgan; persecutusque est eum Iehu et ait: " Etiam hunc percutite! ". Et percusserunt eum in curru suo in ascensu Gaver, qui est iuxta Ieblaam. Qui fugit in Mageddo et mortuus est ibi.
2KGS|9|28|Et imposuerunt eum servi eius super currum suum et tulerunt Ierusalem sepelieruntque in sepulcro cum patribus suis in civitate David.
2KGS|9|29|Anno undecimo Ioram filii Achab regnavit Ochozias super Iudam.
2KGS|9|30|Venit Iehu Iezrahel. Porro Iezabel, introitu eius audito, depinxit oculos suos stibio et ornavit caput suum et respexit per fenestram
2KGS|9|31|ingredientem Iehu per portam et ait: " Numquid pax esse potest Zamri, qui interfecit dominum suum? ".
2KGS|9|32|Levavitque Iehu faciem suam ad fenestram et ait: " Quis est mecum, quisnam? ". Et inclinaverunt se ad eum duo vel tres eunuchi.
2KGS|9|33|At ille dixit eis: " Praecipitate eam deorsum! ". Et praecipitaverunt eam; aspersusque est sanguine paries et equi, qui conculcaverunt eam.
2KGS|9|34|Cumque ingressus esset, ut comederet biberetque, ait: " Ite, videte maledictam illam et sepelite eam, quia filia regis est ".
2KGS|9|35|Cumque issent, ut sepelirent eam, non invenerunt nisi calvariam et pedes et summas manus.
2KGS|9|36|Reversique nuntiaverunt ei. Et ait Iehu: " Sermo Domini est, quem locutus est per servum suum Eliam Thesbiten dicens: In agro Iezrahel comedent canes carnes Iezabel;
2KGS|9|37|et erit cadaver Iezabel sicut stercus super faciem terrae in agro Iezrahel, ita ut non dicatur: "Haeccine est illa Iezabel" ".
2KGS|10|1|Erant autem Achab septuaginta filii in Samaria. Scripsit ergo Iehu litteras et misit in Samariam ad optimates civitatis et ad maiores natu et ad nutricios filiorum Achab dicens:
2KGS|10|2|" Statim ut acceperitis litteras has, qui habetis filios domini vestri et currus et equos et civitatem firmam et arma,
2KGS|10|3|eligite meliorem et iustiorem de filiis domini vestri et ponite eum super solium patris sui et pugnate pro domo domini vestri ".
2KGS|10|4|Timuerunt illi vehementer et dixerunt: " Ecce duo reges non potuerunt stare coram eo, et quomodo nos valebimus resistere? ".
2KGS|10|5|Miserunt ergo praepositus domus et praefectus civitatis et maiores natu et nutricii ad Iehu dicentes: " Servi tui sumus: quaecumque iusseris, faciemus nec constituemus regem; quodcumque tibi placet, fac ".
2KGS|10|6|Rescripsit autem eis litteras secundo dicens: " Si mei estis et oboeditis mihi, tollite capita virorum filiorum domini vestri et venite ad me hac eadem hora cras in Iezrahel ". Porro filii regis, septuaginta viri, apud optimates civitatis nutriebantur.
2KGS|10|7|Cumque venissent litterae ad eos, tulerunt filios regis et occiderunt septuaginta viros et posuerunt capita eorum in cophinis et miserunt ad eum in Iezrahel.
2KGS|10|8|Venit autem nuntius et indicavit ei dicens: " Attulerunt capita filiorum regis". Qui respondit: " Ponite ea duos acervos iuxta introitum portae usque mane ".
2KGS|10|9|Cumque diluxisset, egressus est et stans dixit ad omnem populum: " Vos iusti estis; ecce ego coniuravi contra dominum meum et interfeci eum, sed quis percussit omnes hos?
2KGS|10|10|Videte ergo nunc quoniam non cecidit de sermonibus Domini in terram, quos locutus est Dominus super domum Achab, et Dominus fecit, quod locutus est in manu servi sui Eliae ".
2KGS|10|11|Percussit igitur Iehu omnes, qui reliqui erant de domo Achab in Iezrahel, et universos optimates eius et notos et sacerdotes, donec non remanerent ex eo reliquiae.
2KGS|10|12|Et surrexit et intravit. Deinde profectus est in Samariam; cumque esset ad Betheced Pastorum in via,
2KGS|10|13|invenit fratres Ochoziae regis Iudae dixitque ad eos: " Quinam estis vos? ". At illi responderunt: " Fratres Ochoziae sumus et descendimus ad salutandos filios regis et filios dominae reginae ".
2KGS|10|14|Qui ait: " Comprehendite eos vivos ". Quos cum comprehendissent vivos, iugulaverunt eos iuxta cisternam Betheced, quadraginta duos viros, et non reliquit ex eis quemquam.
2KGS|10|15|Cumque abisset inde, invenit Ionadab filium Rechab in occursum sibi et benedixit ei. Et ait ad eum: " Numquid est cor tuum rectum sicut cor meum cum corde tuo? ". Et ait Ionadab: " Est ". " Si est, inquit, da manum tuam. Qui dedit manum suam. At ille levavit eum ad se in curru
2KGS|10|16|dixitque ad eum: " Veni mecum et vide zelum meum pro Domino ". Et impositum currui suo
2KGS|10|17|duxit in Samariam. Et percussit omnes, qui reliqui fuerant de Achab in Samaria usque ad unum, iuxta verbum Domini, quod locutus est per Eliam.
2KGS|10|18|Congregavit ergo Iehu omnem populum et dixit ad eos: " Achab coluit Baal parum, ego autem colam eum amplius.
2KGS|10|19|Nunc igitur omnes prophetas Baal et universos servos eius et cunctos sacerdotes ipsius vocate ad me; nullus sit qui non veniat. Sacrificium enim grande est mihi Baal; quicumque defuerit, non vivet ". Porro Iehu faciebat hoc insidiose, ut disperderet cultores Baal.
2KGS|10|20|Dixitque: " Sanctificate diem sollemnem Baal ". Vocaveruntque.
2KGS|10|21|Et misit Iehu in universos terminos Israel, et venerunt cuncti servi Baal; non fuit residuus, ne unus quidem qui non veniret. Et ingressi sunt templum Baal, et repleta est domus Baal a summo usque ad summum.
2KGS|10|22|Dixitque ei, qui erat super vestes: " Profer vestimenta universis servis Baal ". Et protulit eis vestes.
2KGS|10|23|Ingressusque Iehu et Ionadab filius Rechab templum Baal ait cultoribus Baal: " Perquirite et videte, ne quis forte vobiscum sit de servis Domini, sed ut sint soli servi Baal ".
2KGS|10|24|Ingressi sunt igitur, ut facerent victimas et holocausta; Iehu autem praeparaverat sibi foris octoginta viros et dixerat eis: " Quicumque permiserit fugere de hominibus his, quos ego adduxero in manus vestras, anima eius erit pro anima illius ".
2KGS|10|25|Factum est ergo cum completum esset holocaustum, praecepit Iehu cursoribus et ducibus suis: " Ingredimini et percutite eos; nullus evadat!. Percusseruntque eos cursores et duces ore gladii et proiecerunt. Tunc ierunt usque in dabir templi Baal.
2KGS|10|26|Et protulerunt lapidem Baal et combusserunt
2KGS|10|27|et comminuerunt eum. Destruxerunt quoque aedem Baal et fecerunt pro ea latrinas usque diem hanc.
2KGS|10|28|Delevit itaque Iehu Baal de Israel.
2KGS|10|29|Verumtamen a peccatis Ieroboam filii Nabat, qui peccare fecerat Israel, non recessit; nec dereliquit vitulos aureos, qui erant in Bethel et in Dan.
2KGS|10|30|Dixit autem Dominus ad Iehu: " Quia studiose fecisti, quod rectum erat in oculis meis et omnia quae erant in corde meo fecisti contra domum Achab, filii tui usque ad quartam generationem sedebunt super thronum Israel ".
2KGS|10|31|Porro Iehu non custodivit, ut ambularet in lege Domini, Dei Israel, in toto corde suo; non enim recessit a peccatis Ieroboam, qui peccare fecerat Israel.
2KGS|10|32|In diebus illis coepit Dominus discindere in Israel; percussitque eos Hazael in universis finibus Israel
2KGS|10|33|a Iordane contra orientalem plagam omnem terram Galaad et Gad et Ruben et Manasse, ab Aroer, quae est super torrentem Arnon, et Galaad et Basan.
2KGS|10|34|Reliqua autem gestorum Iehu et universa, quae fecit, et fortitudo eius, nonne haec scripta sunt in libro annalium regum Israel?
2KGS|10|35|Et dormivit Iehu cum patribus suis, sepelieruntque eum in Samaria; et regnavit Ioachaz filius eius pro eo.
2KGS|10|36|Dies autem, quos regnavit Iehu super Israel, viginti et octo anni sunt, in Samaria.
2KGS|11|1|Athalia vero mater Ochoziae videns mortuum filium suum surrexit et interfecit omne semen regium.
2KGS|11|2|Tollens autem Iosaba filia regis Ioram soror Ochoziae Ioas filium Ochoziae furata est eum de medio filiorum regis, qui interficiebantur, et nutricem eius in cubiculo lectulorum, et absconderunt eum a facie Athaliae, ut non interficeretur.
2KGS|11|3|Eratque cum ea in domo Domini clam sex annis; porro Athalia regnavit super terram.
2KGS|11|4|Anno autem septimo misit Ioiada et assumens centuriones Carum et cursorum introduxit ad se in templum Domini pepigitque cum eis foedus; et adiurans eos in domo Domini ostendit eis filium regis
2KGS|11|5|et praecepit illis dicens: " Hoc est, quod facere debetis: tertia pars vestrum introeat sabbato et observet excubitum domus regis;
2KGS|11|6|tertia autem pars ad portam Sur, et tertia pars sit ad portam, quae est post habitaculum cursorum, et custodietis excubitum domus per vices.
2KGS|11|7|Duae vero partes e vobis omnes egredientes sabbato custodiant excubias domus Domini circum regem.
2KGS|11|8|Et vallabitis eum habentes arma in manibus vestris; si quis autem ingressus fuerit saeptum templi, interficiatur; eritisque cum rege introeunte et egrediente.
2KGS|11|9|Et fecerunt centuriones iuxta omnia, quae praeceperat eis Ioiada sacerdos, et assumentes singuli viros suos, qui ingrediebantur sabbato, cum his, qui egrediebantur sabbato, venerunt ad Ioiada sacerdotem.
2KGS|11|10|Qui dedit centurionibus hastas et peltas regis David, quae erant in domo Domini.
2KGS|11|11|Et steterunt cursores singuli habentes arma in manu sua a parte templi dextera usque ad partem templi sinistram contra altare et aedem circum regem.
2KGS|11|12|Produxitque filium regis et dedit ei diadema et testimonium; feceruntque eum regem et unxerunt et plaudentes manu dixerunt: " Vivat rex! ".
2KGS|11|13|Audivit autem Athalia vocem populi et ingressa ad turbas in templum Domini
2KGS|11|14|vidit regem stantem super tribunal iuxta morem et principes et tubas prope eum omnemque populum terrae laetantem et canentem tubis; et scidit vestimenta sua clamavitque: " Coniuratio, coniuratio! ".
2KGS|11|15|Praecepit autem Ioiada sacerdos centurionibus, qui erant super exercitum, et ait eis: " Educite eam extra consaepta templi, et, quicumque secutus eam fuerit, feriatur gladio ". Dixerat enim sacerdos: " Non occidatur in templo Domini ".
2KGS|11|16|Imposueruntque ei manus et impegerunt eam per viam introitus Equorum in palatium, et interfecta est ibi.
2KGS|11|17|Pepigit igitur Ioiada foedus inter Dominum et inter regem et inter populum, ut esset populus Domini, et inter regem et populum.
2KGS|11|18|Ingressusque est omnis populus terrae templum Baal, et destruxerunt illud et aras eius et imagines contriverunt valide; Matthan quoque sacerdotem Baal occiderunt coram altaribus.Et posuit sacerdos custodias in domo Domini
2KGS|11|19|tulitque centuriones et Cares et cursores et omnem populum terrae; deduxeruntque regem de domo Domini. Et venerunt per viam portae Cursorum in palatium, et sedit super thronum regum.
2KGS|11|20|Laetatusque est omnis populus terrae, et civitas conquievit; Athalia autem occisa est gladio in domo regis.
2KGS|12|1|Septemque annorum erat Ioas, cum regnare coepisset.
2KGS|12|2|Anno septimo Iehu regnavit Ioas; quadraginta annis regnavit in Ierusalem. Nomen matris eius Sebia de Bersabee.
2KGS|12|3|Fecitque Ioas rectum coram Domino cunctis diebus, quibus docuit eum Ioiada sacerdos.
2KGS|12|4|Verumtamen excelsa non abstulit; adhuc populus immolabat et adolebat in excelsis.
2KGS|12|5|Dixitque Ioas ad sacerdotes: " Omnem pecuniam sanctorum, quae illata fuerit in templum Domini a praetereuntibus, quae offertur pro pretio animae, et quam sponte et arbitrio cordis sui inferunt in templum Domini,
2KGS|12|6|accipiant illam singuli sacerdotes a notis suis et instaurent sartatecta domus, si quid necessarium viderint instauratione ".
2KGS|12|7|Igitur usque ad vicesimum tertium annum regis Ioas non instauraverunt sacerdotes sartatecta templi.
2KGS|12|8|Vocavitque rex Ioas Ioiada pontificem et sacerdotes dicens eis: " Quare sartatecta non instauratis templi? Nolite ergo amplius accipere pecuniam a notis vestris, sed ad instaurationem templi reddite eam ".
2KGS|12|9|Acquieveruntque sacerdotes ultra non accipere pecuniam a populo nec instaurare sartatecta domus.
2KGS|12|10|Et tulit Ioiada pontifex gazophylacium unum aperuitque foramen desuper et posuit illud iuxta altare ad dexteram ingredientium domum Domini; mittebantque in eo sacerdotes, qui custodiebant ostia, omnem pecuniam, quae deferebatur ad templum Domini.
2KGS|12|11|Cumque viderent multam pecuniam esse in gazophylacio, ascendebat scriba regis et pontifex, colligebantque et numerabant pecuniam, quae inveniebatur in domo Domini,
2KGS|12|12|et dabant eam iuxta numerum atque mensuram in manu opificum, qui operibus praepositi erant in domo Domini; ipsique impendebant eam in fabris lignorum et in structoribus, qui operabantur in domo Domini,
2KGS|12|13|et in caementariis et in his, qui caedebant saxa, et ut emerent ligna et lapides de lapicidinis, ut instaurarentur sartatecta domus Domini, et pro universis, quae indigebant expensa ad muniendam domum.
2KGS|12|14|Verumtamen non fiebant pelves argenteae templi Domini et cultri et paterae et tubae, omne vas aureum et argenteum, de pecunia, quae inferebatur in templum Domini;
2KGS|12|15|opificibus enim dabatur, ut instauraretur templum Domini.
2KGS|12|16|Et non fiebat ratio his hominibus, qui accipiebant pecuniam, ut distribuerent eam operariis; illi enim in fide agebant.
2KGS|12|17|Pecuniam vero pro delicto et pecuniam pro peccatis non inferebatur in templum Domini, quia sacerdotum erat.
2KGS|12|18|Tunc ascendit Hazael rex Syriae et pugnabat contra Geth; cepitque eam et direxit faciem suam, ut ascenderet in Ierusalem.
2KGS|12|19|Quam ob rem tulit Ioas rex Iudae omnia sanctificata, quae consecraverant Iosaphat et Ioram et Ochozias patres eius reges Iudae, et quae ipse obtulerat, et universum aurum, quod inveniri potuit in thesauris templi Domini et in palatio regis, misitque Hazaeli regi Syriae; et recessit ab Ierusalem.
2KGS|12|20|Reliqua autem gestorum Ioas et universa, quae fecit, nonne haec scripta sunt in libro annalium regum Iudae?
2KGS|12|21|Surrexerunt autem servi eius et coniuraverunt inter se percusseruntque Ioas in domo Mello in descensu Sella.
2KGS|12|22|Iozachar namque filius Semath et Iozabad filius Somer servi eius percusserunt eum, et mortuus est; et sepelierunt eum cum patribus suis in civitate David. Regnavitque Amasias filius eius pro eo.
2KGS|13|1|Anno vicesimo tertio Ioas fi lii Ochoziae regis Iudae re gnavit Ioachaz filius Iehu super Israel in Samaria decem et septem annis.
2KGS|13|2|Et fecit malum coram Domino secutusque est peccatum Ieroboam filii Nabat, qui peccare fecit Israel; non declinavit ab eo.
2KGS|13|3|Iratusque est furor Domini contra Israel et tradidit eos in manu Hazael regis Syriae et in manu Benadad filii Hazael cunctis diebus.
2KGS|13|4|Deprecatus est autem Ioachaz faciem Domini, et audivit eum Dominus; vidit enim angustiam Israel, qua attriverat eos rex Syriae.
2KGS|13|5|Et dedit Dominus Israeli salvatorem, et liberatus est de manu Syriae; habitaveruntque filii Israel in tabernaculis suis sicut heri et nudiustertius.
2KGS|13|6|Verumtamen non recesserunt a peccatis domus Ieroboam, qui peccare fecit Israel; in ipsis ambulaverunt. Siquidem et palus permansit in Samaria.
2KGS|13|7|Et non reliquit Dominus Ioachaz de populo nisi quinquaginta equites et decem currus et decem milia peditum; interfecerat enim eos rex Syriae et redegerat quasi pulverem in tritura areae.
2KGS|13|8|Reliqua autem gestorum Ioachaz et universa, quae fecit, sed et fortitudo eius, nonne haec scripta sunt in libro annalium regum Israel?
2KGS|13|9|Dormivitque Ioachaz cum patribus suis, et sepelierunt eum in Samaria. Regnavitque Ioas filius eius pro eo.
2KGS|13|10|Anno tricesimo septimo Ioas regis Iudae regnavit Ioas filius Ioachaz super Israel in Samaria sedecim annis.
2KGS|13|11|Et fecit, quod malum est in conspectu Domini; non declinavit ab omnibus peccatis Ieroboam filii Nabat, qui peccare fecit Israel; in ipsis ambulavit.
2KGS|13|12|Reliqua autem gestorum Ioas et universa, quae fecit, sed et fortitudo eius, quomodo pugnaverit contra Amasiam regem Iudae, nonne haec scripta sunt in libro annalium regum Israel?
2KGS|13|13|Et dormivit Ioas cum patribus suis; Ieroboam autem sedit super solium eius. Porro Ioas sepultus est in Samaria cum regibus Israel.
2KGS|13|14|Eliseus autem aegrotabat infirmitate, qua et mortuus est; descenditque ad eum Ioas rex Israel et flebat coram eo dicebatque: " Pater mi, pater mi, currus Israel et auriga eius! ".
2KGS|13|15|Et ait illi Eliseus: "Affer arcum et sagittas". Cumque attulisset ad eum arcum et sagittas,
2KGS|13|16|dixit ad regem Israel: " Pone manum tuam super arcum ". Et, cum posuisset ille manum suam, superposuit Eliseus manus suas manibus regis
2KGS|13|17|et ait: " Aperi fenestram orientalem ". Cumque aperuisset, dixit Eliseus: "Iace sagittam!". Et iecit. Et ait Eliseus: " Sagitta salutis Domini, et sagitta salutis contra Syriam. Percutiesque Syriam in Aphec, donec consumas eam ".
2KGS|13|18|Et ait: " Tolle sagittas ". Qui cum tulisset, rursum dixit ei: " Percute iaculo terram!". Et, cum percussisset tribus vicibus et stetisset,
2KGS|13|19|iratus est contra eum vir Dei et ait: " Si percussisses quinquies aut sexies, percussisses Syriam usque ad consummationem; nunc autem tribus vicibus percuties eam ".
2KGS|13|20|Mortuus est ergo Eliseus, et sepelierunt eum. Latrunculi autem de Moab venerunt in terra in ipso anno.
2KGS|13|21|Quidam autem sepelientes hominem viderunt latrunculos et proiecerunt cadaver in sepulcro Elisei et abierunt. Quod cum tetigisset ossa Elisei, revixit homo et stetit super pedes suos.
2KGS|13|22|Igitur Hazael rex Syriae afflixit Israel cunctis diebus Ioachaz.
2KGS|13|23|Et misertus est Dominus eorum et reversus est ad eos propter pactum suum, quod habebat cum Abraham, Isaac et Iacob, et noluit disperdere eos neque proicere penitus usque in praesens tempus.
2KGS|13|24|Mortuus est autem Hazael rex Syriae; et regnavit Benadad filius eius pro eo.
2KGS|13|25|Porro Ioas filius Ioachaz tulit urbes de manu Benadad filii Hazael, quas tulerat de manu Ioachaz patris sui iure proelii; tribus vicibus percussit eum Ioas et reddidit civitates Israeli.
2KGS|14|1|Anno secundo Ioas filii Ioachaz regis Israel regnavit Amasias filius Ioas regis Iudae.
2KGS|14|2|Viginti quinque annorum erat, cum regnare coepisset, viginti autem et novem annis regnavit in Ierusalem. Nomen matris eius Ioaden de Ierusalem.
2KGS|14|3|Et fecit rectum coram Domino, verumtamen non ut David pater eius. Iuxta omnia, quae fecit Ioas pater suus, fecit,
2KGS|14|4|nisi hoc quod excelsa non abstulit; adhuc enim populus immolabat et adolebat in excelsis.
2KGS|14|5|Cumque obtinuisset regnum, percussit servos suos, qui interfecerant regem patrem suum;
2KGS|14|6|filios autem eorum, qui occiderant, non occidit, iuxta quod scriptum est in libro legis Moysi, sicut praecepit Dominus dicens: " Non morientur patres pro filiis, neque filii morientur pro patribus, sed unusquisque in peccato suo morietur ".
2KGS|14|7|Ipse percussit Edom in valle Salinarum decem milia et apprehendit Petram in proelio vocavitque nomen eius Iecethel usque in praesentem diem.
2KGS|14|8|Tunc misit Amasias nuntios ad Ioas filium Ioachaz filii Iehu regem Israel dicens: " Veni, et videamus nos ".
2KGS|14|9|Remisitque Ioas rex Israel ad Amasiam regem Iudae dicens: " Carduus Libani misit ad cedrum, quae est in Libano, dicens: "Da filiam tuam filio meo uxorem". Transieruntque bestiae agri, quae sunt in Libano, et conculcaverunt carduum.
2KGS|14|10|Percutiens invaluisti super Edom, et sublevavit te cor tuum; contentus esto gloria et sede in domo tua. Quare provocas malum, ut cadas tu et Iuda tecum? ".
2KGS|14|11|Et non acquievit Amasias.Ascenditque Ioas rex Israel, et viderunt se ipse et Amasias rex Iudae in Bethsames oppido Iudae.
2KGS|14|12|Percussusque est Iuda coram Israel, et fugerunt unusquisque in tabernacula sua.
2KGS|14|13|Amasiam vero regem Iudae filium Ioas filii Ochoziae cepit Ioas rex Israel in Bethsames et adduxit eum in Ierusalem. Et interrupit murum Ierusalem a porta Ephraim usque ad portam Anguli quadringentis cubitis.
2KGS|14|14|Tulitque omne aurum et argentum et universa vasa, quae inventa sunt in domo Domini et in thesauris regis, et obsides; et reversus est Samariam.
2KGS|14|15|Reliqua autem gestorum Ioas, quae fecit, et fortitudo eius, qua pugnavit contra Amasiam regem Iudae, nonne haec scripta sunt in libro annalium regum Israel?
2KGS|14|16|Dormivitque Ioas cum patribus suis et sepultus est in Samaria cum regibus Israel; et regnavit Ieroboam filius eius pro eo.
2KGS|14|17|Vixit autem Amasias filius Ioas rex Iudae, postquam mortuus est Ioas filius Ioachaz rex Israel, quindecim annis.
2KGS|14|18|Reliqua autem gestorum Amasiae, nonne haec scripta sunt in libro annalium regum Iudae?
2KGS|14|19|Factaque est contra eum coniuratio in Ierusalem, at ille fugit in Lachis; miseruntque post eum in Lachis et interfecerunt eum ibi.
2KGS|14|20|Et asportaverunt eum in equis; sepultusque est in Ierusalem cum patribus suis in civitate David.
2KGS|14|21|Tulit autem universus populus Iudae Azariam annos natum sedecim, et constituerunt eum regem pro patre eius Amasia.
2KGS|14|22|Ipse aedificavit Ailath et restituit eam Iudae, postquam dormivit rex cum patribus suis.
2KGS|14|23|Anno quinto decimo Amasiae filii Ioas regis Iudae regnavit Ieroboam filius Ioas regis Israel in Samaria quadraginta et uno anno.
2KGS|14|24|Et fecit, quod malum est coram Domino; non recessit ab omnibus peccatis Ieroboam filii Nabat, qui peccare fecit Israel.
2KGS|14|25|Ipse restituit terminos Israel ab introitu Emath usque ad mare Arabae iuxta sermonem Domini, Dei Israel, quem locutus est per servum suum Ionam filium Amathi prophetam, qui erat de Gethhepher.
2KGS|14|26|Vidit enim Dominus afflictionem Israel amaram nimis, et quod consumpti essent impuber et puber, et non esset qui auxiliaretur Israel.
2KGS|14|27|Nec locutus est Dominus, ut deleret nomen Israel de sub caelo, sed salvavit eos in manu Ieroboam filii Ioas.
2KGS|14|28|Reliqua autem gestorum Ieroboam et universa, quae fecit, et fortitudo eius, qua proeliatus est, et quomodo restituit, quod de finibus Damasci et Emath fuerat Iudae, Israeli, nonne haec scripta sunt in libro annalium regum Israel?
2KGS|14|29|Dormivitque Ieroboam cum patribus suis regibus Israel; et regnavit Zacharias filius eius pro eo.
2KGS|15|1|Anno vicesimo septimo Ieroboam regis Israel regnavit Azarias filius Amasiae regis Iudae.
2KGS|15|2|Sedecim annorum erat, cum regnare coepisset, et quinquaginta duobus annis regnavit in Ierusalem. Nomen matris eius Iechelia de Ierusalem.
2KGS|15|3|Fecitque, quod erat placitum coram Domino, iuxta omnia, quae fecit Amasias pater eius.
2KGS|15|4|Verumtamen excelsa non est demolitus; adhuc populus sacrificabat et adolebat in excelsis.
2KGS|15|5|Percussit autem Dominus regem, et fuit leprosus usque in diem mortis suae et habitabat in domo separata seorsum; Ioatham vero filius regis gubernabat palatium et iudicabat populum terrae.
2KGS|15|6|Reliqua autem gestorum Azariae et universa, quae fecit, nonne haec scripta sunt in libro annalium regum Iudae?
2KGS|15|7|Et dormivit Azarias cum patribus suis, sepelieruntque eum cum maioribus suis in civitate David; et regnavit Ioatham filius eius pro eo.
2KGS|15|8|Anno tricesimo octavo Azariae regis Iudae regnavit Zacharias filius Ieroboam super Israel in Samaria sex mensibus.
2KGS|15|9|Et fecit, quod malum est coram Domino, sicut fecerant patres eius; non recessit a peccatis Ieroboam filii Nabat, qui peccare fecit Israel.
2KGS|15|10|Coniuravit autem contra eum Sellum filius Iabes percussitque eum in Ieblaam et interfecit; regnavitque pro eo.
2KGS|15|11|Reliqua autem gestorum Zachariae, nonne haec scripta sunt in libro annalium regum Israel?
2KGS|15|12|Iste est sermo Domini, quem locutus est ad Iehu dicens: " Filii usque ad quartam generationem sedebunt de te super thronum Israel ". Factumque est ita.
2KGS|15|13|Sellum filius Iabes regnavit tricesimo nono anno Azariae regis Iudae; regnavit autem uno mense in Samaria.
2KGS|15|14|Et ascendit Manahem filius Gadi de Thersa venitque Samariam et percussit Sellum filium Iabes in Samaria et interfecit eum; regnavitque pro eo.
2KGS|15|15|Reliqua autem gestorum Sellum et coniuratio eius, per quam tetendit insidias, nonne haec scripta sunt in libro annalium regum Israel?
2KGS|15|16|Tunc percussit Manahem Thapsam et omnes, qui erant in ea, et terminos eius de Thersa; noluerant enim aperire ei. Et interfecit omnes praegnantes eius et scidit eas.
2KGS|15|17|Anno tricesimo nono Azariae regis Iudae regnavit Manahem filius Gadi super Israel decem annis in Samaria.
2KGS|15|18|Fecitque, quod erat malum coram Domino; non recessit a peccatis Ieroboam filii Nabat, qui peccare fecit Israel. In diebus eius
2KGS|15|19|venit Phul rex Assyriorum in terram, et dedit Manahem Phul mille talenta argenti, ut esset ei in auxilio et firmaret regnum eius.
2KGS|15|20|Indixitque Manahem argentum super Israel cunctis potentibus, ut daret regi Assyriorum, quinquaginta siclos argenti per singulos. Reversusque est rex Assyriorum et non est moratus in terra.
2KGS|15|21|Reliqua autem gestorum Manahem et universa, quae fecit, nonne haec scripta sunt in libro annalium regum Israel?
2KGS|15|22|Et dormivit Manahem cum patribus suis; regnavitque Phaceia filius eius pro eo.
2KGS|15|23|Anno quinquagesimo Azariae regis Iudae regnavit Phaceia filius Manahem super Israel in Samaria biennio.
2KGS|15|24|Et fecit, quod erat malum coram Domino; non recessit a peccatis Ieroboam filii Nabat, qui peccare fecit Israel.
2KGS|15|25|Coniuravit autem adversus eum Phacee filius Romeliae dux eius et percussit eum in Samaria in turre domus regiae, et cum eo erant quinquaginta viri de filiis Galaaditarum. Et interfecit eum regnavitque pro eo.
2KGS|15|26|Reliqua autem gestorum Phaceia et universa, quae fecit, nonne haec scripta sunt in libro annalium regum Israel?
2KGS|15|27|Anno quinquagesimo secundo Azariae regis Iudae regnavit Phacee filius Romeliae super Israel in Samaria viginti annis.
2KGS|15|28|Et fecit, quod malum erat coram Domino; non recessit a peccatis Ieroboam filii Nabat, qui peccare fecit Israel.
2KGS|15|29|In diebus Phacee regis Israel venit Theglathphalasar rex Assur et cepit Ahion et Abelbethmaacha et Ianoe et Cedes et Asor et Galaad et Galilaeam, universam terram Nephthali, et transtulit eos in Assur.
2KGS|15|30|Coniuravit autem et tetendit insidias Osee filius Ela contra Phacee filium Romeliae; et percussit eum et interfecit regnavitque pro eo vicesimo anno Ioatham filii Oziae.
2KGS|15|31|Reliqua autem gestorum Phacee et universa, quae fecit, nonne haec scripta sunt in libro annalium regum Israel?
2KGS|15|32|Anno secundo Phacee filii Romeliae regis Israel regnavit Ioatham filius Oziae regis Iudae.
2KGS|15|33|Viginti quinque annorum erat, cum regnare coepisset, et sedecim annis regnavit in Ierusalem. Nomen matris eius Ierusa filia Sadoc.
2KGS|15|34|Fecitque, quod erat placitum coram Domino; iuxta omnia, quae fecerat Ozias pater suus, operatus est.
2KGS|15|35|Verumtamen excelsa non abstulit; adhuc populus immolabat et adolebat in excelsis. Ipse aedificavit portam domus Domini superiorem.
2KGS|15|36|Reliqua autem gestorum Ioatham et universa, quae fecit, nonne haec scripta sunt in libro annalium regum Iudae?
2KGS|15|37|In diebus illis coepit Dominus mittere in Iudam Rasin regem Syriae et Phacee filium Romeliae.
2KGS|15|38|Et dormivit Ioatham cum patribus suis sepultusque est cum eis in civitate David patris sui; et regnavit Achaz filius eius pro eo.
2KGS|16|1|Anno septimo decimo Phacee filii Romeliae regnavit Achaz filius Ioatham regis Iudae.
2KGS|16|2|Viginti annorum erat Achaz, cum regnare coepisset, et sedecim annis regnavit in Ierusalem; non fecit, quod erat placitum in conspectu Domini Dei sui, sicut David pater eius,
2KGS|16|3|sed ambulavit in via regum Israel. Insuper et filium suum consecravit transferens per ignem secundum abominationes gentium, quas dissipavit Dominus coram filiis Israel;
2KGS|16|4|immolabat quoque et adolebat in excelsis et in collibus et sub omni ligno frondoso.
2KGS|16|5|Tunc ascendit Rasin rex Syriae et Phacee filius Romeliae rex Israel in Ierusalem ad proeliandum; cumque obsiderent Achaz, non valuerunt superare eum.
2KGS|16|6|In tempore illo restituit Rasin rex Syriae Ailath ad Edom et eiecit Iudaeos de Ailath; et Idumaei venerunt in Ailath et habitaverunt ibi usque in diem hanc.
2KGS|16|7|Misit autem Achaz nuntios ad Theglathphalasar regem Assyriorum dicens: " Servus tuus et filius tuus ego sum. Ascende et salvum me fac de manu regis Syriae et de manu regis Israel, qui consurrexerunt adversum me ".
2KGS|16|8|Et cum collegisset argentum et aurum, quod invenire potuit in domo Domini et in thesauris regis, misit regi Assyriorum munera.
2KGS|16|9|Qui et acquievit voluntati eius. Ascendit enim rex Assyriorum in Damascum et vastavit eam et transtulit habitatores eius in Cir; Rasin autem interfecit.
2KGS|16|10|Perrexitque rex Achaz in occursum Theglathphalasar regis Assyriorum in Damascum. Cumque vidisset altare Damasci, misit rex Achaz ad Uriam sacerdotem exemplar eius et descriptionem omnis operis eius.
2KGS|16|11|Exstruxitque Urias sacerdos altare; iuxta omnia, quae miserat rex Achaz de Damasco, ita fecit Urias sacerdos, donec veniret rex Achaz de Damasco.
2KGS|16|12|Cumque venisset rex de Damasco, vidit altare et accessit ad illud ascenditque
2KGS|16|13|et adolevit holocausta sua et oblationes et libavit libamina et fudit sanguinem pacificorum suorum super altare.
2KGS|16|14|Porro altare aeneum, quod erat coram Domino, transtulit de facie templi et de loco inter altare et templum Domini posuitque illud ex latere altaris ad aquilonem.
2KGS|16|15|Praecepit quoque rex Achaz Uriae sacerdoti dicens: " Super altare maius offer holocaustum matutinum et oblationem vespertinam et holocaustum regis et oblationem eius et holocaustum universi populi terrae et oblationem eorum et libamina eorum; et omnem sanguinem holocausti et universum sanguinem sacrificii super illud effundes. De altari vero aeneo erit mihi deliberandum ".
2KGS|16|16|Fecit igitur Urias sacerdos iuxta omnia, quae praeceperat rex Achaz.
2KGS|16|17|Excidit autem rex Achaz limbos basium et removit luterem, qui erat desuper, et mare deposuit de bobus aeneis, qui sustentabant illud, et posuit super pavimentum stratum lapide.
2KGS|16|18|Musach (id est Porticum) quoque sabbati, quod aedificatum erat in templo, et ingressum regis exterius convertit in templo Domini propter regem Assyriorum.
2KGS|16|19|Reliqua autem gestorum Achaz, quae fecit, nonne haec scripta sunt in libro annalium regum Iudae?
2KGS|16|20|Dormivitque Achaz cum patribus suis et sepultus est cum eis in civitate David; et regnavit Ezechias filius eius pro eo.
2KGS|17|1|Anno duodecimo Achaz regis Iudae regnavit Osee filius Ela in Samaria super Israel novem annis.
2KGS|17|2|Fecitque malum coram Domino, sed non sicut reges Israel, qui ante eum fuerant.
2KGS|17|3|Contra hunc ascendit Salmanasar rex Assyriorum; et factus est ei Osee servus reddebatque illi tributa.
2KGS|17|4|Cumque deprehendisset rex Assyriorum Osee quod rebellare nitens misisset nuntios ad Sua regem Aegypti nec praestaret tributa regi Assyriorum, sicut singulis annis solitus erat, apprehendit eum et vinctum misit in carcerem.
2KGS|17|5|Pervagatusque est omnem terram et ascendens Samariam obsedit eam tribus annis.
2KGS|17|6|Anno autem nono Osee cepit rex Assyriorum Samariam et transtulit Israel in Assur posuitque eos in Hala et iuxta Habor fluvium Gozan et in civitatibus Medorum.
2KGS|17|7|Factum est enim hoc, cum peccassent filii Israel Domino Deo suo, qui eduxerat eos de terra Aegypti, de manu pharaonis regis Aegypti: coluerunt deos alienos.
2KGS|17|8|Et ambulaverunt iuxta ritus gentium, quas consumpserat Dominus in conspectu filiorum Israel et regum Israel, qui similiter fecerant.
2KGS|17|9|Et offenderunt filii Israel operibus non rectis Dominum Deum suum et aedificaverunt sibi excelsa in cunctis urbibus suis a turre custodum usque ad civitatem munitam.
2KGS|17|10|Feceruntque sibi lapides et palos in omni colle sublimi et subter omne lignum nemorosum
2KGS|17|11|et adolebant ibi in omnibus excelsis sicut gentes, quas transtulerat Dominus a facie eorum; feceruntque pessima irritantes Dominum
2KGS|17|12|et coluerunt idola immunda, de quibus praecepit Dominus eis, ne facerent hoc.
2KGS|17|13|Et testificatus est Dominus in Israel et in Iuda per manum omnium prophetarum et videntium dicens: " Revertimini a viis vestris pessimis et custodite mandata mea et praecepta iuxta omnem legem, quam praecepi patribus vestris, et sicut misi ad vos in manu servorum meorum prophetarum.
2KGS|17|14|Qui non audierunt, sed induraverunt cervicem suam iuxta cervicem patrum suorum, qui noluerunt credere in Dominum Deum suum.
2KGS|17|15|Et abiecerunt legitima eius et pactum, quod pepigit cum patribus eorum, et testificationes, quibus contestatus est eos; secutique sunt vanitates et vani facti sunt et secuti sunt gentes, quae erant per circuitum eorum, super quibus praeceperat Dominus eis ut non facerent, sicut et illae faciebant.
2KGS|17|16|Et dereliquerunt omnia praecepta Domini Dei sui feceruntque sibi conflatiles duos vitulos et palum et adoraverunt universam militiam caeli servieruntque Baal
2KGS|17|17|et consecrabant filios suos et filias suas per ignem; et divinationibus inserviebant et auguriis et tradiderunt se, ut facerent malum coram Domino et irritarent eum.
2KGS|17|18|Iratusque est Dominus vehementer Israel et abstulit eos de conspectu suo, et non remansit nisi tribus Iudae tantummodo.
2KGS|17|19|Sed nec ipse Iuda custodivit mandata Domini Dei sui; verum ambulavit in erroribus Israel, quos operatus fuerat.
2KGS|17|20|Proiecitque Dominus omne semen Israel et afflixit eos et tradidit in manu diripientium, donec proiceret eos a facie sua,
2KGS|17|21|ex eo iam tempore, quo scissus est Israel a domo David, et constituerunt sibi regem Ieroboam filium Nabat; separavit enim Ieroboam Israel a Domino et peccare eos fecit peccatum magnum.
2KGS|17|22|Et ambulaverunt filii Israel in universis peccatis Ieroboam, quae fecerat; non recesserunt ab eis,
2KGS|17|23|usquequo auferret Dominus Israel a facie sua, sicut locutus fuerat in manu omnium servorum suorum prophetarum. Translatusque est Israel de terra sua in Assur usque in diem hanc.
2KGS|17|24|Adduxit autem rex Assyriorum de Babylone et de Chutha et de Ava et de Emath et de Sepharvaim et collocavit eos in civitatibus Samariae pro filiis Israel, qui possederunt Samariam et habitaverunt in urbibus eius.
2KGS|17|25|Cumque ibi habitare coepissent, non timebant Dominum. Et immisit eis Dominus leones, qui interficiebant inter eos.
2KGS|17|26|Nuntiatumque est regi Assyriorum et dictum: " Gentes, quas transtulisti et habitare fecisti in civitatibus Samariae, ignorant legitima Dei terrae; et immisit eis leones, et ecce interficiunt eos, eo quod ignorent ritum Dei terrae ".
2KGS|17|27|Praecepit autem rex Assyriorum dicens: " Ducite illuc unum de sacerdotibus, quos inde captivos adduxistis, et vadat et habitet cum eis et doceat eos legitima Dei terrae ".
2KGS|17|28|Igitur cum venisset unus de sacerdotibus his, qui captivi ducti fuerant de Samaria, habitavit in Bethel et docebat eos quomodo colerent Dominum.
2KGS|17|29|Et unaquaeque gens fabricata est deum suum; posueruntque eos in fanis excelsis, quae fecerant Samaritae, gens et gens in urbibus suis, in quibus habitabant.
2KGS|17|30|Viri enim Babylonii fecerunt Socchothbenoth, viri autem Chutheni fecerunt Nergel, et viri de Emath fecerunt Asima;
2KGS|17|31|porro Hevaei fecerunt Nebahaz et Tharthac, hi autem, qui erant de Sepharvaim, comburebant filios suos igne Adramelech et Anamelech diis Sepharvaim.
2KGS|17|32|Et nihilominus colebant Dominum. Fecerunt autem sibi de medio ipsorum sacerdotes excelsorum et ponebant eos in fanis excelsorum;
2KGS|17|33|et, cum Dominum colerent, diis quoque suis serviebant iuxta consuetudinem gentium, de quibus translati fuerant Samariam.
2KGS|17|34|Usque in praesentem diem morem sequuntur antiquum: non timent Dominum neque custodiunt instituta et iudicium ipsorum et legem et mandatum, quod praeceperat Dominus filiis Iacob, quem cognominavit Israel,
2KGS|17|35|et percusserat cum eis pactum et mandaverat eis dicens: " Nolite timere deos alienos et non adoretis eos neque colatis et non immoletis eis,
2KGS|17|36|sed Dominum, qui eduxit vos de terra Aegypti in fortitudine magna et in brachio extento, ipsum timete, illum adorate et ipsi immolate.
2KGS|17|37|Instituta quoque et iudicia et legem et mandatum, quod scripsit vobis, custodite, ut faciatis cunctis diebus; et non timeatis deos alienos.
2KGS|17|38|Et pactum, quod percussi vobiscum, nolite oblivisci nec timeatis deos alienos,
2KGS|17|39|sed Dominum Deum vestrum timete, et ipse eruet vos de manu omnium inimicorum vestrorum ".
2KGS|17|40|Illi vero non audierunt, sed iuxta consuetudinem suam pristinam perpetrabant.
2KGS|17|41|Fuerunt igitur gentes istae timentes quidem Dominum, sed nihilominus et idolis suis servientes; nam et filii eorum et nepotes, sicut fecerunt parentes sui, ita faciunt usque in praesentem diem.
2KGS|18|1|Anno tertio Osee filii Ela regis Israel regnavit Ezechias filius Achaz regis Iudae.
2KGS|18|2|Viginti quinque annorum erat, cum regnare coepisset, et viginti et novem annis regnavit in Ierusalem. Nomen matris eius Abi filia Zachariae.
2KGS|18|3|Fecitque, quod erat bonum coram Domino, iuxta omnia, quae fecerat David pater suus.
2KGS|18|4|Ipse dissipavit excelsa et contrivit lapides et succidit palum confregitque serpentem aeneum, quem fecerat Moyses; siquidem usque ad illud tempus filii Israel adolebant ei; vocabatur Nohestan.
2KGS|18|5|In Domino, Deo Israel, speravit. Itaque post eum non fuit similis ei de cunctis regibus Iudae sed neque in his, qui ante eum fuerunt.
2KGS|18|6|Et adhaesit Domino et non recessit a vestigiis eius fecitque mandata eius, quae praeceperat Dominus Moysi,
2KGS|18|7|unde et erat Dominus cum eo, et in cunctis, ad quae procedebat, prospere agebat.Rebellavit quoque contra regem Assyriorum et non servivit ei.
2KGS|18|8|Ipse percussit Philisthaeos usque Gazam et terminos eius, a turre custodum usque ad civitatem munitam.
2KGS|18|9|Anno quarto regis Ezechiae, qui erat annus septimus Osee filii Ela regis Israel, ascendit Salmanasar rex Assvriorum Samariam et oppugnavit eam
2KGS|18|10|et cepit. Post annos tres, anno sexto Ezechiae, id est nono anno Osee regis Israel, capta est Samaria.
2KGS|18|11|Et transtulit rex Assyriorum Israel in Assur collocavitque eos in Hala et Habor iuxta fluvium Gozan et in civitatibus Medorum,
2KGS|18|12|quia non audierunt vocem Domini Dei sui, sed praetergressi sunt pactum eius; omnia, quae praeceperat Moyses servus Domini, non audierunt neque fecerunt.
2KGS|18|13|Anno quarto decimo regis Ezechiae ascendit Sennacherib rex Assyriorum ad universas civitates Iudae munitas et cepit eas.
2KGS|18|14|Tunc misit Ezechias rex Iudae nuntios ad regem Assyriorum Lachis dicens: " Peccavi. Recede a me, et omne, quod imposueris mihi, feram ". Indixit itaque rex Assyriorum Ezechiae regi Iudae trecenta talenta argenti et triginta talenta auri;
2KGS|18|15|deditque Ezechias omne argentum, quod repertum fuerat in domo Domini et in thesauris regis.
2KGS|18|16|In tempore illo confregit Ezechias valvas templi Domini et postes, quos ipse inauraverat, et dedit aurum regi Assyriorum.
2KGS|18|17|Misit autem rex Assyriorum Tharthan et Rabsaris et Rabsacen de Lachis ad regem Ezechiam cum manu valida Ierusalem. Qui cum ascendissent, venerunt in Ierusalem et steterunt iuxta aquae ductum piscinae superioris, quae est in via agri fullonis,
2KGS|18|18|vocaveruntque regem. Egressus est autem ad eos Eliachim filius Helciae praepositus domus et Sobna scriba et Ioah filius Asaph a commentariis.
2KGS|18|19|Dixitque ad eos Rabsaces: " Loquimini Ezechiae: Haec dicit rex magnus, rex Assyriorum: Quae est ista fiducia, qua niteris?
2KGS|18|20|Forsitan putas verbum labiorum esse consilium et fortitudinem ad proelium? In quo confidis, ut audeas rebellare contra me?
2KGS|18|21|An speras in baculo arundineo atque confracto, Aegypto, super quem, si incubuerit homo, comminutus ingreditur manum eius et perforabit eam? Sic est pharao rex Aegypti omnibus, qui confidunt in eo.
2KGS|18|22|Quod si dixeritis mihi: "In Domino Deo nostro habemus fiduciam", nonne iste est, cuius abstulit Ezechias excelsa et altaria et praecepit Iudae et Ierusalem: "Ante altare hoc adorabitis in Ierusalem?".
2KGS|18|23|Nunc igitur spondete cum domino meo rege Assyriorum; dabo tibi duo milia equorum; et vide an habere valeas ascensores eorum.
2KGS|18|24|Et quomodo potes in fugam vertere unum satrapam de servis domini mei minimis? An fiduciam habes in Aegypto propter currus et equites?
2KGS|18|25|Numquid sine Domini voluntate ascendi ad locum istum, ut demolirer eum? Dominus dixit mihi: "Ascende ad terram hanc et demolire eam" ".
2KGS|18|26|Dixerunt autem Eliachim filius Helciae et Sobna et Ioah Rabsaci: " Precamur, ut loquaris nobis servis tuis Aramaice, siquidem intellegimus hanc linguam, et non loquaris nobis Iudaice, audiente populo, qui est super murum ".
2KGS|18|27|Responditque eis Rabsaces: " Numquid ad dominum tuum et ad te misit me dominus meus, ut loquerer sermones hos, et non ad viros, qui sedent super murum, ut comedant stercora sua et bibant urinam suam vobiscum? ".
2KGS|18|28|Stetit itaque Rabsaces et clamavit voce magna Iudaice et ait: " Audite verba regis magni, regis Assyriorum:
2KGS|18|29|Haec dicit rex: Non vos seducat Ezechias; non enim poterit eruere vos de manu mea!
2KGS|18|30|Neque fiduciam vobis tribuat super Domino dicens: "Eruens liberabit nos Dominus, et non tradetur civitas haec in manu regis Assyriorum".
2KGS|18|31|Nolite audire Ezechiam! Haec enim dicit rex Assyriorum: Facite mecum benedictionem et egredimini ad me, et comedet unusquisque de vinea sua et de ficu sua, et bibetis aquas de cisternis vestris,
2KGS|18|32|donec veniam et transferam vos in terram, quae similis terrae vestrae est, in terram fructiferam et fertilem vini, terram panis et vinearum, terram olivarum olei ac mellis; et vivetis et non moriemini. Nolite audire Ezechiam, qui vos decipit dicens: "Dominus liberabit nos!".
2KGS|18|33|Numquid liberaverunt dii gentium unusquisque terram suam de manu regis Assyriorum?
2KGS|18|34|Ubi sunt dii Emath et Arphad? Ubi sunt dii Sepharvaim, Ana et Ava? Numquid liberaverunt Samariam de manu mea?
2KGS|18|35|Quinam illi sunt in universis diis terrarum, qui eruerunt regionem suam de manu mea, ut possit eruere Dominus Ierusalem de manu mea? ".
2KGS|18|36|Tacuit itaque populus et non respondit ei quidquam; siquidem praeceptum regis acceperant, ut non responderent ei.
2KGS|18|37|Venitque Eliachim filius Helciae praepositus domus et Sobna scriba et Ioah filius Asaph a commentariis ad Ezechiam, scissis vestibus, et nuntiaverunt ei verba Rabsacis.
2KGS|19|1|Quae cum audisset rex Ezechias, scidit vestimenta sua et opertus est sacco ingressusque est domum Domini.
2KGS|19|2|Et misit Eliachim praepositum domus et Sobnam scribam et senes de sacerdotibus opertos saccis ad Isaiam prophetam filium Amos.
2KGS|19|3|Qui dixerunt: " Haec dicit Ezechias: Dies tribulationis et increpationis et blasphemiae dies iste; venerunt filii usque ad partum, et vires non habet parturiens.
2KGS|19|4|Forte audiet Dominus Deus tuus universa verba Rabsacis, quem misit rex Assyriorum dominus suus, ut exprobraret Deum viventem, et puniet verba, quae audivit Dominus Deus tuus; et fac orationem pro reliquiis, quae remanent ".
2KGS|19|5|Venerunt ergo servi regis Ezechiae ad Isaiam.
2KGS|19|6|Dixitque eis Isaias: " Haec dicetis domino vestro: Haec dicit Dominus: Noli timere a facie sermonum, quos audisti, quibus blasphemaverunt pueri regis Assyriorum me;
2KGS|19|7|ecce ego immittam ei spiritum, et audiet nuntium et revertetur in terram suam; et deiciam eum gladio in terra sua ".
2KGS|19|8|Reversus est igitur Rabsaces et invenit regem Assyriorum oppugnantem Lobnam; audierat enim quod recessisset de Lachis.
2KGS|19|9|Cumque audisset de Tharaca rege Aethiopiae dicentes: " Ecce egressus est, ut pugnet adversum te ", iterum misit nuntios ad Ezechiam dicens:
2KGS|19|10|" Haec dicite Ezechiae regi Iudae: Non te seducat Deus tuus, in quo habes fiduciam, neque dicas: "Non tradetur Ierusalem in manu regis Assyriorum".
2KGS|19|11|Tu enim ipse audisti, quae fecerint reges Assyriorum universis terris, quomodo vastaverint eas. Num ergo solus poteris liberari?
2KGS|19|12|Numquid liberaverunt dii gentium singulos, quos vastaverunt patres mei, Gozan videlicet et Charran et Reseph et filios Eden, qui erant in Thelassar?
2KGS|19|13|Ubi est rex Emath et rex Arphad et rex civitatis Sepharvaim, Ana et Ava? ".
2KGS|19|14|Itaque cum accepisset Ezechias litteras de manu nuntiorum et legisset eas, ascendit in domum Domini et expandit eas coram Domino
2KGS|19|15|et oravit in conspectu eius dicens: " Domine, Deus Israel, qui sedes super cherubim! Tu es Deus solus regnorum omnium terrae, tu fecisti caelum et terram.
2KGS|19|16|Inclina aurem tuam et audi; aperi, Domine, oculos tuos et vide et audi omnia verba Sennacherib, qui misit, ut exprobraret Deum viventem.
2KGS|19|17|Vere, Domine, dissipaverunt reges Assyriorum gentes et terras earum
2KGS|19|18|et miserunt deos eorum in ignem; non enim erant dii, sed opera manuum hominum ex ligno et lapide, et perdiderunt eos.
2KGS|19|19|Nunc igitur, Domine Deus noster, salvos nos fac de manu eius, ut sciant omnia regna terrae quia tu, Domine, es Deus solus ".
2KGS|19|20|Misit autem Isaias filius Amos ad Ezechiam dicens: " Haec dicit Dominus, Deus Israel: Quae deprecatus es me super Sennacherib rege Assyriorum, audivi.
2KGS|19|21|Iste est sermo, quem locutus est Dominus de eo:Sprevit te et subsannavit virgo filia Sion;post tergum tuum caputmovit filia Ierusalem.
2KGS|19|22|Cui exprobrasti et quem blasphemasti?Contra quem exaltasti vocemet elevasti in excelsum oculos tuos? Contra Sanctum Israel!
2KGS|19|23|Per manum servorum tuorumexprobrasti Dominoet dixisti: "In multitudine curruum meorumascendi excelsa montium in summitate Libaniet succidi sublimes cedros eius,electas abietes eius,et ingressus sum usque ad terminos eius,silvam condensam.
2KGS|19|24|Ego fodi et bibi aquas alienaset siccavi vestigiis pedum meorum omnes aquas Aegypti".
2KGS|19|25|Numquid non audisti,ab initio quid fecerim?Ex diebus antiquis plasmavi illudet nunc adduxi;eruntque in eradicationem,in acervos ruinarum civitates munitae.
2KGS|19|26|Et, qui sedent in eis breviata manu,contremuerunt et confusi sunt;facti sunt quasi fenum agriet gramen virens, herba tectorum, quae arefacta est, antequam veniret ad maturitatem.
2KGS|19|27|Sessionem tuamet egressum tuum et introitum tuum ego praesciviet furorem tuum contra me;
2KGS|19|28|insanisti in me,et superbia tua ascendit in aures meas.Ponam itaque circulum in naribus tuiset frenum in labris tuiset reducam te in viam,per quam venisti.
2KGS|19|29|Tibi autem, Ezechia, hoc erit signum:Comede hoc anno, quod reppereris, in secundo autem anno, quae sponte nascuntur;porro in anno tertio seminate et metite,plantate vineas et comedite fructum earum.
2KGS|19|30|Et, quodcumque reliquum fuerit de domo Iudae,mittet radicem deorsumet faciet fructum sursum;
2KGS|19|31|de Ierusalem quippe egredientur reliquiae,et, quod relinquetur, de monte Sion.Zelus Domini exercituum faciet hoc.
2KGS|19|32|Quam ob rem haec dicit Dominus de rege Assyriorum:Non ingredietur urbem hancnec mittet in eam sagittamnec occurret ei clipeonec fundet aggerem circa eam.
2KGS|19|33|Per viam, qua venit, reverteturet civitatem hanc non ingredietur, dicit Dominus.
2KGS|19|34|Protegamque urbem hanc et salvabo eampropter me et propter David servum meum ".
2KGS|19|35|Factum est igitur in nocte illa: egressus est angelus Domini et percussit in castris Assyriorum centum octoginta quinque milia. Cumque diluculo surrexissent, viderunt omnia corpora mortuorum.
2KGS|19|36|Et recedens abiit et reversus est Sennacherib rex Assyriorum et mansit in Nineve.
2KGS|19|37|Cumque adoraret in templo Nesroch dei sui, Adramelech et Sarasar filii eius percusserunt eum gladio fugeruntque in terram Armeniorum. Et regnavit Asarhaddon filius eius pro eo.
2KGS|20|1|In diebus illis aegrotavit Ezechias usque ad mortem. Et venit ad eum Isaias filius Amos prophetes dixitque ei: " Haec dicit Dominus: Dispone domui tuae, morieris enim et non vives ".
2KGS|20|2|Qui convertit faciem suam ad parietem et oravit Dominum dicens:
2KGS|20|3|" Obsecro, Domine, memento quomodo ambulaverim coram te in veritate et in corde perfecto et, quod placitum est coram te, fecerim ". Flevit itaque Ezechias fletu magno.
2KGS|20|4|Et antequam egrederetur Isaias mediam partem atrii, factus est sermo Domini ad eum dicens:
2KGS|20|5|" Revertere et dic Ezechiae duci populi mei: Haec dicit Dominus, Deus David patris tui: Audivi orationem tuam, vidi lacrimam tuam, et ecce sano te; die tertio ascendes templum Domini.
2KGS|20|6|Et addam diebus tuis quindecim annos; sed et de manu regis Assyriorum liberabo te et civitatem hanc et protegam urbem istam propter me et propter David servum meum ".
2KGS|20|7|Dixitque Isaias: " Afferte massam ficorum ". Quam cum attulissent et posuissent super ulcus eius, curatus est.
2KGS|20|8|Dixit autem Ezechias ad Isaiam: " Quod erit signum quia Dominus me sanabit et quia ascensurus sum die tertio templum Domini? ".
2KGS|20|9|Cui ait Isaias: " Hoc erit tibi signum a Domino quod facturus sit Dominus sermonem, quem locutus est: Vis ut accedat umbra decem gradibus, an ut revertatur totidem gradibus? ".
2KGS|20|10|Et ait Ezechias: " Facile est umbram descendere decem gradibus, nec hoc volo ut fiat, sed ut revertatur retrorsum decem gradibus ".
2KGS|20|11|Invocavit itaque Isaias propheta Dominum; et reduxit umbram per gradus, quibus iam descenderat in gradibus Achaz, retrorsum decem gradibus.
2KGS|20|12|In tempore illo misit Merodachbaladan filius Baladan rex Babyloniorum litteras et munera ad Ezechiam; audierat enim quod aegrotasset Ezechias.
2KGS|20|13|Laetatus est autem in adventu eorum Ezechias et ostendit eis totam domum thesauri sui, argentum et aurum et aromata et oleum optimum et domum vasorum suorum et omnia, quae inventa sunt in thesauris suis: non fuit, quod non monstraret eis Ezechias in domo sua et in omni potestate sua.
2KGS|20|14|Venit autem Isaias propheta ad regem Ezechiam dixitque ei: " Quid dixerunt viri isti et unde venerunt ad te? ". Cui ait Ezechias: " De terra longinqua venerunt, de Babylone ".
2KGS|20|15|At ille respondit: " Quid viderunt in domo tua? ". Ait Ezechias: " Omnia, quae sunt in domo mea viderunt; nihil est, quod non monstraverim eis in thesauris meis ".
2KGS|20|16|Dixit itaque Isaias Ezechiae: " Audi sermonem Domini:
2KGS|20|17|Ecce dies venient, et auferentur omnia, quae sunt in domo tua, et quae condiderunt patres tui usque in diem hanc, in Babylone; non remanebit quidquam, ait Dominus.
2KGS|20|18|Sed et de filiis tuis, qui egredientur ex te, quos generabis, tollentur et erunt eunuchi in palatio regis Babylonis ".
2KGS|20|19|Dixit Ezechias ad Isaiam: " Bonus sermo Domini, quem locutus es ". Et ait: " Nonne erit pax et securitas in diebus meis? ".
2KGS|20|20|Reliqua autem gestorum Ezechiae et omnis fortitudo eius, et quomodo fecerit piscinam et aquae ductum et introduxerit aquas in civitatem, nonne haec scripta sunt in libro annalium regum Iudae?
2KGS|20|21|Dormivitque Ezechias cum patribus suis; et regnavit Manasses filius eius pro eo.
2KGS|21|1|Duodecim annorum erat Manasses, cum regnare coe pisset, et quinquaginta quinque annis regnavit in Ierusalem. Nomen matris eius Haphsiba.
2KGS|21|2|Fecitque malum in conspectu Domini iuxta abominationes gentium, quas delevit Dominus a facie filiorum Israel.
2KGS|21|3|Conversusque est et aedificavit excelsa, quae dissipaverat Ezechias pater eius, et erexit aras Baal et fecit palum, sicut fecerat Achab rex Israel, et adoravit omnem militiam caeli et coluit eam.
2KGS|21|4|Exstruxitque aras in domo Domini, de qua dixit Dominus: " In Ierusalem ponam nomen meum ".
2KGS|21|5|Et exstruxit altaria universae militiae caeli in duobus atriis templi Domini
2KGS|21|6|et traduxit filium suum per ignem et hariolatus est et observavit auguria et constituit pythones et haruspices multiplicavit, ut faceret malum coram Domino et irritaret eum.
2KGS|21|7|Posuit quoque palum Aserae, quem fecerat, in templo, super quo locutus est Dominus ad David et ad Salomonem filium eius: " In templo hoc et in Ierusalem, quam elegi de cunctis tribubus Israel, ponam nomen meum in sempiternum;
2KGS|21|8|et ultra non faciam commoveri pedem Israel de terra, quam dedi patribus eorum, sic tamen si custodierint opere omnia, quae praecepi eis, et universam legem, quam mandavit eis servus meus Moyses ".
2KGS|21|9|Illi vero non audierunt, sed seducti sunt a Manasse, ut facerent malum plus quam gentes, quas contrivit Dominus a facie filiorum Israel.
2KGS|21|10|Locutusque est Dominus in manu servorum suorum prophetarum dicens:
2KGS|21|11|" Quia fecit Manasses rex Iudae abominationes istas pessimas super omnia, quae fecerunt Amorraei ante eum, et peccare fecit etiam Iudam in idolis suis,
2KGS|21|12|propterea haec dicit Dominus, Deus Israel: Ecce ego inducam mala super Ierusalem et Iudam, ut quicumque audierit, tinniant ambae aures eius.
2KGS|21|13|Et extendam super Ierusalem funiculum Samariae et pondus domus Achab et extergam Ierusalem sicut qui extergit vas, extergit et convertit super faciem eius.
2KGS|21|14|Et proiciam reliquias hereditatis meae et tradam eas in manu inimicorum eius; eruntque in vastitate et rapina cunctis adversariis suis,
2KGS|21|15|eo quod fecerint malum coram me et perseveraverint irritantes me ex die, qua egressi sunt patres eorum ex Aegypto, usque ad diem hanc ".
2KGS|21|16|Insuper et sanguinem innoxium fudit Manasses multum nimis, donec impleret Ierusalem usque ad summum, absque peccatis suis, quibus peccare fecit Iudam, ut faceret malum coram Domino.
2KGS|21|17|Reliqua autem gestorum Manasse et universa, quae fecit, et peccatum eius, quod peccavit, nonne haec scripta sunt in libro annalium regum Iudae?
2KGS|21|18|Dormivitque Manasses cum patribus suis et sepultus est in horto domus suae, in horto Oza; et regnavit Amon filius eius pro eo.
2KGS|21|19|Viginti et duo annorum erat Amon, cum regnare coepisset, duobusque annis regnavit in Ierusalem. Nomen matris eius Mesallemeth filia Harus de Ieteba.
2KGS|21|20|Fecitque malum in conspectu Domini, sicut fecerat Manasses pater eius,
2KGS|21|21|et ambulavit in omni via, per quam ambulaverat pater eius; servivitque idolis, quibus servierat pater suus, et adoravit ea.
2KGS|21|22|Et dereliquit Dominum, Deum patrum suorum et non ambulavit in via Domini.
2KGS|21|23|Tetenderuntque ei insidias servi sui et interfecerunt regem in domo sua;
2KGS|21|24|percussit autem populus terrae omnes, qui coniuraverant contra regem Amon, et constituerunt sibi regem Iosiam filium eius pro eo.
2KGS|21|25|Reliqua autem gestorum Amon, quae fecit, nonne haec scripta sunt in libro annalium regum Iudae?
2KGS|21|26|Sepelieruntque eum in sepulcro suo in horto Oza; et regnavit Iosias filius eius pro eo.
2KGS|22|1|Octo annorum erat Iosias, cum regnare coepisset, et tri ginta et uno anno regnavit in Ierusalem. Nomen matris eius Idida filia Adaia de Bascath.
2KGS|22|2|Fecitque, quod placitum erat coram Domino, et ambulavit per omnes vias David patris sui; non declinavit ad dexteram sive ad sinistram.
2KGS|22|3|Anno autem octavo decimo regis Iosiae misit rex Saphan filium Eseliae filii Mesullam scribam ad templum Domini dicens ei:
2KGS|22|4|" Vade ad Helciam sacerdotem magnum, ut effundatur pecunia, quae illata est in templum Domini, quam collegerunt ianitores a populo,
2KGS|22|5|deturque opificibus praepositis in domo Domini, qui et distribuent eam his, qui operantur in templo Domini ad instauranda sartatecta templi,
2KGS|22|6|tignariis videlicet et caementariis et his, qui interrupta componunt, et ut emantur ligna et lapides de lapicidinis ad instaurandum templum.
2KGS|22|7|Verumtamen non supputetur eis argentum, quod accipiunt, quia in potestate habent et in fide ".
2KGS|22|8|Dixit autem Helcias pontifex ad Saphan scribam: " Librum legis repperi in domo Domini! ". Deditque Helcias volumen Saphan, qui et legit illud.
2KGS|22|9|Venit quoque Saphan scriba ad regem et renuntiavit ei, quod praeceperat, et ait: " Effuderunt servi tui pecuniam, quae reperta est in domo, et dederunt opificibus praefectis operum templi Domini ".
2KGS|22|10|Narravitque Saphan scriba regi dicens: " Librum dedit mihi Helcias sacerdos ".Quem cum legisset Saphan coram rege,
2KGS|22|11|et audisset rex verba libri legis, scidit vestimenta sua
2KGS|22|12|et praecepit Helciae sacerdoti et Ahicam filio Saphan et Achobor filio Micha et Saphan scribae et Asaiae servo regis dicens:
2KGS|22|13|" Ite et consulite Dominum super me et super populo et super omni Iuda de verbis voluminis istius, quod inventum est; magna enim ira Domini succensa est contra nos, quia non audierunt patres nostri verba libri huius, ut facerent omne, quod scriptum est nobis ".
2KGS|22|14|Ierunt itaque Helcias sacerdos et Ahicam et Achobor et Saphan et Asaia ad Holdam propheten uxorem Sellum filii Thecuae filii Haraas custodis vestium, quae habitabat in Ierusalem in secunda, locutique sunt ad eam,
2KGS|22|15|et illa respondit eis: " Haec dicit Dominus, Deus Israel: Dicite viro, qui misit vos ad me:
2KGS|22|16|Haec dicit Dominus: Ecce ego adducam mala super locum hunc et super habitatores eius omnia verba libri, quae legit rex Iudae,
2KGS|22|17|quia dereliquerunt me et sacrificaverunt diis alienis irritantes me in cunctis operibus manuum suarum; et succendetur indignatio mea in loco hoc et non exstinguetur.
2KGS|22|18|Regi autem Iudae, qui misit vos, ut consuleretis Dominum, sic dicetis: Haec dicit Dominus, Deus Israel: Pro eo quod audisti verba voluminis,
2KGS|22|19|et perterritum est cor tuum, et humiliatus es coram Domino, auditis sermonibus contra locum istum et habitatores eius, quo videlicet fierent in stuporem et in maledictum, et scidisti vestimenta tua et flevisti coram me, et ego audivi, ait Dominus;
2KGS|22|20|idcirco colligam te ad patres tuos, et colligeris ad sepulcrum tuum in pace, ut non videant oculi tui omnia mala, quae inducturus sum super locum istum ". Et renuntiaverunt regi, quod dixerat.
2KGS|23|1|Qui misit, et congregati sunt ad eum omnes senes Iudae et Ierusalem;
2KGS|23|2|ascenditque rex templum Domini et omnes viri Iudae universique, qui habitabant in Ierusalem cum eo, sacerdotes et prophetae et omnis populus a parvo usque ad magnum. Legitque, cunctis audientibus, omnia verba libri foederis, qui inventus est in domo Domini.
2KGS|23|3|Stetitque rex super gradum suum et percussit foedus coram Domino, ut ambularent post Dominum et custodirent praecepta eius et testimonia et legitima in omni corde et in tota anima et suscitarent verba foederis huius, quae scripta erant in libro illo. Acquievitque universus populus pacto.
2KGS|23|4|Et praecepit rex Helciae pontifici et sacerdotibus secundi ordinis et ianitoribus, ut proicerent de templo Domini omnia vasa, quae facta fuerant Baal et Aserae et universae militiae caeli; et combussit ea foris Ierusalem in convalle Cedron et tulit pulverem eorum in Bethel.
2KGS|23|5|Et delevit aedituos, quos posuerant reges Iudae ad sacrificandum in excelsis per civitates Iudae et in circuitu Ierusalem, et eos, qui adolebant Baal et soli et lunae et duodecim signis et omni militiae caeli.
2KGS|23|6|Et efferri fecit palum de domo Domini foras Ierusalem in convalle Cedron et combussit eum ibi et redegit in pulverem et proiecit super sepulcrum vulgi.
2KGS|23|7|Destruxit quoque aediculas prostibulorum, quae erant in domo Domini, in quibus mulieres texebant vestes pro Asera.
2KGS|23|8|Congregavitque omnes sacerdotes de civitatibus Iudae et contaminavit excelsa, ubi sacrificabant sacerdotes, de Gabaa usque Bersabee; et destruxit excelsa pilosorum in introitu portae Iosue principis civitatis, ad sinistram ingredientis portam civitatis.
2KGS|23|9|Verumtamen non ascendebant sacerdotes excelsorum ad altare Domini in Ierusalem, sed tantum comedebant azyma in medio fratrum suorum.
2KGS|23|10|Contaminavit quoque Topheth, quod est in convalle Benennom, ut nemo consecraret filium suum aut filiam per ignem Moloch.
2KGS|23|11|Abstulit quoque equos, quos dederant reges Iudae soli in introitu templi Domini iuxta cubiculum Nathanmelech eunuchi, quod erat in Pharurim; currus autem solis combussit igne.
2KGS|23|12|Altaria quoque, quae erant super tectum cenaculi Achaz, quae fecerant reges Iudae, et altaria, quae fecerat Manasses in duobus atriis templi Domini, destruxit rex et contrivit ea ibi et dispersit cinerem eorum in torrentem Cedron.
2KGS|23|13|Excelsa quoque, quae erant ex adverso Ierusalem ad dexteram partem montis Perditionis, quae aedificaverat Salomon rex Israel Astharoth idolo Sidoniorum et Chamos idolo Moab et Melchom idolo filiorum Ammon, polluit rex;
2KGS|23|14|et contrivit lapides et succidit palos replevitque loca eorum ossibus mortuorum.
2KGS|23|15|Insuper et altare, quod erat in Bethel, excelsum, quod fecerat Ieroboam filius Nabat, qui peccare fecit Israel, etiam altare illud et excelsum destruxit atque combussit et comminuit in pulverem succenditque palum.
2KGS|23|16|Et conversus Iosias vidit ibi sepulcra, quae erant in monte, misitque et tulit ossa de sepulcris et combussit ea super altare et polluit illud iuxta verbum Domini, quod clamaverat vir Dei, cum staret Ieroboam in die festo ad altare. Et conversus elevavit oculos in sepulcrum viri Dei, qui clamaverat verba haec,
2KGS|23|17|et ait: " Quis est titulus ille, quem video? ". Responderuntque ei cives illius urbis: " Sepulcrum est hominis Dei, qui venit de Iuda et clamavit verba haec, quae fecisti super altare Bethel ".
2KGS|23|18|Et ait: " Dimittite eum; nemo commoveat ossa eius ". Et intacta manserunt ossa illius cum ossibus prophetae, qui venerat de Samaria.
2KGS|23|19|Insuper et omnia fana excelsorum, quae erant in civitatibus Samariae, quae fecerant reges Israel ad irritandum Dominum, abstulit Iosias et fecit eis secundum omnia opera, quae fecerat in Bethel.
2KGS|23|20|Et immolavit universos sacerdotes excelsorum, qui erant ibi super altaria, et combussit ossa humana super ea; reversusque est Ierusalem.
2KGS|23|21|Et praecepit omni populo dicens: " Facite Pascha Domino Deo vestro secundum quod scriptum est in libro foederis huius ".
2KGS|23|22|Nec enim factum est Pascha tale a diebus iudicum, qui iudicaverunt Israel, et omnibus diebus regum Israel et regum Iudae,
2KGS|23|23|sicut in octavo decimo anno regis Iosiae factum est Pascha istud Domino in Ierusalem.
2KGS|23|24|Sed et pythones et hariolos et theraphim et idola abominationesque omnes, quae erant in terra Iudae et in Ierusalem, abstulit Iosias, ut statueret verba legis, quae scripta sunt in libro, quem invenit Helcias sacerdos in templo Domini.
2KGS|23|25|Similis illi non fuit ante eum rex, qui reverteretur ad Dominum in omni corde suo et in tota anima sua et in universa virtute sua iuxta omnem legem Moysi, neque post eum surrexit similis illi.
2KGS|23|26|Verumtamen non est aversus Dominus ab ira furoris sui magni, quo iratus est furor eius contra Iudam propter omnes irritationes, quibus provocaverat eum Manasses.
2KGS|23|27|Dixit itaque Dominus: " Etiam Iudam auferam a facie mea, sicut abstuli Israel, et proiciam civitatem hanc, quam elegi, Ierusalem et domum, de qua dixi: Erit nomen meum ibi ".
2KGS|23|28|Reliqua autem gestorum Iosiae et universa, quae fecit, nonne haec scripta sunt in libro annalium regum Iudae?
2KGS|23|29|In diebus eius ascendit pharao Nechao rex Aegypti contra regem Assyriorum ad flumen Euphraten. Et abiit Iosias rex in occursum eius, qui occidit eum in Mageddo, cum vidisset eum.
2KGS|23|30|Et portaverunt eum in curru servi sui mortuum de Mageddo et pertulerunt in Ierusalem et sepelierunt eum in sepulcro suo. Tulitque populus terrae Ioachaz filium Iosiae et unxerunt eum et constituerunt eum regem pro patre suo.
2KGS|23|31|Viginti trium annorum erat Ioachaz, cum regnare coepisset, et tribus mensibus regnavit in Ierusalem. Nomen matris eius Amital filia Ieremiae de Lobna.
2KGS|23|32|Et fecit malum coram Domino iuxta omnia, quae fecerant patres eius.
2KGS|23|33|Vinxitque eum pharao Nechao in Rebla, quae est in terra Emath, ne regnaret in Ierusalem; et imposuit multam terrae centum talentis argenti et talento auri;
2KGS|23|34|regemque constituit pharao Nechao Eliachim filium Iosiae pro Iosia patre eius vertitque nomen eius Ioachim. Porro Ioachaz tulit, et venit in Aegyptum et mortuus est ibi.
2KGS|23|35|Argentum autem et aurum dedit Ioachim pharaoni, cum indixisset terrae, ut conferretur argentum iuxta praeceptum pharaonis; et secundum uniuscuiusque aestimationem exegit tam argentum quam aurum de populo terrae, ut daret pharaoni Nechao.
2KGS|23|36|Viginti quinque annorum erat Ioachim, cum regnare coepisset, et undecim annis regnavit in Ierusalem. Nomen matris eius Zebida filia Phadaia de Ruma.
2KGS|23|37|Et fecit malum coram Domino iuxta omnia, quae fecerant patres eius.
2KGS|24|1|In diebus eius ascendit Nabuchodonosor rex Babylonis, et factus est ei Ioachim servus tribus annis et rursum rebellavit contra eum.
2KGS|24|2|Immisitque ei Dominus turmas Chaldaeorum et turmas Syriae, turmas Moab et turmas filiorum Ammon; et immisit eas in Iudam, ut disperderent eum iuxta verbum Domini, quod locutus erat per servos suos prophetas.
2KGS|24|3|Factum est autem hoc propter iram Domini contra Iudam, ut auferret eum de conspectu suo propter peccata Manasse universa, quae fecit,
2KGS|24|4|et propter sanguinem innoxium, quem effudit et implevit Ierusalem cruore innocentium; et ob hanc rem noluit Dominus propitiari.
2KGS|24|5|Reliqua autem gestorum Ioachim et universa, quae fecit, nonne haec scripta sunt in libro annalium regum Iudae? Et dormivit Ioachim cum patribus suis;
2KGS|24|6|regnavitque Ioachin filius eius pro eo.
2KGS|24|7|Et ultra non addidit rex Aegypti ut egrederetur de terra sua; tulerat enim rex Babylonis a rivo Aegypti usque ad fluvium Euphraten omnia, quae fuerant regis Aegypti.
2KGS|24|8|Decem et octo annorum erat Ioachin, cum regnare coepisset, et tribus mensibus regnavit in Ierusalem. Nomen matris eius Naestha filia Elnathan de Ierusalem.
2KGS|24|9|Et fecit malum coram Domino iuxta omnia, quae fecerat pater eius.
2KGS|24|10|In tempore illo ascenderunt servi Nabuchodonosor regis Babylonis in Ierusalem, et venit urbs in obsidione.
2KGS|24|11|Venitque Nabuchodonosor rex Babylonis ad civitatem, cum servi eius oppugnarent eam;
2KGS|24|12|egressusque est Ioachin rex Iudae ad regem Babylonis ipse et mater eius et servi eius et principes eius et eunuchi eius; et cepit eum rex Babylonis anno octavo regni sui.
2KGS|24|13|Et protulit inde omnes thesauros domus Domini et thesauros domus regiae et concidit universa vasa aurea, quae fecerat Salomon rex Israel in templo Domini, iuxta verbum Domini.
2KGS|24|14|Et transtulit omnem Ierusalem et universos principes et omnes fortes exercitus decem milia in captivitatem et omnem artificem et clusorem; nihilque relictum est, exceptis pauperibus populi terrae.
2KGS|24|15|Transtulit quoque Ioachin in Babylonem; et matrem regis et uxores regis et eunuchos eius et cives validos terrae duxit in captivitatem de Ierusalem in Babylonem
2KGS|24|16|et omnes viros robustos septem milia et artifices et clusores mille, omnes viros fortes bellatores; duxitque eos rex Babylonis captivos in Babylonem.
2KGS|24|17|Et constituit Matthaniam patruum eius pro eo; imposuitque nomen ei Sedeciam.
2KGS|24|18|Vicesimum et primum annum aetatis habebat Sedecias, cum regnare coepisset, et undecim annis regnavit in Ierusalem. Nomen matris eius erat Amital filia Ieremiae de Lobna.
2KGS|24|19|Et fecit malum coram Domino iuxta omnia, quae fecerat Ioachim;
2KGS|24|20|irascebatur enim Dominus contra Ierusalem et contra Iudam, donec proiceret eos a facie sua.Recessitque Sedecias a rege Babylonis.
2KGS|25|1|Factum est autem anno nono regni eius, mense decimo, decima die mensis venit Nabuchodonosor rex Babylonis ipse et omnis exercitus eius in Ierusalem; et circumdederunt eam et exstruxerunt in circuitu eius munitiones.
2KGS|25|2|Et clausa est civitas atque vallata usque ad undecimum annum regis Sedeciae.
2KGS|25|3|Nona die mensis quarti praevaluit fames in civitate, nec erat panis populo terrae.
2KGS|25|4|Et interrupta est civitas, et omnes viri bellatores fugerunt exieruntque de civitate nocte per viam portae, quae est inter duplicem murum ad hortum regis, obsidentibus Chaldaeis in circuitu civitatem. Abierunt itaque per viam, quae ducit ad Arabam.
2KGS|25|5|Et persecutus est exercitus Chaldaeorum regem comprehenditque eum in planitie Iericho, et omnis exercitus eius dispersus est et reliquit eum.
2KGS|25|6|Apprehensum ergo regem duxerunt ad regem Babylonis in Rebla, qui locutus est cum eo iudicium.
2KGS|25|7|Filios autem Sedeciae occidit coram eo et oculos eius effodit vinxitque eum catenis aereis et adduxit in Babylonem.
2KGS|25|8|Mense quinto septima die mensis, ipse est annus nonus decimus regis Babylonis, venit Nabuzardan princeps satellitum servus regis Babylonis Ierusalem
2KGS|25|9|et succendit domum Domini et domum regis et omnes domos Ierusalem; omnemque domum combussit igne.
2KGS|25|10|Et muros Ierusalem in circuitu destruxit omnis exercitus Chaldaeorum, qui erat cum principe satellitum.
2KGS|25|11|Reliquam autem populi partem, qui remanserat in civitate, et perfugas, qui transfugerant ad regem Babylonis, et reliquum vulgus transtulit Nabuzardan princeps satellitum;
2KGS|25|12|et de pauperibus terrae reliquit in vinitores et agricolas.
2KGS|25|13|Columnas autem aereas, quae erant in templo Domini, et bases et mare aereum, quod erat in domo Domini, confregerunt Chaldaei et transtulerunt aes omnium in Babylonem.
2KGS|25|14|Ollas quoque et trullas et cultros et phialas et omnia vasa aerea, in quibus ministrabant, tulerunt;
2KGS|25|15|necnon thymiamateria et phialas, quae aurea aurea et quae argentea argentea, tulit princeps satellitum;
2KGS|25|16|columnas duas, mare unum et bases, quas fecerat Salomon templo Domini; non erat pondus aeris omnium horum vasorum.
2KGS|25|17|Decem et octo cubitos altitudinis habebat columna una et capitellum aereum super se altitudinis quinque cubitorum; et reticulum et malogranata super capitellum in circuitu omnia aerea; similem et columna secunda habebat ornatum.
2KGS|25|18|Tulit quoque princeps satellitum Saraiam sacerdotem primum et Sophoniam sacerdotem secundum et tres ianitores
2KGS|25|19|et de civitate eunuchum unum, qui erat praefectus super viros bellatores, et quinque viros de his, qui steterant coram rege, quos repperit in civitate, et scribam principis exercitus, qui probabat tirones de populo terrae, et sexaginta viros e populo terrae, qui inventi fuerant in civitate;
2KGS|25|20|quos tollens Nabuzardan princeps satellitum duxit ad regem Babylonis in Rebla,
2KGS|25|21|percussitque eos rex Babylonis et interfecit in Rebla in terra Emath.Et translatus est Iuda de terra sua.
2KGS|25|22|Populo autem, qui relictus erat in terra Iudae, quem dimiserat Nabuchodonosor rex Babylonis, praefecit Godoliam filium Ahicam filii Saphan.
2KGS|25|23|Quod cum audissent omnes duces militum, videlicet quod constituisset rex Babylonis Godoliam, ipsi et viri, qui erant cum eis, venerunt ad Godoliam in Maspha: Ismael filius Nathaniae et Iohanan filius Caree et Saraia filius Thanehumeth Netophathites et Iezonias filius Maachathitis, ipsi et socii eorum.
2KGS|25|24|Iuravitque eis Godolias et sociis eorum dicens: " Nolite timere a servis Chaldaeorum; manete in terra et servite regi Babylonis, et bene erit vobis ".
2KGS|25|25|Factum est autem in mense septimo venit Ismael filius Nathaniae filii Elisama de semine regio et decem viri cum eo; percusseruntque Godoliam, qui mortuus est, sed et Iudaeos et Chaldaeos, qui erant cum eo in Maspha.
2KGS|25|26|Consurgens autem populus a parvo usque ad magnum et principes militum venerunt in Aegyptum timentes Chaldaeos.
2KGS|25|27|Factum est vero anno tricesimo septimo transmigrationis Ioachin regis Iudae, mense duodecimo vicesima septima die mensis sublevavit Evilmerodach rex Babylonis anno, quo regnare coeperat, caput Ioachin regis Iudae de carcere.
2KGS|25|28|Et locutus est ei benigna et posuit thronum eius super thronos regum, qui erant cum eo in Babylone,
2KGS|25|29|et mutavit vestes eius, quas habuerat in carcere; et comedebat panem semper in conspectu eius cunctis diebus vitae suae.
2KGS|25|30|Annonam quoque constituit ei absque intermissione, quae et dabatur ei a rege per singulos dies omnibus diebus vitae suae.
1CHR|1|1|Adam, Seth, Enos,
1CHR|1|2|Cainan, Malaleel, Iared,
1CHR|1|3|Henoch, Ma thusala, Lamech,
1CHR|1|4|Noe, Sem, Cham et Iapheth.
1CHR|1|5|Filii Iapheth: Gomer, Magog, Madai et Iavan, Thubal, Mosoch, Thiras.
1CHR|1|6|Porro filii Gomer: Aschenez et Riphath et Thogorma.
1CHR|1|7|Filii autem Iavan: Elisa et Tharsis, Getthim et Rodanim.
1CHR|1|8|Filii Cham: Chus et Mesraim, Phut et Chanaan.
1CHR|1|9|Filii autem Chus: Saba et Hevila, Sabatha et Regma et Sabathacha. Porro filii Regma: Saba et Dedan.
1CHR|1|10|Chus autem genuit Nemrod; iste coepit esse potens in terra.
1CHR|1|11|Mesraim vero genuit Ludim et Anamim et Laabim et Nephthuim,
1CHR|1|12|Phetrusim quoque et Chasluim, de quibus egressi sunt Philisthim e Caphtorim.
1CHR|1|13|Chanaan vero genuit Sidonem primogenitum, Heth,
1CHR|1|14|Iebusaeum quoque et Amorraeum et Gergesaeum
1CHR|1|15|Hevaeumque et Aracaeum et Sinaeum,
1CHR|1|16|Aradium quoque et Samaraeum et Emathaeum.
1CHR|1|17|Filii Sem: Elam et Assur et Arphaxad et Lud et Aram. Filii autem Aram: Us et Hul et Gether et Mes.
1CHR|1|18|Arphaxad autem genuit Sala, qui et ipse genuit Heber.
1CHR|1|19|Porro Heber nati sunt duo filii: nomen uni Phaleg, quia in diebus eius divisa est terra, et nomen fratris eius Iectan.
1CHR|1|20|Iectan autem genuit Elmodad et Saleph et Asarmoth et Iare,
1CHR|1|21|Adoram quoque et Uzal et Decla,
1CHR|1|22|Ebal etiam et Abimael et Saba necnon
1CHR|1|23|et Ophir et Hevila et Iobab; omnes isti filii Iectan.
1CHR|1|24|Sem, Arphaxad, Sala,
1CHR|1|25|Heber, Phaleg, Reu,
1CHR|1|26|Seruch, Nachor, Thare,
1CHR|1|27|Abram: iste est Abraham.
1CHR|1|28|Filii autem Abraham: Isaac et Ismael.
1CHR|1|29|Et hae generationes eorum: primogenitus Ismaelis Nabaioth et Cedar et Adbeel et Mabsam,
1CHR|1|30|Masma et Duma, Massa, Hadad et Thema,
1CHR|1|31|Iethur, Naphis, Cedma; hi sunt filii Ismaelis.
1CHR|1|32|Filii autem Ceturae concubinae Abraham, quos genuit: Zamran, Iecsan, Madan, Madian, Iesboc, Sue. Porro filii Iecsan: Saba et Dedan. Filii autem Dedan: Assurim et Latusim et Loommim.
1CHR|1|33|Filii autem Madian: Epha et Opher et Henoch et Abida et Eldaa. Omnes hi filii Ceturae.
1CHR|1|34|Generavit autem Abraham Isaac, cuius fuerunt filii Esau et Israel.
1CHR|1|35|Filii Esau: Eliphaz, Rahuel, Iehus, Ialam, Core.
1CHR|1|36|Filii Eliphaz: Theman, Omar, Sepho, Gatham, Cenez, Thamna, Amalec.
1CHR|1|37|Filii Rahuel: Nahath, Zara, Samma, Meza.
1CHR|1|38|Filii Seir: Lotan, Sobal, Sebeon, Ana, Dison, Eser, Disan.
1CHR|1|39|Filii Lotan: Hori, Hemam; soror autem Lotan fuit Thamna.
1CHR|1|40|Filii Sobal: Alvan et Manahath et Ebal et Sepho et Onam. Filii Sebeon: Aia et Ana.
1CHR|1|41|Filii Ana: Dison. Filii Dison: Hemdan et Eseban et Iethran et Charran.
1CHR|1|42|Filii Eser: Bilhan et Zavan et Iacan. Filii Disan: Us et Aran.
1CHR|1|43|Isti sunt reges, qui imperaverunt in terra Edom, antequam esset rex super filios Israel: Bela filius Beor, et nomen civitatis eius Denaba.
1CHR|1|44|Mortuus est autem Bela, et regnavit pro eo Iobab filius Zarae de Bosra.
1CHR|1|45|Cumque et Iobab fuisset mortuus, regnavit pro eo Husam de terra Themanorum.
1CHR|1|46|Obiit quoque et Husam, et regnavit pro eo Adad filius Badad, qui percussit Madian in terra Moab; et nomen civitatis eius Avith.
1CHR|1|47|Cumque et Adad fuisset mortuus, regnavit pro eo Semla de Masreca.
1CHR|1|48|Sed et Semla mortuus est; et regnavit pro eo Saul de Rohoboth, quae iuxta amnem sita est.
1CHR|1|49|Mortuo quoque Saul, regnavit pro eo Baalhanan filius Achobor.
1CHR|1|50|Sed et hic mortuus est, et regnavit pro eo Adad, cuius urbis fuit nomen Phau; et appellata est uxor eius Meetabel filia Matred filiae Mezaab.
1CHR|1|51|Adad autem mortuo, duces pro regibus in Edom esse coeperunt: dux Thamna, dux Alva, dux Ietheth,
1CHR|1|52|dux Oolibama, dux Ela, dux Phinon,
1CHR|1|53|dux Cenez, dux Theman, dux Mabsar,
1CHR|1|54|dux Magdiel, dux Iram. Hi duces Edom.
1CHR|2|1|Filii autem Israel: Ruben, Simeon, Levi, Iuda, Issachar et Zabulon,
1CHR|2|2|Dan, Ioseph, Beniamin, Nephthali, Gad, Aser.
1CHR|2|3|Filii Iudae: Her, Onan et Sela; hi tres nati sunt ei de filia Sue Chananitide. Fuit autem Her primogenitus Iudae malus coram Domino, et occidit eum.
1CHR|2|4|Thamar autem nurus eius peperit ei Phares et Zara; omnes ergo filii Iudae quinque.
1CHR|2|5|Filii autem Phares: Esrom et Hamul.
1CHR|2|6|Filii quoque Zarae: Zamri et Ethan et Heman, Chalchol quoque et Darda; simul quinque.
1CHR|2|7|Filii Charmi: Achar, qui turbavit Israel et peccavit in furto anathematis.
1CHR|2|8|Filii Ethan: Azarias.
1CHR|2|9|Filii autem Esrom, qui nati sunt ei: Ierameel et Aram et Chaleb.
1CHR|2|10|Porro Aram genuit Aminadab, Aminadab autem genuit Naasson principem filiorum Iudae,
1CHR|2|11|Naasson quoque genuit Salmon, de quo ortus est Booz.
1CHR|2|12|Booz vero genuit Obed, qui et ipse genuit Isai.
1CHR|2|13|Isai autem genuit primogenitum Eliab, secundum Abinadab, tertium Samma,
1CHR|2|14|quartum Nathanael, quintum Raddai,
1CHR|2|15|sextum Asom, septimum David.
1CHR|2|16|Quorum sorores fuerunt: Sarvia et Abigail; filii Sarviae: Abisai, Ioab et Asael, tres.
1CHR|2|17|Abigail autem genuit Amasa, cuius pater fuit Iether Ismaelites.
1CHR|2|18|Chaleb vero filius Esrom genuit de uxore sua nomine Azuba, de qua nati sunt Ierioth, Ieser et Sobab et Ardon.
1CHR|2|19|Cumque mortua fuisset Azuba, accepit uxorem Chaleb Ephratha, quae peperit ei Hur.
1CHR|2|20|Porro Hur genuit Uri, et Uri genuit Beseleel.
1CHR|2|21|Post haec ingressus est Esrom ad filiam Machir patris Galaad et accepit eam, cum ipse esset annorum sexaginta; quae peperit ei Segub.
1CHR|2|22|Sed et Segub genuit Iair, qui possedit viginti tres civitates in terra Galaad.
1CHR|2|23|Cepitque Gesur et Aram oppida Iair ipsis et Canath et viculos eius sexaginta civitates. Omnes isti filii Machir patris Galaad.
1CHR|2|24|Cum autem mortuus esset Esrom, ingressus est Chaleb ad Ephratha uxorem Esrom patris sui. Habuit quoque Esrom uxorem Abia, quae peperit ei Ashur patrem Thecue.
1CHR|2|25|Nati sunt autem filii Ierameel primogeniti Esrom: Ram primogenitus eius et Buna et Aran et Asom et Ahia.
1CHR|2|26|Duxit quoque uxorem alteram Ierameel nomine Atara, quae fuit mater Onam.
1CHR|2|27|Sed et filii Ram primogeniti Ierameel fuerunt: Moos et Iamin et Acar.
1CHR|2|28|Onam autem habuit filios: Sammai et Iada. Filii autem Sammai: Nadab et Abisur.
1CHR|2|29|Nomen vero uxoris Abisur Abiail, quae peperit ei Ahobban et Molid.
1CHR|2|30|Filii autem Nadab fuerunt Saled et Apphaim; mortuus est autem Saled absque liberis.
1CHR|2|31|Filius vero Apphaim: Iesi, qui Iesi genuit Sesan; porro Sesan genuit Oholai.
1CHR|2|32|Filii autem Iada fratris Semmei: Iether et Ionathan; sed et Iether mortuus est absque liberis.
1CHR|2|33|Porro Ionathan genuit Phaleth et Ziza. Isti fuerunt filii Ierameel.
1CHR|2|34|Sesan autem non habuit filios sed filias et servum Aegyptium nomine Ieraa;
1CHR|2|35|deditque ei filiam suam uxorem, quae peperit ei Eththei.
1CHR|2|36|Eththei autem genuit Nathan, et Nathan genuit Zabad;
1CHR|2|37|Zabad quoque genuit Ophlal, et Ophlal genuit Obed.
1CHR|2|38|Obed genuit Iehu, Iehu genuit Azariam;
1CHR|2|39|Azarias genuit Helles, Helles genuit Elasa.
1CHR|2|40|Elasa genuit Sisamoi, Sisamoi genuit Sellum;
1CHR|2|41|Sellum genuit Iecemiam, Iecemias genuit Elisama.
1CHR|2|42|Filii autem Chaleb fratris Ierameel: Mesa primogenitus eius, ipse est pater Ziph; et filius eius Maresa pater Hebron.
1CHR|2|43|Porro filii Hebron: Core et Thapphua et Recem et Samma;
1CHR|2|44|Samma autem genuit Raham patrem Iercaam, et Recem genuit Sammai.
1CHR|2|45|Filius Sammai: Maon, et Maon pater Bethsur.
1CHR|2|46|Epha autem concubina Chaleb peperit Charran et Mosa et Gezez; porro Charran genuit Gezez.
1CHR|2|47|Filii Iahaddai: Regem et Iotham et Gesan et Phalet et Epha et Saaph.
1CHR|2|48|Concubina Chaleb Maacha peperit Saber et Tharana.
1CHR|2|49|Genuit autem Saaph pater Madmena Sue patrem Machbena et patrem Gabaa. Filia vero Chaleb fuit Achsa.
1CHR|2|50|Hi erant filii Chaleb.Filii Hur primogeniti Ephratha: Sobal pater Cariathiarim,
1CHR|2|51|Salmon pater Bethlehem, Hariph pater Bethgader.
1CHR|2|52|Fuerunt autem filii Sobal patris Cariathiarim Raaia, dimidium Manahat
1CHR|2|53|et cognationes Cariathiarim: Iethraei et Phutaei et Sumathaei et Maseraei. Ex his egressi sunt Saraitae et Esthaolitae.
1CHR|2|54|Filii Salmon: Bethlehem et Netophathitae, Atarothbethioab et dimidium Manahat de Saraa,
1CHR|2|55|cognationes quoque de Cariathsepher habitantes in Iabes: Therathaei, Semathaei et Suchathaei. Hi sunt Cinaei, qui orti sunt de Ammath patre domus Rechab.
1CHR|3|1|David vero hos habuit filios, qui ei nati sunt in Hebron: primoge nitum Amnon ex Achinoam Iezrahelitide, secundum Daniel de Abigail de Carmel,
1CHR|3|2|tertium Absalom filium Maacha filiae Tholmai regis Gesur, quartum Adoniam filium Haggith,
1CHR|3|3|quintum Saphatiam ex Abital, sextum Iethraam de Egla uxore sua.
1CHR|3|4|Sex ergo nati sunt ei in Hebron, ubi regnavit septem annis et sex mensibus. Triginta autem et tribus annis regnavit in Ierusalem.
1CHR|3|5|Porro in Ierusalem nati sunt ei filii: Samua et Sobab et Nathan et Salomon, quattuor de Bethsabee filia Ammiel;
1CHR|3|6|Iebahar quoque et Elisama et Eliphalet
1CHR|3|7|et Noga et Napheg et Iaphia
1CHR|3|8|necnon Elisama et Eliada et Eliphalet, novem.
1CHR|3|9|Omnes hi filii David absque filiis concubinarum; habueruntque sororem Thamar.
1CHR|3|10|Filius autem Salomonis Roboam, cuius Abia filius genuit Asa; de hoc quoque natus est Iosaphat
1CHR|3|11|pater Ioram; qui Ioram genuit Ochoziam, ex quo ortus est Ioas.
1CHR|3|12|Et huius Amasias filius genuit Azariam, porro Azariae filius Ioatham
1CHR|3|13|procreavit Achaz patrem Ezechiae, de quo natus est Manasses.
1CHR|3|14|Sed et Manasses genuit Amon patrem Iosiae;
1CHR|3|15|filii autem Iosiae fuerunt: primogenitus Iohanan, secundus Ioachim, tertius Sedecias, quartus Sellum.
1CHR|3|16|Filii Ioachim: Iechonias filius eius, Sedecias filius eius.
1CHR|3|17|Filii Iechoniae captivi fuerunt: Salathiel filius eius,
1CHR|3|18|Melchiram, Phadaia, Senasser et Iecemias, Hosama et Nadabias.
1CHR|3|19|De Phadaia orti sunt Zorobabel et Semei. Zorobabel genuit Mosollam, Hananiam et Salomith sororem eorum
1CHR|3|20|Hasabamque et Ohol et Barachiam et Hasadiam, Iosabhesed, quinque.
1CHR|3|21|Filii autem Hananiae: Pheltias, Iesaias, Raphaia, Arnan, Abdia et Sechenias.
1CHR|3|22|Filii Secheniae: Semeia et Hattus et Igal et Baria et Naaria et Saphat, sex numero.
1CHR|3|23|Filii Naariae: Elioenai et Ezechias et Ezricam, tres.
1CHR|3|24|Filii Elioenai: Odovia et Eliasib et Pheleia et Accub et Iohanan et Dalaia et Anani, septem.
1CHR|4|1|Filii Iudae: Phares, Esrom et Charmi et Hur et Sobal.
1CHR|4|2|Reaia vero filius Sobal genuit Iahath, de quo nati sunt Ahumai et Laad; hae cognationes Saraitarum.
1CHR|4|3|Et ista stirps Etam: Iezrahel et Iesema et Iedebos, nomenque sororis eorum Asalelphuni.
1CHR|4|4|Phanuel autem pater Gedor et Ezer pater Hosa; isti sunt filii Hur primogeniti Ephratha patris Bethlehem.
1CHR|4|5|Ashur vero patris Thecue erant duae uxores: Halaa et Naara.
1CHR|4|6|Peperit autem ei Naara Oozam et Hepher et Themani et Ahasthari; isti sunt filii Naara.
1CHR|4|7|Porro filii Halaa: Sereth et Sohar et Ethnan.
1CHR|4|8|Cos autem genuit Anob et Sobeba et cognationes Aharehel filii Arum.
1CHR|4|9|Fuit autem Iabes inclitus prae fratribus suis; et mater eius vocavit nomen illius Iabes dicens: " Quia peperi eum in dolore ".
1CHR|4|10|Invocavit vero Iabes Deum Israel dicens: " Si benedicens benedixeris mihi et dilataveris terminos meos, et fuerit manus tua mecum, et feceris me a malitia non opprimi! ". Et praestitit Deus quae precatus est.
1CHR|4|11|Chelub autem frater Suaa genuit Mahir, qui fuit pater Esthon.
1CHR|4|12|Porro Esthon genuit Bethrapha et Phasea et Tehinna patrem Hirnaas (id est urbis Naas); hi sunt viri Recha.
1CHR|4|13|Filii autem Cenez: Othoniel et Saraia; porro filii Othoniel: Hathath et Maonathi.
1CHR|4|14|Maonathi genuit Ophra, Saraia autem genuit Ioab patrem Geharasim (id est vallis Artificum); ibi quippe artifices erant.
1CHR|4|15|Filii vero Chaleb filii Iephonne: Hir et Ela et Naham; filius quoque Ela: Cenez.
1CHR|4|16|Filii quoque Iallelel: Ziph et Zipha, Thiria et Asarel.
1CHR|4|17|Et filii Ezra: Iether et Mered et Epher et Ialon. Et genuit Iether Mariam et Sammai et Iesba patrem Esthemo.
1CHR|4|18|Hi autem sunt filii Bethiae filiae pharaonis, quam accepit Mered.
1CHR|4|19|Filii autem uxoris eius Iudaicae sororis Naham patris Ceilae: Dalaia et Simeon pater Ioman. Filii autem Naham patris Ceilae: Garmitae et Esthemo Maachathitarum.
1CHR|4|20|Filii quoque Simon: Ammon et Rinna, Benhanan et Thilon. Et filii Iesi: Zoheth et Benzoheth.
1CHR|4|21|Filii Sela filii Iudae: Her pater Lecha et Laada pater Maresa et cognationes domus operantium byssum in Bethasbea
1CHR|4|22|et Iochim virique Chozeba et Ioas et Saraph, qui principes fuerunt in Moab et qui reversi sunt in Bethlehem; hae autem sunt res veteres.
1CHR|4|23|Hi sunt figuli habitantes Netaim et Gedera; apud regem in operibus eius commorati sunt ibi.
1CHR|4|24|Filii Simeon: Namuel et Iamin, Iarib, Zara, Saul;
1CHR|4|25|Sellum filius eius, Mabsam filius eius, Masma filius eius.
1CHR|4|26|Filii Masma: Hamuel filius eius, Zacchur filius eius, Semei filius eius.
1CHR|4|27|Filii Semei sedecim et filiae sex; fratres autem eius non habuerunt filios multos, et universa cognatio eorum non potuit adaequare summam filiorum Iudae.
1CHR|4|28|Habitaverunt autem in Bersabee et Molada et Asarsual
1CHR|4|29|et in Bilha et in Esem et in Tholad
1CHR|4|30|et in Bathuel et in Horma et in Siceleg
1CHR|4|31|et in Bethmarchaboth et in Asarsusim et in Bethberai et in Saarim; hae civitates eorum usque ad regem David.
1CHR|4|32|Villae quoque eorum: Etam et Ain, Remmon et Thochen et Asan, civitates quinque.
1CHR|4|33|Et universi viculi eorum per circuitum civitatum istarum usque ad Baal; haec est habitatio eorum et genealogia.
1CHR|4|34|Masobab quoque et Iemlech et Iosa filius Amasiae
1CHR|4|35|et Ioel et Iehu filius Iosabiae filii Saraiae filii Asiel
1CHR|4|36|et Elioenai et Iacoba et Isuhaia et Asaia et Adiel et Isimiel et Banaia,
1CHR|4|37|Ziza quoque filius Sephei filii Allon filii Iedaia filii Semri filii Samaia.
1CHR|4|38|Isti nominatim inscripti erant principes in cognationibus suis; et familiae eorum expansae sunt vehementer,
1CHR|4|39|et profecti sunt ad introitum Gedor usque ad orientem vallis, ut quaererent pascua gregibus suis.
1CHR|4|40|Inveneruntque pascuas uberes et valde bonas et terram latissimam et quietam et fertilem, in qua ante habitaverunt de stirpe Cham.
1CHR|4|41|Hi ergo venerunt, qui inscripti erant nominatim, in diebus Ezechiae regis Iudae, et percusserunt tabernacula eorum et Meunitas, qui inventi fuerunt ibi, et deleverunt eos usque in praesentem diem habitaveruntque pro eis, quoniam uberrimas ibidem pascuas reppererunt.
1CHR|4|42|De filiis quoque Simeon abierunt in montem Seir viri quingenti habentes principes Pheltiam et Naariam et Raphaiam et Oziel filios Iesi
1CHR|4|43|et percusserunt reliquias, quae evadere potuerant Amalecitarum, et habitaverunt ibi pro eis usque ad diem hanc.
1CHR|5|1|Filii quoque Ruben primogeniti Israel: ipse quippe fuit primoge nitus eius, sed, cum violasset torum patris sui, data sunt primogenita eius filiis Ioseph filii Israel, ut non computaretur in primogenitum,
1CHR|5|2|quia Iuda erat quidem fortissimus inter fratres suos et de stirpe eius principes germinati sunt, primogenita autem reputata sunt Ioseph.
1CHR|5|3|Filii ergo Ruben primogeniti Israel: Henoch et Phallu, Hesron et Charmi.
1CHR|5|4|Filii Ioel: Semeia filius eius, Gog filius eius, Semei filius eius,
1CHR|5|5|Micha filius eius, Reaia filius eius, Baal filius eius,
1CHR|5|6|Beera filius eius, quem captivum duxit Theglathphalasar rex Assyriorum, et fuit princeps in tribu Ruben.
1CHR|5|7|Fratres autem eius in cognationibus eius, quando numerabantur in genealogiis suis, erant: caput Iehiel, deinde Zacharias;
1CHR|5|8|porro Bela filius Azaz filii Samma filii Ioel, ipse habitavit in Aroer usque ad Nabo et Baalmeon.
1CHR|5|9|Contra orientalem quoque plagam habitavit usque ad introitum eremi, quae est inde a flumine Euphrate; multum quippe gregum eorum numerus creverat in terra Galaad.
1CHR|5|10|In diebus autem Saul proeliati sunt contra Agarenos et interfecerunt illos; habitaveruntque pro eis in tabernaculis eorum in omni plaga, quae respicit ad orientem Galaad.
1CHR|5|11|Filii vero Gad e regione eorum habitaverunt in terra Basan usque Salcha:
1CHR|5|12|Ioel in capite et Sapham secundus, porro Ianai et Saphat in Basan;
1CHR|5|13|fratres vero eorum secundum familias suas: Michael et Mosollam et Seba et Iorai et Iachan et Zie et Heber, septem.
1CHR|5|14|Hi filii Abihail filii Huri filii Iaroe filii Galaad filii Michael filii Iesesi filii Ieddo filii Buz.
1CHR|5|15|Ahi filius Abdiel filii Guni princeps familiarum eorum.
1CHR|5|16|Et habitaverunt in Galaad et in Basan et in viculis eius et in cunctis suburbanis Saron usque ad terminos.
1CHR|5|17|Omnes hi numerati sunt in diebus Ioatham regis Iudae et in diebus Ieroboam regis Israel.
1CHR|5|18|Filii Ruben et Gad et dimidiae tribus Manasse viri bellatores scuta portantes et gladios et tendentes arcum eruditique ad proelia, quadraginta quattuor milia et septingenti sexaginta procedentes ad pugnam;
1CHR|5|19|dimicaverunt contra Agarenos et Ituraeos et Naphisaeos et Nodabaeos.
1CHR|5|20|Et datum est eis auxilium, traditique sunt in manus eorum Agareni et universi, qui fuerant cum eis, quia Deum invocaverunt cum proeliarentur, et exaudivit eos, eo quod credidissent in eum.
1CHR|5|21|Ceperuntque omnia, quae possederant, camelorum quinquaginta milia et ovium ducenta quinquaginta milia, asinos duo milia et animas hominum centum milia;
1CHR|5|22|vulnerati autem multi corruerunt; fuit enim bellum Domini. Habitaveruntque pro eis usque ad transmigrationem.
1CHR|5|23|Filii quoque dimidiae tribus Manasse possederunt terram a Basan usque Baalhermon et Sanir et montem Hermon; ingens quippe numerus erat.
1CHR|5|24|Et hi fuerunt principes familiarum eorum: Epher et Iesi et Eliel et Azriel et Ieremia et Odovia et Iediel; viri bellatores fortissimi et nominati, duces in familiis suis.
1CHR|5|25|Reliquerunt autem Deum patrum suorum et fornicati sunt post deos populorum terrae, quos abstulit Deus coram eis.
1CHR|5|26|Et suscitavit Deus Israel spiritum Phul regis Assyriorum et spiritum Theglathphalasar regis Assur; et transtulit Ruben et Gad et dimidium tribus Manasse et adduxit eos in Hala et Habor et Ara et fluvium Gozan usque ad diem hanc.
1CHR|5|27|Filii Levi: Gerson, Caath, Merari.
1CHR|5|28|Filii Caath: Amram, Isaar, Hebron et Oziel.
1CHR|5|29|Filii Amram: Aaron, Moyses et Maria. Filii Aaron: Nadab et Abiu, Eleazar et Ithamar.
1CHR|5|30|Eleazar genuit Phinees, et Phinees genuit Abisue;
1CHR|5|31|Abisue vero genuit Bocci, et Bocci genuit Ozi.
1CHR|5|32|Ozi genuit Zaraiam, et Zaraias genuit Meraioth,
1CHR|5|33|porro Meraioth genuit Amariam, et Amarias genuit Achitob;
1CHR|5|34|Achitob genuit Sadoc, Sadoc genuit Achimaas,
1CHR|5|35|Achimaas genuit Azariam, Azarias genuit Iohanan;
1CHR|5|36|Iohanan genuit Azariam: ipse est qui sacerdotio functus est in domo, quam aedificavit Salomon in Ierusalem.
1CHR|5|37|Genuit autem Azarias Amariam, et Amarias genuit Achitob,
1CHR|5|38|Achitob genuit Sadoc, et Sadoc genuit Sellum;
1CHR|5|39|Sellum genuit Helciam, et Helcias genuit Azariam.
1CHR|5|40|Azarias genuit Saraiam, et Saraias genuit Iosedec;
1CHR|5|41|porro Iosedec egressus est, quando transtulit Dominus Iudam et Ierusalem per manus Nabuchodonosor.
1CHR|6|1|Filii ergo Levi: Gerson, Caath et Merari.
1CHR|6|2|Et haec nomina filio rum Gerson: Lobni et Semei.
1CHR|6|3|Filii Caath: Amram et Isaar et Hebron et Oziel.
1CHR|6|4|Filii Merari: Moholi et Musi.Hae autem cognationes Levi secundum familias eorum:
1CHR|6|5|Gerson, Lobni filius eius, Iahath filius eius, Zimma filius eius,
1CHR|6|6|Ioah filius eius, Addo filius eius, Zara filius eius, Iethrai filius eius.
1CHR|6|7|Filii Caath: Aminadab filius eius, Core filius eius, Asir filius eius,
1CHR|6|8|Elcana filius eius, Abiasaph filius eius, Asir filius eius,
1CHR|6|9|Thahath filius eius, Uriel filius eius, Ozias filius eius, Saul filius eius.
1CHR|6|10|Filii Elcana: Amasai et Achimoth,
1CHR|6|11|Elcana filius eius, Sophai filius eius, Nahath filius eius,
1CHR|6|12|Eliab filius eius, Ieroham filius eius, Elcana filius eius, Samuel filius eius.
1CHR|6|13|Filii Samuel: primogenitus Ioel et secundus Abia.
1CHR|6|14|Filii autem Merari: Moholi, Lobni filius eius, Semei filius eius, Oza filius eius,
1CHR|6|15|Samaa filius eius, Haggia filius eius, Asaia filius eius.
1CHR|6|16|Isti sunt, quos constituit David super cantum domus Domini, ex quo collocata est arca;
1CHR|6|17|et ministrabant coram habitatione tabernaculi conventus canentes, donec aedificaret Salomon domum Domini in Ierusalem; stabant autem iuxta ordinem suum in ministerio.
1CHR|6|18|Hi vero sunt, qui assistebant cum filiis suis. De filiis Caath: Heman cantor filius Ioel filii Samuel
1CHR|6|19|filii Elcana filii Ieroham filii Eliel filii Thohu
1CHR|6|20|filii Suph filii Elcana filii Mahath filii Amasai
1CHR|6|21|filii Elcana filii Ioel filii Azariae filii Sophoniae
1CHR|6|22|filii Thahath filii Asir filii Abiasaph filii Core
1CHR|6|23|filii Isaar filii Caath filii Levi filii Israel.
1CHR|6|24|Et frater eius Asaph, qui stabat a dextris eius, Asaph filius Barachiae filii Samaa
1CHR|6|25|filii Michael filii Basaiae filii Melchiae
1CHR|6|26|filii Athnai filii Zara filii Adaia
1CHR|6|27|filii Ethan filii Zimma filii Semei
1CHR|6|28|filii Iahath filii Gerson filii Levi.
1CHR|6|29|Filii autem Merari fratres eorum ad sinistram: Ethan filius Cusi filii Abdi filii Melluch
1CHR|6|30|filii Hasabiae filii Amasiae filii Helciae
1CHR|6|31|filii Amsi filii Bani filii Somer
1CHR|6|32|filii Moholi filii Musi filii Merari filii Levi.
1CHR|6|33|Fratres quoque eorum Levitae, qui ordinati sunt in cunctum ministerium habitaculi domus Domini;
1CHR|6|34|Aaron vero et filii eius adolebant super altare holocausti et super altare thymiamatis in omne opus sancti sanctorum, et ut expiarent pro Israel, iuxta omnia quae praecepit Moyses servus Dei.
1CHR|6|35|Hi sunt autem filii Aaron: Eleazar filius eius, Phinees filius eius, Abisue filius eius,
1CHR|6|36|Bocci filius eius, Ozi filius eius, Zaraia filius eius,
1CHR|6|37|Meraioth filius eius, Amarias filius eius, Achitob filius eius,
1CHR|6|38|Sadoc filius eius, Achimaas filius eius.
1CHR|6|39|Et haec habitacula eorum per castra atque confinia, filiorum scilicet Aaron ex cognatione Caathitarum; ipsis enim sorte contigerat.
1CHR|6|40|Dederunt igitur eis Hebron in terra Iudae et suburbana eius per circuitum;
1CHR|6|41|agros autem civitatis et villas Chaleb filio Iephonne.
1CHR|6|42|Porro filiis Aaron dederunt civitatem ad confugiendum: Hebron et Lobna et suburbana eius,
1CHR|6|43|Iether quoque et Esthemo cum suburbanis eius, sed et Helon et Dabir cum suburbanis suis,
1CHR|6|44|Asan quoque et Iutta et Bethsames et suburbana earum;
1CHR|6|45|de tribu autem Beniamin: Gabaon et Gabaa et suburbana earum et Almath cum suburbanis suis, Anathoth quoque cum suburbanis suis: omnes civitates tredecim, singulae per cognationes suas.
1CHR|6|46|Filiis autem Caath residuis de cognatione sua dederunt ex tribu Ephraim et ex tribu Dan et ex dimidia tribu Manasse in possessionem urbes decem.
1CHR|6|47|Porro filiis Gerson per cognationes suas de tribu Issachar et de tribu Aser et de tribu Nephthali et de tribu Manasse in Basan urbes tredecim.
1CHR|6|48|Filiis autem Merari per cognationes suas de tribu Ruben et de tribu Gad et de tribu Zabulon dederunt sorte civitates duodecim.
1CHR|6|49|Dederunt quoque filii Israel Levitis civitates et suburbana earum;
1CHR|6|50|dederuntque per sortem ex tribu filiorum Iudae et ex tribu filiorum Simeon et ex tribu filiorum Beniamin urbes has, quas vocaverunt nominibus suis.
1CHR|6|51|Et his, qui erant ex cognationibus filiorum Caath, fuerunt civitates in terminis eorum de tribu Ephraim.
1CHR|6|52|Dederunt ergo eis urbem ad confugiendum: Sichem cum suburbanis suis in monte Ephraim et Gazer cum suburbanis suis,
1CHR|6|53|Iecmaam quoque cum suburbanis suis et Bethoron similiter;
1CHR|6|54|necnon et Aialon cum suburbanis suis et Gethremmon in eundem modum.
1CHR|6|55|Porro ex dimidia tribu Manasse Thanach et suburbana eius, Ieblaam et suburbana eius, his videlicet qui de cognationibus filiorum Caath reliqui erant.
1CHR|6|56|Filiis autem Gerson de cognationibus dimidiae tribus Manasse: Golan in Basan et suburbana eius et Astharoth cum suburbanis suis.
1CHR|6|57|De tribu Issachar Cedes et suburbana illius et Dabereth cum suburbanis suis,
1CHR|6|58|Ramoth quoque et suburbana illius et Anem cum suburbanis suis.
1CHR|6|59|De tribu vero Aser: Masal cum suburbanis suis et Abdon similiter,
1CHR|6|60|Hucoc quoque et suburbana eius et Rohob cum suburbanis suis.
1CHR|6|61|Porro de tribu Nephthali: Cedes in Galilaea et suburbana eius, Hamon cum suburbanis suis et Cariathaim et suburbana eius.
1CHR|6|62|Filiis autem Merari residuis de tribu Zabulon: Remmon et suburbana eius et Thabor cum suburbanis suis.
1CHR|6|63|Trans Iordanem quoque ex adverso Iericho, contra orientem Iordanis de tribu Ruben: Bosor in solitudine cum suburbanis suis et Iasa cum suburbanis suis,
1CHR|6|64|Cademoth quoque et suburbana eius et Mephaath cum suburbanis suis.
1CHR|6|65|Necnon et de tribu Gad: Ramoth in Galaad et suburbana eius et Mahanaim cum suburbanis suis,
1CHR|6|66|sed et Hesebon cum suburbanis eius, et Iazer cum suburbanis suis.
1CHR|7|1|Porro filii Issachar: Thola et Phua, Iasub et Semron, quat tuor.
1CHR|7|2|Filii Thola: Ozi et Raphaia et Ieriel et Iemai et Iebsem et Samuel, principes familiarum suarum; de stirpe Thola viri fortissimi numerati sunt iuxta genealogias suas in diebus David viginti duo milia sescenti.
1CHR|7|3|Filii Ozi: Izrahia, de quo nati sunt Michael et Obadia et Ioel et Iesia, quinque principes omnes.
1CHR|7|4|Cumque eis erant secundum genealogias familiarum suarum turmae accinctae ad proelium, viri fortissimi, triginta sex milia; multas enim habuere uxores et filios.
1CHR|7|5|Fratresque eorum per omnes cognationes Issachar robustissimi ad pugnandum octoginta septem milia numerati sunt.
1CHR|7|6|Filii Beniamin: Bela et Bochor et Iedihel, tres.
1CHR|7|7|Filii Bela: Esebon et Ozi et Oziel et Ierimoth et Urai, quinque principes familiarum et ad pugnandum robustissimi; numerus autem eorum viginti duo milia et triginta quattuor.
1CHR|7|8|Porro filii Bochor: Zamira et Ioas et Eliezer et Elioenai et Amri et Ierimoth et Abia et Anathoth et Almath; omnes hi filii Bochor.
1CHR|7|9|Numerati sunt autem in genealogiis suis principes familiarum suarum ad bella fortissimi viginti milia et ducenti.
1CHR|7|10|Porro filii Iedihel: Bilhan; filii autem Bilhan: Iehus et Beniamin et Aod et Chanaana et Zethan et Tharsis et Ahisahar;
1CHR|7|11|omnes hi filii Iedihel principes familiarum suarum viri fortissimi decem et septem milia et ducenti ad proelium procedentes.
1CHR|7|12|Suphim quoque et Huphim filii Hir et Husim filii Aher.
1CHR|7|13|Filii autem Nephthali: Iasiel et Guni et Ieser et Sellum, filii Bilhae.
1CHR|7|14|Porro filius Manasse: Asriel, quem peperit concubina eius Syra; peperit quoque Machir patrem Galaad.
1CHR|7|15|Machir autem accepit uxorem de Huphim et Suphim et habuit sororem nomine Maacha; nomen autem secundi Salphaad, nataeque sunt Salphaad filiae.
1CHR|7|16|Et peperit Maacha uxor Machir filium vocavitque nomen eius Phares; porro nomen fratris eius Sares et filii eius Ulam et Recem.
1CHR|7|17|Filius autem Ulam: Badan; hi sunt filii Galaad filii Machir filii Manasse.
1CHR|7|18|Soror autem eius Ammalecheth peperit Isod et Abiezer et Maala.
1CHR|7|19|Erant autem filii Semida: Ahin et Sechem et Leci et Aniam.
1CHR|7|20|Filii autem Ephraim: Suthala, Bared filius eius, Thahath filius eius, Elada filius eius, Thahath filius eius,
1CHR|7|21|et huius filius Zabad et huius filius Suthala et huius filius Ezer et Elad. Occiderunt autem eos viri Geth indigenae, quia descenderant, ut invaderent possessiones eorum.
1CHR|7|22|Luxit igitur Ephraim pater eorum multis diebus, et venerunt fratres eius, ut consolarentur eum;
1CHR|7|23|ingressusque est ad uxorem suam, quae concepit et peperit filium, et vocavit nomen eius Beria, eo quod in malis domus eius ortus esset.
1CHR|7|24|Filia autem eius fuit Sara, quae aedificavit Bethoron inferiorem et superiorem et Ozensara.
1CHR|7|25|Porro filius eius Rapha et Reseph et Thale filius eius, de quo natus est Thaan,
1CHR|7|26|qui genuit Laadan; huius quoque filius Ammiud genuit Elisama,
1CHR|7|27|de quo ortus est Nun, qui habuit filium Iosue.
1CHR|7|28|Possessio autem eorum et habitationes: Bethel cum filiabus suis et contra orientem Noran, ad occidentalem plagam Gazer et filiae eius, Sichem quoque cum filiabus suis usque Hai et filias eius.
1CHR|7|29|Iuxta filios quoque Manasse: Bethsan et filias eius, Thanach et filias eius, Mageddo et filias eius, Dor et filias eius. In his habitaverunt filii Ioseph filii Israel.
1CHR|7|30|Filii Aser: Iemna et Iesua et Isui et Beria et Sara soror eorum.
1CHR|7|31|Filii autem Beria: Heber et Melchiel, ipse est pater Barzaith.
1CHR|7|32|Heber autem genuit Iephlat et Somer et Hotham et Suaa sororem eorum.
1CHR|7|33|Filii Iephlat: Phosech et Bamaal et Asoth; hi filii Iephlat.
1CHR|7|34|Porro filii Somer fratris sui: Roaga et Haba et Aram.
1CHR|7|35|Filii autem Hotham fratris eius: Supha et Iemna et Selles et Amal.
1CHR|7|36|Filii Supha: Sue, Hamapher et Sual et Beri et Iamra,
1CHR|7|37|Bosor et Od et Samma et Salusa et Iethran et Beera.
1CHR|7|38|Filii Iether: Iephonne et Phaspha et Ara.
1CHR|7|39|Filii autem Olla: Area et Hanniel et Resia.
1CHR|7|40|Omnes hi filii Aser, principes familiarum electi atque fortissimi, capita principum; numerus autem eorum, qui inscripti erant in exercitu ad bellum, viginti sex milia.
1CHR|8|1|Beniamin autem genuit Bela primogenitum suum, Asbel se cundum, Ahara tertium,
1CHR|8|2|Nohaa quartum et Rapha quintum.
1CHR|8|3|Fueruntque filii Bela: Addar et Gera pater Aod,
1CHR|8|4|Abisue quoque et Naaman et Ahoe,
1CHR|8|5|sed et Gera et Sephuphan et Huram.
1CHR|8|6|Hi sunt filii Aod principes familiarum habitantium in Gabaa, qui translati sunt in Manahath;
1CHR|8|7|Naaman autem et Ahia et Gera: ipse transtulit eos et genuit Oza et Ahiud.
1CHR|8|8|Porro Saharaim genuit in regione Moab, postquam dimisit Husim et Bara uxores suas;
1CHR|8|9|genuit autem de Hodes uxore sua Iobab et Sebia et Mesa et Melcham,
1CHR|8|10|Iehus quoque et Sechia et Marma; hi sunt filii eius principes in familiis suis.
1CHR|8|11|De Husim vero genuit Abitob et Elphaal;
1CHR|8|12|porro filii Elphaal Heber et Misaam et Samad; hic aedificavit Ono et Lod et filias eius.
1CHR|8|13|Beria autem et Samma principes familiarum habitantium in Aialon; hi fugaverunt habitatores Geth.
1CHR|8|14|Et Ahi et Sesac et Ierimoth
1CHR|8|15|et Zabadia et Arad et Eder,
1CHR|8|16|Michael quoque et Iespha et Ioha filii Beria.
1CHR|8|17|Et Zabadia et Mosollam et Hezeci et Heber
1CHR|8|18|et Iesamari et Iezlia et Iobab filii Elphaal
1CHR|8|19|et Iacim et Zechri et Zabdi
1CHR|8|20|et Elioenai et Selethai et Eliel
1CHR|8|21|et Adaia et Baraia et Samarath filii Semei
1CHR|8|22|et Iesphan et Heber et Eliel
1CHR|8|23|et Abdon et Zechri et Hanan
1CHR|8|24|et Hanania et Elam et Anathothia
1CHR|8|25|et Iephdaia et Phanuel filii Sesac.
1CHR|8|26|Et Samsari et Sohoria et Otholia
1CHR|8|27|et Iersia et Elia et Zechri filii Ieroham.
1CHR|8|28|Hi capita familiarum secundum genealogias, principes qui habitaverunt in Ierusalem.
1CHR|8|29|In Gabaon autem habitaverunt Iehiel pater Gabaon, et nomen uxoris eius Maacha,
1CHR|8|30|filiusque eius primogenitus Abdon et Sur et Cis et Baal et Ner et Nadab,
1CHR|8|31|Gedor quoque et Ahio et Zacher et Macelloth;
1CHR|8|32|et Macelloth genuit Samaa. Habitaveruntque ex adverso fratrum suorum in Ierusalem cum fratribus suis.
1CHR|8|33|Ner autem genuit Cis, et Cis genuit Saul. Porro Saul genuit Ionathan et Melchisua et Abinadab et Isbaal.
1CHR|8|34|Filius autem Ionathan Meribbaal, et Meribbaal genuit Micha;
1CHR|8|35|filii Micha Phithon et Melech et Tharaa et Ahaz.
1CHR|8|36|Et Ahaz genuit Ioada, et Ioada genuit Almath et Azmaveth et Zamri; porro Zamri genuit Mosa.
1CHR|8|37|Et Mosa genuit Banaa, cuius filius fuit Raphaia, de quo ortus est Elasa, qui genuit Asel.
1CHR|8|38|Porro Asel sex filii fuere his nominibus: Ezricam primogenitus eius, Ismael, Saria, Azarias, Obdia et Hanan; omnes hi filii Asel.
1CHR|8|39|Filii autem Esec fratris eius: Ulam primogenitus et Iehus secundus et Eliphalet tertius.
1CHR|8|40|Fueruntque filii Ulam viri robustissimi ad bellum et magno robore tendentes arcum et multos habentes filios ac nepotes usque ad centum quinquaginta. Omnes hi filii Beniamin.
1CHR|9|1|Universus ergo Israel dinume ratus est, et summa eorum scrip ta est in libro regum Israel et Iudae. Translatique sunt in Babylonem propter delictum suum.
1CHR|9|2|Qui autem habitaverunt primi in possessionibus et in urbibus suis: Israel et sacerdotes et Levitae et Nathinaei.
1CHR|9|3|Commorati sunt in Ierusalem de filiis Iudae et de filiis Beniamin, de filiis quoque Ephraim et Manasse.
1CHR|9|4|Uthai filius Ammiud filii Amri filii Imri filii Bani: de filiis Phares filii Iudae;
1CHR|9|5|et de Selanitis: Asaia primogenitus et filii eius;
1CHR|9|6|de filiis autem Zara: Iehuel et fratres eorum sescenti nonaginta.
1CHR|9|7|Porro de filiis Beniamin: Sallu filius Mosollam filii Odovia filii Asana
1CHR|9|8|et Iobania filius Ieroham et Ela filius Ozi filii Mochori et Mosollam filius Saphatiae filii Rahuel filii Iebaniae
1CHR|9|9|et fratres eorum secundum genealogias suas nongenti quinquaginta sex; omnes hi principes familiarum secundum familias suas.
1CHR|9|10|De sacerdotibus autem: Iedaia, Ioiarib et Iachin,
1CHR|9|11|Azarias quoque filius Helciae filii Mosollam filii Sadoc filii Meraioth filii Achitob principes domus Dei.
1CHR|9|12|Porro Adaias filius Ieroham filii Phassur filii Melchiae et Maasai filius Adiel filii Iezra filii Mosollam filii Mosollamoth filii Emmer,
1CHR|9|13|fratres quoque eorum principes per familias suas mille septingenti sexaginta, fortissimi robore ad faciendum opus ministerii in domo Dei.
1CHR|9|14|De Levitis autem: Semeia filius Hassub filii Ezricam filii Hasabia de filiis Merari;
1CHR|9|15|Bacbacar quoque, Hares et Galal et Matthania filius Micha filii Zechri filii Asaph
1CHR|9|16|et Abdia filius Semeiae filii Galal filii Idithun et Barachia filius Asa filii Elcana, qui habitavit in atriis Netophathitarum.
1CHR|9|17|Ianitores autem: Sellum et Accub et Telmon et Ahiman; et frater eorum Sellum princeps
1CHR|9|18|et usque ad hoc tempus est in porta regis ad orientem. Hi erant ianitores castris filiorum Levi.
1CHR|9|19|Sellum vero filius Core filii Abiasaph filii Core cum fratribus suis de domo patris sui: hi Coritae erant super opera ministerii custodes liminum tabernaculi; patres autem eorum super castra Domini custodiebant introitum,
1CHR|9|20|et Phinees filius Eleazari princeps erat super eos olim - Dominus sit cum eo! -
1CHR|9|21|Zacharias filius Mosollamia ianitor portae tabernaculi conventus.
1CHR|9|22|Omnes hi electi in ostiarios liminum ducenti duodecim, et descripti in villis propriis, quos constituerunt David et Samuel videns in munus perpetuum,
1CHR|9|23|tam ipsos quam filios eorum in ostiis domus Domini, domus tabernaculi, in custodias.
1CHR|9|24|Per quattuor ventos erant ostiarii, id est ad orientem et ad occidentem, ad aquilonem et ad austrum.
1CHR|9|25|Fratres autem eorum in viculis suis morabantur et veniebant per septem dies de tempore usque ad tempus, ut essent cum illis.
1CHR|9|26|Nam munus habebant perpetuum hi quattuor principes ianitorum. Hi scilicet Levitae erant super exedras et thesauros domus Domini;
1CHR|9|27|per gyrum quoque templi Domini pernoctabant in custodiis suis, ut et ipsi mane aperirent fores.
1CHR|9|28|De horum genere erant et super vasa ministerii, ad numerum enim et inferebantur vasa et efferebantur;
1CHR|9|29|de ipsis et, qui credita habebant utensilia et omnia utensilia sancta, praeerant similae et vino et oleo et turi et aromatibus.
1CHR|9|30|Filii quidam autem sacerdotum unguenta ex aromatibus conficiebant;
1CHR|9|31|et Matthathias Levites, primogenitus Sellum Coritae, munere perpetuo praefectus erat eorum, quae in sartagine frigebantur.
1CHR|9|32|Porro de filiis Caath fratribus eorum super panes erant propositionis, ut semper novos per singula sabbata praepararent.
1CHR|9|33|Hi sunt cantores, principes per familias Levitarum, qui in exedris vacantes morabantur, ita ut die et nocte iugiter suo ministerio deservirent.
1CHR|9|34|Hi sunt capita Levitarum per familias suas secundum genealogias suas principes; hi habitaverunt in Ierusalem.
1CHR|9|35|In Gabaon autem commorati sunt pater Gabaon Iehiel, et nomen uxoris eius Maacha.
1CHR|9|36|Filius primogenitus eius Abdon et Sur et Cis et Baal et Ner et Nadab,
1CHR|9|37|Gedor quoque et Ahio et Zacharias et Macelloth.
1CHR|9|38|Porro Macelloth genuit Samaam; isti habitaverunt e regione fratrum suorum in Ierusalem cum fratribus suis.
1CHR|9|39|Ner autem genuit Cis, et Cis genuit Saul. Et Saul genuit Ionathan et Melchisua et Abinadab et Isbaal.
1CHR|9|40|Filius autem Ionathan Meribbaal, et Meribbaal genuit Micha;
1CHR|9|41|porro filii Micha: Phithon et Melech et Tharaa et Ahaz.
1CHR|9|42|Ahaz autem genuit Iara, et Iara genuit Almath et Azmaveth et Zamri; Zamri autem genuit Mosa.
1CHR|9|43|Mosa vero genuit Banaa, cuius filius Raphaia genuit Elasa, de quo ortus est Asel.
1CHR|9|44|Porro Asel sex filios habuit his nominibus: Ezricam primogenitus eius, Ismael, Saria, Azarias, Obdia, Hanan; hi filii Asel.
1CHR|10|1|Philisthim autem pugnabant contra Israel, fugeruntque viri Israel a facie Philisthim et ceciderunt vulnerati in monte Gelboe;
1CHR|10|2|cumque appropinquassent Philisthaei persequentes Saul et filios eius, percusserunt Ionathan et Abinadab et Melchisua filios Saul.
1CHR|10|3|Et aggravatum est proelium contra Saul, inveneruntque eum sagittarii et vulneraverunt iaculis;
1CHR|10|4|et dixit Saul ad armigerum suum: " Evagina gladium tuum et interfice me, ne forte veniant incircumcisi isti et illudant mihi ". Noluit autem armiger eius hoc facere timore perterritus. Arripuit igitur Saul ensem et irruit in eum;
1CHR|10|5|quod cum vidisset armiger eius, videlicet mortuum esse Saul, irruit etiam ipse in gladium suum et mortuus est.
1CHR|10|6|Interiit ergo Saul et tres filii eius; omnis domus illius pariter concidit.
1CHR|10|7|Quod cum vidissent omnes viri Israel, qui habitabant in campestribus, quod fugissent, et mortui essent Saul et filii eius, dereliquerunt urbes suas et huc illucque dispersi sunt; veneruntque Philisthim et habitaverunt in eis.
1CHR|10|8|Die igitur altero venerunt Philisthim, ut spoliarent interfectos, et invenerunt Saul et filios eius iacentes in monte Gelboe;
1CHR|10|9|cumque spoliassent eum et amputassent caput armisque nudassent, miserunt in terram suam per circuitum, ut annuntiaretur in idolorum templis et in populis.
1CHR|10|10|Arma autem eius consecraverunt in fano Astharoth et caput affixerunt in templo Dagon.
1CHR|10|11|Hoc cum audissent viri Iabes Galaad, omnia scilicet quae Philisthim fecerunt super Saul,
1CHR|10|12|consurrexerunt omnes viri fortes et tulerunt cadavera Saul et filiorum eius attuleruntque ea in Iabes et sepelierunt ossa eorum subter quercum, quae erat in Iabes, et ieiunaverunt septem diebus.
1CHR|10|13|Mortuus est ergo Saul propter iniquitatem suam, eo quod praevaricatus sit mandatum Domini, quod praeceperat, et non custodierit illud, sed insuper etiam pythonissam consuluerit
1CHR|10|14|nec quaesierit Dominum; propter quod et interfecit eum et transtulit regnum eius ad David filium Isai.
1CHR|11|1|Congregatus est igitur omnis Israel ad David in Hebron dicens: " Os tuum sumus et caro tua.
1CHR|11|2|Heri quoque et nudiustertius, cum adhuc regnaret Saul, tu eras qui educebas et introducebas Israel; tibi enim dixit Dominus Deus tuus: "Tu pasces populum meum Israel et tu eris princeps super eum" ".
1CHR|11|3|Venerunt ergo omnes maiores natu Israel ad regem in Hebron, et iniit David cum eis foedus in Hebron coram Domino; unxeruntque eum regem super Israel iuxta sermonem Domini, quem locutus est in manu Samuel.
1CHR|11|4|Abiit quoque David et omnis Israel in Ierusalem, haec est Iebus, ubi erant Iebusaei habitatores terrae.
1CHR|11|5|Dixeruntque, qui habitabant in Iebus, ad David: " Non ingredieris huc ". Porro David cepit arcem Sion, quae est civitas David;
1CHR|11|6|dixitque: " Omnis, qui percusserit Iebusaeum, in primis erit princeps et dux ". Ascendit igitur primus Ioab filius Sarviae et factus est princeps.
1CHR|11|7|Habitavit autem David in arce, et idcirco appellata est civitas David.
1CHR|11|8|Aedificavitque urbem in circuitu a Mello usque ad gyrum; Ioab autem reliqua urbis instauravit.
1CHR|11|9|Proficiebatque David vadens et crescens, et Dominus exercituum erat cum eo.
1CHR|11|10|Hi principes virorum fortium David, qui adiuverunt eum, ut rex fieret super omnem Israel iuxta verbum Domini, quod locutus est ad Israel;
1CHR|11|11|et iste numerus robustorum David: Iesbaam filius Hachamon filius Hachamonitis princeps inter triginta; iste levavit hastam suam super trecentos, quos occidit impetu uno.
1CHR|11|12|Et post eum Eleazar filius Dodo Ahohites, qui erat inter tres potentes;
1CHR|11|13|iste fuit cum David in Aphesdommim, quando Philisthim congregati sunt ad locum illum in proelium. Et erat ager regionis illius plenus hordeo, fugeratque populus a facie Philisthinorum.
1CHR|11|14|Hic stetit in medio agri et defendit eum; cumque percussisset Philisthaeos, dedit Dominus salutem magnam populo suo.
1CHR|11|15|Descenderunt autem tres de triginta principibus ad petram, in qua erat David, ad speluncam Odollam, quando Philisthim fuerant castrametati in valle Raphaim.
1CHR|11|16|Porro David erat in praesidio, et statio Philisthinorum in Bethlehem;
1CHR|11|17|desideravit igitur David et dixit: " O si quis daret mihi aquam de cisterna Bethlehem, quae est in porta! ".
1CHR|11|18|Tres ergo isti per media castra Philisthinorum perrexerunt et hauserunt aquam de cisterna Bethlehem, quae erat in porta, et attulerunt ad David, ut biberet. Qui noluit, sed magis libavit illam Domino
1CHR|11|19|dicens: " Avertat a me Deus meus, ut hoc faciam et sanguinem virorum istorum bibam, quia in periculo animarum suarum attulerunt mihi aquam ". Et ob hanc causam noluit bibere. Haec fecerunt tres robustissimi.
1CHR|11|20|Abisai quoque frater Ioab; ipse erat princeps inter triginta et ipse levavit hastam suam contra trecentos, quos interfecit, et ipse erat inter tres nominatus,
1CHR|11|21|inter triginta duplici honore eminens et princeps eorum; verumtamen usque ad tres non pervenerat.
1CHR|11|22|Banaias filius Ioiadae vir robustissimus, qui multa opera perpetrarat, de Cabseel; ipse percussit duos Ariel de Moab et ipse descendit et interfecit leonem in media cisterna tempore nivis.
1CHR|11|23|Et ipse percussit virum Aegyptium, cuius statura erat quinque cubitorum, et habebat lanceam ut liciatorium texentium; descendit ergo ad eum cum virga et rapuit hastam, quam tenebat manu, et interfecit eum hasta sua.
1CHR|11|24|Haec fecit Banaias filius Ioiadae, qui erat inter tres robustos nominatus,
1CHR|11|25|inter triginta primus; verumtamen ad tres usque non pervenerat, posuit autem eum David super satellites suos.
1CHR|11|26|Porro fortissimi in exercitu: Asael frater Ioab et Elchanan filius Dodo de Bethlehem,
1CHR|11|27|Sammoth Harodites, Elica Harodites, Heles Phalonites,
1CHR|11|28|Hira filius Acces Thecuites, Abiezer Anathothites,
1CHR|11|29|Sobbochai Husathites, Ilai Ahohites,
1CHR|11|30|Maharai Netophathites, Heled filius Baana Netophathites,
1CHR|11|31|Ithai filius Ribai de Gabaa filiorum Beniamin, Banaia Pharathonites,
1CHR|11|32|Hurai de tor rentibus Gaas, Abiel Arbathites,
1CHR|11|33|Azmaveth Bahurimites, Eliaba Saalbonites,
1CHR|11|34|Asem Gezonites, Ionathan filius Sage Ararites,
1CHR|11|35|Ahiam filius Sachar Ararites, Eliphal filius Ur,
1CHR|11|36|Hepher Mecherathites, Ahia Phelonites,
1CHR|11|37|Hesro de Carmel, Naarai filius Azbai,
1CHR|11|38|Ioel frater Nathan, Mibahar filius Agarai,
1CHR|11|39|Selec Ammonites, Naharai Berothites armiger Ioab filii Sarviae,
1CHR|11|40|Hira Iethraeus, Gareb Iethraeus,
1CHR|11|41|Urias Hetthaeus, Zabad filius Oholai,
1CHR|11|42|Adina filius Siza Rubenites princeps Rubenitarum, et cum eo triginta;
1CHR|11|43|Hanan filius Maacha et Iosaphat Matthanites,
1CHR|11|44|Ozia Astharothites, Sama et Iehiel filii Hotham Aroerites,
1CHR|11|45|Iedihel filius Semri et Ioha frater eius Thosaites,
1CHR|11|46|Eliel Mahumites et Ieribai et Iosaia filii Elnaem et Iethma Moabites,
1CHR|11|47|Eliel et Obed et Iasiel de Soba.
1CHR|12|1|Hi quoque venerunt ad Da vid in Siceleg, cum adhuc fu geret Saul filium Cis; qui erant fortissimi et egregii pugnatores
1CHR|12|2|tendentes arcum et utraque manu fundis saxa iacientes et dirigentes sagittas. De fratribus Saul ex Beniamin:
1CHR|12|3|princeps Ahiezer et Ioas filii Samaa Gabaathites et Iaziel et Phalet filii Azmaveth et Baracha et Iehu Anathothites;
1CHR|12|4|Iesmaias quoque Gabaonites fortissimus inter triginta et super triginta,
1CHR|12|5|Ieremias et Iahaziel et Iohanan et Iozabad Gederothites,
1CHR|12|6|Eluzai et Ierimoth et Baalia et Samaria et Saphatia Haruphites,
1CHR|12|7|Elcana et Iesia et Azareel et Ioezer et Iesbaam Coritae,
1CHR|12|8|Ioela quoque et Zabadia filii Ieroham de Gedor.
1CHR|12|9|Sed et de Gad transfugerunt ad David, cum lateret in deserto, viri robustissimi et pugnatores optimi tenentes clipeum et hastam; facies eorum quasi facies leonis et veloces quasi capreae in montibus:
1CHR|12|10|Ezer princeps, Abdias secundus, Eliab tertius,
1CHR|12|11|Masmana quartus, Ieremias quintus,
1CHR|12|12|Etthei sextus, Eliel septimus,
1CHR|12|13|Iohanan octavus, Elzebad nonus,
1CHR|12|14|Ieremias decimus, Machbanai undecimus.
1CHR|12|15|Hi de filiis Gad principes exercitus, minimus contra centum praevalebat et maximus contra mille.
1CHR|12|16|Isti sunt qui transierunt Iordanem mense primo, quando inundare consuevit super ripas suas, et omnes fugaverunt, qui morabantur in vallibus ad orientalem plagam et occidentalem.
1CHR|12|17|Venerunt autem et de Beniamin et de Iuda ad praesidium, in quo morabatur David.
1CHR|12|18|Egressusque est David obviam eis et ait: " Si pacifice venistis ad me, ut auxiliemini mihi, cor meum iungatur vobis; si autem insidiamini mihi pro adversariis meis, cum ego iniquitatem in manibus non habeam, videat Deus patrum nostrorum et iudicet ".
1CHR|12|19|Spiritus vero induit Amasai principem inter triginta, et ait: Tui sumus, o David,et tecum, fili Isai!Pax, pax tibiet pax adiutoribus tuis;te enim adiuvat Deus tuus ".Suscepit ergo eos David et constituit principes turmae.
1CHR|12|20|Porro de Manasse transfugerunt ad David, quando veniebat cum Philisthim adversus Saul, ut pugnaret; et non dimicavit cum eis, quia inito consilio remiserunt eum principes Philisthinorum dicentes: " Periculo capitis nostri revertetur ad dominum suum Saul ".
1CHR|12|21|Quando igitur reversus est in Siceleg, transfugerunt ad eum de Manasse Ednas et Iozabad et Iedihel et Michael et Iozabad et Eliu et Selathai principes milium in Manasse:
1CHR|12|22|hi praebuerunt auxilium David adversus latrunculos; omnes enim erant viri fortissimi et facti sunt principes in exercitu.
1CHR|12|23|Sed et per singulos dies veniebant ad David ad auxiliandum ei, usque dum fieret grandis numerus quasi exercitus Dei.
1CHR|12|24|Iste quoque est numerus principum exercitus, qui venerunt ad David, cum esset in Hebron, ut transferrent regnum Saul ad eum iuxta verbum Domini.
1CHR|12|25|Filii Iudae portantes clipeum et hastam sex milia octingenti expediti ad proelium.
1CHR|12|26|De filiis Simeon virorum fortissimorum ad pugnandum septem milia centum.
1CHR|12|27|De filiis Levi quattuor milia sescenti;
1CHR|12|28|Ioiada quoque princeps de stirpe Aaron et cum eo tria milia septingenti;
1CHR|12|29|Sadoc etiam iuvenis fortissimus et familia eius principes viginti duo.
1CHR|12|30|De filiis autem Beniamin fratribus Saul tria milia; magna enim pars eorum adhuc sequebatur domum Saul.
1CHR|12|31|Porro de filiis Ephraim viginti milia octingenti, fortissimi robore viri nominati in familiis suis.
1CHR|12|32|Et ex dimidia parte tribus Manasse decem et octo milia; singuli per nomina sua destinati, ut venirent et constituerent regem David.
1CHR|12|33|De filiis quoque Issachar viri eruditi, qui norant singula tempora ad sciendum quid facere deberet Israel, principes ducenti et omnes fratres eorum ad iussa eorum.
1CHR|12|34|Porro de Zabulon, qui egrediebantur ad proelium et stabant in acie instructi omnibus armis bellicis, quinquaginta milia venerunt, ut congregarentur non in corde duplici.
1CHR|12|35|Et de Nephthali principes mille; et cum eis instructa clipeo et hasta triginta septem milia.
1CHR|12|36|De Dan etiam praeparata ad proelium viginti octo milia sescenti.
1CHR|12|37|Et de Aser egredientes ad pugnam et in acie procedentes quadraginta milia.
1CHR|12|38|Trans Iordanem autem de filiis Ruben et de Gad et dimidia parte tribus Manasse, instructi omnibus armis bellicis, centum viginti milia.
1CHR|12|39|Omnes isti viri bellatores expediti ad pugnandum corde perfecto venerunt in Hebron, ut constituerent regem David super universum Israel; sed et omnes reliqui ex Israel uno corde erant, ut rex fieret David.
1CHR|12|40|Fueruntque ibi apud David tribus diebus comedentes et bibentes; praeparaverunt enim eis fratres sui.
1CHR|12|41|Sed et qui iuxta eos erant, usque ad Issachar et Zabulon et Nephthali, afferebant panes in asinis et camelis et mulis et bobus, escam farinae, palathas, uvam passam, vinum, oleum, boves, oves ad omnem copiam; gaudium quippe erat in Israel.
1CHR|13|1|Iniit autem consilium David cum tribunis et centurionibus et universis principibus
1CHR|13|2|et ait ad omnem coetum Israel: " Si placet vobis, et a Domino Deo nostro egreditur sermo, quem loquor, mittamus ad fratres nostros reliquos in universas regiones Israel et ad sacerdotes et Levitas, qui habitant in suburbanis urbium, ut congregentur ad nos,
1CHR|13|3|et reducamus arcam Dei nostri ad nos; non enim requisivimus eam in diebus Saul ".
1CHR|13|4|Et respondit universa multitudo, ut ita fieret; placuerat enim sermo omni populo.
1CHR|13|5|Congregavit ergo David cunctum Israel a Sihor Aegypti usque ad introitum dum ingrediaris Emath, ut adduceret arcam Dei de Cariathiarim.
1CHR|13|6|Et ascendit David et omnis Israel in Baala, in Cariathiarim, quae est in Iuda, ut afferrent inde arcam Dei Domini sedentis super cherubim, ubi invocatum est nomen eius.
1CHR|13|7|Imposueruntque arcam Dei super plaustrum novum de domo Abinadab. Oza autem et Ahio minabant plaustrum.
1CHR|13|8|Porro David et universus Israel ludebant coram Deo omni virtute in canticis et in citharis et psalteriis et tympanis et cymbalis et tubis.
1CHR|13|9|Cum autem pervenissent ad aream Chidon, tetendit Oza manum suam, ut sustentaret arcam; boves quippe lascivientes proruperunt.
1CHR|13|10|Iratus est itaque Dominus contra Ozam et percussit eum, eo quod contigisset arcam; et mortuus est ibi coram Deo.
1CHR|13|11|Contristatusque est David, eo quod dirupisset Dominus Ozam; et vocatus est locus ille Pharesoza (id est Diruptio Ozae) usque in praesentem diem.
1CHR|13|12|Et timuit Deum tunc temporis dicens: " Quomodo possum ad me introducere arcam Dei? ".
1CHR|13|13|Et ob hanc causam non eam adduxit ad se, hoc est in civitatem David, sed avertit in domum Obededom Getthaei.
1CHR|13|14|Mansit ergo arca Dei apud domum Obededom tribus mensibus; et benedixit Dominus domui eius et omnibus quae habebat.
1CHR|14|1|Misit quoque Hiram rex Tyri nuntios ad David et ligna cedrina et artifices parietum lignorumque, ut aedificarent ei domum.
1CHR|14|2|Cognovitque David quod confirmasset eum Dominus in regem super Israel et sublevatum esset regnum suum propter populum eius Israel.
1CHR|14|3|Accepit quoque David alias uxores in Ierusalem genuitque filios et filias;
1CHR|14|4|et haec nomina eorum, qui nati sunt ei in Ierusalem: Samua et Sobab, Nathan et Salomon,
1CHR|14|5|Iebahar et Elisua et Eliphalet,
1CHR|14|6|Noga quoque et Napheg et Iaphia,
1CHR|14|7|Elisama et Beeliada et Eliphalet.
1CHR|14|8|Audientes autem Philisthim quod unctus esset David in regem super universum Israel, ascenderunt omnes, ut quaererent eum; quod cum audisset David, egressus est obviam eis.
1CHR|14|9|Porro Philisthim venientes diffusi sunt in valle Raphaim.
1CHR|14|10|Consuluitque David Deum dicens: " Si ascendam contra Philisthaeos, et si trades eos in manu mea? ". Et dixit ei Dominus: " Ascende, et tradam eos in manu tua ".
1CHR|14|11|Cumque illi ascendissent in Baalpharasim, percussit eos ibi David et dixit: " Dirupit Deus inimicos meos per manum meam sicut dirumpuntur aquae. Et idcirco vocatum est nomen loci illius Baalpharasim (id est Dominus diruptionum).
1CHR|14|12|Dereliqueruntque ibi deos suos, quos David iussit exuri.
1CHR|14|13|Alia etiam vice Philisthim irruerunt et diffusi sunt in valle;
1CHR|14|14|consuluitque rursum David Deum, et dixit ei Deus: " Non ascendas post eos; circumdabis eos et venies contra illos ex adverso arborum celthium;
1CHR|14|15|cumque audieris sonitum gradientis in cacumine arborum celthium, tunc egredieris ad bellum; egressus est enim Deus ante te, ut percutias castra Philisthim ".
1CHR|14|16|Fecit ergo David, sicut praeceperat ei Deus, et percussit castra Philisthinorum de Gabaon usque Gazer.
1CHR|14|17|Divulgatumque est nomen David in universis regionibus, et Dominus dedit pavorem eius super omnes gentes.
1CHR|15|1|Fecit quoque sibi domos in civitate David et praeparavit locum arcae Dei tetenditque ei tabernaculum.
1CHR|15|2|Tunc dixit David: " Illicitum est, ut a quocumque portetur arca Dei, nisi a Levitis, quos elegit Dominus ad portandum eam et ad ministrandum sibi usque in aeternum ".
1CHR|15|3|Congregavitque David universum Israel in Ierusalem, ut afferretur arca Domini in locum suum, quem praeparaverat ei;
1CHR|15|4|necnon et filios Aaron et Levitas.
1CHR|15|5|De filiis Caath Uriel princeps fuit et fratres eius centum viginti;
1CHR|15|6|de filiis Merari Asaia princeps et fratres eius ducenti viginti;
1CHR|15|7|de filiis Gerson Ioel princeps et fratres eius centum triginta;
1CHR|15|8|de filiis Elisaphan Semeias princeps et fratres eius ducenti;
1CHR|15|9|de filiis Hebron Eliel princeps et fratres eius octoginta;
1CHR|15|10|de filiis Oziel Aminadab princeps et fratres eius centum duodecim.
1CHR|15|11|Vocavitque David Sadoc et Abiathar sacerdotes et Levitas Uriel, Asaiam, Ioel, Semeiam, Eliel et Aminadab
1CHR|15|12|et dixit ad eos: " Vos, qui estis principes familiarum Leviticarum, sanctificamini cum fratribus vestris et afferte arcam Domini, Dei Israel, ad locum, quem praeparavi.
1CHR|15|13|Quia a principio non eratis praesentes, fecit Dominus, Deus Israel, diruptionem in nobis; non enim quaesivimus eum, sicut fas erat ".
1CHR|15|14|Sanctificati sunt ergo sacerdotes et Levitae, ut portarent arcam Domini, Dei Israel;
1CHR|15|15|et tulerunt filii Levi arcam Dei, sicut praeceperat Moyses iuxta verbum Domini, umeris suis in vectibus.
1CHR|15|16|Dixitque David principibus Levitarum, ut constituerent de fratribus suis cantores in organis musicorum, nablis videlicet et lyris et cymbalis, ut resonaret fortiter sonitus laetitiae.
1CHR|15|17|Constitueruntque Levitae Heman filium Ioel et de fratribus eius Asaph filium Barachiae, de filiis vero Merari fratribus eorum Ethan filium Casaiae
1CHR|15|18|et cum eis fratres eorum in secundo ordine Zachariam et Bani et Iaziel et Semiramoth et Iahiel et Ani, Eliab et Banaiam et Maasiam et Matthathiam et Eliphalu et Maceniam et Obededom et Iehiel ianitores.
1CHR|15|19|Porro cantores Heman, Asaph et Ethan in cymbalis aeneis bene sonantibus,
1CHR|15|20|Zacharias autem et Oziel et Semiramoth et Iahiel et Ani et Eliab et Maasias et Banaias in nablis secundum " Virgines ".
1CHR|15|21|Porro Matthathias et Eliphalu et Macenias et Obededom et Iehiel et Ozaziu in citharis super octavam, ut dirigerent;
1CHR|15|22|Chonenias autem princeps Levitarum portantium arcam praeerat ad portandum, erat quippe valde sapiens.
1CHR|15|23|Et Barachias et Elcana ianitores pro arca.
1CHR|15|24|Porro Sebania et Iosaphat et Nathanael et Amasai et Zacharias et Banaias et Eliezer sacerdotes clangebant tubis coram arca Dei, et Obededom et Iehias erant ianitores pro arca.
1CHR|15|25|Igitur David et maiores natu Israel et tribuni ierunt ad deportandam arcam foederis Domini de domo Obededom cum laetitia.
1CHR|15|26|Cumque adiuvisset Deus Levitas, qui portabant arcam foederis Domini, immolati sunt septem tauri et septem arietes.
1CHR|15|27|Porro David indutus pallio byssino et universi Levitae, qui portabant arcam, cantoresque et Chonenias princeps pro portanda arca - David autem indutus erat etiam ephod lineo -
1CHR|15|28|universusque Israel deducebant arcam foederis Domini in iubilo et sonitu bucinae et tubis et cymbalis bene sonantibus et nablis et citharis.
1CHR|15|29|Cumque pervenisset arca foederis Domini usque ad civitatem David, Michol filia Saul prospiciens per fenestram vidit regem David saltantem atque ludentem et despexit eum in corde suo.
1CHR|16|1|Attulerunt igitur arcam Dei et constituerunt eam in me dio tabernaculi, quod tetenderat ei David, et obtulerunt holocausta et pacifica coram Deo.
1CHR|16|2|Cumque complesset David offerens holocausta et pacifica, benedixit populo in nomine Domini.
1CHR|16|3|Et divisit unicuique de Israel a viro usque ad mulierem tortam panis et laganum palmarum et palatham.
1CHR|16|4|Constituitque coram arca Domini de Levitis ministros, qui recordarentur operum eius et glorificarent atque laudarent Dominum, Deum Israel:
1CHR|16|5|Asaph principem et secundum eius Zachariam, porro Iehiel et Semiramoth et Iahiel et Matthathiam et Eliab et Banaiam et Obededom et Iehiel in organis psalterii et citharis, Asaph autem, ut cymbalis personaret,
1CHR|16|6|Banaiam vero et Iahaziel sacerdotes, ut canerent tubis iugiter coram arca foederis Dei.
1CHR|16|7|In illo die, tunc fecit David prima vice confiteri Domino per manum Asaph et fratrum eius:
1CHR|16|8|" Confitemini Domino, invocate nomen eius,notas facite in populis opera eius.
1CHR|16|9|Canite ei et psalliteet narrate omnia mirabilia eius.
1CHR|16|10|Laudate nomen sanctum eius,laetetur cor quaerentium Dominum.
1CHR|16|11|Quaerite Dominum et virtutem eius,quaerite faciem eius semper.
1CHR|16|12|Recordamini mirabilium eius, quae fecit,signorum illius et iudiciorum oris eius,
1CHR|16|13|semen Israel, servi eius,filii Iacob, electi illius.
1CHR|16|14|Ipse Dominus Deus noster;in universa terra iudicia eius.
1CHR|16|15|Recordamini in sempiternum pacti eius,sermonis, quem praecepit in mille generationes,
1CHR|16|16|pacti, quod pepigit cum Abraham,et iuramenti illius cum Isaac.
1CHR|16|17|Et constituit illud Iacob in praeceptumet Israel in pactum sempiternum
1CHR|16|18|dicens: "Tibi dabo terram Chanaanfuniculum hereditatis vestrae",
1CHR|16|19|cum essent pauci numero,parvi et coloni in ea.
1CHR|16|20|Et transierunt de gente in gentemet de regno ad populum alterum;
1CHR|16|21|non dimisit quemquam calumniari eos,sed increpuit pro eis reges:
1CHR|16|22|"Nolite tangere christos meoset in prophetis meis nolite malignari".
1CHR|16|23|Canite Domino, omnis terra,annuntiate ex die in diem salutare eius.
1CHR|16|24|Narrate in gentibus gloriam eius,in cunctis populis mirabilia illius.
1CHR|16|25|Quia magnus Dominus et laudabilis nimiset horribilis super omnes deos;
1CHR|16|26|omnes enim dii populorum inania,Dominus autem caelos fecit.
1CHR|16|27|Magnificentia et pulchritudo coram eo,fortitudo et gaudium in loco eius.
1CHR|16|28|Afferte Domino, familiae populorumafferte Domino gloriam et imperium;
1CHR|16|29|date Domino gloriam nominis eius,levate oblationem et venite in conspectu eiuset adorate Dominum in decore sancto.
1CHR|16|30|Commoveatur a facie illius omnis terra;ipse enim fundavit orbem immobilem.
1CHR|16|31|Laetentur caeli, et exsultet terra,et dicant in nationibus: "Dominus regnat!".
1CHR|16|32|Tonet mare et plenitudo eius,exsultent agri et omnia, quae in eis sunt.
1CHR|16|33|Tunc laudabunt ligna saltus coram Domino,quia venit iudicare terram.
1CHR|16|34|Confitemini Domino, quoniam bonus,quoniam in aeternum misericordia eius.
1CHR|16|35|Et dicite: "Salva nos, Deus salvator noster,et congrega nos et erue de gentibus, ut confiteamur nomini sancto tuoet exsultemus in carminibus tuis.
1CHR|16|36|Benedictus Dominus, Deus Israel,ab aeterno usque in aeternum" ".Et dixit omnis populus: " Amen! " et " Laus Domino! ".
1CHR|16|37|Dereliquit itaque ibi coram arca foederis Domini Asaph et fratres eius, ut ministrarent in conspectu arcae iugiter secundum ritum singulorum dierum.
1CHR|16|38|Porro Obededom et fratres eius sexaginta octo et Obededom filium Idithun et Hosa constituit ianitores.
1CHR|16|39|Sadoc autem sacerdotem et fratres illius sacerdotes coram habitaculo Domini in excelso, quod erat in Gabaon,
1CHR|16|40|ut offerrent holocausta Domino super altare holocautomatis iugiter, mane et vespere, iuxta omnia, quae scripta sunt in lege Domini, quam praecepit Israeli.
1CHR|16|41|Et cum eis Heman et Idithun et reliquos electos, qui nominatim memorati sunt ad confitendum Domino: " Quoniam in aeternum misericordia eius ".
1CHR|16|42|Et cum eis Heman et Idithun canentes tuba et quatientes cymbala bene sonantia et omnia musicorum organa ad canendum Deo; filios autem Idithun fecit esse portarios.
1CHR|16|43|Reversusque est omnis populus unusquisque in domum suam et David, ut benediceret etiam domui suae.
1CHR|17|1|Cum autem habitaret David in domo sua, dixit ad Nathan prophetam: " Ecce ego habito in domo cedrina, arca autem foederis Domini sub pellibus est ".
1CHR|17|2|Et ait Nathan ad David: " Omnia, quae in corde tuo sunt, fac; Deus enim tecum est ".
1CHR|17|3|Igitur nocte illa factus est sermo Dei ad Nathan dicens:
1CHR|17|4|" Vade et loquere David servo meo: Haec dicit Dominus: Non aedificabis tu mihi domum ad habitandum;
1CHR|17|5|neque enim mansi in domo ex eo tempore, quo eduxi Israel usque ad hanc diem, sed fui semper migrans de tabernaculo in tabernaculum et de habitatione in habitationem.
1CHR|17|6|Ubicumque ambulabam in omni Israel, numquid locutus sum uni iudicum Israel, quibus praeceperam, ut pascerent populum meum, et dixi: Quare non aedificastis mihi domum cedrinam?
1CHR|17|7|Nunc itaque, sic loqueris ad servum meum David: Haec dicit Dominus exercituum: Ego tuli te, cum in pascuis sequereris gregem, ut esses dux populi mei Israel;
1CHR|17|8|et fui tecum, quocumque perrexisti, et interfeci omnes inimicos tuos coram te fecique tibi nomen quasi unius magnorum, qui celebrantur in terra.
1CHR|17|9|Et dedi locum populo meo Israel et plantavi eum, ut habitaret in eo, et ultra non commovebitur, nec filii iniquitatis atterent eos sicut in principio
1CHR|17|10|et ex diebus, quibus dedi iudices populo meo Israel et humiliavi universos inimicos tuos. Annuntio ergo tibi quod aedificaturus sit domum tibi Dominus.
1CHR|17|11|Cumque impleveris dies tuos, ut vadas ad patres tuos, suscitabo semen tuum post te, quod erit de filiis tuis, et stabiliam regnum eius.
1CHR|17|12|Ipse aedificabit mihi domum, et firmabo solium eius usque in aeternum.
1CHR|17|13|Ego ero ei in patrem, et ipse erit mihi in filium; et misericordiam meam non auferam ab eo, sicut abstuli ab eo, qui ante te fuit.
1CHR|17|14|Et statuam eum in domo mea et in regno meo usque in sempiternum, et thronus eius erit firmissimus in perpetuum ".
1CHR|17|15|Iuxta omnia verba haec et iuxta universam visionem istam, sic locutus est Nathan ad David.
1CHR|17|16|Cumque venisset rex David et sedisset coram Domino, dixit: " Quis ego sum, Domine Deus, et quae domus mea, quia adduxisti me hucusque?
1CHR|17|17|Sed hoc parum visum est in conspectu tuo, Deus; ideoque locutus es super domum servi tui etiam in futurum et aspexisti me excelsum super ordinem hominum, Domine Deus.
1CHR|17|18|Quid ultra addere potest David, cum ita glorificaveris servum tuum et cognoveris eum?
1CHR|17|19|Domine, propter famulum tuum iuxta cor tuum fecisti omnem magnificentiam hanc; et nota esse voluisti universa magnalia.
1CHR|17|20|Domine, non est similis tui, et non est alius deus absque te secundum omnia, quae audivimus auribus nostris.
1CHR|17|21|Quis autem est alius ut populus tuus Israel, gens una in terra, ad quam perrexit Deus, ut liberaret sibi populum, ut faceres tibi nomen magnum et terribile eiciens nationes a facie populi tui, quem de Aegypto liberasti?
1CHR|17|22|Et posuisti populum tuum Israel tibi in populum usque in aeternum; et tu, Domine, factus es Deus eius.
1CHR|17|23|Nunc igitur, Domine, sermo, quem locutus es super famulum tuum et super domum eius, confirmetur in perpetuum; et fac, sicut locutus es.
1CHR|17|24|Permaneatque et magnificetur nomen tuum usque in sempiternum, et dicatur: "Dominus exercituum, Deus Israel, est Deus pro Israel, et domus David servi tui permanens coram te".
1CHR|17|25|Tu enim, Deus meus, revelasti auriculam servi tui, ut aedificares ei domum; et idcirco invenit servus tuus fiduciam, ut oret coram te.
1CHR|17|26|Nunc ergo, Domine, tu es Deus; et locutus es super servum tuum tanta beneficia
1CHR|17|27|et coepisti benedicere domui servi tui, ut sit semper coram te: te enim, Domine, benedicente, benedicta erit in perpetuum ".
1CHR|18|1|Factum est autem post haec, ut percuteret David Phili sthim et humiliaret eos et tolleret Geth et filias eius de manu Philisthim
1CHR|18|2|percuteretque Moab, et fierent Moabitae servi David offerentes ei tributum.
1CHR|18|3|Et percussit David etiam Adadezer regem Soba in regione ad Emath, quando perrexit, ut dilataret imperium suum usque ad flumen Euphraten.
1CHR|18|4|Cepit ergo David mille quadrigas eius et septem milia equites ac viginti milia virorum peditum; subnervavitque omnes equos curruum, exceptis centum quadrigis, quas reservavit sibi.
1CHR|18|5|Supervenit autem et Syrus Damascenus, ut auxilium praeberet Adadezer regi Soba; sed et huius percussit David viginti duo milia virorum
1CHR|18|6|et posuit praesidium in Syria Damasci, ut Syria quoque serviret sibi et offerret tributum. Adiuvitque eum Dominus in cunctis, ad quae perrexerat.
1CHR|18|7|Tulit quoque David arma aurea, quae habuerant servi Adadezer, et attulit ea in Ierusalem;
1CHR|18|8|necnon de Tebah et Chun urbibus Adadezer aeris plurimum, de quo fecit Salomon mare aeneum et columnas et vasa aenea.
1CHR|18|9|Quod cum audisset Thou rex Emath, percussisse videlicet David omnem exercitum Adadezer regis Soba,
1CHR|18|10|misit Adoram filium suum ad regem David, ut salutaret eum et congratularetur, eo quod pugnasset cum Adadezer et percussisset eum; adversarius quippe erat Thou Adadezer.
1CHR|18|11|Sed et omnia vasa aurea et argentea et aenea consecravit rex David Domino cum argento et auro, quod tulerat ex universis gentibus, tam de Idumaea et Moab et filiis Ammon, quam de Philisthim et Amalec.
1CHR|18|12|Abisai vero filius Sarviae percussit Edom in valle Salis decem et octo milia
1CHR|18|13|et constituit in Edom praesidium, ut serviret Idumaea David. Salvavitque Dominus David in cunctis, ad quae perrexerat.
1CHR|18|14|Regnavit ergo David super universum Israel et faciebat iudicium atque iustitiam cuncto populo suo.
1CHR|18|15|Porro Ioab filius Sarviae erat super exercitum, et Iosaphat filius Ahilud a commentariis.
1CHR|18|16|Sadoc autem filius Achitob et Achimelech filius Abiathar sacerdotes et Susa scriba.
1CHR|18|17|Banaias vero filius Ioiadae super legiones Cherethi et Phelethi; porro filii David primi ad manum regis.
1CHR|19|1|Accidit autem post haec, ut moreretur Naas rex filiorum Ammon, et regnaret filius eius pro eo.
1CHR|19|2|Dixitque David: " Faciam misericordiam cum Hanon filio Naas; praestitit enim pater eius mihi gratiam ". Misitque David nuntios ad consolandum eum super morte patris sui. Qui cum pervenissent in terram filiorum Ammon, ut consolarentur Hanon,
1CHR|19|3|dixerunt principes filiorum Ammon ad Hanon: " Tu forsitan putas quod David honoris causa in patrem tuum miserit, qui consolentur te; nec animadvertis quod, ut explorent et investigent et evertant terram tuam, venerint ad te servi eius ".
1CHR|19|4|Igitur Hanon pueros David tulit et rasit et praecidit tunicas eorum a natibus usque ad pedes et dimisit eos.
1CHR|19|5|Qui cum abissent et hoc mandassent David, misit in occursum eorum - grandem enim contumeliam sustinuerant - et praecepit, ut manerent in Iericho, donec cresceret barba eorum, et tunc reverterentur.
1CHR|19|6|Videntes autem filii Ammon quod odiosos se fecissent David, tam Hanon quam reliquus populus miserunt mille talenta argenti, ut conducerent sibi de Mesopotamia et de Syria Maacha et de Soba currus et equites;
1CHR|19|7|conduxeruntque sibi triginta duo milia curruum et regem Maacha cum populo eius. Qui cum venissent, castrametati sunt e regione Medaba; filii quoque Ammon congregati de urbibus suis venerunt ad bellum.
1CHR|19|8|Quod cum audisset David, misit Ioab et omnem exercitum virorum fortium.
1CHR|19|9|Egressique filii Ammon direxerunt aciem iuxta portam civitatis; reges autem, qui ad auxilium venerant, separatim in agro steterunt.
1CHR|19|10|Igitur Ioab intellegens bellum et ex adverso et post tergum contra se fieri elegit viros fortissimos de universo Israel et perrexit contra Syrum;
1CHR|19|11|reliquam autem partem populi dedit sub manu Abisai fratris sui, et perrexerunt contra filios Ammon.
1CHR|19|12|Dixitque: " Si vicerit me Syrus, auxilio eris mihi; si autem superaverint te filii Ammon, ero tibi in praesidium.
1CHR|19|13|Confortare et agamus viriliter pro populo nostro et pro urbibus Dei nostri; Dominus autem, quod in conspectu suo bonum est, faciet ".
1CHR|19|14|Appropinquavit ergo Ioab et populus, qui cum eo erat, contra Syrum ad proelium, et fugerunt a facie eorum.
1CHR|19|15|Porro filii Ammon videntes quod fugisset Syrus, ipsi quoque fugerunt Abisai fratrem eius et ingressi sunt civitatem. Reversusque est etiam Ioab in Ierusalem.
1CHR|19|16|Videns autem Syrus quod cecidisset coram Israel, misit nuntios et adduxit Syrum, qui erat trans fluvium; Sophach autem princeps militiae Adadezer erat dux eorum.
1CHR|19|17|Quod cum nuntiatum esset David, congregavit universum Israel et transivit Iordanem venitque ad eos et direxit ex adverso aciem et pugnavit cum eis.
1CHR|19|18|Fugit autem Syrus Israel, et interfecit David de Syris septem milia curruum et quadraginta milia peditum et Sophach exercitus principem.
1CHR|19|19|Videntes autem servi Adadezer se ab Israel esse superatos, fecerunt pacem cum David et servierunt ei; noluitque ultra Syria auxilium praebere filiis Ammon.
1CHR|20|1|Factum est autem post anni circulum, eo tempore, quo solent reges ad bella procedere, eduxit Ioab robur exercitus et vastavit terram filiorum Ammon; perrexitque et obsedit Rabba. Porro David manebat in Ierusalem, quando Ioab percussit Rabba et destruxit eam.
1CHR|20|2|Tulit autem David coronam Melchom de capite eius et invenit in ea auri pondo talentum et pretiosissimam gemmam, venitque super caput David; manubias quoque urbis plurimas tulit.
1CHR|20|3|Populum autem, qui erat in ea, eduxit et condemnavit ad operam lapicidinarum et ad secures et dolabras ferreas. Sic fecit David cunctis urbibus filiorum Ammon et reversus est cum omni populo suo in Ierusalem.
1CHR|20|4|Post haec initum est bellum in Gazer adversum Philisthaeos, in quo percussit Sobbochai Husathites Saphai de genere Raphaim, et humiliavit eos.
1CHR|20|5|Aliud quoque bellum gestum est adversus Philisthaeos, in quo percussit Elchanan filius Iair Lahmi fratrem Goliath Getthaeum, cuius hastae lignum erat quasi liciatorium texentium.
1CHR|20|6|Sed et aliud bellum accidit in Geth, in quo fuit homo longissimus senos habens digitos, id est simul viginti quattuor, qui et ipse de Rapha fuerat stirpe generatus;
1CHR|20|7|hic blasphemavit Israel, et percussit eum Ionathan filius Samma fratris David. Hi sunt filii Rapha in Geth, qui ceciderunt in manu David et servorum eius.
1CHR|21|1|Consurrexit autem Satan contra Israel et incitavit Da vid, ut numeraret Israel.
1CHR|21|2|Dixitque David ad Ioab et ad principes populi: " Ite et numerate Israel a Bersabee usque Dan et afferte mihi numerum, ut sciam ".
1CHR|21|3|Responditque Ioab: " Augeat Dominus populum suum centuplum quam sunt. Nonne, domine mi rex, omnes servi tui sunt? Quare hoc quaerit dominus meus, quod in peccatum reputetur Israeli? ".
1CHR|21|4|Sed sermo regis magis praevaluit; egressusque est Ioab et circuivit universum Israel et reversus est Ierusalem.
1CHR|21|5|Deditque David numerum census, et inventus est omnis Israel numerus mille milia et centum milia virorum educentium gladium; de Iuda autem quadringenta septuaginta milia bellatorum;
1CHR|21|6|nam Levi et Beniamin non numeravit in medio eorum, eo quod invitus exequeretur regis imperium.
1CHR|21|7|Displicuit autem Deo, quod iussum erat, et percussit Israel.
1CHR|21|8|Dixitque David ad Deum: " Peccavi nimis, ut hoc facerem; obsecro, aufer iniquitatem servi tui, quia valde insipienter egi ".
1CHR|21|9|Et locutus est Dominus ad Gad videntem David dicens:
1CHR|21|10|" Vade et loquere ad David et dic: Haec dicit Dominus: Trium tibi optionem do: unum, quod volueris, elige, et faciam tibi ".
1CHR|21|11|Cumque venisset Gad ad David, dixit ei: " Haec dicit Dominus: Elige, quod volueris:
1CHR|21|12|aut tribus annis famem aut tribus mensibus fugere te hostes tuos et gladium eorum non posse evadere aut tribus diebus gladium Domini et pestilentiam versari in terra et angelum Domini interficere in universis finibus Israel. Nunc igitur vide quid respondeam ei, qui misit me ".
1CHR|21|13|Et dixit David ad Gad: " Ex omni parte me angustiae premunt, sed melius mihi est, ut incidam in manus Domini, quia multae sunt miserationes eius, quam in manus hominum ".
1CHR|21|14|Misit ergo Dominus pestilentiam in Israel, et ceciderunt de Israel septuaginta milia virorum.
1CHR|21|15|Misit quoque Deus angelum in Ierusalem, ut percuteret eam. Cumque percuteretur, vidit Dominus et misertus est super magnitudinem mali et imperavit angelo, qui percutiebat: " Sufficit, iam cesset manus tua ".Porro angelus Domini stabat iuxta aream Ornan Iebusaei.
1CHR|21|16|Levansque David oculos suos vidit angelum Domini stantem inter terram et caelum et evaginatum gladium in manu eius et versum contra Ierusalem; et ceciderunt tam ipse quam maiores natu vestiti ciliciis proni in terram.
1CHR|21|17|Dixitque David ad Deum: " Nonne ego sum, qui iussi, ut numeraretur populus? Ego qui peccavi, ego qui malum feci; iste grex quid commeruit? Domine Deus meus, vertatur, obsecro, manus tua in me et in domum patris mei; populus autem tuus non percutiatur ".
1CHR|21|18|Angelus autem Domini praecepit Gad dicere David, ut ascenderet exstrueretque altare Domino in area Ornan Iebusaei.
1CHR|21|19|Ascendit ergo David iuxta sermonem Gad, quem locutus fuerat ex nomine Domini.
1CHR|21|20|Porro Ornan, cum conversus vidisset angelum, quattuorque filii eius cum eo absconderunt se; nam eo tempore terebat in area triticum.
1CHR|21|21|Igitur, cum veniret David ad Ornan, conspexit eum Ornan et processit ei obviam de area et adoravit illum pronus in terram.
1CHR|21|22|Dixitque ei David: " Da mihi locum areae tuae, ut aedificem in ea altare Domino, ita ut quantum valet argenti accipias, et cesset plaga a populo ".
1CHR|21|23|Dixit autem Ornan ad David: " Tolle, et faciat dominus meus rex, quodcumque ei placet; sed et boves do in holocaustum et tribulas in ligna et triticum in sacrificium; omnia libens praebebo ".
1CHR|21|24|Dixitque ei rex David: " Nequaquam ita fiet, sed argentum dabo quantum valet; neque enim tibi auferre debeo et sic offerre Domino holocausta gratuita ".
1CHR|21|25|Dedit ergo David Ornan pro loco siclos auri iustissimi ponderis sescentos
1CHR|21|26|et aedificavit ibi altare Domino obtulitque holocausta et pacifica et invocavit Dominum. Et exaudivit eum in igne de caelo super altare holocausti,
1CHR|21|27|praecepitque Dominus angelo, et convertit gladium suum in vaginam.
1CHR|21|28|In illo ergo tempore David videns quod exaudisset eum Dominus in area Ornan Iebusaei immolavit ibi victimas.
1CHR|21|29|Tabernaculum autem Domini, quod fecerat Moyses in deserto, et altare holocaustorum ea tempestate erat in excelso Gabaon;
1CHR|21|30|et non praevaluit David ire, ut ibi obsecraret Deum; nimio enim fuerat timore perterritus videns gladium angeli Domini.
1CHR|22|1|Dixitque David: " Haec est domus Domini Dei, et hoc est altare holocausti pro Israel ".
1CHR|22|2|Et praecepit, ut congregarentur omnes advenae de terra Israel, et constituit ex eis latomos ad caedendos lapides et poliendos, ut aedificaretur domus Dei.
1CHR|22|3|Ferrum quoque plurimum ad clavos ianuarum et ad commissuras atque iuncturas praeparavit David et aeris pondus innumerabile.
1CHR|22|4|Ligna quoque cedrina non poterant aestimari, quae Sidonii et Tyrii deportaverant ad David.
1CHR|22|5|Et dixit David: " Salomon filius meus puer parvulus est et tener; domus autem, quae aedificanda est Domino, talis esse debet, ut in cunctis regionibus nominetur et glorificetur. Praeparabo ergo ei necessaria ". Et ob hanc causam ante mortem suam omnes paravit impensas.
1CHR|22|6|Vocavitque Salomonem filium suum et praecepit ei, ut aedificaret domum Domino, Deo Israel;
1CHR|22|7|dixitque David ad Salomonem: " Fili mi, voluntatis meae fuit, ut aedificarem domum nomini Domini Dei mei,
1CHR|22|8|sed factus est ad me sermo Domini dicens: "Multum sanguinem effudisti et magna bella bellasti. Non poteris aedificare domum nomini meo, tanto effuso sanguine coram me.
1CHR|22|9|Filius, qui nascetur tibi, erit vir quietissimus; faciam enim eum requiescere ab omnibus inimicis suis per circuitum et ob hanc causam Salomon vocabitur, et pacem et otium dabo in Israel cunctis diebus eius.
1CHR|22|10|Ipse aedificabit domum nomini meo, et ipse erit mihi in filium, et ego ero ei in patrem; firmaboque solium regni eius super Israel in aeternum".
1CHR|22|11|Nunc ergo, fili mi, sit Dominus tecum; et prosperare et aedifica domum Domino Deo tuo, sicut locutus est de te.
1CHR|22|12|Tantum det tibi Dominus prudentiam et sensum, ut regere possis Israel et custodire legem Domini Dei tui;
1CHR|22|13|tunc enim proficere poteris, si custodieris mandata et iudicia, quae praecepit Dominus Moysi super Israel. Confortare et viriliter age; ne timeas neque paveas.
1CHR|22|14|Ecce ego in labore meo praeparavi impensas domus Domini: auri talenta centum milia et argenti mille milia talentorum, aeris vero et ferri non est pondus, vincitur enim numerus magnitudine. Ligna et lapides praeparavi; tu autem ad ea adicies.
1CHR|22|15|Habes quoque plurimos artifices latomos et caementarios artificesque lignorum et omnium artium ad faciendum opus prudentissimos
1CHR|22|16|in auro et argento et aere et ferro, cuius non est numerus. Surge igitur et fac, et erit Dominus tecum ".
1CHR|22|17|Praecepit quoque David cunctis principibus Israel, ut adiuvarent Salomonem filium suum: "
1CHR|22|18|Cernitis, inquiens, quod Dominus Deus vester vobiscum sit et dederit vobis requiem per circuitum et tradiderit habitatores terrae in manu vestra, et subiecta sit terra coram Domino et coram populo eius.
1CHR|22|19|Praebete igitur corda vestra et animas vestras, ut quaeratis Dominum Deum vestrum; et consurgite et aedificate sanctuarium Domini Dei, ut introducatur arca foederis Domini et vasa Deo consecrata in domum, quae aedificatur nomini Domini ".
1CHR|23|1|Igitur David senex et plenus dierum regem constituit Sa lomonem filium suum super Israel
1CHR|23|2|et congregavit omnes principes Israel et sacerdotes atque Levitas.
1CHR|23|3|Numeratique sunt Levitae a triginta annis et supra, et inventa sunt triginta octo milia virorum.
1CHR|23|4|" Ex his, inquit, praesint ministerio domus Domini viginti quattuor milia, praepositi autem et iudices sex milia;
1CHR|23|5|porro quattuor milia ianitores et totidem psaltae canentes Domino in organis, quae feci ad canendum ".
1CHR|23|6|Et distribuit eos David per vices filiorum Levi Gerson videlicet et Caath et Merari.
1CHR|23|7|Filii Gerson: Ladan et Semei.
1CHR|23|8|Filii Ladan: princeps Iahiel et Zetham et Ioel, tres.
1CHR|23|9|Filii Semei: Salomith et Hoziel et Aran, tres; isti principes familiarum Ladan.
1CHR|23|10|Porro filii Semei: Iahath et Ziza et Iehus et Beria; isti filii Semei, quattuor.
1CHR|23|11|Erat autem Iahath prior, Ziza secundus; porro Iehus et Beria non habuerunt plurimos filios, et idcirco in una familia unaque domo computati sunt.
1CHR|23|12|Filii Caath: Amram et Isaar, Hebron et Oziel, quattuor.
1CHR|23|13|Filii Amram: Aaron et Moyses. Separatusque est Aaron, ut sanctificaret sanctissima, ipse et filii eius in sempiternum, et adoleret Domino et serviret ei ac benediceret in nomine eius in perpetuum.
1CHR|23|14|Moysi quoque hominis Dei filii annumerati sunt in tribu Levi.
1CHR|23|15|Filii Moysi: Gersam et Eliezer.
1CHR|23|16|Filii Gersam: Subael primus.
1CHR|23|17|Fuerunt autem filii Eliezer: Rohobia primus, et non erant Eliezer filii alii; porro filii Rohobia multiplicati sunt nimis.
1CHR|23|18|Filii Isaar: Salomoth primus.
1CHR|23|19|Filii Hebron: Ieriau primus, Amarias secundus, Iahaziel tertius, Iecmaam quartus.
1CHR|23|20|Filii Oziel: Micha primus, Iesia secundus.
1CHR|23|21|Filii Merari: Moholi et Musi. Filii Moholi: Eleazar et Cis;
1CHR|23|22|mortuus est autem Eleazar et non habuit filios sed filias acceperuntque eas filii Cis fratres earum.
1CHR|23|23|Filii Musi: Moholi et Eder et Ierimoth, tres.
1CHR|23|24|Hi filii Levi in familiis suis, principes familiarum per vices et numerum capitum singulorum, qui faciebant opera ministerii domus Domini a viginti annis et supra.
1CHR|23|25|Dixit enim David: " Requiem dedit Dominus, Deus Israel, populo suo et habitat in Ierusalem usque in aeternum;
1CHR|23|26|nec erit officii Levitarum, ut ultra portent tabernaculum et omnia vasa eius ad ministrandum.
1CHR|23|27|Iuxta praecepta igitur David novissima, supputabitur numerus filiorum Levi a viginti annis et supra,
1CHR|23|28|et erunt sub manu filiorum Aaron in cultum domus Domini pro atriis et exedris et in purificationem omnis rei sacrae et in ministerium templi Dei,
1CHR|23|29|pro panibus propositionis et farina oblationis et laganis azymorum et pro sartagine et ad torrendum et super omne pondus atque mensuram.
1CHR|23|30|Et stent mane ad confitendum et canendum Domino similiterque ad vesperam,
1CHR|23|31|tam in oblatione holocaustorum Domini quam in sabbatis et calendis et sollemnitatibus reliquis, iuxta numerum et caeremonias uniuscuiusque rei iugiter coram Domino.
1CHR|23|32|Et custodiant observationes tabernaculi conventus et ritum sanctuarii et observationem filiorum Aaron fratrum suorum, ut ministrent in domo Domini ".
1CHR|24|1|Porro filiis Aaron hae partiones erant.Filii Aaron: Nadab et Abiu et Eleazar et Ithamar.
1CHR|24|2|Mortui sunt autem Nadab et Abiu ante patrem suum absque liberis; sacerdotioque functus est Eleazar et Ithamar.
1CHR|24|3|Et divisit eos David cum Sadoc de filiis Eleazari et cum Achimelech de filiis Ithamar, secundum vices suas et ministerium.
1CHR|24|4|Inventique sunt multo plures filii Eleazar secundum capita virorum quam filii Ithamar; divisit igitur eis, hoc est filiis Eleazar principes per familias sedecim, et filiis Ithamar per familias et domos suas octo.
1CHR|24|5|Porro divisit utrasque inter se familias sortibus; erant enim principes sanctuarii et principes Dei tam de filiis Eleazar quam de filiis Ithamar.
1CHR|24|6|Descripsitque eos Semeias filius Nathanael scriba Levites coram rege et principibus et Sadoc sacerdote et Achimelech filio Abiathar, principibus quoque familiarum sacerdotalium et leviticarum: unam familiam pro Eleazar et unam pro Ithamar.
1CHR|24|7|Exivit autem sors prima Ioiarib, secunda Iedaiae,
1CHR|24|8|tertia Harim, quarta Seorim,
1CHR|24|9|quinta Melchia, sexta Miamin,
1CHR|24|10|septima Accos, octava Abia,
1CHR|24|11|nona Iesua, decima Sechenia,
1CHR|24|12|undecima Eliasib, duodecima Iacim,
1CHR|24|13|tertia decima Hoppha, quarta decima Isbaab,
1CHR|24|14|quinta decima Belga, sexta decima Emmer,
1CHR|24|15|septima decima Hezir, octava decima Aphses,
1CHR|24|16|nona decima Phethahia, vicesima Hezechiel,
1CHR|24|17|vicesima prima Iachin, vicesima secunda Gamul,
1CHR|24|18|vicesima tertia Dalaiau, vicesima quarta Maaziau.
1CHR|24|19|Hae vices eorum secundum ministeria sua, ut ingrediantur domum Domini, et iuxta ritum suum sub manu Aaron patris eorum, sicut praecepit Dominus, Deus Israel.
1CHR|24|20|Porro filiorum Levi, qui reliqui fuerant: de filiis Amram Subael et de filiis Subael Iehedeia.
1CHR|24|21|De filiis quoque Rohobiae princeps Iesias.
1CHR|24|22|De Isaaritis vero Salomoth; de filiis Salomoth Iahath.
1CHR|24|23|De Hebronitis: Ieriau, Amarias secundus, Iahaziel tertius, Iecmaam quartus.
1CHR|24|24|Filius Oziel Micha; de filiis Micha Samir;
1CHR|24|25|frater Micha Iesia; de filiis Iesiae Zacharias.
1CHR|24|26|Filii Merari: Moholi et Musi. Filii eius: Iaziau et Bani.
1CHR|24|27|Filius Merari: de Iaziau filio suo Soam et Zacchur et Hebri.
1CHR|24|28|Porro de Moholi filius Eleazar, qui non habebat liberos.
1CHR|24|29|Filius vero Cis Ierameel;
1CHR|24|30|filii Musi: Moholi, Eder et Ierimoth.Isti filii Levi secundum familias suas.
1CHR|24|31|Ipsi quoque miserunt sortes sicut fratres sui, filii Aaron coram David rege et Sadoc et Achimelech et principibus familiarum sacerdotalium et leviticarum tam maiores quam minores; omnes sors aequaliter dividebat.
1CHR|25|1|Igitur David et magistratus exercitus segregaverunt in ministerium filios Asaph et Heman et Idithun, qui prophetarent in citharis et psalteriis et cymbalis, secundum numerum suum dedicato sibi officio servientes.
1CHR|25|2|De filiis Asaph: Zacchur et Ioseph et Nathania et Asarela filii Asaph erant sub manu Asaph prophetantis sub manu regis.
1CHR|25|3|De Idithun; filii Idithun: Godolias, Sori, Iesaias et Hasabias et Matthathias, sex, sub manu patris sui Idithun, qui in cithara prophetabat ad confitendum et laudandum Dominum.
1CHR|25|4|De Heman quoque; filii Heman: Bocciau, Matthaniau, Oziel, Subael et Ierimoth, Hananias, Hanani, Eliatha, Geddelthi et Romemthiezer et Iesbacasa, Mellothi, Othir, Mahazioth;
1CHR|25|5|omnes isti filii Heman videntis regis iuxta sermones Dei, quod exaltaret cornu eius; deditque Deus Heman filios quattuordecim et filias tres.
1CHR|25|6|Universi sub manu patris sui ad cantandum in templo Domini distributi erant in cymbalis et psalteriis et citharis, in ministeria domus Dei sub manu regis: Asaph et Idithun et Heman.
1CHR|25|7|Fuit autem numerus eorum cum fratribus suis eruditis in cantando Domino, cuncti magistri, ducenti octoginta octo.
1CHR|25|8|Miseruntque sortes pro ministerio ex aequo, tam maior quam minor, magister pariter et discipulus.
1CHR|25|9|Egressaque est sors prima Ioseph, qui erat de Asaph. Secunda Godoliae, ipsi et fratribus eius et filiis eius, duodecim.
1CHR|25|10|Tertia Zacchur, filiis et fratribus eius, duodecim.
1CHR|25|11|Quarta Isari, filiis et fratribus eius, duodecim.
1CHR|25|12|Quinta Nathaniau, filiis et fratribus eius, duodecim.
1CHR|25|13|Sexta Bocciau, filiis et fratribus eius, duodecim.
1CHR|25|14|Septima Isreela, filiis et fratribus eius, duodecim.
1CHR|25|15|Octava Iesaiae, filiis et fratribus eius, duodecim.
1CHR|25|16|Nona Matthaniau, filiis et fratribus eius, duodecim.
1CHR|25|17|Decima Semei, filiis et fratribus eius, duodecim.
1CHR|25|18|Undecima Azareel, filiis et fratribus eius, duodecim.
1CHR|25|19|Duodecima Hasabiae, filiis et fratribus eius, duodecim.
1CHR|25|20|Tertia decima Subael, filiis et fratribus eius, duodecim.
1CHR|25|21|Quarta decima Matthathiae, filiis et fratribus eius, duodecim.
1CHR|25|22|Quinta decima Ierimoth, filiis et fratribus eius, duodecim.
1CHR|25|23|Sexta decima Hananiae, filiis et fratribus eius, duodecim.
1CHR|25|24|Septima decima Iesbacasae, filiis et fratribus eius, duodecim.
1CHR|25|25|Octava decima Hanani, filiis et fratribus eius, duodecim.
1CHR|25|26|Nona decima Mellothi, filiis et fratribus eius, duodecim.
1CHR|25|27|Vicesima Eliatha, filiis et fratribus eius, duodecim.
1CHR|25|28|Vicesima prima Othir, filiis et fratribus eius, duodecim.
1CHR|25|29|Vicesima secunda Geddelthi, filiis et fratribus eius, duodecim.
1CHR|25|30|Vicesima tertia Mahazioth, filiis et fratribus eius, duodecim.
1CHR|25|31|Vicesima quarta Romemthiezer, filiis et fratribus eius, duodecim.
1CHR|26|1|Divisiones autem ianitorum.De Coritis: Meselemia filius Core de filiis Abiasaph.
1CHR|26|2|Filii Meselemiae: Zacharias primogenitus, Iedihel secundus, Zabadias tertius, Iathanael quartus,
1CHR|26|3|Elam quintus, Iohanan sextus, Elioenai septimus.
1CHR|26|4|Filii autem Obededom: Semeias primogenitus, Iozabad secundus, Ioah tertius, Sachar quartus, Nathanael quintus,
1CHR|26|5|Ammiel sextus, Issachar septimus, Phollathi octavus, quia benedixit illi Deus.
1CHR|26|6|Semeiae autem filio eius nati sunt filii praefecti familiarum suarum, erant enim viri fortissimi;
1CHR|26|7|filii ergo Semeiae: Othni et Raphael et Obed, Elzabad, fratres eius viri fortissimi, Eliu quoque et Samachias;
1CHR|26|8|omnes hi de filiis Obededom, ipsi et filii et fratres eorum fortissimi ad ministrandum sexaginta duo de Obededom.
1CHR|26|9|Porro Meselemiae filii et fratres eorum robustissimi decem et octo.
1CHR|26|10|De Hosa autem, de filiis Merari, erant filii: Semri princeps - non enim fuerat primogenitus, et idcirco posuerat eum pater eius in principem -
1CHR|26|11|Helcias secundus, Tabelias tertius, Zacharias quartus; omnes hi filii et fratres Hosa tredecim.
1CHR|26|12|Hae divisiones ianitorum: secundum capita virorum habebant ministeria sicut et fratres eorum ad ministrandum in domo Domini.
1CHR|26|13|Missae sunt ergo sortes ex aequo et parvis et magnis per familias suas in unamquamque portarum.
1CHR|26|14|Cecidit igitur sors orientalis Selemiae; porro Zachariae filio eius consiliario prudentissimo et erudito sortito obtigit plaga septentrionalis;
1CHR|26|15|Obededom vero australis, et filiis eius horreum;
1CHR|26|16|Sephim et Hosa occidentalis iuxta portam Sallecheth apud viam ascensionis. Custodia iuxta custodiam:
1CHR|26|17|ad orientem per diem sex et ad aquilonem quattuor per diem, atque ad meridiem similiter in die quattuor et pro horreo bini et bini,
1CHR|26|18|pro Parbar quoque ad occidentem quattuor in via, duo pro Parbar.
1CHR|26|19|Hae sunt divisiones ianitorum filiorum Core et Merari.
1CHR|26|20|Porro Levitae fratres eorum super thesauros domus Dei ac thesauros rerum consecratarum.
1CHR|26|21|De filiis Ladan Gersonitae principes familiarum Ladan Gersonitae erant Iahielitae.
1CHR|26|22|Filii Iahiel et Zetham et Ioel fratrum eius erant super thesauros domus Domini.
1CHR|26|23|De Amramitis et Isaaritis et Hebronitis et Ozielitis:
1CHR|26|24|Subael filius Gersam filii Moysi praepositus thesauris.
1CHR|26|25|Fratres quoque eius Eliezer, cuius filius Rohobia et huius filius Iesaias; et huius filius Ioram, huius quoque filius Zechri et huius filius Selemith.
1CHR|26|26|Ipse Selemith et fratres eius super omnes thesauros rerum consecratarum, quas sanctificavit David rex et principes familiarum et tribuni et centuriones et duces exercitus
1CHR|26|27|de bellis et manubiis proeliorum, quas consecraverant ad sustentandum templum Domini.
1CHR|26|28|Et universa, quae consecraverant Samuel videns et Saul filius Cis et Abner filius Ner et Ioab filius Sarviae, omnia donaria sacra erant sub manu Selemith et fratrum eius.
1CHR|26|29|De Isaaritis vero erant Chonenias et filii eius ad opera forinsecus super Israel praefecti et iudices.
1CHR|26|30|Porro de Hebronitis Hasabias et fratres eius viri strenui mille septingenti erant magistratus Israel trans Iordanem contra occidentem in cunctis operibus Domini et in ministerium regis;
1CHR|26|31|Hebronitarum autem princeps fuit Ieria secundum cognationes et familias eorum. Quadragesimo anno regni David recensiti sunt et inventi viri fortes in Iazer Galaad
1CHR|26|32|fratresque eius viri strenui duo milia septingenti principes familiarum; praeposuit autem eos David rex Rubenitis et Gadditis et dimidio tribus Manasse in omne ministerium Dei et regis.
1CHR|27|1|Filii autem Israel secundum numerum suum, principes fa miliarum, tribuni et centuriones et praefecti, qui ministrabant regi iuxta turmas suas ingredientes et egredientes per singulos menses in anno, unaquaeque turma viginti quattuor milia.
1CHR|27|2|Primae turmae in primo mense Iesbaam praeerat filius Zabdiel, et sub eo viginti quattuor milia;
1CHR|27|3|erat de filiis Phares princeps cunctorum principum in exercitu mense primo.
1CHR|27|4|Secundi mensis habebat turmam Dudi Ahohites, et sub eo viginti quattuor milia.
1CHR|27|5|Dux quoque turmae tertiae in mense tertio erat Banaias filius Ioiadae sacerdotis, et in divisione sua viginti quattuor milia;
1CHR|27|6|ipse est Banaias fortissimus inter triginta et super triginta; praeerat autem turmae ipsius Amizabad filius eius.
1CHR|27|7|Quartus, mense quarto, Asael frater Ioab et Zabadias filius eius post eum, et in turma eius viginti quattuor milia.
1CHR|27|8|Quintus, mense quinto, princeps Samaoth Zaraita, et in turma eius viginti quattuor milia.
1CHR|27|9|Sextus, mense sexto, Hira filius Acces Thecuites, et in turma eius viginti quattuor milia.
1CHR|27|10|Septimus, mense septimo, Helles Phalonites de filiis Ephraim, et in turma eius viginti quattuor milia.
1CHR|27|11|Octavus, mense octavo, Sobbochai Husathites de stirpe Zara, et in turma eius viginti quattuor milia.
1CHR|27|12|Nonus, mense nono, Abiezer Anathothites de filiis Beniamin, et in turma eius viginti quattuor milia.
1CHR|27|13|Decimus, mense decimo, Maharai Netophathites de stirpe Zara, et in turma eius viginti quattuor milia.
1CHR|27|14|Undecimus, mense undecimo, Banaias Pharathonites de filiis Ephraim, et in turma eius viginti quattuor milia.
1CHR|27|15|Duodecimus, mense duodecimo, Holdai Netophathites de stirpe Othoniel, et in turma eius viginti quattuor milia.
1CHR|27|16|Porro tribubus praeerant Israel: Rubenitis dux Eliezer filius Zechri; Simeonitis Saphatia filius Maacha;
1CHR|27|17|Levitis Hasabias filius Camuel; Aaronitis Sadoc;
1CHR|27|18|Iudae Eliu de fratribus David; Issachar Amri filius Michael;
1CHR|27|19|Zabulon Iesmaias filius Abdiae; Nephthali Ierimoth filius Azriel;
1CHR|27|20|filiis Ephraim Osee filius Ozaziu; dimidio tribus Manasse Ioel filius Phadaiae;
1CHR|27|21|et dimidio tribus Manasse in Galaad Iaddo filius Zachariae; Beniamin autem Iasiel filius Abner;
1CHR|27|22|Dan vero Azareel filius Ieroham: hi principes tribuum Israel.
1CHR|27|23|Noluit autem David numerare eos a viginti annis inferius, quia dixerat Dominus ut multiplicaret Israel quasi stellas caeli.
1CHR|27|24|Ioab filius Sarviae coeperat numerare nec complevit, quia super hoc ira irruerat in Israel, et idcirco numerus non est relatus in librum annalium regis David.
1CHR|27|25|Super thesauros autem regis fuit Azmaveth filius Adiel; his autem thesauris, qui erant in regione, in urbibus et in vicis et in turribus praesidebat Ionathan filius Oziae.
1CHR|27|26|Operi autem rustico et agricolis, qui exercebant terram, praeerat Ezri filius Chelub.
1CHR|27|27|Vinearumque cultoribus Semei Ramathites; cellis autem vinariis in vineis Zabdi Sephamatites.
1CHR|27|28|Nam super oliveta et ficeta, quae erant in Sephela, Baalhanan Gederites; super apothecas autem olei Ioas.
1CHR|27|29|Porro armentis, quae pascebantur in Saron, praepositus fuit Setrai Saronites, et super boves in vallibus Saphat filius Adli.
1CHR|27|30|Super camelos vero Ubil Ismaelites, et super asinas Iehedeia Meronathites;
1CHR|27|31|super oves quoque Iaziz Agarenus: omnes hi principes substantiae regis David.
1CHR|27|32|Ionathan autem patruus David consiliarius, vir prudens et litteratus, ipse et Iahiel filius Hachamonitis erant cum filiis regis.
1CHR|27|33|Achitophel etiam consiliarius regis, et Chusai Arachites amicus regis;
1CHR|27|34|post Achitophel fuit Ioiada filius Banaiae et Abiathar. Princeps autem exercitus regis erat Ioab.
1CHR|28|1|Convocavit igitur David om nes principes Israel, duces tri buum et praepositos turmarum, qui ministrabant regi, tribunos quoque et centuriones et, qui praeerant substantiae et gregibus regis filiorumque suorum, cum eunuchis et fortibus et robustissimis quibusque in exercitu Ierusalem.
1CHR|28|2|Cumque surrexisset rex et stetisset, ait: " Audite me, fratres mei et populus meus. Cogitavi ut aedificarem domum, in qua requiesceret arca foederis Domini et scabellum pedum Dei nostri, et ad aedificandum omnia praeparavi;
1CHR|28|3|Deus autem dixit mihi: "Non aedificabis domum nomini meo, eo quod sis vir bellator et sanguinem fuderis".
1CHR|28|4|Sed elegit Dominus, Deus Israel, me de universa domo patris mei, ut essem rex super Israel in sempiternum; Iudam enim elegit principem, porro in domo Iudae domum patris mei, et in filiis patris mei placuit ei, ut me eligeret regem super cunctum Israel.
1CHR|28|5|Sed et de filiis meis - filios enim multos dedit mihi Dominus - elegit Salomonem filium meum, ut sederet in throno regni Domini super Israel.
1CHR|28|6|Dixitque mihi: "Salomon filius tuus aedificabit domum meam et atria mea; ipsum enim elegi mihi in filium, et ego ero ei in patrem.
1CHR|28|7|Et firmabo regnum eius usque in aeternum, si perseveraverit facere praecepta mea et iudicia, sicut et hodie".
1CHR|28|8|Nunc igitur coram universo Israel coetu Domini, audiente Deo nostro, custodite et perquirite cuncta mandata Domini Dei vestri, ut possideatis terram bonam et relinquatis eam in hereditatem filiis vestris post vos usque in sempiternum.
1CHR|28|9|Tu autem, Salomon, fili mi, scito Deum patris tui et servi ei corde perfecto et animo voluntario; omnia enim corda scrutatur Dominus et universas mentium cogitationes intellegit. Si quaesieris eum, invenies; si autem dereliqueris illum, proiciet te in aeternum.
1CHR|28|10|Nunc ergo vide quia elegit te Dominus, ut aedificares domum sanctuarii; confortare et perfice ".
1CHR|28|11|Dedit autem David Salomoni filio suo descriptionem porticus et templi et cellariorum et cenaculorum et cubiculorum interiorum et domus propitiatorii
1CHR|28|12|necnon et omnium, quae per Spiritum cum eo erant, de atriis domus Domini et de omnibus exedris per circuitum, de thesauris domus Dei et de thesauris rerum consecratarum
1CHR|28|13|et de divisionibus sacerdotalibus et leviticis, de omni opere ministerii domus Domini et de universis vasis ministerii templi Domini,
1CHR|28|14|de auro in pondere per singula vasa ministerii, de omnibus vasis argenteis in pondere per omnia vasa pro operum diversitate;
1CHR|28|15|sed et ad candelabra aurea et ad lucernas eorum aurum pro mensura uniuscuiusque candelabri et lucernarum, similiter et in candelabris argenteis et in lucernis eorum pro diversitate mensurae, pondus argenti indicavit.
1CHR|28|16|Aurum quoque in mensas propositionis pro diversitate mensarum, similiter et argentum in alias mensas argenteas;
1CHR|28|17|ad fuscinulas quoque et phialas et crateras ex auro purissimo et scyphos aureos pro qualitate mensurae pondus distribuit in scyphum et scyphum; similiter et in scyphos argenteos diversum argenti pondus constituit,
1CHR|28|18|altari autem, in quo adoletur incensum, aurum purissimum, et aurum pro structura quadrigae cherubim extendentium alas et velantium arcam foederis Domini.
1CHR|28|19|" Omnia, inquit, venerunt scripta manu Domini ad me, ut intellegerem universa opera exemplaris ".
1CHR|28|20|Dixit quoque David Salomoni filio suo: " Viriliter age et confortare et fac, ne timeas et ne paveas; Dominus enim Deus meus tecum erit et non dimittet te nec derelinquet, donec perficias omne opus ministerii domus Domini.
1CHR|28|21|Ecce divisiones sacerdotum et Levitarum: parati erunt in omne ministerium domus Dei; et assistet tibi in omni opere quisquis in sapientia ad omne ministerium promptus fuerit, principes quoque et universus populus in negotiis tuis ".
1CHR|29|1|Locutusque est David rex ad omnem ecclesiam: " Salomo nem filium meum unum elegit Deus adhuc puerum et tenellum; opus autem grande est: neque enim homini praeparatur habitatio sed Domino Deo.
1CHR|29|2|Ego autem totis viribus meis praeparavi impensas domus Dei mei: aurum ad vasa aurea et argentum in argentea, aes in aenea, ferrum in ferrea, ligna ad lignea, lapides onychinos et ad inserendum, durum caementum et lapides diversorum colorum omnemque pretiosum lapidem et marmor Parium abundantissime.
1CHR|29|3|Et super haec, cum delectarer super domo Dei mei, de peculio meo aurum et argentum do in templum Dei mei, exceptis his, quae paravi in aedem sanctam:
1CHR|29|4|tria milia talenta auri de auro Ophir et septem milia talentorum argenti probatissimi ad operiendos parietes templi;
1CHR|29|5|et ubicumque opus est aurum pro aureis, et ubicumque opus est argentum pro argenteis et pro quolibet opere per manus artificum; et si quis sponte offert, impleat manum suam hodie et offerat, quod voluerit, Domino ".
1CHR|29|6|Sponte obtulerunt itaque principes familiarum et proceres tribuum Israel, tribuni quoque et centuriones et principes operis regis;
1CHR|29|7|dederuntque in opera domus Dei auri talenta quinque milia et solidos decem milia, argenti talenta decem milia et aeris talenta decem et octo milia, ferri quoque centum milia talentorum.
1CHR|29|8|Et apud quemcumque inventi sunt lapides, dederunt in thesaurum domus Domini in manum Iahiel Gersonitis.
1CHR|29|9|Laetatusque est populus super prompto animo eorum, quia corde toto offerebant ea Domino; sed et David rex laetatus est gaudio magno.
1CHR|29|10|Et benedixit Domino coram universa multitudine et ait: Benedictus es, Domine, Deus Israel patris nostri,ab aeterno in aeternum.
1CHR|29|11|Tua est, Domine, magnificentia et potentia,gloria, splendor atque maiestas.Cuncta enim, quae in caelo sunt et in terra, tua sunt.Tuum, Domine, regnum, et tu elevaris ut caput super omnia.
1CHR|29|12|De te sunt divitiae et gloria,tu dominaris omnium.In manu tua virtus et potentia,in manu tua est magnificare et firmare omnia.
1CHR|29|13|Nunc igitur, Deus noster, confitemur tibiet laudamus nomen tuum inclitum.
1CHR|29|14|Quis ego, et quis populus meus, ut possimus haec tibi universa offerre? Tua sunt haec omnia; et, quae de manu tua accepimus, dedimus tibi.
1CHR|29|15|Peregrini enim sumus coram te et advenae, sicut omnes patres nostri; dies nostri quasi umbra super terram, et nulla est spes.
1CHR|29|16|Domine Deus noster, omnis haec copia, quam paravimus, ut aedificaretur domus nomini sancto tuo, de manu tua est, et tua sunt omnia.
1CHR|29|17|Scio, Deus meus, quod probes corda et simplicitatem diligas; unde et ego in simplicitate cordis mei laetus obtuli universa haec et populum tuum, qui hic repertus est, vidi cum ingenti gaudio sponte tibi offerre donaria.
1CHR|29|18|Domine, Deus Abraham et Isaac et Israel patrum nostrorum, custodi in aeternum hanc voluntatem cordis eorum; et semper in venerationem tui mens ista permaneat.
1CHR|29|19|Salomoni quoque filio meo da cor perfectum, ut custodiat mandata tua, testimonia tua et legitima tua et faciat universa et aedificet aedem, cuius impensas paravi ".
1CHR|29|20|Praecepit autem David universae ecclesiae: " Benedicite Domino Deo vestro! ". Et benedixit omnis ecclesia Domino, Deo patrum suorum; et inclinaverunt se et adoraverunt Deum et deinde regem.
1CHR|29|21|Immolaveruntque victimas Domino et obtulerunt holocausta die sequenti, tauros mille, arietes mille, agnos mille cum libaminibus suis et sacrificia abundantissime in omnem Israel.
1CHR|29|22|Et comederunt et biberunt coram Domino in die illo cum grandi laetitia; et fecerunt regem secundo Salomonem filium David atque unxerunt Domino in principem et Sadoc in pontificem.
1CHR|29|23|Seditque Salomon super solium Domini, ut esset rex pro David patre suo, et prosperatus est, et paruit illi omnis Israel.
1CHR|29|24|Sed et universi principes et fortes et cuncti filii regis David dederunt manum subicientes se Salomoni regi.
1CHR|29|25|Magnificavit ergo Dominus Salomonem in excelsum in conspectu omnis Israel et dedit illi gloriam regni, qualem nullus habuit ante eum rex Israel.
1CHR|29|26|Igitur David filius Isai regnavit super universum Israel;
1CHR|29|27|et dies, quibus regnavit super Israel, fuerunt quadraginta anni: in Hebron regnavit septem annis et in Ierusalem annis triginta tribus.
1CHR|29|28|Et mortuus est in senectute bona plenus dierum et divitiis et gloria; et regnavit Salomon filius eius pro eo.
1CHR|29|29|Gesta autem David regis priora et novissima scripta sunt in libro Samuel videntis et in libro Nathan prophetae atque in volumine Gad videntis,
1CHR|29|30|universique regni eius et fortitudinis et temporum, quae transierunt sub eo sive in Israel sive in cunctis regnis terrarum.
2CHR|1|1|Confortatus est ergo Salomon filius David in regno suo, et Dominus Deus eius erat cum eo et magnificavit eum in excelsum.
2CHR|1|2|Praecepitque Salomon universo Israeli, tribunis et centurionibus et iudicibus et ducibus omnis Israel et principibus familiarum
2CHR|1|3|et abiit cum universa multitudine in excelsum Gabaon, ubi erat tabernaculum conventus Dei, quod fecit Moyses famulus Dei in solitudine.
2CHR|1|4|Arcam autem Dei adduxerat David de Cariathiarim in locum, quem praeparaverat ei et ubi fixerat illi tabernaculum, hoc est in Ierusalem;
2CHR|1|5|altare quoque aeneum, quod fabricatus fuerat Beseleel filius Uri filii Hur, ibi erat coram tabernaculo Domini; ibique requisivit eum Salomon et omnis ecclesia.
2CHR|1|6|Ascenditque ibi Salomon ad altare aeneum coram tabernaculo conventus Domini et obtulit in eo mille hostias.
2CHR|1|7|Ecce autem in ipsa nocte apparuit ei Deus dicens: " Postula, quod vis, ut dem tibi ".
2CHR|1|8|Dixitque Salomon Deo: " Tu fecisti cum David patre meo misericordiam magnam et constituisti me regem pro eo.
2CHR|1|9|Nunc ergo, Domine Deus, impleatur sermo tuus, quem pollicitus es David patri meo; tu enim me fecisti regem super populum tuum multum, qui tam innumerabilis est quam pulvis terrae.
2CHR|1|10|Da mihi sapientiam et intellegentiam, ut ingrediar et egrediar coram populo tuo; quis enim potest hunc populum tuum digne, qui tam grandis est, iudicare? ".
2CHR|1|11|Dixit autem Deus ad Salomonem: " Quia hoc magis placuit cordi tuo et non postulasti divitias et substantiam et gloriam neque animas eorum, qui te oderant, sed nec dies vitae plurimos, petisti autem sapientiam et scientiam, ut iudicare possis populum meum, super quem constitui te regem,
2CHR|1|12|sapientia et scientia data sunt tibi; divitias autem et substantiam et gloriam dabo tibi, ita ut nullus in regibus nec ante te nec post te fuerit similis tui ".
2CHR|1|13|Venit ergo Salomon ab excelso Gabaon in Ierusalem coram tabernaculo conventus et regnavit super Israel.
2CHR|1|14|Congregavitque sibi currus et equites, et facti sunt ei mille quadringenti currus et duodecim milia equitum, et fecit eos esse in urbibus quadrigarum et cum rege in Ierusalem.
2CHR|1|15|Praebuitque rex argentum et aurum in Ierusalem quasi lapides et cedros quasi sycomoros, quae nascuntur in Sephela multitudine magna.
2CHR|1|16|Adducebantur autem ei equi de Aegypto et de Coa; negotiatores regis de Coa emebant pretio
2CHR|1|17|et faciebant ascendere et exire de Aegypto quadrigam sescentis argenteis et equum centum quinquaginta; similiter universis regibus Hetthaeorum et Syriae per manus suas educebant.
2CHR|1|18|Decrevit autem Salomon aedificare domum nomini Domini et palatium sibi.
2CHR|2|1|Et numeravit septuaginta milia virorum portantium umeris et octoginta milia, qui caederent lapides in montibus, praepositosque eorum tria milia sescentos.
2CHR|2|2|Misit quoque ad Hiram regem Tyri dicens: " Sicut egisti cum David patre meo et misisti ei ligna cedrina, ut aedificaret sibi domum ad habitandum in ea,
2CHR|2|3|sic fac mecum, ut aedificem domum nomini Domini Dei mei, ut consecrem eam ad adolendum coram illo fumiganda aromata et ad propositionem panum sempiternam et ad holocautomata mane et vespere, sabbatis quoque et neomeniis et sollemnitatibus Domini Dei nostri in sempiternum, quae mandata sunt Israeli.
2CHR|2|4|Domus enim, quam aedificare cupio, magna est; magnus est enim Deus noster super omnes deos.
2CHR|2|5|Quis ergo poterit praevalere, ut aedificet ei dignam domum? Si caelum et caeli caelorum capere eum nequeunt, quantus ego sum, ut possim aedificare ei domum? Sed ad hoc tantum, ut adoleatur incensum coram illo.
2CHR|2|6|Mitte ergo mihi virum eruditum, qui noverit operari in auro et argento, aere et ferro, purpura, coccino et hyacintho, et qui sciat sculpere caelaturas cum his artificibus, quos mecum habeo in Iudaea et Ierusalem, quos praeparavit David pater meus.
2CHR|2|7|Sed et ligna cedrina mitte mihi et arceuthina et pinea de Libano; scio enim quod servi tui noverint caedere ligna de Libano, et erunt servi mei cum servis tuis,
2CHR|2|8|ut parentur mihi ligna plurima; domus enim, quam cupio aedificare, magna erit nimis et inclita.
2CHR|2|9|Praeterea operariis, qui caesuri sunt ligna, servis tuis dabo in cibaria tritici choros viginti milia et hordei choros totidem et vini viginti milia batos, olei quoque batos viginti milia ".
2CHR|2|10|Dixit autem Hiram rex Tyri per litteras, quas miserat Salomoni: " Quia dilexit Dominus populum suum, idcirco te regnare fecit super eum ".
2CHR|2|11|Et addidit dicens: " Benedictus Dominus, Deus Israel, qui fecit caelum et terram, qui dedit David regi filium sapientem et eruditum et sensatum atque prudentem, ut aedificaret domum Domino et palatium sibi.
2CHR|2|12|Misi ergo tibi virum prudentem et scientissimum Hiram magistrum meum,
2CHR|2|13|filium mulieris de filiabus Dan, cuius pater fuit Tyrius, qui novit operari in auro et argento, aere et ferro et lapidibus et lignis, in purpura quoque et hyacintho et bysso et coccino, et qui scit caelare omnem sculpturam et adinvenire prudenter, quodcumque in opere necessarium est, cum artificibus tuis et cum artificibus domini mei David patris tui.
2CHR|2|14|Triticum ergo et hordeum et oleum et vinum, quae pollicitus es, domine mi, mitte servis tuis.
2CHR|2|15|Nos autem caedemus ligna de Libano, quot necessaria habueris, et applicabimus ea ratibus per mare in Ioppe; tuum autem erit transferre ea in Ierusalem ".
2CHR|2|16|Numeravit igitur Salomon omnes viros peregrinos, qui erant in terra Israel post dinumerationem, quam dinumeravit David pater eius; et inventi sunt centum quinquaginta milia et tria milia sescenti.
2CHR|2|17|Fecitque ex eis septuaginta milia, qui umeris onera portarent, et octoginta milia, qui lapides in montibus caederent; tria autem milia et sescentos praepositos operum populi.
2CHR|3|1|Et coepit Salomon aedificare domum Domini in Ierusalem in monte Moria, qui demonstratus fuerat a David patre eius, in loco, quem paraverat David in area Ornan Iebusaei.
2CHR|3|2|Coepit autem aedificare mense secundo anno quarto regni sui.
2CHR|3|3|Et hae sunt mensurae, quas statuit Salomon, ut aedificaret domum Dei: longitudinis cubiti in mensura prima sexaginta, latitudinis cubiti viginti.
2CHR|3|4|Porticum vero ante frontem, quae tendebatur in longum, iuxta mensuram latitudinis domus, cubitorum viginti; porro altitudo centum viginti cubitorum erat. Et deauravit eam intrinsecus auro mundissimo.
2CHR|3|5|Domum quoque maiorem texit tabulis ligneis abiegnis et laminas auri obryzi affixit per totum; scalpsitque in eis palmas et quasi catenulas se invicem complectentes.
2CHR|3|6|Stravit quoque pavimentum templi pretiosissimo marmore decore multo.
2CHR|3|7|Porro aurum erat de Parvaim, de cuius laminis texit domum, et trabes eius et postes et parietes et ostia; et caelavit cherubim in parietibus.
2CHR|3|8|Fecit quoque domum sancti sanctorum: longitudinem iuxta latitudinem domus cubitorum viginti et latitudinem similiter viginti cubitorum; et laminis auri optimi texit eam quasi talentis sescentis.
2CHR|3|9|Sed et pro clavis usus est auro ponderis quinquaginta siclorum. Cenacula quoque texit auro.
2CHR|3|10|Fecit etiam in domo sancti sanctorum cherubim duos opere statuario et texit eos auro.
2CHR|3|11|Alae cherubim viginti cubitis extendebantur, ita ut una ala haberet cubitos quinque et tangeret parietem domus, et altera quinque cubitos habens alam tangeret alterius cherub.
2CHR|3|12|Similiter cherub alterius ala quinque habebat cubitos et tangebat parietem, et ala eius altera quinque cubitorum alam cherub alterius contingebat.
2CHR|3|13|Igitur alae utriusque cherubim expansae erant et extendebantur per cubitos viginti; ipsi autem stabant erectis pedibus, et facies eorum erant versae ad exteriorem domum.
2CHR|3|14|Fecit quoque velum ex hyacintho, purpura, cocco et bysso et intexuit ei cherubim.
2CHR|3|15|Ante fores etiam templi duas columnas, quae triginta et quinque cubitos habebant altitudinis; porro capita earum quinque cubitorum.
2CHR|3|16|Necnon et quasi catenulas in torque, et superposuit eas capitibus columnarum; malogranata etiam centum, quae catenulis interposuit.
2CHR|3|17|Ipsas quoque columnas posuit ante faciem templi, unam a dextris et alteram a sinistris; eam, quae a dextris erat, vocavit Iachin et, quae ad laevam, Booz.
2CHR|4|1|Fecit quoque altare aeneum viginti cubitorum longitudinis et viginti cubitorum latitudinis et decem cubitorum
2CHR|4|2|altitudinis. Mare etiam fusile decem cubitis a labio usque ad labium rotundum per circuitum; quinque cubitos habebat altitudinis, et funiculus triginta cubitorum ambiebat gyrum eius.
2CHR|4|3|Similitudo quoque boum erat subter illud, in circuitu circumdabant illud decem cubitis - duobus versibus alvum maris circuibant boves fusiles in una fusione cum mari.
2CHR|4|4|Et ipsum mare super duodecim boves impositum erat, quorum tres respiciebant aquilonem et alii tres occidentem, porro tres alii meridiem et tres, qui reliqui erant, orientem habentes mare superpositum; posteriora autem boum erant intrinsecus sub mari.
2CHR|4|5|Porro vastitas eius habebat mensuram palmi, et labium illius erat quasi labium calicis vel repandi lilii; capiebatque tria milia batos.
2CHR|4|6|Fecit quoque luteres decem et posuit quinque a dextris et quinque a sinistris, ut lavarent in eis omnia, quae in holocaustum oblaturi erant; porro in mari sacerdotes lavabantur.
2CHR|4|7|Fecit autem et candelabra aurea decem secundum speciem, qua iussa erant fieri, et posuit ea in templo quinque a dextris et quinque a sinistris.
2CHR|4|8|Necnon et mensas decem, et posuit eas in templo quinque a dextris et quinque a sinistris; phialas quoque aureas centum.
2CHR|4|9|Fecit etiam atrium sacerdotum et atrium grande et ostia in atrio, quae texit aere.
2CHR|4|10|Porro mare posuit in latere dextro contra orientem ad meridiem.
2CHR|4|11|Fecit autem Hiram lebetes et vatilla et phialas et complevit omne opus regis Salomonis in domo Dei;
2CHR|4|12|hoc est columnas duas et globos et capitella super caput columnarum duarum et serta duo, quae tegerent globos capitellorum;
2CHR|4|13|malogranata quoque quadringenta et serta duo, ita ut bini ordines malogranatorum singulis sertis iungerentur, quae protegerent globos capitellorum columnarum.
2CHR|4|14|Bases etiam fecit et luteres, quos superposuit basibus,
2CHR|4|15|mare unum, boves quoque duodecim sub mari;
2CHR|4|16|et lebetes et vatilla et fuscinulas: omnia vasa fecit regi Salomoni Hiram magister eius pro domo Domini ex aere mundissimo.
2CHR|4|17|In regione Iordanis fudit ea rex in argillosa terra inter Succoth et Saredatha.
2CHR|4|18|Fecitque Salomon multitudinem vasorum innumerabilem, ita ut ignoraretur pondus aeris.
2CHR|4|19|Fecitque Salomon omnia vasa domus Dei et altare aureum et mensas et super eas panes propositionis;
2CHR|4|20|candelabra quoque cum lucernis suis, ut lucerent ante Dabir iuxta ritum, ex auro purissimo,
2CHR|4|21|et florem et lucernas et forcipes aureos: omnia de auro perfectissimo facta sunt;
2CHR|4|22|cultros quoque et phialas et sartagines et turibula ex auro purissimo. Et ostia templi interiora in sancta sanctorum et ostia templi forinsecus aurea.
2CHR|5|1|Sicque completum est omne opus, quod fecit Salomon in do mo Domini. Intulit igitur Salomon omnia, quae voverat David pater suus, argentum et aurum, et universa vasa posuit in thesauris domus Dei.
2CHR|5|2|Post quae congregavit maiores natu Israel et cunctos principes tribuum et capita familiarum de filiis Israel in Ierusalem, ut adducerent arcam foederis Domini de civitate David, quae est Sion.
2CHR|5|3|Venerunt igitur ad regem omnes viri Israel in die sollemni mensis septimi.
2CHR|5|4|Cumque venissent cuncti seniorum Israel, portaverunt Levitae arcam
2CHR|5|5|et intulerunt eam et tabernaculum conventus et omnem paraturam tabernaculi. Porro omnia vasa sanctuarii, quae erant in tabernaculo, portaverunt sacerdotes levitici generis.
2CHR|5|6|Rex autem Salomon et universus coetus Israel, omnes, qui fuerunt congregati ad eum ante arcam, immolabant oves et boves absque ullo numero: tanta enim erat multitudo victimarum.
2CHR|5|7|Et intulerunt sacerdotes arcam foederis Domini in locum suum ad Dabir templi, in sancta sanctorum subter alas cherubim,
2CHR|5|8|ita ut cherubim expanderent alas suas super locum, in quo posita erat arca, et ipsam arcam tegerent cum vectibus suis ab alto.
2CHR|5|9|Vectium autem, quibus portabatur arca, quia paululum longiores erant, capita parebant ante Dabir; si vero quis erat extrinsecus eos videre non poterat. Fuit itaque arca ibi usque in praesentem diem.
2CHR|5|10|Nihilque erat aliud in arca, nisi duae tabulae, quas posuerat Moyses in Horeb, quando fecit Dominus foedus cum filiis Israel egredientibus ex Aegypto.
2CHR|5|11|Egressis autem sacerdotibus de sanctuario - omnes enim sacerdotes, qui ibi potuerant inveniri, sanctificati sunt, non observantes vices et ministeriorum ordinem,
2CHR|5|12|et Levitae cantores, omnes, qui sub Asaph erant et qui sub Heman et qui sub Idithun, filii et fratres eorum, vestiti byssinis, cymbalis et psalteriis et citharis stabant ad orientalem plagam altaris, et cum eis sacerdotes centum viginti canentes tubis -
2CHR|5|13|igitur cunctis pariter et tubis et voce et cymbalis et organis et diversi generis musicorum concinentibus et vocem in sublime tollentibus, cum una voce Dominum laudare coepissent et dicere: " Confitemini Domino quoniam bonus, quoniam in aeternum misericordia eius ", impleta est domus Dei nube,
2CHR|5|14|nec potuerunt sacerdotes stare et ministrare propter nubem; compleverat enim gloria Domini domum Dei.
2CHR|6|1|Tunc Salomon ait: " Dominus pollicitus est, ut habitaret in ca ligine;
2CHR|6|2|ego autem aedificavi domum in habitaculum tuum, ut habitares ibi in perpetuum ".
2CHR|6|3|Et convertit rex faciem suam et benedixit universae multitudini Israel - nam omnis turba stabat intenta - et ait:
2CHR|6|4|" Benedictus Dominus, Deus Israel, qui, quod locutus est ore suo David patri meo, opere complevit dicens:
2CHR|6|5|"A die qua eduxi populum meum de terra Aegypti non elegi civitatem de cunctis tribubus Israel, ut aedificaretur in ea domus nomini meo, neque elegi quemquam alium virum, ut esset dux in populo meo Israel,
2CHR|6|6|sed elegi Ierusalem, ut sit nomen meum in ea, et elegi David, ut constituerem eum super populum meum Israel".
2CHR|6|7|Cumque fuisset voluntatis David patris mei, ut aedificaret domum nomini Domini, Dei Israel,
2CHR|6|8|dixit Dominus ad eum: "Quia haec fuit voluntas tua, ut aedificares domum nomini meo, bene quidem fecisti huiuscemodi habere voluntatem,
2CHR|6|9|sed non tu aedificabis domum, verum filius tuus, qui egredietur de lumbis tuis, ipse aedificabit domum nomini meo".
2CHR|6|10|Complevit ergo Dominus sermonem suum, quem locutus fuerat, et ego surrexi pro David patre meo et sedi super thronum Israel, sicut locutus est Dominus, et aedificavi domum nomini Domini, Dei Israel;
2CHR|6|11|et posui in ea arcam, in qua est pactum Domini, quod pepigit cum filiis Israel ".
2CHR|6|12|Stetit ergo coram altari Domini ex adverso universae multitudinis Israel et extendit manus suas.
2CHR|6|13|Siquidem fecerat Salomon basim aeneam et posuerat eam in medio atrii habentem quinque cubitos longitudinis et quinque cubitos latitudinis et tres cubitos altitudinis, stetitque super eam; et deinceps, flexis genibus contra universam multitudinem Israel et palmis in caelum levatis,
2CHR|6|14|ait: " Domine, Deus Israel, non est similis tui Deus in caelo et in terra, qui custodis pactum et misericordiam cum servis tuis, qui ambulant coram te in toto corde suo,
2CHR|6|15|qui praestitisti servo tuo David patri meo quaecumque locutus fueras ei, et, quae ore promiseras, opere complesti, sicut et praesens tempus probat.
2CHR|6|16|Nunc ergo, Domine, Deus Israel, imple servo tuo patri meo David, quaecumque locutus es dicens: "Non deficiet ex te vir coram me, qui sedeat super thronum Israel, ita tamen si custodierint filii tui vias suas et ambulaverint in lege mea, sicut et tu ambulasti coram me".
2CHR|6|17|Et nunc, Domine, Deus Israel, firmetur sermo tuus, quem locutus es servo tuo David!
2CHR|6|18|Ergone credibile est, ut habitet Deus cum hominibus super terram? Si caelum et caeli caelorum non te capiunt, quanto magis domus ista, quam aedificavi!
2CHR|6|19|Sed respice orationem servi tui et obsecrationem eius, Domine Deus meus, et audi clamorem et preces, quas fundit famulus tuus coram te,
2CHR|6|20|ut aperias oculos tuos super domum istam diebus ac noctibus, super locum in quo pollicitus es, ut ponas nomen tuum et exaudires orationem, quam servus tuus orat in eo.
2CHR|6|21|Et exaudi preces famuli tui et populi tui Israel, qui oraverint ad locum istum; exaudi de habitaculo tuo, de caelis, exaudi et propitiare!
2CHR|6|22|Si peccaverit quispiam in proximum suum, et ille exegerit ab eo iuramentum, ut se maledicto constringat coram altari in domo ista,
2CHR|6|23|tu audies de caelo et facies iudicium servorum tuorum, ita ut reddas iniquo viam suam in caput proprium et ulciscaris iustum retribuens ei secundum iustitiam suam.
2CHR|6|24|Si superatus fuerit populus tuus Israel ab inimicis, quia peccaturi sunt tibi, et conversi egerint paenitentiam et confitentes nomini tuo oraverint et fuerint deprecati in domo ista,
2CHR|6|25|tu exaudies de caelo, et propitiare peccato populi tui Israel et reduc eos in terram, quam dedisti eis et patribus eorum.
2CHR|6|26|Si clauso caelo pluvia non fluxerit propter peccata populi, et deprecati te fuerint in loco isto et confessi nomini tuo et conversi a peccatis suis, cum eos afflixeris,
2CHR|6|27|exaudi de caelo, Domine, et dimitte peccata servorum tuorum et populi tui Israel, doce eos viam bonam, per quam ingrediantur, et da pluviam terrae, quam dedisti populo tuo ad possidendum.
2CHR|6|28|Fames si orta fuerit in terra et pestilentia, uredo et aurugo et locusta et bruchus et hostes, vastatis regionibus, portas eius obsederint, omnisque plaga et infirmitas presserit,
2CHR|6|29|si quis de populo tuo Israel fuerit deprecatus cognoscens plagam et infirmitatem suam et expanderit manus suas ad domum hanc,
2CHR|6|30|tu exaudi de caelo, de loco habitationis tuae, et propitiare et redde unicuique secundum vias suas, quia nosti cor eius; tu enim solus nosti corda filiorum hominum,
2CHR|6|31|ut timeant te et ambulent in viis tuis cunctis diebus, quibus vivunt super faciem terrae, quam dedisti patribus nostris.
2CHR|6|32|Externum quoque, qui non est de populo tuo Israel, si venerit de terra longinqua propter nomen tuum magnum et propter manum tuam robustam et brachium tuum extentum, et oraverit in loco isto,
2CHR|6|33|tu exaudies de caelo firmissimo habitaculo tuo et facies cuncta, pro quibus invocaverit te ille peregrinus, ut sciant omnes populi terrae nomen tuum et timeant te sicut populus tuus Israel et cognoscant quia nomen tuum invocatum est super domum hanc, quam aedificavi.
2CHR|6|34|Si egressus fuerit populus tuus ad bellum contra adversarios suos per viam, in qua miseris eos, et oraverint te contra viam, in qua civitas haec est, quam elegisti, et domus, quam aedificavi nomini tuo,
2CHR|6|35|tu exaudies de caelo preces eorum et obsecrationem, et facies iudicium eorum.
2CHR|6|36|Si autem peccaverint tibi - neque enim est homo, qui non peccet - et iratus fueris eis et tradideris hostibus, et captivos duxerint eos in terram longinquam vel propinquam,
2CHR|6|37|et conversi in corde suo in terra, ad quam captivi ducti fuerant, egerint paenitentiam et deprecati te fuerint in terra captivitatis suae dicentes: "Peccavimus, inique fecimus, iniuste egimus";
2CHR|6|38|et reversi fuerint ad te in toto corde suo et in tota anima sua in terra captivitatis suae, ad quam ducti sunt, et oraverint te contra viam terrae suae, quam dedisti patribus eorum, et urbis, quam elegisti, et domus, quam aedificavi nomini tuo,
2CHR|6|39|ut exaudias de caelo, de loco habitationis tuae, preces eorum et supplicationes eorum et facias iudicium et dimittas populo tuo, qui peccavit tibi;
2CHR|6|40|tu es enim Deus meus. Aperiantur, quaeso, oculi tui, et aures tuae intentae sint ad orationem, quae fit in loco isto.
2CHR|6|41|Nunc igitur consurge, Domine Deus, in requiem tuam, tu et arca fortitudinis tuae; sacerdotes tui, Domine Deus, induantur salutem, et sancti tui laetentur in bonis.
2CHR|6|42|Domine Deus, ne averteris faciem christi tui; memento misericordiarum David servi tui ".
2CHR|7|1|Cumque complesset Salomon fundens preces, ignis descendit de caelo et devoravit holocaustum et victimas, et maiestas Domini implevit domum.
2CHR|7|2|Nec poterant sacerdotes ingredi templum Domini, eo quod implesset maiestas Domini templum Domini.
2CHR|7|3|Sed et omnes filii Israel videbant descendentem ignem et gloriam Domini super domum et corruentes proni in terram super pavimentum stratum lapide adoraverunt et laudaverunt Dominum: " Quoniam bonus, quoniam in saeculum misericordia eius ".
2CHR|7|4|Rex autem et omnis populus immolabant victimas coram Domino.
2CHR|7|5|Mactavit igitur rex Salomon hostias boum viginti duo milia, ovium centum viginti milia, et dedicavit domum Dei rex et universus populus.
2CHR|7|6|Sacerdotes autem stabant in officiis suis et Levitae in organis carminum Domini, quae fecit David rex ad laudandum Dominum: " Quoniam in aeternum misericordia eius ", hymnos David canentes per manus suas. Porro sacerdotes canebant tubis ante eos, cunctusque Israel stabat.
2CHR|7|7|Sanctificavit quoque Salomon medium atrii ante templum Domini; obtulerat enim ibi holocausta et adipes pacificorum, quia altare aeneum, quod fecerat, non poterat sustinere holocausta et oblationes et adipes.
2CHR|7|8|Fecit ergo Salomon sollemnitatem in tempore illo septem diebus, et omnis Israel cum eo, ecclesia magna valde ab introitu Emath usque ad torrentem Aegypti.
2CHR|7|9|Feceruntque die octavo collectam magnam, eo quod dedicassent altare septem diebus et sollemnitatem celebrassent diebus septem.
2CHR|7|10|Igitur in die vicesimo tertio mensis septimi dimisit populum ad tabernacula sua, laetantem atque gaudentem super bono, quod fecerat Dominus Davidi et Salomoni et Israeli populo suo.
2CHR|7|11|Complevitque Salomon domum Domini et domum regis; et in omnibus, quae disposuerat in corde suo, ut faceret in domo Domini et in domo sua, prosperatus est.
2CHR|7|12|Apparuit autem ei Dominus nocte et ait: " Audivi orationem tuam et elegi locum istum mihi in domum sacrificii.
2CHR|7|13|Si clausero caelum, et pluvia non fluxerit, et mandavero et praecepero locustae, ut devoret terram, et misero pestilentiam in populum meum,
2CHR|7|14|humiliatus autem populus meus, super quos invocatum est nomen meum, deprecatus me fuerit et exquisierit faciem meam et egerit paenitentiam a viis suis pessimis, ego exaudiam de caelo et propitius ero peccatis eorum et sanabo terram eorum.
2CHR|7|15|Nunc oculi mei erunt aperti, et aures meae attentae ad orationem eius, qui in loco isto oraverit;
2CHR|7|16|elegi enim et sanctificavi locum istum, ut sit nomen meum ibi in sempiternum, et permaneant oculi mei et cor meum ibi cunctis diebus.
2CHR|7|17|Tu quoque, si ambulaveris coram me, sicut ambulavit David pater tuus, et feceris iuxta omnia, quae praecepi tibi, et decreta et iudicia mea servaveris,
2CHR|7|18|stabiliam thronum regni tui, sicut pollicitus sum David patri tuo dicens: Non auferetur de stirpe tua vir, qui sit princeps in Israel.
2CHR|7|19|Si autem aversi fueritis et dereliqueritis decreta mea et praecepta mea, quae proposui vobis, et abeuntes servieritis diis alienis et adoraveritis eos,
2CHR|7|20|evellam vos de terra mea, quam dedi vobis, et domum hanc, quam sanctificavi nomini meo, proiciam a facie mea et tradam eam in parabolam et in fabulam cunctis populis.
2CHR|7|21|Et super domo ista, quae erat excelsa, universi transeuntes stupebunt et dicent: "Quare fecit Dominus sic terrae huic et domui huic?".
2CHR|7|22|Respondebuntque: "Quia dereliquerunt Dominum, Deum patrum suorum, qui eduxit eos de terra Aegypti, et apprehenderunt deos alienos et adoraverunt eos et coluerunt, idcirco venerunt super eos universa haec mala" ".
2CHR|8|1|Expletis autem viginti annis, postquam aedificavit Salomon domum Domini et domum suam,
2CHR|8|2|civitates, quas dederat Hiram Salomoni, aedificavit et habitare ibi fecit filios Israel.
2CHR|8|3|Abiit quoque in Emath Soba et obtinuit eam.
2CHR|8|4|Et aedificavit Palmyram in deserto et omnes civitates horreorum, quas aedificavit in Emath.
2CHR|8|5|Exstruxitque Bethoron superiorem et Bethoron inferiorem, civitates munitas habentes muros et portas et vectes,
2CHR|8|6|Baalath etiam et omnes urbes horreorum, quae fuerunt Salomonis, cunctasque urbes quadrigarum et urbes equorum. Omnia quaecumque voluit Salomon atque disposuit, aedificavit in Ierusalem et in Libano et in universa terra potestatis suae.
2CHR|8|7|Omnem populum, qui derelictus fuerat de Hetthaeis et Amorraeis et Pherezaeis et Hevaeis et Iebusaeis, qui non erant de stirpe Israel,
2CHR|8|8|de filiis eorum, qui remanserant post eos in terra, quos non interfecerant filii Israel, subiugavit Salomon in tributarios usque in diem hanc.
2CHR|8|9|Porro de filiis Israel non posuit, ut servirent operibus regis; ipsi enim erant viri bellatores et principes pugnatorum eius et principes quadrigarum et equitum eius.
2CHR|8|10|Omnes autem principes praefectorum regis Salomonis fuerunt ducenti quinquaginta, qui praefuerant populo.
2CHR|8|11|Filiam vero pharaonis transtulit de civitate David in domum, quam aedificaverat ei; dixit enim rex: " Non habitabit mulier mihi in domo David regis Israel, eo quod sanctificata sit, quia ingressa est in eam arca Domini ".
2CHR|8|12|Tunc obtulit Salomon holocausta Domino super altare Domini, quod exstruxerat ante porticum,
2CHR|8|13|ut per singulos dies offerretur in eo iuxta praeceptum Moysi in sabbatis et in calendis et in festis diebus ter per annum, id est in sollemnitate Azymorum et in sollemnitate Hebdomadarum et in sollemnitate Tabernaculorum.
2CHR|8|14|Et constituit iuxta dispositionem David patris sui officia sacerdotum in ministeriis suis et Levitas in ordine suo, ut laudarent et ministrarent coram sacerdotibus iuxta ritum uniuscuiusque diei, et ianitores in divisionibus suis per portam et portam; sic enim praeceperat David homo Dei.
2CHR|8|15|Nec praetergressi sunt mandata regis de sacerdotibus et Levitis in omnibus et in custodiis thesaurorum.
2CHR|8|16|Et firmatum est totum opus Salomonis ex eo die, quo fundavit domum Domini, usque in diem, quo perfecit eam.
2CHR|8|17|Tunc abiit Salomon in Asiongaber et in Ailath ad oram maris Rubri, quae est in terra Edom.
2CHR|8|18|Misit autem ei Hiram per manus servorum suorum naves et nautas gnaros maris; et abierunt cum servis Salomonis in Ophir tuleruntque inde quadringenta quinquaginta talenta auri et attulerunt ad regem Salomonem.
2CHR|9|1|Regina quoque Saba, cum audisset famam Salomonis, venit, ut tentaret eum in aenigmatibus in Ierusalem cum magno comitatu et camelis, qui portabant aromata et auri plurimum gemmasque pretiosas. Cumque venisset ad Salomonem, locuta est ei, quaecumque erant in corde suo.
2CHR|9|2|Et exposuit ei Salomon omnia, quae proposuerat, nec quidquam fuit quod ei non perspicuum fecerit.
2CHR|9|3|Quae postquam vidit, sapientiam scilicet Salomonis et domum, quam aedificaverat,
2CHR|9|4|necnon et cibaria mensae eius et sessionem servorum et officia ministrorum eius et vestimenta eorum, pincernas quoque et vestes eorum et victimas, quas immolabat in domo Domini, non erat prae stupore ultra in ea spiritus.
2CHR|9|5|Dixitque ad regem: " Verus est sermo, quem audieram in terra mea, de rebus tuis et sapientia tua;
2CHR|9|6|non credebam narrantibus, donec ipsa venissem, et vidissent oculi mei, et probassem vix medietatem sapientiae tuae mihi fuisse narratam; vicisti famam, quam audivi.
2CHR|9|7|Beati viri tui et beati servi tui, qui assistunt coram te omni tempore et audiunt sapientiam tuam!
2CHR|9|8|Sit Dominus Deus tuus benedictus, qui voluit te ordinare super thronum suum regem Domini Dei tui! Quia diligit Deus tuus Israel et vult servare eum in aeternum, idcirco posuit te super eum regem, ut facias iudicia atque iustitiam ".
2CHR|9|9|Dedit autem regi centum viginti talenta auri et aromata multa nimis et gemmas pretiosissimas; non fuerunt aromata talia ut haec, quae dedit regina Saba regi Salomoni.
2CHR|9|10|Sed et servi Hiram cum servis Salomonis attulerunt aurum de Ophir et ligna thyina et gemmas pretiosissimas;
2CHR|9|11|et fecit rex de lignis thyinis gradus in domo Domini et in domo regia, citharas quoque et psalteria cantoribus. Numquam visa sunt in terra Iudae ligna talia.
2CHR|9|12|Rex autem Salomon dedit reginae Saba cuncta, quae voluit et quae postulavit, et multo plura quam attulerat ad eum. Quae reversa abiit in terram suam cum servis suis.
2CHR|9|13|Erat autem pondus auri, quod afferebatur Salomoni per singulos annos, sescenta sexaginta sex talenta auri,
2CHR|9|14|excepta ea summa, quae proveniebat ex tributis mercatorum et negotiatorum afferentium et omnium regum Arabiae et ducum terrae, qui comportabant aurum et argentum Salomoni.
2CHR|9|15|Fecit igitur rex Salomon ducenta scuta aurea de summa sescentorum aureorum, qui in singulis scutis expendebantur,
2CHR|9|16|trecentas quoque peltas aureas trecentorum aureorum, quibus tegebantur singulae peltae, posuitque ea rex in domo Saltus Libani.
2CHR|9|17|Fecit quoque rex solium eburneum grande et vestivit illud auro mundissimo;
2CHR|9|18|sex quoque gradus, quibus ascendebatur ad solium, et scabellum aureum et brachiola duo altrinsecus et duos leones stantes iuxta brachiola,
2CHR|9|19|sed et alios duodecim leunculos stantes super sex gradus ex utraque parte; non fuit tale solium in universis regnis.
2CHR|9|20|Omnia quoque vasa convivii regis erant aurea, et vasa domus Saltus Libani ex auro purissimo; argentum enim in diebus Salomonis pro nihilo reputabatur.
2CHR|9|21|Siquidem naves regis ibant in Tharsis cum servis Hiram; semel in annis tribus veniebant naves Tharsis portantes aurum et argentum et ebur et simias et pavos.
2CHR|9|22|Magnificatus est igitur rex Salomon super omnes reges terrae divitiis et sapientia.
2CHR|9|23|Omnesque reges terrarum desiderabant faciem videre Salomonis, ut audirent sapientiam, quam dederat Deus in corde eius,
2CHR|9|24|et deferebant ei munera, vasa argentea et aurea et vestes et arma et aromata, equos et mulos per singulos annos.
2CHR|9|25|Habuit quoque Salomon quattuor milia stabula equorum et curruum equitumque duodecim milia; constituitque eos in urbibus quadrigarum et, ubi erat rex, in Ierusalem.
2CHR|9|26|Exercuit etiam potestatem super cunctos reges, a fluvio Euphrate usque ad terram Philisthinorum et usque ad terminos Aegypti;
2CHR|9|27|tantamque copiam praebuit argenti in Ierusalem quasi lapidum, et cedrorum tantam multitudinem velut sycomororum, quae gignuntur in Sephela.
2CHR|9|28|Adducebantur autem ei equi de Aegypto cunctisque regionibus.
2CHR|9|29|Reliqua vero operum Salomonis priorum et novissimorum scripta sunt in verbis Nathan prophetae et in prophetia Ahiae Silonitis, in visione quoque Addo videntis super Ieroboam filium Nabat.
2CHR|9|30|Regnavit autem Salomon in Ierusalem super omnem Israel quadraginta annis;
2CHR|9|31|dormivitque cum patribus suis, et sepelierunt eum in civitate David patris eius. Regnavitque Roboam filius eius pro eo.
2CHR|10|1|Profectus est autem Roboam in Sichem; illuc enim cunctus Israel convenerat, ut constituerent eum regem.
2CHR|10|2|Quod cum audisset Ieroboam filius Nabat, qui erat in Aegypto - fugerat quippe illuc ante Salomonem - statim reversus est;
2CHR|10|3|vocaveruntque eum, et venit cum universo Israel, et locuti sunt ad Roboam dicentes:
2CHR|10|4|" Pater tuus durissimo iugo nos pressit; tu leviora impera patre tuo, qui nobis gravem imposuit servitutem, et paululum de onere subleva, et serviemus tibi ".
2CHR|10|5|Qui ait: " Post tres dies revertimini ad me ".Cumque abisset populus,
2CHR|10|6|iniit rex Roboam consilium cum senibus, qui steterant coram patre eius Salomone, dum adhuc viveret, dicens: " Quid datis consilii, ut respondeam populo? ".
2CHR|10|7|Qui dixerunt ei: " Si placueris populo huic et lenieris eos verbis clementibus, servient tibi omni tempore ".
2CHR|10|8|At ille reliquit consilium senum et cum iuvenibus tractare coepit, qui cum eo nutriti fuerant et erant in comitatu illius.
2CHR|10|9|Dixitque ad eos: " Quid vobis videtur, vel respondere quid debemus populo huic, qui dixit mihi: "Subleva iugum, quod imposuit nobis pater tuus"? ".
2CHR|10|10|Et responderunt iuvenes, qui nutriti fuerant cum eo, atque dixerunt: " Sic loqueris populo, qui dixit tibi: "Pater tuus aggravavit iugum nostrum, tu subleva", et sic respondebis eis: Minimus digitus meus grossior est lumbis patris mei;
2CHR|10|11|pater meus imposuit vobis iugum grave, et ego maius pondus apponam; pater meus cecidit vos flagellis, ego vero caedam scorpionibus ".
2CHR|10|12|Venit ergo Ieroboam et universus populus ad Roboam die tertio, sicut praeceperat eis rex dicens: "Revertimini ad me die tertio ".
2CHR|10|13|Responditque rex dura, derelicto consilio seniorum;
2CHR|10|14|locutusque est iuxta iuvenum voluntatem: Pater meus grave vobis imposuit iugum,quod ego gravius faciam.Pater meus cecidit vos flagellis,ego vero caedam scorpionibus ".
2CHR|10|15|Et non acquievit populi precibus. Erat enim voluntatis Dei, ut compleretur sermo eius, quem locutus fuerat per manum Ahiae Silonitis ad Ieroboam filium Nabat.
2CHR|10|16|Israel autem universus videns quod noluisset eos audire rex, locutus est ad eum: Non est nobis pars in David,neque hereditas in filio Isai!Revertere in tabernacula tua, Israel!Tu autem vide domum tuam, David! ".Et abiit Israel in tabernacula sua.
2CHR|10|17|Super filios autem Israel, qui habitabant in civitatibus Iudae, regnavit Roboam.
2CHR|10|18|Misitque rex Roboam Adoram, qui praeerat servituti, et lapidaverunt eum filii Israel, et mortuus est. Porro rex Roboam currum festinavit ascendere et fugit in Ierusalem.
2CHR|10|19|Recessitque Israel a domo David usque ad diem hanc.
2CHR|11|1|Venit autem Roboam in Ie rusalem et convocavit univer sam domum Iudae et Beniamin, centum octoginta milia electorum bellantium, ut dimicaret contra Israel et converteret ad se regnum suum.
2CHR|11|2|Factusque est sermo Domini ad Semeiam hominem Dei dicens:
2CHR|11|3|" Loquere ad Roboam filium Salomonis regem Iudae et ad universum Israel, qui est in Iuda et Beniamin:
2CHR|11|4|Haec dicit Dominus: Non ascendetis neque pugnabitis contra fratres vestros. Revertatur unusquisque in domum suam, quia mea hoc gestum est voluntate ". Qui cum audissent sermonem Domini, reversi sunt nec perrexerunt contra Ieroboam.
2CHR|11|5|Habitavit autem Roboam in Ierusalem et aedificavit civitates muratas in Iuda.
2CHR|11|6|Exstruxitque Bethlehem et Etam et Thecue,
2CHR|11|7|Bethsur quoque et Socho et Odollam
2CHR|11|8|necnon Geth et Maresa et Ziph,
2CHR|11|9|sed et Aduram et Lachis et Azeca,
2CHR|11|10|Saraa quoque et Aialon et Hebron, quae erant in Iuda et Beniamin civitates munitissimas.
2CHR|11|11|Cumque clausisset eas muris, posuit in eis principes ciborumque horrea et olei et vini.
2CHR|11|12|Sed et in singulis urbibus fecit armamentarium scutorum et hastarum firmavitque eas summa diligentia et imperavit super Iudam et Beniamin.
2CHR|11|13|Sacerdotes autem et Levitae, qui erant in universo Israel, venerunt ad eum de cunctis sedibus suis.
2CHR|11|14|Levitae relinquentes suburbana et possessiones suas transierunt ad Iudam et Ierusalem, eo quod abiecisset eos Ieroboam et posteri eius, ne sacerdotio Domini fungerentur.
2CHR|11|15|Qui constituit sibi sacerdotes excelsorum et daemoniorum vitulorumque, quos fecerat.
2CHR|11|16|Sed sequentes eos et de cunctis tribubus Israel quicumque dederant cor suum, ut quaererent Dominum, Deum Israel, venerunt Ierusalem ad immolandum victimas Domino, Deo patrum suorum.
2CHR|11|17|Et roboraverunt regnum Iudae et confirmaverunt Roboam filium Salomonis per tres annos; ambulaverunt enim in viis David et Salomonis annis tantum tribus.
2CHR|11|18|Duxit autem Roboam uxorem Mahalath filiam Ierimoth filii David et Abihail filiae Eliab filii Isai,
2CHR|11|19|quae peperit ei filios Iehus et Samariam et Zoom.
2CHR|11|20|Post hanc quoque accepit Maacha filiam Absalom, quae peperit ei Abia et Ethai et Ziza et Salomith.
2CHR|11|21|Amavit autem Roboam Maacha filiam Absalom super omnes uxores suas et concubinas; nam uxores decem et octo duxerat, concubinas autem sexaginta. Et genuit viginti octo filios et sexaginta filias.
2CHR|11|22|Constituit vero in capite Abiam filium Maacha ducem super fratres suos; ipsum enim regem facere cogitabat.
2CHR|11|23|Et sapienter filios suos dispersit in cunctis finibus Iudae et Beniamin in universis civitatibus muratis. Praebuitque eis escas plurimas et multas petivit uxores.
2CHR|12|1|Cumque roboratum fuisset regnum Roboam et conforta tum, dereliquit legem Domini, et omnis Israel cum eo.
2CHR|12|2|Anno autem quinto regni Roboam ascendit Sesac rex Aegypti in Ierusalem - quia peccaverunt Domino -
2CHR|12|3|cum mille ducentis curribus et sexaginta milibus equitum, nec erat numerus vulgi, quod venerat cum eo ex Aegypto, Libyes scilicet et Socciitae et Aethiopes.
2CHR|12|4|Cepitque civitates munitissimas in Iuda et venit usque Ierusalem.
2CHR|12|5|Semeias autem propheta ingressus est ad Roboam et principes Iudae, qui congregati fuerant in Ierusalem fugientes Sesac, dixitque ad eos: " Haec dicit Dominus: Vos reliquistis me, et ego reliqui vos in manu Sesac ".
2CHR|12|6|Humiliatique principes Israel et rex dixerunt: " Iustus est Dominus! ".
2CHR|12|7|Cumque vidisset Dominus quod humiliati essent, factus est sermo Domini ad Semeiam dicens: " Quia humiliati sunt, non disperdam eos daboque eis mox effugium, et non effundetur furor meus super Ierusalem per manum Sesac.
2CHR|12|8|Verumtamen servient ei, ut sciant distantiam servitutis meae et servitutis regni terrarum ".
2CHR|12|9|Ascendit itaque Sesac rex Aegypti in Ierusalem, sublatis thesauris domus Domini et domus regis; omniaque secum tulit et clipeos aureos, quos fecerat Salomon.
2CHR|12|10|Pro quibus fecit rex Roboam aeneos et tradidit illos principibus cursorum, qui custodiebant vestibulum palatii.
2CHR|12|11|Cumque introiret rex domum Domini, veniebant cursores et tollebant eos; iterumque referebant eos ad armamentarium suum.
2CHR|12|12|Verumtamen, quia humiliatus est, aversa est ab eo ira Domini, nec deletus est penitus; siquidem et in Iuda inventa sunt opera bona.
2CHR|12|13|Confortatus est igitur rex Roboam in Ierusalem atque regnavit. Quadraginta autem et unius anni erat, cum regnare coepisset, et decem septemque annis regnavit in Ierusalem urbe, quam elegit Dominus, ut confirmaret nomen suum ibi de cunctis tribubus Israel. Nomenque matris eius Naama Ammanitis.
2CHR|12|14|Fecit autem malum et non praeparavit cor suum, ut quaereret Dominum.
2CHR|12|15|Opera vero Roboam prima et novissima scripta sunt in verbis Semeiae prophetae et Addo videntis, genealogia quoque et bella, quae erant inter Roboam et Ieroboam cunctis diebus.
2CHR|12|16|Et dormivit Roboam cum patribus suis sepultusque est in civitate David; et regnavit Abia filius eius pro eo.
2CHR|13|1|Anno octavo decimo regis Ieroboam regnavit Abia su per Iudam.
2CHR|13|2|Tribus annis regnavit in Ierusalem. Nomenque matris eius Michaia filia Uriel de Gabaa.Et erat bellum inter Abiam et Ieroboam.
2CHR|13|3|Cumque inisset Abia certamen et haberet bellicosissimos viros electorum quadringenta milia, Ieroboam instruxit e contra aciem octingenta milia virorum, qui et ipsi electi erant et ad bella fortissimi.
2CHR|13|4|Stetit igitur Abia super montem Semaraim, qui est in monte Ephraim, et ait: " Audi, Ieroboam et omnis Israel:
2CHR|13|5|Num ignoratis quod Dominus, Deus Israel, dederit regnum David super Israel in sempiternum, ipsi et filiis eius, pactum salis?
2CHR|13|6|Et surrexit Ieroboam filius Nabat servus Salomonis filii David et rebellavit contra dominum suum;
2CHR|13|7|congregatique sunt ad eum viri vanissimi, filii Belial, et praevaluerunt contra Roboam filium Salomonis. Porro Roboam erat iuvenis et corde pavido nec potuit resistere eis.
2CHR|13|8|Nunc ergo vos dicitis quod resistere possitis regno Domini, quod possidet per filios David, habetisque grandem populi multitudinem atque vitulos aureos, quos fecit vobis Ieroboam in deos.
2CHR|13|9|Et eiecistis sacerdotes Domini filios Aaron atque Levitas et fecistis vobis sacerdotes sicut populi terrarum. Quicumque venerit et initiaverit manum suam in tauro de bobus et in arietibus septem, fit sacerdos eorum, qui non sunt dii.
2CHR|13|10|Noster autem Deus Dominus est, quem non reliquimus; sacerdotesque ministrant Domino de filiis Aaron, et Levitae sunt in ordine suo.
2CHR|13|11|Holocausta quoque offerunt Domino per singulos dies, mane et vespere, et thymiama aromatum, et proponuntur panes in mensa mundissima. Estque apud nos candelabrum aureum et lucernae eius, ut accendantur semper ad vesperam; nos quippe custodimus praecepta Domini Dei nostri, quem vos reliquistis.
2CHR|13|12|Ergo in exercitu nostro dux Deus est et sacerdotes eius, qui clangunt tubis et resonant contra vos, filii Israel; nolite pugnare contra Dominum, Deum patrum vestrorum, quia non vobis expedit ".
2CHR|13|13|Ieroboam autem retro moliebatur insidias, ut venirent post eos, et erant ante Iudam, et insidiae post eos.
2CHR|13|14|Respiciensque Iuda vidit instare bellum ex adverso et post tergum et clamavit ad Dominum, ac sacerdotes tubis canere coeperunt,
2CHR|13|15|omnesque viri Iudae vociferati sunt; et ecce, illis clamantibus, perterruit Deus Ieroboam et omnem Israel coram Abia et Iuda.
2CHR|13|16|Fugeruntque filii Israel Iudam, et tradidit eos Deus in manu eorum.
2CHR|13|17|Percussit ergo eos Abia et populus eius plaga magna; et corruerunt vulnerati ex Israel quingenta milia virorum fortium.
2CHR|13|18|Humiliatique sunt filii Israel in tempore illo, et confortati filii Iudae, eo quod sperassent in Domino, Deo patrum suorum.
2CHR|13|19|Persecutus est autem Abia fugientem Ieroboam et cepit civitates eius Bethel et filias eius et Iesana cum filiabus suis, Ephron quoque et filias eius.
2CHR|13|20|Nec invaluit ultra Ieroboam in diebus Abiae. Quem percussit Dominus, et mortuus est.
2CHR|13|21|Abia autem confortatus est et accepit sibi uxores quattuordecim procreavitque viginti duos filios et sedecim filias.
2CHR|13|22|Reliqua autem gestorum Abiae viarumque et sermonum eius scripta sunt in enarratione prophetae Addo.
2CHR|13|23|Dormivit autem Abia cum patribus suis, et sepelierunt eum in civitate David; regnavitque Asa filius eius pro eo. In cuius diebus quievit terra annis decem.
2CHR|14|1|Fecit autem Asa, quod bo num et placitum erat in con spectu Domini Dei sui, et subvertit altaria peregrini cultus et excelsa
2CHR|14|2|et confregit lapides palosque succidit
2CHR|14|3|ac praecepit Iudae, ut quaereret Dominum, Deum patrum suorum, et faceret legem et universa mandata,
2CHR|14|4|et abstulit e cunctis urbibus Iudae excelsa et thymiateria et regnavit in pace.
2CHR|14|5|Aedificavit quoque urbes munitas in Iuda, quia quievit terra, et nulla temporibus eius bella surrexerant, pacem Domino ei largiente.
2CHR|14|6|Dixit autem Iudae: " Aedificemus civitates istas et vallemus muris et roboremus turribus et portis et seris, donec a bellis quieta sunt omnia; quia quaesivimus Dominum Deum nostrum, quaesivit nos et dedit nobis pacem per gyrum ". Aedificaverunt igitur et prosperati sunt.
2CHR|14|7|Habuit autem Asa exercitum portantium scuta et hastas de Iuda trecenta milia, de Beniamin vero scutariorum et sagittariorum ducenta octoginta milia; omnes isti viri fortissimi.
2CHR|14|8|Egressus est autem contra eos Zara Aethiops cum exercitu, decies centena milia et curribus trecentis, et venit usque Maresa.
2CHR|14|9|Porro Asa perrexit obviam ei, et instruxerunt aciem ad bellum in valle, quae est ad septentrionem Maresa,
2CHR|14|10|et invocavit Asa Dominum Deum suum et ait: " Domine, non est apud te ulla distantia, utrum paucis auxilieris an pluribus; adiuva nos, Domine Deus noster. In te enim et in tuo nomine habentes fiduciam venimus contra hanc multitudinem. Domine, Deus noster tu es, non praevaleat contra te homo ".
2CHR|14|11|Exterruit itaque Dominus Aethiopes coram Asa et Iuda; fugeruntque Aethiopes.
2CHR|14|12|Et persecutus est eos Asa et populus, qui cum eo erat, usque Gerar; et ruerunt Aethiopes usque ad internecionem, quia Domino caedente contriti sunt et exercitu illius proeliante. Tulerunt ergo spolia multa
2CHR|14|13|et percusserunt omnes civitates per circuitum Gerarae; terror quippe Domini eos invaserat. Et diripuerunt omnes urbes et multam praedam asportaverunt.
2CHR|14|14|Sed et caulas ovium destruentes tulerunt pecorum infinitam multitudinem et camelorum reversique sunt Ierusalem.
2CHR|15|1|Azarias autem filius Oded, facto in se spiritu Dei,
2CHR|15|2|egressus est in occursum Asa et dixit ei: " Audite me, Asa et omnis Iuda et Beniamin! Dominus vobiscum, quia fuistis cum eo. Si quaesieritis eum, invenietur a vobis; si autem dereliqueritis eum, derelinquet vos.
2CHR|15|3|Transierunt autem multi dies in Israel absque Deo veritatis et absque sacerdote doctore et absque lege.
2CHR|15|4|Cumque reversi essent in angustia sua ad Dominum, Deum Israel, et quaesivissent eum, inventus est ab eis.
2CHR|15|5|In temporibus illis non erat pax egredienti et ingredienti sed perturbatio magna multa in cunctis habitatoribus terrarum;
2CHR|15|6|contundebatur enim gens contra gentem, et civitas contra civitatem, quia Dominus conturbabat eos in omni angustia.
2CHR|15|7|Vos autem confortamini, et non dissolvantur manus vestrae; erit enim merces operi vestro ".
2CHR|15|8|Cum audisset Asa verba haec et prophetiam, confortatus est et abstulit idola de omni terra Iudae et Beniamin et ex urbibus, quas ceperat montis Ephraim, et dedicavit altare Domini, quod erat ante porticum Domini.
2CHR|15|9|Congregavitque universum Iudam et Beniamin et advenas cum eis de Ephraim et de Manasse et de Simeon; plures enim ad eum confugerant ex Israel videntes quod Dominus Deus illius esset cum eo.
2CHR|15|10|Cumque convenissent in Ierusalem mense tertio anno quinto decimo regni Asa,
2CHR|15|11|immolaverunt Domino in die illa de manubiis, quas adduxerant: boves septingentos et oves septem milia.
2CHR|15|12|Et inierunt foedus, ut quaererent Dominum, Deum patrum suorum, in toto corde et in tota anima sua:
2CHR|15|13|si quis autem non quaesierit Dominum, Deum Israel, moriatur a minimo usque ad maximum, a viro usque ad mulierem.
2CHR|15|14|Iuraveruntque Domino voce magna in iubilo et in clangore tubarum et in sonitu bucinarum.
2CHR|15|15|Omnes, qui erant in Iuda, gavisi sunt de iuramento; in omni enim corde suo iuraverant et in tota voluntate quaesierant eum, et inventus fuerat ab eis. Praestititque eis Dominus requiem per circuitum.
2CHR|15|16|Sed et Maacham matrem Asa rex amovit, ne esset domina, eo quod fecisset simulacrum Aserae; quod contrivit Asa et in frusta comminuens combussit in torrente Cedron.
2CHR|15|17|Excelsa autem derelicta sunt in Israel; attamen cor Asa erat perfectum cunctis diebus eius.
2CHR|15|18|Ea quae voverat pater suus et ipse, intulit in domum Dei, argentum et aurum vasorumque diversam supellectilem.
2CHR|15|19|Bellum vero non fuit usque ad tricesimum quintum annum regni Asa.
2CHR|16|1|Anno autem tricesimo sexto regni eius ascendit Baasa rex Israel in Iudam; et muro circumdabat Rama, ut nullus tute posset egredi et ingredi de regno Asa.
2CHR|16|2|Protulit ergo Asa argentum et aurum de thesauris domus Domini et domus regis misitque ad Benadad regem Syriae, qui habitabat in Damasco, dicens:
2CHR|16|3|" Foedus inter me et te est et inter patrem meum et patrem tuum; quam ob rem misi tibi argentum et aurum, ut, rupto foedere, quod habes cum Baasa rege Israel, facias eum a me recedere ".
2CHR|16|4|Acquiescens Benadad regi Asa misit principes exercituum suorum ad urbes Israel, qui percusserunt Ahion et Dan et Abelmaim et universa horrea urbium Nephthali.
2CHR|16|5|Quod cum audisset Baasa, desivit aedificare Rama et intermisit opus suum.
2CHR|16|6|Porro Asa rex assumpsit universum Iudam, et tulerunt lapides Rama et ligna, quibus aedificaverat Baasa, aedificavitque ex eis Gabaa et Maspha.
2CHR|16|7|In tempore illo venit Hanani videns ad Asa regem Iudae et dixit ei: " Quia habuisti fiduciam in rege Syriae et non in Domino Deo tuo, idcirco evasit Syriae regis exercitus de manu tua.
2CHR|16|8|Nonne Aethiopes et Libyes magnus exercitus erant quadrigis et equitibus et multitudine nimia, quos, cum Domino credidisses, tradidit in manu tua?
2CHR|16|9|Oculi enim Domini contemplantur universam terram et praebent fortitudinem his, qui corde perfecto credunt in eum. Stulte igitur egisti in hoc, quia ex praesenti tempore contra te bella consurgent ".
2CHR|16|10|Iratusque Asa adversus videntem iussit eum mitti in nervum, valde quippe super hoc fuerat indignatus; et vexavit Asa quosdam de populo in tempore illo.
2CHR|16|11|Opera autem Asa prima et novissima scripta sunt in libro regum Iudae et Israel.
2CHR|16|12|Aegrotavit etiam Asa anno tricesimo nono regni sui dolore pedum vehementissimo et nec in infirmitate sua quaesivit Dominum, sed magis in medicorum arte confisus est.
2CHR|16|13|Dormivitque Asa cum patribus suis et mortuus est anno quadragesimo primo regni sui.
2CHR|16|14|Et sepelierunt eum in sepulcro suo, quod foderat sibi in civitate David; posueruntque eum super lectum plenum aromatibus et variis unguentis, quae erant pigmentariorum arte confecta, et fecerunt in exsequiis eius combustionem splendidam valde.
2CHR|17|1|Regnavit autem Iosaphat filius eius pro eo et invaluit contra Israel.
2CHR|17|2|Constituitque militum numeros in cunctis urbibus Iudae, quae erant vallatae muris; praesidiaque disposuit in terra Iudae et in civitatibus Ephraim, quas ceperat Asa pater eius.
2CHR|17|3|Et fuit Dominus cum Iosaphat, quia ambulavit in viis patris sui primis et non speravit in Baalim
2CHR|17|4|sed in Deo patris sui et perrexit in praeceptis illius et non iuxta peccata Israel.
2CHR|17|5|Confirmavitque Dominus regnum in manu eius, et dedit omnis Iuda munera Iosaphat; factaeque sunt ei infinitae divitiae et multa gloria.
2CHR|17|6|Cumque sumpsisset cor eius audaciam propter vias Domini, etiam excelsa et palos de Iuda abstulit.
2CHR|17|7|Tertio autem anno regni sui misit principes suos Benhail et Abdiam et Zachariam et Nathanael et Michaiam, ut docerent in civitatibus Iudae,
2CHR|17|8|et cum eis Levitas Semeiam et Nathaniam et Zabadiam, Asael quoque et Semiramoth et Ionathan Adoniamque et Thobiam Levitas et cum eis Elisama et Ioram sacerdotes.
2CHR|17|9|Docebantque in Iuda habentes librum legis Domini et circuibant cunctas urbes Iudae atque erudiebant populum.
2CHR|17|10|Itaque factus est pavor Domini super omnia regna terrarum, quae erant per gyrum Iudae, nec audebant bellare contra Iosaphat.
2CHR|17|11|Sed et de Philisthim Iosaphat munera deferebant et vectigal argenti; Arabes quoque adducebant pecora arietum septem milia septingenta et hircos totidem.
2CHR|17|12|Crevit ergo Iosaphat et magnificatus est usque in sublime atque aedificavit in Iuda castella urbesque horreorum.
2CHR|17|13|Et multae copiae praesto erant ei in urbibus Iudae; viri quoque bellatores et robusti erant in Ierusalem,
2CHR|17|14|quorum iste numerus per familias singulorum: in Iuda principes exercitus, Ednas dux, et cum eo robustissimorum trecenta milia;
2CHR|17|15|et ad latus eius Iohanan princeps et cum eo ducenta octoginta milia;
2CHR|17|16|ad latus quoque istius Amasias filius Zechri consecratus Domino et cum eo ducenta milia virorum fortium;
2CHR|17|17|de Beniamin autem robustus ad proelia Eliada et cum eo tenentium arcum et clipeum ducenta milia;
2CHR|17|18|et ad latus eius Iozabad et cum eo centum octoginta milia expeditorum militum.
2CHR|17|19|Hi omnes erant ad manum regis, exceptis aliis, quos posuerat in urbibus muratis in universo Iuda.
2CHR|18|1|Fuit ergo Iosaphat dives et inclitus multum et affinitate coniunctus est Achab.
2CHR|18|2|Descenditque post annos ad eum in Samariam, ad cuius adventum mactavit Achab oves et boves plurimos ipsi et populo, qui venerat cum eo; persuasitque illi, ut ascenderet in Ramoth Galaad.
2CHR|18|3|Dixitque Achab rex Israel ad Iosaphat regem Iudae: " Veni mecum in Ramoth Galaad ". Cui ille respondit: " Ut ego, et tu; sicut populus tuus, sic et populus meus, tecumque erimus in bello ".
2CHR|18|4|Dixitque Iosaphat ad regem Israel: " Consule, obsecro, impraesentiarum sermonem Domini ".
2CHR|18|5|Congregavitque rex Israel prophetarum quadringentos viros et dixit ad eos: " In Ramoth Galaad ad bellandum ire debemus an quiescere? ". At illi: Ascende, inquiunt, et tradet Deus in manu regis ".
2CHR|18|6|Dixitque Iosaphat: " Numquid non est hic et alius propheta Domini, ut ab illo etiam requiramus? ".
2CHR|18|7|Et ait rex Israel ad Iosaphat: " Adhuc est vir unus, a quo possumus quaerere Domini voluntatem; sed ego odi eum, quia non prophetat mihi bonum sed malum omni tempore: est autem Michaeas filius Iemla ". Dixitque Iosaphat: " Ne loquaris, rex, hoc modo ".
2CHR|18|8|Vocavit ergo rex Israel unum de eunuchis et dixit ei: " Voca cito Michaeam filium Iemla ".
2CHR|18|9|Porro rex Israel et Iosaphat rex Iudae uterque sedebant in solio suo vestiti cultu regio; sedebant autem in area iuxta portam Samariae, omnesque prophetae vaticinabantur coram eis.
2CHR|18|10|Sedecias vero filius Chanaana fecit sibi cornua ferrea et ait: " Haec dicit Dominus: His ventilabis Syriam, donec conteras eam ".
2CHR|18|11|Omnesque prophetae similiter prophetabant atque dicebant: " Ascende in Ramoth Galaad et prosperaberis; et tradet Dominus in manu regis ".
2CHR|18|12|Nuntius autem, qui ierat ad vocandum Michaeam, ait illi: " En verba omnium prophetarum uno ore bona regi annuntiant; quaeso ergo te, ut et sermo tuus ab eis non dissentiat, loquarisque prospera ".
2CHR|18|13|Cui respondit Michaeas: " Vivit Dominus, quia, quodcumque dixerit Deus meus, hoc loquar! ".
2CHR|18|14|Venit ergo ad regem. Cui rex ait: " Michaea, ire debemus in Ramoth Galaad ad bellandum an quiescere? ". Cui ille respondit: " Ascendite et prosperamini, ut tradantur hostes in manus vestras ".
2CHR|18|15|Dixitque rex: " Iterum atque iterum te adiuro, ut non mihi loquaris nisi, quod verum est, in nomine Domini ".
2CHR|18|16|At ille ait: Vidi universum Israeldispersum in montibussicut oves absque pastore.Et dixit Dominus:Non habent isti dominum; revertatur unusquisque in domum suam in pace" ".
2CHR|18|17|Et ait rex Israel ad Iosaphat: " Nonne dixi tibi quod non prophetaret iste mihi quidquam boni sed ea, quae mala sunt? ".
2CHR|18|18|At ille idcirco ait: " Audite verbum Domini: Vidi Dominum sedentem in solio suo et omnem exercitum caeli assistentem ei a dextris et sinistris.
2CHR|18|19|Et dixit Dominus: "Quis decipiet Achab regem Israel, ut ascendat et corruat in Ramoth Galaad?". Cumque diceret unus hoc modo et alter alio,
2CHR|18|20|processit spiritus et stetit coram Domino et ait: "Ego decipiam eum". Cui Dominus: "In quo, inquit, decipies?".
2CHR|18|21|At ille respondit: "Egrediar et ero spiritus mendax in ore omnium prophetarum eius". Dixitque Dominus: "Decipies et praevalebis; egredere et fac ita".
2CHR|18|22|Nunc igitur, ecce dedit Dominus spiritum mendacii in ore omnium prophetarum tuorum et Dominus locutus est de te mala ".
2CHR|18|23|Accessit autem Sedecias filius Chanaana et percussit Michaeae maxillam et ait: " Per quam viam transivit spiritus Domini a me, ut loqueretur tibi? ".
2CHR|18|24|Dixitque Michaeas: " Tu ipse videbis in die illo, quando ingressus fueris cubiculum intra cubiculum, ut abscondaris ".
2CHR|18|25|Praecepit autem rex Israel dicens: " Tollite Michaeam et ducite eum ad Amon principem civitatis et ad Ioas filium regis
2CHR|18|26|et dicetis: "Haec dicit rex: Mittite hunc in carcerem et date ei panis modicum et aquae pauxillum, donec revertar in pace" ".
2CHR|18|27|Dixitque Michaeas: " Si reversus fueris in pace, non est locutus Dominus in me ". Et ait: " Audite, populi omnes! ".
2CHR|18|28|Igitur ascenderunt rex Israel et Iosaphat rex Iudae in Ramoth Galaad.
2CHR|18|29|Dixitque rex Israel ad Iosaphat: " Mutabo habitum et sic ad pugnam vadam; tu autem induere vestibus tuis ". Mutatoque rex Israel habitu venit ad bellum.
2CHR|18|30|Rex autem Syriae praeceperat ducibus curruum suorum dicens: " Ne pugnetis contra minimum aut contra maximum, nisi contra solum regem Israel.
2CHR|18|31|Itaque, cum vidissent principes curruum Iosaphat, dixerunt: " Rex Israel est iste! ". Et circumdederunt eum dimicantes. At ille clamavit ad Dominum, et auxiliatus est ei atque avertit eos Deus ab illo.
2CHR|18|32|Cum enim vidissent duces curruum quod non esset rex Israel, reliquerunt eum.
2CHR|18|33|Accidit autem, ut unus e populo sagittam in incertum iaceret et percuteret regem Israel inter iuncturas et loricam. At ille aurigae suo ait: " Converte manum tuam et educ me de acie, quia vulneratus sum ".
2CHR|18|34|Et aggravata est pugna in die illo; porro rex Israel stabat in curru suo contra Syros usque ad vesperam et mortuus est occidente sole.
2CHR|19|1|Reversus est autem Iosaphat rex Iudae in domum suam pacifice in Ierusalem.
2CHR|19|2|Cui occurrit Iehu filius Hanani videns et ait ad eum: " Impio praebes auxilium et his, qui oderunt Dominum, amicitia iungeris, et idcirco iram quidem Domini merebaris;
2CHR|19|3|sed bona opera inventa sunt in te, eo quod abstuleris palos de terra et praeparaveris cor tuum, ut requireres Deum ".
2CHR|19|4|Habitavit ergo Iosaphat in Ierusalem. Rursumque egressus est ad populum de Bersabee usque ad montem Ephraim et revocavit eos ad Dominum, Deum patrum suorum.
2CHR|19|5|Constituitque iudices terrae in cunctis civitatibus Iudae munitis per singula loca.
2CHR|19|6|Et praecipiens iudicibus: " Videte, ait, quid faciatis. Non enim homini exercetis iudicium sed Domino, qui vobiscum est, quando iudicaveritis.
2CHR|19|7|Sit timor Domini, vobiscum et caute cuncta facite; non est enim apud Dominum Deum nostrum iniquitas nec personarum acceptio nec cupido munerum.
2CHR|19|8|In Ierusalem quoque constituit Iosaphat ex Levitis et sacerdotibus et principibus familiarum Israel pro iudicio Domini et pro causis habitatorum Ierusalem.
2CHR|19|9|Praecepitque eis dicens: " Sic agetis in timore Domini fideliter et corde perfecto.
2CHR|19|10|Omnem causam, quae venerit ad vos fratrum vestrorum, qui habitant in urbibus suis, ubicumque quaestio est de homicidio, de lege, de mandato, de praeceptis et de iustificationibus, commonete eos, ut non peccent in Dominum, et ne veniat ira super vos et super fratres vestros; sic ergo agetis et non peccabitis.
2CHR|19|11|Amarias autem sacerdos princeps super vos in omnibus, quae ad Deum pertinent, praesidebit; porro Zabadias filius Ismael, qui est dux in domo Iudae, super ea opera erit, quae ad regis officium pertinent; habetisque Levitas coram vobis ut scribas. Confortamini et agite diligenter, et sit Dominus cum bonis ".
2CHR|20|1|Post haec congregati sunt filii Moab et filii Ammon et cum eis de Meunitis ad Iosaphat, ut pugnarent contra eum.
2CHR|20|2|Veneruntque nuntii et indicaverunt Iosaphat dicentes: " Venit contra te multitudo magna de his locis, quae trans mare sunt, de Edom, et ecce consistunt in Asasonthamar, quae est Engaddi ".
2CHR|20|3|Iosaphat autem timore perterritus totum se contulit ad rogandum Dominum et praedicavit ieiunium universo Iudae.
2CHR|20|4|Congregatusque est Iuda ad precandum Dominum; sed et de omnibus urbibus suis venerunt ad obsecrandum eum.
2CHR|20|5|Cumque stetisset Iosaphat in medio coetu Iudae et Ierusalem in domo Domini ante atrium novum,
2CHR|20|6|ait: " Domine, Deus patrum nostrorum, tu es Deus in caelo et dominaris cunctis regnis gentium; in manu tua est fortitudo et potentia, nec quisquam tibi potest resistere.
2CHR|20|7|Nonne tu, Deus noster, expulisti habitatores terrae huius coram populo tuo Israel et dedisti eam semini Abraham amici tui in sempiternum?
2CHR|20|8|Habitaveruntque in ea et exstruxerunt in illa sanctuarium nomini tuo dicentes:
2CHR|20|9|"Si irruerint super nos mala, gladius iudicii, pestilentia et fames, stabimus coram domo hac in conspectu tuo, quia nomen tuum est in domo hac, et clamabimus ad te in tribulationibus nostris, et exaudies salvosque facies".
2CHR|20|10|Nunc igitur ecce filii Ammon et Moab et mons Seir, per quos non concessisti Israeli ut transirent, quando egrediebantur de Aegypto, sed declinaverunt ab eis et non interfecerunt illos,
2CHR|20|11|e contrario agunt et nituntur eicere nos de possessione tua, quam tradidisti nobis.
2CHR|20|12|Deus noster, ergo non iudicabis eos? In nobis quidem non tanta est fortitudo, ut possimus huic multitudini resistere, quae irruit super nos; sed, cum ignoremus quid agere debeamus, hoc solum habemus residui, ut oculos nostros dirigamus ad te ".
2CHR|20|13|Omnis vero Iuda stabat coram Domino cum parvulis et uxoribus et liberis suis.
2CHR|20|14|Erat autem Iahaziel filius Zachariae filii Banaiae filii Iehiel filii Matthaniae Levites de filiis Asaph, super quem factus est spiritus Domini in medio congregationis,
2CHR|20|15|et ait: " Attendite, omnis Iuda et qui habitatis Ierusalem et tu rex Iosaphat: Haec dicit Dominus vobis: Nolite timere nec paveatis hanc multitudinem magnam; non est enim vestra pugna sed Dei.
2CHR|20|16|Cras descendetis contra eos; ascensuri enim sunt per clivum nomine Sis, et invenietis illos in summitate torrentis, qui est contra solitudinem Ieruel.
2CHR|20|17|Non eritis vos, qui dimicabitis; sed tantummodo confidenter state et videbitis auxilium Domini super vos, o Iuda et Ierusalem. Nolite timere nec paveatis; cras egredimini contra eos, et Dominus erit vobiscum ".
2CHR|20|18|Iosaphat ergo inclinavit se super faciem suam in terra, et omnis Iuda et habitatores Ierusalem ceciderunt coram Domino et adoraverunt eum.
2CHR|20|19|Porro Levitae de filiis Caath, de filiis Core scilicet, surrexerunt et laudabant Dominum, Deum Israel, voce magna in excelsum.
2CHR|20|20|Cumque mane surrexissent, egressi sunt ad desertum Thecue; profectisque eis, stans Iosaphat in medio eorum dixit: " Audite me, Iuda et habitatores Ierusalem! Credite in Domino Deo vestro et permanebitis; credite prophetis eius, et cuncta evenient vobis prospera ".
2CHR|20|21|Habuitque consilium cum populo et statuit cantores Domini, ut laudarent eum in ornatu sancto et antecederent exercitum ac voce consona dicerent: " Confitemini Domino, quoniam in aeternum misericordia eius ".
2CHR|20|22|Cumque coepissent laudes canere, vertit Dominus insidias eorum contra filios Ammon et Moab et montem Seir, qui egressi fuerant, ut pugnarent contra Iudam, et percussi sunt.
2CHR|20|23|Et filii Ammon et Moab consurrexerunt adversum habitatores montis Seir, ut interficerent et delerent eos; cumque hoc opere perpetrassent, etiam in semetipsos versi mutuis concidere vulneribus.
2CHR|20|24|Porro Iuda, cum venisset ad speculam, quae respicit solitudinem, vidit procul omnem late regionem plenam cadaveribus, nec superesse quemquam, qui necem potuisset evadere.
2CHR|20|25|Venit ergo Iosaphat et omnis populus cum eo ad detrahenda spolia mortuorum inveneruntque iumenta multa et supellectilem, vestes quoque et vasa pretiosissima et diripuerunt, ita ut omnia portare non possent, et per tres dies spolia auferebant pro praedae magnitudine.
2CHR|20|26|Die autem quarto congregati sunt in valle Baracha; etenim, quoniam ibi benedixerant Domino, vocaverunt locum illum vallis Benedictionis usque in praesentem diem.
2CHR|20|27|Reversusque est omnis vir Iudae et Ierusalem et Iosaphat ante eos in Ierusalem cum laetitia magna, eo quod dedisset eis Dominus gaudium de inimicis suis;
2CHR|20|28|ingressique sunt Ierusalem cum psalteriis et citharis et tubis in domum Domini.
2CHR|20|29|Irruit autem pavor Dei super universa regna terrarum, cum audissent quod pugnasset Dominus contra inimicos Israel.
2CHR|20|30|Quievitque regnum Iosaphat, et praebuit ei Deus eius pacem per circuitum.
2CHR|20|31|Regnavit igitur Iosaphat super Iudam. Et erat triginta quinque annorum, cum regnare coepisset; viginti autem et quinque annis regnavit in Ierusalem. Nomen matris eius Azuba filia Selachi.
2CHR|20|32|Et ambulavit in via patris sui Asa nec declinavit ab ea, faciens quod rectum erat coram Domino.
2CHR|20|33|Verumtamen excelsa non ablata sunt; et adhuc populus non direxerat cor suum ad Deum patrum suorum.
2CHR|20|34|Reliqua autem gestorum Iosaphat, priorum et novissimorum, scripta sunt in verbis Iehu filii Hanani, quae digesta sunt in libros regum Israel.
2CHR|20|35|Post haec iniit amicitias Iosaphat rex Iudae cum Ochozia rege Israel, cuius opera fuerunt impiissima,
2CHR|20|36|et particeps fuit, ut facerent naves, quae irent in Tharsis, feceruntque classem in Asiongaber.
2CHR|20|37|Prophetavit autem Eliezer filius Dodiae de Maresa contra Iosaphat dicens: " Quia habuisti foedus cum Ochozia, percussit Dominus opera tua ". Contritaeque sunt naves nec potuerunt ire in Tharsis.
2CHR|21|1|Dormivit autem Iosaphat cum patribus suis et sepultus est cum eis in civitate David; regnavitque Ioram filius eius pro eo.
2CHR|21|2|Qui habuit fratres filios Iosaphat Azariam et Iahiel et Zachariam et Azariam et Michael et Saphatiam: omnes hi filii Iosaphat regis Israel.
2CHR|21|3|Deditque eis pater suus multa munera argenti et auri et res pretiosas cum civitatibus munitissimis in Iuda; regnum autem tradidit Ioram, eo quod esset primogenitus.
2CHR|21|4|Surrexit ergo Ioram super regnum patris sui; cumque se confirmasset, occidit omnes fratres suos gladio et quosdam de principibus Israel.
2CHR|21|5|Triginta duorum annorum erat Ioram, cum regnare coepisset, et octo annis regnavit in Ierusalem.
2CHR|21|6|Ambulavitque in viis regum Israel, sicut egerat domus Achab; filia quippe Achab erat uxor eius. Et fecit malum in conspectu Domini.
2CHR|21|7|Noluit autem Dominus disperdere domum David propter pactum, quod inierat cum eo, et quia promiserat, ut daret ei lucernam et filiis eius omni tempore.
2CHR|21|8|In diebus illis rebellavit Edom, ne esset subditus Iudae, et constituit sibi regem.
2CHR|21|9|Cumque transisset Ioram cum principibus suis et cunctis curribus, qui erant secum, surrexit nocte et percussit Edom, qui eum circumdederat, et omnes duces curruum eius.
2CHR|21|10|Attamen rebellavit Edom, ne esset sub dicione Iudae, usque ad hanc diem. Eo tempore et Lobna recessit, ne esset sub manu illius; dereliquerat enim Dominum, Deum patrum suorum.
2CHR|21|11|Insuper et excelsa fabricatus est in montibus Iudae et fornicari fecit habitatores Ierusalem et praevaricari Iudam.
2CHR|21|12|Allatae sunt autem ei litterae ab Elia propheta, in quibus scriptum erat: "Haec dicit Dominus, Deus David patris tui: Quoniam non ambulasti in viis Iosaphat patris tui et in viis Asa regis Iudae,
2CHR|21|13|sed incessisti per iter regum Israel et fornicari fecisti Iudam et habitatores Ierusalem imitatus fornicationem domus Achab, insuper et fratres tuos domum patris tui meliores te occidisti:
2CHR|21|14|ecce Dominus percutiet plaga magna populum tuum, filios et uxores tuas universamque substantiam tuam;
2CHR|21|15|tu autem aegrotabis pessimo languore uteri tui, donec egrediantur vitalia tua paulatim per singulos dies ".
2CHR|21|16|Suscitavit ergo Dominus contra Ioram spiritum Philisthinorum et Arabum, qui confines sunt Aethiopibus,
2CHR|21|17|et ascenderunt in terram Iudae et irruperunt in eam diripueruntque cunctam substantiam, quae inventa est in domo regis, insuper et filios eius et uxores, nec remansit ei filius nisi Ioachaz, qui minimus natu erat.
2CHR|21|18|Et post haec omnia percussit eum Dominus alvi languore insanabili.
2CHR|21|19|Cumque diei succederet dies, et temporum spatia volverentur, duorum annorum expletus est circulus; et sic longa consumptus tabe, ita ut egereret etiam viscera sua, languore pariter et vita caruit. Mortuusque est in infirmitate pessima, et non fecit ei populus eius secundum morem combustionis exsequias, sicut fecerat maioribus eius.
2CHR|21|20|Triginta duorum annorum fuit, cum regnare coepisset, et octo annis regnavit in Ierusalem. Obiitque nullo relicto desiderio sui; et sepelierunt eum in civitate David, verumtamen non in sepulcro regum.
2CHR|22|1|Constituerunt autem habita tores Ierusalem Ochoziam fi lium eius minimum regem pro eo; omnes enim maiores natu interfecerat turba, quae irruerat cum Arabibus in castra. Regnavitque Ochozias filius Ioram regis Iudae.
2CHR|22|2|Filius viginti duo annorum erat Ochozias, cum regnare coepisset, et uno anno regnavit in Ierusalem. Nomen matris eius Athalia filia Amri.
2CHR|22|3|Sed et ipse ingressus est per vias domus Achab; mater enim eius impulit eum, ut impie ageret.
2CHR|22|4|Fecit igitur malum in conspectu Domini sicut domus Achab; ipsi enim fuerunt ei consiliarii post mortem patris sui in interitum eius.
2CHR|22|5|Ambulavitque in consiliis eorum et perrexit cum Ioram filio Achab rege Israel in bellum contra Hazael regem Syriae in Ramoth Galaad; vulneraveruntque Syri Ioram.
2CHR|22|6|Qui reversus est, ut curaretur in Iezrahel a plagis, quas acceperat in supradicto certamine.Igitur Ochozias filius Ioram rex Iudae descendit, ut inviseret Ioram filium Achab in Iezrahel aegrotantem.
2CHR|22|7|Voluntatis quippe fuit Dei adversum Ochoziam, ut veniret ad Ioram et, cum venisset, egrederetur cum eo adversum Iehu filium Namsi, quem unxit Dominus, ut deleret domum Achab.
2CHR|22|8|Cum ergo iudicium faceret Iehu in domum Achab, invenit principes Iudae et filios fratrum Ochoziae, qui ministrabant ei, et interfecit illos.
2CHR|22|9|Ipsumque perquisivit Ochoziam, et comprehenderunt eum latentem in Samaria; adductumque ad se Iehu occidit. Et sepelierunt eum, eo quod dicebant eum esse filium Iosaphat, qui quaesierat Dominum in toto corde suo.Nec erat aliquis de stirpe Ochoziae, qui posset regnare.
2CHR|22|10|Athalia autem mater eius videns quod mortuus esset filius suus surrexit et interfecit omnem stirpem regiam domus Iudae.
2CHR|22|11|Porro Iosabeth filia regis tulit Ioas filium Ochoziae et furata est eum de medio filiorum regis, cum interficerentur, absconditque cum nutrice sua in cubiculo lectulorum. Iosabeth autem, quae absconderat eum, erat filia regis Ioram, uxor Ioiadae pontificis, soror Ochoziae; et idcirco Athalia non interfecit eum.
2CHR|22|12|Fuit ergo cum eis in domo Dei absconditus sex annis, quibus regnavit Athalia super terram.
2CHR|23|1|Anno autem septimo confor tatus Ioiada assumpsit centu riones, Azariam videlicet filium Ieroham et Ismael filium Iohanan, Azariam quoque filium Obed et Maasiam filium Adaiae et Elisaphat filium Zechri, et iniit cum eis foedus.
2CHR|23|2|Qui circumeuntes Iudam congregaverunt Levitas de cunctis urbibus Iudae et principes familiarum Israel veneruntque in Ierusalem.
2CHR|23|3|Iniit igitur omnis congregatio pactum in domo Dei cum rege. Dixitque ad eos Ioiada: " Ecce filius regis regnabit, sicut locutus est Dominus super filios David.
2CHR|23|4|Hoc est ergo, quod facietis.
2CHR|23|5|Tertia pars vestrum, qui veniunt ad sabbatum sacerdotum et Levitarum et ianitorum, erit in portis, tertia vero pars ad domum regis et tertia in porta, quae appellatur Fundamenti; omne vero reliquum vulgus sit in atriis domus Domini.
2CHR|23|6|Nec quisquam alius ingrediatur domum Domini, nisi sacerdotes et qui ministrant de Levitis; ipsi tantummodo ingrediantur, quia sanctificati sunt. Et omne reliquum vulgus observet observationem Domini.
2CHR|23|7|Levitae autem circumdent regem habentes singuli arma sua in manu. Et si quis alius ingressus fuerit templum, interficiatur. Sintque cum rege et intrante et egrediente ".
2CHR|23|8|Fecerunt igitur Levitae et universus Iuda iuxta omnia, quae praeceperat Ioiada pontifex; et assumpserunt singuli viros suos, qui veniebant sabbato cum his, qui sabbato egressuri erant: siquidem Ioiada pontifex non dimisit abire turmas, quae sibi per singulas hebdomadas succedere consueverant.
2CHR|23|9|Deditque Ioiada sacerdos centurionibus lanceas clipeosque et peltas regis David, quae erant in domo Dei.
2CHR|23|10|Constituitque omnem populum tenentium tela a parte templi dextra usque ad partem templi sinistram coram altari et templo per circuitum regis.
2CHR|23|11|Et eduxerunt filium regis et dederunt ei diadema et testimonium et constituerunt eum regem. Unxerunt quoque illum Ioiada pontifex et filii eius; imprecatique sunt ei atque dixerunt: " Vivat rex! ".
2CHR|23|12|Quod cum audisset Athalia, vocem scilicet currentium atque laudantium regem, ingressa est ad populum in templum Domini.
2CHR|23|13|Cumque vidisset regem stantem super gradum suum in introitu et principes tubasque circa eum omnemque populum terrae gaudentem atque clangentem tubis cantoresque cum diversi generis organis signum dantes ad laudandum, scidit vestimenta sua et ait: " Coniuratio, coniuratio! ".
2CHR|23|14|Praecepit autem Ioiada pontifex centurionibus, qui erant super exercitum, dicens: " Educite illam extra saepta templi! Qui autem sequetur eam, interficiatur foris gladio! ". Dixerat enim sacerdos: " Non occidetis eam in domo Domini! ".
2CHR|23|15|Et imposuerunt ei manus; cumque intrasset portam Equorum domus regis, interfecerunt eam ibi.
2CHR|23|16|Pepigit autem Ioiada foedus inter se universumque populum et regem, ut esset populus Domini.
2CHR|23|17|Itaque ingressus est omnis populus domum Baal et destruxerunt eam et altaria ac simulacra illius confregerunt; Matthan quoque sacerdotem Baal interfecerunt ante aras.
2CHR|23|18|Constituit autem Ioiada praepositos in domo Domini sub manibus sacerdotum et Levitarum, quos distribuit David in domo Domini, ut offerrent holocausta Domino, sicut scriptum est in lege Moysi, in gaudio et canticis iuxta dispositionem David.
2CHR|23|19|Constituit quoque ianitores in portis domus Domini, ut non ingrederetur eam immundus in omni re.
2CHR|23|20|Assumpsitque centuriones et fortissimos viros ac principes populi et omne vulgus terrae, et fecerunt descendere regem de domo Domini et introire per medium portae Superioris in domum regis et collocaverunt eum in solio regali.
2CHR|23|21|Laetatusque est omnis populus terrae, et urbs quievit; porro Athalia interfecta est gladio.
2CHR|24|1|Septem annorum erat Ioas, cum regnare coepisset, et quadraginta annis regnavit in Ierusalem. Nomen matris eius Sebia de Bersabee.
2CHR|24|2|Fecitque, quod bonum est coram Domino, cunctis diebus Ioiadae sacerdotis.
2CHR|24|3|Accepit autem ei Ioiada uxores duas, e quibus genuit filios et filias.
2CHR|24|4|Post quae placuit Ioas, ut instauraret domum Domini.
2CHR|24|5|Congregavitque sacerdotes et Levitas et dixit eis: " Egredimini ad civitates Iudae et colligite de universo Israel pecuniam ad sartatecta templi Dei vestri per singulos annos. Festinatoque hoc facite ". Porro Levitae non festinarunt.
2CHR|24|6|Vocavitque rex Ioiadam principem et dixit ei: " Quare non tibi fuit curae, ut cogeres Levitas inferre de Iuda et de Ierusalem pecuniam, quae constituta est a Moyse servo Domini, ut inferret eam omnis congregatio Israel in tabernaculum testimonii?
2CHR|24|7|Athalia enim impiissima et filii eius dissipaverunt domum Dei et de universis, quae sanctificata fuerant templo Domini, dedicaverunt Baalim ".
2CHR|24|8|Praecepit ergo rex, et fecerunt arcam posueruntque eam iuxta portam domus Domini forinsecus.
2CHR|24|9|Et praedicatum est in Iuda et Ierusalem, ut deferrent singuli pretium Domino, quod constituit Moyses servus Dei super Israel in deserto.
2CHR|24|10|Laetatique sunt cuncti principes et omnis populus et ingressi contulerunt in arcam atque miserunt ita, ut impleretur.
2CHR|24|11|Cumque tempus esset, ut deferrent arcam ad magistratus regis per manus Levitarum, et viderent multam esse pecuniam, ingrediebatur scriba regis et quem primus sacerdos constituerat, effundebantque pecuniam, quae erat in arca; porro arcam reportabant ad locum suum. Sicque faciebant per singula tempora, et congregata est infinita pecunia,
2CHR|24|12|quam dederunt rex et Ioiada his, qui praeerant operibus domus Domini. At illi conducebant ex ea caesores lapidum et artifices operum singulorum, ut instaurarent domum Domini, fabros quoque ferri et aeris, ut domus Dei fulciretur.
2CHR|24|13|Egeruntque operarii, et obducebatur cicatrix operi per manus eorum, ac suscitaverunt domum Domini in statum pristinum et firme eam stare fecerunt.
2CHR|24|14|Cumque haec complessent, detulerunt coram rege et Ioiada reliquam partem pecuniae, de qua facta sunt vasa templi in ministerium et ad holocausta, phialae quoque et cetera vasa aurea et argentea. Et offerebantur holocausta in domo Domini iugiter cunctis diebus Ioiadae.
2CHR|24|15|Senuit autem Ioiada plenus dierum et mortuus est cum centum triginta esset annorum.
2CHR|24|16|Sepelieruntque eum in civitate David cum regibus, eo quod fecisset bonum in Israel cum Deo et cum domo eius.
2CHR|24|17|Postquam autem obiit Ioiada, ingressi sunt principes Iudae et adoraverunt regem, qui delinitus obsequiis eorum acquievit eis.
2CHR|24|18|Et dereliquerunt templum Domini, Dei patrum suorum, servieruntque palis et sculptilibus, et facta est ira contra Iudam et Ierusalem propter hoc peccatum.
2CHR|24|19|Mittebatque eis prophetas, ut reverterentur ad Dominum, quos protestantes illi audire nolebant.
2CHR|24|20|Spiritus itaque Dei induit Zachariam filium Ioiadae sacerdotis; et stetit in conspectu populi et dixit eis: " Haec dicit Deus: Quare transgredimini praecepta Domini, quod vobis non proderit? Quia dereliquistis Dominum, ipse dereliquit vos ".
2CHR|24|21|Qui coniuraverunt adversus eum et lapidaverunt eum iuxta regis imperium in atrio domus Domini.
2CHR|24|22|Et non est recordatus Ioas rex misericordiae, quam fecerat Ioiada pater illius secum, sed interfecit filium eius. Qui cum moreretur, ait: " Videat Dominus et requirat! ".
2CHR|24|23|Cumque evolutus esset annus, ascendit contra eum exercitus Syriae venitque in Iudam et Ierusalem et exterminaverunt cunctos principes populi atque universam praedam miserunt regi Damascum.
2CHR|24|24|Et certe, cum permodicus venisset numerus Syrorum, tradidit Dominus manibus eorum exercitum magnum valde, eo quod reliquissent Dominum, Deum patrum suorum; in Ioas quoque ignominiosa exercuere iudicia.
2CHR|24|25|Et abeuntes dimiserunt eum in languoribus magnis. Coniuraverunt autem contra eum servi sui in ultionem sanguinis filii Ioiadae sacerdotis et occiderunt eum in lectulo suo, et mortuus est. Sepelieruntque eum in civitate David, sed non in sepulcris regum.
2CHR|24|26|Insidiati vero sunt ei Zabad filius Semath Ammanitidis et Iozabad filius Semarith Moabitidis.
2CHR|24|27|Porro de filiis eius, de summa tributi, quod impositum fuerat sub eo, et de instauratione domus Dei scriptum est in commentariis libri regum. Regnavitque Amasias filius eius pro eo.
2CHR|25|1|Viginti quinque annorum erat Amasias, cum regnare coepisset, et viginti novem annis regnavit in Ierusalem. Nomen matris eius Ioaden de Ierusalem.
2CHR|25|2|Fecitque bonum in conspectu Domini, verumtamen non in corde perfecto.
2CHR|25|3|Cumque roboratum sibi videret imperium, iugulavit servos suos, qui occiderant regem patrem suum,
2CHR|25|4|sed filios eorum non interfecit, sicut scriptum est in libro legis Moysi, ubi praecepit Dominus dicens: " Non occidentur patres pro filiis, neque filii pro patribus suis, sed unusquisque in suo peccato morietur ".
2CHR|25|5|Congregavit igitur Amasias Iudam et constituit eos per familias tribunosque et centuriones in universo Iuda et Beniamin. Et recensuit a viginti annis sursum invenitque trecenta milia iuvenum, qui egrederentur ad pugnam et tenerent hastam et clipeum.
2CHR|25|6|Mercede quoque conduxit de Israel centum milia robustorum centum talentis argenti.
2CHR|25|7|Venit autem homo Dei ad illum et ait: " O rex, ne egrediatur tecum exercitus Israel; non est enim Dominus cum Israel, cunctis filiis Ephraim.
2CHR|25|8|Quod si putas in robore exercitus bella consistere, superari te faciet Deus ab hostibus: Dei quippe est et adiuvare et in fugam vertere ".
2CHR|25|9|Dixitque Amasias ad hominem Dei: " Quid ergo fiet de centum talentis, quae dedi militibus Israel? ". Et respondit ei homo Dei: " Habet Dominus, unde tibi dare possit multo his plura ".
2CHR|25|10|Separavit itaque Amasias exercitum, qui venerat ad eum ex Ephraim, ut reverteretur in locum suum; at illi contra Iudam vehementer irati reversi sunt in regionem suam.
2CHR|25|11|Porro Amasias confidenter eduxit populum suum et abiit in vallem Salinarum percussitque filios Seir decem milia.
2CHR|25|12|Et alia decem milia virorum ceperunt filii Iudae et adduxerunt ad praeruptum cuiusdam petrae praecipitaveruntque eos de summo in praeceps, qui universi crepuerunt.
2CHR|25|13|At ille exercitus, quem remiserat Amasias, ne secum iret ad proelium, diffusus est in civitatibus Iudae a Samaria usque Bethoron et, interfectis tribus milibus, diripuit praedam magnam.
2CHR|25|14|Amasias vero, post caedem Idumaeorum et allatos deos filiorum Seir, statuit illos in deos sibi et adorabat eos et illis adolebat.
2CHR|25|15|Quam ob rem iratus Dominus contra Amasiam misit ad illum prophetam, qui diceret ei: " Cur adorasti deos, qui non liberaverunt populum suum de manu tua? ".
2CHR|25|16|Cumque haec ille loqueretur, respondit ei: " Num consiliarium regis fecimus te? Quiesce! Cur interficiam te? ". Discedensque propheta: " Sed scio, inquit, quod decrevit Deus occidere te, quia fecisti hoc et non acquievisti consilio meo ".
2CHR|25|17|Igitur Amasias rex Iudae, inito consilio, misit ad Ioas filium Ioachaz filii Iehu regem Israel dicens: " Veni, videamus nos mutuo! ".
2CHR|25|18|At ille remisit nuntium dicens: " Carduus, qui est in Libano, misit ad cedrum Libani dicens: "Da filiam tuam filio meo uxorem". Et ecce bestiae agri, quae erant in Libano, transierunt et conculcaverunt carduum.
2CHR|25|19|Dixisti: "Percussi Edom!". Et idcirco erigitur cor tuum in superbiam. Sede in domo tua! Cur malum adversum te provocas, ut cadas et tu et Iuda tecum? ".
2CHR|25|20|Noluit audire Amasias, eo quod Domini esset voluntas, ut traderetur in manibus hostium propter cultum deorum Edom.
2CHR|25|21|Ascendit igitur Ioas rex Israel, et mutuos sibi praebuere conspectus: ipse et Amasias rex Iudae in Bethsames Iudae.
2CHR|25|22|Corruitque Iuda coram Israel et fugit in tabernacula sua.
2CHR|25|23|Porro Amasiam regem Iudae filium Ioas filii Ioachaz cepit Ioas rex Israel in Bethsames et adduxit in Ierusalem destruxitque murum eius a porta Ephraim usque ad portam Anguli quadringentis cubitis.
2CHR|25|24|Omne quoque aurum et argentum et universa vasa, quae repererat in domo Dei et apud Obededom in thesauris etiam domus regiae, necnon et obsides reduxit Samariam.
2CHR|25|25|Vixit autem Amasias filius Ioas rex Iudae, postquam mortuus est Ioas filius Ioachaz rex Israel, quindecim annis.
2CHR|25|26|Reliqua vero gestorum Amasiae priorum et novissimorum scripta sunt in libro regum Iudae et Israel.
2CHR|25|27|Qui postquam recessit a Domino, tetenderunt ei insidias in Ierusalem; cumque fugisset Lachis, miserunt post eum in Lachis et interfecerunt eum ibi.
2CHR|25|28|Reportantesque super equos sepelierunt eum cum patribus suis in civitate David.
2CHR|26|1|Omnis autem populus Iudae Oziam annorum sedecim constituit regem pro patre suo Amasia.
2CHR|26|2|Ipse reaedificavit Ailath et restituit eam dicioni Iudae, postquam dormivit rex cum patribus suis.
2CHR|26|3|Sedecim annorum erat Ozias, cum regnare coepisset, et quinquaginta duobus annis regnavit in Ierusalem. Nomen matris eius Iechelia de Ierusalem.
2CHR|26|4|Fecitque, quod erat rectum in oculis Domini iuxta omnia, quae fecerat Amasias pater eius.
2CHR|26|5|Et exquisivit Deum in diebus Zachariae, qui erudivit eum in timore Dei; et quamdiu requirebat Dominum, eum prosperari fecit Deus.
2CHR|26|6|Denique egressus est et pugnavit contra Philisthim et destruxit murum Geth et murum Iabniae murumque Azoti. Aedificavit quoque oppida in regione Azoti et Philisthim.
2CHR|26|7|Et adiuvit eum Deus contra Philisthim et contra Arabas, qui habitabant in Gurbaal, et contra Meunitas.
2CHR|26|8|Pendebantque Ammonitae munera Oziae; et divulgatum est nomen eius usque ad introitum Aegypti, quia confortatus est in excelsum.
2CHR|26|9|Aedificavitque Ozias turres in Ierusalem super portam Anguli et super portam Vallis et super Angulum firmavitque eas.
2CHR|26|10|Exstruxit etiam turres in solitudine et fodit cisternas plurimas, eo quod haberet multa pecora tam in Sephela quam in planitie; agricolas quoque habuit et vinitores in montibus et in campis fertilibus; erat quippe homo agriculturae deditus.
2CHR|26|11|Fuit autem exercitus bellatorum eius, qui procedebant ad proelia in turmis secundum numerum census per manum Iehiel scribae Maasiaeque praefecti sub manu Hananiae, qui erat de ducibus regis.
2CHR|26|12|Omnisque numerus principum per familias virorum fortium duorum milium sescentorum.
2CHR|26|13|Et sub eis universus exercitus trecentorum et septem milium quingentorum, qui erant apti ad bella, ut pro rege contra adversarios dimicarent.
2CHR|26|14|Praeparavit quoque eis Ozias, id est cuncto exercitui, clipeos et hastas et galeas et loricas arcusque et fundas ad iaciendos lapides.
2CHR|26|15|Et fecit in Ierusalem machinas excogitatas arte, quas in turribus collocavit et in angulis murorum, ut mitterent sagittas et saxa grandia; egressumque est nomen eius procul, eo quod mirabiliter auxiliaretur ei Dominus et corroborasset illum.
2CHR|26|16|Sed, cum roboratus esset, elevatum est cor eius in interitum suum, et deliquit contra Dominum Deum suum; ingressusque templum Domini adolere voluit incensum super altare thymiamatis.
2CHR|26|17|Statimque ingressus post eum Azarias sacerdos et cum eo sacerdotes Domini octoginta viri fortissimi;
2CHR|26|18|restiterunt regi atque dixerunt: " Non est tui officii, Ozia, ut adoleas incensum Domino, sed sacerdotum, hoc est filiorum Aaron, qui consecrati sunt ad huiuscemodi ministerium. Egredere de sanctuario, quia praevaricatus es; et non reputabitur tibi in gloriam hoc a Domino Deo ".
2CHR|26|19|Iratusque est Ozias et tenens in manu turibulum, ut adoleret incensum, minabatur sacerdotibus. Statimque orta est lepra in fronte eius coram sacerdotibus in domo Domini super altare thymiamatis.
2CHR|26|20|Cumque respexisset eum Azarias pontifex et omnes reliqui sacerdotes, viderunt lepram in fronte eius et festinato expulerunt eum; sed et ipse acceleravit egredi, eo quod malo afflixisset eum Dominus.
2CHR|26|21|Fuit igitur Ozias rex leprosus usque ad diem mortis suae et habitavit in domo separata plenus lepra, eo quod abscissus fuerat de domo Domini. Porro Ioatham filius eius rexit domum regis et iudicabat populum terrae.
2CHR|26|22|Reliqua autem gestorum Oziae priorum et novissimorum scripsit Isaias filius Amos propheta.
2CHR|26|23|Dormivitque Ozias cum patribus suis, et sepelierunt eum in agro regalium sepulcrorum, eo quod dicebant: " Erat leprosus ". Regnavitque Ioatham filius eius pro eo.
2CHR|27|1|Viginti quinque annorum erat Ioatham, cum regnare coepisset, et sedecim annis regnavit in Ierusalem. Nomen matris eius Ierusa filia Sadoc.
2CHR|27|2|Fecitque, quod rectum erat coram Domino iuxta omnia, quae fecerat Ozias pater suus, excepto quod non est ingressus templum Domini, et adhuc populus delinquebat.
2CHR|27|3|Ipse aedificavit portam domus Domini Superiorem et in muro Ophel multa construxit.
2CHR|27|4|Urbes quoque aedificavit in montibus Iudae et in saltibus castella et turres.
2CHR|27|5|Ipse pugnavit contra regem filiorum Ammon et vicit eos, dederuntque ei filii Ammon in anno illo centum talenta argenti et decem milia choros tritici ac totidem choros hordei; haec ei praebuerunt filii Ammon etiam in anno secundo et tertio.
2CHR|27|6|Corroboratusque est Ioatham, eo quod direxisset vias suas coram Domino Deo suo.
2CHR|27|7|Reliqua autem gestorum Ioatham et omnes pugnae eius et viae scriptae sunt in libro regum Israel et Iudae.
2CHR|27|8|Viginti quinque annorum erat, cum regnare coepisset, et sedecim annis regnavit in Ierusalem.
2CHR|27|9|Dormivitque Ioatham cum patribus suis, et sepelierunt eum in civitate David; et regnavit Achaz filius eius pro eo.
2CHR|28|1|Viginti annorum erat Achaz, cum regnare coepis set, et sedecim annis regnavit in Ierusalem. Non fecit rectum in conspectu Domini sicut David pater eius,
2CHR|28|2|sed ambulavit in viis regum Israel. Insuper et simulacra fudit Baalim.
2CHR|28|3|Ipse est, qui adolevit in valle filii Ennom et lustravit filios suos in igne iuxta abominationes gentium, quas expulit Dominus coram filiis Israel.
2CHR|28|4|Sacrificabat quoque et thymiama succendebat in excelsis et in collibus et sub omni ligno frondoso.
2CHR|28|5|Tradiditque eum Dominus Deus eius in manu regis Syriae, qui percussit eum multosque captivos de eo cepit et adduxit in Damascum. Manibus quoque regis Israel traditus est et percussus plaga grandi.
2CHR|28|6|Occidit enim Phacee filius Romeliae de Iuda centum viginti milia in die uno, omnes viros bellatores, eo quod reliquissent Dominum, Deum patrum suorum.
2CHR|28|7|Eodem tempore occidit Zechri vir potens ex Ephraim Maasiam filium regis et Ezricam praefectum domus, Elcanam quoque secundum a rege.
2CHR|28|8|Ceperuntque filii Israel de fratribus suis ducenta milia mulierum, puerorum et puellarum, et infinitam praedam pertuleruntque eam in Samariam.
2CHR|28|9|Erat autem ibi propheta Domini nomine Oded, qui egressus obviam exercitui venienti in Samariam dixit eis: " Ecce, iratus Dominus, Deus patrum vestrorum, contra Iudam tradidit eos in manibus vestris, et occidistis eos atrociter, ita ut ad caelum pertingeret vestra crudelitas.
2CHR|28|10|Insuper filios Iudae et Ierusalem vultis vobis subicere in servos et ancillas. Attamen nonne vos ipsi estis in culpa coram Domino Deo vestro?
2CHR|28|11|Audite ergo consilium meum et reducite captivos, quos adduxistis de fratribus vestris, quia magnus furor Domini imminet vobis ".
2CHR|28|12|Steterunt itaque viri de principibus filiorum Ephraim, Azarias filius Iohanan, Barachias filius Mosollamoth, Ezechias filius Sellum et Amasa filius Adali, contra eos, qui veniebant de proelio,
2CHR|28|13|et dixerunt eis: " Non introducetis huc captivos, quia ad culpam coram Domino, quae iam est super nos, vultis adicere super peccata nostra et culpam nostram. Grandis quippe culpa est nobis, et ira furoris Domini super Israel ".
2CHR|28|14|Dimiseruntque viri bellatores captivos et universa, quae ceperant, coram principibus et omni multitudine.
2CHR|28|15|Et surrexerunt viri nominatim designati et confortaverunt captivos omnesque, qui nudi erant, vestierunt de spoliis. Cumque vestissent eos et calceassent et refecissent cibo ac potu unxissentque, deduxerunt eos sollicite, et quidem omnes vacillantes in iumentis, et adduxerunt Iericho civitatem Palmarum ad fratres eorum. Ipsique reversi sunt Samariam.
2CHR|28|16|Tempore illo misit rex Achaz ad regem Assyriorum auxilium postulans.
2CHR|28|17|Venerunt enim et Idumaei et percusserunt Iudam et ceperunt captivos.
2CHR|28|18|Philisthim quoque diffusi sunt per urbes Sephelae et Nageb Iudae ceperuntque Bethsames et Aialon et Gederoth, Socho quoque cum viculis eius et Thamnan et Gamzo cum viculis earum et habitaverunt in eis.
2CHR|28|19|Humiliaverat enim Dominus Iudam propter Achaz regem Israel, eo quod relaxasset ei frenum et contemptui habuisset Dominum.
2CHR|28|20|Venitque contra eum Theglathphalasar rex Assyriorum, qui afflixit eum, non autem confortavit.
2CHR|28|21|Achaz enim, spoliata domo Domini et domo regis et principum, dedit regi Assyriorum munera, et tamen nihil ei profuit.
2CHR|28|22|Insuper et in tempore angustiae suae auxit contemptum in Dominum. Ipse rex Achaz
2CHR|28|23|immolavit diis Damasci victimas percussoribus suis et dixit: " Dii regum Syriae auxiliantur eis; quos ego placabo hostiis, et aderunt mihi ", cum e contrario ipsi fuerint ruina ei et universo Israel.
2CHR|28|24|Direptis itaque Achaz omnibus vasis domus Dei atque confractis, clausit ianuas templi Dei et fecit sibi altaria in universis angulis Ierusalem.
2CHR|28|25|In singulis quoque urbibus Iudae exstruxit excelsa ad adolendum diis alienis atque ad iracundiam provocavit Dominum, Deum patrum suorum.
2CHR|28|26|Reliqua autem gestorum eius et omnium operum suorum priorum et novissimorum scripta sunt in libro regum Iudae et Israel.
2CHR|28|27|Dormivitque Achaz cum patribus suis, et sepelierunt eum in civitate Ierusalem; non autem posuerunt eum in sepulcra regum Israel. Regnavitque Ezechias filius eius pro eo.
2CHR|29|1|Igitur Ezechias regnare coepit, cum viginti quinque esset annorum, et viginti novem annis regnavit in Ierusalem. Nomen matris eius Abi filia Zachariae.
2CHR|29|2|Fecitque, quod erat placitum in conspectu Domini, iuxta omnia, quae fecerat David pater eius.
2CHR|29|3|Ipse anno et mense primo regni sui aperuit valvas domus Domini et instauravit eas.
2CHR|29|4|Adduxitque sacerdotes atque Levitas et congregavit eos in plateam orientalem
2CHR|29|5|dixitque ad eos: " Audite me, Levitae! Nunc sanctificamini; mundate domum Domini, Dei patrum vestrorum, et auferte omnem immunditiam de sanctuario.
2CHR|29|6|Peccaverunt patres nostri et fecerunt malum in conspectu Domini Dei nostri derelinquentes eum; averterunt facies suas a tabernaculo Domini et praebuerunt dorsum.
2CHR|29|7|Insuper clauserunt ostia, quae erant in porticu, et exstinxerunt lucernas incensumque non adoleverunt et holocausta non obtulerunt in sanctuario Deo Israel.
2CHR|29|8|Concitatus est itaque furor Domini super Iudam et Ierusalem; tradiditque eos in commotionem et in stuporem et in sibilum, sicut ipsi cernitis oculis vestris.
2CHR|29|9|En, corruerunt patres nostri gladiis, filii nostri et filiae nostrae et coniuges captivae ductae sunt propter hoc scelus.
2CHR|29|10|Nunc igitur placet mihi, ut ineam foedus cum Domino, Deo Israel, et avertat a nobis furorem irae suae.
2CHR|29|11|Filii mei, nolite neglegere; vos enim elegit Dominus, ut stetis coram eo et ministretis illi colatisque eum et adoleatis ".
2CHR|29|12|Surrexerunt ergo Levitae, Mahath filius Amasai et Ioel filius Azariae de filiis Caath; porro de filiis Merari Cis filius Abdi et Azarias filius Iallelel; de filiis autem Gerson Ioah filius Zimma et Eden filius Ioah;
2CHR|29|13|at vero de filiis Elisaphan Semri et Iehiel; de filiis quoque Asaph Zacharias et Matthanias;
2CHR|29|14|necnon de filiis Heman Iahiel et Semei; sed et de filiis Idithun Semeias et Oziel.
2CHR|29|15|Congregaveruntque fratres suos et sanctificati sunt et ingressi iuxta mandatum regis et imperium Domini, ut expiarent domum Dei.
2CHR|29|16|Sacerdotes quoque ingressi intra templum Domini, ut mundarent illud, extulerunt omnem immunditiam, quam intro reppererant in vestibulum domus Domini, quam tulerunt Levitae et asportaverunt ad torrentem Cedron foras.
2CHR|29|17|Coeperunt autem prima die mensis primi sanctificare et in die octava eiusdem mensis ingressi sunt porticum templi Domini et sanctificaverunt templum Domini diebus octo; et in die sexta decima mensis eiusdem, quod coeperant, impleverunt.
2CHR|29|18|Ingressi quoque sunt ad Ezechiam regem et dixerunt ei: " Mundavimus omnem domum Domini et altare holocausti vasaque eius necnon et mensam propositionis cum omnibus vasis suis
2CHR|29|19|cunctamque templi supellectilem, quam removerat rex Achaz in regno suo in praevaricatione sua, restituimus et sanctificavimus. Ecce exposita sunt omnia coram altari Domini ".
2CHR|29|20|Consurgensque diluculo Ezechias rex adunavit principes civitatis et ascendit domum Domini.
2CHR|29|21|Attuleruntque simul tauros septem, arietes septem, agnos septem et hircos septem pro peccato, pro regno, pro sanctuario, pro Iuda; dixit quoque sacerdotibus filiis Aaron, ut offerrent super altare Domini.
2CHR|29|22|Mactaverunt igitur tauros et susceperunt sacerdotes sanguinem et fuderunt illum super altare; mactaverunt etiam arietes et illorum sanguinem super altare fuderunt; immolaverunt agnos et fuderunt super altare sanguinem.
2CHR|29|23|Applicaverunt hircos pro peccato coram rege et universa multitudine imposueruntque manus suas super eos,
2CHR|29|24|et immolaverunt illos sacerdotes et asperserunt sanguinem eorum super altare pro piaculo universi Israelis; pro omni quippe Israel praeceperat rex, ut holocaustum fieret et pro peccato.
2CHR|29|25|Constituit quoque Levitas in domo Domini cum cymbalis et psalteriis et citharis secundum dispositionem David et Gad videntis regis et Nathan prophetae; siquidem Domini praeceptum fuit per manum prophetarum eius.
2CHR|29|26|Steteruntque Levitae tenentes organa David, et sacerdotes tubas.
2CHR|29|27|Et iussit Ezechias, ut offerrent holocaustum super altare; cumque offerretur holocaustum, coeperunt laudes canere Domino et clangere tubis atque in diversis organis David regis Israel concrepare.
2CHR|29|28|Omni autem turba adorante, cantores et ii, qui tenebant tubas, erant in officio suo, donec compleretur holocaustum.
2CHR|29|29|Cumque finita esset oblatio, incurvatus est rex et omnes, qui erant cum eo, et adoraverunt.
2CHR|29|30|Praecepitque Ezechias et principes Levitis, ut laudarent Dominum verbis David et Asaph videntis; qui laudaverunt eum magna laetitia et curvato genu adoraverunt.
2CHR|29|31|Ezechias autem etiam haec addidit: " Nunc, impletis manibus vestris Domino, accedite et afferte victimas et sacrificia pro gratiarum actione in domo Domini ". Attulit ergo universa multitudo hostias et sacrificia pro gratiarum actione, et omnis voluntarius et proni animi holocausta.
2CHR|29|32|Porro numerus holocaustorum, quae attulit multitudo, hic fuit: tauros septuaginta, arietes centum, agnos ducentos, in holocaustum Domino omnia haec.
2CHR|29|33|Sanctificaveruntque Domino boves sescentos et oves tria milia.
2CHR|29|34|Sacerdotes vero pauci erant nec poterant sufficere, ut pelles holocaustorum detraherent; unde et Levitae fratres eorum adiuverunt eos, donec impleretur opus, et sanctificarentur sacerdotes; Levitae quippe recti corde, ut sanctificarentur magis quam sacerdotes.
2CHR|29|35|Fuerunt igitur holocausta plurima, adipes pacificorum et libamina, quae pertinebant ad holocausta.Restitutus est ita cultus domus Domini.
2CHR|29|36|Laetatusque est Ezechias et omnis populus de eo, quod paravit Dominus populo; repente quippe hoc factum est.
2CHR|30|1|Misit quoque Ezechias ad omnem Israel et Iudam scri psitque et epistulas ad Ephraim et Manassen, ut venirent ad domum Domini in Ierusalem et facerent Pascha Domino, Deo Israel.
2CHR|30|2|Inito quoque consilio regis et principum et universi coetus in Ierusalem, decreverunt, ut facerent Pascha mense secundo.
2CHR|30|3|Non enim potuerant facere in tempore suo, quia sacerdotes, qui possent sufficere, sanctificati non fuerant, et populus necdum congregatus erat in Ierusalem.
2CHR|30|4|Placuit ergo sermo regi et omni multitudini,
2CHR|30|5|et decreverunt, ut mitterent nuntios in universum Israel de Bersabee usque Dan, ut venirent et facerent Pascha Domino, Deo Israel, in Ierusalem; in plurima enim multitudine non fecerant, sicut lege praescriptum est.
2CHR|30|6|Perrexeruntque cursores cum epistulis ex regis manu et principum eius in universum Israel et Iudam, iuxta quod rex iusserat, praedicantes: " Filii Israel, revertimini ad Dominum, Deum Abraham et Isaac et Israel, ut revertatur ad reliquias, quae effugerunt manum regum Assyriorum.
2CHR|30|7|Nolite fieri sicut patres vestri et fratres, qui recesserunt a Domino, Deo patrum suorum, et tradidit eos in interitum, ut ipsi cernitis.
2CHR|30|8|Nolite nunc indurare cervices vestras sicut patres vestri. Tradite manus Domino et venite ad sanctuarium eius, quod sanctificavit in aeternum; servite Domino Deo vestro, ut avertatur a vobis ira furoris eius.
2CHR|30|9|Si enim vos reversi fueritis ad Dominum, fratres vestri et filii habebunt misericordiam coram dominis suis, qui illos duxere captivos, et revertentur in terram hanc: misericors enim et clemens est Dominus Deus vester et non avertet faciem suam a vobis, si reversi fueritis ad eum ".
2CHR|30|10|Igitur cursores pergebant de civitate in civitatem per terram Ephraim et Manasse usque Zabulon, illis irridentibus et subsannantibus eos.
2CHR|30|11|Attamen quidam viri ex Aser et Manasse et Zabulon se humiliaverunt et venerunt Ierusalem.
2CHR|30|12|In Iuda quoque facta est manus Domini, ut daret eis cor unum, ut facerent praeceptum regis et principum iuxta verbum Domini.
2CHR|30|13|Congregatus est ergo in Ierusalem populus multus, ut faceret sollemnitatem Azymorum in mense secundo, ecclesia magna valde.
2CHR|30|14|Et surgentes destruxerunt altaria, quae erant in Ierusalem, atque universa thymiamateria subvertentes proiecerunt in torrentem Cedron.
2CHR|30|15|Et mactaverunt Pascha quarta decima die mensis secundi; sacerdotes autem atque Levitae confusi sanctificati sunt et attulerunt holocausta in domum Domini.
2CHR|30|16|Steteruntque in ordine suo iuxta dispositionem et legem Moysi hominis Dei, sacerdotes vero suscipiebant effundendum sanguinem de manibus Levitarum,
2CHR|30|17|eo quod multi in coetu sanctificati non essent; idcirco Levitae mactaverunt victimas Paschae omnibus, qui non erant mundi, ut sanctificarent illas Domino.
2CHR|30|18|Valde magna enim pars populi, de Ephraim et Manasse et Issachar et Zabulon, non erant mundati; et comederunt Pascha non iuxta, quod scriptum est. Et oravit pro eis Eze chias dicens: " Dominus bonus propitietur
2CHR|30|19|cunctis, qui direxerunt cor suum, ut requirerent Dominum, Deum patrum suorum, quamvis non secundum munditiam sanctuarii ".
2CHR|30|20|Quem exaudivit Dominus, et placatus est populo.
2CHR|30|21|Feceruntque filii Israel, qui inventi sunt in Ierusalem, sollemnitatem Azymorum septem diebus in laetitia magna, laudaverunt Dominum et per singulos dies Levitae et sacerdotes per organa benesonantia.
2CHR|30|22|Et locutus est Ezechias ad cor omnium Levitarum, qui habebant intellegentiam bonam super Domino; et compleverunt sollemnitatem septem dierum immolantes victimas pacificorum et laudantes Dominum, Deum patrum suorum.
2CHR|30|23|Placuitque universae multitudini, ut celebrarent etiam alios dies septem, quod et fecerunt cum ingenti gaudio.
2CHR|30|24|Ezechias enim rex Iudae praebuerat multitudini mille tauros et septem milia ovium; principes vero dederant populo tauros mille et oves decem milia; sanctificata est ergo sacerdotum plurima multitudo.
2CHR|30|25|Et hilaritate perfusa est omnis turba Iudae, tam sacerdotum et Levitarum quam universae frequentiae, quae venerat ex Israel, advenae quoque, qui venerant de terra Israel vel habitabant in Iuda.
2CHR|30|26|Factaque est grandis laetitia in Ierusalem, qualis a diebus Salomonis filii David regis Israel in ea urbe non fuerat.
2CHR|30|27|Surrexerunt autem sacerdotes levitici generis benedicentes populo; et exaudita est vox eorum, pervenitque oratio eorum in habitaculum sanctum eius in caelum.
2CHR|31|1|Cumque haec fuissent rite celebrata, egressus est omnis Israel, qui inventus fuerat in urbibus Iudae, et fregerunt simulacra succideruntque palos, demoliti sunt excelsa et altaria destruxerunt non solum de universo Iuda et Beniamin, sed et de Ephraim quoque et Manasse, donec penitus everterent. Reversique sunt omnes filii Israel in possessiones et civitates suas.
2CHR|31|2|Ezechias autem constituit turmas sacerdotales et leviticas per divisiones suas, unumquemque in officio proprio tam sacerdotum videlicet quam Levitarum, ad holocausta et pacifica, ut ministrarent et confiterentur canerentque laudes in portis castrorum Domini.
2CHR|31|3|Pars autem regis erat, ut de propria eius substantia offerretur holocaustum mane semper et vespere, sabbatis quoque et calendis et sollemnitatibus ceteris, sicut scriptum est in lege Moysi.
2CHR|31|4|Praecepit etiam populo habitanti Ierusalem, ut darent partes sacerdotibus et Levitis, ut possent vacare legi Domini.
2CHR|31|5|Quod cum percrebruisset in auribus multitudinis, plurimas obtulere primitias filii Israel frumenti, vini et olei, mellis quoque et omnium, quae gignit humus, et decimas obtulerunt de omnibus abundanter.
2CHR|31|6|Sed et filii Israel et Iudae, qui habitabant in urbibus Iudae, obtulerunt decimas boum et ovium decimasque sanctorum, quae sanctificabant Domino Deo suo; atque universa portantes fecerunt acervos plurimos.
2CHR|31|7|Mense tertio coeperunt acervorum iacere fundamenta et mense septimo compleverunt eos.
2CHR|31|8|Cumque ingressi fuissent Ezechias et principes, viderunt acervos et benedixerunt Domino ac populo Israel.
2CHR|31|9|Interrogavitque Ezechias sacerdotes et Levitas, cur ita iacerent acervi.
2CHR|31|10|Respondit illi Azarias sacerdos primus de stirpe Sadoc dicens: " Ex quo coeperunt offerre donationem in domum Domini, comedimus et saturati sumus, et remanserunt plurima, eo quod benedixerit Dominus populo suo; reliquiarum autem copia est ista, quam cernis ".
2CHR|31|11|Praecepit igitur Ezechias, ut praepararent cellas in domo Domini. Quod cum fecissent,
2CHR|31|12|intulerunt tam donationem quam decimas et quaecumque sanctificaverant fideliter. Fuit autem praefectus eorum Chonenias Levita et Semei frater eius secundus,
2CHR|31|13|post quem Iahiel et Azazias et Nahath et Asael et Ierimoth, Iozabad quoque et Eliel et Iesmachias et Mahath et Banaias praepositi sub manibus Choneniae et Semei fratris eius ex imperio Ezechiae regis et Azariae pontificis domus Dei.
2CHR|31|14|Core vero filius Iemna Levites et ianitor orientalis portae praepositus erat iis, quae sponte offerebantur Domino, ad distribuendum donationem Domini et sanctissima.
2CHR|31|15|Et sub cura eius Eden et Beniamin, Iesua et Semeias, Amarias quoque et Sechenias in civitatibus sacerdotum, ut fideliter distribuerent fratribus suis tam maioribus quam minoribus in divisionibus suis,
2CHR|31|16|dummodo recensiti essent mares ab annis tribus et supra, cuncti qui ingrediebantur templum Domini, ut singulorum dierum ministeria observarent iuxta divisiones suas.
2CHR|31|17|Sacerdotes recensiti erant per familias, et Levitae a vicesimo anno et supra per ministeria et turmas suas.
2CHR|31|18|Et recensita erat universa familia omnis turmae, tam pro uxoribus quam liberis eorum utriusque sexus, quia in fidelitate servitii ipsorum sanctificati erant omnes.
2CHR|31|19|Porro pro filiis Aaron, sacerdotibus in agris et suburbanis urbium singularum dispositi erant nominatim viri, qui partes distribuerent universo sexui masculino de sacerdotibus et omni, qui recensitus erat inter Levitas.
2CHR|31|20|Fecit ergo Ezechias secundum haec in omni Iuda operatusque est bonum et rectum et verum coram Domino Deo suo.
2CHR|31|21|Et in universo opere, quod coepit in servitio domus Dei, et iuxta legem et praeceptum volens requirere Deum suum, in toto corde suo operatus et prosperatus est.
2CHR|32|1|Post quae et huiuscemodi fidem venit Sennacherib rex Assyriorum et ingressus Iudam obsedit civitates munitas volens eas capere.
2CHR|32|2|Quod cum vidisset Ezechias, venisse scilicet Sennacherib et totum belli impetum verti contra Ierusalem,
2CHR|32|3|inito cum principibus consilio virisque fortissimis, ut obturarent capita fontium, qui erant extra urbem, et, hoc omnium decernente sententia,
2CHR|32|4|congregata est plurima multitudo, et obturaverunt cunctos fontes et rivum, qui fluebat in medio terrae, dicentes: " Ne veniant reges Assyriorum et inveniant aquarum abundantiam! ".
2CHR|32|5|Aedificavit quoque agens industrie omnem murum, qui fuerat dissipatus, et exstruxit turres desuper et forinsecus alterum murum instauravitque Mello in civitate David et fecit iacula plurima et clipeos.
2CHR|32|6|Constituitque principes belli super populum et convocavit illos ad se in platea portae civitatis ac locutus est ad cor eorum dicens:
2CHR|32|7|" Viriliter agite et confortamini! Nolite timere nec paveatis regem Assyriorum et universam multitudinem, quae est cum eo. Multo enim plures nobiscum sunt quam cum illo:
2CHR|32|8|cum illo est brachium carneum, nobiscum autem Dominus Deus noster, qui auxiliator est noster pugnatque pro nobis ". Confortatusque est populus huiuscemodi verbis Ezechiae regis Iudae.
2CHR|32|9|Quae postquam gesta sunt, misit Sennacherib rex Assyriorum servos suos Ierusalem - ipse enim cum universo exercitu obsidebat Lachis - ad Ezechiam regem Iudae et ad omnem populum, qui erat in urbe, dicens:
2CHR|32|10|" Haec dicit Sennacherib rex Assyriorum: In quo habentes fiduciam sedetis obsessi in Ierusalem?
2CHR|32|11|Nonne Ezechias decipit vos, ut tradat morti in fame et siti affirmans quod Dominus Deus vester liberet vos de manu regis Assyriorum?
2CHR|32|12|Numquid non iste est Ezechias, qui destruxit excelsa illius et altaria et praecepit Iudae et Ierusalem dicens: "Coram altari uno adorabitis et in ipso comburetis sacrificia"?
2CHR|32|13|An ignoratis quae ego fecerim et patres mei cunctis terrarum populis? Numquid praevaluerunt dii gentium terrarum liberare regionem suam de manu mea?
2CHR|32|14|Quis est de universis diis gentium, quas deleverunt patres mei, qui potuerit eruere populum suum de manu mea, ut possit etiam Deus vester eruere vos de hac manu?
2CHR|32|15|Non vos ergo decipiat Ezechias nec vana persuasione deludat, neque credatis ei! Si enim nullus potuit deus cunctarum gentium atque regnorum liberare populum suum de manu mea et de manu patrum meorum, quanto minus Deus vester poterit eruere vos de manu mea! ".
2CHR|32|16|Sed et alia multa locuti sunt servi eius contra Dominum Deum et contra Ezechiam servum eius.
2CHR|32|17|Epistulas quoque scripsit plenas blasphemiae in Dominum, Deum Israel, et locutus est adversus eum: " Sicut dii gentium terrarum non potuerunt liberare populos suos de manu mea, sic et Deus Ezechiae eruere non poterit populum suum de manu ista ".
2CHR|32|18|Insuper et clamore magno, lingua Iudaica, ad populum Ierusalem, qui sedebat in muro, personabant, ut terrerent et perturbarent eos et caperent civitatem.
2CHR|32|19|Locutusque est Sennacherib contra Deum Ierusalem sicut adversum deos populorum terrae opera manuum hominum.
2CHR|32|20|Oraverunt igitur Ezechias rex et Isaias filius Amos prophetes adversum hanc blasphemiam ac vociferati sunt in caelum.
2CHR|32|21|Et misit Dominus angelum, qui percussit omnem virum robustum et bellatorem et principem in castris regis Assyriorum; reversusque est cum ignominia in terram suam. Cumque ingressus esset domum dei sui, filii, qui egressi fuerant de visceribus eius, interfecerunt eum ibi gladio.
2CHR|32|22|Salvavit ergo Dominus Ezechiam et habitatores Ierusalem de manu Sennacherib regis Assyriorum et de manu omnium et praestitit eis quietem per circuitum.
2CHR|32|23|Multi etiam deferebant munera Domino in Ierusalem et res pretiosas Ezechiae regi Iudae, qui exaltatus est post haec coram cunctis gentibus.
2CHR|32|24|In diebus illis aegrotavit Ezechias usque ad mortem et oravit Dominum; exaudivitque eum et dedit ei signum.
2CHR|32|25|Sed non iuxta beneficia, quae acceperat, retribuit, quia elevatum est cor eius; et facta est contra eum ira et contra Iudam et Ierusalem.
2CHR|32|26|Humiliatusque est postea, eo quod exaltatum fuisset cor eius, tam ipse quam habitatores Ierusalem; et idcirco non venit super eos ira Domini in diebus Ezechiae.
2CHR|32|27|Fuit autem Ezechias dives et inclitus valde; et thesauros sibi plurimos congregavit argenti, auri et lapidis pretiosi, aromatum et clipeorum omnisque generis rerum pretiosarum.
2CHR|32|28|Apothecas quoque frumenti, vini et olei et praesepia omnium iumentorum caulasque pecoribus
2CHR|32|29|et urbes exaedificavit sibi; habebat quippe greges ovium et armentorum innumerabiles, eo quod dedisset ei Deus substantiam multam nimis.
2CHR|32|30|Ipse est Ezechias, qui obturavit superiorem exitum aquarum Gihon et avertit eas subter ad occidentem urbis David. In omnibus operibus suis prosperatus est.
2CHR|32|31|Attamen sic in legatione principum Babylonis, qui missi fuerant ad eum, ut interrogarent de portento, quod acciderat super terram, dereliquit eum Deus, ut tentaretur, et nota fierent omnia, quae erant in corde eius.
2CHR|32|32|Reliqua autem gestorum Ezechiae et misericordiarum eius scripta sunt in visione Isaiae filii Amos prophetae et in libro regum Iudae et Israel.
2CHR|32|33|Dormivitque Ezechias cum patribus suis, et sepelierunt eum in ascensu ad sepulcra filiorum David; et celebravit eius exsequias universus Iuda et omnes habitatores Ierusalem. Regnavitque Manasses filius eius pro eo.
2CHR|33|1|Duodecim annorum erat Manasses, cum regnare coe pisset, et quinquaginta quinque annis regnavit in Ierusalem.
2CHR|33|2|Fecit autem malum coram Domino iuxta abominationes gentium, quas expulit Dominus coram filiis Israel.
2CHR|33|3|Et conversus instauravit excelsa, quae demolitus fuerat Ezechias pater eius, construxitque aras Baalim et fecit palos et adoravit omnem militiam caeli et coluit eam.
2CHR|33|4|Aedificavit quoque altaria in domo Domini, de qua dixerat Dominus: " In Ierusalem erit nomen meum in aeternum ".
2CHR|33|5|Aedificavit autem ea cuncto exercitui caeli in duobus atriis domus Domini.
2CHR|33|6|Transireque fecit filios suos per ignem in valle filii Ennom. Hariolatus est, sectabatur auguria, maleficis artibus inserviebat, habebat secum pythones et aruspices; multaque mala operatus est coram Domino, ut irritaret eum.
2CHR|33|7|Posuit quoque sculptile, idolum, quod fecerat, in domo Dei, de qua locutus est Deus ad David et ad Salomonem filium eius dicens: " In domo hac et in Ierusalem, quam elegi de cunctis tribubus Israel, ponam nomen meum in sempiternum.
2CHR|33|8|Et moveri non faciam pedem Israel de terra, quam tradidi patribus eorum, ita dumtaxat si custodierint facere, quae praecepi eis, cunctamque legem et praecepta atque iudicia, per manum Moysi ".
2CHR|33|9|Igitur Manasses seduxit Iudam et habitatores Ierusalem, ut facerent malum super omnes gentes, quas subverterat Dominus a facie filiorum Israel.
2CHR|33|10|Locutusque est Dominus ad eum et ad populum illius, et attendere noluerunt.
2CHR|33|11|Idcirco superinduxit eis principes exercitus regis Assyriorum; ceperuntque Manassen compedibus et vinctum catenis duxerunt Babylonem.
2CHR|33|12|Qui, postquam coangustatus est, oravit Dominum Deum suum et egit paenitentiam valde coram Deo patrum suorum.
2CHR|33|13|Deprecatusque est eum, et placatus ei exaudivit orationem eius reduxitque eum Ierusalem in regnum suum; et cognovit Manasses quod Dominus ipse esset Deus.
2CHR|33|14|Post haec aedificavit murum extra civitatem David ad occidentem Gihon in convalle et ad introitum portae Piscium per circuitum Ophel et exaltavit illum vehementer; constituitque principes exercitus in cunctis civitatibus Iudae munitis.
2CHR|33|15|Et abstulit deos alienos et idolum de domo Domini, aras quoque, quas fecerat in monte domus Domini et in Ierusalem, et proiecit omnia extra urbem.
2CHR|33|16|Porro instauravit altare Domini et immolavit super illud victimas pacificorum et pro gratiarum actione praecepitque Iudae, ut serviret Domino, Deo Israel.
2CHR|33|17|Attamen adhuc populus immolabat in excelsis Domino Deo suo.
2CHR|33|18|Reliqua autem gestorum Manasse et obsecratio eius ad Deum suum, verba quoque videntium, qui loquebantur ad eum in nomine Domini, Dei Israel, continentur in sermonibus regum Israel.
2CHR|33|19|Oratio quoque eius et exauditio et cuncta peccata atque contemptus, loca etiam, in quibus aedificavit excelsa et fecit palos et statuas, antequam ageret paenitentiam, scripta sunt in sermonibus Hozai.
2CHR|33|20|Dormivit ergo Manasses cum patribus suis, et sepelierunt eum in domo sua. Regnavitque pro eo filius eius Amon.
2CHR|33|21|Viginti duorum annorum erat Amon, cum regnare coepisset, et duobus annis regnavit in Ierusalem.
2CHR|33|22|Fecitque malum in conspectu Domini, sicut fecerat Manasses pater eius, et cunctis idolis, quae Manasses fuerat fabricatus, immolavit atque servivit.
2CHR|33|23|Et non humiliavit se ante faciem Domini, sicut humiliaverat se Manasses pater eius, et multo maiora deliquit.
2CHR|33|24|Cumque coniurassent adversus eum servi sui, interfecerunt eum in domo sua.
2CHR|33|25|Porro populus terrae, caesis omnibus, qui conspiraverant contra regem Amon, consti tuit regem Iosiam filium eius pro eo.
2CHR|34|1|Octo annorum erat Iosias, cum regnare coepisset, et tri ginta et uno annis regnavit in Ierusalem.
2CHR|34|2|Fecitque quod erat rectum in conspectu Domini, et ambulavit in viis David patris sui; non declinavit neque ad dextram neque ad sinistram.
2CHR|34|3|Octavo autem anno regni sui, cum adhuc esset puer, coepit quaerere Deum patris sui David; et duodecimo anno coepit mundare Iudam et Ierusalem ab excelsis et palis sculptilibusque et conflatilibus.
2CHR|34|4|Destruxeruntque coram eo aras Baalim; et thymiamateria, quae eis superposita fuerant, demolitus est; palos etiam et sculptilia et conflatilia succidit atque comminuit et super tumulos eorum, qui eis immolare consueverant, fragmenta dispersit.
2CHR|34|5|Ossa praeterea sacerdotum combussit in altaribus ipsorum; mundavitque Iudam et Ierusalem,
2CHR|34|6|sed et in urbibus Manasse et Ephraim et Simeon usque Nephthali, in plateis eorum undique
2CHR|34|7|dissipavit altaria et palos et sculptilia contrivit in frusta; cunctaque thymiamateria demolitus est de universa terra Israel et reversus est Ierusalem.
2CHR|34|8|Igitur anno octavo decimo regni sui, cum mundaret terram et domum, misit Saphan filium Eseliae et Maasiam principem civitatis et Ioah filium Ioachaz a commentariis, ut instaurarent domum Domini Dei sui.
2CHR|34|9|Qui venerunt ad Helciam sacerdotem magnum acceptamque ab eo pecuniam, quae illata fuerat in domum Domini, et quam congregaverant Levitae ianitores de Manasse et Ephraim et universis reliquiis Israel ab omni quoque Iuda et Beniamin et habitatoribus Ierusalem,
2CHR|34|10|tradiderunt in manibus opificum, qui praeerant in domo Domini, et illi dederunt eam operariis, qui operabantur in domo Domini, ut instaurarent templum et infirma quaeque sarcirent;
2CHR|34|11|dederunt scilicet eam lignariis et caementariis, ut emerent lapides dolatos et ligna ad commissuras aedificii et ad contignationem domorum, quas destruxerant reges Iudae.
2CHR|34|12|Qui fideliter cuncta faciebant. Erant autem praepositi operantium Iahath et Abdias Levitae de filiis Merari, Zacharias et Mosollam de filiis Caath, qui dirigebant opus. Omnes autem Levitae scientes organis canere
2CHR|34|13|erant super eos, qui onera portabant et dirigebant omnes, qui varia opera faciebant. De Levitis quoque erant scribae et praefecti et ianitores.
2CHR|34|14|Cumque efferrent pecuniam, quae illata fuerat in templum Domini, repperit Helcias sacerdos librum legis Domini per manum Moysi
2CHR|34|15|et ait ad Saphan scribam: " Librum legis inveni in domo Domini ". Et tradidit ei.
2CHR|34|16|At ille intulit volumen ad regem et insuper nuntiavit ei dicens: " Omnia, quae dedisti in manu servorum tuorum, ecce complentur.
2CHR|34|17|Argentum, quod repertum est in domo Domini, effuderunt, datum que est praefectis et operariis ".
2CHR|34|18|Et nuntiavit Saphan scriba regi dicens: " Librum tradidit mihi Helcias sacerdos ". Et legebat illum Saphan coram rege.
2CHR|34|19|Et factum est, cum audisset rex verba legis, scidit vestimenta sua
2CHR|34|20|et praecepit Helciae et Ahicam filio Saphan et Abdon filio Micha, Saphan quoque scribae et Asaiae servo regis dicens:
2CHR|34|21|" Ite et consulite Dominum pro me et pro reliquiis Israel et Iudae super sermonibus libri, qui repertus est. Magnus enim furor Domini effusus est super nos, eo quod non custodierint patres nostri verba Domini, ut facerent iuxta omnia, quae scripta sunt in isto volumine ".
2CHR|34|22|Abiit igitur Helcias et hi, qui simul a rege missi fuerant, ad Holdam propheten uxorem Sellum filii Thecuae filii Haraas custodis vestium, quae habitabat in Ierusalem in secunda, et locuti sunt ei iuxta verba haec.
2CHR|34|23|Et illa respondit eis: " Haec dicit Dominus, Deus Israel: Dicite viro, qui misit vos ad me:
2CHR|34|24|Haec dicit Dominus: Ecce ego inducam mala super locum istum et super habitatores eius, cuncta maledicta, quae scripta sunt in libro hoc, quem legerunt coram rege Iudae,
2CHR|34|25|quia dereliquerunt me et sacrificaverunt diis alienis, ut me ad iracundiam provocarent in cunctis operibus manuum suarum; idcirco effundetur furor meus super locum istum et non exstinguetur.
2CHR|34|26|Ad regem autem Iudae, qui misit vos pro Domino consulendo, sic loquimini: Haec dicit Dominus, Deus Israel: Quoniam audisti verba voluminis,
2CHR|34|27|atque emollitum est cor tuum, et humiliatus es in conspectu Dei super his, quae dicta sunt contra locum hunc et habitatores Ierusalem, humiliatusque coram me scidisti vestimenta tua et flevisti coram me, ego quoque audivi, dicit Dominus.
2CHR|34|28|Ecce colligam te ad patres tuos, et infereris in sepulcrum tuum in pace; nec videbunt oculi tui omne malum, quod ego inducturus sum super locum istum et super habitatores eius ".Rettuleruntque itaque regi cuncta, quae dixerat.
2CHR|34|29|At ille, convocatis universis maioribus natu Iudae et Ierusalem,
2CHR|34|30|ascendit domum Domini, unaque omnes viri Iudae et habitatores Ierusalem, sacerdotes et Levitae et cunctus populus a minimo usque ad maximum. Quibus audientibus, in domo Domini legit rex omnia verba voluminis foederis inventi in domo Domini.
2CHR|34|31|Et stans in gradu suo percussit foedus coram Domino, ut ambularet post eum et custodiret praecepta et testimonia et iustificationes eius in toto corde suo et in tota anima sua faceretque verba foederis scripta in hoc libro.
2CHR|34|32|Adiuravit quoque super hoc omnes, qui reperti fuerant in Ierusalem et Beniamin; et fecerunt habitatores Ierusalem iuxta pactum Domini, Dei patrum suorum.
2CHR|34|33|Abstulit ergo Iosias cunctas abominationes de universis regionibus filiorum Israel et fecit omnes, qui inventi erant in Israel, servire Domino Deo suo. Cunctis diebus eius non recesserunt a Domino, Deo patrum suorum.
2CHR|35|1|Fecit autem Iosias in Ierusalem Pascha Domino, quod immolatum est quarta decima die mensis primi.
2CHR|35|2|Et constituit sacerdotes in officiis suis confortavitque eos, ut ministrarent in domo Domini.
2CHR|35|3|Levitis quoque, qui erudiebant omnem Israel et consecrati erant Domino, locutus est: " Ponite arcam sanctam in templum, quod aedificavit Salomon filius David rex Israel; nequaquam eam ultra umeris portabitis. Nunc ministrate Domino Deo vestro et populo eius Israel.
2CHR|35|4|Et praeparate vos per familias vestras in divisionibus singulis, sicut scripsit David rex Israel, et descripsit Salomon filius eius;
2CHR|35|5|et ministrate in sanctuario partibus familiarum fratrum vestrorum, filiorum populi, singulis pars familiae Levitarum.
2CHR|35|6|Mactate ergo Pascha et sanctificamini et praeparate vos pro fratribus vestris, ut faciatis iuxta verbum, quod locu tus est Dominus in manu Moysi.
2CHR|35|7|Dedit praeterea Iosias omni populo, qui ibi inventus fuerat pro Pascha, agnos et haedos de gregibus triginta milia, boumque tria milia; haec de regis universa substantia.
2CHR|35|8|Duces quoque eius sponte obtulerunt, tam populo quam sacerdotibus et Levitis; porro Helcias et Zacharias et Iahiel principes domus Domini dederunt sacerdotibus ad faciendum Pascha pecora commixtim duo milia sescenta et boves trecentos.
2CHR|35|9|Chonenias autem, Semeias etiam et Nathanael fratres eius necnon Hasabias et Iehiel et Iozabad principes Levitarum dederunt ceteris Levitis ad celebrandum Pascha quinque milia pecorum et boves quingentos.
2CHR|35|10|Praeparatumque est ministerium, et steterunt sacerdotes in loco suo, Levitae quoque in turmis iuxta regis imperium.
2CHR|35|11|Et mactatum est Pascha; asperseruntque sacerdotes manu sua sanguinem, et Levitae detraxerunt pelles holocaustorum
2CHR|35|12|et separaverunt holocaustum, ut darent partibus familiarum populi, et offerretur Domino, sicut scriptum est in libro Moysi. De bobus quoque fecere similiter.
2CHR|35|13|Et assaverunt Pascha super ignem, iuxta quod lege praeceptum est; pacificas vero hostias coxerunt in lebetis et caccabis et ollis et festinato distribuerunt universae plebi.
2CHR|35|14|Sibi autem et sacerdotibus postea paraverunt; nam in oblatione holocaustorum et adipum usque ad noctem sacerdotes fuerant occupati, unde Levitae et sibi et sacerdotibus filiis Aaron paraverunt novissimis.
2CHR|35|15|Porro cantores filii Asaph stabant in loco suo, iuxta praeceptum David et Asaph et Heman et Idithun prophetarum regis; ianitores vero per portas singulas observabant, ita ut ne puncto quidem discederent a ministerio, quia fratres eorum Levitae paraverunt eis cibos.
2CHR|35|16|Omnis igitur cultus Domini rite praeparatus est in die illa, ut facerent Pascha et offerrent holocausta super altare Domini, iuxta praeceptum regis Iosiae.
2CHR|35|17|Feceruntque filii Israel, qui reperti fuerant ibi, Pascha in tempore illo et sollemnitatem Azymorum septem diebus.
2CHR|35|18|Non fuit simile huic in Israel a diebus Samuelis prophetae, sed nec quisquam de cunctis regibus Israel fecit Pascha sicut Iosias cum sacerdotibus et Levitis et omni Iuda et Israel, qui repertus fuerat, et habitantibus in Ierusalem.
2CHR|35|19|Octavo decimo anno regni Iosiae hoc Pascha celebratum est.
2CHR|35|20|Postquam instauraverat Iosias templum, ascendit Nechao rex Aegypti ad pugnandum in Charchamis iuxta Euphraten. Et processit in occursum eius Iosias.
2CHR|35|21|At ille, missis ad eum nuntiis, ait: " Quid mihi et tibi est, rex Iudae? Non adversum te hodie venio, sed contra aliam pugno domum, ad quam me Deus festinato ire praecepit. Desine adversum Deum facere, qui mecum est, ne interficiat te ".
2CHR|35|22|Noluit Iosias reverti, sed audacter praeparavit contra eum bellum nec acquievit sermonibus Nechao ex ore Dei; verum perrexit, ut dimicaret in campo Mageddo.
2CHR|35|23|Ibique vulneratus a sagittariis dixit pueris suis: " Educite me de proelio, quia oppido vulneratus sum ".
2CHR|35|24|Qui transtulerunt eum de curru in alterum currum eius et asportaverunt in Ierusalem. Mortuusque est et sepultus in sepulcris patrum suorum; et universus Iuda et Ierusalem luxerunt eum.
2CHR|35|25|Ieremias fecit planctum super Iosiam; et omnes cantores atque cantrices usque in praesentem diem lamentationes super Iosia replicant, et quasi lex obtinuit in Israel; ecce scriptum fertur in Lamentationibus.
2CHR|35|26|Reliqua autem gestorum Iosiae et misericordiae eius, quae lege praecepta sunt Domini,
2CHR|35|27|gesta quoque illius prima et novissima scripta sunt in libro regum Israel et Iudae.
2CHR|36|1|Tulit ergo populus terrae Ioachaz filium Iosiae et con stituit regem pro patre suo in Ierusalem.
2CHR|36|2|Viginti trium annorum erat Ioachaz, cum regnare coepisset, et tribus mensibus regnavit in Ierusalem.
2CHR|36|3|Amovit autem eum rex Aegypti, cum venisset Ierusalem, et condemnavit terram centum talentis argenti et talento auri.
2CHR|36|4|Constituitque regem pro eo Eliachim fratrem eius super Iudam et Ierusalem et vertit nomen eius Ioachim. Ipsum vero Ioachaz tulit secum et adduxit in Aegyptum.
2CHR|36|5|Viginti quinque annorum erat Ioachim, cum regnare coepisset, et undecim annis regnavit in Ierusalem; fecitque malum coram Domino Deo suo.
2CHR|36|6|Contra hunc ascendit Nabuchodonosor rex Chaldaeorum et vinctum catenis duxit in Babylonem,
2CHR|36|7|ad quam et ex vasis Domini transtulit et posuit ea in templo suo.
2CHR|36|8|Reliqua autem gestorum Ioachim et abominationum eius, quas operatus est, et quae inventa sunt contra eum, continentur in libro regum Israel et Iudae. Regnavitque autem Ioachin filius eius pro eo.
2CHR|36|9|Decem et octo annorum erat Ioachin, cum regnare coepisset, et tribus mensibus ac decem diebus regnavit in Ierusalem; fecitque malum in conspectu Domini.
2CHR|36|10|Cumque anni circulus volveretur, misit Nabuchodonosor rex, qui adduxerunt eum in Babylonem, asportatis simul pretiosissimis vasis domus Domini; regem vero constituit Sedeciam fratrem eius super Iudam et Ierusalem.
2CHR|36|11|Viginti et unius anni erat Sedecias, cum regnare coepisset, et undecim annis regnavit in Ierusalem.
2CHR|36|12|Fecitque malum in oculis Domini Dei sui nec humiliavit se coram Ieremia propheta loquente ad se ex ore Domini.
2CHR|36|13|Contra regem quoque Nabuchodonosor rebellavit, qui adiuraverat eum per Deum, et induravit cervicem suam et cor, ut non reverteretur ad Dominum, Deum Israel.
2CHR|36|14|Sed et universi principes sacerdotum et populus multiplicaverunt praevaricationes suas iuxta universas abominationes gentium et polluerunt domum Domini, quam sanctificaverat in Ierusalem.
2CHR|36|15|Mittebat autem Dominus, Deus patrum suorum, ad illos per manum nuntiorum suorum de nocte consurgens et cotidie commonens, eo quod parceret populo et habitaculo suo.
2CHR|36|16|At illi subsannabant nuntios Dei et parvipendebant sermones eius illudebantque prophetis, donec ascenderet furor Domini in populum eius, et esset nulla curatio.
2CHR|36|17|Adduxit enim super eos regem Chaldaeorum et interfecit iuvenes eorum gladio in domo sanctuarii sui; non est misertus adulescentis et virginis et senis nec decrepiti quidem, sed omnes tradidit in manibus eius.
2CHR|36|18|Universaque vasa domus Dei tam maiora quam minora et thesauros templi et regis et principum transtulit in Babylonem.
2CHR|36|19|Incenderunt hostes domum Dei destruxeruntque murum Ierusalem, universa palatia combusserunt et, quidquid pretiosum fuerat, demoliti sunt.
2CHR|36|20|Si quis evaserat gladium, ductus in Babylonem servivit regi et filiis eius, donec imperaret rex Persarum,
2CHR|36|21|ut compleretur sermo Domini ex ore Ieremiae: donec terra acciperet sabbata sua, cunctis diebus devastationis egit sabbatum, usque dum complerentur septuaginta anni.
2CHR|36|22|Anno autem primo Cyri regis Persarum ad explendum sermonem Domini, quem locutus fuerat per os Ieremiae, suscitavit Dominus spiritum Cyri regis Persarum, qui iussit praedicari in universo regno suo etiam per scripturam dicens:
2CHR|36|23|" Haec dicit Cyrus rex Persarum: Omnia regna terrae dedit mihi Dominus, Deus caeli, et ipse praecepit mihi, ut aedificarem ei domum in Ierusalem, quae est in Iudaea. Quis ex vobis est de omni populo eius? Sit Dominus Deus suus cum eo, et ascendat ".
EZRA|1|1|In anno primo Cyri regis Persarum, ut compleretur verbum Domini ex ore Ieremiae, suscitavit Dominus spiritum Cyri regis Persarum, qui emisit edictum in omni regno suo etiam per scripturam dicens:
EZRA|1|2|" Haec dicit Cyrus rex Persarum: Omnia regna terrae dedit mihi Dominus, Deus caeli, et ipse praecepit mihi, ut aedificarem ei domum in Ierusalem, quae est in Iudaea.
EZRA|1|3|Quis ex vobis est de omni populo eius? Sit Dominus Deus suus cum eo, et ascendat in Ierusalem, quae est in Iudaea, et aedificet domum Domini, Dei Israel; ipse est Deus, qui est in Ierusalem.
EZRA|1|4|Et omnes reliqui in cunctis locis, ubicumque habitant, adiuventur a viris de loco suo, argento et auro et substantia et pecore sicut et oblationibus spontaneis pro templo Dei, quod est in Ierusalem ".
EZRA|1|5|Et surrexerunt principes familiarum de Iuda et Beniamin et sacerdotes et Levitae et omnis, cuius Deus suscitavit spiritum, ut ascenderent ad aedificandum templum Domini, quod erat in Ierusalem.
EZRA|1|6|Universique, qui erant in circuitu, confortaverunt manus eorum cum vasis argenteis et aureis, substantia, pecore et pensitationibus, praeter oblationes spontaneas.
EZRA|1|7|Rex quoque Cyrus protulit vasa templi Domini, quae tulerat Nabuchodonosor de Ierusalem et posuerat ea in templo dei sui;
EZRA|1|8|protulit autem ea Cyrus rex Persarum per manum Mithridatis praepositi thesauri, qui enumeravit ea Sasabassar principi Iudae.
EZRA|1|9|Et hic est numerus eorum: phialae aureae triginta, phialae argenteae mille, cultri viginti novem, scyphi aurei triginta,
EZRA|1|10|scyphi quoque argentei quadringenti decem, vasa alia plurima; 11 omnia vasa aurea et argentea quinque milia quadringenta. Universa tulit Sasabassar cum his, qui ascendebant de transmigratione Babylonis in Ierusalem.
EZRA|2|1|Hi sunt autem provinciae filii, qui ascenderunt de captivitate migrantium, quos transtulerat Nabuchodonosor rex Babylonis in Babylonem, et reversi sunt in Ierusalem et Iudam, unusquisque in civitatem suam.
EZRA|2|2|Qui venerunt cum Zorobabel, Iesua, Nehemias, Saraia, Rahelaia, Mardochaeus, Belsan, Mesphar, Beguai, Rehum, Baana.Numerus virorum populi Israel:
EZRA|2|3|filii Pharos duo milia centum septuaginta duo;
EZRA|2|4|filii Saphatia trecenti septuaginta duo;
EZRA|2|5|filii Area septingenti septuaginta quinque;
EZRA|2|6|filii Phahathmoab, hi sunt filii Iesua et Ioab, duo milia octingenti duodecim;
EZRA|2|7|filii Elam mille ducenti quinquaginta quattuor;
EZRA|2|8|filii Zethua nongenti quadraginta quinque;
EZRA|2|9|filii Zachai septingenti sexaginta;
EZRA|2|10|filii Bani sescenti quadraginta duo;
EZRA|2|11|filii Bebai sescenti viginti tres;
EZRA|2|12|filii Azgad mille ducenti viginti duo;
EZRA|2|13|filii Adonicam sescenti sexaginta sex;
EZRA|2|14|filii Beguai duo milia quinquaginta sex;
EZRA|2|15|filii Adin quadringenti quinquaginta quattuor;
EZRA|2|16|filii Ater, qui erant ex Ezechia, nonaginta octo;
EZRA|2|17|filii Besai trecenti viginti tres;
EZRA|2|18|filii Iora centum duodecim;
EZRA|2|19|filii Hasum ducenti viginti tres;
EZRA|2|20|filii Gebbar nonaginta quinque;
EZRA|2|21|filii Bethlehem centum viginti tres;
EZRA|2|22|viri Netopha quinquaginta sex;
EZRA|2|23|viri Anathoth centum viginti octo;
EZRA|2|24|filii Azmaveth quadraginta duo;
EZRA|2|25|filii Cariathiarim, Cephira et Beroth septingenti quadraginta tres;
EZRA|2|26|filii Rama et Gabaa sescenti viginti unus;
EZRA|2|27|viri Machmas centum viginti duo;
EZRA|2|28|viri Bethel et Hai ducenti viginti tres;
EZRA|2|29|filii Nabo quinquaginta duo;
EZRA|2|30|filii Megbis centum quinquaginta sex;
EZRA|2|31|filii Elam alterius mille ducenti quinquaginta quattuor;
EZRA|2|32|filii Harim trecenti viginti;
EZRA|2|33|filii Lod, Hadid et Ono septingenti viginti quinque;
EZRA|2|34|filii Iericho trecenti quadraginta quinque;
EZRA|2|35|filii Senaa tria milia sescenti triginta.
EZRA|2|36|Sacerdotes: filii Iedaia de domo Iesua nongenti septuaginta tres,
EZRA|2|37|filii Emmer mille quinquaginta duo,
EZRA|2|38|filii Phassur mille ducenti quadraginta septem,
EZRA|2|39|filii Harim mille decem et septem.
EZRA|2|40|Levitae: filii Iesua, hi sunt filii Cadmihel, Bennui, Odoviae, septuaginta quattuor.
EZRA|2|41|Cantores: filii Asaph centum viginti octo.
EZRA|2|42|Ianitores: filii Sellum, filii Ater, filii Telmon, filii Accub, filii Hatita, filii Sobai: universi centum triginta novem.
EZRA|2|43|Oblati: filii Siha, filii Hasupha, filii Tabbaoth,
EZRA|2|44|filii Ceros, filii Siaa, filii Phadon,
EZRA|2|45|filii Lebana, filii Hagaba, filii Accub,
EZRA|2|46|filii Hagab, filii Semlai, filii Hanan,
EZRA|2|47|filii Giddel, filii Gaher, filii Raaia,
EZRA|2|48|filii Rasin, filii Necoda, filii Gazam,
EZRA|2|49|filii Oza, filii Phasea, filii Besai,
EZRA|2|50|filii Asena, filii Meunitarum, filii Nephusorum,
EZRA|2|51|filii Bacbuc, filii Hacupha, filii Harhur,
EZRA|2|52|filii Basluth, filii Mahida, filii Harsa,
EZRA|2|53|filii Bercos, filii Sisara, filii Thema,
EZRA|2|54|filii Nasia, filii Hatipha.
EZRA|2|55|Filii servorum Salomonis: filii Sotai, filii Sophereth, filii Pheruda,
EZRA|2|56|filii Iaala, filii Darcon, filii Giddel,
EZRA|2|57|filii Saphatia, filii Hatil, filii Phochereth Hassebaim, filii Ami.
EZRA|2|58|Omnes oblati et filii servorum Salomonis trecenti nonaginta duo.
EZRA|2|59|Et hi, qui ascenderunt de Thelmela, Thelharsa, Cherub et Addon et Emmer et non potuerunt indicare domum patrum suorum et semen suum, utrum ex Israel essent:
EZRA|2|60|filii Dalaia, filii Tobia, filii Necoda, sescenti quinquaginta duo.
EZRA|2|61|Et de filiis sacerdotum: filii Hobia, filii Accos, filii Berzellai, qui accepit de filiabus Berzellai Galaaditis uxorem et vocatus est nomine eorum.
EZRA|2|62|Hi quaesierunt tabulas genealogiae suae et non invenerunt; et eiecti sunt de sacerdotio.
EZRA|2|63|Et dixit praepositus eis, ut non comederent de sanctificatis sanctuarii, donec surgeret sacerdos pro Urim et Tummim.
EZRA|2|64|Omnis multitudo simul quadraginta duo milia trecenti sexaginta,
EZRA|2|65|exceptis servis eorum et ancillis, qui erant septem milia trecenti triginta septem, insuper et cantores atque cantatrices ducenti.
EZRA|2|66|Equi eorum septingenti triginta sex, muli eorum ducenti quadraginta quinque,
EZRA|2|67|cameli eorum quadringenti triginta quinque, asini eorum sex milia septingenti viginti.
EZRA|2|68|Nonnulli autem de principibus familiarum, cum ingrederentur templum domini, quod est in Ierusalem, sponte obtulerunt in domum Dei ad exstruendam eam in loco suo.
EZRA|2|69|Se cundum vires suas dederunt in aerarium operis auri solidos sexaginta milia et mille, argenti minas quinque milia et vestes sacerdotales centum.
EZRA|2|70|Habitaverunt ergo ibi sacerdotes et Levitae et quidam de populo; cantores autem et ianitores et oblati in urbibus suis, universusque Israel in civitatibus suis.
EZRA|3|1|Iamque venerat mensis septi mus, et erant filii Israel in civita tibus suis. Congregatus est ergo populus quasi vir unus in Ierusalem.
EZRA|3|2|Et surrexit Iesua filius Iosedec et fratres eius sacerdotes et Zorobabel filius Salathiel et fratres eius et aedificaverunt altare Dei Israel, ut offerrent in eo holocautomata, sicut scriptum est in lege Moysi viri Dei.
EZRA|3|3|Collocaverunt autem altare super bases suas, deterrentibus eos per circuitum populis terrarum, et obtulerunt super illud holocaustum Domino mane et vespere.
EZRA|3|4|Feceruntque sollemnitatem Tabernaculorum, sicut scriptum est, et holocaustum diebus singulis per ordinem, secundum praeceptum pro singulis diebus;
EZRA|3|5|et praeter holocaustum sempiternum illa etiam pro calendis et universis sollemnitatibus, quae erant consecratae Domino, et pro omnibus, quae ultro offerebantur Domino.
EZRA|3|6|A primo die mensis septimi coeperunt offerre holocaustum Domino; porro templum Dei nondum fundatum erat.
EZRA|3|7|Dederunt autem pecunias latomis et fabris, cibum quoque et potum et oleum Sidoniis Tyriisque, ut deferrent ligna cedrina de Libano ad mare Ioppe, iuxta quod concesserat Cyrus rex Persarum eis.
EZRA|3|8|Anno autem secundo adventus eorum ad templum Dei in Ierusalem mense secundo, coeperunt Zorobabel filius Salathiel et Iesua filius Iosedec et reliqui de fratribus eorum sacerdotes et Levitae et omnes, qui venerant de captivitate in Ierusalem, et constituerunt Levitas a viginti annis et supra, ut dirigerent opus templi Domini.
EZRA|3|9|Stetitque Iesua et filii eius et fratres eius, Cadmihel, Bennui et Odovia quasi vir unus, ut dirigerent eos, qui faciebant opus in templo Dei; itemque filii Henadad et filii eorum et fratres eorum Levitae.
EZRA|3|10|Fundato igitur ab aedificatoribus templo Domini, steterunt sacerdotes in ornatu suo cum tubis, et Levitae filii Asaph in cymbalis, ut laudarent Deum iuxta mandatum David regis Israel.
EZRA|3|11|Et concinebant in hymnis et gratiarum actione Domino: " Quoniam bonus, quoniam in aeternum misericordia eius " super Israel. Omnis quoque populus vociferabatur clamore magno in laudando Dominum, eo quod fundatum esset templum Domini.
EZRA|3|12|Plurimi etiam senes de sacerdotibus et Levitis et principibus familiarum, qui viderant oculis suis prius templum in loco suo, flebant voce magna; et multi vociferantes in laetitia elevabant vocem.
EZRA|3|13|Nec poterat quisquam agnoscere vocem clamoris laetantium et vocem fletus populi, quoniam populus vociferabatur clamore magno, et strepitus audiebatur procul.
EZRA|4|1|Audierunt autem hostes Iudae et Beniamin, quia filii captivita tis aedificarent templum Domino, Deo Israel,
EZRA|4|2|et accedentes ad Zorobabel et ad principes familiarum dixerunt eis: " Aedificemus vobiscum, quia ita ut vos quaerimus Deum vestrum et immolavimus victimas a diebus Asarhaddon regis Assyriae, qui adduxit nos huc ".
EZRA|4|3|Et dixit eis Zorobabel et Iesua et reliqui principes familiarum Israel: Non est vobis et nobis, ut aedificemus domum Deo nostro, sed nos ipsi soli aedificabimus Domino, Deo Israel, sicut praecepit nobis Cyrus rex Persarum ".
EZRA|4|4|Factum est igitur, ut populus terrae impediret manus populi Iudae et turbaret eos in aedificando.
EZRA|4|5|Conduxerunt autem adversus eos consiliatores, ut destruerent consilium eorum omnibus diebus Cyri regis Persarum et usque ad regnum Darii regis Persarum.
EZRA|4|6|In regno autem Asueri, in principio regni eius, scripserunt accusationem adversus habitatores Iudae et Ierusalem.
EZRA|4|7|Et in diebus Artaxerxis scripsit Beselam, Mithridates et Tabel et reliqui, qui erant in consilio eorum, ad Artaxerxem regem Persarum; scriptura autem accusationis erat scripta litteris Syriacis et composita sermone Syro.
EZRA|4|8|Rehum praefectus et Samsai scriba scripserunt epistulam unam de Ierusalem Artaxerxi regi huiuscemodi:
EZRA|4|9|" Rehum praefectus et Samsai scriba et reliqui socii eorum, iudices et duces, magistratus Persae, Erchuaei, Babylonii, Susanechaei, hoc est Elamitae,
EZRA|4|10|et ceteri de gentibus, quas transtulit Asenaphar magnus et gloriosus et habitare fecit in civitatibus Samariae et in reliquis regionibus trans flumen in pace ".
EZRA|4|11|Hoc est exemplar epistulae, quam miserunt ad eum: Artaxerxi regi, servi tui, viri, qui sunt trans fluvium. Igitur
EZRA|4|12|notum sit regi quia Iudaei, qui ascenderunt a te ad nos, venerunt in Ierusalem civitatem rebellem et pessimam, quam aedificant, exstruentes muros eius, fundamenta iam componentes.
EZRA|4|13|Nunc notum sit regi quia, si civitas illa aedificata fuerit, et muri eius instaurati, tributum et annonam et vectigal non dabunt, et ad ultimum regibus noxa erit.
EZRA|4|14|Nos autem, memores salis, quod in palatio comedimus, et quia laesiones regis videre nefas ducimus, idcirco misimus et nuntiavimus regi,
EZRA|4|15|ut recenseas in libris historiarum patrum tuorum, et invenies in his historiis et scies quoniam urbs illa urbs rebellis est et nocens regibus et provinciis, et seditiones concitantur in ea ex diebus antiquis; quam ob rem et civitas ipsa destructa est.
EZRA|4|16|Nuntiamus nos regi quoniam, si civitas illa aedificata fuerit, et muri ipsius instaurati, possessionem trans fluvium non habebis ".
EZRA|4|17|Verbum misit rex ad Rehum praefectum et Samsai scribam et ad reliquos, qui erant in consilio eorum, qui habitabant in Samaria et in regione trans fluvium: " Pax. Nunc igitur scriptura,
EZRA|4|18|quam misistis ad nos, manifeste lecta est coram me.
EZRA|4|19|Et a me praeceptum est, et recensuerunt inveneruntque quoniam civitas illa a diebus antiquis adversum reges rebellabat, et rebelliones et seditiones concitabantur in ea;
EZRA|4|20|nam et reges fortissimi fuerunt in Ierusalem, qui et dominati sunt omni regioni, quae trans fluvium est, tributum quoque et annonam et vectigal accipiebant.
EZRA|4|21|Nunc ergo praecipite, ut desistant isti homines, et urbs illa non aedificetur, donec forte a me iussum fuerit.
EZRA|4|22|Videte, ne negligenter hoc impleatis, et paulatim crescat malum contra reges ".
EZRA|4|23|Itaque exemplum edicti Artaxerxis regis lectum est coram Rehum praefectum et Samsai scriba et consiliariis eorum; et abierunt festini in Ierusalem ad Iudaeos et prohibuerunt eos in brachio et robore.
EZRA|4|24|Tunc intermissum est opus domus Domini in Ierusalem et non fiebat usque ad annum secundum regni Darii regis Persarum.
EZRA|5|1|Prophetae autem Aggaeus et Zacharias filius Addo propheta verunt ad Iudaeos, qui erant in Iudaea et Ierusalem, in nomine Dei Israel, quod erat super eos.
EZRA|5|2|Tunc surrexerunt Zorobabel filius Salathiel et Iesua filius Iosedec et coeperunt aedificare templum Dei in Ierusalem; prophetae autem Dei adiuvabant eos.
EZRA|5|3|In ipso autem tempore venit ad eos Thathanai, qui erat dux trans flumen, et Stharbuzanai et consiliarii eorum, sicque dixerunt eis: " Quis dedit vobis potestatem, ut domum hanc aedificaretis et materiam istam praepararetis?
EZRA|5|4|Quae sunt nomina hominum auctorum aedificationis illius? ".
EZRA|5|5|Oculus autem Dei eorum factus est super senes Iudaeorum, et non obstiterunt eis, usque dum res ad Darium referretur, et tunc sententia de hac re redderetur.
EZRA|5|6|Exemplar epistulae, quam misit Thathanai dux regionis trans flumen et Stharbuzanai et consiliatores eius et duces, qui erant trans flumen, ad Darium regem.
EZRA|5|7|Sermo, quem miserant ei, sic scriptus erat: Dario regi pax omnis.
EZRA|5|8|Notum sit regi isse nos ad Iudaeam provinciam, ad domum Dei magni, quae aedificatur lapide quadrato, et ligna ponuntur in parietibus; opusque illud diligenter exstruitur et crescit in manibus eorum.
EZRA|5|9|Interrogavimus ergo senes illos et ita diximus eis: "Quis dedit vobis potestatem, ut domum hanc aedificaretis et materiam istam praepararetis?".
EZRA|5|10|Sed et nomina eorum quaesivimus ab eis, ut nuntiaremus tibi, scripsimusque nomina eorum virorum, qui sunt principes in eis.
EZRA|5|11|Huiuscemodi autem sermonem responderunt nobis dicentes: "Nos sumus servi Dei caeli et terrae et aedificamus templum, quod erat exstructum ante hos annos multos, quodque rex Israel magnus aedificaverat et exstruxerat.
EZRA|5|12|Postquam autem ad iracundiam provocaverunt patres nostri Deum caeli, tradidit eos in manus Nabuchodonosor regis Babylonis Chaldaei, qui domum hanc destruxit et populum eius transtulit in Babylonem.
EZRA|5|13|Anno autem primo Cyri regis Babylonis, Cyrus rex proposuit edictum, ut domus Dei haec aedificaretur.
EZRA|5|14|Nam et vasa templi Dei aurea et argentea, quae Nabuchodonosor tulerat de templo, quod erat in Ierusalem, et asportaverat ea in templum Babylonis, protulit Cyrus rex de templo Babylonis, et data sunt viro cuidam nomine Sasabassar, quem et principem constituit,
EZRA|5|15|dixitque ei: 'Haec vasa tolle et vade et pone ea in templo, quod est in Ierusalem, et domus Dei aedificetur in loco suo'.
EZRA|5|16|Tunc itaque Sasabassar ille venit et posuit fundamenta templi Dei in Ierusalem, et ex eo tempore usque nunc aedificatur et necdum completum est".
EZRA|5|17|Nunc ergo, si videtur regi bonum, recenseat in aerario regis, quod est in Babylone, utrumnam a Cyro rege potestas data fuerit, ut aedificaretur domus Dei in Ierusalem, et voluntatem regis super hac re mittat ad nos ".
EZRA|6|1|Tunc Darius rex praecepit, et recensuerunt in tabulis aerarii, quod est in Babylone,
EZRA|6|2|et inventum est in Ecbatanis, quod est castrum in Medena provincia, volumen unum, et sic scriptus erat in eo commentarius:
EZRA|6|3|" Anno primo Cyri regis, Cyrus rex decrevit de domo Dei, quae est in Ierusalem: Aedificetur domus, ubi immolent et sacrificent; altitudo eius cubitorum sexaginta et latitudo eius cubitorum sexaginta,
EZRA|6|4|ordines de lapidibus quadratis tres et ordo de lignis unus; sumptus autem de domo regis dabuntur.
EZRA|6|5|Sed et vasa templi Dei aurea et argentea, quae Nabuchodonosor tulerat de templo Ierusalem et attulerat in Babylonem, reddantur et referantur in templum, quod est in Ierusalem, in locum suum, in templo Dei.
EZRA|6|6|Nunc ergo, Thathanai dux regionis, quae est trans flumen, Stharbuzanai et consiliarii eius et duces, qui estis trans flumen, procul recedite ab illo loco,
EZRA|6|7|dimittite fieri templum Dei illud; dux Iudaeorum et seniores eorum aedificent domum Dei illam in loco suo.
EZRA|6|8|Sed et a me praeceptum est quomodo agere debeatis cum senioribus Iudaeorum illis, qui aedificant domum Dei illam: ut de arca regis, id est de tributis, quae dantur de regione trans flumen, studiose sumptus dentur viris illis sine intermissione.
EZRA|6|9|Et si quid necesse fuerit, sive vituli et arietes et agni in holocaustum Deo caeli, sive frumentum, sal, vinum et oleum, secundum ordinationem sacerdotum, qui sunt in Ierusalem, detur eis per singulos dies sine neglegentia.
EZRA|6|10|Et offerant oblationes suaves Deo caeli orentque pro vita regis et filiorum eius.
EZRA|6|11|A me ergo positum est decretum, ut omnis homo, qui hanc mutaverit iussionem, tollatur lignum de domo ipsius et erigatur et configatur in eo; domus autem eius ponatur in sterquilinium.
EZRA|6|12|Deus autem, qui habitare fecit nomen suum ibi, dissipet omnia regna et populum, qui extenderit manum suam, ut contemnat et dissipet domum Dei illam, quae est in Ierusalem. Ego Darius statui decretum, quod studiose impleri volo ".
EZRA|6|13|Igitur Thathanai dux regionis trans flumen et duces et consiliarii eius, secundum quod praeceperat Darius rex, sic diligenter exsecuti sunt.
EZRA|6|14|Seniores autem Iudaeorum prosperabantur in aedificatione iuxta prophetiam Aggaei prophetae et Zachariae filii Addo et perfecerunt aedificationem, iubente Deo Israel et iubente Cyro et Dario et Artaxerxe regibus Persarum,
EZRA|6|15|et compleverunt domum Dei istam die tertia mensis Adar, qui est annus sextus regni Darii regis.
EZRA|6|16|Fecerunt autem filii Israel, sacerdotes et Levitae et reliqui filiorum transmigrationis dedicationem domus Dei illius in gaudio.
EZRA|6|17|Et obtulerunt in dedicationem domus Dei illius boves centum, arietes ducentos, agnos quadringentos, hircos caprarum pro peccato totius Israel duodecim, iuxta numerum tribuum Israel.
EZRA|6|18|Et statuerunt sacerdotes in ordinibus suis et Levitas in vicibus suis in ministerium Dei in Ierusalem, sicut scriptum est in libro Moysi.
EZRA|6|19|Fecerunt autem filii Israel transmigrationis Pascha quarta decima die mensis primi.
EZRA|6|20|Levitae universi se purificaverunt; purificati autem cuncti immolaverunt Pascha universis filiis transmigrationis et fratribus suis sacerdotibus et sibi.
EZRA|6|21|Et comederunt filii Israel, qui reversi fuerant de transmigratione, et omnes, qui a coinquinatione gentium terrae transierunt ad eos, ut quaererent Dominum, Deum Israel.
EZRA|6|22|Et fecerunt sollemnitatem Azymorum septem diebus in laetitia, quoniam laetificaverat eos Dominus et converterat cor regis Assyriae ad eos, ut adiuvaret manus eorum in opere domus Domini, Dei Israel.
EZRA|7|1|Post haec autem in regno Arta xerxis regis Persarum, Esdras fi lius Saraiae filii Azariae filii Helciae
EZRA|7|2|filii Sellum filii Sadoc filii Achitob
EZRA|7|3|filii Amariae filii Azariae filii Meraioth
EZRA|7|4|filii Zaraiae filii Ozi filii Bocci
EZRA|7|5|filii Abisue filii Phinees filii Eleazar filii Aaron summi sacerdotis,
EZRA|7|6|ipse Esdras ascendit de Babylone et ipse scriba velox in lege Moysi, quam dedit Dominus, Deus Israel. Cumque manus Domini Dei eius esset super eum, dedit ei rex omnem petitionem eius.
EZRA|7|7|Et ascenderunt de filiis Israel et de filiis sacerdotum et de filiis Levitarum et de cantoribus et de ianitoribus et de oblatis in Ierusalem, anno septimo Artaxerxis regis.
EZRA|7|8|Venit in Ierusalem mense quinto, ipse est annus septimus regis.
EZRA|7|9|In primo die mensis primi coepit ascendere de Babylone et in primo die mensis quinti venit in Ierusalem, iuxta manum Dei sui bonam super se.
EZRA|7|10|Esdras enim applicavit cor suum, ut investigaret et impleret legem Domini et faceret et doceret in Israel praeceptum et iudicium.
EZRA|7|11|Hoc est autem exemplar epistulae, quam dedit rex Artaxerxes Esdrae sacerdoti, scribae erudito in mandatis Domini et praeceptis eius in Israel.
EZRA|7|12|" Artaxerxes rex regum Esdrae sacerdoti, scribae legis Dei caeli, salutem.
EZRA|7|13|A me decretum est, ut cuicumque placuerit in regno meo de populo Israel et de sacerdotibus eius et de Levitis ire in Ierusalem, tecum vadat.
EZRA|7|14|A facie enim regis et septem consiliatorum eius missus es, ut visites Iudaeam et Ierusalem secundum legem Dei tui, quae est in manu tua,
EZRA|7|15|et ut feras argentum et aurum, quod rex et consiliatores eius sponte obtulerunt Deo Israel, cuius in Ierusalem tabernaculum est.
EZRA|7|16|Et omne argentum et aurum, quodcumque inveneris in universa provincia Babylonis simul cum oblationibus sponte oblatis a populo et a sacerdotibus pro domo Dei sui, quae est in Ierusalem,
EZRA|7|17|igitur studiose eme de hac pecunia boves, arietes, agnos et oblationes et libamina eorum et offer ea super altare templi Dei vestri, quod est in Ierusalem.
EZRA|7|18|Sed et, si quid tibi et fratribus tuis placuerit de reliquo argento et auro ut faciatis iuxta voluntatem Dei vestri, facite.
EZRA|7|19|Vasa quoque, quae dantur tibi in ministerium domus Dei tui, trade in conspectu Dei in Ierusalem.
EZRA|7|20|Sed et cetera, quibus opus fuerit in domum Dei tui, quantumcumque necesse est ut expendas, dabitur ab aerario regis.
EZRA|7|21|Et ego Artaxerxes rex statui atque decrevi omnibus custodibus arcae publicae, qui sunt trans flumen, ut quodcumque petierit a vobis Esdras sacerdos, scriba legis Dei caeli, absque mora detis
EZRA|7|22|usque ad argenti talenta centum et usque ad frumenti coros centum et usque ad vini batos centum et usque ad batos olei centum; sal vero absque mensura.
EZRA|7|23|Omne, quod requirit Deus caeli, tribuatur diligenter in domo Dei caeli, ne forte irascatur contra regnum regis et filiorum eius.
EZRA|7|24|Vobis quoque notum facimus de universis sacerdotibus et Levitis et cantoribus et ianitoribus, oblatis et ministris domus Dei huius, ut tributum et annonas et vectigal non habeatis potestatem imponendi super eos.
EZRA|7|25|Tu autem, Esdra, secundum sapientiam Dei tui, quae est in manu tua, constitue praesides et iudices, ut iudicent omni populo, qui est trans flumen, his videlicet, qui noverunt legem Dei tui; sed et imperitos docete.
EZRA|7|26|Et omnis, qui non fecerit legem Dei tui et legem regis diligenter, iudicium erit de eo, sive in mortem sive in exsilium sive in damnum substantiae eius vel certe in carcerem ".
EZRA|7|27|Benedictus Dominus, Deus patrum nostrorum, qui dedit hoc in corde regis, ut glorificaret domum Domini, quae est in Ierusalem,
EZRA|7|28|et in me inclinavit misericordiam regis et consiliariorum eius et cunctorum principum eius potentium. Et ego confortatus manu Domini Dei mei, quae erat in me, congregavi de Israel principes, qui ascenderent mecum.
EZRA|8|1|Hi sunt ergo principes familiarum et genealogia eorum, qui ascenderunt mecum in regno Artaxerxis regis de Babylone:
EZRA|8|2|De filiis Phinees, Gersom. De filiis Ithamar, Daniel. De filiis David, Hattus filius Secheniae.
EZRA|8|3|De filiis Pharos, Zacharias; et cum eo numerati sunt viri centum quinquaginta.
EZRA|8|4|De filiis Phahathmoab, Elioenai filius Zaraiae, et cum eo ducenti viri.
EZRA|8|5|De filiis Zethua, Sechenia filius Iahaziel, et cum eo trecenti viri.
EZRA|8|6|De filiis Adin, Ebed filius Ionathan, et cum eo quinquaginta viri.
EZRA|8|7|De filiis Elam, Iesaias filius Athaliae, et cum eo septuaginta viri.
EZRA|8|8|De filiis Saphatiae, Zabadia filius Michael, et cum eo octoginta viri.
EZRA|8|9|De filiis Ioab, Abdia filius Iahiel, et cum eo ducenti decem et octo viri.
EZRA|8|10|De filiis Bani, Selomith filius Iosphiae, et cum eo centum sexaginta viri.
EZRA|8|11|De filiis Bebai, Zacharias filius Bebai, et cum eo viginti octo viri.
EZRA|8|12|De filiis Azgad, Iohanan filius Eccetan, et cum eo centum et decem viri.
EZRA|8|13|De filiis Adonicam ascenderunt iuniores, et haec nomina eorum: Eliphalet et Iehiel et Semeias, et cum eis sexaginta viri.
EZRA|8|14|De filiis Beguai, Uthai filius Zabud, et cum eis septuaginta viri.
EZRA|8|15|Congregavi autem eos ad fluvium, qui decurrit ad Ahava, et mansimus ibi tribus diebus. Recensui populum et sacerdotes; de filiis autem Levi non inveni ibi.
EZRA|8|16|Itaque misi Eliezer et Ariel et Semeiam et Ioiarib et Elnathan et Nathan et Zachariam et Mosollam principes sapientes.
EZRA|8|17|Et misi eos ad Eddo, qui est primus in Chasphiae loco, et posui in ore eorum verba, quae loquerentur ad Eddo et fratres eius, ut adducerent nobis ministros domus Dei nostri.
EZRA|8|18|Et adduxerunt nobis per manum Dei nostri bonam super nos virum doctissimum de filiis Moholi filii Levi filii Israel nomine Serebiam et filios eius et fratres eius decem et octo
EZRA|8|19|et Hasabiam et cum eo Iesaiam de filiis Merari filiosque eius et fratres eius viginti
EZRA|8|20|et de oblatis, quos dederant David et principes ad ministeria Levitarum, ducentos viginti viros; omnes hi suis nominibus recensiti sunt.
EZRA|8|21|Et praedicavi ibi ieiunium iuxta fluvium Ahava, ut affligeremur coram Deo nostro et peteremus ab eo iter prosperum nobis et filiis nostris universaeque substantiae nostrae.
EZRA|8|22|Erubui enim petere a rege praesidium et equites, qui defenderent nos ab inimico in via, quia dixeramus regi: " Manus Dei nostri est super omnes, qui quaerunt eum in bonitate, et potentia eius et fortitudo eius super omnes, qui derelinquunt eum ".
EZRA|8|23|Ieiunavimus autem et rogavimus Deum nostrum per hoc, et evenit nobis prospere.
EZRA|8|24|Et separavi de principibus sacerdotum duodecim, Serebiam et Hasabiam et cum eis de fratribus eorum decem,
EZRA|8|25|appendique eis argentum et aurum et vasa: tributum domus Dei nostri, quod obtulerat rex et consiliatores eius et principes eius universusque Israel eorum, qui ibi inveniebantur.
EZRA|8|26|Et appendi in manibus eorum argenti talenta sescenta quinquaginta et vasa argentea centum, quae habebant talenta duo, auri centum talenta,
EZRA|8|27|et crateres aureos viginti, qui habebant solidos millenos, et vasa aeris fulgentis optimi duo pretiosa ut aurum.
EZRA|8|28|Et dixi eis: " Vos sancti Domini, et vasa sancta et argentum et aurum consecrata Domino, Deo patrum nostrorum;
EZRA|8|29|vigilate et custodite, donec appendatis coram principibus sacerdotum et Levitarum et ducibus familiarum Israel in Ierusalem, in habitaculis domus Domini ".
EZRA|8|30|Susceperunt autem sacerdotes et Levitae pondus argenti et auri et vasorum, ut deferrent Ierusalem in domum Dei nostri.
EZRA|8|31|Promovimus ergo a flumine Ahava duodecimo die mensis primi, ut pergeremus Ierusalem; et manus Dei nostri fuit super nos et liberavit nos de manu inimici et insidiatoris in via,
EZRA|8|32|et venimus Ierusalem et mansimus ibi tribus diebus.
EZRA|8|33|Die autem quarta appensum est argentum et aurum et vasa in domo Dei nostri per manum Meremoth filii Uriae sacerdotis et cum eo Eleazar filius Phinees cumque eis Iozabad filius Iesua et Noadia filius Bennui Levitae,
EZRA|8|34|iuxta numerum et pondus omnia; descriptumque est omne pondus. In tempore illo,
EZRA|8|35|qui venerant de captivitate, filii transmigrationis, obtulerunt holocautomata Deo Israel, vitulos duodecim pro omni populo Israel, arietes nonaginta sex, agnos septuaginta septem, hircos pro peccato duodecim: omnia in holocaustum Domino.
EZRA|8|36|Dederunt autem edicta regis satrapis regis et ducibus trans flumen et sublevaverunt populum et domum Dei.
EZRA|9|1|Postquam autem haec completa sunt, accesserunt ad me princi pes dicentes: " Non est separatus populus Israel, sacerdotes et Levitae a populis terrarum et abominationibus eorum, Chananaei videlicet et Hetthaei et Pherezaei et Iebusaei et Ammonitarum et Moabitarum et Aegyptiorum et Amorraeorum.
EZRA|9|2|Tulerunt enim de filiabus eorum sibi et filiis suis et commiscuerunt semen sanctum cum populis terrarum; manus etiam principum et magistratuum fuit in transgressione hac prima ".
EZRA|9|3|Cumque audissem sermonem istum, scidi vestimentum meum et pallium et evelli capillos capitis mei et barbae et sedi maerens.
EZRA|9|4|Convenerunt autem ad me omnes, qui timebant verba Dei Israel pro transgressione eorum, qui de captivitate venerant; et ego sedebam tristis usque ad sacrificium vespertinum.
EZRA|9|5|Et in sacrificio vespertino surrexi de afflictione mea et, scisso vestimento et pallio, curvavi genua mea et expandi manus meas ad Dominum Deum meum.
EZRA|9|6|Et dixi: " Deus meus, confundor et erubesco levare faciem meam ad te, quoniam iniquitates nostrae multiplicatae sunt super caput nostrum, et delicta nostra creverunt usque ad caelum
EZRA|9|7|a diebus patrum nostrorum. Peccavimus graviter usque ad diem hanc, et propter iniquitates nostras traditi sumus, ipsi et reges nostri et sacerdotes nostri, in manum regum terrarum et in gladium et in captivitatem et in rapinam et in confusionem vultus sicut et die hac.
EZRA|9|8|Et nunc ad momentum invenimus gratiam apud Dominum Deum nostrum, ut servaret nobis reliquias et figeret nobis tentorium in loco sancto eius et illuminaret oculos nostros Deus noster et daret nobis solacium modicum in servitute nostra.
EZRA|9|9|Quia servi sumus, et in servitute nostra non dereliquit nos Deus noster, sed inclinavit super nos misericordiam regum Persarum, ut darent nobis solacium, et erigeretur domus Dei nostri, et instaurarentur ruinae eius, et dedit nobis refugium in Iuda et Ierusalem.
EZRA|9|10|Et nunc quid dicemus, Deus noster, post haec? Dereliquimus mandata tua,
EZRA|9|11|quae praecepisti in manu servorum tuorum prophetarum dicens: "Terra, ad quam vos ingredimini, ut possideatis eam, terra immunda est, iuxta immunditiam populorum terrarum et abominationem eorum, qui repleverunt eam a fine usque ad finem coinquinatione sua.
EZRA|9|12|Nunc ergo filias vestras ne detis filiis eorum et filias eorum ne accipiatis filiis vestris et non quaeratis pacem eorum et prosperitatem eorum usque in aeternum, ut confortemini et comedatis, quae bona sunt terrae, et heredes habeatis filios vestros usque in saeculum".
EZRA|9|13|Et post omnia, quae venerunt super nos in operibus nostris pessimis et in delicto nostro magno, quia tu, Deus noster, non iudicasti secundum iniquitates nostras et dedisti nobis salutem, sicut est hodie,
EZRA|9|14|numquid amplius irrita faciemus mandata tua et matrimonia iungemus cum populis abominationum istarum? Numquid iratus es nobis usque ad consummationem, ut non essent reliquiae et salus?
EZRA|9|15|Domine, Deus Israel, tua clementia superstites sumus sicut die hac! Ecce coram te sumus in delicto nostro; non enim stari potest coram te propter hoc ".
EZRA|10|1|Dum ergo oraret Esdras et imploraret flens et prostratus ante templum Dei, collectus est ad eum de Israel coetus grandis nimis virorum et mulierum et puerorum; et flevit populus fletu multo.
EZRA|10|2|Et respondit Sechenias filius Iehiel de filiis Elam et dixit Esdrae: " Nos praevaricati sumus in Deum nostrum et duximus uxores alienigenas de populis terrae. Nunc autem spes est in Israel super hoc:
EZRA|10|3|percutiamus foedus cum Domino Deo nostro, ut proiciamus universas uxores et eos, qui de his nati sunt, iuxta voluntatem Domini et eorum, qui timent praeceptum Domini Dei nostri, et secundum legem fiat.
EZRA|10|4|Surge, tuum est decernere, nosque erimus tecum; confortare et fac ".
EZRA|10|5|Surrexit ergo Esdras et fecit principes sacerdotum et Levitarum et omnem Israel iurare, ut facerent secundum verbum hoc, et iuraverunt.
EZRA|10|6|Et surrexit Esdras ante domum Dei et abiit ad cubiculum Iohanan filii Eliasib et pernoctavit ibi; panem non comedit et aquam non bibit, lugebat enim transgressionem eorum, qui venerant de captivitate.
EZRA|10|7|Et missa est vox in Iuda et in Ierusalem omnibus filiis transmigrationis, ut congregarentur in Ierusalem;
EZRA|10|8|et omnis, qui non venerit in tribus diebus iuxta consilium principum et seniorum, auferetur universa substantia eius, et ipse abicietur de coetu transmigrationis.
EZRA|10|9|Convenerunt igitur omnes viri Iudae et Beniamin in Ierusalem tribus diebus, ipse est mensis nonus vicesimo die mensis, et sedit omnis populus in platea domus Dei, trementes pro peccato et pluviis.
EZRA|10|10|Et surrexit Esdras sacerdos et dixit ad eos: " Vos transgressi estis et duxistis uxores alienigenas, ut adderetis super delictum Israel.
EZRA|10|11|Et nunc date confessionem Domino, Deo patrum vestrorum, et facite placitum eius et separamini a populis terrae et ab uxoribus alienigenis ".
EZRA|10|12|Et respondit universa multitudo dixitque voce magna: " Iuxta verbum tuum ad nos, sic fiat.
EZRA|10|13|Verumtamen quia populus multus est et tempus pluviae, et non sustinemus stare foris, et opus non est diei unius vel duorum - multi quippe peccavimus in sermone isto -
EZRA|10|14|constituantur principes in universa multitudine; et omnes in civitatibus nostris, qui duxerunt uxores alienigenas, veniant in temporibus statutis, et cum his seniores per civitatem et civitatem et iudices eius, donec avertatur ira Dei nostri a nobis super peccato hoc ".
EZRA|10|15|Tantummodo Ionathan filius Asael et Iaasia filius Thecue steterunt contra hoc, et Mosollam et Sabethai Levites adiuverunt eos.
EZRA|10|16|Feceruntque sic filii transmigrationis. Et elegit Esdras sacerdos viros principes familiarum iuxta domus patrum eorum, omnes autem per nomina eorum, et sederunt in die primo mensis decimi, ut quaererent rem.
EZRA|10|17|Et absolverunt causam cunctorum, qui duxerant uxores alienigenas, intra diem primam mensis primi.
EZRA|10|18|Et inventi sunt de filiis sacerdotum, qui duxerant uxores alienigenas. De filiis Iesua filii Iosedec et de fratribus eius: Maasia et Eliezer et Iarib et Godolia;
EZRA|10|19|et dederunt manus suas, ut eicerent uxores suas et pro delicto suo arietem offerrent.
EZRA|10|20|Et de filiis Emmer: Hanani et Zabadia.
EZRA|10|21|Et de filiis Harim: Maasia et Elia et Semeia et Iehiel et Ozias.
EZRA|10|22|Et de filiis Phassur: Elioenai, Maasia, Ismael, Nathanael, Iozabad et Elasa.
EZRA|10|23|Et de filiis Levitarum: Iozabad et Semei et Celaia, ipse est Celita, Phethahia, Iuda et Eliezer.
EZRA|10|24|Et de cantoribus: Eliasib. Et de ianitoribus: Sellum et Telem et Uri.
EZRA|10|25|Et ex Israel de filiis Pharos: Remia et Iezia et Melchia et Miamin et Eleazar et Melchia et Banaia.
EZRA|10|26|Et de filiis Elam: Matthania, Zacharias et Iehiel et Abdi et Ierimoth et Elia.
EZRA|10|27|Et de filiis Zethua: Elioenai, Eliasib, Matthania et Ierimoth et Zabad et Aziza.
EZRA|10|28|Et de filiis Bebai: Iohanan, Hanania, Zabbai, Athalai.
EZRA|10|29|Et de filiis Beguai: Mosollam et Melluch et Adaia, Iasub et Saal et Ramoth.
EZRA|10|30|Et de filiis Phahathmoab: Edna et Chalal, Banaias et Maasias, Matthanias, Beseleel, Bennui et Manasse.
EZRA|10|31|Et de filiis Harim: Eliezer, Iesia, Melchias, Semeias, Simeon,
EZRA|10|32|Beniamin, Melluch, Samarias.
EZRA|10|33|Et de filiis Hasum: Matthanai, Matthatha, Zabad, Eliphalet, Iermai, Manasse, Semei.
EZRA|10|34|De filiis Bani: Maaddi, Amram et Ioel,
EZRA|10|35|Banaia et Badaias, Cheliau,
EZRA|10|36|Vania, Meremoth et Eliasib,
EZRA|10|37|Matthanias, Matthanai et Iasi.
EZRA|10|38|Et de filiis Bennui: Semei
EZRA|10|39|et Selemias et Nathan et Adaias
EZRA|10|40|et Mechnedebai, Sisai, Sarai,
EZRA|10|41|Azareel et Selemias, Samaria,
EZRA|10|42|Sellum, Amaria, Ioseph.
EZRA|10|43|De filiis Nabo: Iehiel, Matthathias, Zabad, Zabina, Ieddu et Ioel et Banaia.
EZRA|10|44|Omnes hi acceperant uxores alienigenas et dimiserunt uxores et filios.
NEH|1|1|Verba Nehemiae filii Hacha liae. Et factum est in mense Ca sleu, anno vicesimo, et ego eram in castro Susan.
NEH|1|2|Et venit Hanani unus de fratribus meis, ipse et viri ex Iuda; et interrogavi eos de Iudaeis, qui salvati erant et supererant de captivitate, et de Ierusalem.
NEH|1|3|Et dixerunt mihi: " Superstites, qui supererant de captivitate ibi in provincia, in afflictione magna sunt et in opprobrio; et murus Ierusalem dissipatus est, et portae eius combustae sunt igne ".
NEH|1|4|Cumque audissem verba huiuscemodi, sedi et flevi et luxi diebus multis; ieiunabam et orabam ante faciem Dei caeli.
NEH|1|5|Et dixi: " Quaeso, Domine, Deus caeli, Deus fortis, magne atque terribilis, qui custodis pactum et misericordiam cum his, qui te diligunt et custodiunt mandata tua;
NEH|1|6|fiat auris tua auscultans, et oculi tui aperti, ut audias orationem servi tui, quam ego oro coram te hodie, die et nocte pro filiis Israel servis tuis, et confiteor pro peccatis filiorum Israel, quibus peccaverunt tibi. Ego quoque et domus patris mei peccavimus,
NEH|1|7|delinquentes deliquimus contra te et non custodivimus praecepta et mandata et iudicia, quae praecepisti Moysi famulo tuo.
NEH|1|8|Memento verbi, quod mandasti Moysi servo tuo dicens: "Cum transgressi fueritis, ego dispergam vos in populos;
NEH|1|9|si autem revertamini ad me et custodiatis praecepta mea et faciatis ea, etiamsi abducti fueritis in extrema caeli, inde congregabo vos et reducam in locum quem elegi, ut habitaret nomen meum ibi".
NEH|1|10|Ipsi enim sunt servi tui et populus tuus, quos redemisti in fortitudine tua magna et in manu tua valida.
NEH|1|11|Obsecro, Domine, sit auris tua attendens ad orationem servi tui et ad orationem servorum tuorum, qui volunt timere nomen tuum; et fac servum tuum prosperari hodie et da ei gratiam ante virum hunc ". Ego enim eram pincerna regis.
NEH|2|1|Factum est autem in mense Nisan, anno vicesimo Artaxerxis regis, dum biberet, levavi vinum et dedi regi; non enim eram ingratus coram eo.
NEH|2|2|Dixitque mihi rex: " Quare vultus tuus tristis est, cum te aegrotum non videam? Nihil est aliud nisi tristitia cordis ". Et timui valde
NEH|2|3|et dixi regi: " Rex, in aeternum vive! Quare non maereat vultus meus, quia civitas sepulcrorum patrum meorum deserta est, et portae eius combustae sunt igne? ".
NEH|2|4|Et ait mihi rex: " Pro qua re postulas? ". Et oravi Deum caeli
NEH|2|5|et dixi ad regem: " Si videtur regi bonum, et si placet servus tuus ante faciem tuam, ut mittas me in Iudaeam ad civitatem sepulcrorum patrum meorum, et aedificabo eam ".
NEH|2|6|Dixitque mihi rex, et regina sedebat iuxta eum: " Usque ad quod tempus erit iter tuum, et quando reverteris? ". Et placuit regi mittere me; et constitui ei tempus.
NEH|2|7|Et dixi regi: " Si regi videtur bonum, epistulae dentur mihi ad duces regionis trans flumen, ut me transire permittant, donec veniam in Iudaeam;
NEH|2|8|et epistulam ad Asaph custodem saltus regis, ut det mihi ligna, ut contignare possim portas turris domus et muri civitatis et domus, in qua habitabo ". Et dedit mihi rex, quia manus Dei mei bona super me.
NEH|2|9|Et veni ad duces regionis trans flumen dedique eis epistulas regis. Miserat autem rex mecum principes militum et equites.
NEH|2|10|Et audierunt Sanaballat Horonites et Thobias servus Ammanites et contristati sunt afflictione magna, quod venisset homo, qui quaereret prosperitatem filiorum Israel.
NEH|2|11|Et veni Ierusalem et eram ibi tribus diebus.
NEH|2|12|Et surrexi nocte ego, et viri pauci mecum, et non indicavi cuiquam quid Deus meus dedisset in corde meo, ut facerem in Ierusalem; et iumentum non erat mecum, nisi animal cui sedebam.
NEH|2|13|Et egressus sum per portam Vallis nocte et ad fontem Draconis et portam Sterquilinii et considerabam murum Ierusalem dissipatum et portas eius consumptas igne.
NEH|2|14|Et transivi ad portam Fontis et ad piscinam Regis, et non erat locus iumento cui sedebam, ut transiret.
NEH|2|15|Et ascendi per torrentem nocte et considerabam murum; et iterum veni ad portam Vallis et reversus sum.
NEH|2|16|Magistratus autem nesciebant quo abissem aut quid ego facerem, sed et Iudaeis et sacerdotibus et optimatibus et magistratibus et reliquis, qui faciebant opus, usque ad id loci nihil indicaveram.
NEH|2|17|Et dixi eis: " Vos nostis afflictionem, in qua sumus, quia Ierusalem deserta est, et portae eius consumptae sunt igne; venite et aedificemus murum Ierusalem et non simus ultra opprobrium ".
NEH|2|18|Et indicavi eis quod manus Dei mei bona esset super me et verba regis, quae locutus esset mihi, et dixerunt: " Surgamus et aedificemus! ". Et confortatae sunt manus eorum in bonum.
NEH|2|19|Audierunt autem Sanaballat Horonites et Thobias servus Ammanites et Gosem Arabs et subsannaverunt nos et despexerunt dixeruntque: " Quae est haec res, quam facitis? Numquid contra regem vos rebellatis? ".
NEH|2|20|Et dedi eis responsum dicens: " Deus caeli ipse nos facit prosperari, et nos servi eius sumus; surgamus et aedificemus. Vobis autem non est pars et ius et memoria in Ierusalem ".
NEH|3|1|Et surrexit Eliasib sacerdos magnus et fratres eius sacerdotes et aedificaverunt portam Gregis; contignaverunt eam et statuerunt valvas eius et usque ad turrim Meah et turrim Hananeel.
NEH|3|2|Et iuxta eos aedificaverunt viri Iericho, et iuxta eos aedificavit Zacchur filius Imri.
NEH|3|3|Portam autem Piscium aedificaverunt filii Asnaa; ipsi contignaverunt eam et statuerunt valvas eius et seras et vectes.
NEH|3|4|Et iuxta eos restauravit Meremoth filius Uriae filii Accos, et iuxta eum restauravit Mosollam filius Barachiae filii Mesezabel, et iuxta eum restauravit Sadoc filius Baana,
NEH|3|5|et iuxta eum restauraverunt Thecueni; optimates autem eorum non supposuerunt colla sua in opere Domini sui.
NEH|3|6|Et portam Veterem restauraverunt Ioiada filius Phasea et Mosollam filius Besodia; ipsi contignaverunt eam et statuerunt valvas eius et seras et vectes.
NEH|3|7|Et iuxta eos restauraverunt Meltias Gabaonites et Iadon Meronathites, viri de Gabaon et Maspha, qui erant ad solium ducis, qui erat in regione trans flumen;
NEH|3|8|et iuxta eos restauravit Oziel filius Araia de aurificibus, et iuxta eum restauravit Hananias de pigmentariis et firmaverunt Ierusalem usque ad murum latiorem.
NEH|3|9|Et iuxta eum restauravit Raphaia filius Hur, princeps dimidiae partis vici Ierusalem;
NEH|3|10|et iuxta eum restauravit Iedaia filius Haromaph contra domum suam, et iuxta eum restauravit Hattus filius Hasabneia.
NEH|3|11|Alteram partem restauravit Melchias filius Harim et Hassub filius Phahathmoab usque ad turrim Furnorum.
NEH|3|12|Et iuxta eos restauravit Sellum filius Alohes, princeps mediae partis vici Ierusalem, ipse et filiae eius.
NEH|3|13|Portam Vallis restauravit Hanun et habitatores Zanoa; ipsi aedificaverunt eam et statuerunt valvas eius et seras et vectes et mille cubitos in muro usque ad portam Sterquilinii.
NEH|3|14|Et portam Sterquilinii restauravit Melchias filius Rechab, princeps vici Bethcharem; ipse aedificavit eam et statuit valvas eius et seras et vectes.
NEH|3|15|Et portam Fontis restauravit Sellum filius Cholhoza princeps pagi Maspha; ipse aedificavit eam et texit et statuit valvas eius et seras et vectes et murum piscinae Siloae iuxta hortum regis et usque ad gradus, qui descendunt de civitate David.
NEH|3|16|Post eum restauravit Nehemias filius Azboc princeps dimidiae partis vici Bethsur usque contra sepulcra David et usque ad piscinam, quae repleta est, et usque ad domum Fortium.
NEH|3|17|Post eum restauraverunt Levitae, Rehum filius Bani; iuxta eum restauravit Hasabias princeps dimidiae partis vici Ceilae pro vico suo;
NEH|3|18|post eum aedificaverunt fratres eorum Bavai filius Henadad princeps dimidiae partis vici Ceilae.
NEH|3|19|Et restauravit iuxta eum Ezer filius Iesua princeps Maspha mensuram alteram contra ascensum armentarii in angulo.
NEH|3|20|Post eum restauravit Baruch filius Zachai mensuram alteram ab angulo usque ad portam domus Eliasib sacerdotis magni.
NEH|3|21|Post eum restauravit Meremoth filius Uriae filii Aecos mensuram secundam a porta domus Eliasib usque ad extremitatem domus Eliasib.
NEH|3|22|Et post eum restauraverunt sacerdotes viri de campestribus.
NEH|3|23|Post eos restauravit Beniamin et Hassub contra domum suam; post eos restauravit Azarias filius Maasiae filii Ananiae iuxta domum suam.
NEH|3|24|Post eum restauravit Bennui filius Henadad mensuram alteram a domo Azariae usque ad angulum et flexuram.
NEH|3|25|Phalel filius Ozi contra angulum turris, quae eminet de domo regis excelsa in atrio carceris; post eum Phadaia filius Pharos restauravit
NEH|3|26|usque contra portam Aquarum ad orientem et turrim, quae prominebat.
NEH|3|27|Post eum restauraverunt Thecueni mensuram alteram a regione contra magnam turrim eminentem usque ad murum templi.
NEH|3|28|Sursum autem a porta Equorum restauraverunt sacerdotes, unusquisque contra domum suam.
NEH|3|29|Post eos restauravit Sadoc filius Emmer contra domum suam; et post eum restauravit Semeia filius Secheniae custos portae orientalis.
NEH|3|30|Post eum restauravit Hanania filius Selemiae et Hanun filius Seleph sextus mensuram alteram. Post eum restauravit Mosollam filius Barachiae contra cellam suam.
NEH|3|31|Post eum restauravit Melchias de aurificibus usque ad domum oblatorum et mercatorum, contra portam Iudicialem, et usque ad cenaculum anguli;
NEH|3|32|et inter cenaculum anguli et portam Gregis restauraverunt aurifices et negotiatores.
NEH|3|33|Factum est autem, cum audisset Sanaballat quod aedificaremus murum, iratus est et indignatus est nimis et subsannavit Iudaeos
NEH|3|34|et dixit coram fratribus suis et optimatibus Samariae: " Quid Iudaei faciunt imbecilles? Num hoc conceditur eis? Num, quia sacrificant, complebunt in una die? Numquid vivificare poterunt lapides de acervis pulveris, qui combusti sunt? ".
NEH|3|35|Sed et Thobias Ammanites, qui erat ad latus eius, ait: " Sine aedificare; si ascenderit vulpes, diruet murum eorum lapideum ".
NEH|3|36|Audi, Deus noster, quia facti sumus irrisio! Converte contumeliam eorum super caput eorum et da eos in irrisionem in terra captivitatis!
NEH|3|37|Ne operias iniquitatem eorum, et peccatum eorum coram facie tua non deleatur, quia offenderunt te coram aedificantibus.
NEH|3|38|Itaque aedificavimus murum, et compositus est totus murus usque ad partem dimidiam, et populus dabat cor suum, ut operaretur.
NEH|4|1|Factum est autem cum audisset Sanaballat et Thobias et Arabes et Ammanitae et Azotii quod prosperaretur restauratio muri Ierusalem et quod coepissent interrupta concludi, irati sunt nimis;
NEH|4|2|et conspiraverunt omnes pariter, ut venirent et pugnarent contra Ierusalem et facerent confusionem.
NEH|4|3|Et oravimus Deum nostrum et posuimus custodiam die ac nocte contra eos.
NEH|4|4|Dixit autem Iudas: " Debilitata est fortitudo portantis, et humus nimia est; et nos non poterimus aedificare murum ".
NEH|4|5|Et dixerunt hostes nostri: " Nesciant et ignorent, donec veniamus in medium eorum et interficiamus eos et cessare faciamus opus ".
NEH|4|6|Factum est autem venientibus Iudaeis, qui habitabant iuxta eos, et dicentibus nobis per decem vices ex omnibus locis, quibus venerant ad nos,
NEH|4|7|statuimus nos in inferioribus post murum in locis apertis, et ordinavi populum secundum familias cum gladiis suis et lanceis suis et arcubus suis.
NEH|4|8|Et perspexi atque surrexi, et aio ad optimates et magistratus et ad reliquam partem vulgi: " Nolite timere a facie eorum; Domini magni et terribilis mementote et pugnate pro fratribus vestris, filiis vestris et filiabus vestris et uxoribus vestris et domibus vestris ".
NEH|4|9|Factum est autem cum audissent inimici nostri nuntiatum esse nobis, dissipavit Deus consilium eorum, et reversi sumus omnes ad murum, unusquisque ad opus suum.
NEH|4|10|Et factum est a die illa, media pars iuvenum meorum faciebat opus, et media tenebat lanceas et scuta et arcus et loricas, et principes post omnem domum Iudae.
NEH|4|11|Aedificantium in muro et portantium onera et imponentium, una manu sua faciebat opus et altera tenebat gladium;
NEH|4|12|aedificantium enim unusquisque gladio erat accinctus renes, et sic aedificabant; et, qui clangebat bucina, iuxta me.
NEH|4|13|Et dixi ad optimates et ad magistratus et ad reliquam partem vulgi: " Opus grande est et latum, et nos separati sumus in muro procul alter ab altero;
NEH|4|14|in loco quocumque audieritis clangorem tubae, illuc concurrite ad nos. Deus noster pugnabit pro nobis ".
NEH|4|15|Et sic nos fecimus opus, et media pars nostrum tenebat lanceas ab ascensu aurorae, donec egrediantur astra.
NEH|4|16|In tempore quoque illo dixi populo: " Unusquisque cum puero suo pernoctet in medio Ierusalem; et erit nobis custodia per noctem, et opus per diem ".
NEH|4|17|Ego autem et fratres mei et pueri mei et custodes, qui erant post me, non deponebamus vestimenta nostra; unusquisque tenebat gladium in dextera sua.
NEH|5|1|Et factus est clamor populi et uxorum eius magnus adversus fratres suos Iudaeos.
NEH|5|2|Et erant qui dicerent: " Filios nostros et filias nostras pignoravimus, ut acciperemus frumentum et comederemus et viveremus! ".
NEH|5|3|Et erant qui dicerent: " Agros nostros et vineas et domos nostras opposuimus, ut acciperemus frumentum in fame! ".
NEH|5|4|Et alii dicebant: " Mutuo sumpsimus pecunias in tributa regis pro agris nostris et vineis nostris.
NEH|5|5|Et nunc sicut caro fratrum nostrorum sic caro nostra est, et sicut filii eorum ita et filii nostri; ecce nos subiugamus filios nostros et filias nostras in servitutem, et de filiabus nostris quaedam iam in servitute subiugatae sunt, nec habemus unde possint redimi, quia agros nostros et vineas nostras alii possident ".
NEH|5|6|Et iratus sum nimis, cum audissem clamorem eorum secundum verba haec.
NEH|5|7|Cogitavique in corde meo et increpavi optimates et magistratus et dixi eis: " Usuras singuli a fratribus vestris exigitis! ". Et congregavi adversum eos contionem magnam
NEH|5|8|et dixi eis: " Nos, ut scitis, redemimus fratres nostros Iudaeos, qui venditi fuerant gentibus, secundum possibilitatem nostram; quin potius et vos vendetis fratres vestros, ut vendentur nobis? ". Et siluerunt nec invenerunt quid responderent.
NEH|5|9|Dixique ad eos: " Non est bona res, quam facitis. Quare non in timore Dei nostri ambulatis, ne exprobretur nobis a gentibus inimicis nostris?
NEH|5|10|Et ego et fratres mei et pueri mei commodavimus plurimis pecuniam et frumentum; non repetamus usuras istas.
NEH|5|11|Reddite eis hodie agros suos et vineas suas et oliveta sua et domos suas et centesimam pecuniae frumenti vini et olei, quam exigere soletis ab eis ".
NEH|5|12|Et dixerunt: " Reddemus et ab eis nihil quaeremus; sicque faciemus, ut loqueris ". Et vocavi sacerdotes et feci eos iurare, ut facerent, sicut dictum erat.
NEH|5|13|Insuper excussi sinum meum et dixi: " Sic excutiat Deus omnem virum, qui non compleverit verbum istud, de domo sua et de laboribus suis; sic excutiatur et vacuus fiat! ". Et dixit universa multitudo: " Amen! ". Et laudaverunt Deum. Fecit ergo populus, sicut erat dictum.
NEH|5|14|A die autem illa, qua praeceperat rex mihi, ut essem dux in terra Iudae, ab anno vicesimo usque ad annum tricesimum secundum Artaxerxis regis, per annos duodecim ego et fratres mei annonas, quae ducibus debebantur, non comedimus.
NEH|5|15|Duces autem priores, qui fuerant ante me, gravaverunt populum et acceperunt ab eis cotidie pro pane siclos argenti quadraginta; sed et ministri eorum depresserunt populum. Ego autem non feci ita propter timorem Dei,
NEH|5|16|quin potius in opere muri restauravi et agrum non emi; et omnes pueri mei congregati ad opus erant.
NEH|5|17|Iudaei quoque et magistratus, centum quinquaginta viri, et qui veniebant ad nos de gentibus, quae in circuitu nostro sunt, in mensa mea erant.
NEH|5|18|Parabatur autem mihi per dies singulos bos unus, arietes sex electi, exceptis volatilibus; et inter dies decem vina diversa multa. Insuper et annonas ducatus mei non quaesivi; gravis enim erat servitus populi huius.
NEH|5|19|Memento mei, Deus meus, in bonum, secundum omnia, quae feci populo huic.
NEH|6|1|Factum est autem cum audisset Sanaballat et Thobias et Gosem Arabs et ceteri inimici nostri, quod aedificassem ego murum, et non esset in ipso residua interruptio - usque ad tempus autem illud valvas non posueram in portis -
NEH|6|2|miserunt Sanaballat et Gosem ad me dicentes: " Veni, et conveniamus in Cephirim in campo Ono ". Ipsi autem cogitabant, ut facerent mihi malum.
NEH|6|3|Misi ergo ad eos nuntios dicens: " Opus grande ego facio et non possum descendere; cur cessare oportet opus, si desistero et descendero ad vos?.
NEH|6|4|Miserunt autem ad me secundum verbum hoc per quattuor vices, et respondi eis iuxta sermonem priorem.
NEH|6|5|Et misit ad me Sanaballat iuxta verbum prius quinta vice puerum suum, et epistulam non obsignatam habebat in manu sua, in qua erat scriptum:
NEH|6|6|" In gentibus auditum est, et Gosem dixit quod tu et Iudaei cogitetis rebellare, et propterea aedifices murum et levare te velis super eos regem; iuxta hanc vocem
NEH|6|7|et prophetas posueris, qui praedicent de te in Ierusalem dicentes: "Rex in Iudaea est!". Nunc autem auditurus est rex verba haec; idcirco nunc veni, ut ineamus consilium pariter ".
NEH|6|8|Et misi ad eum dicens: " Non est factum secundum verba haec, quae tu loqueris; de corde enim tuo tu componis haec ".
NEH|6|9|Omnes enim hi terrebant nos cogitantes: " Fatigabuntur manus eorum ab opere, et non complebitur ". Quam ob causam magis confortavi manus meas.
NEH|6|10|Et ingressus sum domum Semeiae filii Dalaiae filii Meetabel, ubi erat detentus. Qui ait: " Tractemus nobiscum in domo Dei, in medio templi, et claudamus portas aedis, quia venturi sunt, ut interficiant te; utique nocte venturi sunt ad occidendum te".
NEH|6|11|Et dixi: " Num quisquam similis mei fugit? Et quis ut ego ingredietur templum et vivet? Non ingrediar ".
NEH|6|12|Et intellexi quod Deus non misisset eum, sed quasi vaticinans locutus esset ad me, quia Thobias et Sanaballat conduxerant eum.
NEH|6|13|Acceperat enim pretium, ut territus sic agerem et peccarem, et haberent malum, quod exprobrarent mihi.
NEH|6|14|Memento, Deus meus, Thobiae et Sanaballat iuxta opera eorum talia, sed et Noadiae prophetae et ceterorum prophetarum, qui terrebant me!
NEH|6|15|Completus est autem murus vicesimo quinto die mensis Elul, quinquaginta duobus diebus.
NEH|6|16|Factum est ergo, cum audissent omnes inimici nostri, et vidissent universae gentes, quae erant in circuitu nostro, ut conciderent intra semetipsos et scirent quod a Deo factum esset opus hoc.
NEH|6|17|Sed et in diebus illis, multae optimatum Iudaeorum epistulae mittebantur ad Thobiam, et a Thobia veniebant ad eos.
NEH|6|18|Multi enim in Iudaea coniurationem fecerunt cum eo, quia gener erat Secheniae filii Area, et Iohanan filius eius acceperat filiam Mosollam filii Barachiae.
NEH|6|19|Sed et laudabant eum coram me et verba mea nuntiabant ei; et Thobias mittebat epistulas, ut terreret me.
NEH|7|1|Postquam autem aedificatus est murus, et posui valvas et recen sui ianitores et cantores et Levitas,
NEH|7|2|praeposui Hanani fratrem meum et Hananiam principem arcis supra Ierusalem - ipse enim quasi vir verax et timens Deum plus ceteris videbatur -
NEH|7|3|et dixi eis: " Non aperiantur portae Ierusalem usque ad calorem solis. Dum adhuc calor permanet, claudantur portae et oppilentur; et ponant custodes de habitatoribus Ierusalem, singulos per vices suas et unumquemque contra domum suam ".
NEH|7|4|Civitas autem erat lata nimis et grandis, et populus parvus in medio eius, et non erant domus aedificatae.
NEH|7|5|Deus autem meus dedit in corde meo, et congregavi optimates et magistratus et vulgus, ut recenserem eos; et inveni librum census eorum, qui ascenderant primum, et inventum est scriptum in eo:
NEH|7|6|Isti filii provinciae, qui ascenderunt de captivitate migrantium, quos transtulerat Nabuchodonosor rex Babylonis, et reversi sunt in Ierusalem et in Iudaeam unusquisque in civitatem suam.
NEH|7|7|Qui venerunt cum Zorobabel, Iesua, Nehemias, Azarias, Raamias, Nahamani, Mardochaeus, Belsan, Mespharath, Beguai, Nahum, Baana.Numerus virorum populi Israel:
NEH|7|8|filii Pharos duo milia centum septuaginta duo;
NEH|7|9|filii Saphatia trecenti septuaginta duo;
NEH|7|10|filii Area sescenti quinquaginta duo;
NEH|7|11|filii Phahathmoab, hi sunt filii Iesua et Ioab, duo milia octingenti decem et octo;
NEH|7|12|filii Elam mille ducenti quinquaginta quattuor;
NEH|7|13|filii Zethua octingenti quadraginta quinque;
NEH|7|14|filii Zachai septingenti sexaginta;
NEH|7|15|filii Bennui sescenti quadraginta octo;
NEH|7|16|filii Bebai sescenti viginti octo;
NEH|7|17|filii Azgad duo milia trecenti viginti duo;
NEH|7|18|filii Adonicam sescenti sexaginta septem;
NEH|7|19|filii Beguai duo milia sexaginta septem;
NEH|7|20|filii Adin sescenti quinquaginta quinque;
NEH|7|21|filii Ater, qui erant ex Ezechia, nonaginta octo;
NEH|7|22|filii Hasum trecenti viginti octo;
NEH|7|23|filii Besai trecenti viginti quattuor;
NEH|7|24|filii Hareph centum duodecim;
NEH|7|25|filii Gabaon nonaginta quinque;
NEH|7|26|filii Bethlehem et Netopha centum octoginta octo;
NEH|7|27|viri Anathoth centum viginti octo;
NEH|7|28|viri Bethazmaveth quadraginta duo;
NEH|7|29|viri Cariathiarim, Cephira et Beroth septingenti quadraginta tres;
NEH|7|30|viri Rama et Gabaa sescenti viginti unus;
NEH|7|31|viri Machmas centum viginti duo;
NEH|7|32|viri Bethel et Hai centum viginti tres;
NEH|7|33|viri Nabo alterius quinquaginta duo;
NEH|7|34|viri Elam alterius mille ducenti quinquaginta quattuor;
NEH|7|35|filii Harim trecenti viginti;
NEH|7|36|filii Iericho trecenti quadraginta quinque;
NEH|7|37|filii Lod, Hadid et Ono septingenti viginti unus;
NEH|7|38|filii Senaa tria milia nongenti triginta.
NEH|7|39|Sacerdotes: filii Iedaia de domo Iesua nongenti septuaginta tres;
NEH|7|40|filii Emmer mille quinquaginta duo;
NEH|7|41|filii Phassur mille ducenti quadraginta septem;
NEH|7|42|filii Harim mille decem et septem.
NEH|7|43|Levitae: filii Iesua, hi sunt filii Cadmihel, Bennui et Odoviae, septuaginta quattuor.
NEH|7|44|Cantores: filii Asaph centum quadraginta octo.
NEH|7|45|Ianitores: filii Sellum, filii Ater, filii Telmon, filii Accub, filii Hatita, filii Sobai, centum triginta octo.
NEH|7|46|Oblati: filii Siha, filii Hasupha, filii Tabbaoth,
NEH|7|47|filii Ceros, filii Siaa, filii Phadon,
NEH|7|48|filii Lebana, filii Hagaba, filii Selmai,
NEH|7|49|filii Hanan, filii Giddel, filii Gaher,
NEH|7|50|filii Raaia, filii Rasin, filii Necoda,
NEH|7|51|filii Gazam, filii Oza, filii Phasea,
NEH|7|52|filii Besai, filii Meunitarum, filii Nephusorum,
NEH|7|53|filii Bacbuc, filii Hacupha, filii Harhur,
NEH|7|54|filii Basluth, filii Mahida, filii Harsa,
NEH|7|55|filii Bercos, filii Sisara, filii Thema,
NEH|7|56|filii Nasia, filii Hatipha.
NEH|7|57|Filii servorum Salomonis: filii Sotai, filii Sophereth, filii Pheruda,
NEH|7|58|filii Iaala, filii Darcon, filii Giddel,
NEH|7|59|filii Saphatia, filii Hatil, filii Phochereth Hassebaim, filii Amon.
NEH|7|60|Omnes oblati et filii servorum Salomonis trecenti nonaginta duo.
NEH|7|61|Hi sunt autem, qui ascenderunt de Thelmela, Thelharsa, Cherub, Addon et Emmer et non potuerunt indicare domum patrum suorum et semen suum, utrum ex Israel essent:
NEH|7|62|filii Dalaia, filii Thobia, filii Necoda sescenti quadraginta duo.
NEH|7|63|Et de sacerdotibus: filii Hobia, filii Accos, filii Berzellai, qui accepit de filiabus Berzellai Galaaditis uxorem et vocatus est nomine eorum.
NEH|7|64|Hi quaesierunt tabulas genealogiae suae et non invenerunt; et eiecti sunt de sacerdotio;
NEH|7|65|dixitque praepositus eis, ut non manducarent de sanctificatis sanctuarii, donec staret sacerdos pro Urim et Tummim.
NEH|7|66|Omnis multitudo simul quadraginta duo milia trecenti sexaginta,
NEH|7|67|absque servis et ancillis eorum, qui erant septem milia trecenti triginta septem; insuper et cantores et cantatrices ducenti quadraginta quinque.
NEH|7|68|Equi eorum septingenti triginta sex, muli eorum ducenti quadraginta quinque,
NEH|7|69|cameli eorum quadringenti triginta quinque, asini sex milia septingenti viginti.
NEH|7|70|Nonnulli autem de principibus familiarum dederunt in opus: praepositus dedit in thesaurum auri drachmas mille, phialas quinquaginta, tunicas sacerdotales quingentas triginta;
NEH|7|71|et de principibus familiarum dederunt in thesaurum operis auri drachmas viginti milia et argenti minas duo milia ducentas.
NEH|7|72|Et quod dedit reliquus populus, auri drachmas viginti milia et argenti minas duo milia et tunicas sacerdotales sexaginta septem. Habitaverunt autem ibi sacerdotes et Levitae; ianitores autem et cantores et quidam de populo et oblati et omnis Israel habitaverunt in civitatibus suis.Et venerat mensis septimus; filii autem Israel erant in civitatibus suis.
NEH|8|1|Congregatusque est omnis populus quasi vir unus ad plateam, quae est ante portam Aquarum, et dixerunt Esdrae scribae, ut afferret librum legis Moysi, quam praece perat Dominus Israeli.
NEH|8|2|Attulit ergo Esdras sacerdos legem coram multitudine virorum et mulierum cunctisque, qui poterant intellegere, in die prima mensis septimi.
NEH|8|3|Et legit in eo in platea, quae erat ante portam Aquarum, de mane usque ad mediam diem in conspectu virorum et mulierum et eorum, qui intellegere poterant; et aures omnis populi erant erectae ad librum legis.
NEH|8|4|Stetit autem Esdras scriba super gradum ligneum, quem ad hoc fecerant; et steterunt iuxta eum Matthathias et Sema et Anaia et Uria et Helcia et Maasia ad dexteram eius, et ad sinistram Phadaia, Misael et Melchia et Hasum et Hasbadana, Zacharia et Mosollam.
NEH|8|5|Et aperuit Esdras librum coram omni populo - super universum quippe populum eminebat - et, cum aperuisset eum, stetit omnis populus.
NEH|8|6|Et benedixit Esdras Domino, Deo magno; et respondit omnis populus: " Amen, amen ", elevans manus suas. Et incurvati sunt et adoraverunt Deum proni in terram.
NEH|8|7|Porro Iesua et Bani et Serebia, Iamin, Accub, Sabethai, Hodia, Maasia, Celita, Azarias, Iozabad, Hanan, Phalaia et Levitae erudiebant populum in lege; populus autem stabat in gradu suo.
NEH|8|8|Et legerunt in libro legis Dei distincte et aperierunt sensum et explicaverunt lectionem.
NEH|8|9|Dixit autem Nehemias, ipse est praepositus, et Esdras sacerdos et scriba et Levitae instruentes populum universo populo: " Dies iste sanctificatus est Domino Deo nostro! Nolite lugere et nolite flere ". Flebat enim omnis populus, cum audiret verba legis.
NEH|8|10|Et dixit eis: " Ite, comedite pinguia et bibite mulsum et mittite partes his, qui non praeparaverunt sibi, quia sanctus dies Domini nostri est; et nolite contristari, gaudium etenim Domini est fortitudo vestra ".
NEH|8|11|Levitae autem silentium faciebant in omni populo dicentes: " Tacete, quia dies sanctus est, et nolite dolere ".
NEH|8|12|Abiit itaque omnis populus, ut comederet et biberet et mitteret partes et faceret laetitiam magnam, quia intellexerant verba, quae docuerat eos.
NEH|8|13|Et in die secundo congregati sunt principes familiarum universi populi, sacerdotes et Levitae ad Esdram scribam, ut intellegerent verba legis.
NEH|8|14|Et invenerunt scriptum in lege, quam praecepit Dominus per Moysen, ut habitent filii Israel in tabernaculis in die sollemni mense septimo
NEH|8|15|et ut praedicent et divulgent vocem in universis urbibus suis et in Ierusalem dicentes: " Egredimini in montem et afferte frondes olivae et frondes oleastri, frondes myrti et ramos palmarum et frondes ligni nemorosi, ut fiant tabernacula, sicut scriptum est ".
NEH|8|16|Et egressus est populus, et attulerunt feceruntque sibi tabernacula, unusquisque in domate suo et in atriis suis et in atriis domus Dei et in platea portae Aquarum et in platea portae Ephraim.
NEH|8|17|Fecit ergo universa ecclesia eorum, qui redierant de captivitate, tabernacula et habitaverunt in tabernaculis. Non enim fecerant a diebus Iosue filii Nun taliter filii Israel usque ad diem illum; et fuit laetitia magna nimis.
NEH|8|18|Legit autem in libro legis Dei per dies singulos, a die primo usque ad diem novissimum; et fecerunt sollemnitatem septem diebus et in die octavo conventum iuxta ordinationem.
NEH|9|1|In die autem vicesimo quarto mensis huius convenerunt filii Is rael in ieiunio et in saccis, et humus super eos.
NEH|9|2|Et separatum est semen filiorum Israel ab omni alienigena; et steterunt et confitebantur peccata sua et iniquitates patrum suorum.
NEH|9|3|Et consurrexerunt ad standum et legerunt in volumine legis Domini Dei sui per quartam partem diei; et per quartam partem confitebantur et adorabant Dominum Deum suum.
NEH|9|4|Surrexerunt autem super gradum Levitarum Iesua et Bani et Cadmihel, Sebania, Bunni, Serebia, Bani et Chanani et clamaverunt voce magna ad Dominum Deum suum.
NEH|9|5|Et dixerunt Levitae Iesua et Cadmihel, Bani, Hasabneia, Serebia, Hodia, Sebania, Phethahia: Surgite, benedicite Domino Deo vestroab aetemo usque in aeternum,et benedicant nomini gloriae tuae excelsosuper omnem benedictionem et laudem.
NEH|9|6|Tu ipse, Domine, solus;tu fecisti caelum et caelum caelorumet omnem exercitum eorum,terram et universa, quae in ea sunt, maria et omnia, quae in eis sunt;et tu vivificas omnia haec,et exercitus caeli te adorat.
NEH|9|7|Tu ipse, Domine Deus, qui elegisti Abramet eduxisti eum de Ur Chaldaeorumet posuisti nomen eius Abraham.
NEH|9|8|Et invenisti cor eius fidele coram teet percussisti cum eo foedus,ut dares terram Chananaei, Hetthaei et Amorraeiet Pherezaei et Iebusaei et Gergesaei,nempe ut dares semini eius;et implesti verba tua,quoniam iustus es.
NEH|9|9|Et vidisti afflictionem patrum nostrorum in Aegyptoclamoremque eorum audisti iuxta mare Rubrum.
NEH|9|10|Et dedisti signa atque portenta in pharaoneet in universis servis eius et in omni populo terrae illius;cognovisti enim quia superbe egerant contra eos,et fecisti tibi nomen, sicut et in hac die.
NEH|9|11|Et mare divisisti ante eos,et transierunt per medium maris in sicco;persecutores autem eorum proiecisti in profundum,quasi lapidem in aquas validas.
NEH|9|12|Et in columna nubis ductor eorum fuisti per diemet in columna ignis per noctem,ut illuminaret eis viam, per quam ingrediebantur.
NEH|9|13|Ad montem quoque Sinai descendistiet locutus es cum eis de caelo;et dedisti eis iudicia rectaet legem rectam, mandata et praecepta bona.
NEH|9|14|Et sabbatum sanctificatum tuum ostendisti eiset praecepta et mandata et legem praecepisti eisin manu Moysi servi tui.
NEH|9|15|Panem quoque de caelo dedisti eis in fame eorumet aquam de petra eduxisti eis in siti eorum;et dixisti eis, ut ingrederentur et possiderent terram,super quam levasti manum tuam, ut traderes eis.
NEH|9|16|Ipsi vero patres nostri superbe egeruntet induraverunt cervices suas et non audierunt mandata tua.
NEH|9|17|Et noluerunt audireet non sunt recordati mirabilium tuorum, quae feceras eis,et induraverunt cervices suaset posuerunt caput suum,ut reverterentur ad servitutem suam in Aegyptum.Tu autem Deus propitius, clemens et misericors,longanimis et multae miserationis, non dereliquisti eos.
NEH|9|18|Et quidem, cum fecissent sibi vitulum conflatilemet dixissent: "Iste est Deus tuus,qui eduxit te de Aegypto"feceruntque blasphemias magnas;
NEH|9|19|tu autem in misericordiis tuis multisnon dimisisti eos in deserto:columna nubis non recessit ab eis per diem,ut duceret eos in viam;et columna ignis per noctem,ut illuminaret eis iter, per quod ingrederentur.
NEH|9|20|Et spiritum tuum bonum dedisti, qui doceret eos,et manna tuum non prohibuisti ab ore eorumet aquam dedisti eis in siti eorum.
NEH|9|21|Quadraginta annis pavisti eos in deserto,nihilque eis defuit;vestimenta eorum non inveteraverunt,et pedes eorum non intumuerunt.
NEH|9|22|Et dedisti eis regna et populoset partitus es eis sortes;et possederunt terram Sehon et terram regis Hesebonet terram Og regis Basan.
NEH|9|23|Et multiplicasti filios eorum sicut stellas caeli;et adduxisti eos ad terram, de qua dixeras patribus eorum,ut ingrederentur et possiderent.
NEH|9|24|Et venerunt filii et possederunt terram,et humiliasti coram eis habitatores terrae Chananaeos;et dedisti eos in manu eorumet reges eorum et populos terrae,ut facerent eis, sicut placebat illis.
NEH|9|25|Ceperunt itaque urbes munitas et humum pinguem;et possederunt domos plenas cunctis bonis,cisternas ab aliis fabricatas, vineas et olivetaet ligna pomifera multa.Et comederunt et saturati sunt et impinguati suntet delectati sunt in bonitate tua magna.
NEH|9|26|Vexaverunt autem te et rebellaverunt contra teet proiecerunt legem tuam post terga sua;et prophetas tuos occiderunt,qui contestabantur eos, ut reverterentur ad te;feceruntque blasphemias grandes.
NEH|9|27|Et dedisti eos in manu hostium suorum,et afflixerunt eos;et in tempore tribulationis suae clamaverunt ad te,et tu de caelo audistiet secundum miserationes tuas multas dedisti eis salvatores,qui salvarent eos da manu hostium suorum.
NEH|9|28|Cumque requievissent, reversi sunt,ut facerent malum in conspectu tuo;et dereliquisti eos in manu inimicorum suorum,et dominati sunt eis.Conversique sunt et clamaverunt ad te;tu autem de caelo exaudistiet liberasti eos in misericordiis tuis multis vicibus.
NEH|9|29|Et contestatus es eos, ut reduceres eos ad legem tuam;ipsi vero superbe egerunt et non audierunt mandata tuaet in iudicia tua peccaverunt, quae si fecerit homo, vivet in eis, et dederunt umerum rebellemet cervicem suam induraverunt nec audierunt.
NEH|9|30|Et pepercisti eis annos multoset contestatus es eos in spiritu tuoper manum prophetarum tuorum, et non audierunt;et tradidisti eos in manu populorum terrarum.
NEH|9|31|In misericordiis autem tuis plurimisnon fecisti eos in consumptionemnec dereliquisti eos;quoniam Deus misericors et clemens es tu.
NEH|9|32|Nunc itaque, Deus noster magne, fortis et terribilis,custodiens pactum et misericordiam,ne parvipendas omnem laborem,qui invenit nos, reges nostros et principes nostroset sacerdotes nostros et prophetas nostroset patres nostros et omnem populum tuuma diebus regum Assyriae usque in diem hanc.
NEH|9|33|Et tu iustus es in omnibus, quae venerunt super nos,quia recte fecisti,nos autem impie egimus.
NEH|9|34|Reges nostri, principes nostri, sacerdotes nostri et patres nostrinon fecerunt legem tuamet non attenderunt mandata tua et testimonia tua,quae testificatus es in eis.
NEH|9|35|Et ipsi in regnis suis et in bonitate tua multa, quam dederas eis,et in terra latissima et pingui,quam tradideras in conspectu eorum,non servierunt tibi nec reversi sunt a studiis suis pessimis.
NEH|9|36|Ecce nos ipsi hodie servi sumus;et in terra, quam dedisti patribus nostris,ut comederent fructum eius et bona eius, nos ipsi servi sumus.
NEH|9|37|Et fruges eius multiplicantur regibus,quos posuisti super nos propter peccata nostra,et corporibus nostris dominantur et iumentis nostrissecundum voluntatem suam,et in tribulatione magna sumus ".
NEH|10|1|" Super omnibus ergo his nos ipsi percutimus foedus et scribimus, et signant principes nostri, Levitae nostri et sacerdotes nostri ".
NEH|10|2|Signatores autem fuerunt: Nehemias praepositus, filius Hachaliae, et Sedecias,
NEH|10|3|Saraias, Azarias, Ieremias,
NEH|10|4|Phassur, Amarias, Melchias,
NEH|10|5|Hattus, Sebania, Melluch,
NEH|10|6|Harim, Meremoth, Abdias,
NEH|10|7|Daniel, Genthon, Baruch,
NEH|10|8|Mosollam, Abia, Miamin,
NEH|10|9|Maazia, Belgai, Semeia; hi sacerdotes.
NEH|10|10|Porro Levitae: Iesua filius Azaniae, Bennui de filiis Henadad, Cadmihel
NEH|10|11|et fratres eorum Sebania, Hodia, Celita, Phalaia, Hanan,
NEH|10|12|Micha, Rohob, Hasabia,
NEH|10|13|Zacchur, Serebia, Sebania,
NEH|10|14|Hodia, Bani, Baninu.
NEH|10|15|Capita populi: Pharos, Phahathmoab, Elam, Zethua, Bani,
NEH|10|16|Bunni, Azgad, Bebai,
NEH|10|17|Adonia, Beguai, Adin,
NEH|10|18|Ater, Ezechia, Azur,
NEH|10|19|Hodia, Hasum, Besai,
NEH|10|20|Hareph, Anathoth, Nebai,
NEH|10|21|Megphias, Mosollam, Hezir,
NEH|10|22|Mesezabel, Sadoc, Ieddua,
NEH|10|23|Pheltia, Hanan, Anaia,
NEH|10|24|Osee, Hanania, Hassub,
NEH|10|25|Alohes, Phalea, Sobec,
NEH|10|26|Rehum, Hasabna, Maasia,
NEH|10|27|Ahia, Hanan, Anan,
NEH|10|28|Melluch, Harim, Baana.
NEH|10|29|Et reliqui de populo, sacerdotes, Levitae, ianitores et cantores, oblati et omnes, qui se separaverunt de populis terrarum ad legem Dei, uxores eorum, filii eorum et filiae eorum, omnes, qui poterant sapere,
NEH|10|30|adhaeserunt fratribus suis optimatibus pollicentes et iurantes, ut ambularent in lege Dei, quam dederat in manu Moysi servi Dei, et ut facerent et custodirent universa mandata Domini Dei nostri et iudicia eius et praecepta eius,
NEH|10|31|et ut non daremus filias nostras populo terrae et filias eorum non acciperemus filiis nostris.
NEH|10|32|Et si populi terrae importaverint venalia et omnia cibaria per diem sabbati, ut vendant, non accipiemus ab eis in sabbato et in die sanctificato; et dimittemus annum septimum et omnem exactionem.
NEH|10|33|Et statuimus super nos praecepta, ut demus tertiam partem sicli per annum ad opus domus Dei nostri,
NEH|10|34|ad panes propositionis et ad oblationem sempiternam et in holocaustum sempiternum in sabbatis, in calendis, in sollemnitatibus et in sanctificata et in sacrificium pro peccato, ut expietur pro Israel, et in omnem usum domus Dei nostri.
NEH|10|35|Sortes ergo misimus super oblationem lignorum inter sacerdotes et Levitas et populum, ut inferrentur in domum Dei nostri per domos patrum nostrorum, in temporibus constitutis ab anno in annum, ut arderent super altare domini Dei nostri, sicut scriptum est in lege;
NEH|10|36|et ut afferremus primogenita terrae nostrae et primitiva universi fructus omnis ligni ab anno in annum in domo Domini,
NEH|10|37|et primitiva filiorum nostrorum et pecorum nostrorum, sicut scriptum est in lege, et primitiva boum nostrorum et ovium nostrarum, ut afferrentur in domum Dei nostri sacerdotibus, qui ministrant in domo Dei nostri;
NEH|10|38|et primitias ciborum nostrorum et libaminum nostrorum et poma omnis ligni, vindemiae quoque et olei, afferemus sacerdotibus ad gazophylacium Dei nostri, et decimam partem terrae nostrae Levitis. Ipsi Levitae decimas accipient ex omnibus civitatibus agriculturae nostrae.
NEH|10|39|Erit autem sacerdos filius Aaron cum Levitis in decimis Levitarum colligendis, et Levitae offerent decimam partem decimae in domo Dei nostri ad gazophylacium thesauri.
NEH|10|40|Ad gazophylacium enim deportabunt filii Israel et filii Levi primitias frumenti, vini et olei; et ibi erunt vasa sanctificata et sacerdotes, qui ministrabant, et ianitores et cantores. Et non dimittemus domum Dei nostri.
NEH|11|1|Habitaverunt autem princi pes populi in Ierusalem; reli qua vero plebs misit sortem, ut adducerent unum virum de decem ad habitandum in Ierusalem civitate sancta, novem vero partes in civitatibus.
NEH|11|2|Benedixit autem populus omnibus viris, qui se sponte obtulerant, ut habitarent in Ierusalem.
NEH|11|3|Hi sunt itaque principes provinciae, qui habitaverunt in Ierusalem et in civitatibus Iudae. Habitavit autem unusquisque in possessione sua, in urbibus suis, Israel, sacerdotes, Levitae, oblati et filii servorum Salomonis.
NEH|11|4|Et in Ierusalem habitaverunt de filiis Iudae et de filiis Beniamin. De filiis Iudae: Athaias filius Oziam filii Zachariae filii Amariae filii Saphatiae filii Malaleel, de filiis Phares;
NEH|11|5|et Maasia filius Baruch filius Cholhoza filius Hazia filius Adaia filius Ioiarib filius Zachariae filius Silonitis.
NEH|11|6|Omnes filii Phares, qui habitaverunt in Ierusalem, quadringenti sexaginta octo viri fortes.
NEH|11|7|Hi sunt autem filii Beniamin: Sallu filius Mosollam filius Ioed filius Phadaia filius Colaia filius Maasia filius Etheel filius Iesaia;
NEH|11|8|et fratres eius viri fortes, nongenti viginti octo.
NEH|11|9|Et Ioel filius Zechri praepositus eorum, et Iudas filius Asana super civitatem secundus.
NEH|11|10|Et de sacerdotibus: Iedaia filius Ioiarib filius
NEH|11|11|Saraia filius Helciae filius Mosollam filius Sadoc filius Meraioth filius Achitob princeps domus Dei;
NEH|11|12|et fratres eorum facientes opera templi, octingenti viginti duo. Et Adaia filius Ieroham filius Phelelia filius Amsi filius Zachariae filius Phassur filius Melchiae;
NEH|11|13|et fratres eius principes familiarum ducenti quadraginta duo. Et Amassai filius Azareel filius Ahazi filius Mosollamoth filius Emmer;
NEH|11|14|et fratres eorum potentes nimis, centum viginti octo; et praepositus eorum Zabdiel vir nobilis.
NEH|11|15|Et de Levitis: Semeia filius Hassub filius Ezricam filius Hasabia filius Bunni;
NEH|11|16|et Sabethai et Iozabad super omnia opera, quae erant forinsecus in domo Dei, de principibus Levitarum;
NEH|11|17|et Matthania filius Micha filius Zebedaei filius Asaph magister chori incohabat orationem; et Becbecia secundus de fratribus eius, et Abda filius Sammua filius Galal filius Idithun.
NEH|11|18|Omnes Levitae in civitate sancta ducenti octoginta quattuor.
NEH|11|19|Et ianitores: Accub, Telmon et fratres eorum, qui custodiebant ostia, centum septuaginta duo.
NEH|11|20|Et reliqui ex Israel sacerdotes et Levitae in universis civitatibus Iudae, unusquisque in possessione sua.
NEH|11|21|Et oblati habitabant in Ophel; et Siha et Gaspha super oblatos.
NEH|11|22|Et praefectus Levitarum in Ierusalem Ozi filius Bani filius Hasabiae filius Matthaniae filius Michae de filiis Asaph, cantores in ministerio domus Dei.
NEH|11|23|Praeceptum quippe regis super eos erat, et ordo in cantoribus per dies singulos.
NEH|11|24|Et Phethahia filius Mesezabel de filiis Zara filii Iudae, legatus regis in omni negotio populi.
NEH|11|25|Et in viculis per omnes regiones eorum, de filiis Iudae habitaverunt in Cariatharbe et in pagis eius et in Dibon et in pagis eius et in Cabseel et in viculis eius
NEH|11|26|et in Iesua et in Molada et in Bethpheleth
NEH|11|27|et in Asarsual et in Bersabee et in pagis eius
NEH|11|28|et in Siceleg et in Mochona et in pagis eius
NEH|11|29|et in Remmon et in Saraa et in Ierimoth,
NEH|11|30|Zanoa, Odollam et in villis earum, Lachis et regionibus eius et Azeca et pagis eius. Et habitaverunt a Bersabee usque ad vallem Ennom.
NEH|11|31|Filii autem Beniamin in Gabaa, Machmas et Hai et Bethel et pagis eius,
NEH|11|32|Anathoth, Nob, Anania,
NEH|11|33|Asor, Rama, Getthaim,
NEH|11|34|Hadid, Seboim et Neballat,
NEH|11|35|Lod et Ono et valle Artificum.
NEH|11|36|Et de Levitis portiones in Iuda et Beniamin.
NEH|12|1|Hi sunt autem sacerdotes et Levitae, qui ascenderunt cum Zorobabel filio Salathiel et Iesua: Saraia, Ieremias, Esdras,
NEH|12|2|Amaria, Melluch, Hattus,
NEH|12|3|Sechenias, Rehum, Meremoth,
NEH|12|4|Addo, Genthon, Abia,
NEH|12|5|Miamin, Maadia, Belga,
NEH|12|6|Semeia et Ioiarib, Iedaia,
NEH|12|7|Sallu, Amoc, Helcias, Iedaia. Isti principes sacerdotum et fratrum eorum in diebus Iesua.
NEH|12|8|Porro Levitae: Iesua, Bennui, Cadmihel, Serebia, Iuda, Matthanias, super hymnos ipse et fratres eius;
NEH|12|9|et Becbecia atque Hanni fratres eorum coram eis per vices suas.
NEH|12|10|Iesua autem genuit Ioachim, et Ioachim genuit Eliasib, et Eliasib genuit Ioiada,
NEH|12|11|et Ioiada genuit Ionathan, et Ionathan genuit Ieddua.
NEH|12|12|In diebus autem Ioachim erant sacerdotes principes familiarum: Saraiae Maraia, Ieremiae Hanania,
NEH|12|13|Esdrae Mosollam, Amariae Iohanan,
NEH|12|14|Milicho Ionathan, Sebaniae Ioseph,
NEH|12|15|Harim Edna, Meraioth Helci,
NEH|12|16|Adaiae Zacharia, Genthon Mosollam,
NEH|12|17|Abiae Zechri, Miamin Maadiae Phelti,
NEH|12|18|Belgae Sammua, Semeiae Ionathan,
NEH|12|19|Ioiarib Matthanai, Iedaiae Ozi,
NEH|12|20|Sellai Celai, Amoc Heber,
NEH|12|21|Helciae Hasabia, Iedaiae Nathanael.
NEH|12|22|Levitae in diebus Eliasib et Ioiada et Iohanan et Ieddua scripti principes familiarum et sacerdotes usque ad regnurn Darii Persae.
NEH|12|23|Filii Levi principes familiarum scripti in libro Chronicorum usque ad dies Ionathan filii Eliasib.
NEH|12|24|Et principes Levitarum Hasabia, Serebia, Iesua, Bennui et Cadmihel et fratres eorum coram eis, ut laudarent et confiterentur iuxta praeceptum David viri Dei per vices suas;
NEH|12|25|Matthania et Becbecia, Abdia, Mosollam, Telmon, Accub ianitores ad custodiam horreorum iuxta portas.
NEH|12|26|Hi in diebus Ioachim filii Iesua filii Iosedec et in diebus Nehemiae ducis et Esdrae sacerdotis scribaeque.
NEH|12|27|In dedicatione autem muri Ierusalem requisierunt Levitas de omnibus locis suis, ut adducerent eos in Ierusalem et facerent dedicationem in laetitia, in actione gratiarum et cantico et cymbalis, psalteriis et citharis.
NEH|12|28|Congregati sunt autem cantores de campestribus circa Ierusalem et de villis Netophathitarum
NEH|12|29|et de Bethgalgala et de regionibus Gabaa et Azmaveth, quoniam villas aedificaverunt sibi cantores in circuitu Ierusalem.
NEH|12|30|Et mundati sunt sacerdotes et Levitae et mundaverunt populum et portas et murum.
NEH|12|31|Ascendere autem feci principes Iudae super murum et statui duos magnos choros laudantium, quorum unus ivit ad dexteram super murum ad portam Sterquilinii.
NEH|12|32|Et ivit post eos Osaias et media pars principum Iudae
NEH|12|33|et Azarias, Esdras et Mosollam,
NEH|12|34|Iudas et Beniamin et Semeia et Ieremias.
NEH|12|35|Et de sacerdotibus cum tubis et Zacharias filius Ionathan filius Semeiae filius Matthaniae filius Michaiae filius Zacchur filius Asaph;
NEH|12|36|et fratres eius Semeia et Azareel, Malalai, Galalai, Maai, Nathanael et Iudas et Hanani cum musicis David viri Dei; et Esdras scriba ante eos et in porta Fontis.
NEH|12|37|Processerunt per gradus civitatis David in ascensu muri super domum David et usque ad portam Aquarum ad orientem.
NEH|12|38|Et chorus secundus gratias referentium ibat ex adverso, et ego post eum, et media pars populi super murum et super turrim Furnorum et usque ad murum latissimum
NEH|12|39|et super portam Ephraim et super portam Antiquam et super portam Piscium et turrim Hananeel et turrim Meah et usque ad portam Gregis; et steterunt in porta Custodiae.
NEH|12|40|Steteruntque duo chori laudantium in domo Dei, et ego et dimidia pars magistratuum mecum.
NEH|12|41|Et sacerdotes Eliachim, Maasia, Miamin, Michaia, Elioenai, Zacharia, Hanania in tubis;
NEH|12|42|et Maasia et Semeia et Eleazar et Ozi et Iohanan et Melchia et Elam et Ezer. Et clare cecinerunt cantores et Izrahia praepositus.
NEH|12|43|Et obtulerunt in die illa sacrificia magna et laetati sunt; Deus enim laetificaverat eos laetitia magna; sed et uxores eorum et liberi gavisi sunt, et audita est laetitia Ierusalem procul.
NEH|12|44|Praeposuerunt quoque in die illa viros super gazophylacia ad thesaurum, ad libamina et ad primitias et ad decimas, ut colligerent in ea de agris civitatum partes legitimas pro sacerdotibus et Levitis; quia laetificatus est Iuda in sacerdotibus et Levitis, qui adstiterunt
NEH|12|45|et servierunt in ministerio Dei sui et in ministerio purificationis simul cum cantoribus et ianitoribus iuxta praeceptum David et Salomonis filii eius;
NEH|12|46|quia in diebus David et Asaph ab exordio erant catervae cantorum et carmina laudis et actionis gratiarum Deo.
NEH|12|47|Et omnis Israel in diebus Zorobabel et in diebus Nehemiae dabant partes cantoribus et ianitoribus per dies singulos partem suam et partes consecrabant Levitis, et Levitae consecrabant filiis Aaron.
NEH|13|1|In die autem illo lectum est in volumine Moysi, audiente populo, et inventum est scriptum in eo quod non debeant introire Ammonites et Moabites in ecclesiam Dei usque in aeternum,
NEH|13|2|eo quod non occurrerint filiis Israel cum pane et aqua et conduxerint adversum eos Balaam ad maledicendum eis, et convertit Deus noster maledictionem in benedictionem.
NEH|13|3|Factum est autem, cum audissent legem, separaverunt omnem promiscuum ab Israel.
NEH|13|4|Ante hoc autem erat Eliasib sacerdos, qui fuerat praepositus in gazophylacio domus Dei nostri et proximus Thobiae;
NEH|13|5|fecerat ei gazophylacium grande, ubi antea reponebant munera et tus et vasa et decimam frumenti, vini et olei, partes Levitarum et cantorum et ianitorum et tributa sacerdotum.
NEH|13|6|In omnibus autem his non fui in Ierusalem, quia anno tricesimo secundo Artaxerxis regis Babylonis veni ad regem et in fine dierum rogavi, ut abirem a rege,
NEH|13|7|et veni in Ierusalem. Et intellexi malum, quod fecerat Eliasib Thobiae: fecerat enim ei thesaurum in vestibulis domus Dei.
NEH|13|8|Et malum mihi visum est valde, et proieci vasa domus Thobiae foras de gazophylacio;
NEH|13|9|praecepique, et emundaverunt gazophylacia, et rettuli ibi vasa domus Dei, oblationem et tus.
NEH|13|10|Et cognovi quod partes Levitarum non fuissent datae, et fugisset unusquisque in campum suum de Levitis et cantoribus, qui ministrabant.
NEH|13|11|Et egi causam adversus magistratus et dixi: " Quare dereliquimus domum Dei? ". Et congregavi eos et feci stare in stationibus suis.
NEH|13|12|Et omnis Iuda apportabat decimam frumenti, vini et olei in horrea.
NEH|13|13|Et constitui super horrea Selemiam sacerdotem et Sadoc scribam et Phadaiam de Levitis et iuxta eos Hanan filium Zacchur, filium Matthaniae, quoniam fideles comprobati sunt; et ipsi curam habebant distribuendi partes fratribus suis.
NEH|13|14|Memento mei, Deus meus, pro hoc; et ne deleas opera mea bona, quae feci in domo Dei mei et in ministeriis eius!
NEH|13|15|In diebus illis vidi in Iuda calcantes torcularia in sabbato, portantes acervos et onerantes super asinos vinum et uvas et ficus et omne onus et inferentes in Ierusalem die sabbati; et contestatus sum, quando vendebant cibaria.
NEH|13|16|Et ibi Tyrii habitaverunt in ea inferentes pisces et omnia venalia et vendebant in sabbatis filiis Iudae in Ierusalem.
NEH|13|17|Et obiurgavi optimates Iudae et dixi eis: " Quae est haec res mala, quam vos facitis, et profanatis diem sabbati?
NEH|13|18|Numquid non haec fecerunt patres nostri, et adduxit Deus noster super nos omne malum hoc et super civitatem hanc? Et vos additis iracundiam super Israel profanando sabbatum! ".
NEH|13|19|Factum est autem, cum obscuratae essent portae Ierusalem ante diem sabbati, dixi, et clauserunt ianuas; et praecepi, ut non aperirent eas usque post sabbatum. Et de pueris meis constitui super portas, ut nullus inferret onus in die sabbati.
NEH|13|20|Et manserunt negotiatores et vendentes universa venalia foris Ierusalem semel et bis.
NEH|13|21|Et contestatus sum eos et dixi eis: " Quare manetis ex adverso muri? Si iterum hoc feceritis, manum mittam in vos ". Itaque ex tempore illo non venerunt in sabbato.
NEH|13|22|Dixi quoque Levitis, ut mundarentur et venirent ad custodiendas portas et sanctificandam diem sabbati.Et pro hoc ergo memento mei, Deus meus, et parce mihi secundum multitudinem miserationum tuarum!
NEH|13|23|Sed et in diebus illis vidi Iudaeos, qui duxerant uxores Azotidas, Ammonitidas et Moabitidas.
NEH|13|24|Et filii eorum ex media parte loquebantur Azotice et nesciebant loqui Iudaice vel loquebantur iuxta linguam unius vel alterius populi.
NEH|13|25|Et obiurgavi eos et maledixi et cecidi quosdam ex eis et decalvavi eos; et adiuravi in Deo, ut non darent filias suas filiis eorum et non acciperent de filiabus eorum filiis suis et sibimetipsis dicens:
NEH|13|26|" Numquid non in huiuscemodi re peccavit Salomon rex Israel? Et certe in gentibus multis non erat rex similis ei, et dilectus Deo suo erat, et posuit eum Deus regem super omnem Israel; et ipsum ergo duxerunt ad peccatum mulieres alienigenae.
NEH|13|27|Numquid et vobis obsequentes faciemus omne malum grande hoc, ut praevaricemur in Deo nostro et ducamus uxores peregrinas? ".
NEH|13|28|Unus autem de filiis Ioiada filii Eliasib sacerdotis magni gener erat Sanaballat Horonites, quem fugavi a me.
NEH|13|29|Recordare, Domine Deus meus, adversum eos, qui polluunt sacerdotium et pactum sacerdotale et leviticum!
NEH|13|30|Igitur mundavi eos ab omnibus alienigenis et constitui ordines pro sacerdotibus et Levitis, unumquemque in ministerio suo,
NEH|13|31|et pro oblatione lignorum in temporibus constitutis et pro primitiis. Memento mei, Deus meus, in bonum.
ESTH|1|1|Et fuit in diebus Asueri, qui regnavit ab India usque Aethiopiam super centum viginti septem provincias,
ESTH|1|2|quando sedit in solio regni sui in castris Susan,
ESTH|1|3|tertio igitur anno imperii sui, fecit grande convivium cunctis principibus et pueris suis, fortissimis Persarum et Medorum, inclitis et praefectis provinciarum coram se,
ESTH|1|4|ut ostenderet divitias gloriae regni sui ac splendorem atque iactantiam magnitudinis suae multo tempore, centum videlicet et octoginta diebus.
ESTH|1|5|Cumque implerentur dies convivii, invitavit omnem populum, qui inventus est in Susan, a maximo usque ad minimum; et septem diebus iussit convivium praeparari in vestibulo horti palatii regis.
ESTH|1|6|Et pendebant ex omni parte tentoria lintea et carbasina ac hyacinthina sustentata funibus byssinis atque purpureis, qui argenteis circulis inserti erant et columnis marmoreis fulciebantur; lectuli quoque aurei et argentei dispositi erant super pavimentum smaragdino et pario stratum lapide aliisque varii coloris.
ESTH|1|7|Bibebant autem, qui invitati erant, aureis poculis, aliis atque aliis; vinum quoque, ut magnificentia regia dignum erat, abundans et praecipuum ponebatur.
ESTH|1|8|Nec erat qui cogeret ad bibendum, quoniam sic rex statuerat omnibus praepositis domus suae, ut facerent secundum uniuscuiusque voluntatem.
ESTH|1|9|Vasthi quoque regina fecit convivium feminarum in palatio regio, ubi rex Asuerus manere consueverat.
ESTH|1|10|Itaque die septimo, cum rex esset hilarior potione meri, praecepit Mauman et Bazatha et Harbona et Bagatha et Abgatha et Zethar et Charchas, septem eunuchis, qui in conspectu eius ministrabant,
ESTH|1|11|ut introducerent reginam Vasthi coram rege, posito super caput eius diademate regni, ut ostenderet cunctis populis et principibus pulchritudinem illius; erat enim pulchra valde.
ESTH|1|12|Quae renuit et ad regis imperium, quod per eunuchos mandaverat, venire contempsit; unde iratus rex et nimio furore succensus
ESTH|1|13|interrogavit sapientes, qui tempora noverant, et illorum faciebat cuncta consilio scientium leges ac iura maiorum -
ESTH|1|14|erant autem ei proximi Charsena et Sethar et Admatha et Tharsis et Mares et Marsana et Mamuchan, septem duces Persarum atque Medorum, qui videbant faciem regis et primi sedebant in regno C:
ESTH|1|15|" Secundum legem quid oportet fieri Vasthi reginae, quae Asueri regis imperium, quod per eunuchos mandaverat, facere noluit? ".
ESTH|1|16|Responditque Mamuchan, audiente rege atque principibus: " Non solum regem laesit regina Vasthi, sed et omnes principes et populos, qui sunt in cunctis provinciis regis Asueri.
ESTH|1|17|Egredietur enim sermo reginae ad omnes mulieres, ut contemnant viros suos et dicant: "Rex Asuerus iussit, ut regina Vasthi intraret ad eum, et illa noluit".
ESTH|1|18|Atque hac ipsa die dicent omnes principum coniuges Persarum atque Medorum quem audierint sermonem reginae principibus regis; unde despectio et indignatio.
ESTH|1|19|Si tibi, rex, placet, egrediatur edictum a facie tua et scribatur inter leges Persarum atque Medorum, quas immutari illicitum est, ut nequaquam ultra Vasthi ingrediatur ad regem, sed regnum illius altera, quae melior illa est, accipiat.
ESTH|1|20|Et hoc in omne, quod latissimum est, provinciarum tuarum divulgetur imperium, et cunctae uxores, tam maiorum quam minorum, deferent maritis suis honorem ".
ESTH|1|21|Placuit consilium eius regi et principibus, fecitque rex iuxta consilium Mamuchan.
ESTH|1|22|Et misit epistulas ad universas provincias regni sui, ut quaeque gens audire et legere poterat, diversis linguis et litteris, esse viros principes ac maiores in domibus suis et subditas habere omnes mulieres, quae essent cum eis.
ESTH|2|1|His ita gestis, postquam regis Asueri deferbuerat indignatio, recordatus est Vasthi, et quae fecisset vel quae passa esset.
ESTH|2|2|Dixeruntque pueri regis ac ministri eius: " Quaerantur regi puellae virgines ac speciosae,
ESTH|2|3|et constituantur, qui considerent per universas provincias puellas speciosas et virgines et adducant eas ad civitatem Susan et tradant in domum feminarum sub manu Egei eunuchi, qui est praepositus et custos mulierum regiarum; et accipiant mundum muliebrem.
ESTH|2|4|Et, quaecumque inter omnes oculis regis placuerit, ipsa regnet pro Vasthi ". Placuit sermo regi; et ita, ut suggesserant, iussit fieri.
ESTH|2|5|Erat vir Iudaeus in Susan civitate vocabulo Mardochaeus filius Iair filii Semei filii Cis de tribu Beniamin,
ESTH|2|6|qui translatus fuerat de Ierusalem cum captivis, qui ducti fuerant cum Iechonia rege Iudae, quem Nabuchodonosor rex Babylonis transtulerat.
ESTH|2|7|Qui fuit nutricius filiae patrui sui Edissae, quae altero nomine Esther vocabatur et utrumque parentem amiserat: pulchra aspectu et decora facie. Mortuisque patre eius ac matre, Mardochaeus sibi eam adoptavit in filiam.
ESTH|2|8|Et factum est, cum percrebruisset regis imperium, et iuxta mandatum illius multae virgines pulchrae adducerentur Susan et Egeo traderentur, Esther quoque in domum regis in manus Egei custodis feminarum tradita est.
ESTH|2|9|Quae placuit ei et invenit gratiam in conspectu illius; et acceleravit mundum muliebrem et tradidit ei partes suas et septem puellas speciosissimas de domo regis, et tam ipsam quam pedisequas eius transtulit in optimam partem domus feminarum.
ESTH|2|10|Quae non indicaverat ei populum et cognationem suam; Mardochaeus enim praeceperat, ut de hac re omnino reticeret.
ESTH|2|11|Qui deambulabat cotidie ante vestibulum domus, in qua electae virgines servabantur, curam agens salutis Esther et scire volens quid ei accideret.
ESTH|2|12|Cum autem venisset tempus singularum per ordinem puellarum, ut intrarent ad regem, expletis omnibus, quae ad cultum muliebrem pertinebant, per menses duodecim; ita dumtaxat, ut sex mensibus oleo ungerentur myrrhino et aliis sex feminarum pigmentis et aromatibus uterentur,
ESTH|2|13|ingredientesque ad regem, quidquid postulassent, accipiebant, ut portarent secum de triclinio feminarum ad regis cubiculum.
ESTH|2|14|Et, quae intraverat vespere, mane iterum in domum feminarum deducebatur, sub manu Sasagazi eunuchi, qui concubinis praesidebat. Nec habebat potestatem ad regem ultra redeundi, nisi voluisset rex et eam venire iussisset ex nomine.
ESTH|2|15|Evoluto autem tempore per ordinem, instabat dies, quo Esther filia Abihail patrui Mardochaei, quam sibi adoptaverat in filiam, intrare deberet ad regem. Quae non quaesivit quidquam, nisi quae voluit Egeus eunuchus custos feminarum, et omnium oculis gratiosa et amabilis videbatur.
ESTH|2|16|Ducta est itaque ad cubiculum regis Asueri mense decimo, qui vocatur Tebeth, septimo anno regni eius.
ESTH|2|17|Et amavit eam rex plus quam omnes mulieres; habuitque gratiam et favorem coram eo super omnes virgines, et posuit diadema regni in capite eius fecitque eam regnare in loco Vasthi.
ESTH|2|18|Et iussit convivium praeparari magnificum cunctis principibus et servis suis, convivium Esther; et dedit remissionem tributi universis provinciis ac dona largitus est iuxta magnificentiam principalem.
ESTH|2|19|Mardochaeus autem manebat ad regis ianuam,
ESTH|2|20|necdum prodiderat Esther cognationem et populum suum iuxta mandatum eius; quidquid enim ille praecipiebat, observabat Esther, ut eo tempore solita erat, quo eam parvulam nutriebat.
ESTH|2|21|Eo igitur tempore, quo Mardochaeus ad regis ianuam morabatur, irati sunt Bagathan et Thares, duo eunuchi regis, qui ianitores erant volueruntque in regem mittere manus.
ESTH|2|22|Quod Mardochaeum non latuit; statimque nuntiavit reginae Esther, et illa regi ex nomine Mardochaei.
ESTH|2|23|Quaesitum est et inventum, et appensus uterque eorum in patibulo; mandatumque est libro annalium coram rege.
ESTH|3|1|Post haec rex Asuerus exaltavit Aman filium Amadathi, qui erat de stirpe Agag, et posuit solium eius super omnes principes, quos habebat.
ESTH|3|2|Cunctique servi regis, qui in foribus palatii versabantur, flectebant genua et adorabant Aman; sic enim praeceperat rex pro illo. Solus Mardochaeus non flectebat genu neque adorabat eum.
ESTH|3|3|Cui dixerunt pueri regis, qui ad fores palatii praesidebant: " Cur non observas mandatum regis? ".
ESTH|3|4|Cumque hoc crebrius dicerent, et ille nollet audire, nuntiaverunt Aman scire cupientes utrum perseveraret in sententia; dixerat enim eis se esse Iudaeum.
ESTH|3|5|Cumque Aman experimento probasset quod Mardochaeus non sibi flecteret genu nec se adoraret, iratus est valde
ESTH|3|6|et pro nihilo duxit in unum Mardochaeum mittere manus suas - audierat enim quod esset gentis Iudaeae - magisque voluit omnem Iudaeorum, qui erant in regno Asueri, perdere nationem.
ESTH|3|7|Mense primo, cuius vocabulum est Nisan, anno duodecimo regni Asueri, missa est in urnam sors, quae dicitur Phur, coram Aman, quo die et quo mense gens Iudaeorum deberet interfici; et exivit dies tertia decima mensis duodecimi, qui vocatur Adar.
ESTH|3|8|Dixitque Aman regi Asuero: " Est populus per omnes provincias regni tui dispersus, segregatus inter populos alienisque utens legibus, quas ceteri non cognoscunt, insuper et regis scita contemnens; non expedit regi, ut det illis requiem.
ESTH|3|9|Si tibi placet, scriptis decerne, ut pereat, et decem milia talentorum argenti appendam arcariis gazae tuae ".
ESTH|3|10|Tulit ergo rex anulum, quo utebatur, de manu sua et dedit eum Aman filio Amadathi de progenie Agag, hosti Iudaeorum.
ESTH|3|11|Dixitque ad eum: " Argentum, quod polliceris, tuum sit; de populo age, quod tibi placet ".
ESTH|3|12|Vocatique sunt scribae regis mense primo, tertia decima die eius, et scriptum est, ut iusserat Aman, ad omnes satrapas regis et duces provinciarum et principes diversarum gentium, ut quaeque gens legere poterat et audire pro varietate linguarum, ex nomine regis Asueri; et litterae ipsius signatae anulo.
ESTH|3|13|Missae sunt epistulae per cursores ad universas provincias regis, ut perderent, occiderent atque delerent omnes Iudaeos, a puero usque ad senem, parvulos et mulieres uno die, hoc est tertio decimo mensis duodecimi, qui vocatur Adar, et bona eorum diriperent.
ESTH|3|14|Exemplar autem epistularum ut lex in omnibus provinciis promulgandum erat, ut scirent omnes populi et pararent se ad praedictam diem.
ESTH|3|15|Festinabant cursores, qui missi erant, regis imperium explere; statimque in Susan pependit edictum, rege et Aman celebrante convivium, dum civitas ipsa esset conturbata.
ESTH|4|1|Cum comperisset Mardochaeus omnia, quae acciderant, scidit vestimenta sua et indutus est sacco spargens cinerem capiti. Et in platea mediae civitatis voce magna et amara clamabat
ESTH|4|2|usque ad fores palatii gradiens; non enim erat licitum indutum sacco aulam regis intrare.
ESTH|4|3|In omnibus quoque provinciis, quocumque edictum et dogma regis pervenerat, planctus ingens erat apud Iudaeos, ieiunium, ululatus et fletus, sacco et cinere multis pro strato utentibus.
ESTH|4|4|Ingressae sunt autem puellae Esther et eunuchi nuntiaveruntque ei. Quod audiens consternata est valde et misit vestem, ut, ablato sacco, induerent eum; quam accipere noluit.
ESTH|4|5|Accitoque Athach eunucho, quem rex ministrum ei dederat, praecepit ei, ut iret ad Mardochaeum et disceret ab eo cur hoc faceret.
ESTH|4|6|Egressusque Athach ivit ad Mardochaeum stantem in platea civitatis ante ostium palatii.
ESTH|4|7|Qui indicavit ei omnia, quae ei acciderant, quantum Aman promisisset, ut in thesauros regis pro Iudaeorum nece inferret argentum.
ESTH|4|8|Exemplar quoque edicti, quod pendebat in Susan ad perdendum eos, dedit ei, ut reginae ostenderet et moneret eam, ut intraret ad regem et deprecaretur eum et rogaret pro populo suo. 8a " Memor, inquit, dierum humilitatis tuae, quando nutrita sis in manu mea, quia Aman secundus a rege locutus est contra nos in mortem. Et tu, invoca Dominum et loquere regi pro nobis et libera nos de morte ".
ESTH|4|9|Regressus Athach nuntiavit Esther omnia, quae Mardochaeus dixerat.
ESTH|4|10|Quae respondit ei et iussit, ut diceret Mardochaeo:
ESTH|4|11|" Omnes servi regis et cunctae, quae sub dicione eius sunt, norunt provinciae, quod cuique sive viro sive mulieri, qui non vocatus interius atrium regis intraverit, una lex sit, ut statim interficiatur, nisi forte rex auream virgam ad eum tetenderit, ut possit vivere; ego autem triginta iam diebus non sum vocata ad regem ".
ESTH|4|12|Quod cum audisset Mardochaeus,
ESTH|4|13|rursum mandavit Esther dicens: " Ne putes quod animam tuam tantum liberes, quia in domo regis es, prae cunctis Iudaeis.
ESTH|4|14|Si enim nunc silueris, aliunde Iudaeis liberatio et salvatio exsurget, et tu et domus patris tui peribitis; et quis novit utrum idcirco ad regnum veneris, ut in tali tempore parareris? ".
ESTH|4|15|Rursumque Esther haec Mardochaeo verba mandavit:
ESTH|4|16|" Vade et congrega omnes Iudaeos, qui in Susan reperiuntur; et ieiunate pro me. Non comedatis et non bibatis tribus diebus et tribus noctibus, et ego cum ancillis meis similiter ieiunabo; et tunc ingrediar ad regem contra legem faciens; si pereo, pereo ".
ESTH|4|17|Ivit itaque Mardochaeus et fecit omnia, quae ei Esther mandaverat.
ESTH|5|1|Et factum est die tertio, induta Esther regalibus vestimentis ste tit in atrio domus regiae, quod erat interius contra basilicam regis. At ille sedebat super solium suum in consistorio palatii contra ostium domus.
ESTH|5|2|Et factum est, cum vidisset Esther reginam stantem, placuit oculis eius, et extendit contra eam virgam auream, quam tenebat manu; quae accedens tetigit summitatem virgae eius.
ESTH|5|3|Dixitque ad eam rex: " Quid vis, Esther regina? Quae est petitio tua? Etiamsi dimidiam partem regni petieris, dabitur tibi ".
ESTH|5|4|At illa respondit: " Si regi placet, obsecro, ut venias ad me hodie et Aman tecum ad convivium, quod paravi ".
ESTH|5|5|Statimque rex: " Vocate, inquit, cito Aman, ut fiat verbum Esther ".Venerunt itaque rex et Aman ad convivium, quod eis regina paraverat.
ESTH|5|6|Dixitque ei rex, postquam vinum biberat: " Quid petis, ut detur tibi, et pro qua re postulas? Etiamsi dimidiam partem regni mei petieris, impetrabis ".
ESTH|5|7|Cui respondit Esther: " Petitio mea et preces:
ESTH|5|8|Si inveni in conspectu regis gratiam, et si regi placet, ut det mihi, quod postulo, et meam impleat petitionem, veniat rex et Aman ad convivium, quod parabo eis, et cras faciam secundum verbum regis ".
ESTH|5|9|Egressus est itaque illo die Aman laetus et alacer corde. Cumque vidisset Mardochaeum sedentem in foribus palatii, et non solum non assurrexisse sibi, sed nec motum quidem de loco sessionis suae, indignatus est valde.
ESTH|5|10|Et, dissimulata ira, reversus in domum suam convocavit ad se amicos suos et Zares uxorem suam
ESTH|5|11|et exposuit illis magnitudinem divitiarum suarum filiorumque turbam, et quanta eum gloria super omnes principes et servos suos rex elevasset.
ESTH|5|12|Et post haec ait: " Regina quoque Esther nullum alium vocavit ad convivium cum rege praeter me; apud quam etiam cras cum rege pransurus sum.
ESTH|5|13|Et, cum omnia haec habeam, nihil me habere puto, quamdiu videro Mardochaeum Iudaeum sedentem in foribus regis ".
ESTH|5|14|Responderuntque ei Zares uxor eius et ceteri amici: " Iube parari excelsam trabem habentem altitudinis quinquaginta cubitos et dic mane regi, ut appendatur super eam Mardochaeus; et sic ibis cum rege laetus ad convivium ". Placuit ei consilium et iussit excelsam parari trabem.
ESTH|6|1|Noctem illam duxit rex insomnem iussitque afferri sibi librum memorialium, annales priorum temporum. Quae cum illo praesente legerentur,
ESTH|6|2|ventum est ad eum locum, ubi scriptum erat quomodo nuntiasset Mardochaeus insidias Bagathan et Thares duorum eunuchorum ianitorum, qui voluerant manus mittere in regem Asuerum.
ESTH|6|3|Quod cum audisset rex, ait: " Quid pro hac fide honoris ac praemii Mardochaeus consecutus est? ". Dixeruntque ei servi illius ac ministri: " Nihil omnino mercedis accepit ".
ESTH|6|4|Statimque rex: " Quis est, inquit, in atrio? ". Aman quippe exterius atrium domus regiae intraverat, ut suggereret regi, ut iuberet Mardochaeum suspendi in patibulo, quod ei fuerat praeparatum.
ESTH|6|5|Responderunt pueri: " Ecce Aman stat in atrio ". Dixitque rex: " Ingrediatur ".
ESTH|6|6|Cumque esset ingressus, ait illi: " Quid debet fieri viro, quem rex honorare desiderat? ". Cogitans autem in corde suo Aman et reputans quod nullum alium rex nisi se vellet honorare
ESTH|6|7|respondit: " Homo, quem rex honorare cupit,
ESTH|6|8|debet indui vestibus regiis, quibus rex indutus erat, et imponi super equum, qui de sella regis est, et acceperit regium diadema super caput suum;
ESTH|6|9|et primus de regiis principibus nobilissimis induat eum et teneat equum eius et per plateam civitatis incedens clamet et dicat: "Sic honorabitur quemcumque voluerit rex honorare" ".
ESTH|6|10|Dixitque ei rex: " Festina et, sumpta stola et equo, fac, ut locutus es, Mardochaeo Iudaeo, qui sedet in foribus palatii; cave, ne quidquam de his, quae locutus es, praetermittas ".
ESTH|6|11|Tulit itaque Aman stolam et equum; indutumque Mardochaeum et impositum equo praecedebat in platea civitatis atque clamabat: " Hoc honore condignus est quemcumque rex voluerit honorare ".
ESTH|6|12|Reversusque est Mardochaeus ad ianuam palatii; et Aman festinavit ire in domum suam lugens et operto capite.
ESTH|6|13|Narravitque Zares uxori suae et amicis omnia, quae evenissent sibi; cui responderunt sapientes, quos habebat in consilio, et uxor eius: " Si de semine Iudaeorum est Mardochaeus, ante quem cadere coepisti, non poteris praevalere contra eum, sed cades in conspectu eius ".
ESTH|6|14|Adhuc illis loquentibus, venerunt eunuchi regis et cito eum ad convivium, quod regina paraverat, pergere compulerunt.
ESTH|7|1|Intravit itaque rex et Aman, ut biberent cum regina.
ESTH|7|2|Dixitque ei rex etiam in secundo die, postquam vino incaluerat: " Quae est petitio tua, Esther, ut detur tibi, et quid vis fieri? Etiamsi dimidiam regni mei partem petieris, impetrabis ".
ESTH|7|3|Ad quem illa respondit: " Si inveni gratiam in oculis tuis, o rex, et si tibi placet, dona mihi animam meam, pro qua rogo, et populum meum, pro quo obsecro.
ESTH|7|4|Traditi enim sumus, ego et populus meus, ut conteramur, iugulemur et pereamus. Atque utinam in servos et famulas venderemur: tacuissem, quia tribulatio haec non esset digna conturbare regem ".
ESTH|7|5|Respondensque rex Asuerus ait: " Quis est iste et ubi est, ut haec audeat facere? ".
ESTH|7|6|Dixit Esther: " Hostis et inimicus noster pessimus iste est Aman ". Quod ille audiens ilico obstupuit coram rege ac regina.
ESTH|7|7|Rex autem surrexit iratus et de loco convivii intravit in hortum palatii. Aman quoque surrexit, ut rogaret Esther reginam pro anima sua; intellexit enim a rege sibi decretum esse malum.
ESTH|7|8|Qui cum reversus esset de horto et intrasset convivii locum, repperit Aman super lectulum corruisse, in quo iacebat Esther, et ait: " Etiam reginam vult opprimere, me praesente, in domo mea? ". Necdum verbum de ore regis exierat, et statim operuerunt faciem eius.
ESTH|7|9|Dixitque Harbona, unus de eunuchis, qui stabant in ministerio regis: " En etiam lignum, quod paraverat Mardochaeo, qui locutus est bonum pro rege, stat in domo Aman habens altitudinis quinquaginta cubitos ". Cui dixit rex: " Appendite eum in eo ".
ESTH|7|10|Suspensus est itaque Aman in patibulo, quod paraverat Mardochaeo; et regis ira quievit.
ESTH|8|1|Die illo dedit rex Asuerus Esther reginae domum Aman adversarii Iudaeorum, et Mardochaeus ingressus est ante faciem regis; confessa est enim ei Esther quid esset sibi.
ESTH|8|2|Tulitque rex anulum suum, quem ab Aman recipi iusserat, et tradidit Mardochaeo; Esther autem constituit Mardochaeum super domum Aman.
ESTH|8|3|Et adiecit Esther loqui coram rege et procidit ad pedes eius flevitque et locuta ad eum oravit, ut malitiam Aman Agagitae et machinationes eius pessimas, quas excogitaverat contra Iudaeos, iuberet irritas fieri.
ESTH|8|4|At ille ex more sceptrum aureum protendit manu; illaque consurgens stetit ante eum
ESTH|8|5|et ait: " Si placet regi, et si inveni gratiam coram eo, et deprecatio mea non ei videtur esse contraria, et accepta sum in oculis eius, obsecro, ut novis epistulis veteres litterae Aman filii Amadathi, Agagitae, insidiatoris et hostis Iudaeorum, quibus eos in cunctis regis provinciis perire praeceperat, corrigantur.
ESTH|8|6|Quomodo enim potero sustinere malum, quod passurus est populus meus, et interitum cognationis meae? ".
ESTH|8|7|Responditque rex Asuerus Esther reginae et Mardochaeo Iudaeo: " Domum Aman concessi Esther et ipsum iussi appendi in patibulo, quia ausus est manum in Iudaeos mittere.
ESTH|8|8|Scribite ergo Iudaeis sicut vobis placet, ex regis nomine, signantes litteras anulo meo, quia epistulae ex regis nomine scriptae et illius anulo signatae non possunt immutari ".
ESTH|8|9|Accitisque scribis regis - erat autem tempus tertii mensis, qui appellatur Sivan, vicesima et tertia illius die - scriptae sunt epistulae, ut Mardochaeus voluerat, ad Iudaeos et ad satrapas procuratoresque et principes, qui centum viginti septem provinciis ab India usque ad Aethiopiam praesidebant, provinciae atque provinciae, populo et populo, iuxta linguas et litteras suas, et Iudaeis iuxta linguam et litteras suas.
ESTH|8|10|Ipsaeque epistulae, quae ex regis nomine mittebantur, anulo ipsius obsignatae sunt et missae per veredarios electis equis regiis discurrentes.
ESTH|8|11|Quibus permisit rex Iudaeis in singulis civitatibus, ut in unum congregarentur et starent pro animabus suis et omnes inimicos suos cum coniugibus ac liberis interficerent atque delerent et spolia eorum diriperent;
ESTH|8|12|et constituta est per omnes provincias una ultionis dies, id est tertia decima mensis duodecimi, qui vocatur Adar.
ESTH|8|13|Exemplar epistulae in forma legis in omnibus provinciis promulgandum erat, ut omnibus populis notum fieret paratos esse Iudaeos in diem illam ad capiendam vindictam de hostibus suis.
ESTH|8|14|Egressique sunt veredarii celeres nuntios perferentes, et edictum regis pependit in Susan.
ESTH|8|15|Mardochaeus autem de palatio et de conspectu regis egrediens fulgebat vestibus regiis, hyacinthinis videlicet et albis, coronam magnam auream portans in capite et amictus pallio serico atque purpureo; omnisque civitas exsultavit atque laetata est.
ESTH|8|16|Iudaeis autem nova lux oriri visa est, gaudium, honor et tripudium.
ESTH|8|17|Apud omnes populos, urbes atque provincias, quocumque regis iussa veniebant, Iudaeis fuit exsultatio, epulae atque convivia et festus dies, in tantum ut plures alterius gentis et sectae eorum religioni et caeremoniis iungerentur; grandis enim cunctos Iudaici nominis terror invaserat.
ESTH|9|1|Igitur duodecimi mensis - id est Adar - tertia decima die, quando verbum et edictum regis explendum erat, et hostes Iudaeorum sperabant quod dominarentur ipsis, versa vice Iudaei superaverunt adversarios suos.
ESTH|9|2|Congregatique sunt per singulas civitates, ut extenderent manum contra inimicos et persecutores suos; nullusque ausus est resistere, eo quod omnes populos invaserat formido eorum.
ESTH|9|3|Nam et omnes provinciarum principes et satrapae et procuratores omnisque dignitas, quae singulis locis ac operibus praeerat, sustinebant Iudaeos timore Mardochaei,
ESTH|9|4|quem principem esse palatii et plurimum posse cognoverant; fama quoque nominis eius crescebat cotidie et per cunctorum ora volitabat.
ESTH|9|5|Itaque percusserunt Iudaei omnes inimicos suos plaga gladii et necis et interitus, reddentes eis, quod sibi paraverant facere.
ESTH|9|6|In Susan quingentos viros interfecerunt, extra decem filios Aman Agagitae hostis Iudaeorum, quorum ista sunt nomina:
ESTH|9|7|Pharsandatha et Delphon et Esphatha
ESTH|9|8|et Phoratha et Adalia et Aridatha
ESTH|9|9|et Phermesta et Arisai et Aridai et Iezatha.
ESTH|9|10|Quos cum occidissent, praedas de substantiis eorum tangere noluerunt.
ESTH|9|11|Statimque numerus eorum, qui occisi erant in Susan, ad regem relatus est.
ESTH|9|12|Qui dixit reginae: " In urbe Susan interfecerunt et deleverunt Iudaei quingentos viros et decem filios Aman. Quantam putas eos exercuisse caedem in universis provinciis? Quid ultra postulas et quid vis, ut fieri iubeam?.
ESTH|9|13|Cui illa respondit: " Si regi placet, detur potestas Iudaeis, qui in Susan sunt, ut sicut hodie fecerunt, sic et cras faciant, et decem filii Aman in patibulo suspendantur ".
ESTH|9|14|Praecepitque rex, ut ita fieret. Statimque in Susan pependit edictum, et decem filii Aman suspensi sunt.
ESTH|9|15|Congregatis igitur Iudaeis, qui in Susan erant, quarta decima die mensis Adar, interfecti sunt in Susan trecenti viri, nec eorum ab illis direpta substantia est.
ESTH|9|16|Reliqui autem Iudaei per omnes provincias, quae dicioni regis subiacebant, congregati pro animabus suis steterunt, ut requiescerent ab hostibus, ac interfecerunt de persecutoribus suis septuaginta quinque milia, sed nullus de substantiis eorum quidquam contigit.
ESTH|9|17|Dies autem tertius decimus mensis Adar, dies apud omnes interfectionis fuit, et quarta decima die requieverunt. Quem constituerunt esse diem epularum et laetitiae.
ESTH|9|18|At hi, qui in urbe Susan congregati sunt, tertio decimo et quarto decimo die eiusdem mensis in caede versati sunt, quinto decimo autem die requieverunt; et idcirco eundem diem constituerunt sollemnem epularum atque laetitiae.
ESTH|9|19|Hi vero Iudaei, qui in oppidis non muratis ac villis morabantur, quartum decimum diem mensis Adar conviviorum et gaudii decreverunt, ita ut exsultent in eo et mittant sibi mutuo partes epularum. Illi autem, qui in urbibus habitant, agunt etiam quintum decimum diem mensis Adar cum gaudio et convivio et ut diem festum, in quo mittunt sibi mutuo partes epularum.
ESTH|9|20|Scripsit itaque Mardochaeus omnia haec et litteris comprehensa misit ad omnes Iudaeos, qui in omnibus regis provinciis morabantur, tam in vicino positis quam procul,
ESTH|9|21|ut quartam decimam et quintam decimam diem mensis Adar pro festis susciperent et, revertente semper anno, sollemni honore celebrarent
ESTH|9|22|secundum dies, in quibus requieverunt Iudaei ab inimicis suis, et mensem, qui de luctu atque tristitia in hilaritatem gaudiumque ipsis conversus est, essentque istae dies epularum atque laetitiae, et mitterent sibi invicem ciborum partes et pauperibus munuscula largirentur.
ESTH|9|23|Susceperuntque Iudaei in sollemnem ritum cuncta, quae eo tempore facere coeperant, et quae Mardochaeus litteris facienda mandaverat.
ESTH|9|24|Aman enim filius Amadathi stirpis Agag, adversarius omnium Iudaeorum, cogitavit contra eos malum, ut deleret illos, et misit Phur, id est sortem, ut eos conturbaret atque deleret.
ESTH|9|25|Sed postquam ingressa est Esther ad regem, mandavit ille simul cum litteris, ut malum, quod iste contra Iudaeos cogitaverat, reverteretur in caput eius, et suspenderentur ipse et filii eius in patibulo.
ESTH|9|26|Atque ex illo tempore dies isti appellati sunt Phurim propter nomen Phur. Propter cuncta illa, quae in hac epistula continentur,
ESTH|9|27|et propter ea, quae de his viderant et quae eis acciderant, statuerunt et in sollemnem ritum numquam mutandum susceperunt Iudaei super se et semen suum et super cunctos, qui religioni eorum voluerint copulari, ut duos hos dies secundum praeceptum et tempus eorum singulis annis celebrarent.
ESTH|9|28|Isti dies memorarentur et celebrarentur per singulas generationes in singulis cognationibus, provinciis et civitatibus, nec esset ulla civitas, in qua dies Phurim non observarentur a Iudaeis et ab eorum progenie.
ESTH|9|29|Scripseruntque Esther regina filia Abihail et Mardochaeus Iudaeus omni studio ad confirmandam hanc secundam epistulam Phurim.
ESTH|9|30|Et miserunt ad omnes Iudaeos, qui in centum viginti septem provinciis regis Asueri versabantur, verba pacis et veritatis,
ESTH|9|31|statuentes dies Phurim pro temporibus suis, sicut constituerant Mardochaeus et Esther, et sicut illi statuerant pro seipsis et pro semine suo, praecepta ieiuniorum et clamorum.
ESTH|9|32|Et mandatum Esther confirmavit praecepta Phurim et scriptum est in libro.
ESTH|10|1|Rex vero Asuerus terrae et maris insulis imposuit tribu tum.
ESTH|10|2|Cuius fortitudo et imperium et dignitas atque sublimitas, qua exaltavit Mardochaeum, scripta sunt in libro annalium regum Medorum atque Persarum,
ESTH|10|3|et quomodo Mardochaeus Iudaici generis secundus a rege Asuero fuerit et magnus apud Iudaeos et acceptabilis plebi fratrum suorum, quaerens bona populo suo et loquens ea, quae ad pacem seminis sui pertinerent.
JOB|1|1|Vir erat in terra Us nomine Iob, et erat vir ille simplex et rectus ac timens Deum et recedens a malo.
JOB|1|2|Natique sunt ei septem filii et tres filiae.
JOB|1|3|Et fuit possessio eius septem milia ovium et tria milia camelorum, quingenta quoque iuga boum et quingentae asinae ac familia multa nimis; eratque vir ille magnus inter omnes Orientales.
JOB|1|4|Et ibant filii eius et faciebant convivium per domos unusquisque in die suo; et mittentes vocabant tres sorores suas, ut comederent et biberent cum eis.
JOB|1|5|Cumque in orbem transissent dies convivii, mittebat ad eos Iob et sanctificabat illos; consurgensque diluculo offerebat holocausta pro singulis. Dicebat enim: " Ne forte peccaverint filii mei et benedixerint Deo in cordibus suis ". Sic faciebat Iob cunctis diebus.
JOB|1|6|Quadam autem die, cum venissent filii Dei, ut assisterent coram Domino, affuit inter eos etiam Satan.
JOB|1|7|Cui dixit Dominus: " Unde venis? ". Qui respondens ait: " Circuivi terram et perambulavi eam ".
JOB|1|8|Dixitque Dominus ad eum: " Numquid considerasti servum meum Iob, quod non sit ei similis in terra, homo simplex et rectus ac timens Deum et recedens a malo? ".
JOB|1|9|Cui respondens Satan ait: " Numquid Iob frustra timet Deum?
JOB|1|10|Nonne tu vallasti eum ac domum eius universamque substantiam per circuitum, operibus manuum eius benedixisti, et possessio eius crevit in terra?
JOB|1|11|Sed extende paululum manum tuam et tange cuncta, quae possidet, nisi in faciem benedixerit tibi ".
JOB|1|12|Dixit ergo Dominus ad Satan: " Ecce, universa, quae habet, in manu tua sunt; tantum in eum ne extendas manum tuam ". Egressusque est Satan a facie Domini.
JOB|1|13|Cum autem quadam die filii et filiae eius comederent et biberent vinum in domo fratris sui primogeniti,
JOB|1|14|nuntius venit ad Iob, qui diceret: " Boves arabant, et asinae pascebantur iuxta eos;
JOB|1|15|et irruerunt Sabaei tuleruntque eos et pueros percusserunt gladio, et evasi ego solus, ut nuntiarem tibi ".
JOB|1|16|Cumque adhuc ille loqueretur, venit alter et dixit: " Ignis Dei cecidit e caelo et ussit oves puerosque consumpsit, et effugi ego solus, ut nuntiarem tibi ".
JOB|1|17|Sed et illo adhuc loquente, venit alius et dixit: " Chaldaei fecerunt tres turmas et invaserunt camelos et tulerunt eos necnon et pueros percusserunt gladio, et ego fugi solus, ut nuntiarem tibi ".
JOB|1|18|Adhuc loquebatur ille, et ecce alius intravit et dixit: " Filiis tuis et filiabus vescentibus et bibentibus vinum in domo fratris sui primogeniti,
JOB|1|19|repente ventus vehemens irruit a regione deserti et concussit quattuor angulos domus; quae corruens oppressit liberos tuos, et mortui sunt, et effugi ego solus, ut nuntiarem tibi ".
JOB|1|20|Tunc surrexit Iob et scidit vestimenta sua et, tonso capite, corruens in terram adoravit
JOB|1|21|et dixit: Nudus egressus sum de utero matris meaeet nudus revertar illuc.Dominus dedit, Dominus abstulit; sicut Domino placuit, ita factum est:sit nomen Domini benedictum ".
JOB|1|22|In omnibus his non peccavit Iob labiis suis neque stultum quid contra Deum locutus est.
JOB|2|1|Factum est autem, cum quadam die venissent filii Dei, ut starent coram Domino, venit quoque Satan inter eos, ut staret in conspectu eius.
JOB|2|2|Dixit Dominus ad Satan: " Unde venis? ". Qui respondens ait: " Circuivi terram et perambulavi eam ".
JOB|2|3|Et dixit Dominus ad Satan: " Numquid considerasti servum meum Iob, quod non sit ei similis in terra, vir simplex et rectus ac timens Deum et recedens a malo et adhuc retinens innocentiam? Tu autem commovisti me adversus eum, ut affligerem eum frustra ".
JOB|2|4|Cui respondens Satan ait: " Pellem pro pelle et cuncta, quae habet, homo dabit pro anima sua.
JOB|2|5|Alioquin mitte manum tuam et tange os eius et carnem; et tunc videbis, si in faciem benedicet tibi ".
JOB|2|6|Dixit ergo Dominus ad Satan: " Ecce, in manu tua est; verumtamen animam illius serva ".
JOB|2|7|Egressus igitur Satan a facie Domini, percussit Iob ulcere pessimo a planta pedis usque ad verticem eius.
JOB|2|8|Qui testa saniem radebat, sedens in sterquilinio.
JOB|2|9|Dixit autem illi uxor sua: Adhuctu permanes in simplicitate tua?Benedic Deo et morere ".
JOB|2|10|Qui ait ad illam: Quasi una de stultis mulieribuslocuta es!Si bona suscepimus de manu Dei,mala quare non suscipiamus? ".In omnibus his non peccavit Iob labiis suis.
JOB|2|11|Igitur, audientes tres amici Iob omne malum, quod accidisset ei, venerunt singuli de loco suo, Eliphaz Themanites et Baldad Suhites et Sophar Naamathites. Condixerant enim, ut pariter venientes visitarent eum et consolarentur.
JOB|2|12|Cumque elevassent procul oculos suos, non cognoverunt eum et exclamantes ploraverunt; scissisque vestibus, sparserunt pulverem super caput suum in caelum.
JOB|2|13|Et sederunt cum eo in terra septem diebus et septem noctibus, et nemo loquebatur ei verbum; videbant enim dolorem esse vehementem.
JOB|3|1|Post haec aperuit Iob os suum et maledixit diei suo
JOB|3|2|et locutus est:
JOB|3|3|" Pereat dies, in qua natus sum,et nox, in qua dictum est: "Conceptus est homo".
JOB|3|4|Dies ille vertatur in tenebras;non requirat eum Deus desuper,et non illustretur lumine.
JOB|3|5|Obscurent eum tenebrae et umbra mortis;occupet eum caligo,et involvatur amaritudine.
JOB|3|6|Noctem illam tenebrosus turbo possideat;non computetur in diebus anninec numeretur in mensibus.
JOB|3|7|Sit nox illa solitaria nec laude digna;
JOB|3|8|maledicant ei, qui maledicunt diei,qui parati sunt suscitare Leviathan.
JOB|3|9|Obtenebrentur stellae crepusculi eius;exspectet lucem, et non sit,nec videat palpebras aurorae,
JOB|3|10|quia non conclusit ostia ventris, qui portavit me,nec abstulit mala ab oculis meis.
JOB|3|11|Quare non in vulva mortuus sum?Egressus ex utero non statim perii?
JOB|3|12|Quare exceptus genibus?Cur lactatus uberibus?
JOB|3|13|Nunc enim dormiens sileremet somno meo requiescerem
JOB|3|14|cum regibus et consulibus terrae,qui aedificant sibi solitudines,
JOB|3|15|aut cum principibus, qui possident aurumet replent domos suas argento.
JOB|3|16|Aut sicut abortivum absconditum non subsisterem,vel qui concepti non viderunt lucem.
JOB|3|17|Ibi impii cessaverunt a tumultu,et ibi requieverunt fessi robore.
JOB|3|18|Et quondam vincti pariter sine molestianon audierunt vocem exactoris.
JOB|3|19|Parvus et magnus ibi sunt,et servus liber a domino suo.
JOB|3|20|Quare misero data est lux,et vita his, qui in amaritudine animae sunt?
JOB|3|21|Qui exspectant mortem, et non venit,et effodiunt quaerentes illam magis quam thesauros;
JOB|3|22|gaudentque vehementeret laetantur sepulcro.
JOB|3|23|Viro, cuius abscondita est via,et circumdedit eum Deus tenebris.
JOB|3|24|Antequam comedam, suspiro,et quasi inundantes aquae sic rugitus meus.
JOB|3|25|Quia timor, quem timebam, evenit mihi,et, quod verebar, accidit.
JOB|3|26|Non dissimulavi, non silui, non quievi,et venit super me indignatio ".
JOB|4|1|Respondens autem Eliphaz Themanites dixit:
JOB|4|2|" Si coeperimus loqui tibi, forsitan moleste accipies;sed conceptum sermonem tenere quis poterit?
JOB|4|3|Ecce, docuisti multoset manus lassas roborasti;
JOB|4|4|vacillantes confirmaverunt sermones tui,et genua trementia confortasti.
JOB|4|5|Nunc autem venit super te plaga, et defecisti;tetigit te, et conturbatus es.
JOB|4|6|Nonne timor tuus est fiducia tua,spes tua est perfectio viarum tuarum?
JOB|4|7|Recordare, obsecro te, quis umquam innocens periit,aut quando recti deleti sunt?
JOB|4|8|quin potius vidi eos, qui operantur iniquitatemet seminant dolores et metunt eos,
JOB|4|9|flante Deo perisse,et spiritu irae eius esse consumptos.
JOB|4|10|Rugitus leonis et vox leaenaeet dentes catulorum leonum contriti sunt.
JOB|4|11|Leo periit, eo quod non haberet praedam,et catuli leonis dissipati sunt.
JOB|4|12|Porro ad me furtive verbum delatum est,et suscepit auris mea sussurrum eius.
JOB|4|13|In horrore visionis nocturnae,quando solet sopor occupare homines,
JOB|4|14|pavor tenuit me et tremor,et omnia ossa mea perterrita sunt.
JOB|4|15|Et cum spiritus, me praesente, transiret,inhorruerunt pili carnis meae.
JOB|4|16|Stetit quidam, cuius non agnoscebam vultum,imago coram oculis meis,et vocem quasi aurae lenis audivi:
JOB|4|17|"Numquid homo Dei comparatione iustificabitur,aut factore suo purior erit vir?".
JOB|4|18|Ecce, in servis suis fiduciam non habetet in angelis suis reperit pravitatem.
JOB|4|19|Quanto magis hi, qui habitant domos luteas,quorum fundamentum est in pulvere.Consumentur velut tinea!
JOB|4|20|De mane usque ad vesperam succidenturet, quia nullus intellegit, in aeternum peribunt.
JOB|4|21|Nonne evulsum est reliquum eorum ab eis?Morientur, et non in sapientia.
JOB|5|1|Voca ergo, si est qui tibi re spondeat!Ad quem sanctorum converteris?
JOB|5|2|Vere stultum interficit iracundia,et fatuum occidit invidia.
JOB|5|3|Ego vidi stultum firma radiceet maledixi sedi eius statim.
JOB|5|4|Longe fient filii eius a saluteet conterentur in porta, et non erit qui eruat.
JOB|5|5|Cuius messem famelicus comedet,et ipsum rapiet armatus, et bibent sitientes divitias eius.
JOB|5|6|Quia non egreditur ex pulvere nequitia,et de humo non oritur dolor.
JOB|5|7|Sed homo generat laborem,et aves elevant volatum.
JOB|5|8|Quam ob rem ego deprecabor Dominumet ad Deum ponam eloquium meum,
JOB|5|9|qui facit magna et inscrutabiliaet mirabilia absque numero;
JOB|5|10|qui dat pluviam super faciem terraeet irrigat aquis rura;
JOB|5|11|qui ponit humiles in sublimeet maerentes erigit sospitate;
JOB|5|12|qui dissipat cogitationes malignorum,ne possint implere manus eorum, quod coeperant;
JOB|5|13|qui apprehendit sapientes in astutia eorumet consilium pravorum dissipat.
JOB|5|14|Per diem incurrent tenebraset, quasi in nocte, sic palpabunt in meridie.
JOB|5|15|Porro salvum faciet egenum a gladio oris eorumet de manu violenti pauperem;
JOB|5|16|et erit egeno spes,iniquitas autem contrahet os suum.
JOB|5|17|Beatus homo, qui corripitur a Deo;increpationem ergo Omnipotentis ne reprobes.
JOB|5|18|Quia ipse vulnerat et medetur,percutit, et manus eius sanabunt.
JOB|5|19|In sex tribulationibus liberabit te,et in septem non tanget te malum.
JOB|5|20|In fame eruet te de morteet in bello de manu gladii.
JOB|5|21|A flagello linguae absconderiset non timebis vastationem, cum venerit.
JOB|5|22|In vastitate et fame ridebiset bestias terrae non formidabis.
JOB|5|23|Sed cum lapidibus campi pactum tuum,et bestiae terrae pacificae erunt tibi.
JOB|5|24|Et scies quod pacem habeat tabernaculum tuum,et visitans habitationem tuam non falleris.
JOB|5|25|Scies quoque quoniam multiplex erit semen tuum,et progenies tua quasi herba terrae.
JOB|5|26|Ingredieris in abundantia sepulcrum,sicut infertur acervus tritici in tempore suo.
JOB|5|27|Ecce hoc, ut investigavimus, ita est;oboedi illi et tu sapias tibi ".
JOB|6|1|Respondens autem Iob dixit:
JOB|6|2|" Utinam appenderetur aegritu do mea,et calamitatem meam assumerent in statera!
JOB|6|3|Nunc vero arena maris haec gravior apparet,inde verbis meis haesito.
JOB|6|4|Quia sagittae Omnipotentis in me sunt,quarum venenum ebibit spiritus meus;et terrores Dei militant contra me.
JOB|6|5|Numquid rugiet onager, cum habuerit herbam?Aut mugiet bos, cum ante praesepe plenum steterit?
JOB|6|6|Aut poterit comedi insulsum, quod non est sale conditum?Aut poterit gustari herba insulsa?
JOB|6|7|Quae prius nolebat tangere anima mea,nunc prae angustia cibi mei sunt.
JOB|6|8|Quis det, ut veniat petitio mea,et, quod exspecto, tribuat mihi Deus?
JOB|6|9|Utinam Deus me conterat;solvat manum suam et succidat me!
JOB|6|10|Et haec mihi sit consolatio,et exsultabo vel in pavore, qui non parcat,nec celabo sermones Sancti.
JOB|6|11|Quae est enim fortitudo mea, ut sustineam?Aut quis finis meus, ut patienter agam?
JOB|6|12|Num fortitudo lapidum, fortitudo mea?Num caro mea aenea est?
JOB|6|13|An non est auxilium mihi in me,et virtus quoque remota est a me?
JOB|6|14|Qui tollit ab amico suo misericordiam,timorem Omnipotentis derelinquit.
JOB|6|15|Fratres mei mentiti sunt mesicut alveus torrentium, qui evanescunt
JOB|6|16|nigrescentes glacie,cum ingruit super eos nix.
JOB|6|17|Tempore, quo diffluunt, arescuntet, ut incaluerit, solvuntur de loco suo.
JOB|6|18|Deflectunt viatorum turmae de viis suis,ascendentes per desertum pereunt.
JOB|6|19|Commeatus Thema consideraverunt,viatores Saba speraverunt in eis.
JOB|6|20|Confusi sunt, quia speraverunt;venerunt eo usque, et pudore cooperti sunt.
JOB|6|21|Ita nunc vos facti estis mihi;videntes plagam meam, timetis.
JOB|6|22|Numquid dixi: Afferte mihiet de substantia vestra donate mihi?
JOB|6|23|vel: Liberate me de manu hostiset de manu robustorum eruite me?
JOB|6|24|Docete me, et ego tacebo,et, si quid forte ignoravi, instruite me.
JOB|6|25|Quare detraxistis sermonibus veritatis,cum e vobis nullus sit, qui possit arguere me?
JOB|6|26|Ad increpandum tantum eloquia concinnatis,sed in ventum verba desperati.
JOB|6|27|Super pupillum irruitiset subvertere nitimini amicum vestrum.
JOB|6|28|Nunc, quaeso, convertimini ad me,et in faciem vestram non mentiar.
JOB|6|29|Revertite! Nulla erit improbitas.Revertite! Adhuc praesens adest iustitia mea.
JOB|6|30|Estne in lingua mea improbitas?An palatum meum non discernit nequitiam?
JOB|7|1|Nonne militia est vita hominis super terram,et sicut dies mercennarii dies eius?
JOB|7|2|Sicut servus desiderat umbram,et sicut mercennarius praestolatur mercedem suam,
JOB|7|3|sic et ego habui menses vacuoset noctes laboriosas enumeravi mihi.
JOB|7|4|Si dormiero, dicam: Quando consurgam?Et rursum exspectabo vesperamet replebor doloribus usque crepusculum.
JOB|7|5|Induta est caro mea putredine et sordibus pulveris;cutis mea scinditur et diffluit.
JOB|7|6|Dies mei velocius transierunt quam navicula texentiset consumpti sunt deficiente filo.
JOB|7|7|Memento quia ventus est vita mea,et non revertetur oculus meus, ut videat bona.
JOB|7|8|Nec aspiciet me visus hominis;oculi tui in me, et non subsistam.
JOB|7|9|Sicut consumitur nubes et pertransit,sic, qui descenderit ad inferos, non ascendet
JOB|7|10|nec revertetur ultra in domum suam,neque cognoscet eum amplius locus eius.
JOB|7|11|Quapropter et ego non parcam ori meo;loquar in tribulatione spiritus mei, confabulabor cum amaritudine animae meae.
JOB|7|12|Numquid mare ego sum aut cetus,quia posuisti super me custodiam?
JOB|7|13|Si dixero: Consolabitur me lectulus meus,et assumet stratum meum querelam meam,
JOB|7|14|terrebis me per somniaet per visiones horrore concuties.
JOB|7|15|Quam ob rem eligit suspendium anima mea,et mortem ossa mea.
JOB|7|16|Desperavi; nequaquam ultra iam vivam.Parce mihi, nihil enim sunt dies mei.
JOB|7|17|Quid est homo, quia magnificas eum?Aut quid apponis erga eum cor tuum?
JOB|7|18|Visitas eum diluculoet singulis momentis probas illum.
JOB|7|19|Usquequo non avertes oculos a me?Nec dimittis me, ut glutiam salivam meam?
JOB|7|20|Peccavi; quid faciam tibi,o custos hominum?Quare posuisti me contrarium tibi, et factus sum mihimetipsi gravis?
JOB|7|21|Cur non tollis peccatum meumet quare non aufers iniquitatem meam?Ecce, nunc in pulvere dormiam;et, si mane me quaesieris, non subsistam! ".
JOB|8|1|Respondens autem Baldad Suhites dixit:
JOB|8|2|" Usquequo loqueris talia,et spiritus vehemens sermones oris tui?
JOB|8|3|Numquid Deus supplantat iudicium,aut Omnipotens subvertit, quod iustum est?
JOB|8|4|Et si filii tui peccaverunt ei,et dimisit eos in manu iniquitatis suae,
JOB|8|5|tu tamen, si diluculo consurrexeris ad Deumet Omnipotentem fueris deprecatus,
JOB|8|6|si mundus et rectus incesseris,statim evigilabit ad teet pacatum reddet habitaculum iustitiae tuae;
JOB|8|7|in tantum ut, si priora tua fuerint parva,et novissima tua multiplicentur nimis.
JOB|8|8|Interroga enim generationem pristinamet diligenter investiga patrum memoriam.
JOB|8|9|Hesterni quippe sumus et ignoramus,quoniam sicut umbra dies nostri sunt super terram.
JOB|8|10|Nonne ipsi docebunt te, loquentur tibiet de corde suo proferent eloquia?
JOB|8|11|Numquid virere potest scirpus absque umore,aut crescere carectum sine aqua?
JOB|8|12|Cum adhuc sit in flore, nec carpatur manu,ante omnes herbas arescit.
JOB|8|13|Sic viae omnium, qui obliviscuntur Deum,et spes impii peribit.
JOB|8|14|Cuius spes filum tenue,et sicut tela aranearum fiducia eius.
JOB|8|15|Innitetur super domum suam et non stabit;fulciet eam et non consurget.
JOB|8|16|Umectus videtur, antequam veniat sol,et in horto suo germen eius egredietur.
JOB|8|17|Super acervum petrarum radices eius densabuntur,et inter lapides commorabitur.
JOB|8|18|Si absorbuerit eum de loco suo,negabit eum et dicet: "Non novi te".
JOB|8|19|Haec est enim laetitia viae eius,ut rursum de terra alii germinentur.
JOB|8|20|Deus non proiciet simplicemnec porriget manum malignis,
JOB|8|21|donec impleatur risu os tuum,et labia tua iubilo.
JOB|8|22|Qui oderunt te, induentur confusione,et tabernaculum impiorum non subsistet ".
JOB|9|1|Et respondens Iob ait:
JOB|9|2|" Vere scio quod ita sit,et quomodo iustificabitur homo compositus Deo?
JOB|9|3|Si voluerit contendere cum eo,non poterit ei respondere unum pro mille.
JOB|9|4|Sapiens corde est et fortis robore;quis restitit ei, et pacem habuit?
JOB|9|5|Qui transtulit montes, et nescierunt hi, quos subvertit in furore suo.
JOB|9|6|Qui commovet terram de loco suo,et columnae eius concutiuntur.
JOB|9|7|Qui praecipit soli, et non oritur,et stellas claudit quasi sub signaculo.
JOB|9|8|Qui extendit caelos soluset graditur super fluctus maris.
JOB|9|9|Qui facit Arcturum et Orionaet Hyadas et interiora austri.
JOB|9|10|Qui facit magna et incomprehensibiliaet mirabilia, quorum non est numerus.
JOB|9|11|Si venerit ad me, non videbo eum;si abierit, non intellegam.
JOB|9|12|Si repente arripiet, quis eum impediet?Vel quis dicere potest: "Quid facis?".
JOB|9|13|Deus non retinet iram suam,et sub eo curvantur auxilia Rahab.
JOB|9|14|Quantus ergo sum ego, ut respondeam eiet loquar delectis verbis cum eo?
JOB|9|15|Quia, etiamsi iustus essem, non responderem,sed meum iudicem deprecarer;
JOB|9|16|et, cum invocantem exaudierit me,non credam quod audierit vocem meam.
JOB|9|17|In turbine enim conteret meet multiplicabit vulnera mea etiam sine causa.
JOB|9|18|Non concedit requiescere spiritum meumet implet me amaritudinibus.
JOB|9|19|Si fortitudo quaeritur, robustissimus est;si iudicium, quis eum arcesserit?
JOB|9|20|Si iustificare me voluero, os meum condemnabit me;si innocentem ostendero, pravum me comprobabit.
JOB|9|21|Etiamsi simplex fuero, hoc ipsum ignorabit anima mea,et contemnam vitam meam.
JOB|9|22|Unum est, quod locutus sum:Et innocentem et impium ipse consumit.
JOB|9|23|Si subito flagellum occidat,de afflictione innocentium ridebit.
JOB|9|24|Terra data est in manus impii,vultum iudicum eius operit;quod si non ille est, quis ergo est?
JOB|9|25|Dies mei velociores fuerunt cursore:fugerunt et non viderunt bonum;
JOB|9|26|pertransierunt quasi naves arundineae,sicut aquila volans ad escam.
JOB|9|27|Cum dixero: Obliviscar maerorem meum,commutabo faciem meam et hilaris fiam,
JOB|9|28|vereor omnes dolores meos,sciens quod non iustificaveris me.
JOB|9|29|Si autem et sic impius sum,quare frustra laboravi?
JOB|9|30|Si lotus fuero quasi aquis nivis,et lixivo mundavero manus meas,
JOB|9|31|tamen sordibus intinges me,et abominabuntur me vestimenta mea.
JOB|9|32|Neque enim viro, qui similis mei est, respondebo;nec vir, quocum in iudicio contendam.
JOB|9|33|Non est qui utrumque valeat arguereet ponere manum suam in ambobus.
JOB|9|34|Auferat a me virgam suam,et pavor eius non me terreat.
JOB|9|35|Loquar et non timebo eum;quia sic non mecum ipse sum.
JOB|10|1|Taedet animam meam vitae meae;dimittam adversum me eloquium meum,loquar in amaritudine animae meae.
JOB|10|2|Dicam Deo: Noli me condemnare,indica mihi cur me ita iudices.
JOB|10|3|Numquid bonum tibi videtur, si opprimas meet calumnieris me, opus manuum tuarum,et super consilium impiorum arrideas?
JOB|10|4|Numquid oculi carnei tibi sunt,aut, sicut videt homo, et tu videbis?
JOB|10|5|Numquid sicut dies hominis dies tui,et anni tui sicut humana sunt tempora,
JOB|10|6|ut quaeras iniquitatem meamet peccatum meum scruteris,
JOB|10|7|cum scias quia nihil impium fecerim,et sit nemo, qui de manu tua possit eruere?
JOB|10|8|Manus tuae fecerunt meet plasmaverunt me totum in circuitu;et sic repente praecipitas me?
JOB|10|9|Memento, quaeso, quod sicut lutum feceris meet in pulverem reduces me.
JOB|10|10|Nonne sicut lac mulsisti meet sicut caseum me coagulasti?
JOB|10|11|Pelle et carnibus vestisti me;ossibus et nervis compegisti me.
JOB|10|12|Vitam et misericordiam tribuisti mihi,et visitatio tua custodivit spiritum meum.
JOB|10|13|Licet haec celes in corde tuo,tamen scio haec in animo tuo versari.
JOB|10|14|Si peccaverim, observas meet ab iniquitate mea mundum me esse non pateris.
JOB|10|15|Et si impius fuero, vae mihi est;et si iustus, non levabo caput,saturatus afflictione et miseria.
JOB|10|16|Si superbia extollar, quasi catulum leonis capies meet iterum mirabilem te exhibebis in me.
JOB|10|17|Instauras testes tuos contra meet multiplicas iram tuam adversum me,et poenae militant in me.
JOB|10|18|Quare de vulva eduxisti me?Qui utinam consumptus essem, ne oculus me videret!
JOB|10|19|Fuissem quasi non essem,de utero translatus ad tumulum.
JOB|10|20|Numquid non paucitas dierum meorum finietur brevi?Dimitte ergo me, ut refrigerem paululum dolorem meum,
JOB|10|21|antequam vadam, et non revertar,ad terram tenebrarum et umbrae mortis,
JOB|10|22|terram caliginis et tenebrarum,ubi umbra mortis et nullus ordo,sed sempiternus horror inhabitat ".
JOB|11|1|Respondens autem Sophar Naamathites dixit:
JOB|11|2|" Numquid illi, qui multa loquitur, non et respondetur?Aut vir verbosus iustificabitur?
JOB|11|3|Vaniloquium tuum viros tacere faciet,et, cum ceteros irriseris, a nullo confutaberis?
JOB|11|4|Dixisti enim: "Purus est sermo meus,et mundus sum in conspectu tuo".
JOB|11|5|Atque utinam Deus ipse loqueretur tecumet aperiret labia sua tibi,
JOB|11|6|ut ostenderet tibi secreta sapientiaeet arcana consilia eius,et intellegeres quod multo minora quaerat a te,quam meretur iniquitas tua.
JOB|11|7|Forsitan vestigia Dei comprehendeset usque ad perfectum Omnipotentem reperies?
JOB|11|8|Excelsior caelo est, et quid facies?Profundior inferno, et quid cognosces?
JOB|11|9|Longior terra mensura eiuset latior mari.
JOB|11|10|Si subverterit vel concluserit et coarctaverit,quis contradicet ei?
JOB|11|11|Ipse enim novit hominum vanitatem;et videns iniquitatem nonne considerat?
JOB|11|12|Sed et vir vacuus cordatus fit,et homo tamquam pullum onagri nascitur.
JOB|11|13|Tu autem, si cor tuum firmaveriset expanderis ad eum manus tuas,
JOB|11|14|si iniquitatem, quae est in manu tua, abstuleris a te,et non manserit in tabernaculo tuo iniustitia,
JOB|11|15|tunc levare poteris faciem tuam absque maculaet eris stabilis et non timebis.
JOB|11|16|Miseriae quoque oblivisceriset quasi aquarum, quae praeterierunt, recordaberis.
JOB|11|17|Et quasi meridianus fulgor consurget tibi ad vesperam,et, cum te caligine tectum putaveris, orieris ut lucifer.
JOB|11|18|Et habebis fiduciam, proposita tibi spe,et defossus securus dormies.
JOB|11|19|Requiesces, et non erit qui te exterreat;et deprecabuntur faciem tuam plurimi.
JOB|11|20|Oculi autem impiorum deficient,et effugium peribit ab eis;et spes illorum exhalatio animae ".
JOB|12|1|Respondens autem Iob dixit:
JOB|12|2|" Ergo vos estis soli homines,et vobiscum morietur sapientia.
JOB|12|3|Et mihi est cor sicut et vobis,nec inferior vestri sum;quis enim haec, quae nostis, ignorat?
JOB|12|4|Qui deridetur ab amico suo sicut ego,invocabit Deum, et exaudiet eum; deridetur enim iusti integritas.
JOB|12|5|Lampas contempta apud cogitationes eorum, qui securi sunt,parata iis, qui vacillant pede.
JOB|12|6|Tranquilla sunt tabernacula praedonumet secura iis, qui provocant Deum, iis, qui Deum tenent manu sua.
JOB|12|7|Nimirum interroga iumenta, et docebunt te,et volatilia caeli, et indicabunt tibi.
JOB|12|8|Loquere terrae, et docebit te;et narrabunt pisces maris.
JOB|12|9|Quis ignorat in omnibus hisquod manus Domini hoc fecerit?
JOB|12|10|In cuius manu anima omnis viventiset spiritus universae carnis hominis.
JOB|12|11|Nonne auris verba diiudicat,et palatum cibum sibi gustat?
JOB|12|12|In senibus est sapientia,et in longaevis prudentia.
JOB|12|13|Apud ipsum est sapientia et fortitudo;ipse habet consilium et intellegentiam.
JOB|12|14|Si destruxerit, nemo est, qui aedificet;si incluserit hominem, nullus est, qui aperiat.
JOB|12|15|Si continuerit aquas, arescent;et, si emiserit eas, subvertent terram.
JOB|12|16|Apud ipsum est fortitudo et sapientia;ipse novit et decipientem et eum qui decipitur.
JOB|12|17|Inducit consiliarios spoliatoset iudices in stuporem.
JOB|12|18|Balteum regum dissolvitet praecingit fune renes eorum.
JOB|12|19|Inducit sacerdotes spoliatoset optimates supplantat,
JOB|12|20|commutans labium veraciumet doctrinam senum auferens.
JOB|12|21|Effundit despectionem super principeset cingulum fortium relaxat.
JOB|12|22|Qui revelat profunda de tenebriset producit in lucem umbram mortis.
JOB|12|23|Qui multiplicat gentes et perdit easet subversas in integrum restituit.
JOB|12|24|Qui immutat cor principum populi terrae et decipit eoset errare eos faciet per invium desertum.
JOB|12|25|Palpabunt quasi in tenebris et non in luce,et errare eos faciet quasi ebrios.
JOB|13|1|Ecce, omnia haec vidit oculus meus,et audivit auris mea, et intellexi singula.
JOB|13|2|Secundum scientiam vestram, et ego novi;nec inferior vestri sum.
JOB|13|3|Sed tamen ad Omnipotentem loquaret disputare cum Deo cupio;
JOB|13|4|vos autem ostendam fabricatores mendacii,medicos vanos vos omnes.
JOB|13|5|Atque utinam taceretis,ut sit vobis in sapientiam!
JOB|13|6|Audite ergo correptionem meamet contentiones labiorum meorum attendite.
JOB|13|7|Numquid pro Deo profertis mendaciumet pro illo loquimini dolos?
JOB|13|8|Numquid faciem eius accipitiset pro Deo in iudicio contendere nitimini?
JOB|13|9|Aut bonum est quod vos excutiat?Aut, ut illuditur homini, illudetis ei?
JOB|13|10|Ipse vos arguet,cum in abscondito faciem accipitis.
JOB|13|11|Nonne maiestas eius turbabit vos,et terror eius irruet super vos?
JOB|13|12|Sententiae vestrae sunt proverbia cineris;thoraces lutei thoraces vestri.
JOB|13|13|Tacete paulisper, ut loquar ipse,et transeat super me quodcumque.
JOB|13|14|Quare sumam carnes meas dentibus meiset animam meam ponam in manibus meis?
JOB|13|15|Etiamsi occiderit me, in ipso sperabo; verumtamen vias meas in conspectu eius arguam.
JOB|13|16|Et hoc erit salus mea:non enim veniet in conspectu eius omnis impius.
JOB|13|17|Audite sermonem meumet explicationem meam percipite auribus vestris.
JOB|13|18|Ecce iudicium paravi;scio quod iustus inveniar.
JOB|13|19|Quis est qui contendat mecum?Tunc enim tacebo et consummabor.
JOB|13|20|Duo tantum ne facias mihi,et tunc a facie tua non abscondar:
JOB|13|21|Manum tuam longe fac a me,et formido tua non me terreat.
JOB|13|22|Voca me, et ego respondebo tibi;aut ipse loquar, et tu respondebis mihi.
JOB|13|23|Quantas habeo iniquitates et peccata?Scelera mea et delicta ostende mihi.
JOB|13|24|Cur faciem tuam abscondiset arbitraris me inimicum tuum?
JOB|13|25|Contra folium, quod vento rapitur, dure agiset stipulam siccam persequeris.
JOB|13|26|Scribis enim contra me amaritudineset occupatum me vis peccatis adulescentiae meae.
JOB|13|27|Posuisti in nervo pedem meumet observasti omnes semitas measet vestigia pedum meorum considerasti.
JOB|13|28|Qui quasi uter consumendus sum,et quasi vestimentum, quod comeditur a tinea.
JOB|14|1|Homo natus de muliere,brevi vivens tempore, commotione satiatur.
JOB|14|2|Qui quasi flos egreditur et arescitet fugit velut umbra et non permanet.
JOB|14|3|Et dignum ducis super huiuscemodi aperire oculos tuoset adducere eum tecum in iudicium?
JOB|14|4|Quis potest facere mundum de immundo?Ne unus quidem!
JOB|14|5|Si statuti dies hominis sunt,et numerus mensium eius apud te est,et constituti sunt termini eius, quos non praeteribit,
JOB|14|6|averte oculos tuos ab eo, ut quiescat,donec solvat, sicut mercennarius, dies suos.
JOB|14|7|Nam lignum habet spem;si praecisum fuerit, rursum virescet,et rami eius non deficient.
JOB|14|8|Si senuerit in terra radix eius,et in pulvere emortuus fuerit truncus illius,
JOB|14|9|ad odorem aquae germinabitet faciet comam quasi novellae.
JOB|14|10|Homo vero cum mortuus fuerit et debilitatur,exspirat homo et, ubi, quaeso, est?
JOB|14|11|Recedent aquae de mari,et fluvius vacuefactus arescet;
JOB|14|12|sic homo, cum dormierit, non resurget:donec atteratur caelum, non evigilabitnec consurget de somno suo.
JOB|14|13|Quis mihi hoc tribuat, ut in inferno seponas meet abscondas me, donec pertranseat furor tuus,et constituas mihi tempus, in quo recorderis mei?
JOB|14|14|Putasne mortuus homo rursum vivat?Cunctis diebus, quibus nunc milito,exspectarem, donec veniat immutatio mea.
JOB|14|15|Vocares me, et ego responderem tibi;opus manuum tuarum requireres.
JOB|14|16|Tu quidem nunc gressus meos dinumerares,sed parceres peccatis meis.
JOB|14|17|Signares quasi in sacculo delicta mea,sed dealbares iniquitatem meam.
JOB|14|18|Mons cadens decidit,et saxum transfertur de loco suo;
JOB|14|19|lapides excavant aquae,et alluvione terra inundatur:et spem hominis perdes.
JOB|14|20|Praevales adversus eum, et in perpetuum transiet;immutas faciem eius et emittis eum.
JOB|14|21|Sive nobiles fuerint filii eius, non novit;sive ignobiles, non intellegit.
JOB|14|22|Attamen caro eius, dum vivet, dolet,et anima illius super semetipso luget ".
JOB|15|1|Respondens autem Eliphaz Themanites dixit:
JOB|15|2|" Numquid sapiens respondebit sapientia ventosaet implebit vento urente stomachum suum?
JOB|15|3|Arguens verbis, quae nihil prosunt,et sententiis, quae nihil iuvant?
JOB|15|4|Tu autem pietatem dissolviset detrahis meditationi coram Deo.
JOB|15|5|Docet enim iniquitas tua os tuum,et assumis linguam callidorum.
JOB|15|6|Condemnabit te os tuum et non ego,et labia tua respondebunt tibi.
JOB|15|7|Numquid primus homo tu natus eset ante colles formatus?
JOB|15|8|Numquid consilium Dei audistiet tibi attrahis sapientiam?
JOB|15|9|Quid nosti, quod nos ignoremus?Quid intellegis, quod nos nesciamus?
JOB|15|10|Et senes et antiqui sunt inter nos,multo vetustiores quam pater tuus.
JOB|15|11|Numquid parum tibi sunt consolationes Dei?Et verbum lene tecum factum?
JOB|15|12|Quid te elevat cor tuum,et cur attonitos habes oculos?
JOB|15|13|Quid vertis contra Deum spiritum tuumet profers de ore tuo huiuscemodi sermones?
JOB|15|14|Quid est homo, ut immaculatus sit,et ut iustus appareat natus de muliere?
JOB|15|15|Ecce, sanctis suis non fidit,et caeli non sunt mundi in conspectu eius;
JOB|15|16|quanto magis abominabilis et corruptus homo,qui bibit quasi aquam iniquitatem.
JOB|15|17|Ostendam tibi, audi me;quod vidi, narrabo tibi,
JOB|15|18|quod sapientes confitentur,et non celaverunt eos patres eorum:
JOB|15|19|quibus solis data est terra,et non transivit alienus per eos.
JOB|15|20|Cunctis diebus suis impius cruciatur,et numerus annorum incertus est tyranno.
JOB|15|21|Sonitus terroris semper in auribus illius,quasi, cum pax sit, vastator irruat in eum.
JOB|15|22|Non credit quod reverti possit de tenebris,cum sit destinatus gladio.
JOB|15|23|Cum se moverit ad quaerendum panem: "Ubinam?",novit quod paratus sit in manu eius tenebrarum dies.
JOB|15|24|Terrebit eum tribulatio et angustia,vallabit eum sicut regem, qui praeparatur ad proelium.
JOB|15|25|Tetendit enim adversus Deum manum suam,et contra Omnipotentem roboratus est.
JOB|15|26|Cucurrit adversus eum erecto collo,spisso scuto armatus.
JOB|15|27|Operuit faciem eius crassitudo,et de lateribus eius arvina dependet.
JOB|15|28|Habitavit in civitatibus desolatiset in domibus desertis, quae in tumulos sunt redactae.
JOB|15|29|Non ditabitur, nec perseverabit substantia eius;nec mittet in terra radicem suam.
JOB|15|30|Non recedet de tenebris;ramos eius arefaciet flamma,et auferet ventus florem eius.
JOB|15|31|Ne credat vanitati errore deceptus,quia vanitas erit remuneratio eius.
JOB|15|32|Antequam dies eius impleantur, abscindentur,et ramus eius non virescet.
JOB|15|33|Laedetur quasi vinea in primo flore botrus eius,et quasi oliva proiciens florem suum.
JOB|15|34|Cangregatio enim impii sterilis,et ignis devorabit tabernacula eorum, qui munera libenter accipiunt.
JOB|15|35|Concepit dolorem et peperit iniquitatem,et venter eius praeparat dolos.
JOB|16|1|Respondens autem Iob dixit:
JOB|16|2|" Audivi frequenter talia!onsolatores molesti omnes vos estis.
JOB|16|3|Numquid habebunt finem verba ventosa,aut quid te exacerbat, ut respondeas?
JOB|16|4|Poteram et ego similia vestri loqui,si esset anima vestra pro anima mea!Concinnarem super vos sermoneset moverem caput meum super vos.
JOB|16|5|Roborarem vos ore meoet motum labiorum meorum non cohiberem.
JOB|16|6|Si locutus fuero, non quiescet dolor meuset, si tacuero, non recedet a me;
JOB|16|7|nunc autem defatigavit me dolor meus,et tu vastasti omnem coetum meum.
JOB|16|8|Rugae meae testimonium dicunt contra me;et suscitatur falsiloquus adversus faciem meam contradicens mihi,
JOB|16|9|Ira eius discerpsit me et adversata est mihi,et infremuit contra me dentibus suis.Hostis meus acuit oculos suos in me.
JOB|16|10|Aperuerunt super me ora suaet exprobrantes percusserunt maxillam meam,simul conferti contra me.
JOB|16|11|Concludit me Deus apud iniquumet manibus impiorum me tradit.
JOB|16|12|Ego, ille quondam tranquillus, repente contritus sum.Tenuit cervicem meam, confregit meet posuit me sibi quasi in signum.
JOB|16|13|Circumdedit me lanceis suis,scidit lumbos meos, non pepercitet effudit in terra iecur meum.
JOB|16|14|Dirupit me rumpens et diruens,irruit in me quasi gigas.
JOB|16|15|Saccum consui super cutem meamet dimisi in terram cornu meum.
JOB|16|16|Facies mea rubuit a fletu,et palpebrae meae caligaverunt;
JOB|16|17|attamen absque iniquitate manus meae,cum haberem mundas preces.
JOB|16|18|Terra, ne operias sanguinem meum,neque inveniat in te locum latendi clamor meus.
JOB|16|19|Ecce enim in caelo testis meus,et conscius meus in excelsis.
JOB|16|20|Interpretes mei sunt cogitationes meae:ad Deum stillat oculus meus.
JOB|16|21|Atque utinam sic iudicaretur vir cum Deo,sicut iudicatur filius hominis cum collega suo.
JOB|16|22|Ecce enim breves anni transeunt,et semitam, per quam non revertar, ambulo.
JOB|17|1|Spiritus meus attenuatus est,dies mei exstincti,et solum mihi superest sepulcrum.
JOB|17|2|Nonne irrisiones circumdant me,et in amaritudinibus moratur oculus meus?
JOB|17|3|Pone pignus pro me iuxta te;et quis umquam spondens percutiet manum meam?
JOB|17|4|Cor eorum longe fecisti a disciplina;propterea non exaltabuntur.
JOB|17|5|Praedam pollicetur sociis,sed oculi filiorum eius deficient.
JOB|17|6|Posuit me quasi in proverbium vulgiet conspuendum in faciem.
JOB|17|7|Caligavit ab indignatione oculus meus,et membra mea quasi in umbram redacta sunt.
JOB|17|8|Stupebunt iusti super hoc,et innocens contra impium excitabitur.
JOB|17|9|Et tenebit iustus viam suam,et mundus manibus addet fortitudinem.
JOB|17|10|Igitur omnes vos convertimini et venite,et non inveniam in vobis ullum sapientem.
JOB|17|11|Dies mei transierunt, cogitationes meae dissipatae suntet desideria cordis mei.
JOB|17|12|Noctem verterunt in diem;et rursum post tenebras properat lux.
JOB|17|13|Si sustinuero, infernus domus mea est;et in tenebris stravi lectulum meum.
JOB|17|14|Putredini dixi: Pater meus es!;Mater mea et soror mea! vermibus.
JOB|17|15|Ubi est ergo nunc praestolatio mea,et patientiam meam quis considerat?
JOB|17|16|In profundissimum infernum descendent omnia mea;simul in pulvere erit requies mihi? ".
JOB|18|1|Respondens autem Baldad Suhites dixit:
JOB|18|2|" Usque ad quem finem verba iactabitis?Intellegite prius, et sic loquamur.
JOB|18|3|Quare reputati sumus ut iumentaet sorduimus coram vobis?
JOB|18|4|Qui perdis animam tuam in furore tuo,numquid propter te derelinquetur terra,et transferentur rupes de loco suo?
JOB|18|5|Etenim lux impii exstinguetur,nec splendebit flamma ignis eius.
JOB|18|6|Lux obtenebrescet in tabernaculo illius,et lucerna, quae super eum est, exstinguetur.
JOB|18|7|Arctabuntur gressus virtutis eius,et praecipitabit eum consilium suum.
JOB|18|8|Immissi sunt in rete pedes eius,et in reticulo ambulat.
JOB|18|9|Tenet plantam illius laqueus,et firmatur super eum tendiculum.
JOB|18|10|Abscondita est in terra pedica eius,et decipula illius super semitam.
JOB|18|11|Undique terrent eum formidineset involvunt pedes eius.
JOB|18|12|Attenuatur fame robur eius,et pernicies parata costis illius.
JOB|18|13|Devorat partes cutis eius,consumat membra illius primogenitus mortis.
JOB|18|14|Avellitur de tabernaculo suo fiducia eius,et urges eum ad regem formidinum.
JOB|18|15|Habitas in tabernaculo, quod iam non est ei;aspergitur in habitatione eius sulphur.
JOB|18|16|Deorsum radices eius siccantur,sursum autem atteruntur rami eius.
JOB|18|17|Memoria illius periit de terra,et non celebrabitur nomen eius in plateis.
JOB|18|18|Expellent eum de luce in tenebraset de orbe transferent eum.
JOB|18|19|Non erit semen eius neque progenies in populo suo,nec ullae reliquiae in commoratione eius.
JOB|18|20|In die eius stupebunt novissimi,et primos invadet horror.
JOB|18|21|Haec sunt ergo tabernacula iniqui;et iste locus eius, qui ignorat Deum ".
JOB|19|1|Respondens autem Iob dixit:
JOB|19|2|" Usquequo affligitis ani mam meamet atteritis me sermonibus?
JOB|19|3|En decies obiurgatis meet non erubescitis opprimentes me.
JOB|19|4|Nempe, etsi erravi,mecum erit error meus.
JOB|19|5|Si vos contra me erigiminiet arguitis me opprobriis meis,
JOB|19|6|saltem nunc intellegite quia Deus non aequo iudicio afflixerit meet rete suo me cinxerit.
JOB|19|7|Etsi clamo: Vim patior!, non exaudior;si vociferor, non est qui iudicet.
JOB|19|8|Semitam meam circumsaepsit, et transire non possum;et in calle meo tenebras posuit.
JOB|19|9|Spoliavit me gloria meaet abstulit coronam de capite meo.
JOB|19|10|Destruxit me undique, et pereo,et evellit quasi arborem spem meam.
JOB|19|11|Iratus est contra me furor eius,et sic me habuit quasi hostem suum.
JOB|19|12|Simul venerunt turmae eiuset fecerunt sibi viam adversus meet obsederunt in gyro tabernaculum meum.
JOB|19|13|Fratres meos longe fecit a me,et noti mei quasi alieni recesserunt a me.
JOB|19|14|Dereliquerunt me propinqui mei,et, qui me noverant, obliti sunt mei.
JOB|19|15|Inquilini domus meae et ancillae meae sicut alienum habuerunt me,et quasi peregrinus fui in oculis eorum.
JOB|19|16|Servum meum vocavi, et non respondit;ore proprio deprecabar illum.
JOB|19|17|Halitum meum exhorruit uxor mea,et fetui filiis uteri mei.
JOB|19|18|Vel infantes despiciebant meet, cum surgerem, detrahebant mihi.
JOB|19|19|Abominati sunt me quondam consiliarii mei;et, quem maxime diligebam, aversatus est me.
JOB|19|20|Pelli meae, consumptis carnibus, adhaesit os meum,et evanuit cutis mea circa dentes meos.
JOB|19|21|Miseremini mei, miseremini mei, saltem vos, amici mei,quia manus Domini tetigit me.
JOB|19|22|Quare persequimini me sicut Deuset carnibus meis non saturamini?
JOB|19|23|Quis mihi tribuat, ut scribantur sermones mei?Quis mihi det, ut exarentur in libro
JOB|19|24|stilo ferreo et plumbeo,in aeternum sculpantur in silice?
JOB|19|25|Scio enim quod redemptor meus vivitet in novissimo super pulvere stabit;
JOB|19|26|et post pellem meam hanc, quam abstraxerunt,et de carne mea videbo Deum.
JOB|19|27|Quem visurus sum ego ipse,et oculi mei conspecturi sunt, et non alienum.Consumpti sunt renes mei in sinu meo.
JOB|19|28|Si ergo nunc dicitis: "Quomodo persequemur eumet radicem verbi inveniemus contra eum?",
JOB|19|29|timete a facie gladii,quoniam ultor iniquitatum gladius est;et scitote esse iudicium ".
JOB|20|1|Respondens autem Sophar Naamathites dixit:
JOB|20|2|" Idcirco cogitationes meae reducunt me,eo quod intellectus effulsit in me.
JOB|20|3|Doctrinam, qua me arguis, audiam,at spiritus intellegentiae meae respondebit mihi.
JOB|20|4|Scisne hoc a principio,ex quo positus est homo super terram,
JOB|20|5|quod exsultatio iniquorum brevis sit,et gaudium impiorum ad instar puncti?
JOB|20|6|si ascenderit usque ad caelum superbia eius,et caput eius nubes tetigerit,
JOB|20|7|quasi sterquilinium in finem perdetur,et, qui eum viderant, dicent: "Ubi est?".
JOB|20|8|Velut somnium avolans non invenietur,transiet sicut visio nocturna.
JOB|20|9|Oculus, qui eum viderat, non videbit,neque ultra intuebitur eum locus suus.
JOB|20|10|Filii eius satagent complacere pauperibus,et manus illius reddent ei possessionem suam.
JOB|20|11|Ossa eius, quae implebantur adulescentia,cum eo in pulvere dormient.
JOB|20|12|Cum enim dulce fuerit in ore eius malum,abscondet illud sub lingua sua.
JOB|20|13|Parcet illi et non derelinquet illudet celabit in gutture suo.
JOB|20|14|Panis eius in visceribus illiusvertetur in fel aspidum intrinsecus.
JOB|20|15|Divitias, quas devoravit, evomet,et de ventre illius extrahet eas Deus.
JOB|20|16|Venenum aspidum sugebat,et occidet eum lingua viperae.
JOB|20|17|Non videat rivulos olei,torrentes mellis et butyri.
JOB|20|18|Restituet quaestum suum nec deglutiet,de opibus venditionum non laetabitur.
JOB|20|19|Quoniam confringens deseruit pauperes,domum rapuit et non aedificavit eam.
JOB|20|20|Nec est satiatus venter eius;et cum desideriis suis evadere non potuit.
JOB|20|21|Non fuerunt reliquiae de cibo eius,et propterea nihil permanebit de bonis eius.
JOB|20|22|Cum satiatus fuerit, arctabitur;et omnis dolor irruet super eum.
JOB|20|23|Impleat ventrem suum:emittet Deus in eum iram furoris suiet pluet super illum bellum suum.
JOB|20|24|Fugiet arma ferreaet irruet in arcum aereum.
JOB|20|25|Sagitta transverberabit corpus eius,et fulgur iecur eius;vadent et venient super eum horribilia.
JOB|20|26|Omnes tenebrae absconditae sunt in occultis eius,devorabit eum ignis, qui non succenditur;affligetur relictus in tabernaculo suo.
JOB|20|27|Revelabunt caeli iniquitatem eius,et terra consurget adversus eum.
JOB|20|28|Auferetur germen domus illius,detrahetur in die furoris Dei.
JOB|20|29|Haec est pars hominis impii a Deo,et hereditas verborum eius a Domino ".
JOB|21|1|Respondens autem Iob dixit:
JOB|21|2|" Audite, quaeso, sermonesmeos,et sint haec consolationes vestrae.
JOB|21|3|Sustinete me, et ego loquar;et post verba mea ridebitis.
JOB|21|4|Numquid contra hominem disputatio mea est,ut merito non debeam impatiens fieri?
JOB|21|5|Attendite me et obstupesciteet superponite digitum ori vestro.
JOB|21|6|Et ego, quando recordatus fuero, pertimesco,et concutit carnem meam tremor.
JOB|21|7|Quare ergo impii vivunt,senuerunt confortatique sunt divitiis?
JOB|21|8|Semen eorum permanet coram eis,et progenies eorum in conspectu eorum.
JOB|21|9|Domus eorum securae sunt et pacatae,et non est virga Dei super illos.
JOB|21|10|Bos eorum concepit et non abortivit,vacca peperit et non est privata fetu suo.
JOB|21|11|Egrediuntur quasi greges parvuli eorum,et infantes eorum exsultant lusibus.
JOB|21|12|Tenent tympanum et citharamet gaudent ad sonitum organi.
JOB|21|13|Ducunt in bonis dies suoset in puncto ad inferna descendunt.
JOB|21|14|Qui dixerant Deo: "Recede a nobis!Scientiam viarum tuarum nolumus.
JOB|21|15|Quis est Omnipotens, ut serviamus ei,et quid nobis prodest, si oraverimus illum?".
JOB|21|16|Sint in manu eorum bona sua;consilium vero impiorum longe sit a me.
JOB|21|17|Quam saepe lucerna impiorum exstinguitur,et superveniet eis pernicies,et dolores dividet in furore suo?
JOB|21|18|Erunt sicut paleae ante faciem venti,et sicut favilla, quam turbo dispergit.
JOB|21|19|"Servabitne Deus filiis iniquitatem eius?".Retribuat illi, ut sciat.
JOB|21|20|Videbunt oculi eius interfectionem suam,et de furore Omnipotentis bibet.
JOB|21|21|Quid enim ad eum pertinet de domo sua post se,et si numerus mensium eius recidetur?
JOB|21|22|Numquid Deum docebit quispiam scientiam,qui excelsos iudicat?
JOB|21|23|Iste moritur robustus et sanus,dives et felix;
JOB|21|24|viscera eius plena sunt adipe,et medullis ossa illius irrigantur.
JOB|21|25|Alius vero moritur in amaritudine animaeabsque ullis opibus;
JOB|21|26|et tamen simul in pulvere dormient,et vermes operient eos.
JOB|21|27|Certe novi cogitationes vestraset sententias contra me iniquas.
JOB|21|28|Dicitis enim: "Ubi est domus principis,et ubi tabernacula impiorum?".
JOB|21|29|Nonne interrogastis quemlibet de viatoribuset signa eorum non agnovistis?
JOB|21|30|Quia in diem perditionis servatur maluset ad diem furoris abducetur.
JOB|21|31|Quis arguet coram eo viam eius,et, quae fecit, quis reddet illi?
JOB|21|32|Ipse ad sepulcra ducetur,et super tumulum vigilabunt.
JOB|21|33|Dulces erunt ei glebae vallis,et post se omnem hominem trahetet ante se innumerabiles.
JOB|21|34|Quomodo igitur consolamini me frustra,et responsionis vestrae restat perfidia? ".
JOB|22|1|Respondens autem Eliphaz Themanites dixit:
JOB|22|2|" Numquid Deo prodesse potest homo,cum vix intellegens sibi ipse proderit?
JOB|22|3|Quid prodest Omnipotenti, si iustus fueris,aut quid ei confers, si immaculatam feceris viam tuam?
JOB|22|4|Numquid pro tua pietate arguet teet veniet tecum in iudicium?
JOB|22|5|Et non propter malitiam tuam plurimamet infinitas iniquitates tuas?
JOB|22|6|Sumpsisti enim pignori fratres tuos sine causaet nudos spoliasti vestibus.
JOB|22|7|Aquam lasso non dedistiet esurienti cohibuisti panem.
JOB|22|8|Numquid viro forti brachio erit terra,et acceptus sedebit in ea?
JOB|22|9|Viduas dimisisti vacuaset lacertos pupillorum comminuisti.
JOB|22|10|Propterea circumdatus es laqueis,et conturbat te subita formido.
JOB|22|11|Vel tenebras non vides,et impetus aquarum opprimit te.
JOB|22|12|"Nonne Deus excelsior caelo?Et inspice stellarum verticem: quam sublimis!".
JOB|22|13|Et dicis: "Quid enim novit Deuset quasi per caliginem iudicat?
JOB|22|14|Nubes latibulum eius, nec nostra considerat;et circa orbem caeli perambulat".
JOB|22|15|Numquid semitam saeculorum custodire cupis,quam calcaverunt viri iniqui?
JOB|22|16|Qui sublati ante tempus suum,et fluvius subvertit fundamentum eorum.
JOB|22|17|Qui dicebant Deo: "Recede a nobis!"et "Quid faciet Omnipotens nobis?".
JOB|22|18|Cum ille implesset domos eorum bonis,quorum sententia procul erat ab eo.
JOB|22|19|Videbunt iusti et laetabuntur,et innocens subsannabit eos:
JOB|22|20|"Vere succisus est status eorum,et reliquias eorum devoravit ignis".
JOB|22|21|Acquiesce igitur ei, et habeto pacem;et per haec habebis fructus optimos.
JOB|22|22|Suscipe ex ore illius legemet pone sermones eius in corde tuo.
JOB|22|23|Si reversus fueris ad Omnipotentem, aedificaberiset longe facies iniquitatem a tabernaculo tuo.
JOB|22|24|Comparabis tamquam terram aurumet tamquam glaream torrentis Ophir.
JOB|22|25|Eritque Omnipotens metallum tuum,et argentum coacervabitur tibi.
JOB|22|26|Tunc super Omnipotentem deliciis afflueset elevabis ad Deum faciem tuam.
JOB|22|27|Supplex rogabis eum, et exaudiet te,et vota tua reddes.
JOB|22|28|Decernes rem, et veniet tibi,et in viis tuis splendebit lumen.
JOB|22|29|Quia humiliat eum, qui loquitur superba,et demissus oculis ipse salvabitur.
JOB|22|30|Eripiet innocentem,eripietur autem in munditia manuum suarum ".
JOB|23|1|Respondens autem Iob ait:
JOB|23|2|" Nunc quoque in amaritu tudine est querela mea,et manus eius aggravata est super gemitum meum.
JOB|23|3|Quis mihi tribuat, ut cognoscam et inveniam illumet veniam usque ad solium eius?
JOB|23|4|Ponam coram eo iudiciumet os meum replebo increpationibus,
JOB|23|5|ut sciam verba, quae mihi respondeat,et intellegam quid loquatur mihi.
JOB|23|6|Num multa fortitudine contendet mecum?Non! Ipse tantum audiat!
JOB|23|7|Tunc iustus disceptabit cum illo,et ego evaderem in perpetuo a iudice meo.
JOB|23|8|Si ad orientem iero, non apparet;si ad occidentem, non intellegam eum.
JOB|23|9|Si ad sinistram pergam, non apprehendam eum;si me vertam ad dexteram, non videbo illum.
JOB|23|10|Ipse vero scit viam meam,et, si probaverit me, quasi aurum egrediar.
JOB|23|11|Vestigia eius secutus est pes meus,viam eius custodivi et non declinavi ex ea.
JOB|23|12|A mandatis labiorum eius non recessiet in sinu meo abscondi verba oris eius.
JOB|23|13|Ipse enim solus est, et quis repellet eum?Et anima eius, quodcumque voluit, hoc fecit.
JOB|23|14|Cum expleverit in me voluntatem suam,et alia multa similia praesto sunt ei;
JOB|23|15|et idcirco a facie eius turbatus sumet considerans eum timore sollicitor.
JOB|23|16|Deus mollivit cor meum,et Omnipotens conturbavit me.
JOB|23|17|Non enim perii propter imminentes tenebras,nec faciem meam operuit caligo.
JOB|24|1|Cur ab Omnipotente non sunt abscondita tempora,qui autem noverunt eum, ignorant dies illius?
JOB|24|2|Alii terminos transtulerunt,diripuerunt greges et paverunt eos.
JOB|24|3|Asinum pupillorum abegeruntet abstulerunt pro pignore bovem viduae.
JOB|24|4|Subverterunt pauperum viam,et simul se occultare coacti sunt mansueti terrae.
JOB|24|5|Alii, quasi onagri in deserto,egrediuntur ad opus suum:vigilantes ad praedamin terra arida ad panem liberis.
JOB|24|6|Agrum non suum demetuntet vineam peccatoris vindemiant.
JOB|24|7|Nudi pernoctant sine indumento,nec est eis operimentum in frigore.
JOB|24|8|Imbre montium riganturet non habentes refugium adhaerent rupibus.
JOB|24|9|Abripuerunt pupillum ab ubereet pauperem pignori sumpserunt;
JOB|24|10|nudi et incedentes absque vestituet esurientes portant spicas.
JOB|24|11|Inter muros oleum expresseruntet calcatis torcularibus sitiunt.
JOB|24|12|De civitatibus morientes ingemuerunt,et anima vulneratorum clamavit,et Deus non ponit aurem ad precem.
JOB|24|13|Ipsi fuerunt rebelles lumini,nescierunt vias eiusnec morati sunt in semitis eius.
JOB|24|14|Mane primo consurgit homicida,interficit egenum et pauperem;per noctem vero erit quasi fur.
JOB|24|15|Oculus adulteri observat caliginemdicens: "Non me videbit oculus";et operiet vultum suum.
JOB|24|16|Perfodit in tenebris domos, interdiu sese abdideruntet ignoraverunt lucem.
JOB|24|17|Si subito apparuerit aurora, arbitrantur umbram mortis,nam sunt assueti terroribus umbrae mortis.
JOB|24|18|"Levis est super faciem aquae;maledicta est pars eius in terra,nec est qui se dirigat ad vineas eius.
JOB|24|19|Siccitas et calor abstulerunt aquas nivium,et inferi eos, qui peccaverunt.
JOB|24|20|Sinus matris obliviscatur eius,dulcedo illius vermes fiant;non sit in recordatione,sed conteratur quasi lignum iniquitas.
JOB|24|21|Male egit cum sterili, quae non parit,et viduae bene non fecit.
JOB|24|22|Detraxit fortes in fortitudine suaet, cum steterit, ille non credet vitae suae.
JOB|24|23|Dedit ei locum securitatis, quo sustentetur;oculi autem eius sunt in viis illius.
JOB|24|24|Elevati sunt ad modicum et non subsistent,et humiliabuntur sicut omnia et auferenturet sicut summitates spicarum conterentur".
JOB|24|25|Quod si non est ita, quis me potest arguere esse mentitumet ponere in nihilum verba mea? ".
JOB|25|1|Respondens autem Baldad Suhites dixit:
JOB|25|2|" Potestas et terror apud eum est,qui facit pacem in sublimibus suis.
JOB|25|3|Numquid est numerus militum eius?Et super quem non surget lumen illius?
JOB|25|4|Numquid iustificari potest homo comparatus Deo,aut apparere mundus natus de muliere?
JOB|25|5|Ecce luna etiam non splendet,et stellae non sunt mundae in conspectu eius;
JOB|25|6|quanto magis homo putredo,et filius hominis vermis ".
JOB|26|1|Respondens autem Iob dixit:
JOB|26|2|" Quomodo adiuvisti imbecillem?Et sustentas brachium eius, qui non est fortis?
JOB|26|3|Quod dedisti illi consilium, qui non habet sapientiam?Et prudentiam tuam ostendisti plurimam!
JOB|26|4|Quem docere voluisti?Et cuius est spiritus, qui egreditur ex te?
JOB|26|5|Ecce umbrae gemunt sub aquis,et qui habitant cum eis.
JOB|26|6|Nudus est infernus coram illo,et nullum est operimentum Perditioni.
JOB|26|7|Qui extendit aquilonem super vacuumet appendit terram super nihilum.
JOB|26|8|Qui ligat aquas in nubibus suis,ut non erumpant pariter deorsum.
JOB|26|9|Qui operit faciem solii suiexpandens super illud nebulam suam.
JOB|26|10|Terminum circumdedit aquis,usque dum finiantur lux et tenebrae.
JOB|26|11|Columnae caeli contremiscuntet pavent ab increpatione eius.
JOB|26|12|In fortitudine sua terruit mareet prudentia sua percussit Rahab.
JOB|26|13|Spiritus eius serenavit caelos,et manus eius confodit colubrum fugientem.
JOB|26|14|Ecce haec sunt termini viarum eius;et, cum vix parvam stillam sermonis eius audierimus,quis poterit tonitruum magnitudinis illius intueri? ".
JOB|27|1|Addidit quoque Iob assu mens parabolam suam et dixit:
JOB|27|2|" Vivit Deus, qui abstulit ius meum, et Omnipotens, qui ad amaritudinem adduxit animam meam,
JOB|27|3|quia, donec superest halitus in me,et spiritus Dei in naribus meis,
JOB|27|4|non loquentur labia mea iniquitatem,nec lingua mea meditabitur mendacium!
JOB|27|5|Absit a me, ut iustos vos esse iudicem;donec exspirem, non recedam ab innocentia mea.
JOB|27|6|Iustificationem meam, quam coepi tenere, non deseram,neque enim reprehendit me cor meum in omni vita mea.
JOB|27|7|Sit ut impius inimicus meus,et adversarius meus quasi iniquus.
JOB|27|8|Quae est enim spes impii, cum secet,cum rapiat Deus animam eius?
JOB|27|9|Numquid Deus audiet clamorem eius,cum venerit super eum angustia?
JOB|27|10|Aut poterit in Omnipotente delectariet invocare Deum omni tempore?
JOB|27|11|Docebo vos manum Dei,quae Omnipotens habeat, nec abscondam.
JOB|27|12|Ecce vos omnes observastis,et quid sine causa vana loquimini?
JOB|27|13|Haec est pars hominis impii apud Deum,et hereditas violentorum, quam ab Omnipotente suscipient.
JOB|27|14|Si multiplicati fuerint filii eius, in gladio erunt,et nepotes eius non saturabuntur pane.
JOB|27|15|Qui reliqui fuerint ex eo, sepelientur in interitu,et viduae illius non plorabunt.
JOB|27|16|Si comportaverit quasi terram argentumet sicut lutum praeparaverit vestimenta,
JOB|27|17|praeparabit quidem, sed iustus vestietur illis,et argentum innocens dividet.
JOB|27|18|Aedificavit sicut aranea domum suam,et sicut custos fecit umbraculum.
JOB|27|19|Dives, cum dormierit, nihil secum auferet;aperiet oculos suos et nihil inveniet.
JOB|27|20|Apprehendet eum quasi aqua inopia,nocte opprimet eum tempestas.
JOB|27|21|Tollet eum ventus urens et auferet,et velut turbo rapiet eum de loco suo.
JOB|27|22|Et mittet super eum et non parcet;de manu eius fugiens fugiet.
JOB|27|23|Complodet super eum manus suaset sibilabit eum de loco suo.
JOB|28|1|Habet argentum venarum principiaet auro locus est, in quo conflatur.
JOB|28|2|Ferrum de terra tollitur,et lapis solutus calore in aes vertitur.
JOB|28|3|Terminum posuit tenebriset universorum finem ipse scrutatur,lapidem quoque caliginis et umbrae.
JOB|28|4|Aperuit cuniculos gens peregrina,ipsique obliti sunt pedes,penduli haerent plus quam vir nutans.
JOB|28|5|Terra, de qua oriebatur panis,in profundo subversa est sicut per ignem.
JOB|28|6|Locus sapphiri lapides eius,et glebae illius aurum.
JOB|28|7|Semitam ignoravit avis rapax,nec intuitus est eam oculus vulturis.
JOB|28|8|Non calcaverunt eam filii superbiae,nec pertransivit per eam leaena.
JOB|28|9|Ad silicem extendit manum suam,subvertit a radicibus montes.
JOB|28|10|In petris canales excidit,et omne pretiosum vidit oculus eius.
JOB|28|11|Profunda quoque fluviorum scrutatus estet abscondita in lucem produxit.
JOB|28|12|Sapientia vero ubi invenitur?Et quis est locus intellegentiae?
JOB|28|13|Nescit homo structuram eius,nec invenitur in terra viventium.
JOB|28|14|Abyssus dicit: "Non est in me";et mare loquitur: "Non est mecum".
JOB|28|15|Non dabitur aurum obryzum pro ea,nec appendetur argentum in commutatione eius.
JOB|28|16|Non appendetur auro Ophirnec lapidi sardonycho pretiosissimo vel sapphiro.
JOB|28|17|Non adaequabitur ei aurum vel vitrum,nec commutabuntur pro ea vasa auri.
JOB|28|18|Corallia et crystallum non memorabuntur comparatione eius;et possessio sapientiae potior margaritis.
JOB|28|19|Non adaequabitur ei topazius de Aethiopianec auro mundissimo componetur.
JOB|28|20|Unde ergo sapientia venit,et quis est locus intellegentiae?
JOB|28|21|Abscondita est ab oculis omnium viventium,volucres quoque caeli latet.
JOB|28|22|Perditio et mors dixerunt:Auribus nostris audivimus famam eius".
JOB|28|23|Deus intellegit viam eius,et ipse novit locum illius.
JOB|28|24|Ipse enim fines mundi intueturet omnia, quae sub caelo sunt, respicit.
JOB|28|25|Qui fecit ventis ponduset aquas appendit in mensura,
JOB|28|26|quando ponebat pluviis legemet viam procellis sonantibus,
JOB|28|27|tunc vidit illam et enarravitet praeparavit et investigavit.
JOB|28|28|Et dixit homini: "Ecce timor Domini, ipsa est sapientia;et recedere a malo intellegentia" ".
JOB|29|1|Addidit quoque Iob assumens parabolam suam et di xit:
JOB|29|2|" Quis mihi tribuat, ut sim iuxta menses pristinos,secundum dies, quibus Deus custodiebat me?
JOB|29|3|Quando splendebat lucerna eius super caput meum,et ad lumen eius ambulabam in tenebris.
JOB|29|4|Sicut fui in diebus adulescentiae meae,quando familiaris Deus erat in tabernaculo meo,
JOB|29|5|quando erat Omnipotens mecum,et in circuitu meo pueri mei,
JOB|29|6|quando lavabam pedes meos lacte,et petra fundebat mihi rivos olei.
JOB|29|7|Quando procedebam ad portam civitatiset in platea parabam cathedram mihi,
JOB|29|8|videbant me iuvenes et abscondebantur,et senes assurgentes stabant.
JOB|29|9|Principes cessabant loquiet digitum superponebant ori suo.
JOB|29|10|Vocem suam cohibebant duces,et lingua eorum palato suo adhaerebat.
JOB|29|11|Auris audiens beatificabat me,et oculus videns testimonium reddebat mihi,
JOB|29|12|eo quod liberassem pauperem vociferantemet pupillum, cui non esset adiutor.
JOB|29|13|Benedictio perituri super me veniebat,et cor viduae iubilare feci.
JOB|29|14|Iustitia indutus sum et vestivi me,sicut vestimento et diademate, iudicio meo.
JOB|29|15|Oculus fui caecoet pes claudo;
JOB|29|16|pater eram pauperumet causam viri ignoti diligentissime investigabam.
JOB|29|17|Conterebam molas iniquiet de dentibus illius auferebam praedam.
JOB|29|18|Dicebamque: In nidulo meo moriaret sicut palma multiplicabo dies.
JOB|29|19|Radix mea aperta est secus aquas,et ros morabitur in ramis meis.
JOB|29|20|Gloria mea semper innovabitur,et arcus meus in manu mea instaurabitur.
JOB|29|21|Qui me audiebant, blandiebanturet intenti tacebant ad consilium meum.
JOB|29|22|Verbis meis addere nihil audebant,et super illos stillabat eloquium meum.
JOB|29|23|Exspectabant me sicut pluviamet os suum aperiebant quasi ad imbrem serotinum.
JOB|29|24|Si quando ridebam ad eos, non credebant,et lux vultus mei non cadebat in terram.
JOB|29|25|Si voluissem ire ad eos, sedebam primus;cumque sederem quasi rex, circumstante exercitu,eram tamen maerentium consolator.
JOB|30|1|Nunc autem derident meiuniores tempore,quorum non dignabar patresponere cum canibus gregis mei;
JOB|30|2|quorum virtus manuum mihi erat pro nihilo,et robur iuvenile perierat totum.
JOB|30|3|Egestate et fame steriles, qui rodebant in solitudine,serotino tempore fiebant turbo et vastatio;
JOB|30|4|et mandebant herbas et arborum frutices,et radix iuniperorum erat cibus eorum.
JOB|30|5|De medio eiciebantur,clamabant contra eos tamquam fures;
JOB|30|6|ad ripas habitabant torrentiumet in cavernis terrae et petrarum;
JOB|30|7|inter frutices rudebant,sub sentibus se congerebant;
JOB|30|8|filii stultorum et ignobiliumet de terra penitus exturbati.
JOB|30|9|Nunc in eorum canticum versus sumet factus sum eis in proverbium.
JOB|30|10|Abominantur me et longe fugiunt a meet faciem meam conspuere non verentur.
JOB|30|11|Pharetram enim suam aperuit et afflixit meet frenum in os meum immisit.
JOB|30|12|Ad dexteram progenies surrexerunt;pedes meos subverteruntet complanaverunt contra me semitas ruinae.
JOB|30|13|Dissipaverunt itinera mea,insidiati sunt mihi et praevaluerunt,et non fuit qui ferret auxilium.
JOB|30|14|Quasi rupto muro et aperto irruerunt super meet sub ruinis devoluti sunt.
JOB|30|15|Versi sunt contra me in terrores,persequitur quasi ventus principatum meum,et velut nubes pertransiit salus mea.
JOB|30|16|Nunc autem in memetipso effunditur anima mea;et possident me dies afflictionis.
JOB|30|17|Nocte os meum perforatur doloribus;et, qui me comedunt, non dormiunt.
JOB|30|18|In multitudine roboris tenent vestimentum meumet quasi capitio tunicae succinxerunt me.
JOB|30|19|Proiecit me in lutum,et assimilatus sum favillae et cineri.
JOB|30|20|Clamo ad te, et non exaudis me;sto, et non respicis me.
JOB|30|21|Mutatus es mihi in crudelemet in duritia manus tuae adversaris mihi.
JOB|30|22|Elevasti meet quasi super ventum ponens dissolvisti me.
JOB|30|23|Scio quia morti trades me,ubi constituta est domus omni viventi.
JOB|30|24|Verumtamen non ad ruinam mittit manum;et in exitio eius erit salvatio.
JOB|30|25|An non flebam quondam super eo, qui afflictus erat,et compatiebatur anima mea pauperi?
JOB|30|26|Exspectabam bona, et venerunt mihi mala;praestolabar lucem, et eruperunt tenebrae.
JOB|30|27|Interiora mea efferbuerunt absque ulla requie;praevenerunt me dies afflictionis.
JOB|30|28|Taetro vultu incedebam sine consolatione,consurgens in turba clamabam.
JOB|30|29|Frater fui draconumet socius struthionum.
JOB|30|30|Cutis mea denigrata est super me,et ossa mea aruerunt prae caumate.
JOB|30|31|Versa est in luctum cithara mea,et organum meum in vocem flentium.
JOB|31|1|Pepigi foedus cum oculis meisut ne cogitarem quidem de virgine.
JOB|31|2|Quae enim pars mea apud Deum desuper,et quae hereditas apud Omnipotentem in excelsis?
JOB|31|3|Numquid non perditio est iniquo,et alienatio operantibus iniustitiam?
JOB|31|4|Nonne ipse considerat vias measet cunctos gressus meos dinumerat?
JOB|31|5|Si ambulavi in vanitate,et festinavit in dolo pes meus,
JOB|31|6|appendat me in statera iustaet sciat Deus integritatem meam.
JOB|31|7|Si declinavit gressus meus de via,et si secutum est oculos meos cor meum,et si manibus meis adhaesit macula,
JOB|31|8|seram, et alius comedat,et progenies mea eradicetur.
JOB|31|9|Si deceptum est cor meum super muliere,et si ad ostium amici mei insidiatus sum,
JOB|31|10|molat pro alio uxor mea,et super illam incurventur alii.
JOB|31|11|Hoc enim nefas estet iniquitas iudicialis;
JOB|31|12|ignis est usque ad perditionem devoranset omnia eradicans genimina.
JOB|31|13|Si contempsi subire iudicium cum servo meo et ancilla mea,cum disceptarent adversum me,
JOB|31|14|quid enim faciam, cum surrexerit ad iudicandum Deus;et, cum quaesierit, quid respondebo illi?
JOB|31|15|Numquid non in ventre fecit me,qui et illum operatus est,et formavit me in visceribus unus?
JOB|31|16|Si negavi, quod volebant, pauperibuset oculos viduae languescere feci;
JOB|31|17|si comedi buccellam meam solus,et non comedit pupillus ex ea,
JOB|31|18|quia ab infantia mea educavi eum ut pateret de ventre matris meae direxi eam;
JOB|31|19|si despexi pereuntem, eo quod non habuerit indumentum,et absque operimento pauperem;
JOB|31|20|si non benedixerunt mihi latera eius,et de velleribus ovium mearum calefactus est;
JOB|31|21|si levavi super pupillum manum meam,cum viderem in porta adiutorium mihi,
JOB|31|22|umerus meus a iunctura sua cadat,et brachium meum cum ossibus lacertorum confringatur,
JOB|31|23|quia timor super me calamitas a Deo,et contra maiestatem eius nihil valerem!
JOB|31|24|Si putavi aurum securitatem meamet obryzo dixi: Fiducia mea!;
JOB|31|25|si laetatus sum super multis divitiis meis,et quia plurima repperit manus mea;
JOB|31|26|si vidi solem, cum fulgeret,et lunam incedentem clare,
JOB|31|27|et decepit me in abscondito cor meum,et osculatus sum manum meam ore meo,
JOB|31|28|quae est iniquitas iudicialis,eo quod negassem Deum desuper;
JOB|31|29|si gavisus sum ad ruinam eius, qui me oderat,et exsultavi quod invenisset eum malum,
JOB|31|30|cum non dederim ad peccandum guttur meum,ut expeterem maledicens animam eius;
JOB|31|31|si non dixerunt viri tabernaculi mei: "Quis det, qui de carnibus eius non saturatus sit?";
JOB|31|32|foris non mansit peregrinus,ostium meum viatori patuit;
JOB|31|33|si abscondi quasi homo peccatum meumet celavi in sinu meo iniquitatem meam;
JOB|31|34|si expavi ad multitudinem nimiam,et despectio propinquorum terruit me,et magis tacui nec egressus sum ostium.
JOB|31|35|Quis mihi tribuat auditorem?Ecce signum meum! Omnipotens respondeat mihi!Ecce liber, quem scripsit vir litis meae,
JOB|31|36|ut in umero meo portem illumet alligem illum quasi coronam mihi.
JOB|31|37|Numerum graduum meorum pronuntiabo illiet quasi principem adibo eum.
JOB|31|38|Si adversum me terra mea clamat,et cum ipsa sulci eius deflent;
JOB|31|39|si fructus eius comedi absque pecuniaet animam agricolarum eius afflixi,
JOB|31|40|pro frumento oriatur mihi tribulus,et pro hordeo herba foetida! ".Finita sunt verba Iob.
JOB|32|1|Omiserunt autem tres viri isti respondere Iob, eo quod iustus sibi videretur.
JOB|32|2|Et iratus indignatusque est Eliu filius Barachel Buzites de cognatione Ram; iratus est autem adversum Iob, eo quod iustum se esse diceret coram Deo.
JOB|32|3|Porro adversum amicos eius indignatus est, eo quod non invenissent responsionem, sed tantummodo condemnassent Iob.
JOB|32|4|Igitur Eliu exspectavit Iob loquentem, eo quod seniores essent, qui loquebantur;
JOB|32|5|cum autem vidisset Eliu quod tres respondere non potuissent, iratus est vehementer.
JOB|32|6|Respondensque Eliu filius Barachel Buzites dixit: Iunior sum tempore,vos autem antiquiores;idcirco veritus sum et timuivobis indicare meam sententiam.
JOB|32|7|Dixi: Aetas loquetur,et annorum multitudo docebit sapientiam.
JOB|32|8|Sed, ut video, spiritus est in hominibus,et inspiratio Omnipotentis dat intellegentiam.
JOB|32|9|Non sunt longaevi sapientes,nec senes intellegunt iudicium.
JOB|32|10|Ideo dicam: Audite me,ostendam vobis etiam ego meam sapientiam.
JOB|32|11|Exspectavi enim sermones vestros,intendi aurem in prudentiam vestram, donec investigaretis,
JOB|32|12|et ut vos intellegerem nitebar.Sed, ut video, non est qui possit arguere Iobet respondere ex vobis sermonibus eius.
JOB|32|13|Ne forte dicatis: "Invenimus sapientiam;Deus proiecit eum, non homo".
JOB|32|14|Non parabo mihi verba,et ego non secundum sermones vestros respondebo illi.
JOB|32|15|Extimuerunt nec responderunt ultra;abstuleruntque a se eloquia.
JOB|32|16|Quoniam igitur exspectavi, et non sunt locuti,steterunt, nec ultra responderunt,
JOB|32|17|respondebo et ego partem meamet ostendam scientiam meam.
JOB|32|18|Plenus sum enim sermonibus,et coarctat me spiritus pectoris mei;
JOB|32|19|en venter meus quasi mustum absque spiraculo,quod lagunculas novas disrumpit.
JOB|32|20|Loquar et respirabo paululum,aperiam labia mea et respondebo.
JOB|32|21|Non accipiam personam viriet nulli homini blandiar.
JOB|32|22|Nescio enim blandiri,quia in brevi tolleret me Factor meus.
JOB|33|1|Audi igitur, Iob, eloquia meaet omnes sermones meos ausculta.
JOB|33|2|Ecce aperui os meum,loquatur lingua mea in faucibus meis.
JOB|33|3|Ex recto corde sermones mei sunt,et sententiam puram labia mea loquentur.
JOB|33|4|Spiritus Dei fecit me,et spiraculum Omnipotentis vivificavit me.
JOB|33|5|Si potes, responde mihi,praepara te coram me et consiste.
JOB|33|6|Ecce ego sicut tu coram Deo sumet de eodem luto abscissus sum et ego.
JOB|33|7|Verumtamen terror meus non te terreat,et onus meum non sit tibi grave.
JOB|33|8|Dixisti ergo in auribus meis,et vocem verborum tuorum audivi:
JOB|33|9|"Mundus sum ego et absque delicto;immaculatus, et non est iniquitas in me.
JOB|33|10|Quia querelas in me repperit,ideo arbitratus est me inimicum sibi;
JOB|33|11|posuit in nervo pedes meos,custodivit omnes semitas meas".
JOB|33|12|Hoc est ergo, in quo non es iustificatus, respondebo tibi,quia maior est Deus homine.
JOB|33|13|Quare adversus eum contendis,quod non ad omnia verba responderit tibi?
JOB|33|14|Semel loquitur Deus,et secundo idipsum non repetit.
JOB|33|15|Per somnium in visione nocturna,quando irruit sopor super homines,et dormiunt in lectulo,
JOB|33|16|tunc aperit aures virorumet in visionibus terret eos,
JOB|33|17|ut avertat hominem ab his, quae facit,et liberet eum de superbia,
JOB|33|18|eruens animam eius a foveaet vitam illius, ut non transeat canalem mortis.
JOB|33|19|Increpat quoque per dolorem in lectulo,et tremitus ossium eius continuus.
JOB|33|20|Abominabilis ei fit in vita sua panis,et animae illius cibus ante desiderabilis.
JOB|33|21|Tabescet caro eius in conspectu,et ossa, quae non videbantur, nudabuntur.
JOB|33|22|Appropinquavit corruptioni foveae,et vita illius mortiferis sedibus.
JOB|33|23|Si fuerit apud eum angelus, unus de milibus interpres,ut annuntiet homini aequitatem,
JOB|33|24|miserebitur eius et dicet:Libera eum, ut non descendat in foveam;inveni, in quo ei propitier".
JOB|33|25|Revirescet caro eius plus quam in iuventute,revertetur ad dies adulescentiae suae.
JOB|33|26|Deprecabitur Deum, et placabilis ei erit;et videbit faciem eius in iubilo,et reddet homini iustitiam suam.
JOB|33|27|Canit ad homines et dicit: "Peccavi et iustitiam pervertiet non debui satisfacere.
JOB|33|28|Liberavit animam suam, ne pergeret in foveam,sed vivens lucem videret".
JOB|33|29|Ecce haec omnia operatur Deusduobus, tribus vicibus cum homine,
JOB|33|30|ut revocet animas eorum a foveaet illuminet luce viventium.
JOB|33|31|Attende, Iob, et audi meet tace, dum ego loquor.
JOB|33|32|Si autem habes quod loquaris, responde mihi; loquere, volo enim te apparere iustum.
JOB|33|33|Quod si non habes, audi me;tace, et docebo te sapientiam ".
JOB|34|1|Pronuntians itaque Eliu etiam haec locutus est:
JOB|34|2|" Audite, sapientes, verba mea;et eruditi, auscultate me.
JOB|34|3|Auris enim verba probat,et guttur escas gustu diiudicat.
JOB|34|4|Iudicium eligamus nobiset inter nos videamus quid sit melius.
JOB|34|5|Quia dixit Iob: "Iustus sum,et Deus avertit iudicium meum;
JOB|34|6|in iudicando enim me mendacium est,violenta sagitta mea absque ullo peccato".
JOB|34|7|Quis est vir, ut est Iob,qui bibit subsannationem quasi aquam,
JOB|34|8|qui graditur una cum operantibus iniquitatemet ambulat cum viris impiis?
JOB|34|9|Dixit enim: "Non prodest viro,etiamsi cum Deo familiariter agit".
JOB|34|10|Ideo, viri cordati, audite me:Absit a Deo impietas, et ab Omnipotente iniquitas.
JOB|34|11|Opus enim hominis reddet eiet iuxta vias singulorum restituet eis.
JOB|34|12|Vere enim Deus non operatur malum,nec Omnipotens subvertet iudicium.
JOB|34|13|Quis commisit ei terram suam,aut quis posuit totum orbem?
JOB|34|14|Si direxerit ad se cor suum,spiritum illius et halitum ad se trahat,
JOB|34|15|deficiet omnis caro simul,et homo in cinerem revertetur.
JOB|34|16|Si habes ergo intellectum, audi hocet ausculta vocem eloquii mei:
JOB|34|17|Numquid, qui non amat iudicium, reget imperio?Num iustum magnum condemnabis,
JOB|34|18|qui dicet regi: "Nequam!",qui vocabit duces: "Impios!",
JOB|34|19|qui non accipit personas principumnec cognovit opulentum,cum disceptaret contra pauperem?Opus enim manuum eius sunt universi.
JOB|34|20|Subito morientur; et in media nocteturbabuntur populi et pertransibunt,et auferent violentum absque conatu.
JOB|34|21|Oculi enim eius super vias hominum,et omnes gressus eorum considerat.
JOB|34|22|Non sunt tenebrae, et non est umbra mortis,ut abscondantur ibi, qui operantur iniquitatem.
JOB|34|23|Nec enim ultra homini ponit conveniendi locum,ut veniat ad Deum in iudicium.
JOB|34|24|Conteret potentes sine inquisitioneet stare faciet alios pro eis.
JOB|34|25|Novit enim opera eorumet idcirco inducet noctem, et conterentur.
JOB|34|26|Quasi impios percussit eosin loco videntium,
JOB|34|27|qui quasi de industria recesserunt ab eoet omnes vias eius intellegere noluerunt,
JOB|34|28|cum induceret ad se clamorem egeni et audiret vocem pauperum.
JOB|34|29|Ipse enim si quieverit, quis est qui condemnet?Et si absconderit vultum, quis est qui contempletur eum,super gentem et super homines simul?
JOB|34|30|Ne regnet homo impius,ne sint laquei populo.
JOB|34|31|Si enim dixit quispiam Deo:Ferre debui! Iam non perverse agam.
JOB|34|32|Dum videam, tu doce me;si iniquitatem operatus sum, ultra non addam".
JOB|34|33|Numquid pro te Deus satisfaciet,quia respuisti?Tu enim eliges, et non ego;et si quid nosti melius, loquere.
JOB|34|34|Viri intellegentes loquentur mihi,et vir sapiens, qui audiet me:
JOB|34|35|"Iob autem non in sapientia locutus est,et verba illius non sonant disciplinam".
JOB|34|36|Utique, probetur Iob usque ad finemde responsionibus hominum iniquitatis.
JOB|34|37|Quia addit super peccata sua delictum,inter nos plaudit manibuset multiplicat sermones suos contra Deum ".
JOB|35|1|Igitur Eliu haec rursum locutus est:
JOB|35|2|" Numquid aequa tibi videtur tua cogitatio,ut diceres: "Iustificatio mea coram Deo"?
JOB|35|3|Dixisti enim: "Quid ad te?Vel quid tibi proderit, si ego peccavero?".
JOB|35|4|Itaque ego respondebo sermonibus tuiset amicis tuis tecum.
JOB|35|5|Suspice caelum et intuereet contemplare nubes quod altiores te sint.
JOB|35|6|Si peccaveris, quid facies ei?Et si multiplicatae fuerint iniquitates tuae, quid facies contra eum?
JOB|35|7|Porro si iuste egeris, quid donabis ei?Aut quid de manu tua accipiet?
JOB|35|8|Homini, qui similis tui est, nocebit impietas tua,et filium hominis adiuvabit iustitia tua.
JOB|35|9|Propter multitudinem oppressorum clamabuntet eiulabunt propter vim brachii tyrannorum,
JOB|35|10|sed nemo dixit: "Ubi est Deus, qui fecit me,qui dedit carmina in nocte,
JOB|35|11|qui docet nos super iumenta terraeet super volucres caeli erudit nos?".
JOB|35|12|Ibi clamabunt, et non exaudiet,propter superbiam malorum.
JOB|35|13|Etiam, frustra: non audiet Deus,et Omnipotens non intuebitur.
JOB|35|14|Omnino cum dixeris: "Non considerat",iudicium est coram illo, et exspectas eum.
JOB|35|15|Et nunc cum dicis: "Ira eius poenas non infert,nec ulciscitur scelus valde",
JOB|35|16|Iob frustra aperit os suumet absque scientia verba multiplicat ".
JOB|36|1|Addens quoque Eliu haec locutus est:
JOB|36|2|" Sustine me paululum, et indicabo tibi:adhuc enim habeo quod pro Deo loquar.
JOB|36|3|Repetam scientiam meam a longeet Factori meo tribuam iustitiam.
JOB|36|4|Vere enim absque mendacio sermones mei,et perfectus scientia adest tecum.
JOB|36|5|Deus potens est; non abicit,potens virtute cordis.
JOB|36|6|Non vivere faciet impium,sed iudicium pauperibus tribuit.
JOB|36|7|Non auferet a iusto oculos suoset reges in solio collocat in perpetuum,et illi eriguntur.
JOB|36|8|Et si fuerint vincti compedibuset vinciantur funibus paupertatis,
JOB|36|9|indicabit eis opera eorumet scelera eorum, quia violenti fuerunt.
JOB|36|10|Revelabit quoque aurem eorum, ut corripiat,et loquetur, ut revertantur ab iniquitate.
JOB|36|11|Si audierint et observaverint,complebunt dies suos in bonoet annos suos in deliciis.
JOB|36|12|Si autem non audierint, transibunt per canalem mortiset consumentur in stultitia.
JOB|36|13|Impii corde sibi reponent iram Deineque clamabunt, cum vincti fuerint.
JOB|36|14|Morietur in iuventute anima eorum,et vita eorum in adulescentia.
JOB|36|15|Eripiet de angustia sua pauperemet revelabit in tribulatione aurem eius.
JOB|36|16|Igitur salvabit te de ore angusto,amplitudo et non angustiae erunt sub te;requies autem mensae tuae erit plena pinguedine.
JOB|36|17|Causa tua quasi impii iudicata est,causam iudiciumque tenebunt.
JOB|36|18|Cave, ne te seducat abundantia,nec multitudo donorum inclinet te.
JOB|36|19|Nonne proferetur clamor tuus nisi in angustia?Et omnes conatus roboris?
JOB|36|20|Ne inhies nocti,ut ascendat turba pro eis.
JOB|36|21|Cave, ne declines ad iniquitatem;propter hoc enim expertus es miseriam.
JOB|36|22|Ecce, Deus excelsus in fortitudine sua.Quis ei similis doctor?
JOB|36|23|Quis poterit scrutari vias eius,aut quis potest ei dicere: "Operatus es iniquitatem"?
JOB|36|24|Memento, ut magnifices opus eius,de quo cecinerunt viri.
JOB|36|25|Omnes homines vident eum,unusquisque intuetur procul.
JOB|36|26|Ecce, Deus magnus vincens scientiam nostram;numerus annorum eius inaestimabilis.
JOB|36|27|Qui aufert stillas pluviaeet effundit imbres ad instar fluminis,
JOB|36|28|quos nubes effundunt,stillantes super homines multos.
JOB|36|29|Profecto quis intellegit dilatationem nubium,strepitum tabernaculi eius?
JOB|36|30|Ecce extendit circum se lumen suumet fundamenta maris texit.
JOB|36|31|Per haec enim iudicat populoset dat escas copiose.
JOB|36|32|In manibus abscondit lucemet praecipit ei, ut percutiat.
JOB|36|33|Fragor eius de eo annuntiat,zelans ira contra iniquitatem.
JOB|37|1|Super hoc expavit cor meumet emotum est de loco suo.
JOB|37|2|Audite fremitum vocis eiuset murmur de ore illius procedens.
JOB|37|3|Subter omnes caelos ipsum revolvit,et lumen illius super terminos terrae.
JOB|37|4|Post eum rugiet sonitus,tonabit voce magnitudinis suae;et non retardabit, cum audita fuerit vox eius.
JOB|37|5|Tonabit Deus in voce sua mirabiliter,qui facit magna et inscrutabilia.
JOB|37|6|Qui praecipit nivi, ut descendat in terram,et hiemis pluviis et imbri, ut roborentur.
JOB|37|7|Qui in manu omnium hominum signat,ut noverint singuli opera sua.
JOB|37|8|Ingredietur bestia latibulumet in antro suo morabitur.
JOB|37|9|Ab interioribus egredietur tempestas,et ab Arcturo frigus.
JOB|37|10|Flante Deo, datur gelu,et expansio aquarum solidatur.
JOB|37|11|Fulgur proicitur a nube,et nubes spargunt lumen suum;
JOB|37|12|quae lustrant per circuitum,quocumque eas voluntas gubernantis duxerit,ad omne, quod praeceperit illis super faciem orbis terrarum,
JOB|37|13|sive in castigatione terrae suae,sive in misericordia eas iusserit inveniri.
JOB|37|14|Ausculta haec, Iob;sta et considera mirabilia Dei.
JOB|37|15|Numquid scis quando praeceperit Deus,ut ostenderent lucem nubes eius?
JOB|37|16|Numquid nosti semitas nubium magnaset mirabilia perfecti scientia?
JOB|37|17|Nonne vestimenta tua calida sunt,cum quieverit terra austro?
JOB|37|18|Tu forsitan cum eo expandisti caelos,qui solidissimi, quasi aere, fusi sunt?
JOB|37|19|Ostende nobis quid dicamus illi;nos disponere verba nescimus propter tenebras.
JOB|37|20|Quis narrabit ei, quae loquor?Et, si locutus fuerit, homo deglutietur.
JOB|37|21|At nunc non vident lucem:aer offuscatus est nubibus,sed ventus transiens fugabit eas.
JOB|37|22|Ab aquilone splendor auri venit;et circa Deum terribilis maiestas.
JOB|37|23|Omnipotentem attingere non possumus: magnus fortitudine;et iudicium et multam iustitiam deprimere non potest.
JOB|37|24|Ideo timebunt eum homines,non contemplabitur omnes, qui sibi videntur corde sapientes ".
JOB|38|1|Respondens autem Dominus Iob de turbine dixit:
JOB|38|2|" Quis est iste obscurans consiliumsermonibus imperitis?
JOB|38|3|Accinge sicut vir lumbos tuos;interrogabo te, et edoce me.
JOB|38|4|Ubi eras, quando ponebam fundamenta terrae?Indica mihi, si habes intellegentiam.
JOB|38|5|Quis posuit mensuras eius, si nosti?Vel quis tetendit super eam lineam?
JOB|38|6|Super quo bases illius solidatae sunt?Aut quis demisit lapidem angularem eius,
JOB|38|7|cum clamarent simul astra matutina,et iubilarent omnes filii Dei?
JOB|38|8|Quis conclusit ostiis mare,quando erumpebat quasi de visceribus procedens,
JOB|38|9|cum ponerem nubem vestimentum eiuset caligine illud quasi fascia obvolverem?
JOB|38|10|Definivi illud terminis meiset posui vectem et ostia
JOB|38|11|et dixi: Usque huc venies et non procedes ampliuset hic confringes tumentes fluctus tuos.
JOB|38|12|Numquid in diebus tuis praecepisti diluculoet assignasti aurorae locum suum,
JOB|38|13|et, cum extrema terrae teneres,excussi sunt impii ex ea?
JOB|38|14|Vertetur in lutum signatumet stabit sicut vestimentum.
JOB|38|15|Cohibetur ab impiis lux sua,et brachium excelsum confringetur.
JOB|38|16|Numquid ingressus es scaturigines mariset in novissimis abyssi deambulasti?
JOB|38|17|Numquid apertae sunt tibi portae mortis,et ostia tenebrosa vidisti?
JOB|38|18|Numquid considerasti latitudinem terrae?Indica mihi, si nosti omnia:
JOB|38|19|In qua via lux habitet,et tenebrarum quis locus sit;
JOB|38|20|ut ducas unumquodque ad terminos suoset intellegas semitas domus eius?
JOB|38|21|Novisti, nam tunc natus eras,et numerus dierum tuorum multus!
JOB|38|22|Numquid ingressus es thesauros nivisaut thesauros grandinis aspexisti,
JOB|38|23|quae praeparavi in tempus angustiae,in diem pugnae et belli?
JOB|38|24|Per quam viam spargitur lux,diffunditur ventus urens super terram?
JOB|38|25|Quis dedit vehementissimo imbri cursumet viam fulmini tonanti,
JOB|38|26|ut plueret super terram absque homine,in deserto, ubi nullus mortalium commoratur,
JOB|38|27|ut impleret inviam et desolatamet produceret herbas in terra arida?
JOB|38|28|Quis est pluviae pater,vel quis genuit stillas roris?
JOB|38|29|De cuius sinu egressa est glacies,et pruinam de caelo quis genuit?
JOB|38|30|In similitudinem lapidis aquae durantur,et superficies abyssi constringitur.
JOB|38|31|Numquid coniungere valebis nexus stellarum Pleiadumaut funiculum Arcturi poteris solvere?
JOB|38|32|Numquid produces Coronam in tempore suoet Ursam cum filiis ducis tu?
JOB|38|33|Numquid nosti leges caeliet pones scripturam eius in terra?
JOB|38|34|Numquid elevabis in nebula vocem tuam,et impetus aquarum operiet te?
JOB|38|35|Numquid mittes fulgura, et ibuntet dicent tibi: "Adsumus!"?
JOB|38|36|Quis posuit in visceribus ibis sapientiam,vel quis dedit gallo intellegentiam?
JOB|38|37|Quis recensebit nubes in sapientia,et utres caeli quis declinabit,
JOB|38|38|quando funditur pulvis in solidum,et glebae compinguntur?
JOB|38|39|Numquid capies leaenae praedamet animam catulorum eius implebis,
JOB|38|40|quando cubant in antriset in specubus insidiantur?
JOB|38|41|Quis praeparat corvo escam suam,quando pulli eius clamant ad Deum vagantes,eo quod non habeant cibos?
JOB|39|1|Numquid nosti tempus partus ibicum in petrisvel parturientes cervas observasti?
JOB|39|2|Dinumerasti menses conceptus earumet scisti tempus partus earum?
JOB|39|3|Incurvantur ad fetum et pariuntet fetus suos emittunt.
JOB|39|4|Impinguantur filii earum et adolescunt in campo,egrediuntur et non revertuntur ad eas.
JOB|39|5|Quis dimisit onagrum liberum,et vincula ipsius quis solvit?
JOB|39|6|Cui dedi in solitudine domumet tabernacula eius in terra salsuginis.
JOB|39|7|Contemnit multitudinem civitatis,clamorem exactoris non audit.
JOB|39|8|Explorat montes pascuae suaeet virentia quaeque perquirit.
JOB|39|9|Numquid volet taurus ferus servire tibiaut morabitur ad praesepe tuum?
JOB|39|10|Numquid alligabis taurum ferum ad arandum loro tuo,aut confringet glebas vallium post te?
JOB|39|11|Numquid fiduciam habebis in magna fortitudine eiuset derelinques ei labores tuos?
JOB|39|12|Numquid credes illi quod revertaturet sementem in aream tuam congreget?
JOB|39|13|Ala struthionis laeta est,penna vero ciconiae et avolat.
JOB|39|14|Quando derelinquit ova sua in terra,in pulvere calefiunt.
JOB|39|15|Obliviscitur quod pes conculcet ea,aut bestia agri conterat.
JOB|39|16|Duratur ad filios suos quasi non sint sui;frustra laborans nullo timore anxiatur.
JOB|39|17|Privavit enim eam Deus sapientianec dedit illi intellegentiam.
JOB|39|18|Cum tempus fuerit, in altum alas erigit,deridet equum et ascensorem eius.
JOB|39|19|Numquid praebebis equo fortitudinemaut circumdabis collo eius iubam?
JOB|39|20|Numquid suscitabis eum quasi locustas?Gloria hinnitus eius terror;
JOB|39|21|vallem ungula fodit, exsultat audacter,in occursum pergit armatis.
JOB|39|22|Contemnit pavorem nec territurneque cedit gladio.
JOB|39|23|Super ipsum sonabit pharetra,micat hasta et acinaces.
JOB|39|24|Fervens et fremens sorbet terramnec consistet, cum tubae sonaverit clangor.
JOB|39|25|Ubi audierit bucinam, dicit: "Uah!".Procul odoratur bellum,exhortationem ducum et ululatum exercitus.
JOB|39|26|Numquid per sapientiam tuam plumescit accipiter,expandens alas suas ad austrum?
JOB|39|27|Numquid ad praeceptum tuum elevabitur aquilaet in arduis ponet nidum suum?
JOB|39|28|In petris manetet in praeruptis silicibus commoraturatque in culmine et arce.
JOB|39|29|Inde contemplatur escam,et de longe oculi eius prospiciunt.
JOB|39|30|Pulli eius lambent sanguinem;et, ubicumque cadaver fuerit, statim adest ".
JOB|40|1|Et respondens Dominus locutus est ad Iob:
JOB|40|2|" Numquid contendit cum Omnipotente reprehensor?Qui arguit Deum, debet respondere ad ea ".
JOB|40|3|Respondens autem Iob Domino dixit:
JOB|40|4|" Ecce leviter locutus sum, quid respondebo tibi?Manum meam ponam super os meum.
JOB|40|5|Unum locutus sum, quod non repetam,et alterum, quibus ultra non addam ".
JOB|40|6|Respondens autem Dominus Iob de turbine dixit:
JOB|40|7|" Accinge sicut vir lumbos tuos;interrogabo te, et edoce me.
JOB|40|8|Numquid irritum facies iudicium meumet condemnabis me, ut tu iustificeris?
JOB|40|9|Et si habes brachium sicut Deuset si voce simili tonas?
JOB|40|10|Circumda tibi decorem et sublimitatem;gloria et decore induere.
JOB|40|11|Effunde vehementiam furoris tuiet respiciens omnem arrogantem humilia.
JOB|40|12|Respice cunctos superbos et confunde eoset contere impios in loco suo.
JOB|40|13|Absconde eos in pulvere simulet facies eorum claude in fovea;
JOB|40|14|et ego confiteborquod salvare te possit dextera tua.
JOB|40|15|Ecce Behemoth, quem feci tecum;fenum quasi bos comedit.
JOB|40|16|Fortitudo eius in lumbis eius,et virtus illius in umbilico ventris eius.
JOB|40|17|Stringit caudam suam quasi cedrum,nervi femorum eius perplexi sunt.
JOB|40|18|Ossa eius velut fistulae aeris,cartilago illius quasi laminae ferreae.
JOB|40|19|Ipse est principium viarum Dei;qui fecit eum, applicabit gladium eius.
JOB|40|20|Huic montes tributum ferunt,omnes bestiae agri ludunt ibi.
JOB|40|21|Sub lotis silvestribus dormit,in secreto calami et in locis umentibus;
JOB|40|22|loti silvestres umbra eum protegunt,circumdant eum salices torrentis.
JOB|40|23|Si fluvius intumescat, non tremit;securus est, si prorumpat fluctus ad os eius.
JOB|40|24|In oculis eius quis capiet eumet in sudibus perforabit nares eius?
JOB|40|25|An extrahere poteris Leviathan hamoet fune ligabis linguam eius?
JOB|40|26|Numquid pones iuncum in naribus eiusaut spina perforabis maxillam eius?
JOB|40|27|Numquid multiplicabit ad te precesaut loquetur tibi mollia?
JOB|40|28|Numquid feriet tecum pactum,et accipies eum servum sempiternum?
JOB|40|29|Numquid illudes ei quasi aviaut ligabis eum pro puellis tuis?
JOB|40|30|Speculabuntur super eum socii,divident illum negotiatores?
JOB|40|31|Numquid implebis telis pellem eiuset iaculo hamato piscium caput illius?
JOB|40|32|Pone super eum manum tuam;memento belli nec ultra addas.
JOB|41|1|Ecce spes eius frustrabitur eum,et aspectu eius praecipitabitur.
JOB|41|2|Nemo tam audax, ut suscitet eum.Quis enim resistere potest vultui eius?
JOB|41|3|Quis eum aggressus est et salvus fuit?Sub omni caelo quisnam?
JOB|41|4|Non tacebo super membra eiuset eloquar robur et gratiam struis.
JOB|41|5|Quis revelabit faciem indumenti eius,et duplicia mandibulae eius quis intrabit?
JOB|41|6|Portas vultus eius quis aperiet?Per gyrum dentium eius formido.
JOB|41|7|Corpus illius quasi scuta fusilia,compactum sigillo siliceo:
JOB|41|8|unum uni coniungitur,et ne spiraculum quidem incedit per ea;
JOB|41|9|unum alteri adhaeret,et tenentes se nequaquam separantur.
JOB|41|10|Sternutatio eius favillae ignis,et oculi eius ut palpebrae diluculi.
JOB|41|11|De ore eius lampades procedunt,sicut scintillae ignis emittuntur.
JOB|41|12|De naribus eius procedit fumus,sicut ollae succensae atque ferventis.
JOB|41|13|Halitus eius prunas ardere facit,et flamma de ore eius egreditur.
JOB|41|14|In collo eius morabitur fortitudo,et faciem eius praecedit angor.
JOB|41|15|Palearia eius cohaerentia sibicompressa non moventur.
JOB|41|16|Cor eius induratur tamquam lapiset duratur quasi mola inferior.
JOB|41|17|Cum surrexerit, tremunt forteset ab undis retrorsum convertuntur.
JOB|41|18|Qui impegerit in eum, gladius eius non stabitnec hasta neque pilum neque thorax;
JOB|41|19|reputat enim quasi paleas ferrumet quasi lignum putridum aes.
JOB|41|20|Non fugat eum vir sagittarius,in stipulam versi sunt ei lapides fundae.
JOB|41|21|Quasi stipulam aestimat fustemet deridet vibrantem acinacem.
JOB|41|22|Sub ipso acumina testae,et sternit tribula super lutum.
JOB|41|23|Fervescere facit quasi ollam profundumet mare ponit quasi vas unguentarium.
JOB|41|24|Post se illuminat semitam,aestimatur abyssus quasi canescens.
JOB|41|25|Non est super terram potestas, quae comparetur ei,qui factus est, ut nullum timeret.
JOB|41|26|Omne sublime videt:ipse est rex super universos filios superbiae ".
JOB|42|1|Respondens autem Iob Domino dixit:
JOB|42|2|" Scio quia omnia potes,et nulla te latet cogitatio.
JOB|42|3|Quis est iste, qui celat consiliumabsque scientia?Ideo insipienter locutus sumet mirabilia, quae excederent scientiam meam.
JOB|42|4|Audi, et ego loquar;interrogabo te, et responde mihi.
JOB|42|5|Auditu auris audivi te;nunc autem oculus meus videt te.
JOB|42|6|Idcirco ipse me reprehendoet ago paenitentiam in favilla et cinere ".
JOB|42|7|Postquam autem locutus est Dominus verba haec ad Iob, dixit ad Eliphaz Themanitem: " Iratus est furor meus in te et in duos amicos tuos, quoniam non estis locuti coram me rectum sicut servus meus Iob.
JOB|42|8|Sumite ergo vobis septem tauros et septem arietes et ite ad servum meum Iob et offerte holocaustum pro vobis; Iob autem servus meus orabit pro vobis. Faciem eius suscipiam, ut non vobis imputetur stultitia; neque enim locuti estis ad me recta sicut servus meus Iob ".
JOB|42|9|Abierunt ergo Eliphaz Themanites et Baldad Suhites et Sophar Naamathites et fecerunt, sicut locutus fuerat Dominus ad eos, et suscepit Dominus faciem Iob.
JOB|42|10|Dominus vertit sortem Iob, cum oraret ille pro amicis suis; et addidit Dominus omnia, quaecumque fuerant Iob, duplicia.
JOB|42|11|Venerunt autem ad eum omnes fratres sui et universae sorores suae et cuncti, qui noverant eum prius; et comederunt cum eo panem in domo eius et moverunt super eum caput et consolati sunt eum super omni malo, quod intulerat Dominus super eum; et dederunt ei unusquisque argenteum unum et inaurem auream unam.
JOB|42|12|Dominus autem benedixit novissimis Iob magis quam principio eius; et facta sunt ei quattuordecim milia ovium et sex milia camelorum et mille iuga boum et mille asinae.
JOB|42|13|Et fuerunt ei septem filii et tres filiae;
JOB|42|14|et vocavit nomen unius Columbam et nomen secundae Cassiam et nomen tertiae Cornustibii.
JOB|42|15|Non sunt autem inventae mulieres speciosae sicut filiae Iob in universa terra; deditque eis pater suus hereditatem inter fratres earum.
JOB|42|16|Vixit autem Iob post haec centum quadraginta annis et vidit filios suos et filios filiorum suorum usque ad quartam generationem; et mortuus est senex et plenus dierum.
PS|1|1|Beatus vir, qui non abiit in consilio impiorumet in via peccatorum non stetitet in conventu derisorum non sedit,
PS|1|2|sed in lege Domini voluntas eius,et in lege eius meditatur die ac nocte.
PS|1|3|Et erit tamquam lignum plantatum secus decursus aquarum,quod fructum suum dabit in tempore suo;et folium eius non defluet,et omnia, quaecumque faciet, prosperabuntur.
PS|1|4|Non sic impii, non sic,sed tamquam pulvis, quem proicit ventus.
PS|1|5|Ideo non consurgent impii in iudicio,neque peccatores in concilio iustorum.
PS|1|6|Quoniam novit Dominus viam iustorum,et iter impiorum peribit.
PS|2|1|Quare fremuerunt gentes,et populi meditati sunt inania?
PS|2|2|Astiterunt reges terrae,et principes convenerunt in unumadversus Dominum et adversus christum eius:
PS|2|3|" Dirumpamus vincula eorumet proiciamus a nobis iugum ipsorum! ".
PS|2|4|Qui habitat in caelis, irridebit eos,Dominus subsannabit eos.
PS|2|5|Tunc loquetur ad eos in ira suaet in furore suo conturbabit eos:
PS|2|6|" Ego autem constitui regem meum super Sion, montem sanctum meum! ".
PS|2|7|Praedicabo decretum eius.Dominus dixit ad me: " Filius meus es tu;ego hodie genui te.
PS|2|8|Postula a me, et dabo tibi gentes hereditatem tuamet possessionem tuam terminos terrae.
PS|2|9|Reges eos in virga ferreaet tamquam vas figuli confringes eos ".
PS|2|10|Et nunc, reges, intellegite;erudimini, qui iudicatis terram.
PS|2|11|Servite Domino in timoreet exsultate ei cum tremore.
PS|2|12|Apprehendite disciplinam, ne quando irascatur,et pereatis de via,cum exarserit in brevi ira eius.Beati omnes, qui confidunt in eo.
PS|3|1|PSALMUS. David, cum fugit a filio suo Absalom.
PS|3|2|Domine, quid multiplicati sunt, qui tribulant me?Multi insurgunt adversum me,
PS|3|3|multi dicunt animae meae: Non est salus ipsi in Deo ".
PS|3|4|Tu autem, Domine, protector meus es,gloria mea et exaltans caput meum.
PS|3|5|Voce mea ad Dominum clamavi,et exaudivit me de monte sancto suo.
PS|3|6|Ego obdormivi et soporatus sum,exsurrexi, quia Dominus suscepit me.
PS|3|7|Non timebo milia populi circumdantis me.Exsurge, Domine salvum me fac, Deus meus;
PS|3|8|quoniam tu percussisti in maxillam omnes adversantes mihi,dentes peccatorum contrivisti.
PS|3|9|Domini est salus,et super populum tuum benedictio tua.
PS|4|1|Magistro chori. Fidibus. PSALMUS. David.
PS|4|2|Cum invocarem, exaudivit me Deus iustitiae meae.In tribulatione dilatasti mihi;miserere mei et exaudi orationem meam.
PS|4|3|Filii hominum, usquequo gravi corde?Ut quid diligitis vanitatem et quaeritis mendacium?
PS|4|4|Et scitote quoniam mirificavit Dominus sanctum suum;Dominus exaudiet, cum clamavero ad eum.
PS|4|5|Irascimini et nolite peccare;loquimini in cordibus vestris,in cubilibus vestris et conquiescite.
PS|4|6|Sacrificate sacrificium iustitiaeet sperate in Domino.
PS|4|7|Multi dicunt: " Quis ostendit nobis bona? ".Leva in signum super nos lumen vultus tui, Domine!
PS|4|8|Maiorem dedisti laetitiam in corde meo,quam cum multiplicantur frumentum et vinum eorum.
PS|4|9|In pace in idipsum dormiam et requiescam,quoniam tu, Domine, singulariter in spe constituisti me.
PS|5|1|Magistro chori. Ad tibias. PSALMUS. David.
PS|5|2|Verba mea auribus percipe, Domine;intellege gemitum meum.
PS|5|3|Intende voci clamoris mei,rex meus et Deus meus.
PS|5|4|Quoniam ad te orabo, Domine,mane exaudies vocem meam;mane astabo tibi et exspectabo.
PS|5|5|Quoniam non Deus volens iniquitatem tu es;neque habitabit iuxta te malignus,
PS|5|6|neque permanebunt iniusti ante oculos tuos.
PS|5|7|Odisti omnes, qui operantur iniquitatem,perdes omnes, qui loquuntur mendacium;virum sanguinum et dolosum abominabitur Dominus.
PS|5|8|Ego autem in multitudine misericordiae tuaeintroibo in domum tuam;adorabo ad templum sanctum tuum in timore tuo.
PS|5|9|Domine, deduc me in iustitia tua propter inimicos meos,dirige in conspectu meo viam tuam.
PS|5|10|Quoniam non est in ore eorum veritas,cor eorum fovea;sepulcrum patens est guttur eorum,molliunt linguas suas.
PS|5|11|Iudica illos, Deus; decidant a cogitationibus suis;secundum multitudinem impietatum eorum expelle eos,quoniam irritaverunt te, Domine.
PS|5|12|Et omnes, qui sperant in te,laetentur, in aeternum exsultent.Obumbrabis eis, et gloriabuntur in te,qui diligunt nomen tuum;
PS|5|13|quoniam tu benedices iusto, Domine,quasi scuto, bona voluntate coronabis eum.
PS|6|1|Magistro chori. Fidibus. Super octavam. PSALMUS. David.
PS|6|2|Domine, ne in furore tuo arguas meneque in ira tua corripias me.
PS|6|3|Miserere mei, Domine, quoniam infirmus sum;sana me, Domine, quoniam conturbata sunt ossa mea.
PS|6|4|Et anima mea turbata est valde,sed tu, Domine, usquequo?
PS|6|5|Convertere, Domine, eripe animam meam;salvum me fac propter misericordiam tuam.
PS|6|6|Quoniam non est in morte, qui memor sit tui;in inferno autem quis confitebitur tibi?
PS|6|7|Laboravi in gemitu meo,lavabam per singulas noctes lectum meum;lacrimis meis stratum meum rigabam.
PS|6|8|Turbatus est a maerore oculus meus,inveteravi inter omnes inimicos meos.
PS|6|9|Discedite a me, omnes, qui operamini iniquitatem,quoniam exaudivit Dominus vocem fletus mei.
PS|6|10|Exaudivit Dominus deprecationem meam,Dominus orationem meam suscepit.
PS|6|11|Erubescant et conturbentur vehementer omnes inimici mei;convertantur et erubescant valde velociter.
PS|7|1|Lamentatio David, quam cantavit Domino propter Chus Beniaminitam.
PS|7|2|Domine Deus meus, in te speravi;salvum me fac ex omnibus persequentibus me et libera me,
PS|7|3|ne quando rapiat ut leo animam meamdiscerpens, dum non est qui salvum faciat.
PS|7|4|Domine Deus meus, si feci istud,si est iniquitas in manibus meis,
PS|7|5|si reddidi retribuenti mihi malaet exspoliavi inimicum meum dimittens inanem,
PS|7|6|persequatur inimicus animam meam et comprehendatet conculcet in terra vitam meamet gloriam meam in pulverem deducat.
PS|7|7|Exsurge, Domine, in ira tuaet exaltare contra indignationem inimicorum meorumet exsurge, Deus meus, in iudicio, quod mandasti.
PS|7|8|Et synagoga populorum circumdabit te,et super hanc in altum regredere:
PS|7|9|Dominus iudicat populos.Iudica me, Domine, secundum iustitiam meamet secundum innocentiam meam, quae est in me.
PS|7|10|Consumatur nequitia peccatorum;et iustum confirma:scrutans corda et renes Deus iustus.
PS|7|11|Adiutorium meum apud Deum,qui salvos facit rectos corde.
PS|7|12|Deus iudex iustus,fortis, irascens per singulos dies.
PS|7|13|Nonne iterum gladium suum exacuit,arcum suum tetendit et paravit illum?
PS|7|14|Et paravit sibi vasa mortis,sagittas suas ardentes effecit.
PS|7|15|Ecce parturiit iniustitiam,concepit dolorem et peperit iniquitatem;
PS|7|16|lacum aperuit et effodit eumet incidit in foveam, quam fecit.
PS|7|17|Convertetur dolor eius in caput eius,et in verticem ipsius iniquitas eius descendet.
PS|7|18|Confitebor Domino secundum iustitiam eiuset psallam nomini Domini Altissimi.
PS|8|1|Magistro chori. Ad modum cantici " Torcularia... ". PSALMUS. David.
PS|8|2|Domine, Dominus noster,quam admirabile est nomen tuum in universa terra,quoniam elevata est magnificentia tua super caelos.
PS|8|3|Ex ore infantium et lactantium perfecisti laudempropter inimicos tuos,ut destruas inimicum et ultorem.
PS|8|4|Quando video caelos tuos, opera digitorum tuorum,lunam et stellas, quae tu fundasti,
PS|8|5|quid est homo, quod memor es eius,aut filius hominis, quoniam visitas eum?
PS|8|6|Minuisti eum paulo minus ab angelis,gloria et honore coronasti eum
PS|8|7|et constituisti eum super opera manuum tuarum.Omnia subiecisti sub pedibus eius:
PS|8|8|oves et boves universas,insuper et pecora campi,
PS|8|9|volucres caeli et pisces maris,quaecumque perambulant semitas maris.
PS|8|10|Domine, Dominus noster,quam admirabile est nomen tuum in universa terra!
PS|9|1|Magistro chori. Ad modum cantici " Mut labben ". PSALMUS. David.
PS|9|2|ALEPH. Confitebor tibi, Domine, in toto corde meo,narrabo omnia mirabilia tua.
PS|9|3|Laetabor et exsultabo in te,psallam nomini tuo, Altissime.
PS|9|4|BETH. Cum convertuntur inimici mei retrorsum,infirmantur et pereunt a facie tua.
PS|9|5|Quoniam fecisti iudicium meum et causam meam,sedisti super thronum, qui iudicas iustitiam.
PS|9|6|GHIMEL. Increpasti gentes, perdidisti impium;nomen eorum delesti in aeternum et in saeculum saeculi.
PS|9|7|Inimici defecerunt, solitudines sempiternae factae sunt;et civitates destruxisti: periit memoria eorum cum ipsis.
PS|9|8|HE. Dominus autem in aeternum sedebit,paravit in iudicium thronum suum;
PS|9|9|et ipse iudicabit orbem terrae in iustitia,iudicabit populos in aequitate.
PS|9|10|VAU. Et erit Dominus refugium oppresso,refugium in opportunitatibus, in tribulatione.
PS|9|11|Et sperent in te, qui noverunt nomen tuum,quoniam non dereliquisti quaerentes te, Domine.
PS|9|12|ZAIN. Psallite Domino, qui habitat in Sion;annuntiate inter gentes studia eius.
PS|9|13|Quoniam requirens sanguinem recordatus est eorum,non est oblitus clamorem pauperum.
PS|9|14|HETH. Miserere mei, Domine;vide afflictionem meam de inimicis meis,qui exaltas me de portis mortis,
PS|9|15|ut annuntiem omnes laudationes tuas in portis filiae Sion,exsultem in salutari tuo.
PS|9|16|TETH. Infixae sunt gentes in fovea, quam fecerunt;in laqueo isto, quem absconderunt,comprehensus est pes eorum.
PS|9|17|Manifestavit se Dominus iudicium faciens;in operibus manuum suarum comprehensus est peccator.
PS|9|18|IOD. Convertentur peccatores in infernum,omnes gentes, quae obliviscuntur Deum.
PS|9|19|CAPH. Quoniam non in finem oblivio erit pauperis;exspectatio pauperum non peribit in aeternum.
PS|9|20|Exsurge, Domine, non confortetur homo;iudicentur gentes in conspectu tuo.
PS|9|21|Constitue, Domine, terrorem super eos;sciant gentes quoniam homines sunt.
PS|10|1|LAMED. Ut quid, Domine, stas a longe,abscondis te in opportunitatibus, in tribulatione?
PS|10|2|Dum superbit, impius insequitur pauperem;comprehendantur in consiliis, quae cogitant.
PS|10|3|Quoniam gloriatur peccator in desideriis animae suae,et avarus sibi benedicit.
PS|10|4|NUN. Spernit Dominum peccator in arrogantia sua: Non requiret; non est Deus ".
PS|10|5|Hae sunt omnes cogitationes eius;prosperantur viae illius in omni tempore.Excelsa nimis iudicia tua a facie eius;omnes inimicos suos aspernatur.
PS|10|6|Dixit enim in corde suo: " Non movebor;in generationem et generationem ero sine malo ".
PS|10|7|PHE. Cuius maledictione os plenum est et fraudulentia et dolo,sub lingua eius labor et nequitia.
PS|10|8|Sedet in insidiis ad vicos,in occultis interficit innocentem.
PS|10|9|SADE. Oculi eius in pauperem respiciunt;insidiatur in abscondito quasi leo in spelunca sua.Insidiatur, ut rapiat pauperem;rapit pauperem, dum attrahit in laqueum suum.
PS|10|10|Irruit et inclinat se, et miseri caduntin fortitudine brachiorum eius.
PS|10|11|Dixit enim in corde suo: " Oblitus est Deus;avertit faciem suam, non videbit in finem ". -
PS|10|12|COPH. Exsurge, Domine Deus, exalta manum tuam,ne obliviscaris pauperum.
PS|10|13|Propter quid spernit impius Deum?Dixit enim in corde suo: " Non requires ".
PS|10|14|RES. Vidisti: tu laborem et dolorem consideras,ut tradas eos in manus tuas.Tibi derelictus est pauper,orphano tu factus es adiutor.
PS|10|15|SIN. Contere brachium peccatoris et maligni;quaeres peccatum illius et non invenies.
PS|10|16|Dominus rex in aeternum et in saeculum saeculi:perierunt gentes de terra illius.
PS|10|17|TAU. Desiderium pauperum exaudisti, Domine;confirmabis cor eorum, intendes aurem tuam
PS|10|18|iudicare pupillo et humili,ut non apponat ultra inducere timorem homo de terra.
PS|11|1|Magistro chori. David.In Domino confido, quomodo dicitis animae meae: Transmigra in montem sicut passer!
PS|11|2|Quoniam ecce peccatores intenderunt arcum,paraverunt sagittas suas super nervum,ut sagittent in obscuro rectos corde.
PS|11|3|Quando fundamenta evertuntur,iustus quid faciat? ".
PS|11|4|Dominus in templo sancto suo,Dominus, in caelo sedes eius.Oculi eius in pauperem respiciunt,palpebrae eius interrogant filios hominum.
PS|11|5|Dominus interrogat iustum et impium;qui autem diligit iniquitatem, odit anima eius.
PS|11|6|Pluet super peccatores carbones ignis et sulphur;et spiritus procellarum pars calicis eorum.
PS|11|7|Quoniam iustus Dominus et iustitias dilexit,recti videbunt vultum eius.
PS|12|1|Magistro chori. Super octavam. PSALMUS. David.
PS|12|2|Salvum me fac, Domine, quoniam defecit sanctus,quoniam deminuti sunt fideles a filiis hominum.
PS|12|3|Vana locuti sunt unusquisque ad proximum suum;in labiis dolosis, in duplici corde locuti sunt.
PS|12|4|Disperdat Dominus universa labia dolosaet linguam magniloquam.
PS|12|5|Qui dixerunt: " Lingua nostra magnificabimur,labia nostra a nobis sunt;quis noster dominus est? ".
PS|12|6|" Propter miseriam inopum et gemitum pauperum,nunc exsurgam, dicit Dominus;ponam in salutari illum, quem despiciunt ".
PS|12|7|Eloquia Domini eloquia casta,argentum igne examinatum, separatum a terra,purgatum septuplum.
PS|12|8|Tu, Domine, servabis nos et custodies nosa generatione hac in aeternum.In circuitu impii ambulant,cum exaltantur sordes inter filios hominum.
PS|13|1|Magistro chori. PSALMUS. David.
PS|13|2|Usquequo, Domine, oblivisceris me in finem?Usquequo avertes faciem tuam a me?
PS|13|3|Usquequo ponam consilia in anima mea,dolorem in corde meo per diem?Usquequo exaltabitur inimicus meus super me?
PS|13|4|Respice et exaudi me, Domine Deus meus.Illumina oculos meos, ne quando obdormiam in morte,
PS|13|5|ne quando dicat inimicus meus: " Praevalui adversus eum! ";neque exsultent, qui tribulant me, si motus fuero.
PS|13|6|Ego autem in misericordia tua speravi.Exsultabit cor meum in salutari tuo;cantabo Domino, qui bona tribuit mihi.
PS|14|1|Magistro chori. David.Dixit insipiens in corde suo: " Non est Deus ".Corrupti sunt et abominationes operati sunt;non est qui faciat bonum.
PS|14|2|Dominus de caelo prospexit super filios hominum,ut videret si est intellegens aut requirens Deum.
PS|14|3|Omnes declinaverunt, simul corrupti sunt;non est qui faciat bonum, non est usque ad unum.
PS|14|4|Nonne scient omnes, qui operantur iniquitatem,qui devorant plebem meam sicut escam panis?Dominum non invocaverunt;
PS|14|5|illic trepidaverunt timore,quoniam Deus cum generatione iusta est.
PS|14|6|Vos consilium inopis confundetis,Dominus autem spes eius est.
PS|14|7|Quis dabit ex Sion salutare Israel?Cum converterit Dominus captivitatem plebis suae,exsultabit Iacob, et laetabitur Israel.
PS|15|1|PSALMUS. David.Domine, quis habitabit in tabernaculo tuo?Quis requiescet in monte sancto tuo?
PS|15|2|Qui ingreditur sine macula et operatur iustitiam,qui loquitur veritatem in corde suo,
PS|15|3|qui non egit dolum in lingua suanec fecit proximo suo malumet opprobrium non intulit proximo suo.
PS|15|4|Ad nihilum reputatus est in conspectu eius malignus,timentes autem Dominum glorificat.Qui iuravit in detrimentum suum et non mutat,
PS|15|5|qui pecuniam suam non dedit ad usuramet munera super innocentem non accepit.Qui facit haec, non movebitur in aeternum.
PS|16|1|Miktam. David.Conserva me, Deus, quoniam speravi in te.
PS|16|2|Dixi Domino: " Dominus meus es tu, bonum mihi non est sine te ".
PS|16|3|In sanctos, qui sunt in terra, inclitos viros,omnis voluntas mea in eos.
PS|16|4|Multiplicantur dolores eorum, qui post deos alienos acceleraverunt.Non effundam libationes eorum de sanguinibusneque assumam nomina eorum in labiis meis.
PS|16|5|Dominus pars hereditatis meae et calicis mei:tu es qui detines sortem meam.
PS|16|6|Funes ceciderunt mihi in praeclaris;insuper et hereditas mea speciosa est mihi.
PS|16|7|Benedicam Dominum, qui tribuit mihi intellectum;insuper et in noctibus erudierunt me renes mei.
PS|16|8|Proponebam Dominum in conspectu meo semper;quoniam a dextris est mihi, non commovebor.
PS|16|9|Propter hoc laetatum est cor meum,et exsultaverunt praecordia mea;insuper et caro mea requiescet in spe.
PS|16|10|Quoniam non derelinques animam meam in infernonec dabis sanctum tuum videre corruptionem.
PS|16|11|Notas mihi facies vias vitae,plenitudinem laetitiae cum vultu tuo,delectationes in dextera tua usque in finem.
PS|17|1|Precatio. David.Exaudi, Domine, iustitiam meam,intende deprecationem meam.Auribus percipe orationem meam, non in labiis dolosis.
PS|17|2|De vultu tuo iudicium meum prodeat;oculi tui videant aequitates.
PS|17|3|Proba cor meum et visita nocte;igne me examina, et non invenies in me iniquitatem.
PS|17|4|Non transgreditur os meum ad opera hominum,propter verba labiorum tuorum custodivi me a viis violenti.
PS|17|5|Retine gressus meos in semitis tuis,ut non moveantur vestigia mea.
PS|17|6|Ego ad te clamavi, quoniam exaudis me, Deus;inclina aurem tuam mihi et exaudi verba mea.
PS|17|7|Mirifica misericordias tuas,qui salvos facis ab insurgentibussperantes in dextera tua.
PS|17|8|Custodi me ut pupillam oculi,sub umbra alarum tuarum protege me
PS|17|9|a facie impiorum, qui me afflixerunt.Inimici mei in furore circumdederunt me,
PS|17|10|adipem suum concluserunt;os eorum locutum est superbiam.
PS|17|11|Incedentes nunc circumdederunt me,oculos suos statuerunt prosternere in terram.
PS|17|12|Aspectus eorum quasi leonis parati ad praedamet sicut catuli leonis recubantis in abditis.
PS|17|13|Exsurge, Domine, praeveni eum, supplanta eum;eripe animam meam ab impio framea tua,
PS|17|14|a mortuis manu tua, Domine,a mortuis, quorum defecit portio vitae.De reconditis tuis adimpleas ventrem eorum,saturentur filii et dimittant reliquias parvulis suis.
PS|17|15|Ego autem in iustitia videbo faciem tuam;satiabor, cum evigilavero, conspectu tuo.
PS|18|1|Magistro chori. David, servi Domini,qui locutus est ad Dominum verba huius cantici,quando Dominus eum liberaverate potestate omnium inimicorum suorum
PS|18|2|et e manu Saul. Dixit igitur:Diligam te, Domine, fortitudo mea.
PS|18|3|Domine, firmamentum meum et refugium meum et liberator meus;Deus meus, adiutor meus, et sperabo in eum;protector meus et cornu salutis meae et susceptor meus.
PS|18|4|Laudabilem invocabo Dominum,et ab inimicis meis salvus ero.
PS|18|5|Circumdederunt me fluctus mortis,et torrentes Belial conturbaverunt me;
PS|18|6|funes inferni circumdederunt me,praeoccupaverunt me laquei mortis.
PS|18|7|In tribulatione mea invocavi Dominumet ad Deum meum clamavi;exaudivit de templo suo vocem meam,et clamor meus in conspectu eius introivit in aures eius.
PS|18|8|Commota est et contremuit terra;fundamenta montium concussa suntet commota sunt, quoniam iratus est.
PS|18|9|Ascendit fumus de naribus eius,et ignis de ore eius devorans;carbones succensi processerunt ab eo.
PS|18|10|Inclinavit caelos et descendit,et caligo sub pedibus eius.
PS|18|11|Et ascendit super cherub et volavit,ferebatur super pennas ventorum.
PS|18|12|Et posuit tenebras latibulum suum,in circuitu eius tabernaculum eius,tenebrosa aqua, nubes aeris.
PS|18|13|Prae fulgore in conspectu eius nubes transierunt,grando et carbones ignis.
PS|18|14|Et intonuit de caelo Dominus,et Altissimus dedit vocem suam:grando et carbones ignis.
PS|18|15|Et misit sagittas suas et dissipavit eos,fulgura iecit et conturbavit eos.
PS|18|16|Et apparuerunt fontes aquarum,et revelata sunt fundamenta orbis terrarumab increpatione tua, Domine,ab inspiratione spiritus irae tuae.
PS|18|17|Misit de summo et accepit meet assumpsit me de aquis multis;
PS|18|18|eripuit me de inimicis meis fortissimiset ab his, qui oderunt me,quoniam confortati sunt super me.
PS|18|19|Oppugnaverunt me in die afflictionis meae,et factus est Dominus fulcimentum meum;
PS|18|20|et eduxit me in latitudinem,salvum me fecit, quoniam voluit me.
PS|18|21|Et retribuet mihi Dominus secundum iustitiam meamet secundum puritatem manuum mearum reddet mihi,
PS|18|22|quia custodivi vias Domininec impie recessi a Deo meo.
PS|18|23|Quoniam omnia iudicia eius in conspectu meo,et iustitias eius non reppuli a me;
PS|18|24|et fui immaculatus cum eoet observavi me ab iniquitate.
PS|18|25|Et retribuit mihi Dominus secundum iustitiam meamet secundum puritatem manuum mearumin conspectu oculorum eius.
PS|18|26|Cum sancto sanctus eriset cum viro innocente innocens eris
PS|18|27|et cum electo electus eriset cum perverso callidus eris.
PS|18|28|Quoniam tu populum humilem salvum facieset oculos superborum humiliabis.
PS|18|29|Quoniam tu accendis lucernam meam, Domine;Deus meus illuminat tenebras meas.
PS|18|30|Quoniam in te aggrediar hostium turmaset in Deo meo transiliam murum.
PS|18|31|Deus, impolluta via eius,eloquia Domini igne examinata;protector est omnium sperantium in se.
PS|18|32|Quoniam quis Deus praeter Dominum?Aut quae munitio praeter Deum nostrum?
PS|18|33|Deus, qui praecinxit me virtuteet posuit immaculatam viam meam;
PS|18|34|qui perfecit pedes meos tamquam cervorumet super excelsa statuit me;
PS|18|35|qui docet manus meas ad proelium,et tendunt arcum aereum brachia mea.
PS|18|36|Et dedisti mihi scutum salutis tuae,et dextera tua suscepit me,et exauditio tua magnificavit me.
PS|18|37|Dilatasti gressus meos subtus me,et non sunt infirmata vestigia mea.
PS|18|38|Persequebar inimicos meos et comprehendebam illoset non convertebar, donec deficerent.
PS|18|39|Confringebam illos, nec poterant stare,cadebant subtus pedes meos.
PS|18|40|Et praecinxisti me virtute ad bellumet supplantasti insurgentes in me subtus me.
PS|18|41|Et inimicos meos dedisti mihi dorsumet odientes me disperdidisti.
PS|18|42|Clamaverunt, nec erat qui salvos faceret,ad Dominum, nec exaudivit eos.
PS|18|43|Et comminui eos ut pulverem ante faciem venti,ut lutum platearum contrivi eos.
PS|18|44|Eripuisti me de contradictionibus populi,constituisti me in caput gentium.Populus, quem non cognovi, servivit mihi,
PS|18|45|in auditu auris oboedivit mihi.Filii alieni blanditi sunt mihi,
PS|18|46|filii alieni inveterati sunt,contremuerunt in abditis suis.
PS|18|47|Vivit Dominus, et benedictus Adiutor meus,et exaltetur Deus salutis meae.
PS|18|48|Deus, qui das vindictas mihiet subdis populos sub me,liberator meus de inimicis meis iracundis;
PS|18|49|et ab insurgentibus in me exaltas me,a viro iniquo eripis me.
PS|18|50|Propterea confitebor tibi in nationibus, Domine,et nomini tuo psalmum dicam,
PS|18|51|magnificans salutes regis suiet faciens misericordiam christo suoDavid et semini eius usque in saeculum.
PS|19|1|Magistro chori. PSALMUS. David.
PS|19|2|Caeli enarrant gloriam Dei,et opera manuum eius annuntiat firmamentum.
PS|19|3|Dies diei eructat verbum,et nox nocti indicat scientiam.
PS|19|4|Non sunt loquelae neque sermones,quorum non intellegantur voces:
PS|19|5|in omnem terram exivit sonus eorum,et in fines orbis terrae verba eorum.
PS|19|6|Soli posuit tabernaculum in eis,et ipse, tamquam sponsus procedens de thalamo suo,exsultavit ut gigas ad currendam viam.
PS|19|7|A finibus caelorum egressio eius,et occursus eius usque ad fines eorum,nec est quod se abscondat a calore eius.
PS|19|8|Lex Domini immaculata, reficiens animam,testimonium Domini fidele, sapientiam praestans parvulis.
PS|19|9|Iustitiae Domini rectae, laetificantes corda,praeceptum Domini lucidum, illuminans oculos.
PS|19|10|Timor Domini mundus, permanens in saeculum saeculi;iudicia Domini vera, iusta omnia simul,
PS|19|11|desiderabilia super aurum et lapidem pretiosum multum,et dulciora super mel et favum stillantem.
PS|19|12|Etenim servus tuus eruditur in eis;in custodiendis illis retributio multa.
PS|19|13|Errores quis intellegit?Ab occultis munda me
PS|19|14|et a superbia custodi servum tuum, ne dominetur mei,Tunc immaculatus eroet emundabor a delicto maximo.
PS|19|15|Sint ut complaceant eloquia oris mei,et meditatio cordis mei in conspectu tuo.Domine, adiutor meus et redemptor meus.
PS|20|1|Magistro chori. PSALMUS. David.
PS|20|2|Exaudiat te Dominus in die tribulationis,protegat te nomen Dei Iacob.
PS|20|3|Mittat tibi auxilium de sanctoet de Sion tueatur te.
PS|20|4|Memor sit omnis sacrificii tuiet holocaustum tuum pingue habeat.
PS|20|5|Tribuat tibi secundum cor tuumet omne consilium tuum adimpleat.
PS|20|6|Laetabimur in salutari tuoet in nomine Dei nostri levabimus signa;impleat Dominus omnes petitiones tuas.
PS|20|7|Nunc cognovi quoniam salvum fecit Dominus christum suum:exaudivit illum de caelo sancto suo,in virtutibus salutis dexterae eius.
PS|20|8|Hi in curribus, et hi in equis,nos autem nomen Domini Dei nostri invocavimus.
PS|20|9|Ipsi incurvati sunt et ceciderunt,nos autem surreximus et erecti sumus.
PS|20|10|Domine, salvum fac regem,et exaudi nos in die, qua invocaverimus te.
PS|21|1|Magistro chori. PSALMUS. David.
PS|21|2|Domine, in virtute tua laetabitur rexet super salutare tuum exsultabit vehementer.
PS|21|3|Desiderium cordis eius tribuisti eiet voluntatem labiorum eius non denegasti.
PS|21|4|Quoniam praevenisti eum in benedictionibus dulcedinis;posuisti in capite eius coronam de auro purissimo.
PS|21|5|Vitam petiit a te, et tribuisti eilongitudinem dierum in saeculum et in saeculum saeculi.
PS|21|6|Magna est gloria eius in salutari tuo,magnificentiam et decorem impones super eum;
PS|21|7|quoniam pones eum benedictionem in saeculum saeculi,laetificabis eum in gaudio ante vultum tuum.
PS|21|8|Quoniam rex sperat in Dominoet in misericordia Altissimi non commovebitur.
PS|21|9|Inveniet manus tua omnes inimicos tuos,dextera tua inveniet, qui te oderunt.
PS|21|10|Pones eos ut clibanum ignis in tempore vultus tui:Dominus in ira sua deglutiet eos,et devorabit eos ignis.
PS|21|11|Fructum eorum de terra perdeset semen eorum de filiis hominum.
PS|21|12|Quoniam intenderunt in te mala,cogitaverunt consilia: nihil potuerunt.
PS|21|13|Quoniam pones eos dorsum,arcus tuos tendes in vultum eorum.
PS|21|14|Exaltare, Domine, in virtute tua;cantabimus et psallemus virtutes tuas.
PS|22|1|Magistro chori. Ad modum cantici " Cerva diluculo ". PSALMUS. David.
PS|22|2|Deus, Deus meus, quare me dereliquisti?Longe a salute mea verba rugitus mei.
PS|22|3|Deus meus, clamo per diem, et non exaudis,et nocte, et non est requies mihi.
PS|22|4|Tu autem sanctus es,qui habitas in laudibus Israel.
PS|22|5|In te speraverunt patres nostri,speraverunt, et liberasti eos;
PS|22|6|ad te clamaverunt et salvi facti sunt,in te speraverunt et non sunt confusi.
PS|22|7|Ego autem sum vermis et non homo,opprobrium hominum et abiectio plebis.
PS|22|8|Omnes videntes me deriserunt me;torquentes labia moverunt caput:
PS|22|9|" Speravit in Domino: eripiat eum,salvum faciat eum, quoniam vult eum ".
PS|22|10|Quoniam tu es qui extraxisti me de ventre,spes mea ad ubera matris meae.
PS|22|11|In te proiectus sum ex utero,de ventre matris meae Deus meus es tu.
PS|22|12|Ne longe fias a me,quoniam tribulatio proxima est,quoniam non est qui adiuvet.
PS|22|13|Circumdederunt me vituli multi,tauri Basan obsederunt me.
PS|22|14|Aperuerunt super me os suumsicut leo rapiens et rugiens.
PS|22|15|Sicut aqua effusus sum,et dissoluta sunt omnia ossa mea.Factum est cor meum tamquam ceraliquescens in medio ventris mei.
PS|22|16|Aruit tamquam testa palatum meum,et lingua mea adhaesit faucibus meis,et in pulverem mortis deduxisti me.
PS|22|17|Quoniam circumdederunt me canes multi,concilium malignantium obsedit me.Foderunt manus meas et pedes meos,
PS|22|18|et dinumeravi omnia ossa mea.Ipsi vero consideraverunt et inspexerunt me;
PS|22|19|diviserunt sibi vestimenta meaet super vestem meam miserunt sortem.
PS|22|20|Tu autem, Domine, ne elongaveris;fortitudo mea, ad adiuvandum me festina.
PS|22|21|Erue a framea animam meamet de manu canis unicam meam.
PS|22|22|Salva me ex ore leoniset a cornibus unicornium humilitatem meam.
PS|22|23|Narrabo nomen tuum fratribus meis,in medio ecclesiae laudabo te.
PS|22|24|Qui timetis Dominum, laudate eum;universum semen Iacob, glorificate eum.Metuat eum omne semen Israel,
PS|22|25|quoniam non sprevit neque despexit afflictionem pauperisnec avertit faciem suam ab eoet, cum clamaret ad eum, exaudivit.
PS|22|26|Apud te laus mea in ecclesia magna; vota mea reddam in conspectu timentium eum.
PS|22|27|Edent pauperes et saturabuntur;et laudabunt Dominum, qui requirunt eum: Vivant corda eorum in saeculum saeculi! ".
PS|22|28|Reminiscentur et convertentur ad Dominumuniversi fines terrae,et adorabunt in conspectu eiusuniversae familiae gentium.
PS|22|29|Quoniam Domini est regnum,et ipse dominabitur gentium.
PS|22|30|Ipsum solum adorabunt omnes, qui dormiunt in terra;in conspectu eius procident omnes, qui descendunt in pulverem.Anima autem mea illi vivet,
PS|22|31|et semen meum serviet ipsi.Narrabitur de Domino generationi venturae;
PS|22|32|et annuntiabunt iustitiam eiuspopulo, qui nascetur: " Haec fecit Dominus! ".
PS|23|1|PSALMUS. David.Dominus pascit me, et nihil mihi deerit:
PS|23|2|in pascuis virentibus me collocavit,super aquas quietis eduxit me,
PS|23|3|animam meam refecit.Deduxit me super semitas iustitiae propter nomen suum.
PS|23|4|Nam et si ambulavero in valle umbrae mortis,non timebo mala, quoniam tu mecum es.Virga tua et baculus tuus,ipsa me consolata sunt.
PS|23|5|Parasti in conspectu meo mensamadversus eos, qui tribulant me;impinguasti in oleo caput meum,et calix meus redundat.
PS|23|6|Etenim benignitas et misericordia subsequentur meomnibus diebus vitae meae,et inhabitabo in domo Dominiin longitudinem dierum.
PS|24|1|David. PSALMUS.Domini est terra, et plenitudo eius,orbis terrarum, et qui habitant in eo.
PS|24|2|Quia ipse super maria fundavit eumet super flumina firmavit eum. -
PS|24|3|Quis ascendet in montem Domini,aut quis stabit in loco sancto eius?
PS|24|4|Innocens manibus et mundo corde,qui non levavit ad vana animam suamnec iuravit in dolum.
PS|24|5|Hic accipiet benedictionem a Dominoet iustificationem a Deo salutari suo.
PS|24|6|Haec est generatio quaerentium eum,quaerentium faciem Dei Iacob.
PS|24|7|Attollite, portae, capita vestra,et elevamini, portae aeternales,et introibit rex gloriae.
PS|24|8|Quis est iste rex gloriae?Dominus fortis et potens,Dominus potens in proelio.
PS|24|9|Attollite, portae, capita vestra,et elevamini, portae aeternales,et introibit rex gloriae.
PS|24|10|Quis est iste rex gloriae?Dominus virtutum ipse est rex gloriae.
PS|25|1|David.ALEPH. Ad te, Domine, levavi animam meam,
PS|25|2|BETH. Deus meus, in te confido; non erubescam.Neque exsultent super me inimici mei,
PS|25|3|GHIMEL. etenim universi, qui sustinent te, non confundentur.Confundantur infideliter agentes propter vanitatem.
PS|25|4|DALETH. Vias tuas, Domine, demonstra mihiet semitas tuas edoce me.
PS|25|5|HE. Dirige me in veritate tua et doce me,quia tu es Deus salutis meae,VAU. et te sustinui tota die.
PS|25|6|ZAIN. Reminiscere miserationum tuarum, Domine,et misericordiarum tuarum, quoniam a saeculo sunt.
PS|25|7|HETH. Peccata iuventutis meae et delicta mea ne memineris;secundum misericordiam tuam memento mei tu,propter bonitatem tuam, Domine.
PS|25|8|TETH. Dulcis et rectus Dominus,propter hoc peccatores viam docebit;
PS|25|9|IOD. diriget mansuetos in iudicio,docebit mites vias suas.
PS|25|10|CAPH. Universae viae Domini misericordia et veritascustodientibus testamentum eius et testimonia eius.
PS|25|11|LAMED. Propter nomen tuum, Domine,propitiaberis peccato meo: multum est enim.
PS|25|12|MEM. Quis est homo, qui timet Dominum?Docebit eum viam, quam eligat.
PS|25|13|NUN. Anima eius in bonis demorabitur,et semen eius hereditabit terram.
PS|25|14|SAMECH. Familiariter aget Dominus cum timentibus eum,ut testamentum suum manifestet illis.
PS|25|15|AIN. Oculi mei semper ad Dominum,quoniam ipse evellet de laqueo pedes meos.
PS|25|16|PHE. Respice in me et miserere mei,quia unicus et pauper sum ego.
PS|25|17|SADE. Dilata angustias cordis meiet de necessitatibus meis erue me.
PS|25|18|Vide humilitatem meam et laborem meumet dimitte universa delicta mea.
PS|25|19|RES. Respice inimicos meos, quoniam multiplicati suntet odio crudeli oderunt me.
PS|25|20|SIN. Custodi animam meam et erue me;non erubescam, quoniam speravi in te.
PS|25|21|TAU. Innocentia et aequitas custodiant me,quia sustinui te.
PS|25|22|PHE. Libera, Deus, Israelex omnibus tribulationibus suis.
PS|26|1|David.Iudica me, Domine, quoniam ego in innocentia mea ingressus sumet in Domino sperans non infirmabor.
PS|26|2|Proba me, Domine, et tenta me;ure renes meos et cor meum. -
PS|26|3|Quoniam misericordia tua ante oculos meos est,et ambulavi in veritate tua.
PS|26|4|Non sedi cum viris vanitatiset cum occulte agentibus non introibo.
PS|26|5|Odivi ecclesiam malignantiumet cum impiis non sedebo.
PS|26|6|Lavabo in innocentia manus measet circumdabo altare tuum, Domine,
PS|26|7|ut auditas faciam voces laudiset enarrem universa mirabilia tua.
PS|26|8|Domine, dilexi habitaculum domus tuaeet locum habitationis gloriae tuae.
PS|26|9|Ne colligas cum impiis animam meamet cum viris sanguinum vitam meam,
PS|26|10|in quorum manibus iniquitates sunt,dextera eorum repleta est muneribus.
PS|26|11|Ego autem in innocentia mea ingressus sum;redime me et miserere mei.
PS|26|12|Pes meus stetit in directo,in ecclesiis benedicam Domino.
PS|27|1|David.Dominus illuminatio mea et salus mea; quem timebo?Dominus protector vitae meae; a quo trepidabo?
PS|27|2|Dum appropiant super me nocentes,ut edant carnes meas;qui tribulant me et inimici mei,ipsi infirmati sunt et ceciderunt.
PS|27|3|Si consistant adversum me castra,non timebit cor meum;si exsurgat adversum me proelium, in hoc ego sperabo.
PS|27|4|Unum petii a Domino, hoc requiram:ut inhabitem in domo Dominiomnibus diebus vitae meae,ut videam voluptatem Dominiet visitem templum eius.
PS|27|5|Quoniam occultabit me in tentorio suoin die malorum.Abscondet me in abscondito tabernaculi sui,in petra exaltabit me.
PS|27|6|Et nunc exaltatur caput meumsuper inimicos meos in circuitu meo.Immolabo in tabernaculo eius hostias vociferationis,cantabo et psalmum dicam Domino.
PS|27|7|Exaudi, Domine, vocem meam, qua clamavi;miserere mei et exaudi me.
PS|27|8|De te dixit cor meum: " Exquirite faciem meam! ".Faciem tuam, Domine, exquiram.
PS|27|9|Ne avertas faciem tuam a me,ne declines in ira a servo tuo.Adiutor meus es tu, ne me reiciasneque derelinquas me, Deus salutis meae.
PS|27|10|Quoniam pater meus et mater mea dereliquerunt me,Dominus autem assumpsit me.
PS|27|11|Ostende mihi, Domine, viam tuamet dirige me in semitam rectam propter inimicos meos.
PS|27|12|Ne tradideris me in animam tribulantium me,quoniam insurrexerunt in me testes iniqui,et qui violentiam spirant.
PS|27|13|Credo videre bona Domini in terra viventium.
PS|27|14|Exspecta Dominum, viriliter age,et confortetur cor tuum, et sustine Dominum.
PS|28|1|David.Ad te, Domine, clamabo;Deus meus, ne sileas a me.Ne quando taceas a me,et assimilabor descendentibus in lacum.
PS|28|2|Exaudi vocem deprecationis meae, dum clamo ad te,dum extollo manus meas ad templum sanctum tuum.
PS|28|3|Ne simul trahas me cum peccatoribuset cum operantibus iniquitatem.Qui loquuntur pacem cum proximo suo,mala autem in cordibus eorum.
PS|28|4|Da illis secundum opera eorumet secundum nequitiam adinventionum ipsorum.Secundum opus manuum eorum tribue illis,redde retributionem eorum ipsis.
PS|28|5|Quoniam non intellexerunt opera Dominiet opus manuum eius,destruet illos et non aedificabit eos.
PS|28|6|Benedictus Dominus,quoniam exaudivit vocem deprecationis meae;
PS|28|7|Dominus adiutor meus et protector meus,in ipso speravit cor meum, et adiutus sum,et exsultavit cor meum,et in cantico meo confitebor ei.
PS|28|8|Dominus fortitudo plebi suae,et refugium salvationum christi sui est.
PS|28|9|Salvum fac populum tuum et benedic hereditati tuaeet pasce eos et extolle illos usque in aeternum.
PS|29|1|PSALMUS. David.Afferte Domino, filii Dei,afferte Domino gloriam et potentiam,
PS|29|2|afferte Domino gloriam nominis eius,adorate Dominum in splendore sancto.
PS|29|3|Vox Domini super aquas;Deus maiestatis intonuit,Dominus super aquas multas.
PS|29|4|Vox Domini in virtute,vox Domini in magnificentia.
PS|29|5|Vox Domini confringentis cedros;et confringet Dominus cedros Libani.
PS|29|6|Et saltare faciet, tamquam vitulum, Libanum,et Sarion, quemadmodum filium unicornium. -
PS|29|7|Vox Domini intercidentis flammam ignis,
PS|29|8|vox Domini concutientis desertum,et concutiet Dominus desertum Cades.
PS|29|9|Vox Domini properantis partum cervarum,et denudabit condensa;et in templo eius omnes dicent gloriam.
PS|29|10|Dominus super diluvium habitat,et sedebit Dominus rex in aeternum.
PS|29|11|Dominus virtutem populo suo dabit,Dominus benedicet populo suo in pace.
PS|30|1|PSALMUS. Canticum festi Dedicationis Templi. David.
PS|30|2|Exaltabo te, Domine, quoniam extraxisti menec delectasti inimicos meos super me.
PS|30|3|Domine Deus meus, clamavi ad te, et sanasti me.
PS|30|4|Domine, eduxisti ab inferno animam meam,vivificasti me, ut non descenderem in lacum.
PS|30|5|Psallite Domino, sancti eius,et confitemini memoriae sanctitatis eius,
PS|30|6|quoniam ad momentum indignatio eius,et per vitam voluntas eius.Ad vesperum demoratur fletus,ad matutinum laetitia.
PS|30|7|Ego autem dixi in securitate mea: Non movebor in aeternum ".
PS|30|8|Domine, in voluntate tuapraestitisti decori meo virtutem;avertisti faciem tuam a me,et factus sum conturbatus.
PS|30|9|Ad te, Domine, clamabamet ad Deum meum deprecabar.
PS|30|10|Quae utilitas in sanguine meo,dum descendo in corruptionem?Numquid confitebitur tibi pulvisaut annuntiabit veritatem tuam?
PS|30|11|Audivit Dominus et misertus est mei,Dominus factus est adiutor meus.
PS|30|12|Convertisti planctum meum in choros mihi,conscidisti saccum meum et accinxisti me laetitia,
PS|30|13|ut cantet tibi gloria mea et non taceat.Domine Deus meus, in aeternum confitebor tibi.
PS|31|1|Magistro chori. PSALMUS. David.
PS|31|2|In te, Domine, speravi, non confundar in aeternum;in iustitia tua libera me.
PS|31|3|Inclina ad me aurem tuam,accelera, ut eruas me.Esto mihi in rupem praesidiiet in domum munitam, ut salvum me facias.
PS|31|4|Quoniam fortitudo mea et refugium meum es tuet propter nomen tuum deduces me et pasces me.
PS|31|5|Educes me de laqueo, quem absconderunt mihi,quoniam tu es fortitudo mea.
PS|31|6|In manus tuas commendo spiritum meum;redemisti me, Domine, Deus veritatis.
PS|31|7|Odisti observantes vanitates supervacuas,ego autem in Domino speravi.
PS|31|8|Exsultabo et laetabor in misericordia tua,quoniam respexisti humilitatem meam;agnovisti necessitates animae meae
PS|31|9|nec conclusisti me in manibus inimici;statuisti in loco spatioso pedes meos.
PS|31|10|Miserere mei, Domine, quoniam tribulor;conturbatus est in maerore oculus meus,anima mea et venter meus.
PS|31|11|Quoniam defecit in dolore vita mea,et anni mei in gemitibus;infirmata est in paupertate virtus mea,et ossa mea contabuerunt.
PS|31|12|Apud omnes inimicos meos factus sum opprobriumet vicinis meis valde et timor notis meis:qui videbant me foras, fugiebant a me.
PS|31|13|Oblivioni a corde datus sum tamquam mortuus;factus sum tamquam vas perditum.
PS|31|14|Quoniam audivi vituperationem multorum: horror in circuitu;in eo dum convenirent simul adversum me,auferre animam meam consiliati sunt.
PS|31|15|Ego autem in te speravi, Domine;dixi: " Deus meus es tu,
PS|31|16|in manibus tuis sortes meae ".Eripe me de manu inimicorum meorumet a persequentibus me;
PS|31|17|illustra faciem tuam super servum tuum,salvum me fac in misericordia tua.
PS|31|18|Domine, non confundar, quoniam invocavi te;erubescant impii et obmutescant in inferno.
PS|31|19|Muta fiant labia dolosa,quae loquuntur adversus iustum protervain superbia et in abusione.
PS|31|20|Quam magna multitudo dulcedinis tuae, Domine,quam abscondisti timentibus te.Perfecisti eis, qui sperant in te,in conspectu filiorum hominum.
PS|31|21|Abscondes eos in abscondito faciei tuaea conturbatione hominum;proteges eos in tabernaculoa contradictione linguarum.
PS|31|22|Benedictus Dominus,quoniam mirificavit misericordiam suam mihi in civitate munita.
PS|31|23|Ego autem dixi in trepidatione mea: Praecisus sum a conspectu oculorum tuorum ".Verumtamen exaudisti vocem orationis meae,dum clamarem ad te.
PS|31|24|Diligite Dominum, omnes sancti eius:fideles conservat Dominuset retribuit abundanter facientibus superbiam.
PS|31|25|Viriliter agite, et confortetur cor vestrum,omnes, qui speratis in Domino.
PS|32|1|David. Maskil.Beatus, cui remissa est iniquitas,et obtectum est peccatum.
PS|32|2|Beatus vir, cui non imputavit Dominus delictum,nec est in spiritu eius dolus.
PS|32|3|Quoniam tacui, inveteraverunt ossa mea,dum rugirem tota die.
PS|32|4|Quoniam die ac nocte gravata est super me manus tua,immutatus est vigor meus in ardoribus aestatis.
PS|32|5|Peccatum meum cognitum tibi feciet delictum meum non abscondi.Dixi: " Confitebor adversum me iniquitatem meam Domino ".Et tu remisisti impietatem peccati mei.
PS|32|6|Propter hoc orabit ad te omnis sanctus in tempore opportuno.Et in diluvio aquarum multarumad eum non approximabunt.
PS|32|7|Tu es refugium meum, a tribulatione conservabis me;exsultationibus salutis circumdabis me.
PS|32|8|Intellectum tibi dabo et instruam te in via, qua gradieris;firmabo super te oculos meos.
PS|32|9|Nolite fieri sicut equus et mulus,quibus non est intellectus;in camo et freno si accedis ad constringendum,non approximant ad te.
PS|32|10|Multi dolores impii,sperantem autem in Domino misericordia circumdabit.
PS|32|11|Laetamini in Domino et exsultate, iusti;et gloriamini, omnes recti corde.
PS|33|1|Exsultate, iusti, in Domino;rectos decet collaudatio.
PS|33|2|Confitemini Domino in cithara,in psalterio decem chordarum psallite illi.
PS|33|3|Cantate ei canticum novum,bene psallite ei in vociferatione,
PS|33|4|quia rectum est verbum Domini,et omnia opera eius in fide.
PS|33|5|Diligit iustitiam et iudicium;misericordia Domini plena est terra.
PS|33|6|Verbo Domini caeli facti sunt,et spiritu oris eius omnis virtus eorum.
PS|33|7|Congregans sicut in utre aquas maris,ponens in thesauris abyssos.
PS|33|8|Timeat Dominum omnis terra,a facie autem eius formident omnes inhabitantes orbem.
PS|33|9|Quoniam ipse dixit, et facta sunt,ipse mandavit, et creata sunt.
PS|33|10|Dominus dissipat consilia gentium,irritas facit cogitationes populorum.
PS|33|11|Consilium autem Domini in aeternum manet,cogitationes cordis eius in generatione et generationem.
PS|33|12|Beata gens, cui Dominus est Deus,populus, quem elegit in hereditatem sibi.
PS|33|13|De caelo respexit Dominus,vidit omnes filios hominum.
PS|33|14|De loco habitaculi sui respexitsuper omnes, qui habitant terram,
PS|33|15|qui finxit singillatim corda eorum,qui intellegit omnia opera eorum.
PS|33|16|Non salvatur rex per multam virtutem,et gigas non liberabitur in multitudine virtutis suae.
PS|33|17|Fallax equus ad salutem,in abundantia autem virtutis suae non salvabit.
PS|33|18|Ecce oculi Domini super metuentes eum,in eos, qui sperant super misericordia eius,
PS|33|19|ut eruat a morte animas eorumet alat eos in fame.
PS|33|20|Anima nostra sustinet Dominum,quoniam adiutor et protector noster est;
PS|33|21|quia in eo laetabitur cor nostrum,et in nomine sancto eius speravimus.
PS|33|22|Fiat misericordia tua, Domine, super nos,quemadmodum speravimus in te.
PS|34|1|David, quando se mente alienatum simulavitcoram Abimelech et, ab illo dimissus, abiit.
PS|34|2|ALEPH. Benedicam Dominum in omni tempore,semper laus eius in ore meo.
PS|34|3|BETH. In Domino gloriabitur anima mea,audiant mansueti et laetentur.
PS|34|4|GHIMEL. Magnificate Dominum mecum,et exaltemus nomen eius in idipsum.
PS|34|5|DALETH. Exquisivi Dominum, et exaudivit meet ex omnibus terroribus meis eripuit me.
PS|34|6|HE. Respicite ad eum, et illuminamini,et facies vestrae non confundentur.
PS|34|7|ZAIN. Iste pauper clamavit, et Dominus exaudivit eumet de omnibus tribulationibus eius salvavit eum.
PS|34|8|HETH. Vallabit angelus Domini in circuitu timentes eumet eripiet eos.
PS|34|9|TETH. Gustate et videte quoniam suavis est Dominus;beatus vir, qui sperat in eo.
PS|34|10|IOD. Timete Dominum, sancti eius,quoniam non est inopia timentibus eum.
PS|34|11|CAPH. Divites eguerunt et esurierunt,inquirentes autem Dominum non deficient omni bono.
PS|34|12|LAMED. Venite, filii, audite me:timorem Domini docebo vos.
PS|34|13|MEM. Quis est homo, qui vult vitam,diligit dies, ut videat bonum? -
PS|34|14|NUN. Prohibe linguam tuam a malo,et labia tua, ne loquantur dolum.
PS|34|15|SAMECH. Diverte a malo et fac bonum,inquire pacem et persequere eam.
PS|34|16|AIN. Oculi Domini super iustos,et aures eius in clamorem eorum.
PS|34|17|PHE. Vultus autem Domini super facientes mala,ut perdat de terra memoriam eorum.
PS|34|18|SADE. Clamaverunt, et Dominus exaudivitet ex omnibus tribulationibus eorum liberavit eos.
PS|34|19|COPH. Iuxta est Dominus iis, qui contrito sunt corde,et confractos spiritu salvabit.
PS|34|20|RES. Multae tribulationes iustorum,et de omnibus his liberabit eos Dominus.
PS|34|21|SIN. Custodit omnia ossa eorum,unum ex his non conteretur.
PS|34|22|TAU. Interficiet peccatorem malitia;et, qui oderunt iustum, punientur.
PS|34|23|PHE. Redimet Dominus animas servorum suorum;et non punientur omnes, qui sperant in eo.
PS|35|1|David.Iudica, Domine, iudicantes me;impugna impugnantes me.
PS|35|2|Apprehende clipeum et scutumet exsurge in adiutorium mihi.
PS|35|3|Effunde frameam et securimadversus eos, qui persequuntur me.Dic animae meae: " Salus tua ego sum ".
PS|35|4|Confundantur et revereanturquaerentes animam meam;avertantur retrorsum et confundanturcogitantes mihi mala.
PS|35|5|Fiant tamquam pulvis ante ventum,et angelus Domini impellens eos;
PS|35|6|fiat via illorum tenebrae et lubricum,et angelus Domini persequens eos.
PS|35|7|Quoniam gratis absconderunt mihi laqueum suum,gratis foderunt foveam animae meae.
PS|35|8|Veniat illi calamitas, quam ignorat,et captio, quam abscondit, apprehendat eum,et in eandem calamitatem ipse cadat.
PS|35|9|Anima autem mea exsultabit in Dominoet delectabitur super salutari suo.
PS|35|10|Omnia ossa mea dicent: Domine, quis similis tibi?Eripiens inopem de manu fortiorum eius,egenum et pauperem a diripientibus eum ".
PS|35|11|Surgentes testes iniqui,quae ignorabam, interrogabant me;
PS|35|12|retribuebant mihi mala pro bonis,desolatio est animae meae.
PS|35|13|Ego autem, cum infirmarentur,induebar cilicio,humiliabam in ieiunio animam meam;et oratio mea in sinu meo convertebatur.
PS|35|14|Quasi pro proximo et quasi pro fratre meo ambulabam,quasi lugens matrem contristatus incurvabar.
PS|35|15|Cum autem vacillarem, laetati sunt et convenerunt;convenerunt contra me percutientes, et ignoravi.
PS|35|16|Diripuerunt et non desistebant;tentaverunt me, subsannaverunt me subsannatione,frenduerunt super me dentibus suis.
PS|35|17|Domine, quamdiu aspicies?Restitue animam meam a malignitate eorum,a leonibus unicam meam.
PS|35|18|Confitebor tibi in ecclesia magna,in populo multo laudabo te.
PS|35|19|Non supergaudeant mihi inimici mei mendaces,qui oderunt me gratis et annuunt oculis.
PS|35|20|Etenim non pacifice loquebanturet contra mansuetos terrae dolos cogitabant.
PS|35|21|Et dilataverunt super me os suum;dixerunt: " Euge, euge, viderunt oculi nostri ". -
PS|35|22|Vidisti, Domine, ne sileas;Domine, ne discedas a me.
PS|35|23|Exsurge et evigila ad iudicium meum,Deus meus et Dominus meus, ad causam meam.
PS|35|24|Iudica me secundum iustitiam tuam, Domine Deus meus,et non supergaudeant mihi.
PS|35|25|Non dicant in cordibus suis: Euge animae nostrae ";nec dicant: " Devoravimus eum ".
PS|35|26|Erubescant et revereantur simul, qui gratulantur malis meis;induantur confusione et reverentia, qui magna loquuntur super me
PS|35|27|Exsultent et laetentur, qui volunt iustitiam meam,et dicant semper: " Magnificetur Dominus,qui vult pacem servi sui ".
PS|35|28|Et lingua mea meditabitur iustitiam tuam,tota die laudem tuam.
PS|36|1|Magistro chori. David, servi Domini.
PS|36|2|Susurrat iniquitas ad impium in medio cordis eius;non est timor Dei ante oculos eius.
PS|36|3|Quoniam blanditur ipsi in conspectu eius,ut non inveniat iniquitatem suam et oderit.
PS|36|4|Verba oris eius iniquitas et dolus,desiit intellegere, ut bene ageret.
PS|36|5|Iniquitatem meditatus est in cubili suo,astitit omni viae non bonae,malitiam autem non odivit.
PS|36|6|Domine, in caelo misericordia tua,et veritas tua usque ad nubes;
PS|36|7|iustitia tua sicut montes Dei,iudicia tua abyssus multa:homines et iumenta salvabis, Domine.
PS|36|8|Quam pretiosa misericordia tua, Deus!Filii autem hominum in tegmine alarum tuarum sperabunt;
PS|36|9|inebriabuntur ab ubertate domus tuae,et torrente voluptatis tuae potabis eos.
PS|36|10|Quoniam apud te est fons vitae,et in lumine tuo videbimus lumen.
PS|36|11|Praetende misericordiam tuam scientibus teet iustitiam tuam his, qui recto sunt corde.
PS|36|12|Non veniat mihi pes superbiae,et manus peccatoris non moveat me.
PS|36|13|Ibi ceciderunt, qui operantur iniquitatem,expulsi sunt nec potuerunt stare.
PS|37|1|David.ALEPH. Noli aemulari in malignantibusneque zelaveris facientes iniquitatem,
PS|37|2|quoniam tamquam fenum velociter arescentet quemadmodum herba virens decident.
PS|37|3|BETH. Spera in Domino et fac bonitatem,et inhabitabis terram et pasceris in fide.
PS|37|4|Delectare in Domino,et dabit tibi petitiones cordis tui.
PS|37|5|GHIMEL. Committe Domino viam tuam et spera in eo,et ipse faciet;
PS|37|6|et educet quasi lumen iustitiam tuamet iudicium tuum tamquam meridiem.
PS|37|7|DALETH. Quiesce in Domino et exspecta eum;noli aemulari in eo, qui prosperatur in via sua,in homine, qui molitur insidias.
PS|37|8|HE. Desine ab ira et derelinque furorem,noli aemulari, quod vertit ad malum,
PS|37|9|quoniam qui malignantur, exterminabuntur,sustinentes autem Dominum ipsi hereditabunt terram.
PS|37|10|VAU. Et adhuc pusillum et non erit peccator,et quaeres locum eius et non invenies.
PS|37|11|Mansueti autem hereditabunt terramet delectabuntur in multitudine pacis.
PS|37|12|ZAIN. Insidiabitur peccator iustoet stridebit super eum dentibus suis.
PS|37|13|Dominus autem irridebit eum,quoniam prospicit quod veniet dies eius.
PS|37|14|HETH. Gladium evaginaverunt peccatores,intenderunt arcum suum,ut deiciant pauperem et inopem,ut trucident recte ambulantes in via.
PS|37|15|Gladius eorum intrabit in corda ipsorum,et arcus eorum confringetur.
PS|37|16|TETH. Melius est modicum iustosuper divitias peccatorum multas,
PS|37|17|quoniam brachia peccatorum conterentur,confirmat autem iustos Dominus.
PS|37|18|IOD. Novit Dominus dies immaculatorum,et hereditas eorum in aeternum erit.
PS|37|19|Non confundentur in tempore maloet in diebus famis saturabuntur.
PS|37|20|CAPH. Quia peccatores peribunt,inimici vero Domini ut decor camporum deficient,quemadmodum fumus deficient.
PS|37|21|LAMED. Mutuatur peccator et non solvet,iustus autem miseretur et tribuet.
PS|37|22|Quia benedicti eius hereditabunt terram,maledicti autem eius exterminabuntur.
PS|37|23|MEM. A Domino gressus hominis confirmantur,et viam eius volet.
PS|37|24|Cum ceciderit, non collidetur,quia Dominus sustentat manum eius.
PS|37|25|NUN. Iunior fui et senuiet non vidi iustum derelictumnec semen eius quaerens panem.
PS|37|26|Tota die miseretur et commodat,et semen illius in benedictione erit.
PS|37|27|SAMECH. Declina a malo et fac bonum,et inhabitabis in saeculum saeculi,
PS|37|28|quia Dominus amat iudiciumet non derelinquet sanctos suos.AIN. Iniusti in aeternum disperibunt,et semen impiorum exterminabitur.
PS|37|29|Iusti autem hereditabunt terramet inhabitabunt in saeculum saeculi super eam.
PS|37|30|PHE. Os iusti meditabitur sapientiam,et lingua eius loquetur iudicium;
PS|37|31|lex Dei eius in corde ipsius,et non vacillabunt gressus eius.
PS|37|32|SADE. Considerat peccator iustumet quaerit mortificare eum;
PS|37|33|Dominus autem non derelinquet eum in manibus eiusnec damnabit eum, cum iudicabitur illi.
PS|37|34|COPH. Exspecta Dominum et custodi viam eius,et exaltabit te, ut hereditate capias terram;cum exterminabuntur peccatores, videbis.
PS|37|35|RES. Vidi impium superexaltatumet elevatum sicut cedrum virentem;
PS|37|36|et transivi, et ecce non erat,et quaesivi eum, et non est inventus.
PS|37|37|SIN. Observa innocentiam et vide aequitatem,quoniam est posteritas homini pacifico.
PS|37|38|Iniusti autem disperibunt simul,posteritas impiorum exterminabitur.
PS|37|39|TAU. Salus autem iustorum a Domino,et protector eorum in tempore tribulationis.
PS|37|40|Et adiuvabit eos Dominus et liberabit eoset eruet eos a peccatoribus et salvabit eos,quia speraverunt in eo.
PS|38|1|PSALMUS. David. Ad commemorandum.
PS|38|2|Domine, ne in furore tuo arguas meneque in ira tua corripias me,
PS|38|3|quoniam sagittae tuae infixae sunt mihi,et descendit super me manus tua.
PS|38|4|Non est sanitas in carne mea a facie indignationis tuae,non est pax ossibus meis a facie peccatorum meorum.
PS|38|5|Quoniam iniquitates meae supergressae sunt caput meumet sicut onus grave gravant me nimis. -
PS|38|6|Putruerunt et corrupti sunt livores meia facie insipientiae meae.
PS|38|7|Inclinatus sum et incurvatus nimis;tota die contristatus ingrediebar.
PS|38|8|Quoniam lumbi mei impleti sunt ardoribus,et non est sanitas in carne mea.
PS|38|9|Afflictus sum et humiliatus sum nimis,rugiebam a gemitu cordis mei.
PS|38|10|Domine, ante te omne desiderium meum,et gemitus meus a te non est absconditus.
PS|38|11|Palpitavit cor meum, dereliquit me virtus mea,et lumen oculorum meorum, et ipsum non est mecum.
PS|38|12|Amici mei et proximi meiprocul a plaga mea steterunt,et propinqui mei de longe steterunt.
PS|38|13|Et laqueos posuerunt, qui quaerebant animam meam;et, qui requirebant mala mihi, locuti sunt insidiaset dolos tota die meditabantur.
PS|38|14|Ego autem tamquam surdus non audiebamet sicut mutus non aperiens os suum;
PS|38|15|et factus sum sicut homo non audienset non habens in ore suo redargutiones.
PS|38|16|Quoniam in te, Domine, speravi,tu exaudies, Domine Deus meus.
PS|38|17|Quia dixi: "Ne quando supergaudeant mihi;dum commoventur pedes mei,magnificantur super me ".
PS|38|18|Quoniam ego in lapsum paratus sum,et dolor meus in conspectu meo semper.
PS|38|19|Quoniam iniquitatem meam annuntiaboet sollicitus sum de peccato meo.
PS|38|20|Inimici autem mei vivunt et confirmati sunt;et multiplicati sunt, qui oderunt me inique.
PS|38|21|Retribuentes mala pro bonis detrahebant mihi,pro eo quod sequebar bonitatem.
PS|38|22|Ne derelinquas me, Domine;Deus meus, ne discesseris a me.
PS|38|23|Festina in adiutorium meum,Domine, salus mea.
PS|39|1|Magistro chori, Idithun. PSALMUS. David.
PS|39|2|Dixi: " Custodiam vias meas,ut non delinquam in lingua mea;ponam ori meo custodiam,donec consistit peccator adversum me ".
PS|39|3|Tacens obmutui et silui absque ullo bono,et dolor meus renovatus est.
PS|39|4|Concaluit cor meum intra me,et in meditatione mea exarsit ignis.
PS|39|5|Locutus sum in lingua mea: Notum fac mihi, Domine, finem meum;et numerum dierum meorum quis est,ut sciam quam brevis sit vita mea ".
PS|39|6|Ecce paucorum palmorum fecisti dies meos,et spatium vitae meae tamquam nihilum ante te.Etenim universa vanitas omnis homo constitutus est.
PS|39|7|Etenim ut imago pertransit homo.Etenim vanitas est et concitatur;thesaurizat et ignorat quis congregabit ea.
PS|39|8|Et nunc quae est exspectatio mea, Domine?Spes mea apud te est.
PS|39|9|Ab omnibus iniquitatibus meis erue me,opprobrium insipienti ne ponas me.
PS|39|10|Obmutui et non aperiam os meum,quoniam tu fecisti.
PS|39|11|Amove a me plagas tuas:ab ictu manus tuae ego defeci.
PS|39|12|In increpationibus, propter iniquitatem, corripuisti hominem,et tabescere fecisti, sicut tinea, desiderabilia eius.Etenim vanitas omnis homo.
PS|39|13|Exaudi orationem meam, Domine,et clamorem meum auribus percipe.Ad lacrimas meas ne obsurdescas,quoniam advena ego sum apud te,peregrinus sicut omnes patres mei.
PS|39|14|Avertere a me, ut refrigerer,priusquam abeam et non sim amplius.
PS|40|1|Magistro chori. David. PSALMUS.
PS|40|2|Exspectans exspectavi Dominum,et intendit mihi.
PS|40|3|Et exaudivit clamorem meumet eduxit me de lacu miseriae et de luto faecis;et statuit super petram pedes meoset firmavit gressus meos.
PS|40|4|Et immisit in os meum canticum novum,carmen Deo nostro.Videbunt multi et timebuntet sperabunt in Domino.
PS|40|5|Beatus vir, qui posuit Dominum spem suamet non respexit superbos et declinantes in mendacium.
PS|40|6|Multa fecisti tu, Domine Deus meus, mirabilia tua,et cogitationes tuas pro nobis: non est qui similis sit tibi.Si nuntiare et eloqui voluero,multiplicabuntur super numerum.
PS|40|7|Sacrificium et oblationem noluisti,aures autem fodisti mihi.Holocaustum et pro peccato non postulasti,
PS|40|8|tunc dixi: " Ecce venio.In volumine libri scriptum est de me.
PS|40|9|Facere voluntatem tuam,Deus meus, volui;et lex tua in praecordiis meis ".
PS|40|10|Annuntiavi iustitiam tuam in ecclesia magna;ecce labia mea non prohibebo, Domine, tu scisti.
PS|40|11|Iustitiam tuam non abscondi in corde meo,veritatem tuam et salutare tuum dixi.Non abscondi misericordiam tuamet veritatem tuam ab ecclesia magna.
PS|40|12|Tu autem, Domine, ne prohibeas miserationes tuas a me;misericordia tua et veritas tua semper suscipiant me,
PS|40|13|quoniam circumdederunt me mala, quorum non est numerus;comprehenderunt me iniquitates meae,et non potui videre.Multiplicatae sunt super capillos capitis mei,et cor meum dereliquit me.
PS|40|14|Complaceat tibi, Domine, ut eruas me;Domine, ad adiuvandum me festina.
PS|40|15|Confundantur et revereantur simul,qui quaerunt animam meam, ut auferant eam.Avertantur retrorsum et erubescant,qui volunt mihi mala.
PS|40|16|Obstupescant propter confusionem suam,qui dicunt mihi: " Euge, euge ".
PS|40|17|Exsultent et laetentur in te omnes quaerentes te;et dicant semper: " Magnificetur Dominus ",qui diligunt salutare tuum.
PS|40|18|Ego autem egenus et pauper sum;Dominus sollicitus est mei.Adiutor meus et liberator meus tu es;Deus meus, ne tardaveris.
PS|41|1|Magistro chori. PSALMUS. David.
PS|41|2|Beatus, qui intellegit de egeno;in die mala liberabit eum Dominus.
PS|41|3|Dominus servabit eum et vivificabit eumet beatum faciet eum in terraet non tradet eum in animam inimicorum eius.
PS|41|4|Dominus opem feret illi super lectum doloris eius;universum stratum eius versabis in infirmitate eius.
PS|41|5|Ego dixi: " Domine, miserere mei;sana animam meam, quia peccavi tibi ".
PS|41|6|Inimici mei dixerunt mala mihi: Quando morietur, et peribit nomen eius? ".
PS|41|7|Et si ingrediebatur, ut visitaret, vana loquebatur;cor eius congregabat iniquitatem sibi,egrediebatur foras et detrahebat.
PS|41|8|Simul adversum me susurrabant omnes inimici mei;adversum me cogitabant mala mihi:
PS|41|9|" Maleficium effusum est in eo;et, qui decumbit, non adiciet ut resurgat ".
PS|41|10|Sed et homo pacis meae, in quo speravi,qui edebat panem meum, levavit contra me calcaneum.
PS|41|11|Tu autem, Domine, miserere meiet resuscita me, et retribuam eis.
PS|41|12|In hoc cognovi quoniam voluisti me,quia non gaudebit inimicus meus super me;
PS|41|13|me autem propter innocentiam suscepistiet statuisti me in conspectu tuo in aeternum.
PS|41|14|Benedictus Dominus, Deus Israel,a saeculo et usque in saeculum. Fiat, fiat.
PS|42|1|Magistro chori. Maskil. Filiorum Core.
PS|42|2|Quemadmodum desiderat cervus ad fontes aquarum,ita desiderat anima mea ad te, Deus.
PS|42|3|Sitivit anima mea ad Deum, Deum vivum;quando veniam et apparebo ante faciem Dei?
PS|42|4|Fuerunt mihi lacrimae meae panis die ac nocte,dum dicitur mihi cotidie: " Ubi est Deus tuus? ".
PS|42|5|Haec recordatus sum et effudi in me animam meam;quoniam transibam in locum tabernaculi admirabilisusque ad domum Deiin voce exsultationis et confessionismultitudinis festa celebrantis.
PS|42|6|Quare tristis es, anima mea, et quare conturbaris in me?Spera in Deo, quoniam adhuc confitebor illi,salutare vultus mei et Deus meus.
PS|42|7|In meipso anima mea contristata est;propterea memor ero tuide terra Iordanis et Hermonim, de monte Misar.
PS|42|8|Abyssus abyssum invocat in voce cataractarum tuarum;omnes gurgites tui et fluctus tui super me transierunt.
PS|42|9|In die mandavit Dominus misericordiam suam,et nocte canticum eius apud me est: oratio ad Deum vitae meae.
PS|42|10|Dicam Deo: " Susceptor meus es.Quare oblitus es mei,et quare contristatus incedo,dum affligit me inimicus? ".
PS|42|11|Dum confringuntur ossa mea,exprobraverunt mihi, qui tribulant me,dum dicunt mihi quotidie: " Ubi est Deus tuus? ". -
PS|42|12|Quare tristis es, anima mea, et quare conturbaris in me?Spera in Deo, quoniam adhuc confitebor illi,salutare vultus mei et Deus meus.
PS|43|1|Iudica me, Deus, et discerne causam meam de gente non sancta;ab homine iniquo et doloso erue me.
PS|43|2|Quia tu es Deus refugii mei;quare me reppulisti,et quare tristis incedo, dum affligit me inimicus?
PS|43|3|Emitte lucem tuam et veritatem tuam;ipsae me deducant et adducantin montem sanctum tuum et in tabernacula tua.
PS|43|4|Et introibo ad altare Dei,ad Deum laetitiae exsultationis meae.Confitebor tibi in cithara, Deus, Deus meus.
PS|43|5|Quare tristis es, anima mea, et quare conturbaris in me?Spera in Deo, quoniam adhuc confitebor illi,salutare vultus mei et Deus meus.
PS|44|1|Magistro chori. Filiorum Core. Maskil.
PS|44|2|Deus, auribus nostris audivimus;patres nostri annuntiaverunt nobisopus, quod operatus es in diebus eorum, in diebus antiquis.
PS|44|3|Tu manu tua gentes depulisti et plantasti illos,afflixisti populos et dilatasti eos.
PS|44|4|Nec enim in gladio suo possederunt terram,et brachium eorum non salvavit eos;sed dextera tua et brachium tuumet illuminatio vultus tui,quoniam complacuisti in eis.
PS|44|5|Tu es rex meus et Deus meus,qui mandas salutes Iacob.
PS|44|6|In te inimicos nostros proiecimus,et in nomine tuo conculcavimus insurgentes in nos. -
PS|44|7|Non enim in arcu meo sperabo,et gladius meus non salvabit me.
PS|44|8|Tu autem salvasti nos de affligentibus noset odientes nos confudisti.
PS|44|9|In Deo gloriabimur tota dieet in nomine tuo confitebimur in saeculum.
PS|44|10|Nunc autem reppulisti et confudisti noset non egredieris, Deus, cum virtutibus nostris.
PS|44|11|Convertisti nos retrorsum coram inimicis nostris;et, qui oderunt nos, diripuerunt sibi.
PS|44|12|Dedisti nos tamquam oves ad vescendumet in gentibus dispersisti nos.
PS|44|13|Vendidisti populum tuum sine lucronec ditior factus es in commutatione eorum.
PS|44|14|Posuisti nos opprobrium vicinis nostris,subsannationem et derisum his, qui sunt in circuitu nostro.
PS|44|15|Posuisti nos similitudinem in gentibus,commotionem capitis in populis.
PS|44|16|Tota die verecundia mea contra me est,et confusio faciei meae cooperuit me
PS|44|17|a voce exprobrantis et obloquentis,a facie inimici et ultoris.
PS|44|18|Haec omnia venerunt super nos, nec obliti sumus teet inique non egimus in testamentum tuum.
PS|44|19|Et non recessit retro cor nostrum,nec declinaverunt gressus nostri a via tua;
PS|44|20|sed humiliasti nos in loco vulpiumet operuisti nos umbra mortis.
PS|44|21|Si obliti fuerimus nomen Dei nostriet si expanderimus manus nostras ad deum alienum,
PS|44|22|nonne Deus requiret ista?Ipse enim novit abscondita cordis.
PS|44|23|Quoniam propter te mortificamur tota die,aestimati sumus sicut oves occisionis.
PS|44|24|Evigila, quare obdormis, Domine?Exsurge et ne repellas in finem.
PS|44|25|Quare faciem tuam avertis,oblivisceris inopiae nostrae et tribulationis nostrae?
PS|44|26|Quoniam humiliata est in pulvere anima nostra,conglutinatus est in terra venter noster.Exsurge, Domine, adiuva noset redime nos propter misericordiam tuam.
PS|45|1|Magistro chori. Secundum " Lilia... ". Filiorum Core.Maskil. Canticum amoris.
PS|45|2|Eructavit cor meum verbum bonum,dico ego opera mea regi.Lingua mea calamus scribae velociter scribentis.
PS|45|3|Speciosus forma es prae filiis hominum,diffusa est gratia in labiis tuis,propterea benedixit te Deus in aeternum.
PS|45|4|Accingere gladio tuo super femur tuum, potentissime,magnificentia tua et ornatu tuo.
PS|45|5|Et ornatu tuo procede, currum ascendepropter veritatem et mansuetudinem et iustitiam.Et doceat te mirabilia dextera tua:
PS|45|6|sagittae tuae acutae populi sub te cadent -in corda inimicorum regis.
PS|45|7|Sedes tua, Deus, in saeculum saeculi;sceptrum aequitatis sceptrum regni tui.
PS|45|8|Dilexisti iustitiam et odisti iniquitatem,propterea unxit te Deus, Deus tuus, oleo laetitiae prae consortibus tuis.
PS|45|9|Myrrha et aloe et casia omnia vestimenta tua;e domibus eburneis chordae delectant te.
PS|45|10|Filiae regum in pretiosis tuis;astitit regina a dextris tuis ornata auro ex Ophir. -
PS|45|11|Audi, filia, et vide et inclina aurem tuamet obliviscere populum tuum et domum patris tui;
PS|45|12|et concupiscet rex speciem tuam.Quoniam ipse est dominus tuus, et adora eum.
PS|45|13|Filia Tyri cum muneribus;vultum tuum deprecabuntur divites plebis.
PS|45|14|Gloriosa nimis filia regis intrinsecus,texturis aureis circumamicta.
PS|45|15|In vestibus variegatis adducetur regi;virgines post eam, proximae eius, afferuntur tibi.
PS|45|16|Afferuntur in laetitia et exsultatione,adducuntur in domum regis.
PS|45|17|Pro patribus tuis erunt tibi filii;constitues eos principes super omnem terram.
PS|45|18|Memor ero nominis tuiin omni generatione et generatione;propterea populi confitebuntur tibi in aeternumet in saeculum saeculi.
PS|46|1|Magistro chori. Filiorum Core. Secundum " Virgines... ". Canticum.
PS|46|2|Deus est nobis refugium et virtus,adiutorium in tribulationibus inventus est nimis.
PS|46|3|Propterea non timebimus, dum turbabitur terra,et transferentur montes in cor maris.
PS|46|4|Fremant et intumescant aquae eius, conturbentur montes in elatione eius.
PS|46|5|Fluminis rivi laetificant civitatem Dei,sancta tabernacula Altissimi.
PS|46|6|Deus in medio eius, non commovebitur;adiuvabit eam Deus mane diluculo.
PS|46|7|Fremuerunt gentes, commota sunt regna;dedit vocem suam, liquefacta est terra.
PS|46|8|Dominus virtutum nobiscum,refugium nobis Deus Iacob.
PS|46|9|Venite et videte opera Domini,quae posuit prodigia super terram.Auferet bella usque ad finem terrae,
PS|46|10|arcum conteret et confringet armaet scuta comburet igne.
PS|46|11|Vacate et videte quoniam ego sum Deus:exaltabor in gentibus et exaltabor in terra.
PS|46|12|Dominus virtutum nobiscum,refugium nobis Deus Iacob.
PS|47|1|Magistro chori. Filiorum Core. PSALMUS.
PS|47|2|Omnes gentes, plaudite manibus,iubilate Deo in voce exsultationis,
PS|47|3|quoniam Dominus Altissimus, terribilis,rex magnus super omnem terram.
PS|47|4|Subiecit populos nobiset gentes sub pedibus nostris.
PS|47|5|Elegit nobis hereditatem nostram,gloriam Iacob, quem dilexit.
PS|47|6|Ascendit Deus in iubilo,et Dominus in voce tubae.
PS|47|7|Psallite Deo, psallite;psallite regi nostro, psallite.
PS|47|8|Quoniam rex omnis terrae Deus,psallite sapienter.
PS|47|9|Regnavit Deus super gentes,Deus sedet super sedem sanctam suam.
PS|47|10|Principes populorum congregati suntcum populo Dei Abraham,quoniam Dei sunt scuta terrae:vehementer elevatus est.
PS|48|1|Canticum. PSALMUS. Filiorum Core.
PS|48|2|Magnus Dominus et laudabilis nimisin civitate Dei nostri.
PS|48|3|Mons sanctus eius collis speciosus,exsultatio universae terrae.Mons Sion, extrema aquilonis,civitas regis magni.
PS|48|4|Deus in domibus eius notusfactus est ut refugium.
PS|48|5|Quoniam ecce reges congregati sunt,convenerunt in unum.
PS|48|6|Ipsi cum viderunt, sic admirati sunt,conturbati sunt, diffugerunt;
PS|48|7|illic tremor apprehendit eos,dolores ut parturientis.
PS|48|8|In spiritu orientisconteres naves Tharsis.
PS|48|9|Sicut audivimus, sic vidimusin civitate Domini virtutum,in civitate Dei nostri;Deus fundavit eam in aeternum.
PS|48|10|Recogitamus, Deus, misericordiam tuamin medio templi tui.
PS|48|11|Secundum nomen tuum, Deus,sic et laus tua in fines terrae;iustitia plena est dextera tua.
PS|48|12|Laetetur mons Sion, et exsultent filiae Iudaepropter iudicia tua.
PS|48|13|Circumdate Sion et complectimini eam,numerate turres eius.
PS|48|14|Ponite corda vestra in virtute eiuset percurrite domos eius,ut enarretis in progenie altera.
PS|48|15|Quoniam hic est Deus, Deus nosterin aeternum et in saeculum saeculi;ipse ducet nos in saecula.
PS|49|1|Magistro chori. Filiorum Core. PSALMUS.
PS|49|2|Audite haec, omnes gentes;auribus percipite, omnes, qui habitatis orbem:
PS|49|3|quique humiles et viri nobiles,simul in unum dives et pauper!
PS|49|4|Os meum loquetur sapientiam,et meditatio cordis mei prudentiam.
PS|49|5|Inclinabo in parabolam aurem meam,aperiam in psalterio aenigma meum.
PS|49|6|Cur timebo in diebus malis,cum iniquitas supplantantium circumdabit me?
PS|49|7|Qui confidunt in virtute suaet in multitudine divitiarum suarum gloriantur.
PS|49|8|Etenim seipsum non redimet homo;non dabit Deo propitiationem suam.
PS|49|9|Nimium est pretium redemptionis animae eius:ad ultimum deficiet,
PS|49|10|ut vivat usque in finem nec videat interitum.
PS|49|11|Et videbit sapientes morientes;simul insipiens et stultus peribuntet relinquent alienis divitias suas.
PS|49|12|Sepulcra eorum domus illorum in aeternum;tabernacula eorum in progeniem et progeniem,etsi vocaverunt nominibus suis terras suas.
PS|49|13|Et homo, cum sit in honore, non permanebit;comparatus est iumentis, quae pereunt,et similis factus est illis.
PS|49|14|Haec via illorum, quorum fiducia in semetipsis,et finis eorum, qui complacent in ore suo.
PS|49|15|Sicut oves in inferno positi sunt,mors depascet eos;descendent praecipites ad sepulcrum,et figura eorum erit in consumptionem:infernus habitaculum eorum.
PS|49|16|Verumtamen Deus redimet animam meam,de manu inferi vere suscipiet me.
PS|49|17|Ne timueris, cum dives factus fuerit homo,et cum multiplicata fuerit gloria domus eius,
PS|49|18|quoniam, cum interierit, non sumet omnia,neque descendet cum eo gloria eius.
PS|49|19|Cum animae suae in vita ipsius benedixerit: Laudabunt te quod benefecisti tibi ",
PS|49|20|tamen introibit ad progeniem patrum suorum,qui in aeternum non videbunt lumen.
PS|49|21|Homo, cum in honore esset, non intellexit;comparatus est iumentis, quae pereunt,et similis factus est illis.
PS|50|1|PSALMUS. Asaph.Deus deorum, Dominus, locutus estet vocavit terram a solis ortu usque ad occasum.
PS|50|2|Ex Sion speciosa decore Deus illuxit,
PS|50|3|Deus noster veniet et non silebit:ignis consumens est in conspectu eius,et in circuitu eius tempestas valida.
PS|50|4|Advocabit caelum desursumet terram discernere populum suum:
PS|50|5|" Congregate mihi sanctos meos,qui disposuerunt testamentum meum in sacrificio ".
PS|50|6|Et annuntiabunt caeli iustitiam eius,quoniam Deus iudex est.
PS|50|7|" Audi, populus meus, et loquar,Israel, et testificabor adversum te:Deus, Deus tuus, ego sum.
PS|50|8|Non in sacrificiis tuis arguam te;holocausta enim tua in conspectu meo sunt semper.
PS|50|9|Non accipiam de domo tua vitulosneque de gregibus tuis hircos.
PS|50|10|Quoniam meae sunt omnes ferae silvarum,iumentorum mille in montibus.
PS|50|11|Cognovi omnia volatilia caeli;et, quod movetur in agro, meum est.
PS|50|12|Si esuriero non dicam tibi;meus est enim orbis terrae et plenitudo eius.
PS|50|13|Numquid manducabo carnes taurorumaut sanguinem hircorum potabo?
PS|50|14|Immola Deo sacrificium laudiset redde Altissimo vota tua;
PS|50|15|et invoca me in die tribulationis:eruam te, et honorificabis me ".
PS|50|16|Peccatori autem dixit Deus: Quare tu enarras praecepta meaet assumis testamentum meum in os tuum?
PS|50|17|Tu vero odisti disciplinamet proiecisti sermones meos retrorsum.
PS|50|18|Si videbas furem, currebas cum eo;et cum adulteris erat portio tua.
PS|50|19|Os tuum dimittebas ad malitiam,et lingua tua concinnabat dolos.
PS|50|20|Sedens adversus fratrem tuum loquebariset adversus filium matris tuae proferebas opprobrium.
PS|50|21|Haec fecisti, et tacui.Existimasti quod eram tui similis.Arguam te et statuam illa contra faciem tuam.
PS|50|22|Intellegite haec, qui obliviscimini Deum,ne quando rapiam, et non sit qui eripiat.
PS|50|23|Qui immolabit sacrificium laudis, honorificabit me;et, qui immaculatus est in via, ostendam illi salutare Dei ".
PS|51|1|Magistro chori. PSALMUS. David,
PS|51|2|cum venit ad eum Nathan propheta,postquam cum Bethsabee peccavit.
PS|51|3|Miserere mei, Deus, secundum misericordiam tuam;et secundum multitudinem miserationum tuarumdele iniquitatem meam.
PS|51|4|Amplius lava me ab iniquitate meaet a peccato meo munda me.
PS|51|5|Quoniam iniquitatem meam ego cognosco,et peccatum meum contra me est semper.
PS|51|6|Tibi, tibi soli peccavi et malum coram te feci,ut iustus inveniaris in sententia tua et aequus in iudicio tuo.
PS|51|7|Ecce enim in iniquitate generatus sum,et in peccato concepit me mater mea.
PS|51|8|Ecce enim veritatem in corde dilexistiet in occulto sapientiam manifestasti mihi.
PS|51|9|Asperges me hyssopo, et mundabor;lavabis me, et super nivem dealbabor.
PS|51|10|Audire me facies gaudium et laetitiam,et exsultabunt ossa, quae contrivisti.
PS|51|11|Averte faciem tuam a peccatis meiset omnes iniquitates meas dele.
PS|51|12|Cor mundum crea in me, Deus,et spiritum firmum innova in visceribus meis.
PS|51|13|Ne proicias me a facie tuaet spiritum sanctum tuum ne auferas a me.
PS|51|14|Redde mihi laetitiam salutaris tuiet spiritu promptissimo confirma me.
PS|51|15|Docebo iniquos vias tuas,et impii ad te convertentur.
PS|51|16|Libera me de sanguinibus, Deus, Deus salutis meae,et exsultabit lingua mea iustitiam tuam.
PS|51|17|Domine, labia mea aperies,et os meum annuntiabit laudem tuam.
PS|51|18|Non enim sacrificio delectaris;holocaustum, si offeram, non placebit.
PS|51|19|Sacrificium Deo spiritus contribulatus;cor contritum et humiliatum, Deus, non despicies.
PS|51|20|Benigne fac, Domine, in bona voluntate tua Sion,ut aedificentur muri Ierusalem.
PS|51|21|Tunc acceptabis sacrificium iustitiae, oblationes et holocausta;tunc imponent super altare tuum vitulos.
PS|52|1|Magistro chori. Maskil. David,
PS|52|2|postquam Doeg Edomita ad Saul veniteique narravit dicens: David intravit in domum Abimelech ".
PS|52|3|Quid gloriaris in malitia,qui potens es iniquitate?
PS|52|4|Tota die insidias cogitasti;lingua tua sicut novacula acuta, qui facis dolum.
PS|52|5|Dilexisti malitiam super benignitatem,mendacium magis quam loqui aequitatem.
PS|52|6|Dilexisti omnia verba perditionis, lingua dolosa.
PS|52|7|Propterea Deus destruet te in finem;evellet te et emigrabit te de tabernaculoet radicem tuam de terra viventium.
PS|52|8|Videbunt iusti et timebuntet super eum ridebunt:
PS|52|9|" Ecce homo, qui non posuit Deum refugium suum,sed speravit in multitudine divitiarum suarumet praevaluit in insidiis suis ".
PS|52|10|Ego autem sicut virens oliva in domo Dei.Speravi in misericordia Deiin aeternum et in saeculum saeculi.
PS|52|11|Confitebor tibi in saeculum, quia fecisti;et exspectabo nomen tuum,quoniam bonum est, in conspectu sanctorum tuorum.
PS|53|1|Magistro chori. Secundum " Mahalat ". Maskil. David.Dixit insipiens in corde suo: " Non est Deus ".
PS|53|2|Corrupti sunt et abominationes operati sunt;non est qui faciat bonum.
PS|53|3|Deus de caelo prospexit super filios hominum,ut videat si est intellegens, aut requirens Deum.
PS|53|4|Omnes declinaverunt, simul corrupti sunt;non est qui faciat bonum, non est usque ad unum.
PS|53|5|Nonne scient omnes, qui operantur iniquitatem,qui devorant plebem meam ut cibum panis?Deum non invocaverunt;
PS|53|6|illic trepidaverunt timore, et non erat timor.Quoniam Deus dissipavit ossa eorum, qui te obsidebant,confusi sunt, quoniam Deus sprevit eos. -
PS|53|7|Quis dabit ex Sion salutare Israel?Cum converterit Deus captivitatem plebis suae,exsultabit Iacob, et laetabitur Israel.
PS|54|1|Magistro chori. Fidibus. Maskil. David,
PS|54|2|postquam Ziphaei ad Saul venerunt dicentes: Ecce David apud nos abditus latet ".
PS|54|3|Deus, in nomine tuo salvum me facet in virtute tua iudica me.
PS|54|4|Deus, exaudi orationem meam,auribus percipe verba oris mei!
PS|54|5|Quoniam superbi insurrexerunt adversum me,et fortes quaesierunt animam meamet non proposuerunt Deum ante conspectum suum.
PS|54|6|Ecce enim Deus adiuvat me,et Dominus susceptor est animae meae.
PS|54|7|Converte mala super inimicos meos et in veritate tua disperde illos.
PS|54|8|Voluntarie sacrificabo tibi,confitebor nomini tuo, Domine, quoniam bonum est;
PS|54|9|quoniam ex omni tribulatione eripuit me,et super inimicos meos despexit oculus meus.
PS|55|1|Magistro chori. Fidibus. Maskil. David.
PS|55|2|Auribus percipe, Deus, orationem meamet ne abscondaris a deprecatione mea;
PS|55|3|intende mihi et exaudi me.Excussus sum in meditatione mea et conturbatus sum
PS|55|4|a voce inimici et a tribulatione peccatoris.Quoniam devolverunt in me iniquitatemet in ira molesti erant mihi.
PS|55|5|Cor meum torquetur intra me,et formido mortis cecidit super me.
PS|55|6|Timor et tremor venerunt super me, et contexit me pavor. -
PS|55|7|Et dixi: " Quis dabit mihi pennas sicut columbae,et volabo et requiescam?
PS|55|8|Ecce elongabo fugienset manebo in solitudine.
PS|55|9|Exspectabo eum, qui salvum me faciata spiritu procellae et tempestate ".
PS|55|10|Dissipa, Domine, divide linguas eorum,quoniam vidi violentiam et contentionem in civitate.
PS|55|11|Die ac nocte circumeunt eam super muros eius,
PS|55|12|iniquitas et labor et insidiae in medio eius;et non defecit de plateis eius fraudulentia et dolus.
PS|55|13|Quoniam si inimicus meus maledixisset mihi,sustinuissem utique;et si is qui oderat me, super me magnificatus fuisset,abscondissem me forsitan ab eo.
PS|55|14|Tu vero, homo coaequalis meus,familiaris meus et notus meus,
PS|55|15|qui simul habuimus dulce consortium:in domo Dei ambulavimus in concursu.
PS|55|16|Veniat mors super illos,et descendant in infernum viventes,quoniam nequitiae in habitaculis eorum,in medio eorum.
PS|55|17|Ego autem ad Deum clamabo,et Dominus salvabit me.
PS|55|18|Vespere et mane et meridie meditabor et ingemiscam,et exaudiet vocem meam.
PS|55|19|Redimet in pace animam meam ab his, qui impugnant me,quoniam in multis sunt adversum me.
PS|55|20|Exaudiet Deus et humiliabit illos,qui est ante saecula.Non enim est illis commutatio,et non timuerunt Deum.
PS|55|21|Extendit manum suam in socios;contaminavit foedus suum.
PS|55|22|Lene super butyrum est os eius,pugna autem cor illius:molliti sunt sermones eius super oleum,et ipsi sunt gladii destricti. -
PS|55|23|Iacta super Dominum curam tuam,et ipse te enutriet;non dabit in aeternum fluctuationem iusto.
PS|55|24|Tu vero, Deus, deduces eos in puteum interitus.Viri sanguinum et dolosi non dimidiabunt dies suos;ego autem sperabo in te, Domine.
PS|56|1|Magistro chori. Secundum " Ionat elem rehoqim ".David. Miktam. Cum Gath Philistaei eum tenerent.
PS|56|2|Miserere mei, Deus, quoniam conculcavit me homo,tota die impugnans oppressit me.
PS|56|3|Conculcaverunt me inimici mei tota die,quoniam multi pugnant adversum me, Altissime.
PS|56|4|In quacumque die timebo,ego in te sperabo.
PS|56|5|In Deo, cuius laudabo sermonem,in Deo speravi;non timebo: quid faciet mihi caro?
PS|56|6|Tota die rem meam perturbabant,adversum me omnes cogitationes eorum in malum.
PS|56|7|Concitabant iurgia, insidiabantur,ipsi calcaneum meum observabant.Sicut quaesierunt animam meam,
PS|56|8|ita pro iniquitate retribue illis,in ira populos prosterne, Deus.
PS|56|9|Peregrinationes meas tu numerasti:pone lacrimas meas in utre tuo;nonne in supputatione tua?
PS|56|10|Tunc convertentur inimici mei retrorsum,in quacumque die invocavero:ecce cognovi quoniam Deus meus es.
PS|56|11|In Deo, cuius laudabo sermonem,in Domino, cuius laudabo sermonem,
PS|56|12|in Deo speravi;non timebo: quid faciet mihi homo?
PS|56|13|Super me sunt, Deus, vota tua;reddam laudationes tibi,
PS|56|14|quoniam eripuisti animam meam de morteet pedes meos de lapsu,ut ambulem coram Deo in lumine viventium.
PS|57|1|Magistro chori. Secundum " Ne destruxeris ". David.Miktam. Quando a Saul in cavernam fugit.
PS|57|2|Miserere mei, Deus, miserere mei,quoniam in te confugit anima mea;et in umbra alarum tuarum confugiam,donec transeant insidiae.
PS|57|3|Clamabo ad Deum Altissimum,Deum, qui benefecit mihi.
PS|57|4|Mittet de caelo et liberabit me;dabit in opprobrium conculcantes me.Mittet Deus misericordiam suam et veritatem suam.
PS|57|5|Anima mea recumbit in medio catulorum leonumdevorantium filios hominum.Dentes eorum arma et sagittae,et lingua eorum gladius acutus.
PS|57|6|Exaltare super caelos, Deus,super omnem terram gloria tua.
PS|57|7|Laqueum paraverunt pedibus meis,et incurvavit se anima mea;foderunt ante faciem meam foveam,et ipsi inciderunt in eam.
PS|57|8|Paratum cor meum, Deus,paratum cor meum;
PS|57|9|cantabo et psalmum dicam.Exsurge, gloria mea;exsurge, psalterium et cithara,excitabo auroram.
PS|57|10|Confitebor tibi in populis, Domine,et psalmum dicam tibi in nationibus,
PS|57|11|quoniam magnificata est usque ad caelos misericordia tua,et usque ad nubes veritas tua.
PS|57|12|Exaltare super caelos, Deus,super omnem terram gloria tua.
PS|58|1|Magistro chori. Secundum " Ne destruxeris ".David. Miktam.
PS|58|2|Numquid vere, potentes, iustitiam loquimini,recte iudicatis filios hominum?
PS|58|3|Etenim in corde iniquitates operamini,in terra violentiam manus vestrae concinnant.
PS|58|4|Alienati sunt peccatores ab utero;erraverunt a ventre, qui loquuntur falsa.
PS|58|5|Venenum illis in similitudinem serpentis,sicut aspidis surdae et obturantis aures suas,
PS|58|6|quae non exaudiet vocem incantantiumet venefici incantantis sapienter.
PS|58|7|Deus, contere dentes eorum in ore ipsorum;molas leonum confringe, Domine.
PS|58|8|Diffluant tamquam aqua decurrens,sicut fenum conculcatum arescant.
PS|58|9|Sicut limax, quae tabescens transit, sicut abortivum mulieris, quod non vidit solem.
PS|58|10|Priusquam sentiant ollae vestrae rhamnum,sicut viventes, sicut ardor irae absorbet eos.
PS|58|11|Laetabitur iustus, cum viderit vindictam,pedes suos lavabit in sanguine peccatoris.
PS|58|12|Et dicet homo: " Utique est fructus iusto,utique est Deus iudicans eos in terra ".
PS|59|1|Magistro chori. Secundum " Ne destruxeris ".David. Miktam. Quando Saul viros misit,qui domum observarent et eum occiderent.
PS|59|2|Eripe me de inimicis meis, Deus meus,et ab insurgentibus in me protege me.
PS|59|3|Eripe me de operantibus iniquitatemet de viris sanguinum salva me.
PS|59|4|Quia ecce insidiati sunt animae meae,irruerunt in me fortes.
PS|59|5|Neque delictum neque peccatum in me est, Domine;sine iniquitate mea currunt et praeparantur.Exsurge in occursum meum et vide;
PS|59|6|et tu, Domine, Deus virtutum, Deus Israel,evigila ad visitandas omnes gentes; non miserearis omnibus, qui infideliter operantur.
PS|59|7|Revertentur ad vesperam et latrabunt ut caneset circuibunt civitatem.
PS|59|8|Ecce eructabunt ore suo,et gladius in labiis eorum: " Quis enim audit? ".
PS|59|9|Et tu, Domine, deridebis eos,subsannabis omnes gentes.
PS|59|10|Fortitudo mea, tibi attendam,quia, Deus, praesidium meum es.
PS|59|11|Deus meus, misericordia eius praeveniet me.Deus faciet, ut despiciam inimicos meos.
PS|59|12|Ne occidas eos, ne quando obliviscatur populus meus;disperge illos in virtute tuaet prosterne eos, protector meus, Domine.
PS|59|13|Peccatum oris eorum, sermo labiorum ipsorum,et comprehendantur in superbia sua.Propter exsecrationem et mendacium, quod loquuntur,
PS|59|14|consume eos in furore,consume, et non erunt;et scient quia Deus dominabitur Iacob et finium terrae.
PS|59|15|Revertentur ad vesperam et latrabunt ut caneset circuibunt civitatem.
PS|59|16|Ipsi errabunt ad manducandum;si vero non fuerint saturati, murmurabunt.
PS|59|17|Ego autem cantabo fortitudinem tuamet exsultabo mane misericordiam tuam,quia factus es praesidium meumet refugium meum in die tribulationis meae.
PS|59|18|Fortitudo mea, tibi psallam,quia, Deus, praesidium meum es:Deus meus misericordia mea.
PS|60|1|Magistro chori. Secundum " Lilium praecepti ".Miktam. David. Ad docendum.
PS|60|2|Quando contra Aram Naharaim et Aram Soba egressus est,et quando Ioab reversus devicit Edom in valle Salis:duodecim milia (hominum).
PS|60|3|Deus, reppulisti nos, destruxisti nos.Iratus es. Convertere ad nos!
PS|60|4|Concussisti terram, confregisti eam;sana contritiones eius, quia commota est.
PS|60|5|Ostendisti populo tuo dura,potasti nos vino vertiginis.
PS|60|6|Dedisti metuentibus te signum,ut fugiant a facie arcus.
PS|60|7|Ut liberentur dilecti tui,salvos fac dextera tua et exaudi nos.
PS|60|8|Deus locutus est in sancto suo: Laetabor et partibor Sichimamet convallem Succoth metibor.
PS|60|9|Meus est Galaad, et meus est Manasses,et Ephraim fortitudo capitis mei.Iuda sceptrum meum,
PS|60|10|Moab olla lavacri mei.Super Idumaeam extendam calceamentum meum,super Philistaeam vociferabor ".
PS|60|11|Quis adducet me in civitatem munitam?Quis deducet me usque in Idumaeam?
PS|60|12|Nonne tu, Deus, qui reppulisti nos;et non egredieris, Deus, in virtutibus nostris?Da nobis auxilium de tribulatione, quia vana salus hominis.
PS|60|13|In Deo faciemus virtutem,et ipse conculcabit tribulantes nos.
PS|61|1|Magistro chori. Fidibus. David.
PS|61|2|Exaudi, Deus, deprecationem meam,intende orationi meae.
PS|61|3|A finibus terrae ad te clamavi,dum anxiaretur cor meum.In petram inaccessam mihi deduc me!
PS|61|4|Quia factus es spes mea,turris fortitudinis a facie inimici.
PS|61|5|Inhabitabo in tabernaculo tuo in saecula,protegar in velamento alarum tuarum,
PS|61|6|quoniam tu, Deus meus, exaudisti vota mea,dedisti hereditatem timentium nomen tuum.
PS|61|7|Dies super dies regis adicies,annos eius usque in diem generationis et generationis.
PS|61|8|Sedeat in aeternum in conspectu Dei;misericordia et veritas servent eum.
PS|61|9|Sic psalmum dicam nomini tuo in saeculum saeculi,ut reddam vota mea de die in diem.
PS|62|1|Magistro chori. Secundum Iduthun. PSALMUS. David.
PS|62|2|In Deo tantum quiesce, anima mea,ab ipso enim salutare meum.
PS|62|3|Verumtamen ipse refugium meum et salutare meum,praesidium meum; non movebor amplius.
PS|62|4|Quousque irruitis in hominem, contunditis universi vostamquam parietem inclinatum et maceriam depulsam?
PS|62|5|Verumtamen de excelso suo cogitaverunt depellere;delectabantur mendacio.Ore suo benedicebant et corde suo maledicebant.
PS|62|6|In Deo tantum quiesce, anima mea, quoniam ab ipso patientia mea.
PS|62|7|Verumtamen ipse Deus meus et salutare meum,praesidium meum; non movebor.
PS|62|8|In Deo salutare meum et gloria mea; Deus fortitudinis meae, et refugium meum in Deo est.
PS|62|9|Sperate in eo, omnis congregatio populi,effundite coram illo corda vestra;Deus refugium nobis.
PS|62|10|Verumtamen vanitas filii Adam,mendacium filii hominum.In stateram si conscendant,super fumum leves sunt omnes.
PS|62|11|Nolite sperare in violentiaet in rapina nolite decipi;divitiae si affluant, nolite cor apponere.
PS|62|12|Semel locutus est Deus,duo haec audivi:quia potestas Deo est,
PS|62|13|et tibi, Domine, misericordia;quia tu reddes unicuique iuxta opera sua.
PS|63|1|PSALMUS. David, cum in deserto Iudae commoraretur.
PS|63|2|Deus, Deus meus es tu, ad te de luce vigilo.Sitivit in te anima mea,te desideravit caro mea.In terra deserta et arida et inaquosa,
PS|63|3|sic in sancto apparui tibi,ut viderem virtutem tuam et gloriam tuam.
PS|63|4|Quoniam melior est misericordia tua super vitas,labia mea laudabunt te.
PS|63|5|Sic benedicam te in vita meaet in nomine tuo levabo manus meas.
PS|63|6|Sicut adipe et pinguedine repleatur anima mea,et labiis exsultationis laudabit os meum.
PS|63|7|Cum memor ero tui super stratum meum,in matutinis meditabor de te,
PS|63|8|quia fuisti adiutor meus,et in velamento alarum tuarum exsultabo.
PS|63|9|Adhaesit anima mea post te,me suscepit dextera tua.
PS|63|10|Ipsi vero in ruinam quaesierunt animam meam,introibunt in inferiora terrae,
PS|63|11|tradentur in potestatem gladii,partes vulpium erunt.
PS|63|12|Rex vero laetabitur in Deo;gloriabuntur omnes, qui iurant in eo,quia obstructum est os loquentium iniqua.
PS|64|1|Magistro chori. PSALMUS. David.
PS|64|2|Exaudi, Deus, vocem meam in meditatione mea;a timore inimici custodi animam meam.
PS|64|3|Protege me a conventu malignantium,a multitudine operantium iniquitatem.
PS|64|4|Qui exacuerunt ut gladium linguas suas,intenderunt sagittas suas, venefica verba,
PS|64|5|ut sagittent in occultis immaculatum.Subito sagittabunt eum et non timebunt,
PS|64|6|firmaverunt sibi consilium nequam.Disputaverunt, ut absconderent laqueos,dixerunt: " Quis videbit eos? ".
PS|64|7|Excogitaverunt iniqua, perfecerunt excogitata consilia.Interiora hominis et cor eius abyssus.
PS|64|8|Et sagittavit illos Deus;subito factae sunt plagae eorum,
PS|64|9|et infirmavit eos lingua eorum.Caput movebunt omnes, qui videbunt eos,
PS|64|10|et timebit omnis homo;et annuntiabunt opera Deiet facta eius intellegent.
PS|64|11|Laetabitur iustus in Domino et sperabit in eo,et gloriabuntur omnes recti corde.
PS|65|1|Magistro chori. PSALMUS. David. Canticum.
PS|65|2|Te decet hymnus, Deus, in Sion;et tibi reddetur votum in Ierusalem.
PS|65|3|Qui audis orationem,ad te omnis caro veniet propter iniquitatem.
PS|65|4|Etsi praevaluerunt super nos impietates nostrae,tu propitiaberis eis.
PS|65|5|Beatus, quem elegisti et assumpsisti; inhabitabit in atriis tuis.Replebimur bonis domus tuae,sanctitate templi tui.
PS|65|6|Mirabiliter in aequitateexaudies nos, Deus salutis nostrae,spes omnium finium terrae et maris longinqui.
PS|65|7|Firmans montes in virtute tua,accinctus potentia.
PS|65|8|Compescens sonitum maris,sonitum fluctuum eiuset tumultum populorum.
PS|65|9|Et timebunt, qui habitant terminos terrae, a signis tuis;exitus orientis et occidentis delectabis.
PS|65|10|Visitasti terram et inebriasti eam;multiplicasti locupletare eam.Flumen Dei repletum est aquis;parasti frumenta illorum,quoniam ita parasti eam.
PS|65|11|Sulcos eius irrigans, glebas eius complanans;imbribus emollis eam, benedicis germini eius.
PS|65|12|Coronasti annum benignitate tua,et vestigia tua stillabunt pinguedinem.
PS|65|13|Stillabunt pascua deserti,et exsultatione colles accingentur.
PS|65|14|Induta sunt ovibus prata,et valles abundabunt frumento;clamabunt, etenim hymnum dicent.
PS|66|1|Magistro chori. Canticum. PSALMUS.Iubilate Deo, omnis terra,
PS|66|2|psalmum dicite gloriae nominis eius,glorificate laudem eius.
PS|66|3|Dicite Deo: " Quam terribilia sunt opera tua.Prae multitudine virtutis tuae blandientur tibi inimici tui.
PS|66|4|Omnis terra adoret te et psallat tibi,psalmum dicat nomini tuo ".
PS|66|5|Venite et videte opera Dei,terribilis in adinventionibus super filios hominum.
PS|66|6|Convertit mare in aridam,et in flumine pertransibunt pede;ibi laetabimur in ipso.
PS|66|7|Qui dominatur in virtute sua in aeternum,oculi eius super gentes respiciunt;rebelles non exaltentur in semetipsis.
PS|66|8|Benedicite, gentes, Deum nostrumet auditam facite vocem laudis eius;
PS|66|9|qui posuit animam nostram ad vitamet non dedit in commotionem pedes nostros.
PS|66|10|Quoniam probasti nos, Deus;igne nos examinasti, sicut examinatur argentum.
PS|66|11|Induxisti nos in laqueum,posuisti tribulationes in dorso nostro.
PS|66|12|Imposuisti homines super capita nostra,transivimus per ignem et aquam,et eduxisti nos in refrigerium.
PS|66|13|Introibo in domum tuam in holocaustis;reddam tibi vota mea,
PS|66|14|quae protulerunt labia mea,et locutum est os meum in tribulatione mea.
PS|66|15|Holocausta medullata offeram tibi cum incenso arietum,offeram tibi boves cum hircis.
PS|66|16|Venite, audite, et narrabo, omnes, qui timetis Deum,quanta fecit animae meae.
PS|66|17|Ad ipsum ore meo clamaviet exaltavi in lingua mea.
PS|66|18|Iniquitatem si aspexi in corde meo,non exaudiet Dominus.
PS|66|19|Propterea exaudivit Deus,attendit voci deprecationis meae.
PS|66|20|Benedictus Deus, qui non amovit orationem meamet misericordiam suam a me.
PS|67|1|Magistro chori. Fidibus. PSALMUS. Canticum.
PS|67|2|Deus misereatur nostri et benedicat nobis;illuminet vultum suum super nos,
PS|67|3|ut cognoscatur in terra via tua,in omnibus gentibus salutare tuum.
PS|67|4|Confiteantur tibi populi, Deus;confiteantur tibi populi omnes.
PS|67|5|Laetentur et exsultent gentes,quoniam iudicas populos in aequitateet gentes in terra dirigis.
PS|67|6|Confiteantur tibi populi, Deus;confiteantur tibi populi omnes.
PS|67|7|Terra dedit fructum suum;benedicat nos Deus, Deus noster,
PS|67|8|benedicat nos Deus,et metuant eum omnes fines terrae.
PS|68|1|Magistro chori. David. PSALMUS. Canticum.
PS|68|2|Exsurgit Deus, et dissipantur inimici eius;et fugiunt, qui oderunt eum, a facie eius.
PS|68|3|Sicut dissipatur fumus, tu dissipas;sicut fluit cera a facie ignis,sic pereunt peccatores a facie Dei.
PS|68|4|Et iusti laetentur et exsultent in conspectu Deiet delectentur in laetitia.
PS|68|5|Cantate Deo, psalmum dicite nomini eius;iter facite ei, qui fertur super nubes:Dominus nomen illi.Iubilate in conspectu eius;
PS|68|6|pater orphanorum et iudex viduarum,Deus in habitaculo sancto suo.
PS|68|7|Deus, qui inhabitare facit desolatos in domo,qui educit vinctos in prosperitatem;verumtamen rebelles habitabunt in arida terra. -
PS|68|8|Deus, cum egredereris in conspectu populi tui,cum pertransires in deserto,
PS|68|9|terra mota est, etiam caeli distillaverunta facie Dei Sinai, a facie Dei Israel.
PS|68|10|Pluviam voluntariam effundebas, Deus;hereditatem tuam infirmatam, tu refecisti eam.
PS|68|11|Animalia tua habitabant in ea,parasti in bonitate tua pauperi, Deus.
PS|68|12|Dominus dat verbum;virgines annuntiantes bona sunt agmen ingens:
PS|68|13|" Reges exercituum fugiunt, fugiunt,et species domus dividit spolia.
PS|68|14|Et vos dormitis inter medias caulas:alae columbae nitent argento,et pennae eius pallore auri.
PS|68|15|Dum dispergit Omnipotens reges super eam,nive dealbatur Selmon ".
PS|68|16|Mons Dei mons Basan,mons cacuminum mons Basan.
PS|68|17|Ut quid invidetis, montes cacuminum,monti, in quo beneplacitum est Deo inhabitare?Etenim Dominus habitabit in finem.
PS|68|18|Currus Dei decem milia milium:Dominus venit de Sinai in sancta.
PS|68|19|Ascendisti in altum, captivam duxisti captivitatem;accepisti in donum homines,ut etiam rebelles habitent apud Dominum Deum.
PS|68|20|Benedictus Dominus die cotidie;portabit nos Deus salutarium nostrorum.
PS|68|21|Deus noster, Deus ad salvandum;et Domini, Domini exitus mortis.
PS|68|22|Verumtamen Deus confringet capita inimicorum suorum,verticem capillatum perambulantium in delictis suis.
PS|68|23|Dixit Dominus: " Ex Basan reducam,reducam de profundo maris,
PS|68|24|ut intingatur pes tuus in sanguine,lingua canum tuorum ex inimicis portionem inveniat ".
PS|68|25|Viderunt ingressus tuos, Deus,ingressus Dei mei, regis mei in sancta.
PS|68|26|Praecedunt cantores, postremi veniunt psallentes.in medio iuvenculae tympanistriae.
PS|68|27|" In ecclesiis benedicite Deo,Domino, vos de fontibus Israel ".
PS|68|28|Ibi Beniamin adulescentulus ducens eos,principes Iudae cum turma sua,principes Zabulon, principesNephthali.
PS|68|29|Manda, Deus, virtuti tuae;confirma hoc, Deus, quod operatus es in nobis.
PS|68|30|A templo tuo in Ierusalemtibi afferent reges munera.
PS|68|31|Increpa feram arundinis,congregationem taurorum in vitulis populorum:prosternant se cum laminis argenti.Dissipa gentes, quae bella volunt.
PS|68|32|Venient optimates ex Aegypto,Aethiopia praeveniet manus suas Deo.
PS|68|33|Regna terrae, cantate Deo,psallite Domino, psallite Deo,
PS|68|34|qui fertur super caelum caeli ad orientem;ecce dabit vocem suam, vocem virtutis.
PS|68|35|Tribuite virtutem Deo.Super Israel magnificentia eius,et virtus eius in nubibus.
PS|68|36|Mirabilis, Deus, de sanctuario tuo!Deus Israel ipse tribuet virtutem et fortitudinem plebi suae.Benedictus Deus!
PS|69|1|Magistro chori. Secundum " Lilia... ". David.
PS|69|2|Salvum me fac, Deus,quoniam venerunt aquae usque ad guttur meum.
PS|69|3|Infixus sum in limo profundi, et non est substantia;veni in profunda aquarum, et fluctus demersit me.
PS|69|4|Laboravi clamans, raucae factae sunt fauces meae;defecerunt oculi mei, dum spero in Deum meum.
PS|69|5|Multiplicati sunt super capillos capitis mei,qui oderunt me gratis.Confortati sunt, qui persecuti sunt me inimici mei mendaces;quae non rapui, tunc exsolvebam.
PS|69|6|Deus, tu scis insipientiam meam,et delicta mea a te non sunt abscondita.
PS|69|7|Non erubescant in me, qui exspectant te,Domine, Domine virtutum.Non confundantur super me,qui quaerunt te, Deus Israel.
PS|69|8|Quoniam propter te sustinui opprobrium,operuit confusio faciem meam;
PS|69|9|extraneus factus sum fratribus meiset peregrinus filiis matris meae.
PS|69|10|Quoniam zelus domus tuae comedit me,et opprobria exprobrantium tibi ceciderunt super me.
PS|69|11|Et flevi in ieiunio animam meam,et factum est in opprobrium mihi.
PS|69|12|Et posui vestimentum meum cilicium,et factus sum illis in parabolam.
PS|69|13|Adversum me loquebantur, qui sedebant in porta,et in me canebant, qui bibebant vinum.
PS|69|14|Ego vero orationem meam ad te, Domine,in tempore beneplaciti, Deus.In multitudine misericordiae tuae exaudi me,in veritate salutis tuae.
PS|69|15|Eripe me de luto, ut non infigar,eripiar ab iis, qui oderunt me,et de profundis aquarum.
PS|69|16|Non me demergat fluctus aquarum,neque absorbeat me profundum,neque urgeat super me puteus os suum.
PS|69|17|Exaudi me, Domine, quoniam benigna est misericordia tua;secundum multitudinem miserationum tuarum respice in me.
PS|69|18|Et ne avertas faciem tuam a puero tuo;quoniam tribulor, velociter exaudi me.
PS|69|19|Accede ad animam meam, vindica eam,propter inimicos meos redime me.
PS|69|20|Tu scis opprobrium meumet confusionem meam et reverentiam meam. -In conspectu tuo sunt omnes, qui tribulant me;
PS|69|21|opprobrium contrivit cor meum, et elangui.Et sustinui, qui simul contristaretur, et non fuit,et qui consolaretur, et non inveni.
PS|69|22|Et dederunt in escam meam felet in siti mea potaverunt me aceto.
PS|69|23|Fiat mensa eorum coram ipsis in laqueumet in retributiones et in scandalum.
PS|69|24|Obscurentur oculi eorum, ne videant,et lumbos eorum semper infirma.
PS|69|25|Effunde super eos iram tuam,et furor irae tuae comprehendat eos.
PS|69|26|Fiat commoratio eorum deserta,et in tabernaculis eorum non sit qui inhabitet.
PS|69|27|Quoniam, quem tu percussisti, persecuti sunt,et super dolorem eius, quem vulnerasti, addiderunt.
PS|69|28|Appone iniquitatem super iniquitatem eorum,et non veniant ad iustitiam tuam.
PS|69|29|Deleantur de libro viventiumet cum iustis non scribantur.
PS|69|30|Ego autem sum pauper et dolens;salus tua, Deus, suscipit me.
PS|69|31|Laudabo nomen Dei cum canticoet magnificabo eum in laude.
PS|69|32|Et placebit Domino super taurum,super vitulum cornua producentem et ungulas.
PS|69|33|Videant humiles et laetentur;quaerite Deum, et vivet cor vestrum,
PS|69|34|quoniam exaudivit pauperes Dominuset vinctos suos non despexit.
PS|69|35|Laudent illum caeli et terra,maria et omnia reptilia in eis.
PS|69|36|Quoniam Deus salvam faciet Sionet aedificabit civitates Iudae;et inhabitabunt ibi et possidebunt eam.
PS|69|37|Et semen servorum eius hereditabunt eam;et, qui diligunt nomen eius, habitabunt in ea.
PS|70|1|Magistro chori. David. Ad commemorandum.
PS|70|2|Deus, in adiutorium meum intende;Domine, ad adiuvandum me festina.
PS|70|3|Confundantur et revereantur,qui quaerunt animam meam.Avertantur retrorsum et erubescant,qui volunt mihi mala.
PS|70|4|Convertantur propter confusionem suam,qui dicunt mihi: " Euge, euge ".
PS|70|5|Exsultent et laetentur in te omnes, qui quaerunt te;et dicant semper: " Magnificetur Deus ",qui diligunt salutare tuum.
PS|70|6|Ego vero egenus et pauper sum;Deus, ad me festina.Adiutor meus et liberator meus es tu;Domine, ne moreris.
PS|71|1|In te, Domine, speravi,non confundar in aeternum.
PS|71|2|In iustitia tua libera me et eripe me;inclina ad me aurem tuam et salva me.
PS|71|3|Esto mihi in rupem praesidiiet in domum munitam, ut salvum me facias,quoniam fortitudo mea et refugium meum es tu.
PS|71|4|Deus meus, eripe me de manu peccatoriset de manu contra legem agentis et iniqui.
PS|71|5|Quoniam tu es exspectatio mea, Domine;Domine, spes mea a iuventute mea.
PS|71|6|Super te innixus sum ex utero,de ventre matris meae tu es susceptor meus;in te laus mea semper.
PS|71|7|Tamquam prodigium factus sum multis,et tu adiutor fortis. -
PS|71|8|Repleatur os meum laude tua,tota die magnitudine tua.
PS|71|9|Ne proicias me in tempore senectutis;cum defecerit virtus mea, ne derelinquas me.
PS|71|10|Quia dixerunt inimici mei mihi,et, qui observabant animam meam,consilium fecerunt in unum
PS|71|11|dicentes: " Deus dereliquit eum!Persequimini et comprehenditeeum,quia non est qui eripiat ".
PS|71|12|Deus, ne elongeris a me;Deus meus, in auxilium meum festina.
PS|71|13|Confundantur et deficiant adversantes animae meae;operiantur confusione et pudore, qui quaerunt mala mihi.
PS|71|14|Ego autem semper speraboet adiciam super omnem laudem tuam.
PS|71|15|Os meum annuntiabit iustitiam tuam,tota die salutare tuum:quae dinumerare nescivi.
PS|71|16|Veniam ad potentias Domini;Domine, memorabor iustitiae tuae solius.
PS|71|17|Deus, docuisti me a iuventute mea;et usque nunc annuntiabo mirabilia tua.
PS|71|18|Et usque in senectam et senium,Deus, ne derelinquas me,donec annuntiem brachium tuumgenerationi omni, quae ventura est.Potentia tua
PS|71|19|et iustitia tua, Deus,usque in altissima, qui fecisti magnalia:Deus, quis similis tibi?
PS|71|20|Quantas ostendisti mihi tribulationes multas et malas;iterum vivificasti meet de abyssis terrae iterum reduxisti me.
PS|71|21|Multiplicabis magnitudinem meam et conversus consolaberis me.
PS|71|22|Nam et ego confitebor tibiin psalterio veritatem tuam, Deus meus;psallam tibi in cithara, Sanctus Israel.
PS|71|23|Exsultabunt labia mea, cum cantavero tibi,et anima mea, quam redemisti;
PS|71|24|sed et lingua mea tota die meditabitur iustitiam tuam,cum confusi et reveriti fuerint, qui quaerunt mala mihi.
PS|72|1|Salomonis. Deus, iudicium tuum regi daet iustitiam tuam filio regis;
PS|72|2|iudicet populum tuum in iustitiaet pauperes tuos in iudicio.
PS|72|3|Afferant montes pacem populo,et colles iustitiam.
PS|72|4|Iudicabit pauperes populiet salvos faciet filios inopiset humiliabit calumniatorem.
PS|72|5|Et permanebit cum sole et ante lunamin generatione et generationem.
PS|72|6|Descendet sicut pluvia in gramen,et sicut imber irrigans terram.
PS|72|7|Florebit in diebus eius iustitia et abundantia pacis,donec auferatur luna.
PS|72|8|Et dominabitur a mari usque ad mareet a flumine usque ad terminos orbis terrarum.
PS|72|9|Coram illo procident incolae deserti,et inimici eius terram lingent.
PS|72|10|Reges Tharsis et insulae munera offerent,reges Arabum et Saba dona adducent.
PS|72|11|Et adorabunt eum omnes reges, omnes gentes servient ei.
PS|72|12|Quia liberabit inopem clamantemet pauperem, cui non erat adiutor.
PS|72|13|Parcet pauperi et inopiet animas pauperum salvas faciet.
PS|72|14|Ex oppressione et violentia redimet animas eorum,et pretiosus erit sanguis eorum coram illo. -
PS|72|15|Et vivet, et dabitur ei de auro Arabiae, et orabunt pro ipso semper; tota die benedicent ei.
PS|72|16|Et erit ubertas frumenti in terra, in summis montium fluctuabit, sicut Libanus fructus eius;et florebunt de civitate sicut fenum terrae.
PS|72|17|Sit nomen eius benedictum in saecula,ante solem permanebit nomen eius.Et benedicentur in ipso omnes tribus terrae,omnes gentes magnificabunt eum.
PS|72|18|Benedictus Dominus Deus, Deus Israel,qui facit mirabilia solus.
PS|72|19|Et benedictum nomen maiestatis eius in aeternum;et replebitur maiestate eius omnis terra. Fiat, fiat.
PS|73|1|PSALMUS. Asaph.Quam bonus rectis est Deus,Deus his, qui mundo sunt corde!
PS|73|2|Mei autem paene moti sunt pedes,paene effusi sunt gressus mei,
PS|73|3|quia zelavi super gloriantes,pacem peccatorum videns.
PS|73|4|Quia non sunt eis impedimenta,sanus et pinguis est venter eorum.
PS|73|5|In labore mortalium non suntet cum hominibus non flagellantur.
PS|73|6|Ideo quasi torques est eis superbia,et tamquam indumentum operuit eos violentia.
PS|73|7|Prodit quasi ex adipe iniquitas eorum,erumpunt cogitationes cordis.
PS|73|8|Subsannaverunt et locuti sunt nequitiam,iniquitatem ab excelso locuti sunt.
PS|73|9|Posuerunt in caelo os suum,et lingua eorum transivit in terra.
PS|73|10|Ideo in alto sedent,et aquae plenae non pervenient ad eos.
PS|73|11|Et dixerunt: " Quomodo scit Deus,et si est scientia in Excelso? ".
PS|73|12|Ecce ipsi peccatores et abundantes in saeculomultiplicaverunt divitias.
PS|73|13|Et dixi: " Ergo sine causa mundavi cor meumet lavi in innocentia manus meas;
PS|73|14|et fui flagellatus tota die,et castigatio mea in matutinis ".
PS|73|15|Si dixissem: " Loquar ut illi ",ecce generationem filiorum tuorum prodidissem.
PS|73|16|Et cogitabam, ut cognoscerem hoc;labor erat in oculis meis,
PS|73|17|donec intravi in sanctuarium Deiet intellexi novissima eorum.
PS|73|18|Verumtamen in lubrico posuisti eos,deiecisti eos in ruinas.
PS|73|19|Quomodo facti sunt in desolationem!Subito defecerunt, perierunt prae horrore.
PS|73|20|Velut somnium evigilantis, Domine,surgens imaginem ipsorum contemnes.
PS|73|21|Quia exacerbatum est cor meum,et renes mei compuncti sunt;
PS|73|22|et ego insipiens factus sum et nescivi:ut iumentum factus sum apud te.
PS|73|23|Ego autem semper tecum;tenuisti manum dexteram meam.
PS|73|24|In consilio tuo deduces meet postea cum gloria suscipies me.
PS|73|25|Quis enim mihi est in caelo?Et tecum nihil volui super terram.
PS|73|26|Defecit caro mea et cor meum;Deus cordis mei, et pars mea Deus in aeternum.
PS|73|27|Quia ecce, qui elongant se a te, peribunt;perdidisti omnes, qui fornicantur abs te.
PS|73|28|Mihi autem adhaerere Deo bonum est,ponere in Domino Deo spem meam,ut annuntiem omnes operationes tuasin portis filiae Sion.
PS|74|1|Maskil. Asaph.Ut quid, Deus, reppulisti in finem,iratus est furor tuus super oves pascuae tuae?
PS|74|2|Memor esto congregationis tuae,quam possedisti ab initio.Redemisti virgam hereditatis tuae: mons Sion, in quo habitasti.
PS|74|3|Leva gressus tuos in ruinas sempiternas:omnia vastavit inimicus in sancto.
PS|74|4|Rugierunt, qui oderunt te,in medio congregationis tuae;posuerunt signa sua in signa.
PS|74|5|Visi sunt quasi in altum securim vibrantesin silva condensa.
PS|74|6|Exciderunt ianuas eius in idipsum;in securi et ascia deiecerunt.
PS|74|7|Incenderunt igni sanctuarium tuum,in terram polluerunt tabernaculum nominis tui;
PS|74|8|dixerunt in corde suo: " Opprimamus eos simul ".Combusserunt omnes congregationes Dei in terra.
PS|74|9|Signa nostra non vidimus;iam non est propheta,et apud nos non est qui cognoscat amplius.
PS|74|10|Usquequo, Deus, improperabit inimicus,spernet adversarius nomen tuum in finem?
PS|74|11|Ut quid avertis manum tuamet tenes dexteram tuam in medio sinu tuo?
PS|74|12|Deus autem rex noster ante saecula,operatus est salutes in medio terrae.
PS|74|13|Tu conscidisti in virtute tua mare,contribulasti capita draconum in aquis.
PS|74|14|Tu confregisti capita Leviathan,dedisti eum escam monstris maris.
PS|74|15|Tu dirupisti fontes et torrentes;tu siccasti fluvios perennes.
PS|74|16|Tuus est dies, et tua est nox,tu fabricatus es luminaria et solem.
PS|74|17|Tu statuisti omnes terminos terrae,aestatem et hiemem, tu plasmasti ea.
PS|74|18|Memor esto huius:inimicus improperavit Domino,et populus insipiens sprevit nomen tuum.
PS|74|19|Ne tradas bestiis animas confitentes tibiet animas pauperum tuorum ne obliviscaris in finem.
PS|74|20|Respice in testamentum,quia repleta sunt latibula terrae tentoriis violentiae.
PS|74|21|Ne revertatur humilis factus confusus;pauper et inops laudabunt nomen tuum.
PS|74|22|Exsurge, Deus, iudica causam tuam;memor esto improperiorum tuorum,quae ab insipiente fiunt tota die.
PS|74|23|Ne obliviscaris voces inimicorum tuorum;tumultus adversariorum tuorum ascendit semper.
PS|75|1|Magistro chori. Secundum " Ne destruxeris ".PSALMUS. Asaph. Canticum.
PS|75|2|Confitebimur tibi, Deus;confitebimur et invocabimus nomen tuum:narrabimus mirabilia tua.
PS|75|3|Cum statuero tempus,ego iustitias iudicabo.
PS|75|4|Si liquefacta est terra et omnes, qui habitant in ea,ego confirmavi columnas eius.
PS|75|5|Dixi gloriantibus: " Nolite gloriari! "et delinquentibus: "Nolite exaltare cornu!
PS|75|6|Nolite exaltare in altum cornu vestrum;nolite loqui adversus Deum proterva ".
PS|75|7|Quia neque ab oriente neque ab occidenteneque a desertis exaltatio.
PS|75|8|Quoniam Deus iudex est:hunc humiliat et hunc exaltat.
PS|75|9|Quia calix in manu Dominivini meri plenus mixto.Et inclinavit ex hoc in hoc;verumtamen usque ad faeces epotabunt,bibent omnes peccatores terrae.
PS|75|10|Ego autem annuntiabo in saeculum,cantabo Deo Iacob.
PS|75|11|Et omnia cornua peccatorum confringam,et exaltabuntur cornua iusti.
PS|76|1|Magistro chori. Fidibus. PSALMUS. Asaph. Canticum.
PS|76|2|Notus in Iudaea Deus,in Israel magnum nomen eius.
PS|76|3|Et est in Salem tabernaculum eius,et habitatio eius in Sion.
PS|76|4|Ibi confregit coruscationes arcus,scutum, gladium et bellum.
PS|76|5|Illuminans tu, Mirabilis,a montibus direptionis.
PS|76|6|Spoliati sunt potentes corde, dormierunt somnum suum,et non invenerunt omnes viri fortes manus suas.
PS|76|7|Ab increpatione tua, Deus Iacob,dormitaverunt auriga et equus.
PS|76|8|Tu terribilis es, et quis resistet tibi?Ex tunc ira tua.
PS|76|9|De caelo auditum fecisti iudicium;terra tremuit et quievit,
PS|76|10|cum exsurgeret in iudicium Deus,ut salvos faceret omnes mansuetos terrae.
PS|76|11|Quoniam furor hominis confitebitur tibi,et reliquiae furoris diem festum agent tibi.
PS|76|12|Vovete et reddite Domino Deo vestro;omnes in circuitu eius afferant munera Terribili,
PS|76|13|ei, qui aufert spiritum principum,terribili apud reges terrae.
PS|77|1|Magistro chori. Secundum Idithun. Asaph. PSALMUS.
PS|77|2|Voce mea ad Dominum clamavi;voce mea ad Deum, et intendit mihi.
PS|77|3|In die tribulationis meae Deum exquisivi,manus meae nocte expansae suntet non fatigantur.Renuit consolari anima mea;
PS|77|4|memor sum Dei et ingemisco,exerceor, et deficit spiritus meus.
PS|77|5|Vigiles tenuisti palpebras oculi mei; turbatus sum et non sum locutus.
PS|77|6|Cogitavi dies antiquoset annos aeternos in mente habui.
PS|77|7|Meditatus sum nocte cum corde meoet exercitabar et scobebam spiritum meum.
PS|77|8|Numquid in aeternum proiciet Deus,aut non apponet, ut complacitior sit adhuc?
PS|77|9|Aut deficiet in finem misericordia sua,cessabit verbum a generatione in generationem?
PS|77|10|Aut obliviscetur misereri Deus,aut continebit in ira sua misericordias suas?
PS|77|11|Et dixi: " Hoc vulnus meum:mutatio dexterae Excelsi ".
PS|77|12|Memor ero operum Domini,memor ero ab initio mirabilium tuorum.
PS|77|13|Et meditabor in omnibus operibus tuiset in adinventionibus tuis exercebor.
PS|77|14|Deus, in sancto via tua;quis deus magnus sicut Deus noster?
PS|77|15|Tu es Deus, qui facis mirabilia,notam fecisti in populis virtutem tuam.
PS|77|16|Redemisti in brachio tuo populum tuum,filios Iacob et Ioseph.
PS|77|17|Viderunt te aquae, Deus,viderunt te aquae et doluerunt;etenim commotae sunt abyssi.
PS|77|18|Effuderunt aquas nubila,vocem dederunt nubes,etenim sagittae tuae transeunt.
PS|77|19|Vox tonitrui tui in rota;illuxerunt coruscationes tuae orbi terrae,commota est et contremuit terra.
PS|77|20|In mari via tua, et semitae tuae in aquis multis;et vestigia tua non cognoscuntur.
PS|77|21|Deduxisti sicut oves populum tuumin manu Moysi et Aaron.
PS|78|1|Maskil. Asaph.Attendite, popule meus, doctrinam meam;inclinate aurem vestram in verba oris mei.
PS|78|2|Aperiam in parabolis os meum,eloquar arcana aetatis antiquae.
PS|78|3|Quanta audivimus et cognovimus ea,et patres nostri narraverunt nobis,
PS|78|4|non occultabimus a filiis eorum,generationi alteri narranteslaudes Domini et virtutes eiuset mirabilia eius, quae fecit.
PS|78|5|Constituit testimonium in Iacobet legem posuit in Israel;quanta mandaverat patribus nostrisnota facere ea filiis suis,
PS|78|6|ut cognoscat generatio altera,filii, qui nascentur.Exsurgent et narrabunt filiis suis,
PS|78|7|ut ponant in Deo spem suamet non obliviscantur operum Deiet mandata eius custodiant.
PS|78|8|Ne fiant sicut patres eorum,generatio rebellis et exasperans;generatio, quae non firmavit cor suum,et non fuit fidelis Deo spiritus eius.
PS|78|9|Filii Ephraim, intendentes et mittentes arcum,conversi sunt in die belli.
PS|78|10|Non custodierunt testamentum Deiet in lege eius renuerunt ambulare.
PS|78|11|Et obliti sunt factorum eiuset mirabilium eius, quae ostendit eis.
PS|78|12|Coram patribus eorum fecit mirabiliain terra Aegypti, in campo Taneos.
PS|78|13|Scidit mare et perduxit eoset statuit aquas quasi in utre.
PS|78|14|Et deduxit eos in nube per diemet per totam noctem in illuminatione ignis.
PS|78|15|Scidit petram in eremoet adaquavit eos velut abyssus multa.
PS|78|16|Et eduxit rivulos de petraet deduxit tamquam flumina aquas.
PS|78|17|Et apposuerunt adhuc peccare ei,in iram excitaverunt Excelsum in inaquoso.
PS|78|18|Et tentaverunt Deum in cordibus suis,petentes escas animabus suis;
PS|78|19|et contra Deum locuti sunt,dixerunt: " Numquid poterit Deus parare mensam in deserto? ".
PS|78|20|Ecce percussit petram, et fluxerunt aquae,et torrentes inundaverunt. Numquid et panem poterit dareaut parare carnes populo suo? ".
PS|78|21|Ideo audivit Dominus et exarsit,et ignis accensus est in Iacob,et ira ascendit in Israel.
PS|78|22|Quia non crediderunt in Deonec speraverunt in salutari eius.
PS|78|23|Verumtamen mandavit nubibus desuperet ianuas caeli aperuit;
PS|78|24|et pluit illis manna ad manducandumet panem caeli dedit eis:
PS|78|25|panem angelorum manducavit homo;cibaria misit eis ad abundantiam.
PS|78|26|Excitavit austrum in caeloet induxit in virtute sua africum;
PS|78|27|et pluit super eos sicut pulverem carneset sicut arenam maris volatilia pennata:
PS|78|28|et ceciderunt in medio castrorum eorum,circa tabernacula eorum.
PS|78|29|Et manducaverunt et saturati sunt nimis,et desiderium eorum attulit eis.
PS|78|30|Nondum recesserant a desiderio suo,adhuc escae eorum erant in ore ipsorum,
PS|78|31|et ira Dei ascendit super eoset occidit pingues eorumet electos Israel prostravit.
PS|78|32|In omnibus his peccaverunt adhucet non crediderunt in mirabilibus eius;
PS|78|33|et consumpsit in halitu dies eorumet annos eorum cum festinatione.
PS|78|34|Cum occideret eos, quaerebant eumet conversi veniebant diluculo ad eum;
PS|78|35|et rememorati sunt quia Deus adiutor est eorum,et Deus Excelsus redemptor eorum est.
PS|78|36|Et suaserunt ei in ore suoet lingua sua mentiti sunt ei;
PS|78|37|cor autem eorum non erat rectum cum eo,nec fideles erant in testamento eius.
PS|78|38|Ipse autem est misericorset propitiatur iniquitati et non disperdit.Saepe avertit iram suamet non accendit omnem furorem suum.
PS|78|39|Et recordatus est quia caro sunt,spiritus vadens et non rediens.
PS|78|40|Quoties exacerbaverunt eum in deserto,in iram concitaverunt eum in inaquoso!
PS|78|41|Et reversi sunt et tentaverunt Deumet Sanctum Israel exacerbaverunt.
PS|78|42|Non sunt recordati manus eius,diei, qua redemit eos de manu tribulantis.
PS|78|43|Cum posuit in Aegypto signa suaet prodigia sua in campo Taneos.
PS|78|44|Convertit in sanguinem flumina eorumet rivulos eorum, ne biberent.
PS|78|45|Misit in eos coenomyiam et comedit eos,ranam et perdidit eos.
PS|78|46|Dedit brucho fructus eorum,labores eorum locustae.
PS|78|47|Occidit in grandine vineas eorum,moros eorum in pruina.
PS|78|48|Tradidit grandini iumenta eorumet greges eorum flammae ignis.
PS|78|49|Misit in eos ardorem irae suae,indignationem et comminationem et angustiam,immissionem angelorum malorum.
PS|78|50|Complanavit semitam irae suae;non pepercit a morte animabus eorumet vitam eorum in peste conclusit.
PS|78|51|Percussit omne primogenitum in terra Aegypti,primitias roboris eorum in tabernaculis Cham.
PS|78|52|Abstulit sicut oves populum suumet perduxit eos tamquam gregem in deserto.
PS|78|53|Deduxit eos in spe, et non timuerunt,et inimicos eorum operuit mare.
PS|78|54|Et induxit eos in fines sanctificationis suae,in montem, quem acquisivit dextera eius.
PS|78|55|Et eiecit a facie eorum genteset divisit eis terram in funiculo hereditatiset habitare fecit in tabernaculis eorum tribus Israel.
PS|78|56|Et tentaverunt et exacerbaverunt Deum Excelsumet testimonia eius non custodierunt.
PS|78|57|Recesserunt et praevaricati sunt,quemadmodum patres eorum;conversi sunt retro ut arcus pravus.
PS|78|58|In iram concitaverunt eum in collibus suiset in sculptilibus suis ad aemulationem eum provocaverunt.
PS|78|59|Audivit Deus et exarsitet sprevit valde Israel.
PS|78|60|Et reppulit habitaculum Silo,tabernaculum, ubi habitavit in hominibus.
PS|78|61|Et tradidit in captivitatem virtutem suamet pulchritudinem suam in manus inimici.
PS|78|62|Et conclusit in gladio populum suumet in hereditatem suam exarsit.
PS|78|63|Iuvenes eorum comedit ignis,et virgines eorum non sunt desponsatae.
PS|78|64|Sacerdotes eorum in gladio ceciderunt,et viduae eorum non plorabantur.
PS|78|65|Et excitatus est tamquam dormiens Dominus,tamquam potens crapulatus a vino.
PS|78|66|Et percussit inimicos suos in posteriora,opprobrium sempiternum dedit illis.
PS|78|67|Et reppulit tabernaculum Iosephet tribum Ephraim non elegit,
PS|78|68|sed elegit tribum Iudae,montem Sion, quem dilexit.
PS|78|69|Et aedificavit sicut excelsum sanctuarium suum,sicut terram, quam fundavit in saecula.
PS|78|70|Et elegit David servum suumet sustulit eum de gregibus ovium,
PS|78|71|de post fetantes accepit eum:pascere Iacob populum suumet Israel hereditatem suam.
PS|78|72|Et pavit eos in innocentia cordis suiet in prudentia manuum suarum deduxit eos.
PS|79|1|PSALMUS. Asaph.Deus, venerunt gentes in hereditatem tuam,polluerunt templum sanctum tuum,posuerunt Ierusalem in ruinas.
PS|79|2|Dederunt morticina servorum tuorum escas volatilibus caeli,carnes sanctorum tuorum bestiis terrae.
PS|79|3|Effuderunt sanguinem eorum tamquam aquamin circuitu Ierusalem, et non erat qui sepeliret.
PS|79|4|Facti sumus opprobrium vicinis nostris,subsannatio et illusio his, qui in circuitu nostro sunt.
PS|79|5|Usquequo, Domine? Irasceris in finem?Accendetur velut ignis zelus tuus?
PS|79|6|Effunde iram tuam in gentes, quae te non noverunt,et in regna, quae nomen tuum non invocaverunt,
PS|79|7|quia comederunt Iacobet sedem eius desolaverunt.
PS|79|8|Ne memineris iniquitatum patrum nostrorum,cito anticipent nos misericordiae tuae,quia pauperes facti sumus nimis.
PS|79|9|Adiuva nos, Deus salutaris nostri,propter gloriam nominis tui et libera nos;et propitius esto peccatis nostris propter nomen tuum.
PS|79|10|Quare dicent in gentibus: " Ubi est Deus eorum? ".Innotescat in nationibus coram oculis nostrisultio sanguinis servorum tuorum, qui effusus est.
PS|79|11|Introeat in conspectu tuo gemitus compeditorum;secundum magnitudinem brachii tuisuperstites relinque filios mortis.
PS|79|12|Et redde vicinis nostris septuplum in sinu eorum,improperium ipsorum, quod exprobraverunt tibi, Domine.
PS|79|13|Nos autem, populus tuus et oves pascuae tuae,confitebimur tibi in saeculum;in generationem et generationem annuntiabimus laudem tuam.
PS|80|1|Magistro chori. Secundum " Lilium praecepti ".Asaph. PSALMUS.
PS|80|2|Qui pascis Israel, intende,qui deducis velut ovem Ioseph.Qui sedes super cherubim, effulge
PS|80|3|coram Ephraim, Beniamin et Manasse.Excita potentiam tuam et veni,ut salvos facias nos.
PS|80|4|Deus, converte nos,illustra faciem tuam, et salvi erimus.
PS|80|5|Domine, Deus virtutum,quousque irasceris super orationem populi tui?
PS|80|6|Cibasti nos pane lacrimarumet potum dedisti nobis in lacrimis copiose.
PS|80|7|Posuisti nos in contradictionem vicinis nostris,et inimici nostri subsannaverunt nos.
PS|80|8|Deus virtutum, converte nos,illustra faciem tuam, et salvi erimus.
PS|80|9|Vineam de Aegypto transtulisti,eiecisti gentes et plantasti eam.
PS|80|10|Purgasti locum in conspectu eius,plantasti radices eius, et implevit terram.
PS|80|11|Operti sunt montes umbra eius,et ramis eius cedri Dei;
PS|80|12|extendit palmites suos usque ad mareet usque ad flumen propagines suas.
PS|80|13|Ut quid destruxisti maceriam eius,et vindemiant eam omnes, qui praetergrediuntur viam?
PS|80|14|Exterminavit eam aper de silva,et singularis ferus depastus est eam.
PS|80|15|Deus virtutum, convertere,respice de caelo et vide et visita vineam istam.
PS|80|16|Et protege eam, quam plantavit dextera tua,et super filium hominis, quem confirmasti tibi.
PS|80|17|Incensa est igni et suffossa;ab increpatione vultus tui peribunt.
PS|80|18|Fiat manus tua super virum dexterae tuae,super filium hominis, quem confirmasti tibi.
PS|80|19|Et non discedemus a te, vivificabis nos,et nomen tuum invocabimus.
PS|80|20|Domine, Deus virtutum, converte noset illustra faciem tuam, et salvi erimus.
PS|81|1|Magistro chori. Secundum " Torcularia... ". Asaph.
PS|81|2|Exsultate Deo adiutori nostro;iubilate Deo Iacob.
PS|81|3|Sumite psalmum et date tympanum,psalterium iucundum cum cithara.
PS|81|4|Bucinate in neomenia tuba,in die plenae lunae, in sollemnitate nostra.
PS|81|5|Quia praeceptum in Israel est,et iudicium Deo Iacob.
PS|81|6|Testimonium in Ioseph posuit illud,cum exiret de terra Aegypti;sermonem, quem non noveram, audivi:
PS|81|7|" Diverti ab oneribus dorsum eius;manus eius a cophino recesserunt.
PS|81|8|In tribulatione invocasti me, et liberavi te,exaudivi te in abscondito tempestatis,probavi te apud aquam Meriba.
PS|81|9|Audi, populus meus, et contestabor te;Israel, utinam audias me!
PS|81|10|Non erit in te deus alienus,neque adorabis deum extraneum.
PS|81|11|Ego enim sum Dominus Deus tuus,qui eduxi te de terra Aegypti;dilata os tuum, et implebo illud.
PS|81|12|Et non audivit populus meus vocem meam,et Israel non intendit mihi.
PS|81|13|Et dimisi eos secundum duritiam cordis eorum,ibunt in adinventionibus suis.
PS|81|14|Si populus meus audisset me,Israel si in viis meis ambulasset!
PS|81|15|In brevi inimicos eorum humiliassemet super tribulantes eos misissem manum meam.
PS|81|16|Inimici Domini blandirentur ei,et esset sors eorum in saecula;
PS|81|17|et cibarem eos ex adipe frumentiet de petra melle saturarem eos ".
PS|82|1|PSALMUS. Asaph.Deus stetit in concilio divino,in medio deorum iudicat.
PS|82|2|" Usquequo iudicabitis iniqueet facies peccatorum sumetis?
PS|82|3|Iudicate egeno et pupillo,humilem et pauperem iustificate.
PS|82|4|Eripite pauperemet egenum de manu peccatoris liberate ".
PS|82|5|Nescierunt neque intellexerunt, in tenebris ambulant;movebuntur omnia fundamenta terrae.
PS|82|6|Ego dixi: " Dii estis,et filii Excelsi omnes ".
PS|82|7|Vos autem sicut homines morieminiet sicut unus de principibus cadetis.
PS|82|8|Surge, Deus, iudica terram,quoniam tu hereditabis in omnibus gentibus.
PS|83|1|Canticum. PSALMUS. Asaph.
PS|83|2|Deus, ne quiescas, ne taceasneque compescaris, Deus,
PS|83|3|quoniam ecce inimici tui fremuerunt,et, qui oderunt te, extulerunt caput.
PS|83|4|Adversus populum tuum malignaverunt consiliumet cogitaverunt adversus eos, quos abscondisti tibi.
PS|83|5|Dixerunt: " Venite, et disperdamus eos de gente,et non memoretur nomen Israel ultra! ".
PS|83|6|Quoniam cogitaverunt unanimiter,adversum te testamentum statuerunt:
PS|83|7|tabernacula Idumaeorum et Ismaelitae,Moab et Agareni,
PS|83|8|Gebal et Ammon et Amalec,Philistaea cum habitantibus Tyrum.
PS|83|9|Etenim Assur sociabatur cum illis;facti sunt in adiutorium filiis Lot.
PS|83|10|Fac illis sicut Madian et Sisarae,sicut Iabin in torrente Cison.
PS|83|11|Disperierunt in Endor,facti sunt ut stercus super terram.
PS|83|12|Pone duces eorum sicut Oreb et Zebet Zebee et Salmana, omnes principes eorum,
PS|83|13|qui dixerunt: Hereditate possideamus pascua Dei! ".
PS|83|14|Deus meus, pone illos ut rotamet sicut stipulam ante ventum.
PS|83|15|Sicut ignis, qui comburit silvam,et sicut flamma devorans montes,
PS|83|16|ita persequeris illos in tempestate tuaet in procella tua turbabis eos.
PS|83|17|Imple facies eorum ignominia,et quaerent nomen tuum, Domine.
PS|83|18|Erubescant et conturbentur in saeculum saeculiet confundantur et pereant;
PS|83|19|et cognoscant quia nomen tibi Dominus:tu solus Altissimus super omnem terram.
PS|84|1|Magistro chori. Secundum " Torcularia ".Filiorum Core. PSALMUS.
PS|84|2|Quam dilecta tabernacula tua, Domine virtutum!
PS|84|3|Concupiscit et deficit anima mea in atria Domini.Cor meum et caro mea exsultaverunt in Deum vivum.
PS|84|4|Etenim passer invenit sibi domum,et turtur nidum sibi, ubi ponat pullos suos:altaria tua, Domine virtutum, rex meus et Deus meus.
PS|84|5|Beati, qui habitant in domo tua:in perpetuum laudabunt te.
PS|84|6|Beatus vir, cuius est auxilium abs te,ascensiones in corde suo disposuit.
PS|84|7|Transeuntes per vallem sitientemin fontem ponent eam,etenim benedictionibus vestiet eam pluvia matutina.
PS|84|8|Ibunt de virtute in virtutem,videbitur Deus deorum in Sion.
PS|84|9|Domine, Deus virtutum, exaudi orationem meam;auribus percipe, Deus Iacob.
PS|84|10|Protector noster aspice, Deus,et respice in faciem christi tui.
PS|84|11|Quia melior est dies una in atriis tuis super milia,elegi ad limen esse in domo Dei meimagis quam habitare in tabernaculis peccatorum.
PS|84|12|Quia sol et scutum est Dominus Deus,gratiam et gloriam dabit Dominus;non privabit bonis eos,qui ambulant in innocentia.
PS|84|13|Domine virtutum, beatus homo, qui sperat in te.
PS|85|1|Magistro chori. Filiorum Core. PSALMUS.
PS|85|2|Complacuisti tibi, Domine, in terra tua,convertisti captivitatem Iacob.
PS|85|3|Remisisti iniquitatem plebis tuae,operuisti omnia peccata eorum.
PS|85|4|Contraxisti omnem iram tuam,revertisti a furore indignationis tuae.
PS|85|5|Converte nos, Deus, salutaris noster,et averte iram tuam a nobis.
PS|85|6|Numquid in aeternum irasceris nobisaut extendes iram tuam a generatione in generationem?
PS|85|7|Nonne tu conversus vivificabis nos,et plebs tua laetabitur in te?
PS|85|8|Ostende nobis, Domine, misericordiam tuamet salutare tuum da nobis.
PS|85|9|Audiam, quid loquatur Dominus Deus,quoniam loquetur pacem ad plebem suam et sanctos suoset ad eos, qui convertuntur corde.
PS|85|10|Vere prope timentes eum salutare ipsius,ut inhabitet gloria in terra nostra.
PS|85|11|Misericordia et veritas obviaverunt sibi,iustitia et pax osculatae sunt.
PS|85|12|Veritas de terra orta est,et iustitia de caelo prospexit.
PS|85|13|Etenim Dominus dabit benignitatem,et terra nostra dabit fructum suum.
PS|85|14|Iustitia ante eum ambulabitet ponet in via gressus suos.
PS|86|1|Precatio. David.Inclina, Domine, aurem tuam et exaudi me,quoniam inops et pauper sum ego.
PS|86|2|Custodi animam meam, quoniam sanctus sum;salvum fac servum tuum, Deus meus, sperantem in te
PS|86|3|Miserere mei, Domine, quoniam ad te clamavi tota die.
PS|86|4|Laetifica animam servi tui,quoniam ad te, Domine, animam meam levavi.
PS|86|5|Quoniam tu, Domine, suavis et mitiset multae misericordiae omnibus invocantibus te. -
PS|86|6|Auribus percipe, Domine, orationem meamet intende voci deprecationis meae.
PS|86|7|In die tribulationis meae clamavi ad te,quia exaudies me.
PS|86|8|Non est similis tui in diis, Domine,et nihil sicut opera tua.
PS|86|9|Omnes gentes, quascumque fecisti, venientet adorabunt coram te, Domine,et glorificabunt nomen tuum,
PS|86|10|quoniam magnus es tu et faciens mirabilia:tu es Deus solus.
PS|86|11|Doce me, Domine, viam tuam,et ingrediar in veritate tua;simplex fac cor meum,ut timeat nomen tuum.
PS|86|12|Confitebor tibi, Domine Deus meus, in toto corde meoet glorificabo nomen tuum in aeternum,
PS|86|13|quia misericordia tua magna est super me,et eruisti animam meam ex inferno inferiori.
PS|86|14|Deus, superbi insurrexerunt super me,et synagoga potentium quaesierunt animam meamet non proposuerunt te in conspectu suo.
PS|86|15|Et tu, Domine, Deus miserator et misericors,patiens et multae misericordiae et veritatis,
PS|86|16|respice in me et miserere mei;da fortitudinem tuam puero tuoet salvum fac filium ancillae tuae.
PS|86|17|Fac mecum signum in bonum,ut videant, qui oderunt me, et confundantur,quoniam tu, Domine, adiuvisti me et consolatus es me.
PS|87|1|Filiorum Core. PSALMUS. Canticum.Fundamenta eius in montibus sanctis;
PS|87|2|diligit Dominus portas Sionsuper omnia tabernacula Iacob.
PS|87|3|Gloriosa dicta sunt de te, civitas Dei! -
PS|87|4|Memor ero Rahab et Babylonis inter scientes me;ecce Philistaea et Tyrus cum Aethiopia:hi nati sunt illic.
PS|87|5|Et de Sion dicetur: " Hic et ille natus est in ea;et ipse firmavit eam Altissimus ".
PS|87|6|Dominus referet in librum populorum: Hi nati sunt illic ".
PS|87|7|Et cantant sicut choros ducentes: Omnes fontes mei in te ".
PS|88|1|Canticum. PSALMUS. Filiorum Core. Magistro chori.Secundum " Mahalat ". Ad cantandum. Maskil. Heman Ezrahitae.
PS|88|2|Domine, Deus salutis meae,in die clamavi et nocte coram te.
PS|88|3|Intret in conspectu tuo oratio mea;inclina aurem tuam ad precem meam.
PS|88|4|Quia repleta est malis anima mea,et vita mea inferno appropinquavit.
PS|88|5|Aestimatus sum cum descendentibus in lacum,factus sum sicut homo sine adiutorio.
PS|88|6|Inter mortuos liber,sicut vulnerati dormientes in sepulcris;quorum non es memor amplius,et ipsi de manu tua abscissi sunt.
PS|88|7|Posuisti me in lacu inferiori,in tenebrosis et in umbra mortis.
PS|88|8|Super me gravatus est furor tuus,et omnes fluctus tuos induxisti super me.
PS|88|9|Longe fecisti notos meos a me,posuisti me abominationem eis;conclusus sum et non egrediar.
PS|88|10|Oculi mei languerunt prae afflictione.Clamavi ad te, Domine, tota die,expandi ad te manus meas. -
PS|88|11|Numquid mortuis facies mirabilia,aut surgent umbrae et confitebuntur tibi?
PS|88|12|Numquid narrabit aliquis in sepulcro misericordiam tuamet veritatem tuam in loco perditionis?
PS|88|13|Numquid cognoscentur in tenebris mirabilia tua,et iustitia tua in terra oblivionis?
PS|88|14|Et ego ad te, Domine, clamavi,et mane oratio mea praeveniet te.
PS|88|15|Ut quid, Domine, repellis animam meam,abscondis faciem tuam a me?
PS|88|16|Pauper sum ego et moriens a iuventute mea;portavi pavores tuos et conturbatus sum.
PS|88|17|Super me transierunt irae tuae,et terrores tui exciderunt me.
PS|88|18|Circuierunt me sicut aqua tota die,circumdederunt me simul.
PS|88|19|Elongasti a me amicum et proximum,et noti mei sunt tenebrae.
PS|89|1|Maskil. Ethan Ezrahitae.
PS|89|2|Misericordias Domini in aeternum cantabo;in generationem et generationemannuntiabo veritatem tuam in ore meo.
PS|89|3|Quoniam dixisti: " In aeternum misericordia aedificabitur ",in caelis firmabitur veritas tua.
PS|89|4|" Disposui testamentum electo meo,iuravi David servo meo:
PS|89|5|Usque in aeternum confirmabo semen tuumet aedificabo in generationem et generationem sedem tuam ".
PS|89|6|Confitebuntur caeli mirabilia tua, Domine,etenim veritatem tuam in ecclesia sanctorum.
PS|89|7|Quoniam quis in nubibus aequabitur Domino,similis erit Domino in filiis Dei?
PS|89|8|Deus, metuendus in consilio sanctorum,magnus et terribilis super omnes, qui in circuitu eius sunt.
PS|89|9|Domine, Deus virtutum, quis similis tibi?Potens es, Domine, et veritas tua in circuitu tuo.
PS|89|10|Tu dominaris superbiae maris,elationes fluctuum eius tu mitigas.
PS|89|11|Tu conculcasti sicut vulneratum Rahab,in brachio virtutis tuae dispersisti inimicos tuos.
PS|89|12|Tui sunt caeli, et tua est terra,orbem terrae et plenitudinem eius tu fundasti;
PS|89|13|Aquilonem et austrum tu creasti,Thabor et Hermon in nomine tuo exsultabunt.
PS|89|14|Tibi brachium cum potentia;firma est manus tua, et exaltata dextera tua.
PS|89|15|Iustitia et iudicium firmamentum sedis tuae.Misericordia et veritas praecedent faciem tuam.
PS|89|16|Beatus populus, qui scit iubilationem.Domine, in lumine vultus tui ambulabunt
PS|89|17|et in nomine tuo exsultabunt tota die et in iustitia tua exaltabuntur,
PS|89|18|quoniam decor virtutis eorum tu es,et in beneplacito tuo exaltabitur cornu nostrum.
PS|89|19|Quia Domini est scutum nostrum,et Sancti Israel rex noster.
PS|89|20|Tunc locutus es in visione sanctis tuis et dixisti: Posui adiutorium in potenteet exaltavi electum de plebe.
PS|89|21|Inveni David servum meum;oleo sancto meo unxi eum.
PS|89|22|Manus enim mea firma erit cum eo, et brachium meum confortabit eum.
PS|89|23|Nihil proficiet inimicus in eo,et filius iniquitatis non opprimet eum.
PS|89|24|Et concidam a facie ipsius inimicos eiuset odientes eum percutiam.
PS|89|25|Et veritas mea et misericordia mea cum ipso,et in nomine meo exaltabitur cornu eius.
PS|89|26|Et ponam super mare manum eiuset super flumina dexteram eius.
PS|89|27|Ipse invocabit me: "Pater meus es tu,Deus meus et refugium salutis meae".
PS|89|28|Et ego primogenitum ponam illum,excelsum prae regibus terrae.
PS|89|29|In aeternum servabo illi misericordiam meam;et testamentum meum fidele ipsi.
PS|89|30|Et ponam in saeculum saeculi semen eius;et thronum eius sicut dies caeli.
PS|89|31|Si autem dereliquerint filii eius legem meamet in iudiciis meis non ambulaverint,
PS|89|32|si iustificationes meas profanaverintet mandata mea non custodierint,
PS|89|33|visitabo in virga delictum eorumet in verberibus iniquitatem eorum.
PS|89|34|Misericordiam autem meam non avertam ab eoneque mentiar in veritate mea.
PS|89|35|Non profanabo testamentum meum et, quae procedunt de labiis meis, non faciam irrita.
PS|89|36|Semel iuravi in sancto meo: David non mentiar.
PS|89|37|Semen eius in aeternum manebit,et thronus eius sicut sol in conspectu meo
PS|89|38|et sicut luna firmus stabit in aeternumet testis in caelo fidelis ".
PS|89|39|Tu vero reppulisti et reiecisti,iratus es contra christum tuum;
PS|89|40|evertisti testamentum servi tui,profanasti in terram diadema eius.
PS|89|41|Destruxisti omnes muros eius,posuisti munitiones eius in ruinas.
PS|89|42|Diripuerunt eum omnes transeuntes viam,factus est opprobrium vicinis suis.
PS|89|43|Exaltasti dexteram deprimentium eum,laetificasti omnes inimicos eius.
PS|89|44|Avertisti aciem gladii eiuset non es auxiliatus ei in bello.
PS|89|45|Finem posuisti splendori eiuset sedem eius in terram collisisti.
PS|89|46|Minorasti dies iuventutis eius,perfudisti eum confusione.
PS|89|47|Usquequo, Domine, absconderis in finem,exardescet sicut ignis ira tua?
PS|89|48|Memorare, quam brevis mea substantia.Ad quam vanitatem creasti omnes filios hominum?
PS|89|49|Quis est homo, qui vivet et non videbit mortem,eruet animam suam de manu inferi?
PS|89|50|Ubi sunt misericordiae tuae antiquae, Domine,sicut iurasti David in veritate tua?
PS|89|51|Memor esto, Domine, opprobrii servorum tuorum,quod continui in sinu meo, multarum gentium,
PS|89|52|quo exprobraverunt inimici tui, Domine,quo exprobraverunt vestigia christi tui.
PS|89|53|Benedictus Dominus in aeternum. Fiat, fiat.
PS|90|1|Precatio. Moysis viri Dei. Domine, refugium factus es nobisa generatione in generationem.
PS|90|2|Priusquam montes nascerentur, aut gigneretur terra et orbis,a saeculo et usque in saeculum tu es Deus.
PS|90|3|Reducis hominem in pulverem;et dixisti: " Revertimini, filii hominum ".
PS|90|4|Quoniam mille anni ante oculos tuostamquam dies hesterna, quae praeteriit,et custodia in nocte.
PS|90|5|Auferes eos, somnium erunt:
PS|90|6|mane sicut herba succrescens,mane floret et crescit,vespere decidit et arescit.
PS|90|7|Quia defecimus in ira tuaet in furore tuo turbati sumus.
PS|90|8|Posuisti iniquitates nostras in conspectu tuo,occulta nostra in illuminatione vultus tui.
PS|90|9|Quoniam omnes dies nostri evanuerunt in ira tua,consumpsimus ut suspirium annos nostros.
PS|90|10|Dies annorum nostrorum sunt septuaginta anniaut in valentibus octoginta anni,et maior pars eorum labor et dolor,quoniam cito transeunt, et avolamus.
PS|90|11|Quis novit potestatem irae tuaeet secundum timorem tuum indignationem tuam?
PS|90|12|Dinumerare dies nostros sic doce nos, ut inducamus cor ad sapientiam.
PS|90|13|Convertere, Domine, usquequo?Et deprecabilis esto super servos tuos.
PS|90|14|Reple nos mane misericordia tua,et exsultabimus et delectabimur omnibus diebus nostris.
PS|90|15|Laetifica nos pro diebus, quibus nos humiliasti,pro annis, quibus vidimus mala.
PS|90|16|Appareat servis tuis opus tuum,et decor tuus filiis eorum.
PS|90|17|Et sit splendor Domini Dei nostri super nos,et opera manuum nostrarum confirma super noset opus manuum nostrarum confirma.
PS|91|1|Qui habitat in protectione Altissimi,sub umbra Omnipotentis commorabitur.
PS|91|2|Dicet Domino: " Refugium meumet fortitudo mea, Deus meus, sperabo in eum ".
PS|91|3|Quoniam ipse liberabit te de laqueo venantiumet a verbo maligno.
PS|91|4|Alis suis obumbrabit tibi,et sub pennas eius confugies;scutum et lorica veritas eius.
PS|91|5|Non timebis a timore nocturno,a sagitta volante in die,
PS|91|6|a peste perambulante in tenebris,ab exterminio vastante in meridie.
PS|91|7|Cadent a latere tuo milleet decem milia a dextris tuis;ad te autem non appropinquabit.
PS|91|8|Verumtamen oculis tuis considerabiset retributionem peccatorum videbis.
PS|91|9|Quoniam tu es, Domine, refugium meum.Altissimum posuisti habitaculum tuum.
PS|91|10|Non accedet ad te malum,et flagellum non appropinquabit tabernaculo tuo,
PS|91|11|quoniam angelis suis mandabit de te,ut custodiant te in omnibus viis tuis.
PS|91|12|In manibus portabunt te,ne forte offendas ad lapidem pedem tuum.
PS|91|13|Super aspidem et basiliscum ambulabiset conculcabis leonem et draconem.
PS|91|14|Quoniam mihi adhaesit, liberabo eum;suscipiam eum, quoniam cognovit nomen meum.
PS|91|15|Clamabit ad me, et ego exaudiam eum;cum ipso sum in tribulatione;eripiam eum et glorificabo eum.
PS|91|16|Longitudine dierum replebo eumet ostendam illi salutare meum.
PS|92|1|PSALMUS. Canticum. Pro die Sabbati.
PS|92|2|Bonum est confiteri Dominoet psallere nomini tuo, Altissime,
PS|92|3|annuntiare mane misericordiam tuamet veritatem tuam per noctem
PS|92|4|in decachordo et psalterio,cum cantico in cithara.
PS|92|5|Quia delectasti me, Domine, in factura tua,et in operibus manuum tuarum exsultabo.
PS|92|6|Quam magnificata sunt opera tua, Domine:nimis profundae factae sunt cogitationes tuae.
PS|92|7|Vir insipiens non cognoscet,et stultus non intelleget haec.
PS|92|8|Cum germinaverint peccatores sicut fenum,et floruerint omnes, qui operantur iniquitatem,hoc tamen erit ad interitum in saeculum saeculi;
PS|92|9|tu autem altissimus in aeternum, Domine.
PS|92|10|Quoniam ecce inimici tui, Domine,quoniam ecce inimici tui peribunt,et dispergentur omnes, qui operantur iniquitatem.
PS|92|11|Exaltabis sicut unicornis cornu meum,perfusus sum oleo uberi.
PS|92|12|Et despiciet oculus meus inimicos meos,et in insurgentibus in me malignantibus audiet auris mea. -
PS|92|13|Iustus ut palma florebit,sicut cedrus Libani succrescet.
PS|92|14|Plantati in domo Domini,in atriis Dei nostri florebunt.
PS|92|15|Adhuc fructus dabunt in senecta,uberes et bene virentes erunt,
PS|92|16|ut annuntient quoniam rectus Dominus,refugium meum, et non est iniquitas in eo.
PS|93|1|Dominus regnavit! Decorem indutus est;indutus est Dominus, fortitudine praecinxit se.Etenim firmavit orbem terrae, qui non commovebitur.
PS|93|2|Firmata sedes tua ex tunc,a saeculo tu es.
PS|93|3|Elevaverunt flumina, Domine.elevaverunt flumina vocem suam,elevaverunt flumina fragorem suum.
PS|93|4|Super voces aquarum multarum,super potentes elationes maris,potens in altis Dominus.
PS|93|5|Testimonia tua credibilia facta sunt nimis;domum tuam decet sanctitudo Domine,in longitudinem dierum.
PS|94|1|Deus ultionum, Domine,Deus ultionum, effulge.
PS|94|2|Exaltare, qui iudicas terram,redde retributionem superbis.
PS|94|3|Usquequo peccatores, Domine,usquequo peccatores exsultabunt?
PS|94|4|Effabuntur et loquentur proterva,gloriabuntur omnes, qui operantur iniquitatem. -
PS|94|5|Populum tuum, Domine, humiliantet hereditatem tuam vexant.
PS|94|6|Viduam et advenam interficiuntet pupillos occidunt.
PS|94|7|Et dixerunt: " Non videbit Dominus,nec intelleget Deus Iacob ".
PS|94|8|Intellegite, insipientes in populo;et stulti, quando sapietis?
PS|94|9|Qui plantavit aurem, non audiet,aut qui finxit oculum, non respiciet?
PS|94|10|Qui corripit gentes, non arguet,qui docet hominem scientiam?
PS|94|11|Dominus scit cogitationes hominum,quoniam vanae sunt.
PS|94|12|Beatus homo, quem tu erudieris, Domine,et de lege tua docueris eum,
PS|94|13|ut mitiges ei a diebus malis,donec fodiatur peccatori fovea.
PS|94|14|Quia non repellet Dominus plebem suamet hereditatem suam non derelinquet.
PS|94|15|Quia ad iustitiam revertetur iudicium,et sequentur illam omnes, qui recto sunt corde.
PS|94|16|Quis consurget mihi adversus malignantes,aut quis stabit mecum adversus operantes iniquitatem?
PS|94|17|Nisi quia Dominus adiuvit me,paulo minus habitasset in loco silentii anima mea.
PS|94|18|Si dicebam: " Motus est pes meus ", misericordia tua, Domine, sustentabat me.
PS|94|19|In multitudine sollicitudinum mearum in corde meo,consolationes tuae laetificaverunt animam meam.
PS|94|20|Numquid sociabitur tibi sedes iniquitatis,quae fingit molestiam contra praeceptum?
PS|94|21|Irruunt in animam iustiet sanguinem innocentem condemnant.
PS|94|22|Et factus est mihi Dominus in praesidium,et Deus meus in rupem refugii mei;
PS|94|23|et reddet illis iniquitatem ipsorumet in malitia eorum disperdet eos,
PS|94|24|disperdet illos Dominus Deus noster.
PS|95|1|Venite, exsultemus Domino;iubilemus Deo salutari nostro.
PS|95|2|Praeoccupemus faciem eius in confessioneet in psalmis iubilemus ei.
PS|95|3|Quoniam Deus magnus Dominus,et rex magnus super omnes deos.
PS|95|4|Quia in manu eius sunt profunda terrae,et altitudines montium ipsius sunt.
PS|95|5|Quoniam ipsius est mare, et ipse fecit illud,et siccam manus eius formaverunt.
PS|95|6|Venite, adoremus et procidamuset genua flectamus ante Dominum, qui fecit nos,
PS|95|7|quia ipse est Deus noster,et nos populus pascuae eius et oves manus eius.
PS|95|8|Utinam hodie vocem eius audiatis: Nolite obdurare corda vestra,
PS|95|9|sicut in Meriba, secundum diem Massa in deserto,ubi tentaverunt me patres vestri:probaverunt me, etsi viderunt opera mea.
PS|95|10|Quadraginta annis taeduit me generationis illiuset dixi: Populus errantium corde sunt isti.
PS|95|11|Et ipsi non cognoverunt vias meas;ideo iuravi in ira mea:Non introibunt in requiem meam ".
PS|96|1|Cantate Domino canticum novum,cantate Domino, omnis terra.
PS|96|2|Cantate Domino, benedicite nomini eius,annuntiate de die in diem salutare eius.
PS|96|3|Annuntiate inter gentes gloriam eius,in omnibus populis mirabilia eius.
PS|96|4|Quoniam magnus Dominus et laudabilis nimis,terribilis est super omnes deos.
PS|96|5|Quoniam omnes dii gentium inania,Dominus autem caelos fecit.
PS|96|6|Magnificentia et pulchritudo in conspectu eius,potentia et decor in sanctuario eius.
PS|96|7|Afferte Domino, familiae populorum,afferte Domino gloriam et potentiam,
PS|96|8|afferte Domino gloriam nominis eius.Tollite hostias et introite in atria eius,
PS|96|9|adorate Dominum in splendore sancto.Contremiscite a facie eius, universa terra;
PS|96|10|dicite in gentibus: " Dominus regnavit! ".Etenim correxit orbem terrae, qui non commovebitur;iudicabit populos in aequitate.
PS|96|11|Laetentur caeli, et exsultet terra,sonet mare et plenitudo eius;
PS|96|12|gaudebunt campi et omnia, quae in eis sunt.Tunc exsultabunt omnia ligna silvarum
PS|96|13|a facie Domini, quia venit,quoniam venit iudicare terram.Iudicabit orbem terrae in iustitiaet populos in veritate sua.
PS|97|1|Dominus regnavit! Exsultet terra,laetentur insulae multae.
PS|97|2|Nubes et caligo in circuitu eius,iustitia et iudicium firmamentum sedis eius.
PS|97|3|Ignis ante ipsum praecedetet inflammabit in circuitu inimicos eius.
PS|97|4|Illustrarunt fulgura eius orbem terrae:vidit et contremuit terra.
PS|97|5|Montes sicut cera fluxerunt a facie Domini,a facie Domini omnis terra.
PS|97|6|Annuntiaverunt caeli iustitiam eius,et viderunt omnes populi gloriam eius.
PS|97|7|Confundantur omnes, qui adorant sculptilia,et qui gloriantur in simulacris suis.Adorate eum, omnes angeli eius.
PS|97|8|Audivit et laetata est Sion,et exsultaverunt filiae Iudaepropter iudicia tua, Domine.
PS|97|9|Quoniam tu Dominus, Altissimus super omnem terram,nimis exaltatus es super omnes deos.
PS|97|10|Qui diligitis Dominum, odite malum;custodit ipse animas sanctorum suorum,de manu peccatoris liberabit eos.
PS|97|11|Lux orta est iusto,et rectis corde laetitia.
PS|97|12|Laetamini, iusti, in Dominoet confitemini memoriae sanctitatis eius.
PS|98|1|PSALMUS.Cantate Domino canticum novum,quia mirabilia fecit.Salvavit sibi dextera eius,et brachium sanctum eius.
PS|98|2|Notum fecit Dominus salutare suum,in conspectu gentium revelavit iustitiam suam.
PS|98|3|Recordatus est misericordiae suaeet veritatis suae domui Israel.Viderunt omnes termini terraesalutare Dei nostri.
PS|98|4|Iubilate Deo, omnis terra;erumpite, exsultate et psallite.
PS|98|5|Psallite Domino in cithara,in cithara et voce psalmi;
PS|98|6|in tubis ductilibus et voce tubae corneae,iubilate in conspectu regis Domini.
PS|98|7|Sonet mare et plenitudo eius,orbis terrarum et qui habitant in eo.
PS|98|8|Flumina plaudent manu,simul montes exsultabunt
PS|98|9|a conspectu Domini, quoniam venit iudicare terram.Iudicabit orbem terrarum in iustitiaet populos in aequitate.
PS|99|1|Dominus regnavit! Commoveantur populisedet super cherubim, moveatur terra.
PS|99|2|Dominus in Sion magnuset excelsus super omnes populos.
PS|99|3|Confiteantur nomini tuo magno et terribili,quoniam sanctum est.
PS|99|4|Rex potens iudicium diligit:tu statuisti, quae recta sunt,iudicium et iustitiam in Iacob tu fecisti.
PS|99|5|Exaltate Dominum Deum nostrumet adorate ad scabellum pedum eius,quoniam sanctus est.
PS|99|6|Moyses et Aaron in sacerdotibus eius,et Samuel inter eos, qui invocant nomen eius.Invocabant Dominum, et ipse exaudiebat eos,
PS|99|7|in columna nubis loquebatur ad eos.Custodiebant testimonia eiuset praeceptum, quod dedit illis.
PS|99|8|Domine Deus noster, tu exaudiebas eos;Deus, tu propitius fuisti eis,ulciscens autem adinventiones eorum.
PS|99|9|Exaltate Dominum Deum nostrumet adorate ad montem sanctum eius,quoniam sanctus Dominus Deus noster.
PS|100|1|PSALMUS. Ad gratiarum actionem.
PS|100|2|Iubilate Domino, omnis terra,servite Domino in laetitia;introite in conspectu eius in exsultatione.
PS|100|3|Scitote quoniam Dominus ipse est Deus;ipse fecit nos, et ipsius sumus,populus eius et oves pascuae eius.
PS|100|4|Introite portas eius in confessione,atria eius in hymnis,confitemini illi, benedicite nomini eius.
PS|100|5|Quoniam suavis est Dominus;in aeternum misericordia eius,et usque in generationem et generationem veritas eius.
PS|101|1|David. PSALMUS.Misericordiam et iudicium cantabo;tibi, Domine, psallam.
PS|101|2|Intellegam in via immaculata;quando venies ad me?Perambulabo in innocentia cordis mei,in medio domus meae.
PS|101|3|Non proponam ante oculos meos rem iniustam;facientem praevaricationes odio habebo,non adhaerebit mihi.
PS|101|4|Cor pravum recedet a me,malignum non cognoscam.
PS|101|5|Detrahentem secreto proximo suo,hunc cessare faciam;superbum oculo et inflatum corde,hunc non sustinebo.
PS|101|6|Oculi mei ad fideles terrae, ut sedeant mecum;qui ambulat in via immaculata, hic mihi ministrabit.
PS|101|7|Non habitabit in medio domus meae, qui facit superbiam;qui loquitur iniqua, non stabit in conspectu oculorum meorum.
PS|101|8|In matutino cessare faciam omnes peccatores terrae,ut disperdam de civitate Domini omnes operantes iniquitatem.
PS|102|1|Preces afflicti, qui defessusangorem suum ante Dominum profundit.
PS|102|2|Domine, exaudi orationem meam,et clamor meus ad te veniat.
PS|102|3|Non abscondas faciem tuam a me;in quacumque die tribulor,inclina ad me aurem tuam.In quacumque die invocavero te,velociter exaudi me.
PS|102|4|Quia defecerunt sicut fumus dies mei,et ossa mea sicut cremium aruerunt.
PS|102|5|Percussum est ut fenum et aruit cor meum,etenim oblitus sum comedere panem meum.
PS|102|6|A voce gemitus meiadhaesit os meum carni meae.
PS|102|7|Similis factus sum pellicano solitudinis,factus sum sicut nycticorax in ruinis.
PS|102|8|Vigilavi et factus sum sicut passer solitarius in tecto.
PS|102|9|Tota die exprobrabant mihi inimici mei,exardescentes in me per me iurabant.
PS|102|10|Quia cinerem tamquam panem manducabamet potum meum cum fletu miscebam,
PS|102|11|a facie irae et increpationis tuae,quia elevans allisisti me.
PS|102|12|Dies mei sicut umbra declinaverunt,et ego sicut fenum arui.
PS|102|13|Tu autem, Domine, in aeternum permanes,et memoriale tuum in generationem et generationem.
PS|102|14|Tu exsurgens misereberis Sion,quia tempus miserendi eius,quia venit tempus,
PS|102|15|quoniam placuerunt servis tuis lapides eius,et pulveris eius miserentur.
PS|102|16|Et timebunt gentes nomen tuum, Domine,et omnes reges terrae gloriam tuam,
PS|102|17|quia aedificavit Dominus Sionet apparuit in gloria sua.
PS|102|18|Respexit in orationem inopumet non sprevit precem eorum.
PS|102|19|Scribantur haec pro generatione altera,et populus, qui creabitur, laudabit Dominum.
PS|102|20|Quia prospexit de excelso sanctuario suo,Dominus de caelo in terram aspexit,
PS|102|21|ut audiret gemitus compeditorum, ut solveret filios mortis;
PS|102|22|ut annuntient in Sion nomen Dominiet laudem eius in Ierusalem,
PS|102|23|cum congregati fuerint populi in unumet regna, ut serviant Domino.
PS|102|24|Humiliavit in via virtutem meam,abbreviavit dies meos.Dicam: " Deus meus,
PS|102|25|ne auferas me in dimidio dierum meorum;in generationem et generationem sunt anni tui.
PS|102|26|Initio terram fundasti;et opera manuum tuarum sunt caeli.
PS|102|27|Ipsi peribunt, tu autem permanes;et omnes sicut vestimentum veterascent,et sicut opertorium mutabis eos, et mutabuntur.
PS|102|28|Tu autem idem ipse es, et anni tui non deficient.
PS|102|29|Filii servorum tuorum habitabunt,et semen eorum in conspectu tuo firmabitur ".
PS|103|1|David.Benedic, anima mea, Domino,et omnia, quae intra me sunt, nomini sancto eius.
PS|103|2|Benedic, anima mea, Dominoet noli oblivisci omnes retributiones eius.
PS|103|3|Qui propitiatur omnibus iniquitatibus tuis,qui sanat omnes infirmitates tuas;
PS|103|4|qui redimit de interitu vitam tuam,qui coronat te in misericordia et miserationibus;
PS|103|5|qui replet in bonis aetatem tuam:renovabitur ut aquilae iuventus tua.
PS|103|6|Faciens iustitias Dominuset iudicium omnibus iniuriam patientibus.
PS|103|7|Notas fecit vias suas Moysi,filiis Israel adinventiones suas. -
PS|103|8|Miserator et misericors Dominus,longanimis et multae misericordiae.
PS|103|9|Non in perpetuum contendetneque in aeternum irascetur.
PS|103|10|Non secundum peccata nostra fecit nobisneque secundum iniquitates nostras retribuit nobis.
PS|103|11|Quoniam, quantum exaltatur caelum a terra,praevaluit misericordia eius super timentes eum;
PS|103|12|quantum distat ortus ab occidente,longe fecit a nobis iniquitates nostras.
PS|103|13|Quomodo miseretur pater filiorum,misertus est Dominus timentibus se.
PS|103|14|Quoniam ipse cognovit figmentum nostrum,recordatus est quoniam pulvis sumus.
PS|103|15|Homo: sicut fenum dies eius,tamquam flos agri sic efflorebit.
PS|103|16|Spirat ventus in illum, et non subsistet,et non cognoscet eum amplius locus eius.
PS|103|17|Misericordia autem Domini ab aeternoet usque in aeternum super timentes eum;et iustitia illius in filios filiorum,
PS|103|18|in eos, qui servant testamentum eiuset memores sunt mandatorum ipsius ad faciendum ea.
PS|103|19|Dominus in caelo paravit sedem suam,et regnum ipsius omnibus dominabitur.
PS|103|20|Benedicite Domino, omnes angeli eius, potentes virtute, facientes verbum illiusin audiendo vocem sermonum eius.
PS|103|21|Benedicite Domino, omnes virtutes eius,ministri eius, qui facitis voluntatem eius.
PS|103|22|Benedicite Domino, omnia opera eius,in omni loco dominationis eius.Benedic, anima mea, Domino.
PS|104|1|Benedic, anima mea, Domino.Domine Deus meus, magnificatus es vehementer!Maiestatem et decorem induisti,
PS|104|2|amictus lumine sicut vestimento.Extendens caelum sicut velum,
PS|104|3|qui exstruis in aquis cenacula tua.Qui ponis nubem ascensum tuum,qui ambulas super pennas ventorum.
PS|104|4|Qui facis angelos tuos spirituset ministros tuos ignem urentem.
PS|104|5|Qui fundasti terram super stabilitatem suam,non inclinabitur in saeculum saeculi.
PS|104|6|Abyssus sicut vestimentum operuit eam,super montes stabant aquae.
PS|104|7|Ab increpatione tua fugiunt,a voce tonitrui tui formidant.
PS|104|8|Ascendunt in montes et descendunt in valles,in locum, quem statuisti eis.
PS|104|9|Terminum posuisti, quem non transgredientur,neque convertentur operire terram.
PS|104|10|Qui emittis fontes in torrentes;inter medium montium pertransibunt,
PS|104|11|potabunt omnes bestias agri,exstinguent onagri sitim suam.
PS|104|12|Super ea volucres caeli habitabunt,de medio ramorum dabunt voces.
PS|104|13|Rigas montes de cenaculis tuis,de fructu operum tuorum satias terram.
PS|104|14|Producis fenum iumentiset herbam servituti hominum,educens panem de terra
PS|104|15|et vinum, quod laetificat cor hominis;exhilarans faciem in oleo,panis autem cor hominis confirmat.
PS|104|16|Saturabuntur ligna Dominiet cedri Libani, quas plantavit.
PS|104|17|Illic passeres nidificabunt,erodii domus in vertice earum.
PS|104|18|Montes excelsi cervis,petrae refugium hyracibus.
PS|104|19|Fecit lunam ad tempora signanda,sol cognovit occasum suum.
PS|104|20|Posuisti tenebras, et facta est nox:in ipsa reptabunt omnes bestiae silvae,
PS|104|21|catuli leonum rugientes, ut rapiantet quaerant a Deo escam sibi.
PS|104|22|Oritur sol, et congreganturet in cubilibus suis recumbunt.
PS|104|23|Exit homo ad opus suumet ad operationem suam usque ad vesperum.
PS|104|24|Quam multiplicata sunt opera tua, Domine!Omnia in sapientia fecisti,impleta est terra creatura tua.
PS|104|25|Hoc mare magnum et spatiosum et latum:illic reptilia, quorum non est numerus,animalia pusilla cum magnis;
PS|104|26|illic naves pertransibunt,Leviathan, quem formasti ad ludendum cum eo.
PS|104|27|Omnia a te exspectant,ut des illis escam in tempore suo.
PS|104|28|Dante te illis, colligent,aperiente te manum tuam, implebuntur bonis.
PS|104|29|Avertente autem te faciem, turbabuntur;auferes spiritum eorum, et deficientet in pulverem suum revertentur.
PS|104|30|Emittes spiritum tuum, et creabuntur,et renovabis faciem terrae.
PS|104|31|Sit gloria Domini in saeculum;laetetur Dominus in operibus suis.
PS|104|32|Qui respicit terram et facit eam tremere,qui tangit montes, et fumigant.
PS|104|33|Cantabo Domino in vita mea,psallam Deo meo quamdiu sum.
PS|104|34|Iucundum sit ei eloquium meum,ego vero delectabor in Domino.
PS|104|35|Deficiant peccatores a terraet iniqui, ita ut non sint.Benedic, anima mea, Domino.
PS|105|1|ALLELUIA.Confitemini Domino et invocate nomen eius,annuntiate inter gentes opera eius.
PS|105|2|Cantate ei et psallite ei,meditamini in omnibus mirabilibus eius.
PS|105|3|Laudamini in nomine sancto eius,laetetur cor quaerentium Dominum.
PS|105|4|Quaerite Dominum et potentiam eius,quaerite faciem eius semper.
PS|105|5|Mementote mirabilium eius, quae fecit,prodigia eius et iudicia oris eius,
PS|105|6|semen Abraham, servi eius,filii Iacob, electi eius.
PS|105|7|Ipse Dominus Deus noster;in universa terra iudicia eius.
PS|105|8|Memor fuit in saeculum testamenti sui,verbi, quod mandavit in mille generationes,
PS|105|9|quod disposuit cum Abraham,et iuramenti sui ad Isaac.
PS|105|10|Et statuit illud Iacob in praeceptumet Israel in testamentum aeternum
PS|105|11|dicens: " Tibi dabo terram Chanaanfuniculum hereditatis vestrae ".
PS|105|12|Cum essent numero brevi,paucissimi et peregrini in ea,
PS|105|13|et pertransirent de gente in gentemet de regno ad populum alterum,
PS|105|14|non permisit hominem nocere eiset corripuit pro eis reges:
PS|105|15|" Nolite tangere christos meoset in prophetis meis nolite malignari ".
PS|105|16|Et vocavit famem super terramet omne baculum panis contrivit.
PS|105|17|Misit ante eos virum,in servum venumdatus est Ioseph.
PS|105|18|Strinxerunt in compedibus pedes eius,in ferrum intravit collum eius,
PS|105|19|donec veniret verbum eius,eloquium Domini purgaret eum.
PS|105|20|Misit rex et solvit eum,princeps populorum, et dimisit eum;
PS|105|21|constituit eum dominum domus suaeet principem omnis possessionis suae,
PS|105|22|ut erudiret principes eius sicut semetipsumet senes eius prudentiam doceret.
PS|105|23|Et intravit Israel in Aegyptum,et Iacob peregrinus fuit in terra Cham.
PS|105|24|Et auxit populum suum vehementeret confortavit eum super inimicos eius.
PS|105|25|Convertit cor eorum, ut odirent populum eiuset dolum facerent in servos eius.
PS|105|26|Misit Moysen servum suum,Aaron, quem elegit.
PS|105|27|Posuit in eis verba signorum suorumet prodigiorum in terra Cham.
PS|105|28|Misit tenebras et obscuravit,et restiterunt sermonibus eius.
PS|105|29|Convertit aquas eorum in sanguinemet occidit pisces eorum.
PS|105|30|Edidit terra eorum ranasin penetralibus regum ipsorum.
PS|105|31|Dixit, et venit coenomyiaet scinifes in omnibus finibus eorum.
PS|105|32|Posuit pluvias eorum grandinem,ignem comburentem in terra ipsorum.
PS|105|33|Et percussit vineas eorum et ficulneas eorumet contrivit lignum finium eorum.
PS|105|34|Dixit, et venit locustaet bruchus, cuius non erat numerus,
PS|105|35|et comedit omne fenum in terra eorumet comedit fructum terrae eorum.
PS|105|36|Et percussit omne primogenitum in terra eorum,primitias omnis roboris eorum.
PS|105|37|Et eduxit eos cum argento et auro;et non erat in tribubus eorum infirmus.
PS|105|38|Laetata est Aegyptus in profectione eorum,quia incubuit timor eorum super eos.
PS|105|39|Expandit nubem in protectionemet ignem, ut luceret eis per noctem.
PS|105|40|Petierunt, et venit coturnix,et pane caeli saturavit eos.
PS|105|41|Dirupit petram, et fluxerunt aquae,abierunt in sicco flumina.
PS|105|42|Quoniam memor fuit verbi sancti suiad Abraham puerum suum.
PS|105|43|Et eduxit populum suum in exsultatione,electos suos in laetitia.
PS|105|44|Et dedit illis regiones gentium,et labores populorum possederunt,
PS|105|45|ut custodiant iustificationes eiuset leges eius servent.ALLELUIA.
PS|106|1|ALLELUIA.Confitemini Domino, quoniam bonus,quoniam in saeculum misericordia eius.
PS|106|2|Quis loquetur potentias Domini,auditas faciet omnes laudes eius?
PS|106|3|Beati, qui custodiunt iudiciumet faciunt iustitiam in omni tempore.
PS|106|4|Memento nostri, Domine, in beneplacito populi tui,visita nos in salutari tuo,
PS|106|5|ut videamus bona electorum tuorum,ut laetemur in laetitia gentis tuae,ut gloriemur cum hereditate tua.
PS|106|6|Peccavimus cum patribus nostris,iniuste egimus, iniquitatem fecimus.
PS|106|7|Patres nostri in Aegypto non intellexerunt mirabilia tua,non fuerunt memores multitudinis misericordiarum tuarumet irritaverunt ascendentes in mare, mare Rubrum.
PS|106|8|Et salvavit eos propter nomen suum,ut notam faceret potentiam suam. -
PS|106|9|Et increpuit mare Rubrum, et exsiccatum est,et deduxit eos in abyssis sicut in deserto.
PS|106|10|Et salvavit eos de manu odientiset redemit eos de manu inimici.
PS|106|11|Et operuit aqua tribulantes eos:unus ex eis non remansit.
PS|106|12|Et crediderunt verbis eiuset cantaverunt laudem eius.
PS|106|13|Cito obliti sunt operum eiuset non sustinuerunt consilium eius;
PS|106|14|et concupierunt concupiscentiam in desertoet tentaverunt Deum in inaquoso.
PS|106|15|Et dedit eis petitionem ipsorumet misit saturitatem in animas eorum.
PS|106|16|Et zelati sunt Moysen in castris,Aaron sanctum Domini.
PS|106|17|Aperta est terra et deglutivit Dathanet operuit super congregationem Abiram.
PS|106|18|Et exarsit ignis in synagoga eorum,flamma combussit peccatores.
PS|106|19|Et fecerunt vitulum in Horebet adoraverunt sculptile;
PS|106|20|et mutaverunt gloriam suamin similitudinem tauri comedentis fenum.
PS|106|21|Obliti sunt Deum, qui salvavit eos,qui fecit magnalia in Aegypto,
PS|106|22|mirabilia in terra Cham,terribilia in mari Rubro.
PS|106|23|Et dixit quia disperderet eos,nisi affuisset Moyses electus eius:stetit in confractione in conspectu eius,ut averteret iram eius, ne destrueret eos.
PS|106|24|Et pro nihilo habuerunt terram desiderabilem,non crediderunt verbo eius.
PS|106|25|Et murmuraverunt in tabernaculis suis,non exaudierunt vocem Domini.
PS|106|26|Et elevavit manum suam super eos,ut prosterneret eos in deserto
PS|106|27|et ut deiceret semen eorum in nationibuset dispergeret eos in regionibus.
PS|106|28|Et adhaeserunt Baalphegoret comederunt sacrificia mortuorum;
PS|106|29|et irritaverunt eum in adinventionibus suis,et irrupit in eos ruina.
PS|106|30|Et stetit Phinees et fecit iudicium,et cessavit quassatio,
PS|106|31|et reputatum est ei in iustitiamin generationem et generationem usque in sempiternum.
PS|106|32|Et irritaverunt eum ad aquas Meriba,et vexatus est Moyses propter eos,
PS|106|33|quia exacerbaverunt spiritum eius,et temere locutus est in labiis suis.
PS|106|34|Non disperdiderunt gentes,quas dixit Dominus illis.
PS|106|35|Et commixti sunt inter genteset didicerunt opera eorum.
PS|106|36|Et servierunt sculptilibus eorum,et factum est illis in scandalum.
PS|106|37|Et immolaverunt filios suoset filias suas daemoniis.
PS|106|38|Et effuderunt sanguinem innocentem,sanguinem filiorum suorum et filiarum suarum,quas sacrificaverunt sculptilibus Chanaan.Et infecta est terra in sanguinibus,
PS|106|39|et contaminati sunt in operibus suiset fornicati sunt in adinventionibus suis.
PS|106|40|Et exarsit ira Dominus in populum suumet abominatus est hereditatem suam
PS|106|41|et tradidit eos in manus gentium,et dominati sunt eorum, qui oderunt eos.
PS|106|42|Et tribulaverunt eos inimici eorum,et humiliati sunt sub manibus eorum.
PS|106|43|Saepe liberavit eos;ipsi autem exacerbaverunt eum in consilio suoet corruerunt in iniquitatibus suis.
PS|106|44|Et vidit tribulationem eorum,cum audivit clamorem eorum. -
PS|106|45|Et memor fuit testamenti suiet paenituit eum secundum multitudinem misericordiae suae.
PS|106|46|Et dedit eos in miserationesin conspectu omnium, qui captivos duxerant eos.
PS|106|47|Salvos nos fac, Domine Deus noster,et congrega nos de nationibus,ut confiteamur nomini sancto tuoet gloriemur in laude tua.
PS|106|48|Benedictus Dominus, Deus Israel, a saeculo et usque in saeculum.Et dicet omnis populus: "Fiat, fiat".
PS|107|1|ALLELUIA. Confitemini Domino, quoniam bonus, quoniam in saeculum misericordia eius.
PS|107|2|Dicant, qui redempti sunt a Domino,quos redemit de manu adversarii
PS|107|3|et de regionibus congregavit eos,a solis ortu et occasu,ab aquilone et mari.
PS|107|4|Erraverunt in solitudine, in inaquoso,viam civitatis habitationis non invenerunt.
PS|107|5|Esurientes et sitientes,anima eorum in ipsis defecit.
PS|107|6|Et clamaverunt ad Dominum, cum tribularentur,et de necessitatibus eorum eripuit eos.
PS|107|7|Et deduxit eos in viam rectam,ut irent in civitatem habitationis.
PS|107|8|Confiteantur Domino propter misericordiam eiuset mirabilia eius in filios hominum,
PS|107|9|quia satiavit animam sitientemet animam esurientem replevit bonis.
PS|107|10|Sedentes in tenebris et umbra mortis,vincti in mendicitate et ferro,
PS|107|11|quia exacerbaverunt eloquia Deiet consilium Altissimi spreverunt.
PS|107|12|Et humiliavit in laboribus cor eorum,infirmati sunt, nec fuit qui adiuvaret.
PS|107|13|Et clamaverunt ad Dominum, cum tribularentur,et de necessitatibus eorum liberavit eos.
PS|107|14|Et eduxit eos de tenebris et umbra mortiset vincula eorum dirupit.
PS|107|15|Confiteantur Domino propter misericordiam eiuset mirabilia eius in filios hominum,
PS|107|16|quia contrivit portas aereaset vectes ferreos confregit.
PS|107|17|Stulti facti sunt in via iniquitatis suaeet propter iniustitias suas afflicti sunt;
PS|107|18|omnem escam abominata est anima eorum,et appropinquaverunt usque ad portas mortis.
PS|107|19|Et clamaverunt ad Dominum, cum tribularentur,et de necessitatibus eorum liberavit eos.
PS|107|20|Misit verbum suum et sanavit eoset eripuit eos de interitionibus eorum.
PS|107|21|Confiteantur Domino propter misericordiam eiuset mirabilia eius in filios hominum;
PS|107|22|et sacrificent sacrificium laudiset annuntient opera eius in exsultatione.
PS|107|23|Qui descendunt mare in navibus,facientes operationem in aquis multis,
PS|107|24|ipsi viderunt opera Dominiet mirabilia eius in profundo.
PS|107|25|Dixit et excitavit spiritum procellae,et exaltati sunt fluctus eius.
PS|107|26|Ascendunt usque ad caeloset descendunt usque ad abyssos;anima eorum in malis tabescebat.
PS|107|27|Turbati sunt et moti sunt sicut ebrius,et omnis sapientia eorum devorata est.
PS|107|28|Et clamaverunt ad Dominum, cum tribularentur,et de necessitatibus eorum eduxit eos.
PS|107|29|Et statuit procellam eius in auram,et tacuerunt fluctus eius.
PS|107|30|Et laetati sunt, quia siluerunt,et deduxit eos in portum voluntatis eorum.
PS|107|31|Confiteantur Domino propter misericordiam eiuset mirabilia eius in filios hominum;
PS|107|32|et exaltent eum in ecclesia plebiset in conventu seniorum laudent eum.
PS|107|33|Posuit flumina in desertumet exitus aquarum in sitim,
PS|107|34|terram fructiferam in salsuginema malitia inhabitantium in ea.
PS|107|35|Posuit desertum in stagna aquarumet terram sine aqua in exitus aquarum.
PS|107|36|Et collocavit illic esurientes,et constituerunt civitatem habitationis.
PS|107|37|Et seminaverunt agros et plantaverunt vineas,et fecerunt fructum in proventum suum.
PS|107|38|Et benedixit eis, et multiplicati sunt nimis,et iumenta eorum non minoravit.
PS|107|39|Et pauci facti sunt et vexati sunta tribulatione malorum et dolore.
PS|107|40|Effudit contemptionem super principeset errare fecit eos in deserto invio.
PS|107|41|Et suscepit pauperem de inopiaet posuit sicut oves familias.
PS|107|42|Videbunt recti et laetabuntur,et omnis iniquitas oppilabit os suum.
PS|107|43|Quis sapiens, et custodiet haecet intelleget misericordias Domini?.
PS|108|1|Canticum. PSALMUS. David.
PS|108|2|Paratum cor meum, Deus,paratum cor meum,cantabo et psallam. Euge, gloria mea!
PS|108|3|Exsurge, psalterium et cithara,excitabo auroram.
PS|108|4|Confitebor tibi in populis, Domine,et psallam tibi in nationibus,
PS|108|5|quia magna est usque ad caelos misericordia tua,et usque ad nubes veritas tua.
PS|108|6|Exaltare super caelos, Deus,et super omnem terram gloria tua.
PS|108|7|Ut liberentur dilecti tui,salvum fac dextera tua et exaudi me.
PS|108|8|Deus locutus est in sancto suo: Exsultabo et dividam Sichimamet convallem Succoth dimetiar;
PS|108|9|meus est Galaad, et meus est Manasses,et Ephraim fortitudo capitis mei,Iuda sceptrum meum.
PS|108|10|Moab lebes lavacri mei;super Idumaeam extendam calceamentum meum,super Philistaeam vociferabor ".
PS|108|11|Quis deducet me in civitatem munitam?Quis deducet me usque in Idumaeam?.
PS|108|12|Nonne, Deus, qui reppulisti nos?Et non exibis, Deus, in virtutibus nostris?
PS|108|13|Da nobis auxilium de tribulatione,quia vana salus hominis.
PS|108|14|In Deo faciemus virtutem,et ipse conculcabit inimicos nostros.
PS|109|1|Magistro chori. David. PSALMUS.Deus laudis meae, ne tacueris,
PS|109|2|quia os peccatoris et os dolosi super me apertum est.Locuti sunt adversum me lingua dolosa
PS|109|3|et sermonibus odii circumdederunt meet expugnaverunt me gratis.
PS|109|4|Pro dilectione mea adversabantur mihi;ego autem orabam.
PS|109|5|Et posuerunt adversum me mala pro boniset odium pro dilectione mea.
PS|109|6|Constitue super eum peccatorem,et adversarius stet a dextris eius.
PS|109|7|Cum iudicatur, exeat condemnatus,et oratio eius fiat in peccatum.
PS|109|8|Fiant dies eius pauci,et ministerium eius accipiat alter.
PS|109|9|Fiant filii eius orphani,et uxor eius vidua.
PS|109|10|Instabiles vagentur filii eius et mendicentet eiciantur de ruinis suis. -
PS|109|11|Scrutetur fenerator omnem substantiam eius,et diripiant alieni labores eius.
PS|109|12|Non sit qui praebeat illi misericordiam,nec sit qui misereatur pupillis eius.
PS|109|13|Fiant nati eius in interitum,in generatione una deleatur nomen eorum.
PS|109|14|In memoriam redeat iniquitas patrum eius in conspectu Domini,et peccatum matris eius non deleatur.
PS|109|15|Fiant contra Dominum semper,et disperdat de terra memoriam eorum.
PS|109|16|Pro eo quod non est recordatus facere misericordiamet persecutus est hominem inopem et mendicumet compunctum corde, ut mortificaret.
PS|109|17|Et dilexit maledictionem: et veniat ei;et noluit benedictionem: et elongetur ab eo.
PS|109|18|Et induit maledictionem sicut vestimentum:et intret sicut aqua in interiora eius,et sicut oleum in ossa eius.
PS|109|19|Fiat ei sicut indumentum, quo operitur,et sicut zona, qua semper praecingitur.
PS|109|20|Haec retributio eorum, qui adversantur mihi apud Dominum,et qui loquuntur mala adversus animam meam.
PS|109|21|Et tu, Domine, Domine, fac mecum propter nomen tuum,quia suavis est misericordia tua;libera me,
PS|109|22|quia egenus et pauper ego sum,et cor meum vulneratum est intra me.
PS|109|23|Sicut umbra, cum declinat, pertransii,excussus sum sicut locustae.
PS|109|24|Genua mea infirmata sunt ieiunio,et caro mea contabuit absque oleo.
PS|109|25|Et ego factus sum opprobrium illis:viderunt me et moverunt capita sua.
PS|109|26|Adiuva me, Domine Deus meus,salvum me fac secundum misericordiam tuam.
PS|109|27|Et sciant quia manus tua haec:tu, Domine, hoc fecisti.
PS|109|28|Maledicant illi, et tu benedicas;qui insurgunt in me, confundantur,servus autem tuus laetabitur.
PS|109|29|Induantur, qui detrahunt mihi, pudoreet operiantur sicut diploide confusione sua.
PS|109|30|Confitebor Domino nimis in ore meoet in medio multorum laudabo eum,
PS|109|31|quia astitit a dextris pauperis,ut salvam faceret a iudicantibus animam eius.
PS|110|1|David. PSALMUS.Dixit Dominus Domino meo: " Sede a dextris meis,donec ponam inimicos tuos scabellum pedum tuorum ".
PS|110|2|Virgam potentiae tuae emittet Dominus ex Sion:dominare in medio inimicorum tuorum.
PS|110|3|Tecum principatus in die virtutis tuae,in splendoribus sanctis,ex utero ante luciferum genui te.
PS|110|4|Iuravit Dominus et non paenitebit eum: Tu es sacerdos in aeternum secundum ordinem Melchisedech ".
PS|110|5|Dominus a dextris tuis,conquassabit in die irae suae reges.
PS|110|6|Iudicabit in nationibus: cumulantur cadavera,conquassabit capita in terra spatiosa.
PS|110|7|De torrente in via bibet,propterea exaltabit caput.
PS|111|1|ALLELUIA.ALEPH. Confitebor Domino in toto corde meo,BETH. in consilio iustorum et congregatione.
PS|111|2|GHIMEL. Magna opera Domini,DALETH. exquirenda omnibus, qui cupiunt ea.
PS|111|3|HE. Decor et magnificentia opus eius,VAU. et iustitia eius manet in saeculum saeculi.
PS|111|4|ZAIN. Memoriam fecit mirabilium suorum,HETH. misericors et miserator Dominus.
PS|111|5|TETH. Escam dedit timentibus se;IOD. memor erit in saeculum testamenti sui.
PS|111|6|CAPH. Virtutem operum suorum annuntiavit populo suo,LAMED. ut det illis hereditatem gentium;
PS|111|7|MEM. opera manuum eius veritas et iudicium.NUN. Fidelia omnia mandata eius,
PS|111|8|SAMECH. confirmata in saeculum saeculi,AIN. facta in veritate et aequitate.
PS|111|9|PHE. Redemptionem misit populo suo,SADE. mandavit in aeternum testamentum suum.COPH. Sanctum et terribile nomen eius.
PS|111|10|RES. Initium sapientiae timor Domini,SIN. intellectus bonus omnibus facientibus ea;TAU. laudatio eius manet in saeculum saeculi.
PS|112|1|ALLELUIA.ALEPH. Beatus vir, qui timet Dominum,BETH. in mandatis eius cupit nimis.
PS|112|2|GHIMEL. Potens in terra erit semen eius,DALETH. generatio rectorum benedicetur.
PS|112|3|HE. Gloria et divitiae in domo eius,VAU. et iustitia eius manet in saeculum saeculi.
PS|112|4|ZAIN. Exortum est in tenebris lumen rectis,HETH. misericors et miserator et iustus.
PS|112|5|TETH. Iucundus homo, qui miseretur et commodat,IOD. disponet res suas in iudicio,
PS|112|6|CAPH. quia in aeternum non commovebitur.LAMED. In memoria aeterna erit iustus,
PS|112|7|MEM. ab auditione mala non timebit.NUN. Paratum cor eius, sperans in Domino,
PS|112|8|SAMECH. confirmatum est cor eius, non timebit,AIN. donec despiciat inimicos suos.
PS|112|9|PHE. Distribuit, dedit pauperibus;SADE. iustitia eius manet in saeculum saeculi,COPH. cornu eius exaltabitur in gloria.
PS|112|10|RES. Peccator videbit et irascetur,SIN. dentibus suis fremet et tabescet.TAU. Desiderium peccatorum peribit.
PS|113|1|ALLELUIA.Laudate, pueri Domini,laudate nomen Domini.
PS|113|2|Sit nomen Domini benedictumex hoc nunc et usque in saeculum.
PS|113|3|A solis ortu usque ad occasumlaudabile nomen Domini.
PS|113|4|Excelsus super omnes gentes Dominus,super caelos gloria eius.
PS|113|5|Quis sicut Dominus Deus noster,qui in altis habitat
PS|113|6|et se inclinat, ut respiciatin caelum et in terram?
PS|113|7|Suscitans de terra inopem,de stercore erigens pauperem,
PS|113|8|ut collocet eum cum principibus,cum principibus populi sui.
PS|113|9|Qui habitare facit sterilem in domo,matrem filiorum laetantem.
PS|114|1|ALLELUIA.In exitu Israel de Aegypto,domus Iacob de populo barbaro,
PS|114|2|factus est Iuda sanctuarium eius,Israel potestas eius.
PS|114|3|Mare vidit et fugit,Iordanis conversus est retrorsum;
PS|114|4|montes saltaverunt ut arietes,et colles sicut agni ovium. -
PS|114|5|Quid est tibi, mare, quod fugisti?Et tu, Iordanis, quia conversus es retrorsum?
PS|114|6|Montes, quod saltastis sicut arietes,et colles, sicut agni ovium?
PS|114|7|A facie Domini contremisce, terra,a facie Dei Iacob,
PS|114|8|qui convertit petram in stagna aquarumet silicem in fontes aquarum.
PS|115|1|Non nobis, Domine, non nobis,sed nomini tuo da gloriamsuper misericordia tua et veritate tua.
PS|115|2|Quare dicent gentes: Ubi est Deus eorum? ".
PS|115|3|Deus autem noster in caelo;omnia, quaecumque voluit, fecit.
PS|115|4|Simulacra gentium argentum et aurum,opera manuum hominum.
PS|115|5|Os habent et non loquentur,oculos habent et non videbunt.
PS|115|6|Aures habent et non audient,nares habent et non odorabunt.
PS|115|7|Manus habent et non palpabunt,pedes habent et non ambulabunt;non clamabunt in gutture suo.
PS|115|8|Similes illis erunt, qui faciunt ea,et omnes, qui confidunt in eis.
PS|115|9|Domus Israel speravit in Domino:adiutorium eorum et scutum eorum est.
PS|115|10|Domus Aaron speravit in Domino:adiutorium eorum et scutum eorum est.
PS|115|11|Qui timent Dominum, speraverunt in Domino:adiutorium eorum et scutum eorum est.
PS|115|12|Dominus memor fuit nostriet benedicet nobis:benedicet domui Israel,benedicet domui Aaron,
PS|115|13|benedicet omnibus, qui timent Dominum,pusillis cum maioribus.
PS|115|14|Adiciat Dominus super vos,super vos et super filios vestros.
PS|115|15|Benedicti vos a Domino,qui fecit caelum et terram.
PS|115|16|Caeli, caeli sunt Domino,terram autem dedit filiis hominum.
PS|115|17|Non mortui laudabunt te, Domine,neque omnes, qui descendunt in silentium,
PS|115|18|sed nos, qui vivimus, benedicimus Dominoex hoc nunc et usque in saeculum.
PS|116|1|ALLELUIA.Dilexi, quoniam exaudit Dominusvocem deprecationis meae.
PS|116|2|Quia inclinavit aurem suam mihi,cum in diebus meis invocabam.
PS|116|3|Circumdederunt me funes mortis,et angustiae inferni invenerunt me. Tribulationem et dolorem inveni
PS|116|4|et nomen Domini invocabam: O Domine, libera animam meam ".
PS|116|5|Misericors Dominus et iustus,et Deus noster miseretur.
PS|116|6|Custodiens parvulos Dominus;humiliatus sum, et salvum me faciet.
PS|116|7|Convertere, anima mea, in requiem tuam,quia Dominus benefecit tibi;
PS|116|8|quia eripuit animam meam de morte,oculos meos a lacrimis,pedes meos a lapsu.
PS|116|9|Ambulabo coram Dominoin regione vivorum. -
PS|116|10|Credidi, etiam cum locutus sum: " Ego humiliatus sum nimis ".
PS|116|11|Ego dixi in trepidatione mea: " Omnis homo mendax ".
PS|116|12|Quid retribuam Dominopro omnibus, quae retribuit mihi?
PS|116|13|Calicem salutaris accipiamet nomen Domini invocabo.
PS|116|14|Vota mea Domino reddamcoram omni populo eius.
PS|116|15|Pretiosa in conspectu Dominimors sanctorum eius.
PS|116|16|O Domine, ego servus tuus,ego servus tuus et filius ancillae tuae.Dirupisti vincula mea:
PS|116|17|tibi sacrificabo hostiam laudiset nomen Domini invocabo.
PS|116|18|Vota mea Domino reddamcoram omni populo eius
PS|116|19|in atriis domus Domini,in medio tui, Ierusalem.
PS|117|1|ALLELUIA.Laudate Dominum, omnes gentes;collaudate eum, omnes populi.
PS|117|2|Quoniam confirmata est super nos misericordia eius,et veritas Domini manet in aeternum.
PS|118|1|ALLELUIA.Confitemini Domino, quoniam bonus,quoniam in saeculum misericordia eius.
PS|118|2|Dicat nunc Israel, quoniam bonus,quoniam in saeculum misericordia eius.
PS|118|3|Dicat nunc domus Aaron,quoniam in saeculum misericordia eius.
PS|118|4|Dicant nunc, qui timent Dominum,quoniam in saeculum misericordia eius.
PS|118|5|De tribulatione invocavi Dominum,et exaudivit me educens in latitudinem Dominus.
PS|118|6|Dominus mecum,non timebo, quid faciat mihi homo.
PS|118|7|Dominus mecum adiutor meus,et ego despiciam inimicos meos.
PS|118|8|Bonum est confugere ad Dominumquam confidere in homine.
PS|118|9|Bonum est confugere ad Dominumquam confidere in principibus.
PS|118|10|Omnes gentes circuierunt me,et in nomine Domini excidi eos.
PS|118|11|Circumdantes circumdederunt me,et in nomine Domini excidi eos.
PS|118|12|Circumdederunt me sicut apeset exarserunt sicut ignis in spinis,et in nomine Domini excidi eos.
PS|118|13|Impellentes impulerunt me, ut caderem,et Dominus adiuvit me.
PS|118|14|Fortitudo mea et laus mea Dominuset factus est mihi in salutem.
PS|118|15|Vox iubilationis et salutisin tabernaculis iustorum: Dextera Domini fecit virtutem!
PS|118|16|Dextera Domini exaltata est;dextera Domini fecit virtutem! ".
PS|118|17|Non moriar, sed vivamet narrabo opera Domini.
PS|118|18|Castigans castigavit me Dominuset morti non tradidit me.
PS|118|19|Aperite mihi portas iustitiae;ingressus in eas confitebor Domino.
PS|118|20|Haec porta Domini;iusti intrabunt in eam. -
PS|118|21|Confitebor tibi, quoniam exaudisti meet factus es mihi in salutem.
PS|118|22|Lapidem quem reprobaverunt aedificantes,hic factus est in caput anguli;
PS|118|23|a Domino factum est istudet est mirabile in oculis nostris.
PS|118|24|Haec est dies, quam fecit Dominus:exsultemus et laetemur in ea.
PS|118|25|O Domine, salvum me fac;o Domine, da prosperitatem!
PS|118|26|Benedictus, qui venit in nomine Domini.Benedicimus vobis de domo Domini.
PS|118|27|Deus Dominus et illuxit nobis.Instruite sollemnitatem in ramis condensisusque ad cornua altaris.
PS|118|28|Deus meus es tu, et confitebor tibi,Deus meus, et exaltabo te.
PS|118|29|Confitemini Domino, quoniam bonus,quoniam in saeculum misericordia eius.
PS|119|1|ALLELUIA.ALEPH. Beati immaculati in via,qui ambulant in lege Domini.
PS|119|2|Beati, qui servant testimonia eius,in toto corde exquirunt eum.
PS|119|3|Non enim operati sunt iniquitatem,in viis eius ambulaverunt.
PS|119|4|Tu mandastimandata tua custodiri nimis.
PS|119|5|Utinam dirigantur viae meaead custodiendas iustificationes tuas!
PS|119|6|Tunc non confundar,cum perspexero in omnibus praeceptis tuis.
PS|119|7|Confitebor tibi in directione cordis,in eo quod didici iudicia iustitiae tuae.
PS|119|8|Iustificationes tuas custodiam,non me derelinquas usquequaque.
PS|119|9|BETH. In quo mundabit adulescentior viam suam?In custodiendo sermones tuos.
PS|119|10|In toto corde meo exquisivi te;ne errare me facias a praeceptis tuis.
PS|119|11|In corde meo abscondi eloquia tua,ut non peccem tibi.
PS|119|12|Benedictus es, Domine;doce me iustificationes tuas.
PS|119|13|In labiis meisnumeravi omnia iudicia oris tui.
PS|119|14|In via testimoniorum tuorum delectatus sumsicut in omnibus divitiis.
PS|119|15|In mandatis tuis exerceboret considerabo vias tuas.
PS|119|16|In iustificationibus tuis delectabor,non obliviscar sermonem tuum.
PS|119|17|GHIMEL. Benefac servo tuo, et vivamet custodiam sermonem tuum.
PS|119|18|Revela oculos meos,et considerabo mirabilia de lege tua.
PS|119|19|Incola ego sum in terra,non abscondas a me praecepta tua.
PS|119|20|Defecit anima mea in desiderando iudicia tuain omni tempore.
PS|119|21|Increpasti superbos;maledicti, qui errant a praeceptis tuis.
PS|119|22|Aufer a me opprobrium et contemptum,quia testimonia tua servavi.
PS|119|23|Etsi principes sedent et adversum me loquuntur,servus tamen tuus exercetur in iustificationibus tuis.
PS|119|24|Nam et testimonia tua delectatio mea,et consilium meum iustificationes tuae.
PS|119|25|DALETH. Adhaesit pulveri anima mea;vivifica me secundum verbum tuum.
PS|119|26|Vias meas enuntiavi, et exaudisti me;doce me iustificationes tuas.
PS|119|27|Viam mandatorum tuorum fac me intellegere,et exercebor in mirabilibus tuis.
PS|119|28|Lacrimata est anima mea prae maerore;erige me secundum verbum tuum.
PS|119|29|Viam mendacii averte a meet legem tuam da mihi benigne.
PS|119|30|Viam veritatis elegi,iudicia tua proposui mihi.
PS|119|31|Adhaesi testimoniis tuis, Domine;noli me confundere.
PS|119|32|Viam mandatorum tuorum curram,quia dilatasti cor meum.
PS|119|33|HE. Legem pone mihi, Domine, viam iustificationum tuarum,et servabo eam semper.
PS|119|34|Da mihi intellectum, et servabo legem tuamet custodiam illam in toto corde meo.
PS|119|35|Deduc me in semitam praeceptorum tuorum,quia ipsam volui.
PS|119|36|Inclina cor meum in testimonia tuaet non in avaritiam.
PS|119|37|Averte oculos meos, ne videant vanitatem;in via tua vivifica me.
PS|119|38|Suscita servo tuo eloquium tuum,quod est ad timorem tuum.
PS|119|39|Amove opprobrium meum, quod suspicatus sum,quia iudicia tua iucunda.
PS|119|40|Ecce concupivi mandata tua;in iustitia tua vivifica me.
PS|119|41|VAU. Et veniat super me misericordia tua, Domine,salutare tuum secundum eloquium tuum.
PS|119|42|Et respondebo exprobrantibus mihi verbum,quia speravi in sermonibus tuis.
PS|119|43|Et ne auferas de ore meo verbum veritatis usquequaque,quia in iudiciis tuis supersperavi.
PS|119|44|Et custodiam legem tuam semper,in saeculum et in saeculum saeculi.
PS|119|45|Et ambulabo in latitudine,quia mandata tua exquisivi.
PS|119|46|Et loquar de testimoniis tuis in conspectu regumet non confundar.
PS|119|47|Et delectabor in praeceptis tuis,quae dilexi.
PS|119|48|Et levabo manus meas ad praecepta tua, quae dilexi;et exercebor in iustificationibus tuis. -
PS|119|49|ZAIN. Memor esto verbi tui servo tuo,in quo mihi spem dedisti.
PS|119|50|Hoc me consolatum est in humiliatione mea,quia eloquium tuum vivificavit me.
PS|119|51|Superbi deriserunt me vehementer;a lege autem tua non declinavi.
PS|119|52|Memor fui iudiciorum tuorum a saeculo, Domine,et consolatus sum.
PS|119|53|Indignatio tenuit mepropter peccatores derelinquentes legem tuam.
PS|119|54|Cantica factae sunt mihi iustificationes tuaein loco peregrinationis meae.
PS|119|55|Memor fui nocte nominis tui, Domine,et custodiam legem tuam.
PS|119|56|Hoc factum est mihi,quia mandata tua servavi.
PS|119|57|HETH. Portio mea Dominus:dixi custodire verba tua.
PS|119|58|Deprecatus sum faciem tuam in toto corde meo;miserere mei secundum eloquium tuum.
PS|119|59|Cogitavi vias measet converti pedes meos in testimonia tua.
PS|119|60|Festinavi et non sum moratus,ut custodiam praecepta tua.
PS|119|61|Funes peccatorum circumplexi sunt me,et legem tuam non sum oblitus.
PS|119|62|Media nocte surgebam ad confitendum tibisuper iudicia iustitiae tuae.
PS|119|63|Particeps ego sum omnium timentium teet custodientium mandata tua.
PS|119|64|Misericordia tua, Domine, plena est terra;iustificationes tuas doce me.
PS|119|65|TETH. Bonitatem fecisti cum servo tuo, Domine,secundum verbum tuum.
PS|119|66|Bonitatem et prudentiam et scientiam doce me,quia praeceptis tuis credidi.
PS|119|67|Priusquam humiliarer ego erravi;nunc autem eloquium tuum custodiam.
PS|119|68|Bonus es tu et benefaciens,doce me iustificationes tuas.
PS|119|69|Excogitaverunt contra me dolosa superbi,ego autem in toto corde meo servabo mandata tua.
PS|119|70|Incrassatum est sicut adeps cor eorum,ego vero in lege tua delectatus sum.
PS|119|71|Bonum mihi quia humiliatus sum,ut discam iustificationes tuas.
PS|119|72|Bonum mihi lex oris tuisuper milia auri et argenti.
PS|119|73|IOD. Manus tuae fecerunt me et plasmaverunt me;da mihi intellectum, et discam praecepta tua.
PS|119|74|Qui timent te, videbunt me et laetabuntur,quia in verba tua supersperavi.
PS|119|75|Cognovi, Domine, quia aequitas iudicia tua,et in veritate humiliasti me.
PS|119|76|Fiat misericordia tua, ut consoletur me,secundum eloquium tuum servo tuo.
PS|119|77|Veniant mihi miserationes tuae, et vivam,quia lex tua delectatio mea est.
PS|119|78|Confundantur superbi, quoniam dolose incurvaverunt me,ego autem exercebor in mandatis tuis.
PS|119|79|Convertantur mihi timentes te,et qui noverunt testimonia tua.
PS|119|80|Fiat cor meum immaculatum in iustificationibus tuis,ut non confundar.
PS|119|81|CAPH. Defecit in salutare tuum anima mea,et in verbum tuum supersperavi.
PS|119|82|Defecerunt oculi mei in eloquium tuum,dicentes: " Quando consolaberis me? ".
PS|119|83|Quia factus sum sicut uter in fumo;iustificationes tuas non sum oblitus.
PS|119|84|Quot sunt dies servi tui?Quando facies de persequentibus me iudicium?
PS|119|85|Foderunt mihi foveas superbi,qui non sunt secundum legem tuam.
PS|119|86|Omnia praecepta tua veritas;dolose persecuti sunt me; adiuva me.
PS|119|87|Paulo minus consummaverunt me in terra,ego autem non dereliqui mandata tua.
PS|119|88|Secundum misericordiam tuam vivifica me,et custodiam testimonia oris tui. -
PS|119|89|LAMED. In aeternum, Domine,verbum tuum constitutum est in caelo.
PS|119|90|In generationem et generationem veritas tua;firmasti terram, et permanet.
PS|119|91|Secundum iudicia tua permanent hodie,quoniam omnia serviunt tibi.
PS|119|92|Nisi quod lex tua delectatio mea est,tunc forte periissem in humilia tione mea.
PS|119|93|In aeternum non obliviscar man data tua,quia in ipsis vivificasti me.
PS|119|94|Tuus sum ego: salvum me fac,quoniam mandata tua exqui sivi.
PS|119|95|Me exspectaverunt peccatores, ut perderent me;testimonia tua intellexi.
PS|119|96|Omni consummationi vidi finem,latum praeceptum tuum nimis.
PS|119|97|MEM. Quomodo dilexi legem tuam, Domine;tota die meditatio mea est.
PS|119|98|Super inimicos meos sapientem me fecit praeceptum tuum,quia in aeternum mihi est.
PS|119|99|Super omnes docentes me prudens factus sum,quia testimonia tua meditatio mea est.
PS|119|100|Super senes intellexi,quia mandata tua servavi.
PS|119|101|Ab omni via mala prohibui pedes meos,ut custodiam verba tua.
PS|119|102|A iudiciis tuis non declinavi,quia tu legem posuisti mihi.
PS|119|103|Quam dulcia faucibus meis eloquia tua,super mel ori meo.
PS|119|104|A mandatis tuis intellexi;propterea odivi omnem viam mendacii.
PS|119|105|NUN. Lucerna pedibus meis verbum tuumet lumen semitis meis.
PS|119|106|Iuravi et statuicustodire iudicia iustitiae tuae.
PS|119|107|Humiliatus sum usquequaque, Domine;vivifica me secundum verbum tuum.
PS|119|108|Voluntaria oris mei beneplacita sint, Domine,et iudicia tua doce me.
PS|119|109|Anima mea in manibus meis semper,et legem tuam non sum oblitus.
PS|119|110|Posuerunt peccatores laqueum mihi,et de mandatis tuis non erravi.
PS|119|111|Hereditas mea testimonia tua in aeternum,quia exsultatio cordis mei sunt.
PS|119|112|Inclinavi cor meum ad faciendas iustificationes tuasin aeternum, in finem.
PS|119|113|SAMECH. Duplices corde odio habuiet legem tuam dilexi.
PS|119|114|Tegmen et scutum meum es tu,et in verbum tuum supersperavi.
PS|119|115|Declinate a me, maligni,et servabo praecepta Dei mei.
PS|119|116|Suscipe me secundum eloquium tuum, et vivam;et non confundas me ab exspectatione mea.
PS|119|117|Sustenta me, et salvus eroet delectabor in iustificationibus tuis semper.
PS|119|118|Sprevisti omnes discedentes a iustificationibus tuis,quia mendacium cogitatio eorum.
PS|119|119|Quasi scoriam delesti omnes peccatores terrae;ideo dilexi testimonia tua.
PS|119|120|Horruit a timore tuo caro mea;a iudiciis enim tuis timui.
PS|119|121|AIN. Feci iudicium et iustitiam;non tradas me calumniantibus me.
PS|119|122|Sponde pro servo tuo in bonum;non calumnientur me superbi.
PS|119|123|Oculi mei defecerunt in desiderio salutaris tuiet eloquii iustitiae tuae.
PS|119|124|Fac cum servo tuo secundum misericordiam tuamet iustificationes tuas doce me.
PS|119|125|Servus tuus sum ego;da mihi intellectum, ut sciam testimonia tua.
PS|119|126|Tempus faciendi Domino;dissipaverunt legem tuam.
PS|119|127|Ideo dilexi praecepta tuasuper aurum et obryzum.
PS|119|128|Propterea ad omnia mandata tua dirigebar,omnem viam mendacii odio habui. -
PS|119|129|PHE. Mirabilia testimonia tua,ideo servavit ea anima mea.
PS|119|130|Declaratio sermonum tuorum illuminatet intellectum dat parvulis.
PS|119|131|Os meum aperui et attraxi spiritum,quia praecepta tua desiderabam.
PS|119|132|Convertere in me et miserere meisecundum iudicium tuum cum diligentibus nomen tuum.
PS|119|133|Gressus meos dirige secundum eloquium tuum,et non dominetur mei omnis iniquitas.
PS|119|134|Redime me a calumniis hominum,ut custodiam mandata tua.
PS|119|135|Faciem tuam illumina super servum tuumet doce me iustificationes tuas.
PS|119|136|Rivulos aquarum deduxerunt oculi mei,quia non custodierunt legem tuam.
PS|119|137|SADE. Iustus es, Domine,et rectum iudicium tuum.
PS|119|138|Mandasti in iustitia testimonia tuaet in veritate nimis.
PS|119|139|Consumpsit me zelus meus,quia obliti sunt verba tua inimici mei.
PS|119|140|Ignitum eloquium tuum vehementer,et servus tuus dilexit illud.
PS|119|141|Adulescentulus sum ego et contemptus;mandata tua non sum oblitus.
PS|119|142|Iustitia tua iustitia in aeternum,et lex tua veritas.
PS|119|143|Tribulatio et angustia invenerunt me;praecepta tua delectatio mea est.
PS|119|144|Iustitia testimonia tua in aeternum;intellectum da mihi, et vivam.
PS|119|145|COPH. Clamavi in toto corde, exaudi me, Domine;iustificationes tuas servabo.
PS|119|146|Clamavi ad te, salvum me fac,ut custodiam testimonia tua.
PS|119|147|Praeveni diluculo et clamavi,in verba tua supersperavi.
PS|119|148|Praevenerunt oculi mei vigilias,ut meditarer eloquia tua.
PS|119|149|Vocem meam audi secundum misericordiam tuam, Domine,secundum iudicium tuum vivifica me.
PS|119|150|Appropinquaverunt persequentes me in malitia,a lege autem tua longe facti sunt.
PS|119|151|Prope es tu, Domine,et omnia praecepta tua veritas.
PS|119|152|Ab initio cognovi de testimoniis tuis,quia in aeternum fundasti ea.
PS|119|153|RES. Vide humiliationem meam et eripe me,quia legem tuam non sum oblitus.
PS|119|154|Iudica causam meam et redime me;propter eloquium tuum vivifica me.
PS|119|155|Longe a peccatoribus salus,quia iustificationes tuas non exquisierunt.
PS|119|156|Misericordiae tuae multae, Domine;secundum iudicia tua vivifica me.
PS|119|157|Multi, qui persequuntur me et tribulant me;a testimoniis tuis non declinavi.
PS|119|158|Vidi praevaricantes, et taeduit me,quia eloquia tua non custodierunt.
PS|119|159|Vide quoniam mandata tua dilexi, Domine;secundum misericordiam tuam vivifica me.
PS|119|160|Principium verborum tuorum veritas,in aeternum omnia iudicia iustitiae tuae.
PS|119|161|SIN. Principes persecuti sunt me gratis,et a verbis tuis formidavit cor meum.
PS|119|162|Laetabor ego super eloquia tua,sicut qui invenit spolia multa.
PS|119|163|Mendacium odio habui et abominatus sum;legem autem tuam dilexi.
PS|119|164|Septies in die laudem dixi tibisuper iudicia iustitiae tuae.
PS|119|165|Pax multa diligentibus legem tuam, et non est illis scandalum.
PS|119|166|Exspectabam salutare tuum, Domine,et praecepta tua feci.
PS|119|167|Custodivit anima mea testimonia tua,et dilexi ea vehementer.
PS|119|168|Servavi mandata tua et testimonia tua,quia omnes viae meae in conspectu tuo.
PS|119|169|TAU. Appropinquet deprecatio mea in conspectu tuo, Domine;iuxta verbum tuum da mihi intellectum.
PS|119|170|Intret postulatio mea in conspectu tuo;secundum eloquium tuum libera me.
PS|119|171|Eructabunt labia mea hymnum,cum docueris me iustificationes tuas.
PS|119|172|Cantet lingua mea eloquium tuum,quia omnia praecepta tua iustitia.
PS|119|173|Fiat manus tua, ut adiuvet me,quoniam mandata tua elegi.
PS|119|174|Concupivi salutare tuum, Domine,et lex tua delectatio mea est.
PS|119|175|Vivet anima mea et laudabit te,et iudicia tua adiuvabunt me.
PS|119|176|Erravi sicut ovis, quae periit;quaere servum tuum, quia praecepta tua non sum oblitus.
PS|120|1|Canticum ascensionum.Ad Dominum, cum tribularer, clamavi,et exaudivit me.
PS|120|2|Domine, libera animam meam a labiis mendacii,a lingua dolosa.
PS|120|3|Quid detur tibi aut quid apponatur tibi,lingua dolosa?
PS|120|4|Sagittae potentis acutaecum carbonibus iuniperorum.
PS|120|5|Heu mihi, quia peregrinatus sum in Mosoch,habitavi ad tabernacula Cedar!
PS|120|6|Multum incola fuit anima meacum his, qui oderunt pacem.
PS|120|7|Ego eram pacificus;cum loquebar, illi impugnabant me.
PS|121|1|Canticum ascensionum.Levabo oculos meos in montes:unde veniet auxilium mihi?
PS|121|2|Auxilium meum a Domino,qui fecit caelum et terram.
PS|121|3|Non dabit in commotionem pedem tuumneque dormitabit, qui custodit te.
PS|121|4|Ecce non dormitabit neque dormiet,qui custodit Israel.
PS|121|5|Dominus custodit te,Dominus umbraculum tuumad manum dexteram tuam.
PS|121|6|Per diem sol non percutiet te,neque luna per noctem.
PS|121|7|Dominus custodiet te ab omni malo;custodiet animam tuam Dominus.
PS|121|8|Dominus custodiet introitum tuum et exitum tuumex hoc nunc et usque in saeculum.
PS|122|1|Canticum ascensionum. David.Laetatus sum in eo, quod dixerunt mihi: In domum Domini ibimus ".
PS|122|2|Stantes iam sunt pedes nostriin portis tuis, Ierusalem.
PS|122|3|Ierusalem, quae aedificata est ut civitas,sibi compacta in idipsum.
PS|122|4|Illuc enim ascenderunt tribus, tribus Domini,testimonium Israel, ad confitendum nomini Domini.
PS|122|5|Quia illic sederunt sedes ad iudicium,sedes domus David.
PS|122|6|Rogate, quae ad pacem sunt Ierusalem: Securi sint diligentes te!
PS|122|7|Fiat pax in muris tuis,et securitas in turribus tuis! ".
PS|122|8|Propter fratres meos et proximos meosloquar: " Pax in te! ".
PS|122|9|Propter domum Domini Dei nostriexquiram bona tibi.
PS|123|1|Canticum ascensionum.Ad te levavi oculos meos,qui habitas in caelis.
PS|123|2|Ecce sicut oculi servorum ad manus dominorum suorum,sicut oculi ancillae ad manus dominae suae,ita oculi nostri ad Dominum Deum nostrum,donec misereatur nostri.
PS|123|3|Miserere nostri, Domine, miserere nostri,quia multum repleti sumus despectione;
PS|123|4|quia multum repleta est anima nostraderisione abundantium et despectione superborum.
PS|124|1|Canticum ascensionum. David.Nisi quia Dominus erat in nobis,dicat nunc Israel,
PS|124|2|nisi quia Dominus erat in nobis,cum exsurgerent homines in nos:
PS|124|3|forte vivos deglutissent nos,cum irasceretur furor eorum in nos.
PS|124|4|Forsitan aqua absorbuisset nos,torrens pertransisset animam nostram;
PS|124|5|forsitan pertransissent animam nostramaquae intumescentes.
PS|124|6|Benedictus Dominus,qui non dedit nos in direptionem dentibus eorum.
PS|124|7|Anima nostra sicut passer erepta estde laqueo venantium:laqueus contritus est,et nos erepti sumus.
PS|124|8|Adiutorium nostrum in nomine Domini,qui fecit caelum et terram.
PS|125|1|Canticum ascensionum.Qui confidunt in Domino, sicut mons Sion:non commovebitur, in aeternum manet.
PS|125|2|Ierusalem, montes in circuitu eius,et Dominus in circuitu populi suiex hoc nunc et usque in saeculum.
PS|125|3|Quia non requiescet virga iniquitatis super sortem iustorum,ut non extendant iusti ad iniquitatem manus suas.
PS|125|4|Benefac, Domine, boniset rectis corde.
PS|125|5|Declinantes autem per vias pravasadducet Dominus cum operantibus iniquitatem.Pax super Israel!
PS|126|1|Canticum ascensionum.In convertendo Dominus captivitatem Sion,facti sumus quasi somniantes.
PS|126|2|Tunc repletum est gaudio os nostrum,et lingua nostra exsultatione.Tunc dicebant inter gentes: Magnificavit Dominus facere cum eis ".
PS|126|3|Magnificavit Dominus facere nobiscum;facti sumus laetantes.
PS|126|4|Converte, Domine, captivitatem nostram,sicut torrentes in austro.
PS|126|5|Qui seminant in lacrimis,in exsultatione metent.
PS|126|6|Euntes ibant et flebantsemen spargendum portantes;venientes autem venient in exsultationeportantes manipulos suos.
PS|127|1|Canticum ascensionum. Salomonis.Nisi Dominus aedificaverit domum,in vanum laborant, qui aedificant eam.Nisi Dominus custodierit civitatem,frustra vigilat, qui custodit eam.
PS|127|2|Vanum est vobis ante lucem surgere et sero quiescere,qui manducatis panem laboris,quia dabit dilectis suis somnum.
PS|127|3|Ecce hereditas Domini filii,merces fructus ventris.
PS|127|4|Sicut sagittae in manu potentis,ita filii iuventutis.
PS|127|5|Beatus vir, qui implevit pharetram suam ex ipsis:non confundetur, cum loquetur inimicis suis in porta.
PS|128|1|Canticum ascensionum.Beatus omnis, qui timet Dominum,qui ambulat in viis eius.
PS|128|2|Labores manuum tuarum manducabis,beatus es, et bene tibi erit.
PS|128|3|Uxor tua sicut vitis fructiferain lateribus domus tuae;filii tui sicut novellae olivarumin circuitu mensae tuae.
PS|128|4|Ecce sic benedicetur homo,qui timet Dominum.
PS|128|5|Benedicat tibi Dominus ex Sion,et videas bona Ierusalemomnibus diebus vitae tuae;
PS|128|6|et videas filios filiorum tuorum.Pax super Israel!
PS|129|1|Canticum ascensionum.Saepe expugnaverunt me a iuventute mea,dicat nunc Israel,
PS|129|2|saepe expugnaverunt me a iuventute mea,etenim non potuerunt adversum me.
PS|129|3|Supra dorsum meum araverunt aratores,prolongaverunt sulcos suos.
PS|129|4|Dominus autem iustusconcidit cervices peccatorum.
PS|129|5|Confundantur et convertantur retrorsumomnes, qui oderunt Sion.
PS|129|6|Fiant sicut fenum tectorum,quod, priusquam evellatur, exaruit;
PS|129|7|de quo non implevit manum suam, qui metit,et sinum suum, qui manipulos colligit.
PS|129|8|Et non dixerunt, qui praeteribant: Benedictio Domini super vos,benedicimus vobis in nomine Domini ".
PS|130|1|Canticum ascensionum.De profundis clamavi ad te, Domine;
PS|130|2|Domine, exaudi vocem meam.Fiant aures tuae intendentesin vocem deprecationis meae.
PS|130|3|Si iniquitates observaveris, Domine,Domine, quis sustinebit?
PS|130|4|Quia apud te propitiatio est,ut timeamus te.
PS|130|5|Sustinui te, Domine,sustinuit anima mea in verbo eius;speravit
PS|130|6|anima mea in Dominomagis quam custodes auroram.Magis quam custodes auroram
PS|130|7|speret Israel in Domino,quia apud Dominum misericordia,et copiosa apud eum redemptio.
PS|130|8|Et ipse redimet Israelex omnibus iniquitatibus eius.
PS|131|1|Canticum ascensionum. David.Domine, non est exaltatum cor meum,neque elati sunt oculi mei,neque ambulavi in magnisneque in mirabilibus super me.
PS|131|2|Vere pacatam et quietamfeci animam meam;sicut ablactatus in sinu matris suae,sicut ablactatus, ita in me est anima mea.
PS|131|3|Speret Israel in Dominoex hoc nunc et usque in saeculum.
PS|132|1|Canticum ascensionum.Memento, Domine, Davidet omnis mansuetudinis eius,
PS|132|2|quia iuravit Domino,votum vovit Potenti Iacob:
PS|132|3|" Non introibo in tabernaculum domus meae,non ascendam in lectum strati mei,
PS|132|4|non dabo somnum oculis meiset palpebris meis dormitationem,
PS|132|5|donec inveniam locum Domino,tabernaculum Potenti Iacob ".
PS|132|6|Ecce audivimus eam esse in Ephratha,invenimus eam in campis Iaar.
PS|132|7|Ingrediamur in tabernaculum eius,adoremus ad scabellum pedum eius. -
PS|132|8|Surge, Domine, in requiem tuam,tu et arca fortitudinis tuae.
PS|132|9|Sacerdotes tui induantur iustitiam,et sancti tui exsultent.
PS|132|10|Propter David servum tuumnon avertas faciem christi tui.
PS|132|11|Iuravit Dominus David veritatemet non recedet ab ea: De fructu ventris tuiponam super sedem tuam.
PS|132|12|Si custodierint filii tui testamentum meumet testimonia mea, quae docebo eos,filii eorum usque in saeculumsedebunt super sedem tuam ".
PS|132|13|Quoniam elegit Dominus Sion,desideravit eam in habitationem sibi:
PS|132|14|" Haec requies mea in saeculum saeculi;hic habitabo, quoniam desideravi eam.
PS|132|15|Cibaria eius benedicens benedicam,pauperes eius saturabo panibus.
PS|132|16|Sacerdotes eius induam salutari,et sancti eius exsultatione exsultabunt.
PS|132|17|Illic germinare faciam cornu David,parabo lucernam christo meo.
PS|132|18|Inimicos eius induam confusione,super ipsum autem efflorebit diadema eius ".
PS|133|1|Canticum ascensionum. David.Ecce quam bonum et quam iucundumhabitare fratres in unum:
PS|133|2|sicut unguentum optimum in capite,quod descendit in barbam, barbam Aaron,quod descendit in oram vestimenti eius;
PS|133|3|sicut ros Hermon, qui descendit in montes Sion,quoniam illic mandavit Dominus benedictionem,vitam usque in saeculum.
PS|134|1|Canticum ascensionum.Ecce benedicite Dominum,omnes servi Domini,qui statis in domo Domini per noctes.
PS|134|2|Extollite manus vestras ad sanctuariumet benedicite Dominum.
PS|134|3|Benedicat te Dominus ex Sion,qui fecit caelum et terram.
PS|135|1|ALLELUIA.Laudate nomen Domini,laudate, servi Domini,
PS|135|2|qui statis in domo Domini,in atriis domus Dei nostri.
PS|135|3|Laudate Dominum, quia bonus Dominus;psallite nomini eius, quoniam suave.
PS|135|4|Quoniam Iacob elegit sibi Dominus,Israel in peculium sibi.
PS|135|5|Quia ego cognovi quod magnus est Dominus,et Deus noster prae omnibus diis.
PS|135|6|Omnia, quaecumque voluit,Dominus fecit in caelo et in terra,in mari et in omnibus abyssis.
PS|135|7|Adducens nubes ab extremo terrae,fulgura in pluviam facit,producit ventos de thesauris suis.
PS|135|8|Qui percussit primogenita Aegyptiab homine usque ad pecus.
PS|135|9|Misit signa et prodigia in medio tui, Aegypte,in pharaonem et in omnes servos eius.
PS|135|10|Qui percussit gentes multaset occidit reges fortes:
PS|135|11|Sehon regem Amorraeorumet Og regem Basanet omnia regna Chanaan.
PS|135|12|Et dedit terram eorum hereditatem,hereditatem Israel populo suo.
PS|135|13|Domine, nomen tuum in aeternum;Domine, memoriale tuum in generationem et generationem.
PS|135|14|Quia iudicabit Dominus populum suumet servorum suorum miserebitur.
PS|135|15|Simulacra gentium argentum et aurum,opera manuum hominum.
PS|135|16|Os habent et non loquentur,oculos habent et non videbunt.
PS|135|17|Aures habent et non audient;neque enim est spiritus in ore ipsorum.
PS|135|18|Similes illis erunt, qui faciunt ea,et omnes, qui confidunt in eis.
PS|135|19|Domus Israel, benedicite Domino;domus Aaron, benedicite Domino;
PS|135|20|domus Levi, benedicite Domino;qui timetis Dominum, benedicite Domino.
PS|135|21|Benedictus Dominus ex Sion,qui habitat in Ierusalem. ALLELUIA.
PS|136|1|ALLELUIA.Confitemini Domino, quoniam bonus,quoniam in aeternum misericordia eius.
PS|136|2|Confitemini Deo deorum,quoniam in aeternum misericordia eius.
PS|136|3|Confitemini Domino dominorum,quoniam in aeternum misericordia eius.
PS|136|4|Qui facit mirabilia magna solus,quoniam in aeternum misericordia eius.
PS|136|5|Qui fecit caelos in intellectu,quoniam in aeternum misericordia eius.
PS|136|6|Qui expandit terram super aquas,quoniam in aeternum misericordia eius.
PS|136|7|Qui fecit luminaria magna,quoniam in aeternum misericordia eius:
PS|136|8|solem, ut praeesset diei,quoniam in aeternum misericordia eius;
PS|136|9|lunam et stellas, ut praeessent nocti, quoniam in aeternum misericordia eius.
PS|136|10|Qui percussit Aegyptum in primogenitis eorum,quoniam in aeternum misericordia eius.
PS|136|11|Qui eduxit Israel de medio eorum,quoniam in aeternum misericordia eius,
PS|136|12|in manu potenti et brachio extento,quoniam in aeternum misericordia eius.
PS|136|13|Qui divisit mare Rubrum in divisiones,quoniam in aeternum misericordia eius.
PS|136|14|Et traduxit Israel per medium eius,quoniam in aeternum misericordia eius.
PS|136|15|Et excussit pharaonem et virtutem eius in mari Rubro,quoniam in aeternum misericordia eius.
PS|136|16|Qui traduxit populum suum per desertum,quoniam in aeternum misericordia eius.
PS|136|17|Qui percussit reges magnos,quoniam in aeternum misericordia eius;
PS|136|18|et occidit reges potentes,quoniam in aeternum misericordia eius:
PS|136|19|Sehon regem Amorraeorum,quoniam in aeternum misericordia eius;
PS|136|20|et Og regem Basan,quoniam in aeternum misericordia eius.
PS|136|21|Et dedit terram eorum hereditatem,quoniam in aeternum misericordia eius,
PS|136|22|hereditatem Israel servo suo,quoniam in aeternum misericordia eius.
PS|136|23|Qui in humilitate nostra memor fuit nostri,quoniam in aeternum misericordia eius;
PS|136|24|et redemit nos ab inimicis nostris,quoniam in aeternum misericordia eius.
PS|136|25|Qui dat escam omni carni,quoniam ìn aeternum misericordia eius.
PS|136|26|Confitemini Deo caeli,quoniam in aeternum misericordia eius.
PS|137|1|Super flumina Babylonis,illic sedimus et flevimus,cum recordaremur Sion.
PS|137|2|In salicibus in medio eiussuspendimus citharas nostras.
PS|137|3|Quia illic rogaverunt nos,qui captivos duxerunt nos,verba cantionum,et, qui affligebant nos, laetitiam: Cantate nobis de canticis Sion ".
PS|137|4|Quomodo cantabimus canticum Dominiin terra aliena?
PS|137|5|Si oblitus fuero tui, Ierusalem,oblivioni detur dextera mea;
PS|137|6|adhaereat lingua mea faucibus meis,si non meminero tui,si non praeposuero Ierusalemin capite laetitiae meae.
PS|137|7|Memor esto, Domine, adversus filios Edomdiei Ierusalem;qui dicebant: " Exinanite, exinaniteusque ad fundamentum in ea ".
PS|137|8|Filia Babylonis devastans,beatus, qui retribuet tibi retributionem tuam,quam retribuisti nobis;
PS|137|9|beatus, qui tenebitet allidet parvulos tuos ad petram.
PS|138|1|David.Confitebor tibi, Domine, in toto corde meo,quoniam audisti verba oris mei.In conspectu angelorum psallam tibi,
PS|138|2|adorabo ad templum sanctum tuum;et confitebor nomini tuopropter misericordiam tuam et veritatem tuam,quoniam magnificasti super omne nomen eloquium tuum.
PS|138|3|In quacumque die invocavero te, exaudi me;multiplicabis in anima mea virtutem.
PS|138|4|Confitebuntur tibi, Domine, omnes reges terrae,quia audierunt eloquia oris tui.
PS|138|5|Et cantabunt vias Domini,quoniam magna est gloria Domini;
PS|138|6|quoniam excelsus Dominus et humilem respicitet superbum a longe cognoscit.
PS|138|7|Si ambulavero in medio tribulationis, vivificabis me;et contra iram inimicorum meorum extendes manum tuam,et salvum me faciet dextera tua.
PS|138|8|Dominus perficiet pro me;Domine, misericordia tua in saeculum:opera manuum tuarum ne despicias.
PS|139|1|Magistro chori. David. PSALMUS.Domine, scrutatus es et cognovisti me,
PS|139|2|tu cognovisti sessionem meam et resurrectionem meam.Intellexisti cogitationes meas de longe,
PS|139|3|semitam meam et accubitum meum investigasti.Et omnes vias meas perspexisti,
PS|139|4|quia nondum est sermo in lingua mea,et ecce, Domine, tu novisti omnia.
PS|139|5|A tergo et a fronte coartasti meet posuisti super me manum tuam.
PS|139|6|Mirabilis nimis facta est scientia tua super me,sublimis, et non attingam eam.
PS|139|7|Quo ibo a spiritu tuoet quo a facie tua fugiam?
PS|139|8|Si ascendero in caelum, tu illic es;si descendero in infernum, ades.
PS|139|9|Si sumpsero pennas auroraeet habitavero in extremis maris,
PS|139|10|etiam illuc manus tua deducet me,et tenebit me dextera tua.
PS|139|11|Si dixero: " Forsitan tenebrae compriment me,et nox illuminatio erit circa me ",
PS|139|12|etiam tenebrae non obscurabuntur a te,et nox sicut dies illuminabiturC sicut tenebrae eius ita et lumen eius -.
PS|139|13|Quia tu formasti renes meos,contexuisti me in utero matris meae.
PS|139|14|Confitebor tibi, quia mirabiliter plasmatus sum;mirabilia opera tua,et anima mea cognoscit nimis.
PS|139|15|Non sunt abscondita ossa mea a te,cum factus sum in occulto,contextus in inferioribus terrae.
PS|139|16|Imperfectum adhuc me viderunt oculi tui,et in libro tuo scripti erant omnes dies:ficti erant, et nondum erat unus ex eis.
PS|139|17|Mihi autem nimis pretiosae cogitationes tuae, Deus;nimis gravis summa earum.
PS|139|18|Si dinumerabo eas, super arenam multiplicabuntur;si ad finem pervenerim, adhuc sum tecum.
PS|139|19|Utinam occidas, Deus, peccatores;viri sanguinum, declinate a me.
PS|139|20|Qui loquuntur contra te maligne:exaltantur in vanum contra te.
PS|139|21|Nonne, qui oderunt te, Domine, oderamet insurgentes in te abhorrebam?
PS|139|22|Perfecto odio oderam illos,et inimici facti sunt mihi.
PS|139|23|Scrutare me, Deus, et scito cor meum;proba me et cognosce semitas meas
PS|139|24|et vide, si via vanitatis in me est,et deduc me in via aeterna.
PS|140|1|Magistro chori. PSALMUS. David.
PS|140|2|Eripe me, Domine, ab homine malo, a viro violentiae serva me.
PS|140|3|Qui cogitaverunt mala in corde,tota die constituebant proelia.
PS|140|4|Acuerunt linguas suas sicut serpentis, venenum aspidum sub labiis eorum.
PS|140|5|Custodi me, Domine, de manu peccatoriset a viro violentiae serva me,qui cogitaverunt supplantare gressus meos.
PS|140|6|Absconderunt superbi laqueum mihiet funes extenderunt in rete,iuxta iter offendicula posuerunt mihi.
PS|140|7|Dixi Domino: " Deus meus es tu;auribus percipe, Domine, vocem deprecationis meae ".
PS|140|8|Domine, Domine, virtus salutis meae,obumbrasti caput meum in die belli.
PS|140|9|Ne concedas, Domine, desideria impii;consilia eius ne perficias.
PS|140|10|Exaltant caput, qui circumdant me;malitia labiorum ipsorum operiat eos.
PS|140|11|Cadant super eos carbones ignis,in foveas deicias eos, et non exsurgant.
PS|140|12|Vir linguosus non firmabitur in terra,virum violentiae mala capient in interitu.
PS|140|13|Cognovi quia faciet Dominus iudicium inopiset vindictam pauperum.
PS|140|14|Verumtamen iusti confitebuntur nomini tuo,et habitabunt recti in conspectu tuo.
PS|141|1|PSALMUS. David.Domine, clamavi ad te, ad me festina;intende voci meae, cum clamo ad te.
PS|141|2|Dirigatur oratio mea sicut incensum in conspectu tuo,elevatio manuum mearum ut sacrificium vespertinum. -
PS|141|3|Pone, Domine, custodiam ori meoet vigiliam ad ostium labiorum meorum.
PS|141|4|Non declines cor meum in verbum malitiaead machinandas machinationes in impietatecum hominibus operantibus iniquitatem;et non comedam ex deliciis eorum.
PS|141|5|Percutiat me iustus in misericordia et increpet me;oleum autem peccatoris non impinguet caput meum,quoniam adhuc et oratio mea in malitiis eorum.
PS|141|6|Deiecti in manus duras iudicum eorum,audient verba mea, quoniam suavia erant.
PS|141|7|Sicut frusta dolantis et dirumpentis in terra,dissipata sunt ossa eorum ad fauces inferni.
PS|141|8|Quia ad te, Domine, Domine, oculi mei;ad te confugi, non effundas animam meam.
PS|141|9|Custodi me a laqueo, quem statuerunt mihi,et a scandalis operantium iniquitatem.
PS|141|10|Cadent in retiacula sua peccatores simul,ego autem ultra pertranseam.
PS|142|1|Maskil. David, cum esset in caverna. Precatio.
PS|142|2|Voce mea ad Dominum clamo,voce mea ad Dominum deprecor;
PS|142|3|effundo in conspectu eius lamentationem meam,et tribulationem meam ante ipsum pronuntio.
PS|142|4|Cum deficit in me spiritus meus,tu nosti semitas meas.In via, qua ambulabam,absconderunt laqueum mihi.
PS|142|5|Considerabam ad dexteram et videbam,et non erat qui cognosceret me.Periit fuga a me,et non est qui requirat animam meam. -
PS|142|6|Clamavi ad te, Domine;dixi: " Tu es refugium meum,portio mea in terra viventium.
PS|142|7|Intende ad deprecationem meam,quia humiliatus sum nimis.Libera me a persequentibus me,quia confortati sunt super me.
PS|142|8|Educ de custodia animam meamad confitendum nomini tuo;me circumdabunt iusti,cum retribueris mihi ".
PS|143|1|PSALMUS. David.Domine, exaudi orationem meam, auribus percipe obsecrationem meam in veritate tua;exaudi me in tua iustitia.
PS|143|2|Et non intres in iudicium cum servo tuo,quia non iustificabitur in conspectu tuo omnis vivens.
PS|143|3|Quia persecutus est inimicus animam meam,contrivit in terra vitam meam,collocavit me in obscuris sicut mortuos a saeculo.
PS|143|4|Et anxiatus est in me spiritus meus,in medio mei obriguit cor meum.
PS|143|5|Memor fui dierum antiquorum,meditatus sum in omnibus operibus tuis,in factis manuum tuarum recogitabam.
PS|143|6|Expandi manus meas ad te,anima mea sicut terra sine aqua tibi.
PS|143|7|Velociter exaudi me, Domine;defecit spiritus meus.Non abscondas faciem tuam a me,ne similis fiam descendentibus in lacum.
PS|143|8|Auditam fac mihi mane misericordiam tuam,quia in te speravi.Notam fac mihi viam, in qua ambulem,quia ad te levavi animam meam.
PS|143|9|Eripe me de inimicis meis,Domine, ad te confugi.
PS|143|10|Doce me facere voluntatem tuam,quia Deus meus es tu.Spiritus tuus bonus deducet me in terram rectam;
PS|143|11|propter nomen tuum, Domine, vivificabis me.In iustitia tua educes de tribulatione animam meam
PS|143|12|et in misericordia tua disperdes inimicos meos;et perdes omnes, qui tribulant animam meam,quoniam ego servus tuus sum.
PS|144|1|David.Benedictus Dominus, adiutor meus,qui docet manus meas ad proeliumet digitos meos ad bellum.
PS|144|2|Misericordia mea et fortitudo mea,refugium meum et liberator meus;scutum meum, et in ipso speravi,qui subdit populum meum sub me.
PS|144|3|Domine, quid est homo, quod agnoscis eum,aut filius hominis, quod reputas eum?
PS|144|4|Homo vanitati similis factus est,dies eius sicut umbra praeteriens.
PS|144|5|Domine, inclina caelos tuos et descende;tange montes, et fumigabunt.
PS|144|6|Fulgura coruscationem et dissipa eos;emitte sagittas tuas et conturba eos.
PS|144|7|Emitte manum tuam de alto;eripe me et libera me de aquis multis,de manu filiorum alienigenarum,
PS|144|8|quorum os locutum est vanitatem,et dextera eorum dextera mendacii.
PS|144|9|Deus, canticum novum cantabo tibi,in psalterio decachordo psallam tibi,
PS|144|10|qui das salutem regibus,qui redimis David servum tuum de gladio maligno.
PS|144|11|Eripe me et libera mede manu filiorum alienigenarum,quorum os locutum est vanitatem,et dextera eorum dextera mendacii.
PS|144|12|Filii nostri sicut novellae crescentesin iuventute sua;filiae nostrae sicut columnae angulares,sculptae ut structura templi.
PS|144|13|Promptuaria nostra plena,redundantia omnibus bonis;oves nostrae in milibusinnumerabiles in campis nostris,
PS|144|14|boves nostrae crassae.Non est ruina maceriae neque egressusneque clamor in plateis nostris.
PS|144|15|Beatus populus, cui haec sunt;beatus populus, cui Dominus est Deus.
PS|145|1|Laudes. David.ALEPH. Exaltabo te, Deus meus, rex,et benedicam nomini tuoin saeculum et in saeculum saeculi.
PS|145|2|BETH. Per singulos dies benedicam tibiet laudabo nomen tuumin saeculum et in saeculum saeculi.
PS|145|3|GHIMEL. Magnus Dominus et laudabilis nimis,et magnitudinis eius non est investigatio.
PS|145|4|DALETH. Generatio generationi laudabit opera tua,et potentiam tuam pronuntiabunt.
PS|145|5|HE. Magnificentiam gloriae maiestatis tuae loquenturet mirabilia tua enarrabunt.
PS|145|6|VAU. Et virtutem terribilium tuorum dicentet magnitudinem tuam narrabunt.
PS|145|7|ZAIN. Memoriam abundantiae suavitatis tuae eructabuntet iustitia tua exsultabunt.
PS|145|8|HETH. Miserator et misericors Dominus,longanimis et multae misericordiae.
PS|145|9|TETH. Suavis Dominus universis,et miserationes eius super omnia opera eius.
PS|145|10|IOD. Confiteantur tibi, Domine, omnia opera tua;et sancti tui benedicant tibi.
PS|145|11|CAPH. Gloriam regni tui dicantet potentiam tuam loquantur,
PS|145|12|LAMED. ut notas faciant filiis hominum potentias tuaset gloriam magnificentiae regni tui.
PS|145|13|MEM. Regnum tuum regnum omnium saeculorum,et dominatio tua in omnem generationem et generationem.NUN. Fidelis Dominus in omnibus verbis suiset sanctus in omnibus operibus suis.
PS|145|14|SAMECH. Allevat Dominus omnes, qui corruunt,et erigit omnes depressos.
PS|145|15|AIN. Oculi omnium in te sperant,et tu das illis escam in tempore opportuno.
PS|145|16|PHE. Aperis tu manum tuamet imples omne animal in beneplacito.
PS|145|17|SADE. Iustus Dominus in omnibus viis suiset sanctus in omnibus operibus suis.
PS|145|18|COPH. Prope est Dominus omnibus invocantibus eum,omnibus invocantibus eum in veritate.
PS|145|19|RES. Voluntatem timentium se facietet deprecationem eorum exaudiet et salvos faciet eos.
PS|145|20|SIN. Custodit Dominus omnes diligentes seet omnes peccatores disperdet.
PS|145|21|TAU. Laudationem Domini loquetur os meum,et benedicat omnis caro nomini sancto eiusin saeculum et in saeculum saeculi.
PS|146|1|ALLELUIA.Lauda, anima mea, Dominum;
PS|146|2|laudabo Dominum in vita mea,psallam Deo meo, quamdiu fuero.
PS|146|3|Nolite confidere in principibus,in filiis hominum, in quibus non est salus.
PS|146|4|Exibit spiritus eius, et revertetur in terram suam;in illa die peribunt cogitationes eorum.
PS|146|5|Beatus, cuius Deus Iacob est adiutor,cuius spes in Domino Deo suo,
PS|146|6|qui fecit caelum et terram,mare et omnia, quae in eis sunt;qui custodit veritatem in saeculum,
PS|146|7|facit iudicium oppressis,dat escam esurientibus.Dominus solvit compeditos,
PS|146|8|Dominus illuminat caecos,Dominus erigit depressos,Dominus diligit iustos,
PS|146|9|Dominus custodit advenas,pupillum et viduam sustentatet viam peccatorum disperdit.
PS|146|10|Regnabit Dominus in saecula,Deus tuus, Sion,in generationem et generationem.
PS|147|1|ALLELUIA.Laudate Dominum, quoniam bonum est psallere Deo nostro,quoniam iucundum est celebrare laudem.
PS|147|2|Aedificans Ierusalem Dominus,dispersos Israelis congregabit.
PS|147|3|Qui sanat contritos cordeet alligat plagas eorum;
PS|147|4|qui numerat multitudinem stellarumet omnibus eis nomina vocat.
PS|147|5|Magnus Dominus noster et magnus virtute,sapientiae eius non est numerus.
PS|147|6|Sustentat mansuetos Dominus,humilians autem peccatores usque ad terram.
PS|147|7|Praecinite Domino in confessione,psallite Deo nostro in cithara.
PS|147|8|Qui operit caelum nubibuset parat terrae pluviam.Qui producit in montibus fenumet herbam servituti hominum.
PS|147|9|Qui dat iumentis escam ipsorumet pullis corvorum invocantibus eum.
PS|147|10|Non in fortitudine equi delectatur,nec in tibiis viri beneplacitum est ei.
PS|147|11|Beneplacitum est Domino super timentes eumet in eis, qui sperant super misericordia eius.
PS|147|12|Lauda, Ierusalem, Dominum;collauda Deum tuum, Sion.
PS|147|13|Quoniam confortavit seras portarum tuarum,benedixit filiis tuis in te.
PS|147|14|Qui ponit fines tuos pacemet adipe frumenti satiat te.
PS|147|15|Qui emittit eloquium suum terrae,velociter currit verbum eius.
PS|147|16|Qui dat nivem sicut lanam,pruinam sicut cinerem spargit.
PS|147|17|Mittit crystallum suam sicut buccellas;ante faciem frigoris eius quis sustinebit?
PS|147|18|Emittet verbum suum et liquefaciet ea,flabit spiritus eius, et fluent aquae.
PS|147|19|Qui annuntiat verbum suum Iacob,iustitias et iudicia sua Israel.
PS|147|20|Non fecit taliter omni nationiet iudicia sua non manifestavit eis. ALLELUIA.
PS|148|1|ALLELUIA.Laudate Dominum de caelis,laudate eum in excelsis.
PS|148|2|Laudate eum, omnes angeli eius,laudate eum, omnes virtutes eius.
PS|148|3|Laudate eum, sol et luna,laudate eum, omnes stellae lucentes.
PS|148|4|Laudate eum, caeli caelorumet aquae omnes, quae super caelos sunt. -
PS|148|5|Laudent nomen Domini,quia ipse mandavit, et creata sunt;
PS|148|6|statuit ea in aeternum et in saeculum saeculi;praeceptum posuit, et non praeteribit.
PS|148|7|Laudate Dominum de terra,dracones et omnes abyssi,
PS|148|8|ignis, grando, nix, fumus,spiritus procellarum, qui facit verbum eius,
PS|148|9|montes et omnes colles,ligna fructifera et omnes cedri,
PS|148|10|bestiae et universa pecora,serpentes et volucres pennatae.
PS|148|11|Reges terrae et omnes populi,principes et omnes iudices terrae,
PS|148|12|iuvenes et virgines,senes cum iunioribus
PS|148|13|laudent nomen Domini,quia exaltatum est nomen eius solius.Magnificentia eius super caelum et terram,
PS|148|14|et exaltavit cornu populi sui.Hymnus omnibus sanctis eius,filiis Israel, populo, qui propinquus est ei. ALLELUIA.
PS|149|1|ALLELUIA.Cantate Domino canticum novum;laus eius in ecclesia sanctorum.
PS|149|2|Laetetur Israel in eo, qui fecit eum,et filii Sion exsultent in rege suo.
PS|149|3|Laudent nomen eius in choro,in tympano et cithara psallant ei,
PS|149|4|quia beneplacitum est Domino in populo suo,et honorabit mansuetos in salute.
PS|149|5|Iubilent sancti in gloria,laetentur in cubilibus suis.
PS|149|6|Exaltationes Dei in gutture eorum,et gladii ancipites in manibus eorum,
PS|149|7|ad faciendam vindictam in nationibus,castigationes in populis,
PS|149|8|ad alligandos reges eorum in compedibuset nobiles eorum in manicis ferreis,
PS|149|9|ad faciendum in eis iudicium conscriptum.Gloria haec est omnibus sanctis eius. ALLELUIA.
PS|150|1|ALLELUIA.Laudate Dominum in sanctuario eius,laudate eum in firmamento virtutis eius.
PS|150|2|Laudate eum in magnalibus eius,laudate eum secundum multitudinem magnitudinis eius.
PS|150|3|Laudate eum in sono tubae,laudate eum in psalterio et cithara,
PS|150|4|laudate eum in tympano et choro,laudate eum in chordis et organo,
PS|150|5|laudate eum in cymbalis benesonantibus,laudate eum in cymbalis iubilationis:omne quod spirat, laudet Dominum. ALLELUIA.
PROV|1|1|Parabolae Salomonis filii David regis Israel
PROV|1|2|ad sciendam sapientiam et disciplinam,ad intellegenda verba prudentiae;
PROV|1|3|ad suscipiendam eruditionem doctrinae,iustitiam et iudicium et aequitatem,
PROV|1|4|ut detur parvulis astutia,adulescenti scientia et recogitatio.
PROV|1|5|Audiat sapiens et addet doctrinam,et intellegens dispositiones possidebit:
PROV|1|6|animadvertet parabolam et allegoriam,verba sapientium et aenigmata eorum.
PROV|1|7|Timor Domini principium scientiae.Sapientiam atque doctrinam stulti despiciunt.
PROV|1|8|Audi, fili mi, disciplinam patris tuiet ne reicias legem matris tuae,
PROV|1|9|quia diadema gratiae sunt capiti tuo,et torques collo tuo.
PROV|1|10|Fili mi, si te lactaverint peccatores,ne acquiescas eis.
PROV|1|11|Si dixerint: " Veni nobiscum, insidiemur sanguini,abscondamus tendiculas contra insontem frustra;
PROV|1|12|deglutiamus eos sicut infernus viventeset integros quasi descendentes in lacum:
PROV|1|13|omnem pretiosam substantiam reperiemus,implebimus domos nostras spoliis;
PROV|1|14|sortem mitte nobiscum,marsupium unum sit omnium nostrum ";
PROV|1|15|fili mi, ne ambules cum eis,prohibe pedem tuum a semitis eorum.
PROV|1|16|Pedes enim illorum ad malum curruntet festinant, ut effundant sanguinem.
PROV|1|17|Frustra autem iacitur rete ante oculos pinnatorum.
PROV|1|18|Ipsique contra sanguinem suum insidianturet moliuntur fraudes contra animas suas.
PROV|1|19|Sic semitae omnis ad rapinam intenti:animam ipsius possidentis rapiunt.
PROV|1|20|Sapientia foris praedicat,in plateis dat vocem suam,
PROV|1|21|in capite viarum frequentium clamitat,in foribus portarum urbis profert verba sua:
PROV|1|22|" Usquequo, parvuli, diligitis infantiam,et derisores sibi derisionem cupient,et imprudentes odibunt scientiam?
PROV|1|23|Convertimini ad correptionem meam;en proferam vobis spiritum meumet ostendam vobis verba mea.
PROV|1|24|Quia vocavi, et renuistis,extendi manum meam, et non fuit qui aspiceret;
PROV|1|25|despexistis omne consilium meumet increpationes meas neglexistis.
PROV|1|26|Ego quoque in interitu vestro rideboet subsannabo, cum terror vobis advenerit,
PROV|1|27|cum irruerit ut procella terror,et interitus quasi tempestas ingruerit,quando venerit super vos tribulatio et angustia ".
PROV|1|28|Tunc invocabunt me, et non exaudiam,instanter quaerent me et non invenient me,
PROV|1|29|eo quod exosam habuerint disciplinamet timorem Domini non elegerint
PROV|1|30|nec acquieverint consilio meoet despexerint universam correptionem meam.
PROV|1|31|Comedent igitur fructus viae suaesuisque consiliis saturabuntur.
PROV|1|32|Aversio parvulorum interficiet eos,et securitas stultorum perdet illos.
PROV|1|33|Qui autem me audierit, absque terrore requiescetet tranquillus erit timore malorum sublato.
PROV|2|1|Fili mi, si susceperis sermones meoset mandata mea absconderis penes te,
PROV|2|2|intendens ad sapientiam aurem tuam,inclinans cor tuum ad cognoscendam prudentiam;
PROV|2|3|si enim sapientiam invocaveriset dederis vocem tuam prudentiae,
PROV|2|4|si quaesieris eam quasi pecuniamet sicut thesauros conquisieris illam,
PROV|2|5|tunc intelleges timorem Dominiet scientiam Dei invenies.
PROV|2|6|Quia Dominus dat sapientiam,et ex ore eius scientia et prudentia.
PROV|2|7|Thesaurizabit rectis sollertiamet clipeus erit gradientibus simpliciter
PROV|2|8|servans semitas iustitiaeet vias sanctorum custodiens.
PROV|2|9|Tunc intelleges iustitiam et iudiciumet aequitatem et omnem semitam bonam,
PROV|2|10|quia intrabit sapientia cor tuum,et scientia animae tuae placebit.
PROV|2|11|Consilium custodiet te,et prudentia servabit te,
PROV|2|12|ut eruaris a via malaet ab homine, qui perversa loquitur;
PROV|2|13|qui relinquunt iter rectum,ut ambulent per vias tenebrosas;
PROV|2|14|qui laetantur, cum malefecerint,et exsultant in rebus pessimis:
PROV|2|15|quorum viae perversae sunt,et pravi gressus eorum.
PROV|2|16|Ut eruaris a muliere alienaet ab extranea, quae mollit sermones suos
PROV|2|17|et relinquit ducem pubertatis suaeet pacti Dei sui oblita est.
PROV|2|18|Inclinata est enim ad mortem domus eius,et ad inferos semitae ipsius;
PROV|2|19|omnes, qui ingrediuntur ad eam, non revertenturnec apprehendent semitas vitae.
PROV|2|20|Ut ambules in via bonorumet calles iustorum custodias:
PROV|2|21|qui enim recti sunt, habitabunt in terra,et simplices permanebunt in ea;
PROV|2|22|impii vero de terra perdentur,et, qui inique agunt, auferentur ex ea.
PROV|3|1|Fili mi, ne obliviscaris legis meae,et praecepta mea cor tuum custodiat;
PROV|3|2|longitudinem enim dierum et annos vitaeet pacem apponent tibi.
PROV|3|3|Misericordia et veritas te non deserant;circumda eas gutturi tuoet describe in tabulis cordis tui,
PROV|3|4|et invenies gratiam et successum bonumcoram Deo et hominibus.
PROV|3|5|Habe fiduciam in Domino ex toto corde tuoet ne innitaris prudentiae tuae.
PROV|3|6|In omnibus viis tuis cogita illum,et ipse diriget gressus tuos.
PROV|3|7|Ne sis sapiens apud temetipsum;time Dominum et recede a malo.
PROV|3|8|Sanitas quippe erit umbilico tuo,et irrigatio ossibus tuis.
PROV|3|9|Honora Dominum de tua substantiaet de primitiis omnium frugum tuarum,
PROV|3|10|et implebuntur horrea tua frumento,et vino torcularia tua redundabunt.
PROV|3|11|Disciplinam Domini, fili mi, ne abiciasnec asperneris, cum ab eo corriperis:
PROV|3|12|quem enim diligit, Dominus corripitet quasi pater in filio complacet sibi.
PROV|3|13|Beatus homo, qui invenit sapientiamet qui affluit prudentia:
PROV|3|14|melior est acquisitio eius negotiatione argenti,et auro primo fructus eius.
PROV|3|15|Pretiosior est cunctis gemmis,et omnia pretiosa tua huic non valent comparari;
PROV|3|16|longitudo dierum in dextera eius,et in sinistra illius divitiae et gloria.
PROV|3|17|Viae eius viae pulchrae,et omnes semitae illius pacificae.
PROV|3|18|Lignum vitae est his, qui apprehenderint eam;et, qui tenuerit eam, beatus.
PROV|3|19|Dominus sapientia fundavit terram,stabilivit caelos prudentia;
PROV|3|20|sapientia illius eruperunt abyssi,et nubes rorem stillant.
PROV|3|21|Fili mi, ne effluant haec ab oculis tuis;custodi prudentiam atque consilium,
PROV|3|22|et erit vita animae tuae,et gratia collo tuo;
PROV|3|23|tunc ambulabis fiducialiter in via tua,et pes tuus non impinget.
PROV|3|24|Si dormieris, non timebis;quiesces, et suavis erit somnus tuus.
PROV|3|25|Ne paveas repentino terroreet irruentem tibi turbinem impiorum, cum venerit.
PROV|3|26|Dominus enim erit in latere tuoet custodiet pedem tuum, ne capiaris.
PROV|3|27|Noli prohibere beneficium ab eo, cui debetur,si in potestate manus tuae est, ut facias.
PROV|3|28|Ne dicas amico tuo: " Vade et revertere,cras dabo tibi ", cum statim possis dare.
PROV|3|29|Ne moliaris amico tuo malum,cum ille apud te sedeat cum fiducia.
PROV|3|30|Ne contendas adversus hominem frustra,cum ipse tibi nihil mali fecerit.
PROV|3|31|Ne aemuleris hominem iniustumnec imiteris omnes vias eius,
PROV|3|32|quia abominatio Domini est omnis pravus,et cum simplicibus societas eius.
PROV|3|33|Maledictio a Domino in domo impii,habitacula autem iustorum benedicentur.
PROV|3|34|Ipse deludet illusoreset mansuetis dabit gratiam;
PROV|3|35|gloriam sapientes possidebunt,stultorum exaltatio ignominia.
PROV|4|1|Audite, filii, disciplinam patriset attendite, ut sciatis prudentiam;
PROV|4|2|quoniam doctrinam bonam tribuam vobis,legem meam ne derelinquatis.
PROV|4|3|Nam et ego filius fui patris mei,tenellus et unigenitus coram matre mea;
PROV|4|4|et docebat me atque dicebat: Suscipiat verba mea cor tuum,custodi praecepta mea et vives.
PROV|4|5|Posside sapientiam, posside prudentiam,ne obliviscaris neque declines a verbis oris mei.
PROV|4|6|Ne dimittas eam, et custodiet te,dilige eam, et servabit te.
PROV|4|7|Principium sapientiae: posside sapientiamet in omni possessione tua acquire prudentiam.
PROV|4|8|Arripe illam, et exaltabit te,glorificaberis ab ea, cum eam fueris amplexatus.
PROV|4|9|Dabit capiti tuo diadema gratiae,et corona inclita proteget te ".
PROV|4|10|Audi, fili mi, et suscipe verba mea,ut multiplicentur tibi anni vitae.
PROV|4|11|Viam sapientiae monstravi tibi;duxi te per semitas aequitatis,
PROV|4|12|quas cum ingressus fueris, non arctabuntur gressus tui,et currens non habebis offendiculum.
PROV|4|13|Tene disciplinam nec laxes;custodi illam, quia ipsa est vita tua.
PROV|4|14|Ne ingrediaris in semitas impiorumnec procedas in malorum via.
PROV|4|15|Fuge ab ea nec transeas per illam;declina et desere eam.
PROV|4|16|Non enim dormiunt, nisi malefecerint,et rapitur somnus ab eis, nisi supplantaverint.
PROV|4|17|Comedunt enim panem impietatiset vinum iniquitatis bibunt.
PROV|4|18|Iustorum autem semita quasi lux splendensprocedit et crescit usque ad perfectam diem.
PROV|4|19|Via impiorum tenebrosa;nesciunt, ubi corruant.
PROV|4|20|Fili mi, ausculta sermones meoset ad eloquia mea inclina aurem tuam;
PROV|4|21|ne recedant ab oculis tuis,custodi ea in medio cordis tui:
PROV|4|22|vita enim sunt invenientibus ea,et universae carni sanitas.
PROV|4|23|Omni custodia serva cor tuum,quia ex ipso vita procedit.
PROV|4|24|Remove a te os pravum,et detrahentia labia sint procul a te.
PROV|4|25|Oculi tui recta videant,et palpebrae tuae dirigantur coram te.
PROV|4|26|Observa semitam pedum tuorum,et omnes viae tuae stabilientur.
PROV|4|27|Ne declines ad dexteram neque ad sinistram,averte pedem tuum a malo.
PROV|5|1|Fili mi, attende ad sapientiam meam,et prudentiae meae inclina aurem tuam,
PROV|5|2|ut custodias cogitationes,et disciplinam labia tua conservent.
PROV|5|3|Favum enim stillant labia meretricis,et nitidius oleo guttur eius;
PROV|5|4|novissima autem illius amara quasi absinthiumet acuta quasi gladius biceps.
PROV|5|5|Pedes eius descendunt in mortem,et ad inferos gressus illius tendunt;
PROV|5|6|cum non observet semitam vitae,vagi sunt gressus eius, et ipsa nescit.
PROV|5|7|Nunc ergo, fili mi, audi meet ne recedas a verbis oris mei.
PROV|5|8|Longe fac ab ea viam tuamet ne appropinques foribus domus eius.
PROV|5|9|Ne des alienis honorem tuumet annos tuos crudeli,
PROV|5|10|ne forte impleantur extranei viribus tuis,et labores tui sint in domo aliena,
PROV|5|11|et gemas in novissimis,quando consumpseris carnes tuas et corpus tuum
PROV|5|12|et dicas: " Cur detestatus sum disciplinam,et increpationes renuit cor meum,
PROV|5|13|nec audivi vocem docentium meet magistris non inclinavi aurem meam?
PROV|5|14|Paene fui in omni malo,in medio ecclesiae et synagogae ".
PROV|5|15|Bibe aquam de cisterna tuaet fluenta putei tui,
PROV|5|16|ne deriventur fontes tui foras,et in plateis rivi aquarum;
PROV|5|17|habeto eas solus,nec sint alieni participes tui.
PROV|5|18|Sit vena tua benedicta,et laetare cum muliere adulescentiae tuae;
PROV|5|19|cerva carissima et gratissimus hinnulus,blanditiae eius inebrient te in omni tempore,in amore eius delectare iugiter.
PROV|5|20|Quare seduceris, fili mi, ab alienaet foveris in sinu extraneae?
PROV|5|21|Quoniam ante Dominum viae hominis,et omnes gressus eius considerat.
PROV|5|22|Iniquitates suae capient impium,et funibus peccatorum suorum constringetur.
PROV|5|23|Ipse morietur, quia non habuit disciplinam,et in multitudine stultitiae suae decipietur.
PROV|6|1|Fili mi, si spoponderis pro amico tuo,defixisti apud extraneum manum tuam;
PROV|6|2|illaqueatus es verbis oris tuiet captus propriis sermonibus.
PROV|6|3|Fac ergo, quod dico, fili mi, et temetipsum libera,quia incidisti in manum proximi tui;discurre, prosternere, insta amico tuo.
PROV|6|4|Ne dederis somnum oculis tuisnec palpebris tuis dormitationem.
PROV|6|5|Eruere quasi dammula de rete,et quasi avis de manu aucupis.
PROV|6|6|Vade ad formicam, o piger,et considera vias eius et disce sapientiam.
PROV|6|7|Quae, cum non habeat ducemnec praeceptorem nec principem,
PROV|6|8|parat in aestate cibum sibiet congregat in messe, quod comedat.
PROV|6|9|Usquequo, piger, dormies?Quando consurges e somno tuo?
PROV|6|10|Paululum dormis, paululum dormitas,paululum conseres manus, ut dormias;
PROV|6|11|et veniet tibi quasi viator egestas,et pauperies quasi vir armatus.
PROV|6|12|Homo iniquus, vir inutilis,graditur ore perverso;
PROV|6|13|annuit oculis, terit pede,digito loquitur.
PROV|6|14|Prava in corde suo machinatur,malum in omni tempore, iurgia seminat.
PROV|6|15|Ideo extemplo veniet perditio sua,et subito conteretur nec habebit medicinam.
PROV|6|16|Sex sunt, quae odit Dominus,et septem detestatur anima eius:
PROV|6|17|oculos sublimes, linguam mendacem,manus effundentes innoxium sanguinem,
PROV|6|18|cor machinans cogitationes pravas,pedes veloces ad currendum in malum,
PROV|6|19|proferentem mendacia, testem fallacemet eum, qui seminat inter fratres discordias.
PROV|6|20|Conserva, fili mi, praecepta patris tuiet ne reicias legem matris tuae;
PROV|6|21|liga ea in corde tuo iugiteret circumda gutturi tuo.
PROV|6|22|Cum ambulaveris, dirigent te,cum dormieris, custodient teet, cum evigilaveris, colloquentur tecum.
PROV|6|23|Quia mandatum lucerna est, et lex lux,et via vitae increpatio disciplinae,
PROV|6|24|ut custodiant te a muliere malaet a blanda lingua extraneae;
PROV|6|25|non concupiscat pulchritudinem eius cor tuum,nec capiaris nutibus illius:
PROV|6|26|pretium enim scorti vix est torta panis,mulier autem viri pretiosam animam capit.
PROV|6|27|Numquid potest homo abscondere ignem in sinu suo,et vestimenta illius non ardebunt?
PROV|6|28|Aut ambulare super prunas,et non comburentur plantae eius?
PROV|6|29|Sic qui ingreditur ad mulierem proximi sui;non erit mundus, quicumque tetigerit eam.
PROV|6|30|Non contemptui erit fur, cum furatus fuerit,ut esurientem impleat animam.
PROV|6|31|Deprehensus quoque reddet septuplumet omnem substantiam domus suae tradet.
PROV|6|32|Qui autem adulter est cum muliere, vecors est;perdet animam suam, qui hoc fecerit.
PROV|6|33|Plagam et ignominiam congregat sibi,et opprobrium illius non delebitur.
PROV|6|34|Quia zelus est furor viri,et non parcet in die vindictae
PROV|6|35|nec accipiet personam tuam in piaculumnec suscipiet dona plurima.
PROV|7|1|Fili mi, custodi sermones meoset praecepta mea reconde tibi.
PROV|7|2|Serva mandata mea et vives,et legem meam quasi pupillam oculi tui.
PROV|7|3|Liga ea in digitis tuis,scribe illa in tabulis cordis tui.
PROV|7|4|Dic sapientiae: " Soror mea es "et prudentiam voca Amicam,
PROV|7|5|ut custodiat te a muliere extraneaet ab aliena, quae verba sua dulcia facit.
PROV|7|6|De fenestra enim domus meaeper cancellos prospexi
PROV|7|7|et video inter parvulos;considero inter filios vecordem iuvenem,
PROV|7|8|qui transit per plateam iuxta angulumet prope viam domus illius graditur
PROV|7|9|in obscuro advesperascente die,in mediis tenebris et caligine.
PROV|7|10|Et ecce, occurrit illi mulier ornatu meretricio,cauta corde, garrula et rebellans,
PROV|7|11|quietis impatiensnec valens in domo consistere pedibus suis:
PROV|7|12|nunc foris, nunc in plateiset iuxta angulos insidians.
PROV|7|13|Apprehensumque deosculatur iuvenemet procaci vultu blanditur dicens:
PROV|7|14|" Victimas pro salute vovi,hodie reddidi vota mea;
PROV|7|15|idcirco egressa sum in occursum tuumdesiderans te videre et repperi.
PROV|7|16|Stragulatis vestibus lectulum meum stravi,linteis pictis ex Aegypto;
PROV|7|17|aspersi cubile meum myrrhaet aloe et cinnamomo.
PROV|7|18|Veni, inebriemur voluptatibus,usque mane fruamur amoribus.
PROV|7|19|Non est enim vir in domo sua;abiit via longissima,
PROV|7|20|sacculum pecuniae secum tulit,in die plenae lunae reversurus est in domum suam ".
PROV|7|21|Irretivit eum multis sermonibuset blanditiis labiorum protraxit illum.
PROV|7|22|Stultus eam sequitur quasi bos ductus ad victimam,sicut irretitur vinculo cervus,
PROV|7|23|donec transfigat sagitta iecur eius;velut si avis festinet ad laqueumet nescit quod de periculo animae illius agitur.
PROV|7|24|Nunc ergo, fili mi, audi meet attende verbis oris mei.
PROV|7|25|Ne abstrahatur in viis illius mens tua,neque decipiaris semitis eius.
PROV|7|26|Multos enim vulneratos deiecit,et fortissimi quique interfecti sunt ab ea:
PROV|7|27|viae inferi domus eiuspenetrantes in interiora mortis.
PROV|8|1|Numquid non sapientia clamitat,et prudentia dat vocem suam?
PROV|8|2|In summis verticibussupra viam in mediis semitis stans,
PROV|8|3|iuxta portas ad introitum civitatis,in ipsis foribus conclamat:
PROV|8|4|" O viri, ad vos clamito,et vox mea ad filios hominum.
PROV|8|5|Intellegite, parvuli, astutiam;et insipientes, animadvertite.
PROV|8|6|Audite, quoniam de rebus magnis locutura sum,et aperientur labia mea, ut recta praedicent.
PROV|8|7|Veritatem meditabitur guttur meum,et labia mea detestabuntur impium.
PROV|8|8|Iusti sunt omnes sermones oris mei,non est in eis pravum quid neque perversum;
PROV|8|9|omnes recti sunt intellegentibuset aequi invenientibus scientiam.
PROV|8|10|Accipitc disciplinam meam et non pecuniam,doctrinam magis quam aurum electum.
PROV|8|11|Melior est enim sapientia gemmis,et omne desiderabile ei non potest comparari ".
PROV|8|12|Ego sapientia habito cum prudentiaet artem excogitandi invenio.
PROV|8|13|Timor Domini odisse malum;arrogantiam et superbiam et viam pravamet os bilingue detestor.
PROV|8|14|Meum est consilium et prudentia,mea est intellegentia, mea est fortitudo.
PROV|8|15|Per me reges regnant,et principes iusta decernunt;
PROV|8|16|per me duces imperant,et potentes decernunt iustitiam.
PROV|8|17|Ego diligentes me diligo;et, qui mane vigilant ad me, invenient me.
PROV|8|18|Mecum sunt divitiae et gloria,opes superbae et iustitia.
PROV|8|19|Melior est enim fructus meus auro et obryzo,et genimina mea argento electo.
PROV|8|20|In viis iustitiae ambulo,in medio semitarum iudicii,
PROV|8|21|ut ditem diligentes meet thesauros eorum repleam.
PROV|8|22|Dominus possedit me in initio viarum suarum,antequam quidquam faceret a principio;
PROV|8|23|ab aeterno ordinata sumet ex antiquis, antequam terra fieret.
PROV|8|24|Nondum erant abyssi, et ego iam concepta eram,necdum fontes graves aquis,
PROV|8|25|priusquam montes demergerentur,ante colles ego parturiebar.
PROV|8|26|Adhuc terram non fecerat et camposet initium glebae orbis terrae.
PROV|8|27|Quando praeparabat caelos, aderam,quando certa lege et gyro vallabat abyssos,
PROV|8|28|quando nubes firmabat sursum,et praevaluerunt fontes abyssi,
PROV|8|29|quando circumdabat mari terminum suumet aquis, ne transirent fines suos,quando iecit fundamenta terrae,
PROV|8|30|cum eo eram ut artifex:delectatio eius per singulos dies,ludens coram eo omni tempore,
PROV|8|31|ludens in orbe terrarum,et deliciae meae esse cum filiis hominum.
PROV|8|32|Nunc ergo, filii, audite me:beati, qui custodiunt vias meas;
PROV|8|33|audite disciplinam et estote sapienteset nolite abicere eam.
PROV|8|34|Beatus homo, qui audit meet qui vigilat ad fores meas cotidieet observat ad postes ostii mei.
PROV|8|35|Qui me invenerit, inveniet vitamet hauriet delicias a Domino.
PROV|8|36|Qui autem in me peccaverit, laedet animam suam:omnes, qui me oderunt, diligunt mortem.
PROV|9|1|Sapientia aedificavit sibi domum,excidit columnas septem;
PROV|9|2|immolavit victimas suas, miscuit vinumet proposuit mensam suam.
PROV|9|3|Misit ancillas suas, ut vocarentad arcem et ad excelsa civitatis:
PROV|9|4|" Si quis est parvulus, veniat ad me ".Et vecordi locuta est:
PROV|9|5|" Venite, comedite panem meumet bibite vinum, quod miscui vobis;
PROV|9|6|relinquite infantiam et viviteet ambulate per vias prudentiae ".
PROV|9|7|Qui erudit derisorem, ipse iniuriam sibi facit;et, qui arguit impium, sibi maculam generat.
PROV|9|8|Noli arguere derisorem, ne oderit te;argue sapientem, et diliget te.
PROV|9|9|Da sapienti, et sapientior fiet;doce iustum, et addet doctrinam.
PROV|9|10|Principium sapientiae timor Domini,et scientia Sancti est prudentia.
PROV|9|11|Per me enim multiplicabuntur dies tui,et addentur tibi anni vitae.
PROV|9|12|Si sapiens fueris, tibimetipsi eris;si autem illusor, solus portabis malum.
PROV|9|13|Mulier stulta est clamosa,fatua et nihil sciens;
PROV|9|14|sedit in foribus domus suaesuper sellam in excelsis urbis,
PROV|9|15|ut vocaret transeuntes per viamet pergentes itinere suo:
PROV|9|16|" Qui est parvulus, declinet ad me ".Et vecordi locuta est:
PROV|9|17|" Aquae furtivae dulciores sunt,et panis in abscondito suavior ".
PROV|9|18|Et ignoravit quod ibi sint umbrae,et in profundis inferni convivae eius.
PROV|10|1|Parabolae Salomonis.Filius sapiens laetificat pa trem,filius vero stultus maestitia est matris suae.
PROV|10|2|Nil proderunt thesauri impietatis,iustitia vero liberabit a morte.
PROV|10|3|Non affliget Dominus fame animam iustiet cupiditatem impiorum subvertet.
PROV|10|4|Egestatem operata est manus remissa,manus autem fortium divitias parat.
PROV|10|5|Qui congregat in messe, filius sapiens est;qui autem stertit aestate, filius confusionis.
PROV|10|6|Benedictiones Domini super caput iusti,os autem impiorum operit violentiam.
PROV|10|7|Memoria iusti in benedictione erit,et nomen impiorum putrescet.
PROV|10|8|Sapiens corde praecepta suscipit,et stultus labiis corruet.
PROV|10|9|Qui ambulat simpliciter, ambulat confidenter;qui autem depravat vias suas, manifestus erit.
PROV|10|10|Qui annuit oculo, dabit dolorem,et stultus labiis corruet.
PROV|10|11|Vena vitae os iusti,et os impiorum operit violentiam.
PROV|10|12|Odium suscitat rixas,et universa delicta operit caritas.
PROV|10|13|In labiis sapientis invenitur sapientia,et virga in dorso eius, qui indiget corde.
PROV|10|14|Sapientes recondunt scientiam,os autem stulti ruinae proximum est.
PROV|10|15|Substantia divitis urbs fortitudinis eius,ruina pauperum egestas eorum.
PROV|10|16|Opus iusti ad vitam,fructus autem impii ad peccatum.
PROV|10|17|Graditur ad vitam, qui custodit disciplinam;qui autem increpationes relinquit, errat.
PROV|10|18|Abscondunt odium labia mendacia;qui profert contumeliam, insipiens est.
PROV|10|19|In multiloquio non deerit peccatum;qui autem moderatur labia sua, prudentissimus est.
PROV|10|20|Argentum electum lingua iusti,cor autem impiorum pro nihilo.
PROV|10|21|Labia iusti erudiunt plurimos;qui autem indocti sunt, in cordis egestate morientur.
PROV|10|22|Benedictio Domini divites facit,nec addet ei labor quidquam.
PROV|10|23|Quasi per risum stultus operatur scelus,sapientia autem est viro prudentiae.
PROV|10|24|Quod timet impius, veniet super eum;desiderium suum iustis dabitur.
PROV|10|25|Quasi tempestas transiens non erit impius,iustus autem quasi fundamentum sempiternum.
PROV|10|26|Sicut acetum dentibus et fumus oculis,sic piger his, qui miserunt eum.
PROV|10|27|Timor Domini apponet dies,et anni impiorum breviabuntur.
PROV|10|28|Exspectatio iustorum laetitia,spes autem impiorum peribit.
PROV|10|29|Fortitudo simplici via Dominiet ruina his, qui operantur malum.
PROV|10|30|Iustus in aeternum non commovebitur,impii autem non habitabunt super terram.
PROV|10|31|Os iusti germinabit sapientiam,lingua prava abscindetur.
PROV|10|32|Labia iusti considerant placita,et os impiorum perversa.
PROV|11|1|Statera dolosa abominatio est apud Dominum,et pondus aequum voluntas eius.
PROV|11|2|Venit superbia, veniet et contumelia;apud humiles autem sapientia.
PROV|11|3|Simplicitas iustorum diriget eos,et supplantatio perversorum vastabit illos.
PROV|11|4|Non proderunt divitiae in die ultionis,iustitia autem liberabit a morte.
PROV|11|5|Iustitia simplicis diriget viam eius,et in impietate sua corruet impius.
PROV|11|6|Iustitia rectorum liberabit eos,et in insidiis suis capientur iniqui.
PROV|11|7|Mortuo homine impio, nulla erit ultra spes;et exspectatio divitiarum peribit.
PROV|11|8|Iustus de angustia liberatus est,et tradetur impius pro eo.
PROV|11|9|Simulator ore decipit amicum suum,iusti autem liberabuntur scientia.
PROV|11|10|In bonis iustorum exsultabit civitas,et in perditione impiorum erit laudatio.
PROV|11|11|Benedictione iustorum exaltabitur civitaset ore impiorum subvertetur.
PROV|11|12|Qui despicit amicum suum, indigens corde est,vir autem prudens tacebit.
PROV|11|13|Qui ambulat susurrans, revelat arcana;qui autem fidelis est animi, celat commissum.
PROV|11|14|Ubi non adsunt dispositiones, populus corruet;salus autem, ubi multa consilia.
PROV|11|15|Affligetur malo, qui fidem facit pro extraneo;qui autem odit sponsores, securus erit.
PROV|11|16|Mulier gratiosa inveniet gloriam,et robusti habebunt divitias.
PROV|11|17|Benefacit animae suae vir misericors;qui autem crudelis est, carnem suam affligit.
PROV|11|18|Impius facit opus fallax,seminanti autem iustitiam merces fidelis.
PROV|11|19|Firmus in iustitia praeparat vitam,et sectator malorum mortem.
PROV|11|20|Abominabile Domino cor pravum,et voluntas eius in iis, qui simpliciter ambulant.
PROV|11|21|Manus in manu, non erit impunitus malus,semen autem iustorum salvabitur.
PROV|11|22|Circulus aureus in naribus suismulier pulchra et fatua.
PROV|11|23|Desiderium iustorum omne bonum est,praestolatio impiorum furor.
PROV|11|24|Alii dividunt propria et ditiores fiunt,alii parciores iusto semper in egestate sunt.
PROV|11|25|Anima, quae benedicit, impinguabitur;et, qui inebriat, ipse quoque inebriatur.
PROV|11|26|Qui abscondit frumenta, maledicetur in populis,benedictio autem super caput vendentium.
PROV|11|27|Qui instanter quaerit bonum, quaerit beneplacitum;qui autem investigator malorum est, haec advenient ei.
PROV|11|28|Qui confidit in divitiis suis, corruet,iusti autem quasi virens folium germinabunt.
PROV|11|29|Qui conturbat domum suam, possidebit ventos;et, qui stultus est, serviet sapienti.
PROV|11|30|Fructus iusti lignum vitae;et suscipit animas, qui sapiens est.
PROV|11|31|Si iustus in terra rependitur,quanto magis impius et peccator.
PROV|12|1|Qui diligit disciplinam, diligit scientiam;qui autem odit increpationes, insipiens est.
PROV|12|2|Qui bonus est, hauriet gratiam a Domino,virum autem versutum ipse condemnabit.
PROV|12|3|Non roborabitur homo ex impietate,et radix iustorum non commovebitur.
PROV|12|4|Mulier diligens corona est viro suo,et quasi putredo in ossibus eius, quae est inhonesta.
PROV|12|5|Cogitationes iustorum iudicia,et consilia impiorum fraudulentia.
PROV|12|6|Verba impiorum insidiantur sanguini,os iustorum liberabit eos.
PROV|12|7|Subvertuntur impii et iam non sunt,domus autem iustorum permanebit.
PROV|12|8|Ad doctrinam suam laudabitur vir;qui autem perversus corde est, patebit contemptui.
PROV|12|9|Melior est pauper, qui ministrat sibi,quam gloriosus et indigens pane.
PROV|12|10|Curat iustus iumentorum suorum animas,viscera autem impiorum crudelia.
PROV|12|11|Qui operatur terram suam, satiabitur panibus;qui autem sectatur vana, vecors est.
PROV|12|12|Desiderat impius laqueum pessimorum,radix autem iustorum proficiet.
PROV|12|13|Propter peccata labiorum irretitur malus,effugiet autem iustus de angustia.
PROV|12|14|De fructu oris sui unusquisque replebitur bonis,et iuxta opera manuum suarum retribuetur ei.
PROV|12|15|Via stulti recta in oculis eius;qui autem sapiens est, audit consilia.
PROV|12|16|Fatuus statim indicat iram suam,dissimulat autem iniuriam callidus.
PROV|12|17|Qui spirat veritatem, index iustitiae est,testis autem mendax, fraudulentiae.
PROV|12|18|Est qui temere loquitur et quasi gladio pungit,lingua autem sapientium sanitas est.
PROV|12|19|Labium veritatis firmum erit in perpetuum,ad momentum autem lingua mendacii.
PROV|12|20|Dolus in corde cogitantium mala;qui autem pacis ineunt consilia, sequitur eos gaudium.
PROV|12|21|Nulla calamitas obveniet iusto,impii autem replebuntur malo.
PROV|12|22|Abominatio est Domino labia mendacia,qui autem fideliter agunt, placent ei.
PROV|12|23|Homo versutus celat scientiam,et cor insipientium provocat stultitiam.
PROV|12|24|Manus fortium dominabitur,quae autem remissa est, tributis serviet.
PROV|12|25|Maeror in corde viri humiliabit illum,et sermo bonus laetificabit eum.
PROV|12|26|In rectum ducit amicum iustus,iter autem impiorum decipiet eos.
PROV|12|27|Non assabit ignavia praedam suam,sed substantia pretiosa erit viro industrio.
PROV|12|28|In semita iustitiae vita,est autem etiam iter apertum ad mortem.
PROV|13|1|Filius sapiens disciplina patris;qui autem illusor est, non audit, cum arguitur.
PROV|13|2|De fructu oris sui homo satiabitur bonis,anima autem praevaricatorum violentia.
PROV|13|3|Qui custodit os suum, custodit animam suam;qui autem incautus est eloquio, ruina est ei.
PROV|13|4|Vult et non habet piger,anima autem operantium impinguabitur.
PROV|13|5|Verbum mendax iustus detestabitur,impius autem confundit et dehonestat.
PROV|13|6|Iustitia custodit innocentem in via,impietas autem peccatorem supplantat.
PROV|13|7|Est qui quasi dives habetur, cum nihil habeat;et est qui quasi pauper, cum in multis divitiis sit.
PROV|13|8|Redemptio animae viri divitiae suae;qui autem pauper est, increpationem non sustinet.
PROV|13|9|Lux iustorum laetificat,lucerna autem impiorum exstinguetur.
PROV|13|10|Inter superbos tantum iurgia sunt,et apud humiles sapientia.
PROV|13|11|Substantia festinata minuetur;qui autem colligit manu, multiplicat.
PROV|13|12|Spes, quae differtur, affligit animam,lignum vitae desiderium veniens.
PROV|13|13|Qui contemnit verbum, ipse se obligat;qui autem timet praeceptum, retribuetur ei.
PROV|13|14|Lex sapientis fons vitae,ut declinet a laqueis mortis.
PROV|13|15|Intellegentia bona dabit gratiam,in itinere infidelium vorago.
PROV|13|16|Omnis astutus agit cum consilio;qui autem fatuus est, aperit stultitiam.
PROV|13|17|Nuntius impius cadet in malum,legatus autem fidelis sanitas.
PROV|13|18|Egestas et ignominia ei, qui deserit disciplinam;qui autem acquiescit arguenti, glorificabitur.
PROV|13|19|Desiderium, si compleatur, delectat animam;detestantur stulti fugere mala.
PROV|13|20|Qui cum sapientibus graditur, sapiens erit;amicus stultorum malus efficietur.
PROV|13|21|Peccatores persequitur malum,et iustis retribuentur bona.
PROV|13|22|Bonus relinquit heredes filios et nepotes;et custoditur iusto substantia peccatoris.
PROV|13|23|Multi cibi in novalibus pauperum,et est qui perit, deficiente iudicio.
PROV|13|24|Qui parcit virgae, odit filium suum;qui autem diligit illum, instanter erudit.
PROV|13|25|Iustus comedit et replet animam suam,venter autem impiorum insaturabilis.
PROV|14|1|Sapientia mulierum aedificat domum suam,insipientia eam manibus destruet.
PROV|14|2|Ambulans recto itinere timet Deum;despicit illum, qui infami graditur via.
PROV|14|3|In ore stulti virga superbiae,labia autem sapientium custodiunt eos.
PROV|14|4|Ubi non sunt boves, praesepe vacuum est;plurimae autem segetes in fortitudine bovis.
PROV|14|5|Testis fidelis non mentitur,profert autem mendacium dolosus testis.
PROV|14|6|Quaerit derisor sapientiam et non invenit;doctrina prudentibus facilis.
PROV|14|7|Cede coram viro stulto,quia nescies labia prudentiae.
PROV|14|8|Sapientia callidi est intellegere viam suam,et imprudentia stultorum errans.
PROV|14|9|Stulti parvipendent peccatum,et inter iustos morabitur gratia.
PROV|14|10|Cor novit amaritudinem animae suae,in gaudio eius non miscebitur extraneus.
PROV|14|11|Domus impiorum delebitur,tabernacula vero iustorum germinabunt.
PROV|14|12|Est via, quae videtur homini recta,novissima autem eius deducunt ad mortem.
PROV|14|13|Etiam in risu cor dolore miscebitur,et extrema gaudii luctus occupat.
PROV|14|14|Viis suis replebitur stultus,et super eum erit vir bonus.
PROV|14|15|Simplex credit omni verbo,astutus considerat gressus suos.
PROV|14|16|Sapiens timet et declinat a malo,stultus transilit et confidit.
PROV|14|17|Impatiens operabitur stultitiam,et vir versutus odiosus est.
PROV|14|18|Possidebunt simplices stultitiam,et astuti coronabuntur scientia.
PROV|14|19|Procumbunt mali ante bonos,et impii ante portas iustorum.
PROV|14|20|Etiam proximo suo pauper odiosus erit,amici vero divitum multi.
PROV|14|21|Qui despicit proximum suum, peccat;qui autem miseretur pauperis, beatus erit.
PROV|14|22|Nonne errant, qui operantur malum?Misericordia et veritas iis, qui praeparant bona.
PROV|14|23|In omni labore erit abundantia;verbum autem labiorum tendit tantummodo ad egestatem.
PROV|14|24|Corona sapientium divitiae eorum,fatuitas stultorum fatuitas est.
PROV|14|25|Liberat animas testis fidelis,et profert mendacia versipellis.
PROV|14|26|In timore Domini fiducia fortis,et filiis eius erit spes.
PROV|14|27|Timor Domini fons vitae,declinans a laqueis mortis.
PROV|14|28|In multitudine populi dignitas regis,et in paucitate plebis ruina principis.
PROV|14|29|Qui patiens est, multa gubernatur prudentia;qui autem impatiens est, exaltat stultitiam.
PROV|14|30|Vita carnium sanitas cordis,putredo ossium invidia.
PROV|14|31|Qui calumniatur egentem, exprobrat Factori eius;honorat autem eum, qui miseretur pauperis.
PROV|14|32|In malitia sua impelletur impius,sperat autem iustus in integritate sua.
PROV|14|33|In corde prudentis requiescit sapientia,at in medio stultorum agnoscetur?
PROV|14|34|Iustitia elevat gentem,vituperium autem populorum est peccatum.
PROV|14|35|Acceptus est regi minister intellegens,et iracundia ei, qui turpiter agit.
PROV|15|1|Responsio mollis frangit iram,sermo durus suscitat furorem.
PROV|15|2|Lingua sapientium stillat scientiam,os fatuorum ebullit stultitiam.
PROV|15|3|In omni loco oculi Dominicontemplantur malos et bonos.
PROV|15|4|Lingua placabilis lignum vitae,sed obliquitas in ea conteret spiritum.
PROV|15|5|Stultus irridet disciplinam patris sui;qui autem custodit increpationes, astutior fiet.
PROV|15|6|In domo iusti divitiae plurimae,et in fructibus impii conturbatio.
PROV|15|7|Labia sapientium disseminabunt scientiam;cor stultorum non rectum erit.
PROV|15|8|Victimae impiorum abominabiles Domino;vota iustorum grata sunt ei.
PROV|15|9|Abominatio est Domino via impii;qui sequitur iustitiam, diligetur.
PROV|15|10|Admonitio mala deserenti viam;qui increpationes odit, morietur.
PROV|15|11|Infernus et Perditio coram Domino,quanto magis corda filiorum hominum!
PROV|15|12|Non amat derisor eum, qui se corripit,nec ad sapientes graditur.
PROV|15|13|Cor gaudens exhilarat faciem,in maerore animi deicitur spiritus.
PROV|15|14|Cor sapientis quaerit doctrinam,et os stultorum pascitur stultitia.
PROV|15|15|Omnes dies pauperis mali;hilaris autem corde quasi iuge convivium.
PROV|15|16|Melius est parum cum timore Dominiquam thesauri magni cum sollicitudine.
PROV|15|17|Melius est demensum holerum cum caritatequam vitulus saginatus cum odio.
PROV|15|18|Vir iracundus provocat rixas;qui patiens est, mitigat lites.
PROV|15|19|Iter pigrorum quasi saepes spinarum,via sollertium complanata.
PROV|15|20|Filius sapiens laetificat patrem,et stultus homo despicit matrem suam.
PROV|15|21|Stultitia gaudium sensu carenti;et vir prudens dirigit gressus suos.
PROV|15|22|Dissipantur cogitationes, ubi non est consilium;ubi vero sunt plures consiliarii, confirmantur.
PROV|15|23|Laetatur homo in responsione oris sui,et sermo opportunus est optimus.
PROV|15|24|Semita vitae sursum est viro erudito,ut declinet de inferno deorsum.
PROV|15|25|Domum superborum demolietur Dominuset firmos faciet terminos viduae.
PROV|15|26|Abominatio Domini cogitationes malae,et purus sermo pulcherrimus.
PROV|15|27|Conturbat domum suam, qui sectatur avaritiam;qui autem odit munera, vivet.
PROV|15|28|Mens iusti meditatur, ut respondeat;os impiorum redundat malis.
PROV|15|29|Longe est Dominus ab impiiset orationes iustorum exaudiet.
PROV|15|30|Lux oculorum laetificat animam,fama bona impinguat ossa.
PROV|15|31|Auris, quae audit increpationes vitae,in medio sapientium commorabitur.
PROV|15|32|Qui abicit disciplinam, despicit animam suam;qui autem acquiescit increpationibus, possessor est cordis.
PROV|15|33|Timor Domini disciplina sapientiae,et gloriam praecedit humilitas.
PROV|16|1|Hominis est animum praeparare,et Domini est responsio linguae.
PROV|16|2|Omnes viae hominis purae sunt oculis eius,spirituum ponderator est Dominus.
PROV|16|3|Revela Domino opera tua,et dirigentur cogitationes tuae.
PROV|16|4|Universa secundum proprium finem operatus est Dominus;impium quoque ad diem malum.
PROV|16|5|Abominatio Domini est omnis arrogans;manus in manu, non erit innocens.
PROV|16|6|Misericordia et veritate redimitur iniquitas,et in timore Domini declinatur a malo.
PROV|16|7|Cum placuerint Domino viae hominis,inimicos quoque eius convertet ad pacem.
PROV|16|8|Melius est parum cum iustitiaquam multi fructus sine aequitate.
PROV|16|9|Cor hominis disponit viam suam,sed Domini est dirigere gressus eius.
PROV|16|10|Divinatio in labiis regis,in iudicio non errabit os eius.
PROV|16|11|Pondus et statera iusta Domini sunt,et opera eius omnes lapides sacculi.
PROV|16|12|Abominantur reges agere impie,quoniam iustitia firmatur solium.
PROV|16|13|Voluntas regum labia iusta;qui recta loquitur, diligetur.
PROV|16|14|Indignatio regis nuntii mortis,et vir sapiens placabit eam.
PROV|16|15|In lumine vultus regis vita,et voluntas eius quasi imber serotinus.
PROV|16|16|Possidere sapientiam quanto melius est auro;et acquirere prudentiam pretiosius est argento.
PROV|16|17|Semita iustorum declinare a malo;custos animae suae, qui servat viam suam.
PROV|16|18|Contritionem praecedit superbia,et ante ruinam exaltatio spiritus.
PROV|16|19|Melius est humiliari cum mitibusquam dividere spolia cum superbis.
PROV|16|20|Eruditus in verbo reperiet bona;et, qui sperat in Domino, beatus est.
PROV|16|21|Qui sapiens est corde, appellabitur prudens;et dulcedo labiorum addet doctrinam.
PROV|16|22|Fons vitae eruditio possidentis;poena stultorum stultitia.
PROV|16|23|Cor sapientis erudiet os eiuset labiis eius addet doctrinam.
PROV|16|24|Favus mellis composita verba,dulcedo animae et sanitas ossium.
PROV|16|25|Est via, quae videtur homini recta,et novissima eius ducunt ad mortem.
PROV|16|26|Anima laborantis laborat sibi,quia compulit eum os suum.
PROV|16|27|Vir impius fodit malum,et in labiis eius quasi ignis ardens.
PROV|16|28|Homo perversus suscitat lites,et mussitator separat familiares.
PROV|16|29|Vir iniquus lactat amicum suumet ducit eum per viam non bonam.
PROV|16|30|Qui attonitis oculis cogitat prava,comprimens labia sua perficit malum.
PROV|16|31|Corona dignitatis canities,quae in viis iustitiae reperietur.
PROV|16|32|Melior est patiens viro forti,et, qui dominatur animo suo, expugnatore urbium.
PROV|16|33|Sortes mittuntur in sinum,sed a Domino temperantur.
PROV|17|1|Melior est buccella sicca cum pacequam domus plena victimis cum iurgio.
PROV|17|2|Servus sapiens dominabitur filiis inhonestiset inter fratres hereditatem dividet.
PROV|17|3|Sicut igne probatur argentum et aurum camino,ita corda probat Dominus.
PROV|17|4|Malus oboedit labio iniquo,et fallax obtemperat linguae mendaci.
PROV|17|5|Qui despicit pauperem, exprobrat Factori eius;et, qui in ruina laetatur alterius, non erit impunitus.
PROV|17|6|Corona senum filii filiorum,et gloria filiorum patres eorum.
PROV|17|7|Non decent stultum verba composita,nec principem labium mentiens.
PROV|17|8|Gemma gratissima munus in oculis domini eius;quocumque se verterit, prospere aget.
PROV|17|9|Qui celat delictum, quaerit amicitias;qui sermone repetit, separat foederatos.
PROV|17|10|Plus proficit correptio apud prudentemquam centum plagae apud stultum.
PROV|17|11|Semper iurgia quaerit malus;angelus autem crudelis mittetur contra eum.
PROV|17|12|Expedit magis ursae occurrere, raptis fetibus,quam fatuo confidenti in stultitia sua.
PROV|17|13|Qui reddit mala pro bonis,non recedet malum de domo eius.
PROV|17|14|Aquarum proruptio initium est iurgiorum;et, antequam exacerbetur contentio, desere.
PROV|17|15|Qui iustificat impium et qui condemnat iustum,abominabilis est uterque apud Dominum.
PROV|17|16|Ad quid pretium in manu stulti?Ad emendam sapientiam, cum careat corde?
PROV|17|17|Omni tempore diligit, qui amicus est,et frater ad angustiam natus est.
PROV|17|18|Stultus homo iungit manus,cum spoponderit pro amico suo.
PROV|17|19|Qui diligit delictum, diligit rixas;et, qui exaltat ostium, quaerit effracturam.
PROV|17|20|Qui perversi cordis est, non inveniet bonum;et, qui vertit linguam, incidet in malum.
PROV|17|21|Qui generat stultum, maerorem generat sibi,sed nec pater in fatuo laetabitur.
PROV|17|22|Animus gaudens aetatem floridam facit,spiritus tristis exsiccat ossa.
PROV|17|23|Munera de sinu impius accipit,ut pervertat semitas iudicii.
PROV|17|24|In facie prudentis lucet sapientia,oculi stultorum in finibus terrae.
PROV|17|25|Ira patris filius stultuset dolor matris, quae genuit eum.
PROV|17|26|Non est bonum multam inferre iustonec percutere principem contra rectitudinem.
PROV|17|27|Qui moderatur sermones suos, novit scientiam,et lenis spiritu est vir prudens.
PROV|17|28|Stultus quoque, si tacuerit, sapiens reputabituret, si compresserit labia sua, intellegens.
PROV|18|1|Occasiones quaerit, qui vult recedere ab amico;omni consilio exacerbatur.
PROV|18|2|Non delectatur stultus prudentiased in revelatione cordis sui.
PROV|18|3|Cum venerit impius, veniet et contemptio,et cum ignominia opprobrium.
PROV|18|4|Aqua profunda verba ex ore viri,et torrens redundans fons sapientiae.
PROV|18|5|Accipere personam impii non est bonum,ut declines iustum in iudicio.
PROV|18|6|Labia stulti miscent se rixis,et os eius plagas provocat.
PROV|18|7|Os stulti ruina eius,et labia ipsius laqueus animae eius.
PROV|18|8|Verba susurronis quasi dulcia,et ipsa perveniunt usque ad interiora ventris.
PROV|18|9|Qui mollis et dissolutus est in opere suo,frater est viri dissipantis.
PROV|18|10|Turris fortissima nomen Domini;ad ipsum currit iustus et exaltabitur.
PROV|18|11|Substantia divitis urbs roboris eiuset quasi murus excelsus in cogitatione eius.
PROV|18|12|Antequam conteratur, exaltatur cor hominis;et, antequam glorificetur, humiliatur.
PROV|18|13|Qui prius respondet quam audiat,stultitia est ei et contumelia.
PROV|18|14|Spiritus viri sustentat imbecillitatem suam;spiritum vero confractum, quis poterit sustinere?
PROV|18|15|Cor prudens possidebit scientiam,et auris sapientium quaerit doctrinam.
PROV|18|16|Donum hominis dilatat viam eiuset ante principes deducit eum.
PROV|18|17|Qui prior in contentione loquitur, putatur iustus;venit amicus eius et arguet eum.
PROV|18|18|Lites comprimit sorset inter potentes quoque diiudicat.
PROV|18|19|Frater, qui offenditur, durior est civitate firma,et lites quasi vectes urbium.
PROV|18|20|De fructu oris viri replebitur venter eius,et genimina labiorum ipsius saturabunt eum.
PROV|18|21|Mors et vita in manu linguae;qui diligunt eam, comedent fructus eius.
PROV|18|22|Qui invenit mulierem bonam, invenit bonumet hausit gratiam a Domino.
PROV|18|23|Cum obsecrationibus loquetur pauper,et dives effabitur rigide.
PROV|18|24|Vir cum amicis concuti potest,sed est amicus, qui adhaereat magis quam frater.
PROV|19|1|Melior est pauper, qui ambulat in simplicitate sua,quam qui torquet labia et est insipiens.
PROV|19|2|Ubi non est scientia animae, non est bonum;et, qui festinus est pedibus, offendit.
PROV|19|3|Stultitia hominis supplantat gressus eius,et contra Deum fervet animo suo.
PROV|19|4|Divitiae addunt amicos plurimos;pauper autem ab amico suo separatur.
PROV|19|5|Testis falsus non erit impunitus;et, qui mendacia loquitur, non effugiet.
PROV|19|6|Multi blandiuntur faciei potentis,et omnes amici sunt dona tribuenti.
PROV|19|7|Omnes fratres hominis pauperis oderunt eum,insu7per et amici procul recesserunt ab eo;qui tantum verba sectatur, nihil habebit.
PROV|19|8|Qui autem possessor est mentis, diligit animam suam,et custos prudentiae inveniet bona.
PROV|19|9|Falsus testis non erit impunitus;et, qui loquitur mendacia, peribit.
PROV|19|10|Non decent stultum deliciae,nec servum dominari principibus.
PROV|19|11|Doctrina viri mitigat iram eius,et gloria eius est iniqua praetergredi.
PROV|19|12|Sicut fremitus leonis ita et regis ira,et sicut ros super herbam ita et gratia eius.
PROV|19|13|Calamitas patris filius stultus;et tecta iugiter perstillantia litigiosa mulier.
PROV|19|14|Domus et divitiae hereditas patrum,a Domino autem uxor prudens.
PROV|19|15|Pigredo immittit soporem,et anima dissoluta esuriet.
PROV|19|16|Qui custodit mandatum, custodit animam suam;qui autem neglegit viam suam, mortificabitur.
PROV|19|17|Feneratur Domino, qui miseretur pauperis,et vicissitudinem suam reddet ei.
PROV|19|18|Erudi filium tuum, dum spes est;ad interfectionem autem eius ne ponas animam tuam.
PROV|19|19|Qui impatiens est, sustinebit multam;et, si eum abripere vis, aliud appones.
PROV|19|20|Audi consilium et suscipe disciplinam,ut sis sapiens in novissimis tuis.
PROV|19|21|Multae cogitationes in corde viri,voluntas autem Domini permanebit.
PROV|19|22|Desiderabile in homine est misericordia eius;et melior est pauper quam vir mendax.
PROV|19|23|Timor Domini ad vitam,et in plenitudine commorabitur absque visitatione mali.
PROV|19|24|Abscondit piger manum suam in catinonec ad os suum applicat eam.
PROV|19|25|Derisore flagellato vel parvulus sapientior erit;si autem corripueris sapientem, intelleget disciplinam.
PROV|19|26|Qui affligit patrem et fugat matrem,filius inhonestus et ignominiosus.
PROV|19|27|Acquiesce, fili, ut audias doctrinamnec erres a sermonibus scientiae.
PROV|19|28|Testis iniquus deridet iudicium,et os impiorum devorat iniquitatem.
PROV|19|29|Paratae sunt derisoribus virgae,et plagae stultorum corporibus.
PROV|20|1|Luxuriosa res vinum, et tumultuosa sicera;quicumque his delectatur, non erit sapiens.
PROV|20|2|Sicut rugitus leonis ita et terror regis:qui provocat eum, peccat in animam suam.
PROV|20|3|Honor est homini separari a contentionibus;omnes autem stulti miscentur contumeliis.
PROV|20|4|Propter frigus piger arare noluit;mendicabit ergo aestate, et non dabitur illi.
PROV|20|5|Sicut aqua profunda consilium in corde viri,sed homo sapiens exhauriet illud.
PROV|20|6|Multi homines misericordes vocantur;virum autem fidelem quis inveniet?
PROV|20|7|Iustus, qui ambulat in simplicitate sua,beatos post se filios derelinquet.
PROV|20|8|Rex, qui sedet in solio iudicii,dissipat omne malum intuitu suo.
PROV|20|9|Quis potest dicere: " Mundavi cor meum,purus sum a peccato "?
PROV|20|10|Pondus et pondus, mensura et mensura,utrumque abominabile est apud Dominum.
PROV|20|11|Ex studiis suis intellegitur puer,si munda et recta sint opera eius.
PROV|20|12|Aurem audientem et oculum videntem,Dominus fecit utrumque.
PROV|20|13|Noli diligere somnum, ne te egestas opprimat;aperi oculos tuos et saturare panibus.
PROV|20|14|" Malum est, malum est! " dicit omnis emptoret, cum recesserit, tunc gloriabitur.
PROV|20|15|Est aurum et multitudo gemmarumet vas pretiosum labia scientiae.
PROV|20|16|Tolle vestimentum eius, quia fideiussor exstitit alieni,et pro extraneis aufer pignus ab eo.
PROV|20|17|Suavis est homini panis mendacii,et postea implebitur os eius calculo.
PROV|20|18|Cogitationes consiliis firmantur,et dispensationibus tractanda sunt bella.
PROV|20|19|Ei, qui revelat mysteria et calumniaturet dilatat labia sua, ne commiscearis.
PROV|20|20|Qui maledicit patri suo et matri,exstinguetur lucerna eius in mediis tenebris.
PROV|20|21|Hereditas, ad quam festinatur in principio,in novissimo benedictione carebit.
PROV|20|22|Ne dicas: " Reddam malum ";exspecta Dominum, et liberabit te.
PROV|20|23|Abominatio est apud Dominum pondus et pondus;statera dolosa non est bona in oculis eius.
PROV|20|24|A Domino diriguntur gressus viri;quis autem hominum intellegere potest viam suam?
PROV|20|25|Laqueus est homini inconsulte dicere: " Sanctum! "et post vota retractare.
PROV|20|26|Ventilat impios rex sapienset incurvat super eos rotam.
PROV|20|27|Lucerna Domini spiraculum hominis,quae investigat omnia secreta ventris.
PROV|20|28|Misericordia et veritas custodiunt regem,et roboratur clementia thronus eius.
PROV|20|29|Ornamentum iuvenum fortitudo eorum,et honor senum canities.
PROV|20|30|Livor vulneris absterget mala,et plagae in secretioribus ventris.
PROV|21|1|Sicut rivi aquarum cor regis in manu Domini:quocumque voluerit, inclinabit illud.
PROV|21|2|Omnis via viri recta sibi videtur;appendit autem corda Dominus.
PROV|21|3|Facere misericordiam et iudiciummagis placet Domino quam victimae.
PROV|21|4|Exaltatio oculorum et dilatatio cordis,lucerna impiorum: peccatum.
PROV|21|5|Cogitationes sollertis semper in abundantiam;omnis autem festinus semper in egestate est.
PROV|21|6|Qui congregat thesauros lingua mendacii,vento impingetur ad laqueos mortis.
PROV|21|7|Violentia impiorum detrahet eos,quia noluerunt facere iudicium.
PROV|21|8|Perversa via viri aliena est;qui autem mundus est, rectum opus eius.
PROV|21|9|Melius est sedere in angulo domatisquam cum muliere litigiosa et in domo communi.
PROV|21|10|Anima impii desiderat malum;non miserebitur proximo suo.
PROV|21|11|Multato derisore sapientior erit parvulus;et, si instruatur sapiens, sumet scientiam.
PROV|21|12|Excogitat Iustus de domo impii,ut praecipitet impios in malum.
PROV|21|13|Qui obturat aurem suam ad clamorem pauperis,et ipse clamabit, et non exaudietur.
PROV|21|14|Munus absconditum exstinguit iras,et donum in sinu indignationem maximam.
PROV|21|15|Gaudium iusto est facere iudicium,et ruina operantibus iniquitatem.
PROV|21|16|Vir, qui erraverit a via prudentiae,in coetu umbrarum commorabitur.
PROV|21|17|Qui diligit convivia, in egestate erit;qui amat vinum et pinguia, non ditabitur.
PROV|21|18|Redemptio pro iusto impius,et pro rectis iniquus.
PROV|21|19|Melius est habitare in terra desertaquam cum muliere rixosa et iracunda.
PROV|21|20|Thesaurus desiderabilis et pinguis in habitaculo sapientis,et imprudens homo dissipabit illum.
PROV|21|21|Qui sequitur iustitiam et misericordiam,inveniet vitam et iustitiam et gloriam.
PROV|21|22|Civitatem fortium ascendit sapienset destruit robur fiduciae eius.
PROV|21|23|Qui custodit os suum et linguam suam,custodit ab angustiis animam suam.
PROV|21|24|Superbus et arrogans vocatur derisor,qui operatur in ira superbiae.
PROV|21|25|Desideria occidunt pigrum;noluerunt enim quidquam manus eius operari:
PROV|21|26|tota die concupiscit et desiderat;qui autem iustus est, tribuet et non parcit.
PROV|21|27|Hostiae impiorum abominabiles,eo magis quia offeruntur ex scelere.
PROV|21|28|Testis mendax peribit;vir oboediens loquetur in victoriam.
PROV|21|29|Vir impius obfirmat vultum suum;qui autem rectus est, corrigit viam suam.
PROV|21|30|Non est sapientia, non est prudentia,non est consilium contra Dominum.
PROV|21|31|Equus paratur ad diem belli,Dominus autem salutem tribuit.
PROV|22|1|Melius est nomen bonum quam divitiae multae,super argentum et aurum gratia bona.
PROV|22|2|Dives et pauper obviaverunt sibi:utriusque operator est Dominus.
PROV|22|3|Callidus vidit malum et abscondit se;simplices pertransierunt et afflicti sunt damno.
PROV|22|4|Praemium modestiae timor Domini,divitiae et gloria et vita.
PROV|22|5|Spinae et laquei in via perversi,custos autem animae suae longe recedit ab eis.
PROV|22|6|Institue adulescentem iuxta viam suam;etiam cum senuerit, non recedet ab ea.
PROV|22|7|Dives pauperibus imperat;et, qui accipit mutuum, servus est fenerantis.
PROV|22|8|Qui seminat iniquitatem, metet malaet virga irae suae consummabitur.
PROV|22|9|Qui bono oculo est, benedicetur,de panibus enim suis dedit pauperi.
PROV|22|10|Eice derisorem, et exibit cum eo iurgium;cessabuntque causae et contumeliae.
PROV|22|11|Qui diligit cordis munditiam,propter gratiam labiorum suorum habebit amicum regem.
PROV|22|12|Oculi Domini custodiunt scientiam,et supplantantur verba iniqui.
PROV|22|13|Dicit piger: " Leo est foris,in medio platearum occidendus sum ".
PROV|22|14|Fovea profunda os alienae;cui iratus est Dominus, incidet in eam.
PROV|22|15|Stultitia colligata est in corde pueri,et virga disciplinae fugabit eam.
PROV|22|16|Opprimis pauperem? Ipse augebit divitias suas.Donas ditiori? Ipse egebis.
PROV|22|17|Inclina aurem tuam et audi verba sapientium,appone autem cor ad doctrinam meam,
PROV|22|18|quia pulchra erunt, cum servaveris ea in ventre tuo,et redundabunt in labiis tuis.
PROV|22|19|Ut sit in Domino fiducia tua,ostendi ea tibi hodie.
PROV|22|20|Nonne descripsi ea tibi nudiustertiusin cogitationibus et scientia,
PROV|22|21|ut ostenderem tibi firmitatem verborum veritatis,ut respondeas illi, qui misit te?
PROV|22|22|Non facias violentiam pauperi, quia pauper est,neque conteras egenum in porta,
PROV|22|23|quia iudicabit Dominus causam eorum,et anima spoliabit spoliatores.
PROV|22|24|Noli esse amicus homini iracundoneque ambules cum viro furioso,
PROV|22|25|ne forte discas semitas eiuset sumas scandalum animae tuae.
PROV|22|26|Noli esse cum his, qui iungunt manus suaset qui vades se offerunt pro debitis:
PROV|22|27|si enim non habes unde restituas,quid causae est ut tollat lectum tuum subter te?
PROV|22|28|Ne transferas terminos antiquos,quos posuerunt patres tui.
PROV|22|29|Vidisti virum velocem in opere suo:coram regibus stabit nec erit ante ignobiles.
PROV|23|1|Quando sederis, ut comedas cum principe,diligenter attende, quae apposita sunt ante faciem tuam,
PROV|23|2|et statue cultrum in gutture tuo,si avidus es.
PROV|23|3|Ne desideres de cibis eius,quia est panis mendacii.
PROV|23|4|Noli laborare, ut diteris,sed in prudentia tua acquiesce.
PROV|23|5|Si erigas oculos tuos ad opes, iam non sunt;quia facient sibi pennas quasi aquilae et volabunt in caelum.
PROV|23|6|Ne comedas cum homine invidoet ne desideres cibos eius;
PROV|23|7|quoniam sicut aestimavit in animo suo,ita ipse est. Comede et bibe " dicet tibi,et mens eius non est tecum.
PROV|23|8|Buccellam, quam comederas, evomeset perdes pulchros sermones tuos.
PROV|23|9|In auribus insipientium ne loquaris,quia despicient doctrinam eloquii tui.
PROV|23|10|Ne attingas terminos viduaeet agrum pupillorum ne introeas:
PROV|23|11|redemptor enim illorum fortis est,et ipse iudicabit contra te causam illorum.
PROV|23|12|Introduc ad doctrinam cor tuumet aures tuas ad verba scientiae.
PROV|23|13|Noli subtrahere a puero disciplinam;si enim percusseris eum virga, non morietur:
PROV|23|14|tu virga percuties eumet animam eius de inferno liberabis.
PROV|23|15|Fili mi, si sapiens fuerit cor tuum,gaudebit tecum et cor meum,
PROV|23|16|et exsultabunt renes mei,cum locuta fuerint rectum labia tua.
PROV|23|17|Non aemuletur cor tuum peccatores,sed in timore Domini esto tota die,
PROV|23|18|quia est tibi posteritas,et praestolatio tua non auferetur.
PROV|23|19|Audi, fili mi, et esto sapienset dirige in via animum tuum.
PROV|23|20|Noli esse in conviviis potatorumnec in comissationibus carnis,
PROV|23|21|quia vacantes potibus et comissatores consumentur,et vestietur pannis dormitatio.
PROV|23|22|Audi patrem tuum, qui genuit te,et ne contemnas, cum senuerit mater tua.
PROV|23|23|Veritatem eme et noli vendere;sapientiam eme et doctrinam et intellegentiam.
PROV|23|24|Exsultat gaudio pater iusti;qui sapientem genuit, laetabitur in eo;
PROV|23|25|gaudeat pater tuus et mater tua,et exsultet, quae genuit te.
PROV|23|26|Praebe, fili mi, cor tuum mihi,et oculi tui vias meas custodiant.
PROV|23|27|Fovea enim profunda est meretrix,et puteus angustus aliena,
PROV|23|28|nam insidiatur ipsa in via quasi latroet iniquos in hominibus addet.
PROV|23|29|Cui " Vae "? Cui " Eheu "?Cui rixae? Cui querela?Cui sine causa vulnera? Cui suffusio oculorum?
PROV|23|30|His, qui commorantur in vinoet eunt, ut scrutentur mixtum.
PROV|23|31|Ne intuearis vinum, quando flavescit,cum splenduerit in calice color eius:ingreditur blande,
PROV|23|32|sed in novissimo mordebit ut coluberet sicut regulus vulnerat.
PROV|23|33|Oculi tui videbunt extranea,et cor tuum loquetur perversa;
PROV|23|34|et eris sicut dormiens in medio mariet quasi sopitus ad malum navis:
PROV|23|35|" Verberaverunt me, sed non dolui,percusserunt me, et ego non sensi;quando evigilabo et rursus illud requiram? ".
PROV|24|1|Ne aemuleris viros malosnec desideres esse cum eis,
PROV|24|2|quia rapinas meditatur mens eorum,et perniciem labia eorum loquuntur.
PROV|24|3|Sapientia aedificabitur domus,et prudentia roborabitur.
PROV|24|4|In doctrina replebuntur cellaria,universa substantia pretiosa et pulcherrima.
PROV|24|5|Vir sapiens fortis est,et vir doctus firmat robur.
PROV|24|6|Quia cum dispositione parabis tibi bellum,et erit salus, ubi multa consilia sunt.
PROV|24|7|Excelsa stulto sapientia,in porta non aperiet os suum.
PROV|24|8|Qui cogitat mala facere,vir perniciosus vocabitur.
PROV|24|9|Cogitatio stulti peccatum est,et abominatio hominum detractor.
PROV|24|10|Si fueris lassus in die angustiae,coartabitur fortitudo tua.
PROV|24|11|Erue eos, qui ducuntur ad mortem;et, qui trahuntur ad interitum, retine.
PROV|24|12|Si dixeris: " Nesciebamus hoc ";nonne qui ponderator est cordis, ipse intellegit,et servatorem animae tuae nihil fallitreddetque homini iuxta opera sua?
PROV|24|13|Comede, fili mi, mel, quia bonum estet favum dulcissimum gutturi tuo.
PROV|24|14|Sic, scito, est sapientia animae tuae;quam cum inveneris, erit tibi posteritas,et spes tua non peribit.
PROV|24|15|Ne insidieris, o nequam, domui iustineque vastes requiem eius.
PROV|24|16|Septies enim cadet iustus et resurget;impii autem corruent in malum.
PROV|24|17|Cum ceciderit inimicus tuus, ne gaudeas,et in ruina eius ne exsultet cor tuum,
PROV|24|18|ne forte videat Dominus, et displiceat eiet auferat ab eo iram suam.
PROV|24|19|Ne succendas ira in pessimosnec aemuleris impios,
PROV|24|20|quoniam non erit posteritas maligno,et lucerna impiorum exstinguetur.
PROV|24|21|Time Dominum, fili mi, et regemet cum nova sectantibus non commiscearis,
PROV|24|22|quoniam repente consurget perditio eorum,et ruinam utriusque quis novit?
PROV|24|23|Haec quoque sapientibus:Dignoscere personam in iudicio non est bonum.
PROV|24|24|Qui dicit impio: " Iustus es ",maledicent ei populi, et detestabuntur eum tribus.
PROV|24|25|Qui vero arguunt eum, laudabuntur,et super ipsos veniet benedictio boni.
PROV|24|26|Labia deosculatur,qui recta verba respondet.
PROV|24|27|Praepara foris opus tuumet diligenter exerce illud in agro tuo,ut postea aedifices domum tuam.
PROV|24|28|Ne sis testis frustra contra proximum tuumnec decipias quemquam labiis tuis.
PROV|24|29|Ne dicas: " Quomodo fecit mihi, sic faciam ei,reddam viro secundum opus suum ".
PROV|24|30|Per agrum hominis pigri transiviet per vineam viri sensu carentis:
PROV|24|31|et ecce totum repleverant urticae,et operuerant superficiem eius spinae,et maceria lapidum destructa erat;
PROV|24|32|quod cum vidissem, posui in corde meo,vidi, didici disciplinam:
PROV|24|33|" Parum dormies, modicum dormitabis,pauxillum manus conseres, ut quiescas,
PROV|24|34|et veniet tibi quasi cursor egestas,et mendicitas quasi vir armatus ".
PROV|25|1|Hae quoque parabolae Salomonis, quas transcripse runt viri Ezechiae regis Iudae.
PROV|25|2|Gloria Dei est celare verbum,et gloria regum investigare sermonem.
PROV|25|3|Caelum prae altitudine et terra prae profunditate,et cor regum inscrutabile.
PROV|25|4|Aufer scorias de argento,et egredietur vas pro argentario.
PROV|25|5|Aufer impium de conspectu regis,et firmabitur iustitia thronus eius.
PROV|25|6|Ne gloriosus appareas coram regeet in loco magnorum ne steteris.
PROV|25|7|Melius est enim ut dicatur tibi: " Ascende huc ",quam ut humilieris coram principe.
PROV|25|8|Quae viderunt oculi tui,ne proferas in iurgio cito,quoniam quid facies postea,cum dehonestaverit te amicus tuus?
PROV|25|9|Causam tuam tracta cum amico tuoet secretum extranei ne reveles,
PROV|25|10|ne forte insultet tibi, cum audierit,et contumelia tua revocari non poterit.
PROV|25|11|Mala aurea in ornatibus argenteis,verbum prolatum in tempore suo.
PROV|25|12|Inauris aurea et margaritum fulgenssapiens, qui arguit super aurem audientem.
PROV|25|13|Sicut frigus nivis in die messis,ita legatus fidelis ei, qui misit eum:animam ipsius recreat.
PROV|25|14|Nubes et ventus et pluviae non sequentesvir gloriosus et promissa non complens.
PROV|25|15|Patientia lenietur princeps,et lingua mollis confringet ossa.
PROV|25|16|Mel invenisti? Comede, quod sufficit tibi,ne forte satiatus evomas illud.
PROV|25|17|Subtrahe pedem tuum de domo proximi tui,ne quando satiatus oderit te.
PROV|25|18|Malleus et gladius et sagitta acutahomo, qui loquitur contra proximum suum falsum testimonium.
PROV|25|19|Dens putridus et pes vacillans,qui sperat super infideli in die angustiae.
PROV|25|20|Sicut exuens pallium in die frigoris,sicut acetum in nitro,qui cantat carmina cordi tristi.
PROV|25|21|Si esurierit inimicus tuus, ciba illum;si sitierit, pota illum:
PROV|25|22|prunas enim congregabis super caput eius,et Dominus reddet tibi.
PROV|25|23|Ventus aquilo parturit pluvias,et faciem tristem lingua detrahens.
PROV|25|24|Melius est sedere in angulo domatisquam cum muliere litigiosa et in domo communi.
PROV|25|25|Aqua frigida animae sitientiet nuntius bonus de terra longinqua.
PROV|25|26|Fons turbatus pede et vena corruptaiustus cadens coram impio.
PROV|25|27|Mel nimium comedere non est bonum,nec quaestus gloriae est gloria.
PROV|25|28|Urbs diruta et absque murovir, qui non potest cohibere spiritum suum.
PROV|26|1|Quomodo nix in aestate et pluvia in messe,sic indecens est stulto gloria.
PROV|26|2|Sicut avis ad alia transvolans et hirundo volitans,sic maledictum frustra prolatum non superveniet.
PROV|26|3|Flagellum equo et camus asinoet virga dorso stultorum.
PROV|26|4|Ne respondeas stulto iuxta stultitiam suam,ne tu quoque efficiaris ei similis;
PROV|26|5|responde stulto iuxta stultitiam suam,ne sibi sapiens esse videatur.
PROV|26|6|Amputat sibi pedes et iniuriam bibit,qui mittit verba per manum stulti.
PROV|26|7|Quomodo molles claudo tibiae,sic in ore stultorum parabola.
PROV|26|8|Sicut qui celat lapidem in acervo,ita qui tribuit insipienti honorem.
PROV|26|9|Spina crescens in manu temulenti,sic parabola in ore stultorum.
PROV|26|10|Sagittarius, qui conicit ad omnia,ita qui stultum conducit et qui vagos conducit.
PROV|26|11|Sicut canis, qui revertitur ad vomitum suum,sic stultus, qui iterat stultitiam suam.
PROV|26|12|Vidisti hominem sapientem sibi videri?Magis illo spem habebit stultus.
PROV|26|13|Dicit piger: " Leaena est in via,et leo in plateis ".
PROV|26|14|Ostium vertitur in cardine suo,et piger in lectulo suo.
PROV|26|15|Abscondit piger manum in catinoet laborat, si ad os suum eam converterit.
PROV|26|16|Sapientior sibi piger videturseptem viris respondentibus sententias.
PROV|26|17|Apprehendit auribus canem,qui transiens commiscetur rixae alterius.
PROV|26|18|Sicut insanit, qui mittit sagittaset lanceas in mortem,
PROV|26|19|ita vir, qui decipit amicum suumet dicit: " Nonne ludens feci? ".
PROV|26|20|Cum defecerint ligna, exstinguetur ignis,et, susurrone subtracto, iurgia conquiescent.
PROV|26|21|Sicut carbones ad prunas et ligna ad ignem,sic homo litigiosus ad inflammandas rixas.
PROV|26|22|Verba susurronis quasi dulciaet ipsa perveniunt ad intima ventris.
PROV|26|23|Sicut argentum sordidum ornans vas fictile,sic labia levia et cor malum.
PROV|26|24|Labiis suis se dissimulabit inimicus,cum in corde tractaverit dolos:
PROV|26|25|quando mollierit vocem suam, ne credideris ei,quoniam septem abominationes sunt in corde illius;
PROV|26|26|operiet odium fraudulenter,revelabitur autem malitia eius in concilio.
PROV|26|27|Qui fodit foveam, incidet in eam;et, qui volvit lapidem, revertetur ad eum.
PROV|26|28|Lingua fallax non amat veritatem,et os lubricum operatur ruinas.
PROV|27|1|Ne glorieris in crastinumignorans, quid superventura pariat dies.
PROV|27|2|Laudet te alienus et non os tuum,extraneus et non labia tua.
PROV|27|3|Grave est saxum et onerosa arena,sed ira stulti utroque gravior.
PROV|27|4|Saevitas et erumpens furor,et coram zelo consistere quis poterit?
PROV|27|5|Melior est manifesta correptioquam amor absconditus.
PROV|27|6|Veriora sunt vulnera diligentisquam fraudulenta oscula odientis.
PROV|27|7|Anima saturata calcabit favum,et anima esuriens etiam amarum pro dulci sumet.
PROV|27|8|Sicut avis transmigrans de nido suo,sic vir errans longe a loco suo.
PROV|27|9|Unguento et ture delectatur coret dulcedine amici in consilio ex animo.
PROV|27|10|Amicum tuum et amicum patris tui ne dimiseriset domum fratris tui ne ingrediaris in die afflictionis tuae.Melior est vicinus iuxta quam frater procul.
PROV|27|11|Stude sapientiae, fili mi, et laetifica cor meum,ut possim exprobranti mihi respondere sermonem.
PROV|27|12|Astutus videns malum absconditus est;simplices transeuntes multati sunt.
PROV|27|13|Tolle vestimentum eius, qui spopondit pro extraneo,et pro alienis aufer ei pignus.
PROV|27|14|Qui benedicit proximo suo voce grandi mane consurgens,maledictio reputabitur ei.
PROV|27|15|Tecta perstillantia in die frigoriset litigiosa mulier comparantur;
PROV|27|16|qui retinet eam, quasi qui ventum teneat,et oleum dextera sua tenere reperietur.
PROV|27|17|Ferrum ferro exacuitur,et homo exacuit faciem amici sui.
PROV|27|18|Qui servat ficum, comedet fructus eius;et, qui custos est domini sui, glorificabitur.
PROV|27|19|Quomodo in aqua facies prospicit ad faciem,sic cor hominis ad hominem.
PROV|27|20|Infernus et Perditio numquam implentur,similiter et oculi hominum insatiabiles.
PROV|27|21|Quomodo probatur in conflatorio argentum et in fornace aurum,sic probatur homo ore laudantis.
PROV|27|22|Si pilo contuderis stultum in pila quasi ptisanas,non auferetur ab eo stultitia eius.
PROV|27|23|Diligenter agnosce vultum pecoris tui;appone cor tuum ad greges,
PROV|27|24|non enim habebis iugiter divitias.Num corona tribuetur in generationem et generationem?
PROV|27|25|Nudata sunt prata, et apparuerunt herbae virentes,et collecta sunt fena de montibus;
PROV|27|26|agni ad vestimentum tuum,et haedi ad agri pretium;
PROV|27|27|sufficiat tibi lac caprarum in cibum tuumet in cibum domus tuae et ad victum ancillis tuis.
PROV|28|1|Fugit impius, nemine persequente;iustus autem quasi leo confidens.
PROV|28|2|Propter peccata terrae multi principes eius;et propter hominem intellegentem et sapientemrectus ordo longior erit.
PROV|28|3|Vir pauper et calumnians pauperessimilis est imbri vehementi, in quo paratur fames.
PROV|28|4|Qui derelinquunt legem, laudant impium;qui custodiunt, succenduntur contra eum.
PROV|28|5|Viri mali non intellegunt iudicium;qui autem requirunt Dominum, animadvertunt omnia.
PROV|28|6|Melior est pauper ambulans in simplicitate suaquam perversus in viis suis, quamquam dives.
PROV|28|7|Qui custodit legem, filius sapiens est;qui autem comissatores pascit, confundit patrem suum.
PROV|28|8|Qui coacervat divitias suas usuris et fenore,liberali in pauperes congregat eas.
PROV|28|9|Qui declinat aures suas, ne audiat legem,oratio quoque eius erit exsecrabilis.
PROV|28|10|Qui decipit iustos in via mala, in interitu suo corruet,et simplices possidebunt bona eius.
PROV|28|11|Sapiens sibi videtur vir dives,pauper autem prudens scrutabitur eum.
PROV|28|12|In exsultatione iustorum multa gloria est,et, cum exaltantur impii, abscondit se homo.
PROV|28|13|Qui abscondit scelera sua, non prosperabit;qui autem confessus fuerit et reliquerit ea,misericordiam consequetur.
PROV|28|14|Beatus homo, qui semper est pavidus;qui vero indurat cor suum, corruet in malum.
PROV|28|15|Leo rugiens et ursus esuriensprinceps impius super populum pauperem.
PROV|28|16|Dux indigens prudentia multos opprimet;qui autem odit avaritiam, longi fient dies eius.
PROV|28|17|Hominem, animae cuiusdam sanguine gravatum,si usque ad lacum fugerit, nemo sustineat.
PROV|28|18|Qui ambulat simpliciter, salvus erit;qui perversis graditur viis, subito concidet.
PROV|28|19|Qui operatur terram suam, satiabitur panibus;qui autem sectatur otium, replebitur egestate.
PROV|28|20|Vir fidelis multum laudabitur;qui autem festinat ditari, non erit innocens.
PROV|28|21|Qui dignoscit in iudicio faciem, non benefacit;et pro buccella panis praevaricatur homo.
PROV|28|22|Festinat ditari vir invidus,ignorat quod egestas superveniet ei.
PROV|28|23|Qui corripit hominem, gratiam postea invenietmagis quam ille, qui lingua blanditur.
PROV|28|24|Qui abripit aliquid a patre suo et a matreet dicit: " Hoc non est peccatum ",particeps homicidae est.
PROV|28|25|Qui desiderium dilatat, iurgia concitat;qui vero sperat in Domino, impinguabitur.
PROV|28|26|Qui confidit in corde suo, stultus est;qui autem graditur sapienter, ipse salvabitur.
PROV|28|27|Qui dat pauperi, non indigebit;qui autem occultat oculos, abundabit maledictis.
PROV|28|28|Cum surrexerint impii, abscondentur homines;cum illi perierint, multiplicabuntur iusti.
PROV|29|1|Vir, qui correptiones dura cervice contemnit,subito conteretur absque sanatione.
PROV|29|2|In multiplicatione iustorum laetabitur vulgus;et in dominatione impii gemet populus.
PROV|29|3|Vir, qui amat sapientiam, laetificat patrem suum;qui autem nutrit scorta, perdet substantiam.
PROV|29|4|Rex in iustitia erigit terram;vir acceptor donorum destruet eam.
PROV|29|5|Homo, qui blanditur amico suo,rete expandit gressibus eius.
PROV|29|6|In peccato vir iniquus irretitur laqueo,et iustus exsultabit atque gaudebit.
PROV|29|7|Novit iustus causam pauperum,impius ignorat scientiam.
PROV|29|8|Homines pestilentes dissipant civitatem;sapientes vero avertunt furorem.
PROV|29|9|Vir sapiens, si cum stulto iudicio contenderit,sive irascatur sive rideat, non inveniet requiem.
PROV|29|10|Viri sanguinum oderunt simplicem;iusti autem quaerunt animam eius.
PROV|29|11|Totum spiritum suum profert stultus;sapiens mitigat eum in posterum.
PROV|29|12|Princeps, qui libenter audit verba mendacii,omnes ministros habet impios.
PROV|29|13|Pauper et oppressor obviaverunt sibi,utriusque oculorum illuminator est Dominus.
PROV|29|14|Rex, qui iudicat in veritate pauperes,thronus eius in aeternum firmabitur.
PROV|29|15|Virga atque correptio tribuit sapientiam;puer autem, qui dimittitur voluntati suae, confundit matrem suam.
PROV|29|16|In multiplicatione impiorum multiplicabuntur scelera,et iusti ruinas eorum videbunt.
PROV|29|17|Erudi filium tuum, et refrigerabit teet dabit delicias animae tuae.
PROV|29|18|Cum visio defecerit, dissipabitur populus;qui vero custodit legem, beatus est.
PROV|29|19|Servus verbis non potest erudiri,quia intellegit et respondere contemnit.
PROV|29|20|Vidisti hominem velocem ad loquendum?Magis illo spem habebit insipiens.
PROV|29|21|Qui delicate a pueritia nutrit servum suum,postea sentiet eum contumacem.
PROV|29|22|Vir iracundus provocat rixas;et, qui ad indignandum facilis est, erit ad peccandum proclivior.
PROV|29|23|Superbia hominis humiliabit eum,et humilis spiritu suscipiet gloriam.
PROV|29|24|Qui cum fure participat, odit animam suam;adiuramentum audit et non indicat.
PROV|29|25|Timor hominis inducit laqueum;qui sperat in Domino, sublevabitur.
PROV|29|26|Multi requirunt faciem principis;et iudicium a Domino egreditur singulorum.
PROV|29|27|Abominantur iusti virum impium;et abominantur impii eos, qui recta sunt via.
PROV|30|1|Verba Agur filii Iaces ex Massa.Oraculum hominis ad Itiel,ad Itiel et Ucal.
PROV|30|2|Quoniam stultissimus sum virorum,et sapientia hominum non est mecum;
PROV|30|3|et non didici sapientiamet scientiam sanctorum non novi.
PROV|30|4|Quis ascendit in caelum atque descendit?Quis continuit spiritum in manibus suis?Quis colligavit aquas quasi in vestimento?Quis statuit omnes terminos terrae?Quod nomen est eius, et quod nomen filii eius, si nosti?
PROV|30|5|Omnis sermo Dei probatusclipeus est sperantibus in eum.
PROV|30|6|Ne addas quidquam verbis illius:et arguaris inveniarisque mendax.
PROV|30|7|Duo rogavi te,ne deneges mihi, antequam moriar:
PROV|30|8|vanitatem et verba mendacia longe fac a me,mendicitatem et divitias ne dederis mihi,tribue tantum victum demensum mihi,
PROV|30|9|ne forte satiatus illiciar ad negandumet dicam: " Quis est Dominus? "aut egestate compulsus fureret periurem nomen Dei mei.
PROV|30|10|Ne calumnieris servum ad dominum suum,ne forte maledicat tibi, et puniaris.
PROV|30|11|Generatio, quae patri suo maledicitet quae matri suae non benedicit.
PROV|30|12|Generatio, quae sibi munda videturet non est lota a sordibus suis.
PROV|30|13|Generatio, cuius oculi quam excelsi sunt,et palpebrae eius in alta surrectae!
PROV|30|14|Generatio, quae pro dentibus gladios habet,et cultri molares eius,ut comedat inopes de terraet pauperes ex hominibus.
PROV|30|15|Sanguisugae duae sunt filiae: Affer, affer! ".Tria sunt insaturabilia,et quattuor, quae numquam dicunt: " Sufficit! ":
PROV|30|16|infernus et venter sterilis,terra, quae non satiatur aqua,ignis, qui numquam dicit: " Sufficit! ".
PROV|30|17|Oculum, qui subsannat patremet qui despicit obsequium matris suae,effodiant eum corvi de torrente,et comedant eum filii aquilae.
PROV|30|18|Tria sunt nimis difficilia mihi,et quattuor penitus ignoro:
PROV|30|19|viam aquilae in caelo,viam colubri super petram,viam navis in medio mariet viam viri in adulescentula.
PROV|30|20|Talis est et via mulieris adulterae,quae comedit et tergens os suum dicit: Non sum operata malum ".
PROV|30|21|Per tria movetur terra,et quattuor non potest sustinere:
PROV|30|22|per servum, cum regnaverit,per stultum, cum saturatus fuerit cibo,
PROV|30|23|per odiosam mulierem, cum in matrimonio fuerit assumpta,et per ancillam, cum fuerit heres dominae suae.
PROV|30|24|Quattuor sunt minima terrae,et ipsa sunt sapientiora sapientibus:
PROV|30|25|formicae populus infirmus,quae praeparant in messe cibum sibi;
PROV|30|26|hyraces plebs invalida,qui collocant in petra cubile suum;
PROV|30|27|regem locusta non habetet egreditur universa per turmas suas;
PROV|30|28|stellio manibus nitituret moratur in aedibus regis.
PROV|30|29|Tria sunt, quae bene gradiuntur,et quattuor, quae incedunt feliciter:
PROV|30|30|leo fortissimus bestiarumad nullius pavebit occursum,
PROV|30|31|gallus succinctus lumbos et arieset rex, qui secum habet exercitum.
PROV|30|32|Si stultum te praebuisti, postquam elevatus es in sublime,et si considerasti, ori impone manum.
PROV|30|33|Qui enim fortiter premit lac, exprimit butyrum,et, qui vehementer emungit nares, elicit sanguinem,et, qui provocat iras, producit discordias.
PROV|31|1|Verba Lamuelis regis Massa, quae erudivit eum mater eius.
PROV|31|2|Quid, fili mi? Quid, fili uteri mei?Quid, fili votorum meorum?
PROV|31|3|Ne dederis mulieribus substantiam tuamet vias tuas illis, quae delent reges.
PROV|31|4|Non decet reges, o Lamuel, non decet reges bibere vinum,nec magistratus desiderare siceram,
PROV|31|5|ne forte bibant et obliviscantur iudiciorumet mutent causam omnium filiorum pauperis.
PROV|31|6|Date siceram pereuntiet vinum his, qui amaro sunt animo:
PROV|31|7|bibat et obliviscatur egestatis suaeet doloris sui non recordetur amplius.
PROV|31|8|Aperi os tuum pro mutoet causis omnium filiorum, qui pereunt;
PROV|31|9|aperi os tuum, decerne, quod iustum est,et iudica inopem et pauperem.
PROV|31|10|ALEPH. Mulierem fortem quis inveniet?Longe super gemmas pretium eius.
PROV|31|11|BETH. Confidit in ea cor viri sui et spoliis non indigebit.
PROV|31|12|GHIMEL. Reddet ei bonum et non malum omnibus diebus vitae suae.
PROV|31|13|DALETH. Quaesivit lanam et linumet operata est delectatione manuum suarum.
PROV|31|14|HE. Facta est quasi navis institorisde longe portans panem suum.
PROV|31|15|VAU. Et de nocte surrexitdeditque praedam domesticis suiset cibaria ancillis suis.
PROV|31|16|ZAIN. Consideravit agrum et emit eum;de fructu manuum suarum plantavit vineam.
PROV|31|17|HETH. Accinxit fortitudine lumbos suoset roboravit brachium suum.
PROV|31|18|TETH. Gustavit et vidit quia bona est negotiatio eius;non exstinguetur in nocte lucerna eius.
PROV|31|19|IOD. Manum suam misit ad colos,et digiti eius apprehenderunt fusum.
PROV|31|20|CAPH. Palmas suas aperuit inopiet manum suam extendit ad pauperem.
PROV|31|21|LAMED. Non timebit domui suae a frigoribus nivis:omnes enim domestici eius vestiti sunt duplicibus.
PROV|31|22|MEM. Stragulatam vestem fecit sibi;byssus et purpura indumentum eius.
PROV|31|23|NUN. Nobilis in portis vir eius,quando sederit cum senatoribus terrae.
PROV|31|24|SAMECH. Sindonem fecit et vendiditet cingulum tradidit Chananaeo.
PROV|31|25|Ain. Fortitudo et decor indumentum eius,et ridebit in die novissimo.
PROV|31|26|PHE. Os suum aperuit sapientiae,et lex clementiae in lingua eius.
PROV|31|27|SADE. Consideravit semitas domus suaeet panem otiosa non comedit.
PROV|31|28|COPH. Surrexerunt filii eius et beatissimam praedicaverunt,vir eius et laudavit eam:
PROV|31|29|RES. " Multae filiae fortiter operatae sunt,tu supergressa es universas ".
PROV|31|30|SIN. Fallax gratia et vana est pulchritudo;mulier timens Dominum ipsa laudabitur.
PROV|31|31|TAU. Date ei de fructu manuum suarum,et laudent eam in portis opera eius.
ECCL|1|1|Verba Ecclesiastes filii David regis Ierusalem."
ECCL|1|2|" Vanitas vanitatum,dixit Ecclesiastes,vanitas vanitatum et omnia vanitas ".
ECCL|1|3|Quid lucri est hominide universo labore suo, quo laborat sub sole?
ECCL|1|4|Generatio praeterit, et generatio advenit,terra autem in aeternum stat.
ECCL|1|5|Oritur sol, et occidit solet ad locum suum anhelat ibique renascitur.
ECCL|1|6|Gyrat per meridiem et flectitur ad aquilonem,lustrans universa in circuitu pergit spirituset in circulos suos revertitur.
ECCL|1|7|Omnia flumina pergunt ad mare, et mare non redundat;ad locum, unde exeunt, flumina illuc revertuntur in cursu suo.
ECCL|1|8|Cunctae res difficiles;non potest eas homo explicare sermone.Non saturatur oculus visu,nec auris auditu impletur.
ECCL|1|9|Quod fuit,ipsum est, quod futurum est.Quod factum est,ipsum est, quod faciendum est:
ECCL|1|10|nihil sub sole novum.Si de quadam re dicitur: " Ecce hoc novum est ",iam enim praecessit in saeculis, quae fuerunt ante nos.
ECCL|1|11|Non est priorum memoria,sed nec eorum quidem, qui postea futuri sunt,erit recordatio apud eos,qui futuri sunt in novissimo.
ECCL|1|12|Ego Ecclesiastes fui rex Israel in Ierusalem
ECCL|1|13|et proposui in animo meo quaerere et investigare sapienter de omnibus, quae fiunt sub sole. Hanc occupationem pessimam dedit Deus filiis hominum, ut occuparentur in ea.
ECCL|1|14|Vidi cuncta, quae fiunt sub sole; et ecce universa vanitas et afflictio spiritus.
ECCL|1|15|Quod est curvum, rectum fieri non potest;et, quod deficiens est, numerari non potest.
ECCL|1|16|Locutus sum ego in corde meo dicens: " Ecce ego magnificavi et apposui sapientiam super omnes, qui fuerunt ante me in Ierusalem; et mens mea contemplata est multam sapientiam et scientiam ".
ECCL|1|17|Dedique cor meum, ut scirem sapientiam et scientiam, insipientiam et stultitiam. Et agnovi quod in his quoque esset afflictio spiritus, eo quod
ECCL|1|18|in multa sapientia multus sit maeror;et, qui addit scientiam, addit et laborem.
ECCL|2|1|Dixi ego in corde meo: " Veni, tentabo te gaudio: fruere bo nis "; et ecce hoc quoque vanitas.
ECCL|2|2|De risu dixi: " Insania "et de gaudio: " Quid prodest? ".
ECCL|2|3|Tractavi in corde meo detinere in vino carnem meam, cum cor meum duceretur in sapientia, et amplecti stultitiam, donec viderem quid esset utile filiis hominum, ut faciant sub sole paucis diebus vitae suae.
ECCL|2|4|Magnificavi opera mea: aedificavi mihi domos et plantavi vineas,
ECCL|2|5|feci hortos et pomaria et consevi ea arboribus cuncti generis fructuum
ECCL|2|6|et exstruxi mihi piscinas aquarum, ut irrigarem silvam lignorum germinantium.
ECCL|2|7|Possedi servos et ancillas et habui multam familiam, habui armenta quoque et magnos ovium greges ultra omnes, qui fuerunt ante me in Ierusalem.
ECCL|2|8|Coacervavi mihi etiam argentum et aurum et substantias regum ac provinciarum, feci mihi cantores et cantatrices et delicias filiorum hominum, scyphos et urceos in ministerio ad vina fundenda
ECCL|2|9|et crevi, supergressus sum omnes, qui ante me fuerunt in Ierusalem; sapientia quoque mea perseveravit mecum.
ECCL|2|10|Et omnia, quae desideraverunt oculi mei, non negavi eis nec prohibui cor meum ab omni voluptate, et oblectatum est ex omnibus laboribus, et hanc ratus sum partem meam ab omnibus aerumnis meis.
ECCL|2|11|Cumque me convertissem ad universa opera, quae fecerant manus meae, et ad labores, in quibus sudaveram, et ecce in omnibus vanitas et afflictio spiritus, et nihil lucri esse sub sole.
ECCL|2|12|Verti me ad contemplandam sapientiam et insipientiam et stultitiam: " Quid faciet, inquam, homo, qui veniet post regem? Id quod antea fecerunt.
ECCL|2|13|Et vidi quod tantum praecederet sapientia stultitiam, quantum lux praecedit tenebras.
ECCL|2|14|" Sapientis oculi in capite eius,stultus in tenebris ambulat ";et didici quod unus utriusqueesset interitus.
ECCL|2|15|Et dixi in corde meo: " Si unus et stulti et meus occasus erit, quid mihi prodest quod maiorem sapientiae dedi operam? ". Locutusque cum mente mea, animadverti quod hoc quoque esset vanitas.
ECCL|2|16|Non enim erit memoria sapientis similiter ut stulti in perpetuum; siquidem futura tempora oblivione cuncta pariter operient: moritur doctus similiter ut indoctus.
ECCL|2|17|Et idcirco taeduit me vitae meae, quia malum mihi est, quod sub sole fit; cuncta enim vanitas et afflictio spiritus.
ECCL|2|18|Rursus detestatus sum omnem laborem meum, quo sub sole laboravi, quem relicturus sum homini, qui erit post me;
ECCL|2|19|et quis scit utrum sapiens an stultus futurus sit? Et dominabitur in laboribus meis, quibus desudavi et sollicitus fui sub sole. Hoc quoque vanitas.
ECCL|2|20|Verti me exasperans cor meum de omni labore, quo laboravi sub sole.
ECCL|2|21|Nam est qui laborat in sapientia et doctrina et sollicitudine, et homini, qui non laboraverit, dabit portionem suam; et hoc ergo vanitas et magnum malum.
ECCL|2|22|Quid enim proderit homini de universo labore suo et afflictione cordis, qua sub sole laboravit?
ECCL|2|23|Cuncti dies eius dolores sunt, et aerumnae occupatio eius, nec per noctem cor eius requiescit; et hoc quoque vanitas est.
ECCL|2|24|Nihil melius est homini quam comedere et bibere et ostendere animae suae bona de laboribus suis. Et hoc vidi de manu Dei esse.
ECCL|2|25|Quis enim comedet et deliciis affluet sine eo?
ECCL|2|26|Quia homini bono in conspectu suo dedit sapientiam et scientiam et laetitiam; peccatori autem dedit afflictionem colligendi et congregandi, ut tradat ei, qui placuit Deo; sed et hoc vanitas est et afflictio spiritus.
ECCL|3|1|Omnia tempus habent,et momentum suum cuique negotio sub caelo:
ECCL|3|2|tempus nascendi et tempus moriendi,tempus plantandi et tempus evellendi quod plantatum est,
ECCL|3|3|tempus occidendi et tempus sanandi,tempus destruendi et tempus aedificandi,
ECCL|3|4|tempus flendi et tempus ridendi,tempus plangendi et tempus saltandi,
ECCL|3|5|tempus spargendi lapides et tempus eos colligendi,tempus amplexandi et tempus longe fieri ab amplexibus,
ECCL|3|6|tempus quaerendi et tempus perdendi,tempus custodiendi et tempus abiciendi,
ECCL|3|7|tempus scindendi et tempus consuendi,tempus tacendi et tempus loquendi,
ECCL|3|8|tempus dilectionis et tempus odii,tempus belli et tempus pacis.
ECCL|3|9|Quid lucri habet, qui operatur, de labore suo?
ECCL|3|10|Vidi occupationem, quam dedit Deus filiis hominum, ut occuparentur in ea.
ECCL|3|11|Cuncta fecit bona in tempore suo; et mundum tradidit cordi eorum, et non inveniet homo opus, quod operatus est Deus ab initio usque ad finem.
ECCL|3|12|Cognovi quod nihil boni esset in eis nisi laetari et facere bene in vita sua.
ECCL|3|13|Omnis enim homo, qui comedit et bibit et videt bonum de labore suo, hoc donum Dei est.
ECCL|3|14|Didici quod omnia opera, quae fecit Deus, perseverent in perpetuum; non possumus eis quidquam addere nec auferre, quae fecit Deus, ut timeatur.
ECCL|3|15|Quod iam fuit, ipsum est; et, quod futurum est, iam fuit; et Deus requirit, quod abiit.
ECCL|3|16|Et adhuc vidi sub sole: in loco iudicii ibi impietas, et in loco iustitiae ibi iniquitas;
ECCL|3|17|et dixi in corde meo: " Iustum et impium iudicabit Deus, quia tempus omni rei et omnibus occasio ".
ECCL|3|18|Dixi in corde meo de filiis hominum, ut probaret eos Deus et ostenderet eos in semetipsis similes esse bestiis.
ECCL|3|19|Quoniam sors filiorum hominis et iumentorum una est atque eadem: sicut moritur homo, sic et illa moriuntur; et idem spiritus omnibus: nihil habet homo iumento amplius, quia omnia vanitas.
ECCL|3|20|Et omnia pergunt ad unum locum:de terra facta sunt omnia,et in terram omnia pariter revertuntur.
ECCL|3|21|Quis novit, si spiritus filiorum hominis ascendat sursum, et si spiritus iumentorum descendat deorsum in terram?
ECCL|3|22|Et deprehendi nihil esse melius quam laetari hominem in opere suo; nam haec est pars illius. Quis enim eum adducet, ut post se futura cognoscat?
ECCL|4|1|Verti me ad alia et vidi calumnias, quae sub sole geruntur, et ecce lacrimae oppressorum, et nemo consolator; et ex parte opprimentium violentia, et nemo consolator.
ECCL|4|2|Et laudavi magis mortuos, qui iam defuncti sunt, quam viventes, qui adhuc vitam agunt,
ECCL|4|3|et feliciorem utroque iudicavi, qui necdum natus est nec vidit opera mala, quae sub sole fiunt.
ECCL|4|4|Rursum contemplatus sum omnes labores et omnem successum operis, et hoc esse zelum in proximum suum. Et in hoc ergo vanitas et afflictio spiritus.
ECCL|4|5|Stultus complicat manus suaset comedit carnes suas.
ECCL|4|6|Melior est pugillus cum requiequam plena utraque manus cum labore et afflictione spiritus.
ECCL|4|7|Iterum repperi et aliam vanitatem sub sole:
ECCL|4|8|unus est et secundum non habet, non filium, non fratrem, et tamen laborare non cessat, nec satiantur oculi eius divitiis, nec recogitat dicens: " Cui laboro et fraudo animam meam bonis?". In hoc quoque vanitas est et occupatio pessima.
ECCL|4|9|Melius est duos esse simul quam unum: habent enim emolumentum in labore suo,
ECCL|4|10|quia si unus ceciderit, ab altero fulcietur. Vae soli! Cum ceciderit, non habet sublevantem se.
ECCL|4|11|Insuper, si dormierint duo, fovebuntur mutuo; unus quomodo calefiet?
ECCL|4|12|Et, si quispiam praevaluerit contra unum, duo resistent ei. Et fu niculus triplex non cito rumpitur.
ECCL|4|13|Melior est puer pauper et sapiensrege sene et stulto,qui iam nescit erudiri.
ECCL|4|14|Ille enim de domo carceris exivit, ut regnaret, etiamsi in regno istius natus sit pauper.
ECCL|4|15|Vidi cunctos viventes, qui ambulant sub sole, cum adulescente illo secundo, qui consurgebat pro eo.
ECCL|4|16|Infinitus numerus erat populi, omnium, quos ipse praecedebat; sed qui postea futuri sunt, non laetabuntur in eo. Et hoc vanitas et afflictio spiritus.
ECCL|4|17|Custodi pedem tuum ingrediens domum Dei, nam accedere, ut audias, melius est quam cum stulti offerunt victimas: multo enim melior est oboedientia quam stultorum victimae, qui nesciunt se malum facere.
ECCL|5|1|Ne temere quid loquaris, neque cor tuum sit velox ad proferen dum sermonem coram Deo; Deus enim in caelo, et tu super terram: idcirco sint pauci sermones tui.
ECCL|5|2|Multas curas sequuntur somnia,et in multis sermonibus invenietur stultitia.
ECCL|5|3|Si quid vovisti Deo, ne moreris reddere: displicet enim ei stulta promissio; sed, quodcumque voveris, redde.
ECCL|5|4|Multoque melius est non vovere, quam post votum promissa non reddere.
ECCL|5|5|Ne dederis os tuum, ut peccare faciat carnem tuam, neque dicas coram angelo: " Error fuit "; ne forte iratus Deus contra sermones tuos dissipet opera manuum tuarum.
ECCL|5|6|Ubi multa sunt somnia, plurimae sunt vanitates et sermones innumeri; tu vero Deum time.
ECCL|5|7|Si videris calumnias egenorum et subreptionem iudicii et iustitiae in provincia, non mireris super hoc negotio, quia excelso excelsior vigilat, et super hos quoque eminentiores sunt alii;
ECCL|5|8|et terrae lucrum in omnibus est rex, cuius agri culti sunt.
ECCL|5|9|Qui diligit pecuniam, pecunia non implebitur; et, qui amat divitias, fructum non capiet ex eis; et hoc ergo vanitas.
ECCL|5|10|Ubi multae sunt opes, multi et qui comedunt eas; et quid prodest possessori, nisi quod cernit divitias oculis suis?
ECCL|5|11|Dulcis est somnus operanti,sive parum sive multum comedat;saturitas autem divitisnon sinit eum dormire.
ECCL|5|12|Est et infirmitas pessima, quam vidi sub sole: divitiae conservatae in malum domini sui.
ECCL|5|13|Perierunt enim in negotio pessimo; si generavit filium, in summa egestate erit.
ECCL|5|14|Sicut egressus est de utero matris suae, nudus iterum abibit, sicut venit, et nihil auferet secum de labore suo, quod tollat in manu sua.
ECCL|5|15|Miserabilis prorsus infirmitas: quomodo venit, sic revertetur. Quid ergo prodest ei quod laboravit in ventum?
ECCL|5|16|Cunctis enim diebus vitae suae comedit in tenebris et in curis multis et in aerumna atque tristitia.
ECCL|5|17|Ecce quod ego vidi bonum, quod pulchrum, ut comedat quis et bibat et fruatur laetitia ex labore suo, quo laboravit ipse sub sole, numero dierum vitae suae, quos dedit ei Deus; haec enim est pars illius.
ECCL|5|18|Et quidem omni homini, cui dedit Deus divitias atque substantiam, potestatemque ei tribuit, ut comedat ex eis et tollat partem suam et laetetur de labore suo: hoc est donum Dei.
ECCL|5|19|Non enim satis recordabitur dierum vitae suae, eo quod Deus occupet deliciis cor eius.
ECCL|6|1|Est et aliud malum, quod vidi sub sole, et quidem grave apud homines:
ECCL|6|2|vir, cui dedit Deus divitias et substantiam et honorem, et nihil deest animae suae ex omnibus, quae desiderat; nec tribuit ei potestatem Deus, ut comedat ex eo, sed homo extraneus vorabit illud: hoc vanitas et miseria mala est.
ECCL|6|3|Si genuerit quispiam centum liberos et vixerit multos annos et plures dies aetatis habuerit, et anima illius non sit satiata bonis substantiae suae, immo et sepultura careat, de hoc ego pronuntio quod melior illo sit abortivus.
ECCL|6|4|Frustra enim venit et pergit ad tenebras, et in tenebris abscondetur nomen eius.
ECCL|6|5|Etsi non vidit solem neque cognovit, maior est requies isti quam illi.
ECCL|6|6|Etiamsi duobus milibus annis vixerit et non fuerit perfruitus bonis, nonne ad unum locum properant omnes?
ECCL|6|7|" Omnis labor hominis est ad os eius,sed anima eius non implebitur ".
ECCL|6|8|Quid habet amplius sapiens prae stulto? Et quid pauper, qui sciat ambulare coram vivis?
ECCL|6|9|" Melior est oculorum visio quam vana persequi desideria "; sed et hoc vanitas est et afflictio spiritus.
ECCL|6|10|Quidquid est, iam vocatum est nomen eius; et scitur quod homo sit et non possit contra fortiorem se in iudicio contendere.
ECCL|6|11|Ubi verba sunt plurima, multiplicant vanitatem; quid lucri habet homo?
ECCL|6|12|Quoniam quis scit quid homini bonum sit in vita, in paucis diebus vanitatis suae, quos peragit velut umbra? Aut quis ei poterit indicare quid post eum futurum sub sole sit?
ECCL|7|1|Melius est nomen bonum quam unguenta pretiosa,et dies mortis die nativitatis.
ECCL|7|2|Melius est ire ad domum luctusquam ad domum convivii;in illa enim finis cunctorum hominum,et vivens hoc conferet in corde.
ECCL|7|3|Melior est tristitia risu,quia per tristitiam vultus corrigitur animus.
ECCL|7|4|Cor sapientium in domo luctus,et cor stultorum in domo laetitiae.
ECCL|7|5|Melius est a sapiente corripiquam laetari stultorum canticis,
ECCL|7|6|quia sicut sonitus spinarum ardentium sub olla,sic risus stulti.Sed et hoc vanitas.
ECCL|7|7|Quia calumnia stultum facit sapientem,et munus cor insanire facit.
ECCL|7|8|" Melior est finis negotii quam principium,melior est patiens arrogante ".
ECCL|7|9|Ne sis velox in animo ad irascendum, quia ira in sinu stulti requiescit.
ECCL|7|10|Ne dicas: "Quid, putas, causae est quod priora tempora meliora fuere quam nunc sunt? ". Non enim ex sapientia interrogas de hoc.
ECCL|7|11|Bona est sapientia cum divitiis et prodest videntibus solem.
ECCL|7|12|Sicut enim protegit sapientia, sic protegit pecunia; hoc autem plus habet eruditio, quod sapientia vitam tribuit possessori suo.
ECCL|7|13|Considera opera Dei: quod nemo possit corrigere, quod ille curvum fecerit.
ECCL|7|14|In die bona fruere bonis et in die mala considera: sicut hanc, sic et illam fecit Deus, ita ut non inveniat homo quidquam de futuro.
ECCL|7|15|Cuncta vidi in diebus vanitatis meae: est iustus, qui perit in iustitia sua, et impius, qui multo vivit tempore in malitia sua.
ECCL|7|16|Noli esse nimis iustusneque sapiens supra modum!Cur te perdere vis?
ECCL|7|17|Ne agas nimis impieet noli esse stultus!Cur mori debeas in tempore non tuo?
ECCL|7|18|Bonum est ut, quod habes, teneas, sed et ab illo ne subtrahas manum tuam, quia qui timet Deum, utrumque devitat.
ECCL|7|19|Sapientia confortabit sapientem super decem principes civitatis.
ECCL|7|20|Nullus enim homo iustus in terra, qui faciat bonum et non peccet.
ECCL|7|21|Sed et cunctis sermonibus, qui dicuntur, ne accommodes cor tuum, ne forte audias servum tuum maledicentem tibi;
ECCL|7|22|scit enim conscientia tua, quia et tu crebro maledixisti aliis.
ECCL|7|23|Cuncta tentavi in sapientia, dixi: " Sapiens efficiar ".
ECCL|7|24|Et ipsa longius recessit a me. Longe est, quod fuit; et alta est profunditas. Quis inveniet eam?
ECCL|7|25|Lustravi universa animo meo, ut scirem et considerarem et quaererem sapientiam et rationem et ut cognoscerem impietatem esse stultitiam et errorem imprudentiam.
ECCL|7|26|Et invenio amariorem morte mulierem, quae laqueus venatorum est, et sagena cor eius, vincula sunt manus illius. Qui placet Deo, effugiet eam; qui autem peccator est, capietur ab illa.
ECCL|7|27|Ecce hoc inveni, dixit Ecclesiastes, unum et alterum, ut invenirem rationem,
ECCL|7|28|quam adhuc quaerit anima mea, et non inveni:Hominem de mille unum repperi,mulierem ex omnibus non inveni.
ECCL|7|29|Ecce solummodo hoc inveni:Quod fecerit Deus hominem rectum,et ipsi quaesierint infinitas quaestiones.
ECCL|8|1|Quis talis, ut sapiens est?Et quis cognovit solutionem re rum?Sapientia hominis illuminat vultum eius,et durities faciei illius commutatur.
ECCL|8|2|Os regis observa et propter iuramenta Dei
ECCL|8|3|ne festines recedere a facie eius neque permaneas in re mala, quia omne, quod voluerit, faciet.
ECCL|8|4|Quia sermo illius potestate plenus est, nec dicere ei quisquam potest: " Quare ita facis? ".
ECCL|8|5|Qui custodit praeceptum, non experietur quidquam mali; tempus et iudicium cor sapientis intellegit.
ECCL|8|6|Omni enim negotio tempus est et iudicium, et multa hominis afflictio;
ECCL|8|7|ignorat enim quid futurum sit, nam quomodo sit futurum, quis nuntiabit ei?
ECCL|8|8|Non est in hominis potestate dominari super spiritum nec cohibere spiritum, nec habet potestatem supra diem mortis, nec ulla remissio est ingruente bello, neque salvabit impietas impium.
ECCL|8|9|Omnia haec consideravi et dedi cor meum cunctis operibus, quae fiunt sub sole, quo tempore dominatur homo homini in malum suum.
ECCL|8|10|Et ita vidi impios sepultos, discedentes de loco sancto; in oblivionem cadere in civitate, quod ita egerunt: sed et hoc vanitas est.
ECCL|8|11|Etenim, quia non profertur cito sententia contra opera mala, ideo cor filiorum hominum repletur, ut perpetrent mala.
ECCL|8|12|Nam peccator centies facit malum et prolongat sibi dies; verumtamen novi quod erit bonum timentibus Deum, qui verentur faciem eius.
ECCL|8|13|Non sit bonum impio, nec prolongabit dies suos quasi umbram, qui non timet faciem Domini.
ECCL|8|14|Est vanitas, quae fit super terram: sunt iusti, quibus mala proveniunt, quasi opera egerint impiorum, et sunt impii, quibus bona proveniunt, quasi iustorum facta habeant; sed et hoc vanissimum iudico.
ECCL|8|15|Laudavi igitur laetitiam quod non esset homini bonum sub sole, nisi quod comederet et biberet atque gauderet et hoc solum secum auferret de labore suo in diebus vitae suae, quos dedit ei Deus sub sole.
ECCL|8|16|Cum apposui cor meum, ut scirem sapientiam et intellegerem occupationem, quae versatur in terra, quod diebus et noctibus somnum non capit oculis,
ECCL|8|17|ecce intellexi quod omnium operum Dei nullam possit homo invenire rationem eorum, quae fiunt sub sole; et quanto plus laboraverit homo ad quaerendum, tanto minus inveniet; etiamsi dixerit sapiens se nosse, non poterit reperire.
ECCL|9|1|Omnia haec contuli in corde meo, ut curiose intellegerem quod iusti atque sapientes et opera eorum sunt in manu Dei. Utrum amor sit an odium, omnino nescit homo: coram illis omnia.
ECCL|9|2|Sicut omnibus sors una:iusto et impio,bono et malo,mundo et immundo,immolanti victimas et non immolanti.Sicut bonus sic et peccator;ut qui iurat, ita et ille qui iuramentum timet.
ECCL|9|3|Hoc est pessimum inter omnia, quae sub sole fiunt, quia sors eadem cunctis; unde et corda filiorum hominum implentur malitia et stultitia in vita sua, et novissima eorum apud mortuos.
ECCL|9|4|Qui enim sociatur omnibus viventibus, habet fiduciam: melior est canis vivus leone mortuo.
ECCL|9|5|Viventes enim sciunt se esse morituros; mortui vero nihil noverunt amplius nec habent ultra mercedem, quia oblivioni tradita est memoria eorum.
ECCL|9|6|Amor quoque eorum et odium et invidiae simul perierunt, nec iam habent partem in hoc saeculo et in opere, quod sub sole geritur.
ECCL|9|7|Vade ergo et comede in laetitia panem tuumet bibe cum gaudio vinum tuum,etenim iam diu placuerunt Deo opera tua.
ECCL|9|8|Omni tempore sint vestimenta tua candida,et oleum de capite tuo non deficiat.
ECCL|9|9|Perfruere vita cum uxore, quam diligis, cunctis diebus vitae instabilitatis tuae, qui dati sunt tibi sub sole omni tempore vanitatis tuae: haec est enim pars in vita et in labore tuo, quo laboras sub sole.
ECCL|9|10|Quodcumque facere potest manus tua, instanter operare, quia nec opus nec ratio nec sapientia nec scientia erunt apud inferos, quo tu properas.
ECCL|9|11|Verti me ad aliud et vidi sub sole nec velocium esse cursum nec fortium bellum nec sapientium panem nec doctorum divitias nec prudentium gratiam, sed tempus casumque in omnibus.
ECCL|9|12|Insuper nescit homo finem suum, sed sicut pisces capiuntur sagena mala, et sicut aves laqueo comprehenduntur, sic capiuntur homines in tempore malo, cum eis extemplo supervenerit.
ECCL|9|13|Hanc quoque sub sole vidi sapientiam et probavi maximam:
ECCL|9|14|civitas parva, et pauci in ea viri; venit contra eam rex magnus et vallavit eam exstruxitque munitiones magnas per gyrum.
ECCL|9|15|Inventusque est in ea vir pauper et sapiens et liberavit urbem per sapientiam suam; et nullus deinceps recordatus est hominis illius pauperis.
ECCL|9|16|Et dicebam ego meliorem esse sapientiam fortitudine,sed sapientia pauperis contemnitur,et verba eius non sunt audita.
ECCL|9|17|Verba sapientium cum lenitate audiunturplus quam clamor principis inter stultos.
ECCL|9|18|Melior est sapientia quam arma bellica;sed unus, qui peccaverit, multa bona perdet.
ECCL|10|1|Muscae morientes perdunt et corrumpunt oleum unguentarii.Gravior quam sapientia et gloria est parva stultitia.
ECCL|10|2|Cor sapientis in dextera eius,et cor stulti in sinistra illius.
ECCL|10|3|Sed et in via stultus ambulans, cum ipse insipiens sit, omnes stultos aestimat.
ECCL|10|4|Si spiritus potestatem habentis ascenderit contra te, locum tuum ne dimiseris, quia lenitas faciet cessare peccata maxima.
ECCL|10|5|Est malum, quod vidi sub sole quasi errorem egredientem a facie principis:
ECCL|10|6|positum stultum in dignitate sublimi et divites sedere deorsum.
ECCL|10|7|Vidi servos in equis et principes ambulantes super terram quasi servos.
ECCL|10|8|Qui fodit foveam, incidet in eam;et, qui dissipat murum, mordebit eum coluber.
ECCL|10|9|Qui excidit lapides, affligetur in eis;et, qui scindit ligna, periclitabitur ex eis.
ECCL|10|10|Si retusum fuerit ferrum, et aciem eius non exacueris, labor multiplicabitur, sed lucrum industriae erit sapientia.
ECCL|10|11|Si mordeat serpens incantatione neglecta, nihil lucri habet incantator.
ECCL|10|12|Verba oris sapientis gratia,et labia insipientis praecipitabunt eum.
ECCL|10|13|Initium verborum eius stultitia,et novissimum oris illius insipientia mala.
ECCL|10|14|Stultus verba multiplicat: Ignorat homo quid futurum sit;et, quid post se futurum sit, quis ei poterit indicare?".
ECCL|10|15|Labor stultorum affliget eos,qui nesciunt in urbem pergere.
ECCL|10|16|Vae tibi, terra, cuius rex puer est,et cuius principes mane comedunt.
ECCL|10|17|Beata terra, cuius rex nobilis est,et cuius principes vescuntur in tempore suoad reficiendum et non ad luxuriam.
ECCL|10|18|In pigris manibus humiliabitur contignatio,et in remissis perstillabit domus.
ECCL|10|19|In risum faciunt epulas;vinum laetificat vitam,et pecunia praestat omnia.
ECCL|10|20|In cogitatione tua regi ne detrahaset in secreto cubiculi tui ne maledixeris diviti,quia et aves caeli portabunt vocem tuam,et, qui habet pennas, annuntiabit sententiam.
ECCL|11|1|Mitte panem tuum super transeuntes aquas, quia post tempora multa invenies illum.
ECCL|11|2|Da partem septem necnon et octo, quia ignoras, quid futurum sit mali super terram.
ECCL|11|3|Si repletae fuerint nubes,imbrem super terram effundent;si ceciderit lignum ad austrum aut ad aquilonem,in quocumque loco ceciderit, ibi erit.
ECCL|11|4|Qui observat ventum, non seminat, et, qui considerat nubes, numquam metet.
ECCL|11|5|Quomodo ignoras, quae sit via spiritus, et qua ratione compingantur ossa in ventre praegnantis, sic nescis opera Dei, qui fabricator est omnium.
ECCL|11|6|Mane semina semen tuum,et vespere ne cesset manus tua,quia nescis quid magis prosit,hoc aut illud,et si utrumque simul melius erit.
ECCL|11|7|Dulce lumen,et delectabile est oculis videre solem.
ECCL|11|8|Si annis multis vixerit homoet in his omnibus laetatus fuerit,meminisse debet tenebrosi temporis, quod multum erit:omne, quod venerit, vanitas.
ECCL|11|9|Laetare ergo, iuvenis, in adulescentia tua,et in bono sit cor tuum in diebus iuventutis tuae,et ambula in viis cordis tuiet in intuitu oculorum tuorumet scito quod pro omnibus hisadducet te Deus in iudicium.
ECCL|11|10|Aufer curam a corde tuoet amove malum a carne tua;adulescentia enim et iuventus vanae sunt.
ECCL|12|1|Memento Creatoris tuiin diebus iuventutis tuae,antequam veniat tempus afflictionis,et appropinquent anni, de quibus dicas: Non mihi placent ";
ECCL|12|2|antequam tenebrescatsol et lumen et luna et stellae,et revertantur nubes post pluviam;
ECCL|12|3|quando commovebuntur custodes domus,et nutabunt viri fortissimi,et otiosae erunt molentes imminuto numero,et tenebrescent videntes per foramina,
ECCL|12|4|et claudentur ostia in plateasubmissa voce molentis,et consurgent ad vocem volucris,et subsident omnes filiae carminis;
ECCL|12|5|excelsa quoque timebuntet formidabunt in via.Florebit amygdalus,reptabit locusta,et dissipabitur capparis,quoniam ibit homo in domum aeternitatis suae,et circuibunt in platea plangentes,
ECCL|12|6|antequam rumpatur funiculus argenteus,et frangatur lecythus aureus,et conteratur hydria super fontem,et confringatur rota super cisternam,
ECCL|12|7|et revertatur pulvis in terram suam, unde erat,et spiritus redeat ad Deum, qui dedit illum.
ECCL|12|8|Vanitas vanitatum,dixit Ecclesiastes,et omnia vanitas.
ECCL|12|9|Cumque esset sapientissimus, Ecclesiastes docuit insuper populum scientiam; ponderavit et investigans composuit parabolas multas.
ECCL|12|10|Quaesivit Ecclesiastes verba delectabilia et conscripsit sermones rectissimos ac veritate plenos.
ECCL|12|11|Verba sapientium sicut stimuli, et quasi clavi defixi sunt magistri collationum; data sunt a pastore uno.
ECCL|12|12|His amplius, fili mi, ne requiras: faciendi plures libros nullus est finis, frequensque meditatio carnis afflictio est.
ECCL|12|13|Finis loquendi, omnibus auditis: Deum time et mandata eius observa; hoc est enim omnis homo.
ECCL|12|14|Et cuncta, quae fiunt, adducet Deus in iudicium circa omne occultum, sive bonum sive malum.
SONG|1|1|Canticum Canticorum Salomonis.
SONG|1|2|Osculetur me osculo oris sui!Nam meliores sunt amores tui vino:
SONG|1|3|in fragrantiam unguentorum tuorum optimorum.Oleum effusum nomen tuum;ideo adulescentulae dilexerunt te.
SONG|1|4|Trahe me post te. Curramus!Introducat me rex in cellaria sua;exsultemus et laetemur in tememores amorum tuorum super vinum;recte diligunt te.
SONG|1|5|Nigra sum sed formosa,filiae Ierusalem,sicut tabernacula Cedar,sicut pelles Salma.
SONG|1|6|Nolite me considerare quod fusca sim,quia decoloravit me sol.Filii matris meae irati sunt mihi;posuerunt me custodem in vineis,vineam meam non custodivi.
SONG|1|7|Indica mihi, tu, quem diligit anima mea,ubi pascas,ubi cubes in meridie,ne vagari incipiampost greges sodalium tuorum.
SONG|1|8|Si ignoras,o pulcherrima inter mulieres,egredere et abi post vestigia gregumet pasce haedos tuosiuxta tabernacula pastorum.
SONG|1|9|Equae in curribus pharaonisassimilavi te, amica mea.
SONG|1|10|Pulchrae sunt genae tuae inter inaures,collum tuum inter monilia.
SONG|1|11|Inaures aureas faciemus tibivermiculatas argento.
SONG|1|12|Dum esset rex in accubitu suo,nardus mea dedit odorem suum.
SONG|1|13|Fasciculus myrrhae dilectus meus mihi,qui inter ubera mea commoratur.
SONG|1|14|Botrus cypri dilectus meus mihiin vineis Engaddi.
SONG|1|15|Ecce tu pulchra es, amica mea,ecce tu pulchra es:oculi tui columbarum.
SONG|1|16|Ecce tu pulcher es, dilecte mi,et decorus.Lectulus noster floridus,
SONG|1|17|tigna domorum nostrarum cedrina,laquearia nostra cupressina.
SONG|2|1|Ego flos campiet lilium convallium.
SONG|2|2|Sicut lilium inter spinas,sic amica mea inter filias.
SONG|2|3|Sicut malus inter ligna silvarum,sic dilectus meus inter filios.Sub umbra illius, quem desideraveram, sedi,et fructus eius dulcis gutturi meo.
SONG|2|4|Introduxit me in cellam vinariam,et vexillum eius super me est caritas.
SONG|2|5|Fulcite me uvarum placentis,stipate me malis,quia amore langueo.
SONG|2|6|Laeva eius sub capite meo,et dextera illius amplexatur me.
SONG|2|7|Adiuro vos, filiae Ierusalem,per capreas cervasque camporum,ne suscitetis neque evigilare faciatis dilectam,quoadusque ipsa velit.
SONG|2|8|Vox dilecti mei!Ecce iste venitsaliens in montibus,transiliens colles.
SONG|2|9|Similis est dilectus meus capreaehinnuloque cervorum.En ipse statpost parietem nostrumrespiciens per fenestras,prospiciens per cancellos.
SONG|2|10|En dilectus meus loquitur mihi: Surge, amica mea,columba mea, formosa mea, et veni.
SONG|2|11|Iam enim hiems transiit,imber abiit et recessit.
SONG|2|12|Flores apparuerunt in terra,tempus putationis advenit;vox turturis audita estin terra nostra,
SONG|2|13|ficus protulit grossos suos,vineae florentes dederunt odorem suum;surge, amica mea,speciosa mea, et veni,
SONG|2|14|columba mea, in foraminibus petrae,in caverna abrupta.Ostende mihi faciem tuam,sonet vox tua in auribus meis;vox enim tua dulcis,et facies tua decora ".
SONG|2|15|Capite nobis vulpes, vulpes parvulas,quae demoliuntur vineas,nam vineae nostrae florescunt.
SONG|2|16|Dilectus meus mihi, et ego illi,qui pascitur inter lilia,
SONG|2|17|antequam aspiret dies,et festinent umbrae.Revertere; similis esto,dilecte mi, capreaehinnuloque cervorum super montes Bether.
SONG|3|1|In lectulo meo per noctesquaesivi, quem diligit anima mea;quaesivi illum et non inveni.
SONG|3|2|" Surgam et circuibo civitatem;per vicos et plateasquaeram, quem diligit anima mea".Quaesivi illum et non inveni.
SONG|3|3|Invenerunt me vigiles,qui circumeunt civitatem: Num, quem diligit anima mea, vidistis? ".
SONG|3|4|Paululum cum pertransissem eos,inveni, quem diligit anima mea;tenui eum nec dimittam,donec introducam illum in domum matris meaeet in cubiculum genetricis meae.
SONG|3|5|Adiuro vos, filiae Ierusalem,per capreas cervasque camporum,ne suscitetis neque evigilare faciatis dilectam,donec ipsa velit.
SONG|3|6|Quid hoc, quod ascendit per desertumsicut virgula fumi,aromatizans tus et myrrhamet universum pulverem pigmentarii?
SONG|3|7|En lectulum Salomonis.Sexaginta fortes ambiunt illumex fortissimis Israel,
SONG|3|8|omnes tenentes gladioset ad bella doctissimi,uniuscuiusque ensis super femur suumpropter timores nocturnos.
SONG|3|9|Ferculum fecit sibi rex Salomonde lignis Libani;
SONG|3|10|columnas eius fecit argenteas,reclinatorium aureum,sedile purpureum:medium eius stratum ebeneum.Filiae Ierusalem,
SONG|3|11|egredimini et videte,filiae Sion,regem Salomonemin diademate, quo coronavit illum mater suain die desponsationis illiuset in die laetitiae cordis eius.
SONG|4|1|Quam pulchra es, amica mea,quam pulchra es:oculi tui columbarumper velamen tuum.Capilli tui sicut grex caprarum,quae descenderunt de monte Galaad;
SONG|4|2|dentes tui sicut grex tonsarum,quae ascenderunt de lavacro:omnes gemellis fetibus,et sterilis non est inter eas.
SONG|4|3|Sicut vitta coccinea labia tua,et eloquium tuum dulce;sicut fragmen mali punici, ita genae tuaeper velamen tuum.
SONG|4|4|Sicut turris David collum tuum,quae aedificata est cum propugnaculis:mille clipei pendent ex ea,omnis armatura fortium.
SONG|4|5|Duo ubera tua sicut duo hinnuli,capreae gemelli,qui pascuntur in liliis.
SONG|4|6|Antequam aspiret dies,et festinent umbrae,vadam ad montem myrrhaeet ad collem turis.
SONG|4|7|Tota pulchra es, amica mea,et macula non est in te.
SONG|4|8|Veni de Libano, sponsa,veni de Libano,ingredere;respice de capite Amana,de vertice Sanir et Hermon,de cubilibus leonum,de montibus pardorum.
SONG|4|9|Vulnerasti cor meum, soror mea, sponsa,vulnerasti cor meum in uno oculorum tuorumet in uno monili torquis tui.
SONG|4|10|Quam pulchri sunt amores tui, soror, mea sponsa;meliores sunt amores tui vino,et odor unguentorum tuorum super omnia aromata.
SONG|4|11|Favus distillans labia tua, sponsa;mel et lac sub lingua tua,et odor vestimentorum tuorumsicut odor Libani.
SONG|4|12|Hortus conclusus, soror mea, sponsa,hortus conclusus, fons signatus;
SONG|4|13|propagines tuae paradisus malorum punicorumcum optimis fructibus,cypri cum nardo.
SONG|4|14|Nardus et crocus,fistula et cinnamomumcum universis lignis turiferis,myrrha et aloecum omnibus primis unguentis.
SONG|4|15|Fons hortorum,puteus aquarum viventium,quae fluunt impetu de Libano.
SONG|4|16|Surge, aquilo,et veni, auster;perfla hortum meum,et fluant aromata illius.
SONG|5|1|Veniat dilectus meus in hortum suumet comedat fructus eius optimos.Veni in hortum meum, soror mea, sponsa;messui myrrham meam cum aromatibus meis,comedi favum cum melle,bibi vinum cum lacte meo.Comedite, amici, et bibiteet inebriamini, carissimi.
SONG|5|2|Ego dormio, et cor meum vigilat.Vox dilecti mei pulsantis: Aperi mihi, soror mea, amica mea,columba mea, immaculata mea,quia caput meum plenum est rore, et cincinni mei guttis noctium ".
SONG|5|3|" Exspoliavi me tunica mea,quomodo induar illa?Lavi pedes meos,quomodo inquinabo illos?".
SONG|5|4|Dilectus meus misit manum suam per foramen,et venter meus ilico intremuit.
SONG|5|5|Surrexi, ut aperirem dilecto meo;manus meae stillaverunt myrrham,et digiti mei pleni myrrha probatissimasuper ansam pessuli.
SONG|5|6|Aperui dilecto meo;at ille declinaverat atque transierat.Anima mea liquefacta est, quia discesserat.Quaesivi et non inveni illum;vocavi, et non respondit mihi.
SONG|5|7|Invenerunt me custodes,qui circumeunt civitatem;percusserunt me et vulneraverunt me,tulerunt pallium meum mihicustodes murorum.
SONG|5|8|Adiuro vos, filiae Ierusalem:si inveneritis dilectum meum,quid nuntietis ei? Quia amore langueo ".
SONG|5|9|Quid est dilecto tuo prae ceteris,o pulcherrima mulierum?Quid est dilecto tuo prae ceteris,quia sic adiurasti nos?
SONG|5|10|Dilectus meus candidus et rubicundusdignoscitur ex milibus.
SONG|5|11|Caput eius aurum optimum,cincinni eius sicut racemi palmarum,nigri quasi corvus.
SONG|5|12|Oculi eius sicut columbaesuper rivulos aquarum,quae lacte sunt lotaeet resident iuxta fluenta plenissima.
SONG|5|13|Genae illius sicut areolae aromatum,turriculae unguentorum;labia eius liliadistillantia myrrham primam.
SONG|5|14|Manus illius tornatiles aureae,plenae hyacinthis;venter eius opus eburneumdistinctum sapphiris.
SONG|5|15|Crura illius columnae marmoreae,quae fundatae sunt super bases aureas;species eius ut Libani,electus ut cedri.
SONG|5|16|Guttur illius suavissimum,et totus desiderabilis.Talis est dilectus meus, et ipse est amicus meus,filiae Ierusalem.
SONG|6|1|Quo abiit dilectus tuus,o pulcherrima mulierum?Quo declinavit dilectus tuus,et quaeremus eum tecum?
SONG|6|2|Dilectus meus descendit in hortum suumad areolam aromatum,ut pascatur in hortiset lilia colligat.
SONG|6|3|Ego dilecto meo, et dilectus meus mihi,qui pascitur inter lilia.
SONG|6|4|Pulchra es, amica mea, sicut Thersa,decora sicut Ierusalem,terribilis ut castrorum acies ordinata.
SONG|6|5|Averte oculos tuos a me,quia ipsi me conturbant.Capilli tui sicut grex caprarum,quae descenderunt de Galaad.
SONG|6|6|Dentes tui sicut grex ovium,quae ascenderunt de lavacro:omnes gemellis fetibus,et sterilis non est in eis.
SONG|6|7|Sicut fragmen mali punici, sic genae tuaeper velamen tuum.
SONG|6|8|Sexaginta sunt reginae,et octoginta concubinae,et adulescentularum non est numerus;
SONG|6|9|una est columba mea, perfecta mea,una est matri suae,electa genetrici suae.Viderunt eam filiae et beatissimam praedicaverunt;reginae et concubinae, et laudaverunt eam:
SONG|6|10|" Quae est ista, quae progreditur quasi aurora consurgens,pulchra ut luna,electa ut sol,terribilis ut castrorum acies ordinata? ".
SONG|6|11|Descendi in hortum nucum,ut viderem poma convalliumet inspicerem, si floruisset vinea,et germinassent mala punica.
SONG|6|12|Non advertit animus meus,cum posuit me in quadrigas principis populi mei.
SONG|7|1|Convertere, convertere, Sula mitis;convertere, convertere, ut intueamur te.Quid aspicitis in Sulamitem,cum saltat inter binos choros?
SONG|7|2|Quam pulchri sunt pedes tui in calceamentis,filia principis!Flexurae femorum tuorum sicut monilia,quae fabricata sunt manu artificis.
SONG|7|3|Gremium tuum crater tornatilis:numquam indigeat vino mixto;venter tuus sicut acervus triticivallatus liliis.
SONG|7|4|Duo ubera tua sicut duo hinnuli,gemelli capreae,
SONG|7|5|collum tuum sicut turris eburnea.Oculi tui sicut piscinae in Hesebon,quae sunt ad portam Bathrabbim;nasus tuus sicut turris Libani,quae respicit contra Damascum.
SONG|7|6|Caput tuum ut Carmelus,et comae capitis tui sicut purpura;rex vincitur cincinnis.
SONG|7|7|Quam pulchra es et quam decora,carissima, in deliciis!
SONG|7|8|Statura tua assimilata est palmae,et ubera tua botris.
SONG|7|9|Dixi: " Ascendam in palmamet apprehendam fructus eius ".Et erunt ubera tua sicut botri vineae,et odor oris tui sicut malorum.
SONG|7|10|Guttur tuum sicut vinum optimum,dignum dilecto meo ad potandum,labiisque et dentibus illius ad ruminandum.
SONG|7|11|Ego dilecto meo,et ad me appetitus eius.
SONG|7|12|Veni, dilecte mi, egrediamur in agrum,commoremur in villis;
SONG|7|13|mane properabimus ad vineas,videbimus; si floruit vinea,si flores aperiuntur,si floruerunt mala punica;ibi dabo tibi amores meos.
SONG|7|14|Mandragorae dederunt odorem;in portis nostris omnia poma optima,nova et vetera,dilecte mi, servavi tibi.
SONG|8|1|Quis mihi det te fratrem meum,sugentem ubera matris meae,ut inveniam te foris et deosculer te,et iam me nemo despiciat?
SONG|8|2|Apprehenderem te et ducerem in domum matris meae;ibi me doceres,et darem tibi poculum ex vino conditoet mustum malorum granatorum meorum.
SONG|8|3|Laeva eius sub capite meo,et dextera illius amplexatur me.
SONG|8|4|Adiuro vos, filiae Ierusalem,ne suscitetis neque evigilare faciatis dilectam,donec ipsa velit.
SONG|8|5|Quae est ista, quae ascendit de desertoinnixa super dilectum suum?Sub arbore malo suscitavi te;ibi parturivit te mater tua,ibi parturivit te genetrix tua.
SONG|8|6|Pone me ut signaculum super cor tuum,ut signaculum super brachium tuum,quia fortis est ut mors dilectio,dura sicut infernus aemulatio;lampades eius lampades ignisatque flammae divinae.
SONG|8|7|Aquae multae non potuerunt exstinguere caritatem,nec flumina obruent illam;si dederit homo omnem substantiam domus suae pro dilectione,quasi nihil despicient eum.
SONG|8|8|Soror nostra parvaet ubera non habet;quid faciemus sorori nostraein die, quando alloquenda est?
SONG|8|9|Si murus est,aedificemus super eum propugnacula argentea;si ostium est,compingamus illud tabulis cedrinis.
SONG|8|10|Ego murus,et ubera mea sicut turris;ex quo facta sum coram eoquasi pacem reperiens.
SONG|8|11|Vinea fuit Salomoniin Baalhamon.Tradidit eam custodibus;vir affert pro fructu eiusmille argenteos.
SONG|8|12|Vinea mea coram me est;mille tibi, Salomon,et ducenti his, qui custodiunt fructus eius.
SONG|8|13|Quae habitas in hortis,amici auscultant,fac me audire vocem tuam.
SONG|8|14|Fuge, dilecte mi,et assimilare capreaehinnuloque cervorumsuper montes aromatum.
ISA|1|1|Visio Isaiae filii Amos, quam vidit super Iudam et Ierusalem in diebus Oziae, Ioatham, Achaz, Ezechiae regum Iudae.
ISA|1|2|Audite, caeli, et auribus percipe, terra,quoniam Dominus locutus est: Filios enutrivi et exaltavi,ipsi autem spreverunt me.
ISA|1|3|Cognovit bos possessorem suum,et asinus praesepe domini sui;Israel non cognovit,populus meus non intellexit ".
ISA|1|4|Vae genti peccatrici,populo gravi iniquitate,semini nequam, filiis sceleratis!Dereliquerunt Dominum,blasphemaverunt Sanctum Israel,abalienati sunt retrorsum.
ISA|1|5|Super quo percutiemini vos ultra,addentes praevaricationem?Omne caput languidum,et omne cor maerens.
ISA|1|6|A planta pedis usque ad verticemnon est in eo sanitas;vulnus et livor et plaga tumensnon est circumligatanec curata medicamine neque fota oleo.
ISA|1|7|Terra vestra deserta,civitates vestrae succensae igni;regionem vestram coram vobis alieni devorant,et desolabitur sicut in vastitate hostili.
ISA|1|8|Et derelinquetur filia Sionut umbraculum in vinea,sicut tugurium in cucumerario,sicut civitas, quae obsessa est.
ISA|1|9|Nisi Dominus exercituum reliquisset nobis semen,quasi Sodoma fuissemuset quasi Gomorra similes essemus.
ISA|1|10|Audite verbum Domini,principes Sodomorum;percipite auribus legem Dei nostri, populus Gomorrae.
ISA|1|11|" Quo mihi multitudinem victimarum vestrarum?,dicit Dominus.Plenus sum holocaustis arietumet adipe pinguium;et sanguinem vitulorumet agnorum et hircorum nolui.
ISA|1|12|Cum veneritis ante conspectum meum,quis quaesivit haec de manibus vestris,ut ambularetis in atriis meis?
ISA|1|13|Ne afferatis ultra sacrificium vanum;abominatio mihi incensum,neomenia et sabbatum et conventus;non feram scelus cum coetu sollemni;
ISA|1|14|calendas vestras et sollemnitates vestras odivit anima mea,facta sunt mihi molesta, laboravi sustinens.
ISA|1|15|Et cum extenderitis manus vestras,avertam oculos meos a vobis;et cum multiplicaveritis orationem,non exaudiam:manus enim vestrae sanguine plenae sunt.
ISA|1|16|Lavamini, mundi estote,auferte malum cogitationum vestrarum ab oculis meis;quiescite agere perverse,
ISA|1|17|discite benefacere:quaerite iudicium, subvenite oppresso,iudicate pupillo, defendite viduam.
ISA|1|18|Et venite, et iudicio contendamus,dicit Dominus.Si fuerint peccata vestra ut coccinum,quasi nix dealbabuntur;et, si fuerint rubra quasi vermiculus,velut lana erunt.
ISA|1|19|Si volueritis et audieritis,bona terrae comedetis;
ISA|1|20|quod si nolueritis et me ad iracundiam provocaveritis,gladius devorabit vos,quia os Domini locutum est ".
ISA|1|21|Quomodo facta est meretrixcivitas fidelis, plena iudicii?Iustitia habitavit in ea,nunc autem homicidae.
ISA|1|22|Argentum tuum versum est in scoriam,vinum tuum mixtum est aqua;
ISA|1|23|principes tui infideles, socii furum:omnes diligunt munera, sequuntur retributiones,pupillo non iudicant, et causa viduae non ingreditur ad illos.
ISA|1|24|Propter hoc ait Dominus, Deus exercituum, Fortis Israel: Heu, consolabor super hostibus meiset vindicabor de inimicis meis.
ISA|1|25|Et convertam manum meam ad teet excoquam ad purum scoriam tuamet auferam omne stannum tuum.
ISA|1|26|Et restituam iudices tuos, ut fuerunt prius,et consiliarios tuos sicut antiquitus;post haec vocaberis Civitas iustitiae, Urbs fidelis ".
ISA|1|27|Sion in iudicio redimeturet, qui in ea reversi sunt, in iustitia.
ISA|1|28|Erit autem ruina scelestis et peccatoribus simul;et, qui dereliquerunt Dominum, consumentur.
ISA|1|29|Confundemini enim terebinthis, in quibus delectati estis,et erubescetis super hortis, quos elegistis.
ISA|1|30|Nam eritis velut quercus, defluentibus foliis,et velut hortus absque aqua;
ISA|1|31|et erit fortitudo vestra ut favilla stuppae,et opus eius quasi scintilla,et succendetur utrumque simul, et non erit qui exstinguat.
ISA|2|1|Verbum, quod vidit Isaias filius Amos super Iudam et Ieru salem.
ISA|2|2|Et erit in novissimis diebuspraeparatus mons domus Domini in vertice montium,et elevabitur super colles;et fluent ad eum omnes gentes.
ISA|2|3|Et ibunt populi multi et dicent: Venite, et ascendamus ad montem Domini,ad domum Dei Iacob,ut doceat nos vias suas,et ambulemus in semitis eius ";quia de Sion exibit lex,et verbum Domini de Ierusalem.
ISA|2|4|Et iudicabit genteset arguet populos multos;et conflabunt gladios suos in vomereset lanceas suas in falces;non levabit gens contra gentem gladium,nec exercebuntur ultra ad proelium.
ISA|2|5|Domus Iacob, venite,et ambulemus in lumine Domini.
ISA|2|6|Proiecisti enim populum tuum, domum Iacob,quia repleti sunt hariolis orientalibuset augures habuerunt ut Philisthimet manus alienis porrigunt.
ISA|2|7|Repleta est terra eius argento et auro,et non est finis thesaurorum eius;
ISA|2|8|et repleta est terra eius equis,et innumerabiles quadrigae eius;et repleta est terra eius idolis:opus manuum suarum adoraverunt,quod fecerunt digiti eorum.
ISA|2|9|Et incurvavit se homo,et humiliatus est vir:ne dimittas eis.
ISA|2|10|Ingredere in petram, abscondere in pulverea facie timoris Domini et a gloria maiestatis eius.
ISA|2|11|Oculi sublimes hominis humiliabuntur,et incurvabitur altitudo virorum;exaltabitur autem Dominus solus in die illa.
ISA|2|12|Quia dies Domini exercituumsuper omnem superbum et excelsumet super omnem arrogantem, et humiliabitur;
ISA|2|13|et super omnes cedros Libani sublimes et erectaset super omnes quercus Basan
ISA|2|14|et super omnes montes excelsoset super omnes colles elevatos
ISA|2|15|et super omnem turrim excelsamet super omnem murum munitum
ISA|2|16|et super omnes naves Tharsiset super omnia navigia pulchra.
ISA|2|17|Et incurvabitur sublimitas hominum,et humiliabitur altitudo virorum;et elevabitur Dominus solus in die illa,
ISA|2|18|et idola penitus conterentur.
ISA|2|19|Et introibunt in speluncas petrarumet in voragines terraea facie formidinis Domini et a gloria maiestatis eius,cum surrexerit percutere terram.
ISA|2|20|In die illa proiciet homo idola sua argentea et simulacra sua aurea, quae fecerat sibi, ut adoraret, ad talpas et vespertiliones.
ISA|2|21|Et ingredietur scissuras petrarum et cavernas saxorum a facie formidinis Domini et a gloria maiestatis eius, cum surrexerit percutere terram.
ISA|2|22|Quiescite ergo ab homine, cuius spiritus in naribus eius. Quanti enim aestimabitur ipse?
ISA|3|1|Ecce enim Dominator, Dominus exercituum,aufert a Ierusalem et a Iuda robur et praesidium,omne robur panis et omne robur aquae,
ISA|3|2|fortem et virum bellatorem,iudicem et prophetam et hariolum et senem,
ISA|3|3|principem super quinquaginta et honorabilem vultuet consiliarium et sapientem magumet prudentem incantatorem.
ISA|3|4|Et dabo pueros principes eorum;et infantes dominabuntur eis.
ISA|3|5|Et irruet populus, vir ad virum,unusquisque ad proximum suum:tumultuabitur puer contra senem,et ignobilis contra nobilem.
ISA|3|6|Apprehendet enim vir fratrem suumin domo patris sui: Vestimentum tibi est,princeps esto noster,ruina autem haec sub manu tua ".
ISA|3|7|Clamabit in die illa dicens: Non sum medicus,et in domo mea non est panis neque vestimentum;nolite constituere me principem populi ".
ISA|3|8|Ruit enim Ierusalem, et Iudas concidit,quia lingua eorum et adinventiones eorum contra Dominum,ut provocarent oculos maiestatis eius.
ISA|3|9|Procacitas vultus eorum accusat eos,et peccatum suum quasi Sodomapraedicaverunt nec absconderunt;vae animae eorum,quoniam reddita sunt eis mala!
ISA|3|10|Dicite iusto: " Bene! ",quoniam fructum adinventionum suarum comedet.
ISA|3|11|Vae impio in malum:retributio enim manuum eius fiet ei!
ISA|3|12|Populum meum opprimit infans,et mulieres dominantur ei.Popule meus, qui te beatum dicunt, ipsi te decipiuntet viam gressuum tuorum dissipant.
ISA|3|13|Surgit ad arguendum Dominuset stat ad iudicandos populos.
ISA|3|14|Dominus ad iudicium venietcum senibus populi sui et principibus eius: Vos enim depasti estis vineam,et rapina pauperis in domibus vestris.
ISA|3|15|Quare atteritis populum meumet facies pauperum commolitis? ",dicit Dominus, Deus exercituum.
ISA|3|16|Et dixit Dominus: Pro eo quod elevatae sunt filiae Sionet ambulaverunt extento collo et nutibus oculorum,parvis passibus incedebantet catenulis pedum tinniebant,
ISA|3|17|decalvabit Dominus verticem filiarum Sionet Dominus crinem earum nudabit ".
ISA|3|18|In die illa auferet Dominusornamentum calceamentorum et torques
ISA|3|19|et lunulas et inaureset armillas et mitras,
ISA|3|20|discriminalia et periscelidaset fascias et olfactoriola
ISA|3|21|et anulos et ornamenta narium,
ISA|3|22|mutatoria et palliolaet linteamina et marsupia,
ISA|3|23|specula et sindoneset vittas et pallia.
ISA|3|24|Et erit pro suavi odore foetor,et pro zona funiculus,et pro crispante crine calvitium,et pro fascia pectorali cilicium,stigma pro pulchritudine.
ISA|3|25|Viri tui gladio cadent,et fortes tui in proelio,
ISA|3|26|et maerebunt atque lugebunt portae eius,et desolata in terra sedebit.
ISA|4|1|Et apprehendent septem mulieresvirum unum in die illa dicentes: Panem nostrum comedemuset vestimentis nostris operiemur,tantummodo vocetur nomen tuum super nos:aufer opprobrium nostrum ".
ISA|4|2|In die illa erit germen Domini in splendorem et gloriam,et fructus terrae sublimis et exsultatiohis, qui salvati fuerint de Israel.
ISA|4|3|Et erit: omnis, qui relictus fuerit in Sion,et residuus in Ierusalem, sanctus vocabitur,omnis, qui scriptus est ad vitam in Ierusalem.
ISA|4|4|Cum abluerit Dominus sordem filiarum Sionet sanguinem Ierusalem laverit de medio eiusspiritu iudicii et spiritu ardoris,
ISA|4|5|et creabit Dominus super omnem locum montis Sionet super coetum eiusnubem per diemet fumum et splendorem ignis flammantis in nocte:super omnem enim gloriam protectio,
ISA|4|6|et tabernaculum erit in umbraculum diei ab aestuet in securitatem et absconsionem a turbine et a pluvia.
ISA|5|1|Cantabo dilecto meocanticum amici mei de vinea sua:Vinea facta est dilecto meoin colle pingui;
ISA|5|2|et saepivit eamet lapides elegit ex illaet plantavit in ea vites electaset aedificavit turrim in medio eiuset torcular exstruxit in ea;et exspectavit, ut faceret uvas,et fecit labruscas.
ISA|5|3|Nunc ergo, habitator Ierusalemet vir Iudae,iudicate inter me et vineam meam.
ISA|5|4|Quid est quod debui ultra facere vineae meaeet non feci ei?Cur exspectavi, ut faceret uvas,et fecit labruscas?
ISA|5|5|Et nunc ostendam vobisquid ego faciam vineae meae:auferam saepem eius,et erit in direptionem;diruam maceriam eius,et erit in conculcationem.
ISA|5|6|Et ponam eam desertam:non putabitur et non fodietur,et ascendent vepres et spinae;et nubibus mandabo, ne pluant super eam imbrem.
ISA|5|7|Vinea enim Domini exercituum domus Israel est,et vir Iudae germen eius delectabile;et exspectavi, ut faceret iudicium, et ecce iniquitas,et iustitiam, et ecce nequitia.
ISA|5|8|Vae, qui coniungunt domum ad domumet agrum agro copulant usque ad terminum loci!Numquid habitabitis vos soli in medio terrae?
ISA|5|9|In auribus meis iuravit Dominus exercituum: Certe domus multae desertae erunt,grandes et pulchrae absque habitatore ".
ISA|5|10|Decem enim iugera vinearum facient lagunculam unam,et triginta modii sementis facient modios tres.
ISA|5|11|Vae, qui consurgunt mane ad ebrietatem sectandamet ad potandum usque ad vesperam,ut vinum inflammet eos!
ISA|5|12|Cithara et lyraet tympanum et tibiaet vinum in conviviis eorum,et opus Domini non respiciunt,nec opera manuum eius considerant.
ISA|5|13|Propterea captivus ductus est populus meus,quia non habuit scientiam,et nobiles eius interierunt fame,et multitudo eius siti exaruit.
ISA|5|14|Propterea dilatavit infernus fauces suaset aperuit os suum absque ullo termino;et descendunt fortes Ierusalem, et populus eius,et sublimes et tripudiantes in ea.
ISA|5|15|Et incurvabitur homo, et humiliabitur vir,et oculi sublimium deprimentur;
ISA|5|16|et exaltabitur Dominus exercituum in iudicio,et Deus sanctus sanctificabitur in iustitia,
ISA|5|17|et pascentur agni iuxta ordinem suum velut in prato suo,et alieni comedent in ruinis pinguium.
ISA|5|18|Vae, qui trahunt iniquitatem in funiculis vanitatiset quasi vinculum plaustri peccatum!
ISA|5|19|Qui dicunt: " Festinetet cito veniat opus eius, ut videamus;et appropiet et veniat consilium Sancti Israel,et sciemus illud! ".
ISA|5|20|Vae, qui dicunt malum bonum et bonum malum,ponentes tenebras in lucem et lucem in tenebras,ponentes amarum in dulce et dulce in amarum!
ISA|5|21|Vae, qui sapientes sunt in oculis suiset coram ipsis prudentes!
ISA|5|22|Vae, qui potentes sunt ad bibendum vinum,et viri fortes ad miscendam ebrietatem!
ISA|5|23|Qui absolvunt impium pro muneribuset iustitiam iusti auferunt ab eo!
ISA|5|24|Propter hoc, sicut devorat stipulam lingua ignis,et palea flamma consumitur,sic radix eorum quasi tabes erit,et flos eorum sicut putredo ascendet;abiecerunt enim legem Domini exercituumet eloquium Sancti Israel blasphemaverunt.
ISA|5|25|Ideo exarsit furor Domini in populum suum,et extendit manum suam super eum et percussit eum,et conturbati sunt montes;et facta sunt morticina eorum quasi stercus in medio platearum.In his omnibus non est aversus furor eius,sed adhuc manus eius extenta.
ISA|5|26|Et levabit signum nationibus procul;et sibilabit ad eum de finibus terrae;et ecce festinus velociter veniet.
ISA|5|27|Non est deficiens neque laborans in eo,non dormitabit neque dormiet;neque solvetur cingulum renum eius,nec rumpetur corrigia calceamenti eius.
ISA|5|28|Sagittae eius acutae, et omnes arcus eius extenti;ungulae equorum eius ut silex reputantur,et rotae eius quasi impetus tempestatis.
ISA|5|29|Rugitus eius ut leonis:rugiet ut catuli leonum et frendet;et arripiet praedam et in tuto collocabit,et non erit qui eruat.
ISA|5|30|Et sonabit super eum in die illa sicut sonitus maris.Aspiciet in terram: et ecce tenebrae tribulationis,et lux obtenebrata est in caligine eius.
ISA|6|1|In anno, quo mortuus est rex Ozias, vidi Dominum edentem super solium excelsum et elevatum; et fimbriae eius replebant templum.
ISA|6|2|Seraphim stabant iuxta eum; sex alae uni et sex alae alteri: duabus velabat faciem suam et duabus velabat pedes suos et duabus volabat.
ISA|6|3|Et clamabat alter ad alterum et dicebat: Sanctus, Sanctus, Sanctus Dominus exercituum;plena est omnis terra gloria eius ".
ISA|6|4|Et commota sunt superliminaria cardinum a voce clamantis, et domus repleta est fumo.
ISA|6|5|Et dixi: Vae mihi, quia perii!Quia vir pollutus labiis ego sumet in medio populi polluta labia habentis ego habitoet regem, Dominum exercituum, vidi oculis meis ".
ISA|6|6|Et volavit ad me unus de seraphim, et in manu eius calculus, quem forcipe tulerat de altari,
ISA|6|7|et tetigit os meum et dixit: Ecce tetigit hoc labia tua,et auferetur iniquitas tua,et peccatum tuum mundabitur ".
ISA|6|8|Et audivi vocem Domini dicentis: " Quem mittam? Et quis ibit nobis? ". Et dixi: " Ecce ego, mitte me ".
ISA|6|9|Et dixit: " Vade, et dices populo huic:Audientes audite et nolite intellegere,et videntes videte et nolite cognoscere".
ISA|6|10|Pingue redde cor populi huiuset aures eius aggravaet oculos eius excaeca,ne forte videat oculis suiset auribus suis audiatet corde suo intellegat et convertaturet sanetur ".
ISA|6|11|Et dixi: " Usquequo, Domine? ". Et dixit: Donec desolenturcivitates absque habitatore,et domus sine homine,et terra relinquatur deserta ".
ISA|6|12|Et longe adducet Dominus homines,et magna erit desolatio in medio terrae;
ISA|6|13|et adhuc in ea decimatio,et rursus excisioni tradetursicut terebinthus et sicut quercus,in quibus deiectis manebit aliquid stabile.Semen sanctum erit id quod steterit in ea.
ISA|7|1|Et factum est in diebus Achaz filii Ioatham filii Oziae regis Iu dae, ascendit Rasin rex Syriae et Phacee filius Romeliae rex Israel in Ierusalem ad proeliandum contra eam; et non potuerunt debellare eam.
ISA|7|2|Et nuntiaverunt domui David dicentes: " Requievit Syria super Ephraim ". Et commotum est cor eius et cor populi eius, sicut moventur ligna silvarum a facie venti.
ISA|7|3|Et dixit Dominus ad Isaiam: " Egredere in occursum Achaz, tu et Seariasub (id est Reliquiae revertentur) filius tuus, ad extremum aquaeductus piscinae superioris in viam agri fullonis;
ISA|7|4|et dices ad eum: Vide, ut sileas; noli timere, et cor tuum ne formidet a duabus caudis titionum fumigantium istorum, ob ardorem irae Rasin et Syriae et filii Romeliae,
ISA|7|5|eo quod consilium malum inierit contra te Syria, Ephraim et filius Romeliae dicentes:
ISA|7|6|"Ascendamus ad Iudam et terrorem iniciamus ei et avellamus eum ad nos et ponamus regem in medio eius filium Tabeel" ".
ISA|7|7|Haec dicit Dominus Deus: Non stabit et non erit!
ISA|7|8|Caput enim Syriae Damascus,et caput Damasci Rasin;et adhuc sexaginta et quinque anniet desinet Ephraim esse populus;
ISA|7|9|et caput Ephraim Samaria,et caput Samariae filius Romeliae.Si non credideritis, non permanebitis ".
ISA|7|10|Et adiecit Dominus loqui ad Achaz dicens:
ISA|7|11|" Pete tibi signum a Domino Deo tuo in profundum inferni sive in excelsum supra ".
ISA|7|12|Et dixit Achaz: " Non petam et non tentabo Dominum ".
ISA|7|13|Et dixit: " Audite ergo, domus David; numquid parum vobis est molestos esse hominibus, quia molesti estis et Deo meo?
ISA|7|14|Propter hoc dabit Dominus ipse vobis signum. Ecce, virgo concipiet et pariet filium et vocabit nomen eius Emmanuel;
ISA|7|15|butyrum et mel comedet, ut ipse sciat reprobare malum et eligere bonum.
ISA|7|16|Quia antequam sciat puer reprobare malum et eligere bonum, desolabitur terra, cuius tu formidas duos reges;
ISA|7|17|adducet Dominus super te et super populum tuum et super domum patris tui dies, qui non venerunt a diebus separationis Ephraim a Iuda, regem Assyriorum ".
ISA|7|18|Et erit in die illa:sibilabit Dominus muscae,quae est in extremo fluminum Aegypti,et api, quae est in terra Assur;
ISA|7|19|et venient et requiescent omnesin vallibus praeruptiset in cavernis petrarumet in omnibus frutetiset in omnibus pascuis.
ISA|7|20|In die illa radet Dominusin novacula conducta e regione trans flumenC in rege Assyriorum Ccaput et pilos pedumet barbam quoque abradet.
ISA|7|21|Et erit in die illa:nutriet homo vitulam et duas oves
ISA|7|22|et prae ubertate lactiscomedet butyrum;butyrum enim et mel manducabit omnis,qui relictus fuerit in medio terrae.
ISA|7|23|Et erit in die illa:omnis locus, ubi fuerint mille vites mille argenteis,spinae et vepres erunt.
ISA|7|24|Cum sagittis et arcu ingredientur illuc,vepres enim et spinae erit universa terra.
ISA|7|25|Et in omnes montes, qui in sarculo sarriebantur,nemo veniet prae terrore spinarum et veprium,et erit in pascua bovis et in conculcationem pecoris.
ISA|8|1|Et dixit Dominus ad me: " Sume tibi tabulam grandem et scribe in ea stilo hominis: Maher Salal Has Baz (id est Velociter spolia detrahe, cito praedare).
ISA|8|2|Et adhibui mihi testes fideles, Uriam sacerdotem et Zachariam filium Barachiae;
ISA|8|3|et accessi ad prophetissam, et concepit et peperit filium. Et dixit Dominus ad me: " Voca nomen eius Maher Salal Has Baz,
ISA|8|4|quia antequam sciat puer clamare: "Pater mi" et "Mater mea", afferentur opes Damasci et spolia Samariae coram rege Assyriorum ".
ISA|8|5|Et adiecit Dominus loqui ad me adhuc dicens:
ISA|8|6|" Pro eo quod abiecit populus iste aquas Siloae,quae vadunt cum silentio,et defecit coram Rasin et filio Romeliae,
ISA|8|7|propter hoc ecce Dominus adducet super eosaquas Fluminis fortes et multas,regem Assyriorum et omnem gloriam eius,et ascendet super omnes rivos eiuset fluet super universas ripas eius;
ISA|8|8|et ibit per Iudam inundans et diffluens,usque ad collum veniet.Et erit extensio alarum eiusimplens latitudinem terrae tuae, o Emmanuel ".
ISA|8|9|Clamorem tollite, populi, et consternemini;et audite, universae procul terrae:accingimini et perterremini,accingimini et perterremini.
ISA|8|10|Inite consilium, et dissipabitur;loquimini verbum, et non fiet,quia nobiscum Deus.
ISA|8|11|Haec enim ait Dominus ad me, cum apprehendit me manu et monuit, ne irem in via populi huius, dicens:
ISA|8|12|" Ne vocetis coniurationem,quodcumque populus iste vocat coniurationem,et timorem eius ne timeatis neque paveatis ".
ISA|8|13|Dominum exercituum ipsum sanctificate:ipse pavor vester, et ipse terror vester;
ISA|8|14|et erit in sanctuarium,in lapidem offensionis et in petram scandaliduabus domibus Israel,in laqueum et in insidias habitantibus Ierusalem.
ISA|8|15|Et offendent ex eis plurimiet cadent et conterenturet irretientur et capientur.
ISA|8|16|Liga testimonium, signa legem in discipulis meis.
ISA|8|17|Et exspectabo Dominum, qui abscondit faciem suam a domo Iacob, et praestolabor eum.
ISA|8|18|Ecce ego et pueri, quos dedit mihi Dominus in signum et in portentum Israel a Domino exercituum, qui habitat in monte Sion.
ISA|8|19|Et cum dixerint ad vos: " Quaerite a pythonibus et a divinis, qui susurrant et murmurant; numquid non populus a deo suo requiret, pro vivis a mortuis? ".
ISA|8|20|Ad legem et ad testimonium! Quod si non dixerint iuxta verbum hoc, non erit eis matutina lux.
ISA|8|21|Et transibit per eam afflictus et esuriens;et, cum esurierit, irasceturet maledicet regi suo et deo suoet suspiciet sursum
ISA|8|22|et ad terram intuebitur:et ecce tribulatio et tenebrae,caligo opprimens et obscuritas diffusa.
ISA|8|23|Non erit enim amplius caligo,ubi erat oppressio.Primo tempore contemptibilem reddidit terram Zabulon et terram Nephthali; et novissimo glorificavit viam maris, trans Iordanem, Galilaeam gentium.
ISA|9|1|Populus, qui ambulabat in tenebris,vidit lucem magnam;habitantibus in regione umbrae mortislux orta est eis.
ISA|9|2|Multiplicasti exsultationemet magnificasti laetitiam;laetantur coram tesicut laetantes in messe,sicut exsultant, quando dividunt spolia.
ISA|9|3|Iugum enim oneris eiuset virgam umeri eiuset sceptrum exactoris eiusfregisti, sicut in die Madian.
ISA|9|4|Quia omnis caliga incedentis cum tumultuet vestimentum mixtum sanguineerit in combustionem, cibus ignis.
ISA|9|5|Parvulus enim natus est nobis,filius datus est nobis;et factus est principatus super umerum eius;et vocabitur nomen eiusadmirabilis Consiliarius, Deus fortis,Pater aeternitatis, Princeps pacis.
ISA|9|6|Magnum erit eius imperium,et pacis non erit finissuper solium David et super regnum eius,ut confirmet illud et corroboret in iudicio et iustitiaamodo et usque in sempiternum:zelus Domini exercituum faciet hoc.
ISA|9|7|Verbum misit Dominus in Iacob, et cecidit in Israel.
ISA|9|8|Et sciet omnis populus Ephraim et habitantes Samariamin superbia et magnitudine cordis dicentes:
ISA|9|9|" Lateres ceciderunt, sed quadris lapidibus aedificabimus;sycomori succisae sunt, sed cedris commutabimus ".
ISA|9|10|Et elevavit Dominus hostes super eumet inimicos eius excitavit,
ISA|9|11|Syriam ab oriente et Philisthim ab occidente,qui devoraverunt Israel toto ore.In omnibus his non est aversus furor eius,sed adhuc manus eius extenta.
ISA|9|12|Et populus non est reversus ad percutientem se,et Dominum exercituum non inquisierunt.
ISA|9|13|Et succidit Dominus ab Israel caput et caudam,palmam et arundinem die una:
ISA|9|14|longaevus et honorabilis vultu ipse est caput,et propheta docens mendacium ipse est cauda;
ISA|9|15|rectores populi istius seducenteset, qui regebantur, perierunt.
ISA|9|16|Propter hoc super adulescentulis eius non laetabitur Dominuset pupillorum eius et viduarum non miserebitur,quia omnis impius est et nequam,et universum os loquitur stultitiam.In omnibus his non est aversus furor eius,sed adhuc manus eius extenta.
ISA|9|17|Succensa est enim quasi ignis impietas,veprem et spinam vorat,et succenditur in densitate saltus,et convolvuntur columnae fumi.
ISA|9|18|In ira Domini exercituum incenditur terra;et est populus quasi esca ignis:vir fratri suo non parcit.
ISA|9|19|Et devorat ad dexteram et esuritet comedit ad sinistram et non saturatur;unusquisque carnem proximi sui vorat:
ISA|9|20|Manasses Ephraim, et Ephraim Manassen,simul ipsi contra Iudam.In omnibus his non est aversus furor eius,sed adhuc manus eius extenta.
ISA|10|1|Vae, qui condunt leges iniquaset scribentes iniustitiam scribunt,
ISA|10|2|ut opprimant in iudicio paupereset vim faciant causae humilium populi mei,ut fiant viduae praeda eorum,et pupillos diripiant!
ISA|10|3|Quid facietis in die visitationiset calamitatis de longe venientis?Ad cuius confugietis auxiliumet ubi derelinquetis gloriam vestram?
ISA|10|4|Nam incurvabimini subter captivoset infra occisos cadetis.In omnibus his non est aversus furor eius,sed adhuc manus eius extenta.
ISA|10|5|Vae Assur, virga furoris meiet baculus in manu mea, indignatio mea!
ISA|10|6|Ad gentem impiam mitto eumet contra populum furoris mei mando illi,ut auferat spolia et diripiat praedamet ponat illum in conculcationemquasi lutum platearum.
ISA|10|7|Ipse autem non sic arbitratur,et cor eius non ita existimat;sed in corde suo ad conterendumet ad internecionem gentium non paucarum.
ISA|10|8|Dicet enim: " Numquid non principes mei omnes reges sunt?
ISA|10|9|Numquid non ut Charcamis sic Chalano?Numquid non ut Arphad sic Emath?Numquid non ut Damascus sic Samaria?
ISA|10|10|Quomodo apprehendit manus mea regna idololatra,quorum simulacra plura sunt quam in Ierusalem et in Samaria,
ISA|10|11|numquid non sicut feci Samariae et idolis eius,sic faciam Ierusalem et simulacris eius? ".
ISA|10|12|Et erit: cum impleverit Dominus cuncta opera sua in monte Sion et in Ierusalem, visitabo super fructum superbiae cordis regis Assyriae et super arrogantiam altitudinis oculorum eius.
ISA|10|13|Dixit enim: In fortitudine manus meae feciet in sapientia mea, prudens sum enim;et abstuli terminos populorumet scrinia eorum depraedatus sumet detraxi quasi potens in sublimi sedentes;
ISA|10|14|et apprehendit quasi nidum manus mea fortitudinem populorum;et sicut colliguntur ova derelicta,sic universam terram ego congregavi,et non fuit qui moveret pennam aut aperiret os et ganniret ".
ISA|10|15|Numquid gloriabitur securiscontra eum, qui secat in ea?Aut exaltabitur serracontra eum, qui trahit eam?Quomodo si agitet virga elevantem eam,et exaltet baculus eum, qui non est lignum.
ISA|10|16|Propter hoc mittet Dominator, Dominus exercituum,in pingues eius tenuitatem;et subtus gloriam eiusardor ardebit quasi combustio ignis.
ISA|10|17|Et erit Lumen Israel ignis,et Sanctus eius flamma;et succendetur et devorabit spinas eiuset vepres in die una.
ISA|10|18|Et gloriam saltus eius et horti eiusab anima usque ad carnem consumet,et erit sicut aeger tabescens;
ISA|10|19|et reliquiae ligni saltus eiustam paucae erunt,ut puer scribat ea.
ISA|10|20|Et erit in die illa:non adiciet residuum Israelet, qui effugerint de domo Iacob,inniti super eo, qui percutit eos,sed innitentur super Dominum,Sanctum Israel, in veritate.
ISA|10|21|Reliquiae revertentur,reliquiae, inquam, Iacob, ad Deum fortem.
ISA|10|22|Si enim fuerit populus tuus, Israel, quasi arena maris,reliquiae revertentur ex eo;consummatio decreta redundat in iustitia:
ISA|10|23|interitum enim, qui decretus est,Dominus, Deus exercituum, faciet in medio omnis terrae.
ISA|10|24|Propter hoc haec dicit Dominus, Deus exercituum: " Noli timere, populus meus habitator Sion, ab Assur; in virga percutiet te et baculum suum levabit super te sicut Aegyptus.
ISA|10|25|Adhuc enim paululum modicumque, et consummabitur indignatio et furor meus ad destructionem eorum ".
ISA|10|26|Et suscitabit super eum Dominus exercituum flagellum iuxta plagam Madian in Petra Oreb et virgam suam super mare et levabit eam sicut in Aegypto.
ISA|10|27|Et erit in die illa:auferetur onus eius de umero tuo,et iugum eius de collo tuo.Et vastator ascendit a Remmon.
ISA|10|28|Veniet in Aiath, transibit per Magron,apud Machmas deponit sarcinas suas;
ISA|10|29|transeunt vadum cursim; in Geba pernoctabimus;trepidat Rama, Gabaa Saulis fugit.
ISA|10|30|Hinni voce tua, Bathgallim;attende, Laisa; responde, Anathoth.
ISA|10|31|Migrat Medemena, habitatores Gabim fugiunt;
ISA|10|32|hodie in Nob stabit:agitabit manum suam ad montem filiae Sion,collem Ierusalem.
ISA|10|33|Ecce Dominator, Dominus exercituum,amputat ramos in terrore,et extrema acumina succiduntur,et sublimes humiliantur;
ISA|10|34|et caeduntur condensa saltus ferro,et Libanus cum excelsis suis cadet.
ISA|11|1|Et egredietur virga de stirpe Iesse,et flos de radice eius ascendet;
ISA|11|2|et requiescet super eum spiritus Domini:spiritus sapientiae et intellectus,spiritus consilii et fortitudinis,spiritus scientiae et timoris Domini;
ISA|11|3|et deliciae eius in timore Domini.Non secundum visionem oculorum iudicabitneque secundum auditum aurium decernet;
ISA|11|4|sed iudicabit in iustitia paupereset decernet in aequitate pro mansuetis terrae;et percutiet terram virga oris suiet spiritu labiorum suorum interficiet impium.
ISA|11|5|Et erit iustitia cingulum lumborum eius,et fides cinctorium renum eius.
ISA|11|6|Habitabit lupus cum agno,et pardus cum haedo accubabit;vitulus et leo simul saginabuntur,et puer parvulus minabit eos.
ISA|11|7|Vitula et ursus pascentur,simul accubabunt catuli eorum;et leo sicut bos comedet paleas.
ISA|11|8|Et ludet infans ab uberesuper foramine aspidis;et in cavernam reguli,qui ablactatus fuerit, manum suam mittet.
ISA|11|9|Non nocebunt et non occidentin universo monte sancto meo,quia plena erit terra scientia Domini, sicut aquae mare operiunt.
ISA|11|10|In die illa radix Iessestat in signum populorum;ipsam gentes requirent,et erit sedes eius gloriosa.
ISA|11|11|Et erit in die illa: rursus extendet Dominus manum suamad possidendum residuum populi sui,quod relictum erit ab Assyria et ab Aegyptoet a Phatros et ab Aethiopiaet ab Elam et a Sennaaret ab Emath et ab insulis maris;
ISA|11|12|et levabit signum in nationeset congregabit profugos Israelet dispersos Iudae colliget a quattuor plagis terrae.
ISA|11|13|Et auferetur zelus Ephraim,et hostes Iudae abscindentur;Ephraim non aemulabitur Iudam, et Iudas non pugnabit contra Ephraim.
ISA|11|14|Et volabunt in umeros Philisthim ad mare,simul praedabuntur filios orientis:in Edom et Moab extendent manus suas,et filii Ammon oboedient eis.
ISA|11|15|Et exsiccabit Dominus linguam maris Aegyptiet levabit manum suam super flumen in fortitudine spiritus suiet percutiet illud in septem rivos,ita ut transire faciat eos calceatos.
ISA|11|16|Et erit via residuo populo meo,qui relinquetur ab Assyria,sicut fuit Israeli in die illa,qua ascendit de terra Aegypti.
ISA|12|1|Et dices in die illa: Confitebor tibi, Domine,quoniam cum iratus eras mihi,conversus est furor tuus, et consolatus es me.
ISA|12|2|Ecce Deus salutis meae;fiducialiter agam et non timebo,quia fortitudo mea et laus mea Dominus,et factus est mihi in salutem ".
ISA|12|3|Et haurietis aquas in gaudio de fontibus salutis.
ISA|12|4|Et dicetis in die illa: Confitemini Domino et invocate nomen eius,notas facite in populis adinventiones eius;mementote quoniam excelsum est nomen eius.
ISA|12|5|Cantate Domino, quoniam magnifice fecit;notum sit hoc in universa terra.
ISA|12|6|Exsulta et lauda, quae habitas in Sion,quia magnus in medio tui Sanctus Israel ".
ISA|13|1|Oraculum Babylonis, quod vidit Isaias filius Amos.
ISA|13|2|Super montem decalvatum levate signum,exaltate vocem, levate manum,et ingrediantur portas ducum.
ISA|13|3|Ego mandavi sanctificatis meiset vocavi fortes meos ad iram meam,exsultantes in gloria mea.
ISA|13|4|Vox multitudinis in montibus quasi populi ingentis,vox sonitus regnorum gentium congregatarum.Dominus exercituum recenset militiam belli;
ISA|13|5|veniunt de terra procul a termino caeli,Dominus et vasa furoris eius,ut disperdat omnem terram.
ISA|13|6|Ululate, quia prope est dies Domini;quasi vastitas a Domino veniet.
ISA|13|7|Propter hoc omnes manus dissolventur,et omne cor hominis tabescet.
ISA|13|8|Perterrebuntur.Torsiones et dolores tenebunt eos,quasi parturiens dolebunt;unusquisque ad proximum suum stupebit:facies combustae vultus eorum.
ISA|13|9|Ecce dies Domini venit,crudelis et indignationis plenuset irae furorisque,ad ponendam terram in solitudinem,et peccatores eius conteret de ea.
ISA|13|10|Quoniam stellae caeli et sidera eiusnon expandent lumen suum;obtenebratus est sol in ortu suo,et luna non splendebit in lumine suo.
ISA|13|11|Et visitabo super orbem propter malaet super impios propter iniquitatem eorum;et quiescere faciam superbiam protervorumet arrogantiam fortium humiliabo.
ISA|13|12|Pretiosior erit vir auro,et homo mundo obryzo.
ISA|13|13|Super hoc caelum turbabo,et movebitur terra de loco suoin indignatione Domini exercituumet in die irae furoris eius.
ISA|13|14|Et erit quasi damula fugiens et quasi ovis,et non erit qui congreget;unusquisque ad populum suum convertetur,et singuli ad terram suam fugient.
ISA|13|15|Omnis, qui inventus fuerit, occidetur,et omnis, qui captus fuerit, cadet in gladio;
ISA|13|16|infantes eorum allidentur in oculis eorum,diripientur domus eorum,et uxores eorum violabuntur.
ISA|13|17|Ecce ego suscitabo super eos Medos,qui argentum non quaerant nec aurum velint;
ISA|13|18|sed arcus pueros prosternentet fructui uteri non miserebuntur.
ISA|13|19|Et erit Babylon, splendor regnorum,inclita superbia Chaldaeorum,sicut cum subvertit Dominus Sodomam et Gomorram.
ISA|13|20|Non habitabitur usque in finemet non fundabitur usque ad generationem et generationem,nec ponet ibi tentoria Arabs,nec pastores accubare facient ibi,
ISA|13|21|sed accubabunt ibi bestiae,et replebunt domus eorum ululae,et habitabunt ibi struthiones,et pilosi saltabunt ibi;
ISA|13|22|et respondebunt ibi hyaenae in aedibus eius,et thoes in delubris voluptatis.Prope est ut veniat tempus eius,et dies eius non elongabuntur.
ISA|14|1|Miserebitur enim Dominus Iacobet eliget adhuc de Israelet requiescere eos faciet super humum suam;adiungetur advena ad eoset adhaerebit domui Iacob.
ISA|14|2|Et tenebunt eos populiet adducent eos in locum suum;et possidebit eos domus Israelsuper terram Domini in servos et ancillas;et erunt capientes eos, qui se ceperant,et subicient exactores suos.
ISA|14|3|Et erit in die illa:cum requiem dederit tibi Dominusa labore tuo et a concussione tuaet a servitute dura, qua ante servisti,
ISA|14|4|proferes parabolam istam contra regem Babylonis et dices: Quomodo cessavit exactor, quievit oppressio?
ISA|14|5|Contrivit Dominus baculum impiorum,virgam dominantium,
ISA|14|6|caedentem populos in indignatione plaga sine remissione,subicientem in furore gentes persecutione sine fine.
ISA|14|7|Conquievit et siluit omnis terra,gavisa est, et exsultaverunt.
ISA|14|8|Abietes quoque laetatae sunt super te, et cedri Libani:Ex quo dormisti, non ascendit, qui succidat nos".
ISA|14|9|Infernus subter conturbatus estin occursum adventus tui;suscitat tibi umbras, omnes principes terraesurgere fecit de soliis suis,omnes reges nationum.
ISA|14|10|Universi respondebunt et dicent tibi:Et tu vulneratus es sicut nos,nostri similis effectus es".
ISA|14|11|Detracta est ad inferos superbia tua,sonitus nablorum tuorum;subter te sternitur tinea,et operimentum tuum sunt vermes.
ISA|14|12|Quomodo cecidisti de caelo, lucifer, fili aurorae?Deiectus es in terram, qui deiciebas gentes,
ISA|14|13|qui dicebas in corde tuo:In caelum conscendam,super astra Dei exaltabo solium meum,sedebo in monte conventusin lateribus aquilonis;
ISA|14|14|ascendam super altitudinem nubium,similis ero Altissimo".
ISA|14|15|Verumtamen ad infernum detractus es,in profundum laci.
ISA|14|16|Qui te viderint, te intuenturteque prospicient:Numquid iste est vir, qui conturbavit terram,qui concussit regna,
ISA|14|17|qui posuit orbem desertumet urbes eius destruxit,vinctis eius non aperuit carcerem?
ISA|14|18|Omnes reges gentium universi dormiunt in gloria,vir in domo sua;
ISA|14|19|tu autem proiectus es de sepulcro tuoquasi stirps abominabilis,obvolutus cum his, qui interfecti sunt gladioet descenderunt ad lapides sepulcri,quasi cadaver conculcatum.
ISA|14|20|Non habebis consortium cum eis in sepultura;tu enim terram tuam disperdidisti,tu populum tuum occidisti:non vocabitur in aeternum semen malefactorum.
ISA|14|21|Praeparate filios eius occisioniob iniquitatem patrum suorum;ne consurgant, ut hereditent terram,neque impleant faciem orbis civitatum" ".
ISA|14|22|" Et consurgam contra eos,dicit Dominus exercituum;et perdam Babylonis nomen et reliquiaset germen et progeniem, dicit Dominus;
ISA|14|23|et ponam eam in possessionem ericiiet in paludes aquarum,et scopabo eam in scopa destructionis ",dicit Dominus exercituum.
ISA|14|24|Iuravit Dominus exercituum dicens: Profecto, ut putavi, ita erit;et quomodo mente tractavi, sic eveniet.
ISA|14|25|Conteram Assyrium in terra meaet in montibus meis conculcabo eum;et auferetur ab eis iugum eius,et onus illius ab umero eorum tolletur ".
ISA|14|26|Hoc consilium, quod initum estsuper omnem terram,et haec est manus extentasuper universas gentes.
ISA|14|27|Dominus enim exercituum decrevit,et quis poterit infirmare?Et manus eius extenta,et quis avertet eam?
ISA|14|28|In anno, quo mortuus est rex Achaz, factum est oraculum istud:
ISA|14|29|" Ne laeteris, Philisthaea omnis tu,quoniam comminuta est virga percussoris tui;de radice enim colubri egredietur regulus,et semen eius draco volans.
ISA|14|30|Et pascentur primogeniti egenorum,et pauperes fiducialiter requiescent;et interire faciam in fame radicem tuamet reliquias tuas interficiam.
ISA|14|31|Ulula, porta! Clama, civitas!Contremisce, Philisthaea omnis;ab aquilone enim fumus venit,et non est fugitivus in agminibus eius ".
ISA|14|32|Et quid respondebitur nuntiis gentis? Quia Dominus fundavit Sion,et in ipsam confugiunt pauperes populi eius ".
ISA|15|1|Oraculum Moab.Quia nocte vastata est Ar moab, conticuit;quia nocte vastata est Cirmoab, conticuit.
ISA|15|2|Ascendit filia Dibon ad excelsa in planctum;super Nabo et super Medaba Moab ululavit;in cunctis capitibus eius calvitium, omnis barba rasa.
ISA|15|3|In triviis eius accincti sunt sacco;super tecta eius et in plateis eiusomnes ululant, prorumpunt in fletum.
ISA|15|4|Clamat Hesebon et Eleale,usque Iasa auditur vox eorum;super hoc expediti Moab fremunt,anima eius fremit sibi.
ISA|15|5|Cor meum super Moab clamat,vectes eius usque ad Segor, Eglatselisiam;per ascensum enim Luith flentes ascenduntet in via Oronaim clamorem contritionis levant.
ISA|15|6|Aquae enim Nemrim desertae erunt,quia aruit herba, defecit germen,viror omnis interiit.
ISA|15|7|Ideo supellectiles colligunt, copias divitiarum suastrans torrentem Salicum ducunt.
ISA|15|8|Quoniam circuivit clamor terminum Moab;usque ad Eglaim ululatus eius,et usque ad Beerelim clamor eius.
ISA|15|9|Quia aquae Dimon repletae sunt sanguine;ponam enim super Dimon additamentahis, qui fugerint de Moab leonem, et reliquiis terrae.
ISA|16|1|Emittite agnum dominatori terraede Petra deserti ad montem filiae Sion.
ISA|16|2|Et erit: sicut avis fugiens,et pulli de nido avolantes,sic erunt filiae Moabad vada Arnon.
ISA|16|3|Affer consilium, fac iudicium;pone quasi noctem umbram tuam in meridie,absconde fugientes et vagos ne prodas.
ISA|16|4|Habitent apud te profugi Moab;esto latibulum eorum a facie vastatoris;finitus est enim exactor,consummata est devastatio,defecit calcator a terra.
ISA|16|5|Et firmabitur in misericordia solium;et sedebit super illud in veritate,in tabernaculo David, iudicans et quaerens iudiciumet velociter reddens, quod iustum est.
ISA|16|6|Audivimus superbiam MoabC superbus est valde Csuperbiam eius et arrogantiam eius et indignationem eiuset iactantiam eius non rectam.
ISA|16|7|Idcirco ululabit Moab super Moab,omnes ululabunt;super placentas Cirharesethlamentantur percussi.
ISA|16|8|Quoniam suburbana Hesebon deserta sunt et vinea Sabama;dominos gentium perdiderunt uvae eius;usque ad Iazer pervenerunt,erraverunt in deserto:propagines eius diffusae sunt,transierunt mare.
ISA|16|9|Super hoc plorabo in fletu Iazer vineam Sabama;inebriabo te lacrima mea, Hesebon et Eleale,quoniam super vindemiam tuam et super messem tuamclamor cecidit.
ISA|16|10|Et ablata est laetitia et exsultatio de hortis,et in vineis non exsultant neque iubilant.Vinum in torculari non calcabit, qui calcare consueverat;clamor cessavit.
ISA|16|11|Ideo venter meus super Moab quasi cithara fremit,et viscera mea super Cirhareseth.
ISA|16|12|Et erit: cum apparueritet laboraverit Moab super excelsis,ingredietur ad sancta sua, ut obsecret,et non valebit.
ISA|16|13|Et hoc verbum, quod locutus est Dominus ad Moab ex tunc;
ISA|16|14|nunc autem loquitur Dominus dicens: " In tribus annis, quasi anni mercennarii, auferetur gloria Moab cum omni populo multo, et residuum parvum et modicum nequaquam ingens erit ".
ISA|17|1|Oraculum Damasci. Ecce Damascus desinet esse civitaset erit sicut acervus ruinarum.
ISA|17|2|Derelictae civitates Aroer gregibus erunt;et requiescent ibi, et non erit qui exterreat.
ISA|17|3|Et auferetur munimentum ab Ephraimet regnum a Damasco,et reliquiae Syriae sicut gloria filiorum Israel erunt,dicit Dominus exercituum.
ISA|17|4|Et erit in die illa: attenuabitur gloria Iacob,et pinguedo carnis eius marcescet;
ISA|17|5|et erit, sicut cum messor arripit culmos,et brachium eius spicas legit;et erit, sicut cum quis quaerit spicas in valle Raphaim.
ISA|17|6|Et relinquetur in eo racemus,et sicut cum excutitur olea:duae vel tres olivae in summitate ramisive quattuor aut quinque in cacuminibus arboris fructiferae ",dicit Dominus Deus Israel.
ISA|17|7|In die illa attendet homo ad factorem suum,et oculi eius ad Sanctum Israel respicient;
ISA|17|8|et non attendet ad altaria,quae fecerunt manus eius,et quae operati sunt digiti eius;non respiciet lucos et thymiateria.
ISA|17|9|In die illa erunt civitates fortitudinis eius derelictae,sicut civitates, quas dereliquerunt Hevaei et Amorraeia facie filiorum Israel;et erit desolatio,
ISA|17|10|quia oblita es Dei salutis tuaeet petrae fortitudinis tuae non es recordata:propterea plantabis plantationes iucundaset germen alienum seminabis.
ISA|17|11|In ipso die plantationis tuae saepies easet mane semen tuum florere facies;evanescet messis in die penuriae,et dolor insanabilis erit.
ISA|17|12|Heu!, strepitus populorum multorum;strepunt quasi strepitu maris,et tumultus turbarumquasi sonitu aquarum sonabunt.
ISA|17|13|Sonabunt populi sicut sonitus aquarum inundantium,et increpabit eum, et fugiet procul;et rapietur sicut pulvis montium a facie ventiet sicut turbo coram tempestate.
ISA|17|14|In tempore vespere, et ecce turbatio,ante matutinum non subsistet:haec est pars eorum, qui vastaverunt nos,et sors diripientium nos.
ISA|18|1|Vae terrae alarum strepitantium,quae est trans flumina Aethiopiae!
ISA|18|2|Quae mittit in mari legatoset in vasis papyri super aquas: Ite, nuntii veloces,ad gentem proceram et lucidam,ad populum terribilem,prope et procul,gentem robustam et conculcantem,cuius flumina scindunt terram ".
ISA|18|3|Omnes habitatores orbiset in terra commorantes,cum elevatum fuerit signum in montibus, videbitiset, cum clanguerit tuba, audietis.
ISA|18|4|Quia haec dixit Dominus ad me: Quiescam et considerabo in loco meo,sicut calor torrens orta iam luceet sicut nubes roris in aestu messis ".
ISA|18|5|Etenim ante vindemiam, cum consummatus fuerit flos,et uva germinans maturescens erit,praecidet ramusculos falcibuset propagines abscindet et proiciet;
ISA|18|6|et relinquentur simul avibus montiumet bestiis terrae;et aestate erunt super ea volucres,et omnes bestiae terrae super illa hiemabunt.
ISA|18|7|In tempore illo deferetur munus Domino exercituum a populo procero et lucido, a populo terribili, prope et procul, a gente robusta et conculcante, cuius terram flumina scindunt, ad locum nominis Domini exercituum, montem Sion.
ISA|19|1|Oraculum Aegypti.Ecce Dominus vehitur super nubem levemet ingreditur Aegyptum;et commovebuntur simulacra Aegypti a facie eius,et cor Aegypti tabescet in medio eius.
ISA|19|2|" Et concurrere faciam Aegyptios adversus Aegyptios;et pugnabit vir contra fratrem suum,et vir contra amicum suum,civitas adversus civitatem,regnum adversus regnum.
ISA|19|3|Et dirumpetur spiritus Aegypti in visceribus eius,et consilium eius confundam;et interrogabunt simulacra et divinoset pythones et hariolos.
ISA|19|4|Et tradam Aegyptios in manu domini crudelis,et rex fortis dominabitur eorum ",ait Dominus, Deus exercituum.
ISA|19|5|Et arescet aqua de mari,et fluvius desolabitur atque siccabitur,
ISA|19|6|et putrida fient flumina;attenuabuntur et siccabuntur rivi Aegypti,calamus et iuncus marcescent;
ISA|19|7|nudabuntur ripae Nili,et omnis planta Nili siccabitur;arescet et non erit.
ISA|19|8|Et maerebunt piscatores,et lugebunt omnes mittentes in flumen hamum;et expandentes rete super faciem aquarum languebunt.
ISA|19|9|Confundentur, qui operantur linum,pectentes et texentes byssum.
ISA|19|10|Et opifices eius deprimentur,omnes mercennarii omnino deficient.
ISA|19|11|Quam stulti principes Taneos!Sapientes consiliarii pharaonis dederunt consilium insipiens;quomodo dicetis pharaoni: Filius sapientium ego, filius regum antiquorum "?
ISA|19|12|Ubi nunc sunt sapientes tui?Annuntient tibi et indicentquid cogitaverit Dominus exercituum super Aegyptum.
ISA|19|13|Stulti facti sunt principes Taneos,decepti sunt principes Mempheos,deceperunt Aegyptum anguli tribuum eius.
ISA|19|14|Dominus miscuit in medio eius spiritum vertiginis,et errare fecerunt Aegyptum in omni opere suo,sicut errat ebrius in vomitu suo;
ISA|19|15|et non erit Aegypto opus,quod faciat, caput vel cauda, palma vel arundo.
ISA|19|16|In die illa erunt Aegyptii quasi mulieres et stupebunt et timebunt a facie commotionis manus Domini exercituum, quam ipse movebit super eam.
ISA|19|17|Et erit terra Iudae Aegypto in pavorem: omnis, qui illius fuerit recordatus, pavebit a facie consilii Domini exercituum, quod ipse cogitavit super eam.
ISA|19|18|In die illa erunt quinque civitates in terra Aegypti loquentes lingua Chanaan et iurantes per Dominum exercituum. Civitas Solis vocabitur una.
ISA|19|19|In die illa erit altare Domino in medio terrae Aegypti, et titulus iuxta terminum eius Domino.
ISA|19|20|Et erit in signum et in testimonium Domino exercituum in terra Aegypti. Clamabunt enim ad Dominum a facie tribulantium, et mittet eis salvatorem et propugnatorem, qui liberet eos.
ISA|19|21|Et cognoscetur Dominus ab Aegypto, et cognoscent Aegyptii Dominum in die illa; et colent eum in hostiis et in muneribus et vota vovebunt Domino et solvent.
ISA|19|22|Et percutiet Dominus Aegyptum plaga et sanabit; et revertentur ad Dominum, et placabitur eis et sanabit eos.
ISA|19|23|In die illa erit via de Aegypto in Assyriam; et intrabit Assyrius Aegyptum, et Aegyptius in Assyriam, et servient Aegyptii cum Assyriis.
ISA|19|24|In die illa erit Israel tertius cum Aegypto et Assyria; benedictio in medio terrae,
ISA|19|25|cui benedicet Dominus exercituum dicens: " Benedictus populus meus Aegyptius, et opus manuum mearum Assyrius, et hereditas mea Israel ".
ISA|20|1|In anno quo ingressus est Tharthan in Azotum, cum misisset eum Sargon rex Assyriorum, et pugnasset contra Azotum et cepisset eam,
ISA|20|2|in tempore illo locutus est Dominus in manu Isaiae filii Amos dicens: " Vade et solve saccum de lumbis tuis et calceamenta tua tolle de pedibus tuis ". Et fecit sic, vadens nudus et discalceatus.
ISA|20|3|Et dixit Dominus: " Sicut ambulavit servus meus Isaias nudus et discalceatus tribus annis signum et portentum super Aegyptum et super Aethiopiam,
ISA|20|4|sic minabit rex Assyriorum captivos Aegypti et exsules Aethiopiae, iuvenes et senes, nudos et discalceatos, discoopertis natibus ad ignominiam Aegypti.
ISA|20|5|Et timebunt et confundentur ab Aethiopia spe sua et ab Aegypto gloria sua.
ISA|20|6|Et dicet habitator maritimae regionis huius in die illa: "Ecce, haec erat spes nostra, quo confugimus in auxilium, ut liberaremur a facie regis Assyriorum; et quomodo effugere poterimus nos?" ".
ISA|21|1|Oraculum deserti maris.Sicut turbines per austrum transeuntes,de deserto venit, de terra horribili.
ISA|21|2|Visio dura nuntiata est mihi:praedo praedatur,et vastator vastat.Ascende, Elam;obside, Media;omnem gemitum eius cessare feci.
ISA|21|3|Propterea repleti sunt lumbi mei tremore,angustia possedit me sicut angustia parientis;corrui, cum audirem;conturbatus sum, cum viderem.
ISA|21|4|Vacillat cor meum,pavor invadit me:crepusculum optatumposuit mihi in terrorem.
ISA|21|5|Ponunt mensam,stragulum pandunt, comedunt, bibunt.Surgite, principes,ungite clipeum.
ISA|21|6|Haec enim dixit mihi Dominus: Vade et pone speculatorem;quodcumque viderit, annuntiet.
ISA|21|7|Si viderit currum, bigam equitum,ascensorem asini et ascensorem cameli,intueatur diligenter multo intuitu ".
ISA|21|8|Et clamavit speculator: Super specula, Domine,ego sum stans iugiter per diem,et super custodiam meamego sum stans totis noctibus.
ISA|21|9|Ecce, huc venit agmen virorum,biga equitum ".Et respondit et dixit: Cecidit, cecidit Babylon,et omnia sculptilia deorum eiuscontrita sunt in terram ".
ISA|21|10|Tritura mea et fili areae meae,quae audivi a Domino exercituum, Deo Israel,annuntiavi vobis.
ISA|21|11|Oraculum Duma.Ad me clamat ex Seir: Custos, quid de nocte?Custos, quid de nocte? ".
ISA|21|12|Dixit custos: Venit mane, sed etiam nox;si quaeritis, quaerite,revertimini, venite ".
ISA|21|13|Oraculum in solitudine.In saltu, in solitudine dormietis,turmae Dedanim.
ISA|21|14|Occurrentes sitienti ferte aquam,qui habitatis terram Thema;cum panibus occurrite fugienti:
ISA|21|15|a facie enim gladiorum fugerunt,a facie gladii nudati,a facie arcus extenti,a facie gravis proelii.
ISA|21|16|Quoniam haec dicit Dominus ad me: " Adhuc anno sicut anni mercennarii, et auferetur omnis gloria Cedar;
ISA|21|17|et reliquiae numeri arcuum fortium filiorum Cedar imminuentur; Dominus enim, Deus Israel, locutus est ".
ISA|22|1|Oraculum vallis Visionis.Quidnam tibi est,quia ascendisti omnis in tecta,
ISA|22|2|clamoris plena, urbs tumultuans,civitas exsultans?Interfecti tui non interfecti gladionec mortui in bello;
ISA|22|3|cuncti principes tui fugeruntsimul sine arcu capti;omnes, qui inventi sunt, capti sunt simul,procul fugerunt.
ISA|22|4|Propterea dixi: " Recedite a me,amare flebo;nolite incumbere, ut consolemini mesuper vastitate filiae populi mei ".
ISA|22|5|Dies enim confusioniset conculcationis et fletusDomino, Deo exercituum, in valle Visionis,eversio murorum et vociferatio ad montem.
ISA|22|6|Et Elam sumpsit pharetram,in agmine hominum equitum,et Cir nudavit clipeum.
ISA|22|7|Et electae valles tuaeplenae sunt quadrigarum,et equites ponunt sedes suas in porta.
ISA|22|8|Et revelatum est operimentum Iudae,et respexisti in die illa armamentarium domus Saltus;
ISA|22|9|et scissuras civitatis David vidistis,quia multiplicatae sunt;et congregastis aquas piscinae inferioris.
ISA|22|10|Et domos Ierusalem numerastiset destruxistis domosad muniendum murum;
ISA|22|11|et lacum fecistis inter duos murospro aqua piscinae veteris;sed non suspexistis ad eum, qui fecit haec,et eum, qui haec de longe formavit, non vidistis.
ISA|22|12|Et vocavit Dominus, Deus exercituum, in die illaad fletum et ad planctum,ad calvitium et ad cingendum saccum;
ISA|22|13|et ecce gaudium et laetitia,occidere boves et iugulare pecus,comedere carnes et bibere vinum: Comedamus et bibamus,cras enim moriemur ".
ISA|22|14|Et revelatum est in auribus meisa Domino exercituum: Certe non dimittetur iniquitas haec vobis, donec moriamini! ",dicit Dominus, Deus exercituum.
ISA|22|15|Haec dicit Dominus, Deus exercituum: Vade, ingredere ad procuratorem istum,ad Sobnam praepositum palatii:
ISA|22|16|"Quid tibi hic? Aut quis tibi hic,quia excidisti tibi hic sepulcrum?".Effodiens in excelso sepulcrum suum,excavabat in petra tabernaculum sibi.
ISA|22|17|Ecce Dominus vehementer proiciet te, homo,violenter te apprehendens.
ISA|22|18|In globum te convolvet glomerans;quasi pilam mittet tein terram latam et spatiosam:ibi morieris,et ibi erunt currus gloriae tuae,ignominia domus domini tui.
ISA|22|19|Et expellam te de statione tuaet de ministerio tuo deponam te.
ISA|22|20|Et erit in die illa:vocabo servum meum Eliachim filium Helciae
ISA|22|21|et induam illum tunicam tuamet cingulo tuo cingam eumet potestatem tuam dabo in manu eius;et erit in patrem habitantibus Ierusalemet domui Iudae.
ISA|22|22|Et dabo clavem domus Davidsuper umerum eius;et aperiet, et non erit qui claudat;et claudet, et non erit qui aperiat.
ISA|22|23|Et figam illum paxillum in loco securo,et erit in solium gloriae domui patris sui.
ISA|22|24|Et suspendent super eum omnem gloriam domus patris sui, propagines et stirpes, omne vas parvulum, a pelvibus ad amphoras.
ISA|22|25|In die illa, dicit Dominus exercituum, auferetur paxillus, qui fixus fuerat in loco securo, et frangetur et cadet; et peribit, quod pependerat in eo, quia Dominus locutus est ".
ISA|23|1|Oraculum Tyri.Ululate, naves Tharsis,quia vastatum est refugium vestrum;cum redirent de terra Cetthim, revelatum est eis.
ISA|23|2|Obstupescite, qui habitatis in insula;negotiatores Sidonistransfretantes mare repleverunt te.
ISA|23|3|In aquis multis semen Nili,messis fluminis fruges eius;et facta est negotiatio gentium.
ISA|23|4|Erubesce, Sidon, ait enim mare,fortitudo maris, dicens: Non parturivi et non peperi;et non enutrivi iuvenesnec virgines educavi ".
ISA|23|5|Cum auditum fuerit in Aegypto,dolebunt cum audierint de Tyro.
ISA|23|6|Transite ad Tharsis,ululate, qui habitatis in insula.
ISA|23|7|Estne vestra haec, quae gloriabatur?A diebus pristinis antiquitas eius.Ducebant eam pedes sui longead peregrinandum.
ISA|23|8|Quis cogitavit hocsuper Tyrum quondam coronatam,cuius negotiatores principes,institores eius incliti terrae?
ISA|23|9|Dominus exercituum cogitavit hoc,ut detraheret superbiam omnis gloriaeet viles faceret universos inclitos terrae.
ISA|23|10|Excole terram tuam sicut litus Nili,filia Tharsis, iam non est portus.
ISA|23|11|Manum suam extendit super mare,conturbavit regna.Dominus mandavit adversus Chanaan,ut contereret munimenta eius,
ISA|23|12|et dixit: " Non adicies ultra ut glorieris,violata virgo filia Sidonis;in Cetthim consurgens transfreta:ibi quoque non erit requies tibi ".
ISA|23|13|Ecce terra Chaldaeorum:talis populus non fuit;Assyria fundavit eam pro feris.Erexerunt turres suas;suffoderunt domos eius,posuerunt eam in ruinam.
ISA|23|14|Ululate, naves Tharsis,quia devastatum est praesidium vestrum.
ISA|23|15|Et erit in die illa: in oblivione erit Tyrus septuaginta annis, sicut dies regis unius. Post septuaginta autem annos erit Tyro iuxta canticum meretricis:
ISA|23|16|" Sume citharam, circui civitatem,meretrix oblivioni tradita;bene cane, frequenta canticum,ut memoria tui sit ".
ISA|23|17|Et erit: post septuaginta annos visitabit Dominus Tyrum, et redibit ad mercedes suas et rursum fornicabitur cum universis regnis terrae super faciem terrae.
ISA|23|18|Et erunt negotiatio eius et merces eius sanctificatae Domino; non condentur neque reponentur, quia his, qui habitaverint coram Domino, erit negotiatio eius, ut manducent in saturitate et vestiantur splendide.
ISA|24|1|Ecce Dominus dissipat terram et frangit eamet conturbat faciem eiuset dispergit habitatores eius.
ISA|24|2|Et erit sicut populus sic sacerdos,et sicut servus sic dominus eius,sicut ancilla sic domina eius,sicut emens sic ille qui vendit,sicut fenerator sic is qui mutuum accipit,sicut qui repetit sic qui debet.
ISA|24|3|Dissipatione dissipabitur terraet direptione praedabitur:Dominus enim locutus est verbum hoc.
ISA|24|4|Luget, languet terra,marcescit, languet orbis,marcescit altitudo simul cum terra.
ISA|24|5|Et terra infecta est sub habitatoribus suis,quia transgressi sunt leges,violaverunt mandatum,dissipaverunt foedus sempiternum.
ISA|24|6|Propter hoc maledictio voravit terram,et poenas exsolverunt habitatores eius;ideoque imminuti sunt cultores eius,et relicti sunt homines pauci.
ISA|24|7|Luget mustum,emarcuit vitis,ingemiscunt omnes, qui laetabantur corde.
ISA|24|8|Cessavit gaudium tympanorum,quievit sonitus laetantium,cessavit gaudium citharae;
ISA|24|9|cum cantico non bibent vinum,amara erit potio bibentibus illam.
ISA|24|10|Attrita est civitas inanitatis,clausa est omnis domus, ut nemo introeat;
ISA|24|11|clamor est super vino in plateis,occidit omnis laetitia,translatum est gaudium terrae.
ISA|24|12|Relicta est in urbe solitudo,et in ruinam confracta est porta;
ISA|24|13|quia haec erunt in medio terrae,in medio populorum,quomodo si olivae excutiantur,et finita vindemia colligantur racemi.
ISA|24|14|Hi levabunt vocem suam,laudabunt maiestatem Domini,hinnient de mari.
ISA|24|15|Propter hoc in regionibus lucis glorificate Dominum,in insulis maris nomen Domini, Dei Israel.
ISA|24|16|A finibus terrae laudes audivimus: Gloria iusto ".Et dixi: " Secretum meum mihi,secretum meum mihi.Vae mihi! ".Praevaricantes praevaricati suntet praevaricatione praevaricantium praevaricati sunt.
ISA|24|17|Formido et fovea et laqueus super te,habitator terrae.
ISA|24|18|Et erit: qui fugerit a voce formidinis, cadet in foveam;et, qui ascenderit de fovea,tenebitur laqueo,quia cataractae de excelsis apertae sunt,et concussa sunt fundamenta terrae.
ISA|24|19|Confractione confracta est terra,contritione contrita est terra,commotione commota est terra,
ISA|24|20|agitatione agitabitur terra sicut ebriuset fluctuabit quasi tabernaculum;et gravis erit super eam iniquitas eius,et corruet et non adiciet ut resurgat.
ISA|24|21|Et erit in die illa:visitabit Dominus super militiam caeli in excelsoet super reges terrae super terram;
ISA|24|22|et congregabuntur et vincientur in lacuet claudentur in carcere;et post multos dies visitabuntur.
ISA|24|23|Et erubescet luna, et confundetur sol,quia regnavit Dominus exercituum in monte Sion et in Ierusalemet in conspectu senum suorum glorificabitur.
ISA|25|1|Domine, Deus meus es tu;exaltabo te, confitebor no mini tuo,quoniam fecisti mirabilia,cogitationes antiquas, fideles, veraces.
ISA|25|2|Quia posuisti civitatem in tumulum,urbem munitam in ruinam:arx superborum non amplius est civitas,in sempiternum non reaedificabitur.
ISA|25|3|Super hoc glorificabit te populus fortis,civitas gentium robustarum timebit te;
ISA|25|4|quia factus es fortitudo pauperi,fortitudo egeno in tribulatione sua,protectio a turbine,umbraculum ab aestu:spiritus enim robustorumquasi imber hiemalis.
ISA|25|5|Sicut aestus in aridatumultum superborum humiliabis; sicut aestus in umbra nubiscanticum fortium reprimes.
ISA|25|6|Et faciet Dominus exercituumomnibus populis in monte hocconvivium pinguium,convivium vini meri,pinguium medullatorum,vini deliquati.
ISA|25|7|Et praecipitabit in monte istofaciem vinculi colligati super omnes populoset telam, quam orditus est super omnes nationes.
ISA|25|8|Praecipitabit mortem in sempiternumet absterget Dominus Deus lacrimam ab omni facieet opprobrium populi sui auferet de universa terra,quia Dominus locutus est.
ISA|25|9|Et dicetur in die illa: " Ecce Deus noster iste,exspectavimus eum, ut salvaret nos;iste Dominus, sustinuimus eum:exsultabimus et laetabimur in salutari eius.
ISA|25|10|Quia requiescet manus Domini in monte isto ".Et triturabitur Moab in loco suo,sicuti teruntur paleae in sterquilinio;
ISA|25|11|et extendet manus suas in medio eius,sicut extendit natans ad natandum;et humiliabitur superbia eiuscum allisione manuum eius.
ISA|25|12|Et firmum munimentum murorum tuorum evertit,deiecit, prostravit in terram usque ad pulverem.
ISA|26|1|In die illa cantabitur canticum istud in terra Iudae: Urbs fortis nobis in salutem;posuit muros et antemurale.
ISA|26|2|Aperite portas, et ingrediatur gens iusta,quae servat fidem.
ISA|26|3|Propositum eius est firmum;servabis pacem,quia in te speravit.
ISA|26|4|Sperate in Dominum in saeculis aeternis,Dominus est petra aeterna.
ISA|26|5|Quia evertit habitantes in excelso,civitatem sublimem humiliabit;humiliabit eam usque ad terram,detrahet eam usque ad pulverem.
ISA|26|6|Conculcabit eam pes, pedes pauperis,gressus egenorum.
ISA|26|7|Semita iusti recta est;rectum callem iusti complanas.
ISA|26|8|Et in semita iudiciorum tuorum, Domine, speravimus in te;ad nomen tuum et ad memoriale tuum desiderium animae.
ISA|26|9|Anima mea desiderat te in nocte,sed et spiritu meo in praecordiis meis te quaero.Cum resplenduerint iudicia tua in terra,iustitiam discent habitatores orbis.
ISA|26|10|Fit misericordia impio,non discet iustitiam;in terra probitatis inique geritet non videt maiestatem Domini.
ISA|26|11|Domine, exaltata est manus tua, et non vident;videant confusi zelum tuum in populum,et ignis hostium tuorum devorabit eos.
ISA|26|12|Domine, dabis pacem nobis;omnia enim opera nostra operatus es nobis.
ISA|26|13|Domine Deus noster, possederunt nos domini absque te;tantum in te recordemur nominis tui.
ISA|26|14|Mortui non reviviscent,defuncti non resurgent;propterea visitasti et contrivisti eos et perdidisti omnem memoriam eorum.
ISA|26|15|Auxisti gentem, Domine,auxisti gentem, glorificatus es;elongasti omnes terminos terrae.
ISA|26|16|Domine, in angustia quaesierunt te,fuderunt incantationem, castigatio tua in eis.
ISA|26|17|Sicut quae concipit, cum appropinquaverit ad partumdolens clamat in doloribus suis,sic facti sumus a facie tua, Domine.
ISA|26|18|Concepimus et parturivimus,quasi peperimus ventum.Salutes non fecimus in terra,ideo non nati sunt habitatores terrae.
ISA|26|19|Reviviscent mortui tui, interfecti mei resurgent.Expergiscimini et laudate, qui habitatis in pulvere,quia ros lucis ros tuus,et terra defunctos suos edet in lucem.
ISA|26|20|Vade, populus meus, intra in cubicula tua,claude ostia tua super te,abscondere modicum ad momentum,donec pertranseat indignatio.
ISA|26|21|Ecce enim Dominus egredietur de loco suo,ut visitet iniquitatem habitatoris terrae contra eum;et revelabit terra sanguinem suumet non operiet ultra interfectos suos ".
ISA|27|1|In die illa visitabit Dominusin gladio suo duro et forti et grandisuper Leviathan serpentem fugacemet super Leviathan serpentem tortuosumet occidet draconem, qui in mari est.
ISA|27|2|In die illa vinea erit iucunda;cantate ei.
ISA|27|3|Ego Dominus, qui servo eam;per singula momenta irrigabo eam.Ne forte visitetur contra eam,nocte et die servo eam.
ISA|27|4|Indignatio non est mihi.Quis dabit mihi spinam et veprem?In proelio gradiar super eam,succendam eam pariter,
ISA|27|5|nisi forte protectionem meam apprehendat,faciat pacem mecum,pacem faciat mecum.
ISA|27|6|Diebus futuris radices mittet Iacob,florebit et germinabit Israel,et implebunt faciem orbis fructibus.
ISA|27|7|Numquid iuxta plagam percutientis eum percussit eum?Aut, sicut occiduntur occisi eius, occisus est?
ISA|27|8|In mensura punit eum deiciens eum,impellit in spiritu suo duro, tempore quo spirat eurus.
ISA|27|9|Idcirco super hoc dimittetur iniquitas Iacob,et hic erit omnis fructus ablationis peccati eius:ut scilicet ponat omnes lapides altarissicut lapides calcis comminutos,ne exstent luci et thymiateria.
ISA|27|10|Civitas enim munita desolata est,habitaculum derelictum et dimissum quasi desertum;ibi pascetur vitulus et ibi accubabitet consumet arbusta eius.
ISA|27|11|In siccitate frondes illius conterentur;mulieres venient et comburent eas.Ipse enim non est populus sapiens,propterea non miserebitur eius, qui fecit eum,et, qui formavit eum, non parcet ei.
ISA|27|12|Et erit: in die illa percutiet spicas Dominusa Flumine usque ad torrentem Aegypti;et vos congregabiminiunus et unus, filii Israel.
ISA|27|13|Et erit: in die illa clangetur in tuba magna;et venient, qui perditi fuerant de terra Assyriorum,et qui eiecti erant in terra Aegypti,et adorabunt Dominumin monte sancto in Ierusalem.
ISA|28|1|Vae coronae superbiae ebriorum Ephraimet flori decidenti gloriae maiestatis eius,qui erant in vertice vallis pinguissimae,errantes a vino!
ISA|28|2|Ecce validus et fortis Dominosicut impetus grandinis, turbo confringens,sicut impetus aquarum multarum inundantium,et deiciet in terram violenter.
ISA|28|3|Pedibus conculcabiturcorona superbiae ebriorum Ephraim;
ISA|28|4|et erit flos decidens gloriae maiestatis eius,qui est super verticem vallis pinguium,quasi ficus praecox ante messem,quam quis, ut viderit,manu statim arreptam devorabit.
ISA|28|5|In die illa erit Dominus exercituumcorona gloriaeet sertum maiestatisresiduo populi sui
ISA|28|6|et spiritus iudiciisedenti ad iudicandumet fortitudovertentibus proelium usque ad portam.
ISA|28|7|Verum hi quoque prae vino vacillantet prae ebrietate nutant;sacerdos et propheta vacillant prae ebrietate,absorpti sunt a vino,nutant in ebrietate,vacillant in visione,fluctuant in iudicio.
ISA|28|8|Omnes enim mensae repletae sunt vomitu sordiumque,ita ut non esset ultra locus.
ISA|28|9|Quem docebit scientiam?Et quem intellegere faciet auditum?Ablactatos a lacte,avulsos ab uberibus.
ISA|28|10|Etenim praeceptum ad praeceptum, praeceptum ad praeceptum,regula ad regulam, regula ad regulam,modicum ibi, modicum ibi.
ISA|28|11|Balbis enim labiis et lingua alteraloquetur ad populum istum,
ISA|28|12|cui dixerat: " Haec requies, reficite lassum;et hoc est refrigerium ".Et noluerunt audire.
ISA|28|13|Et erit eis verbum Domini: Praeceptum ad praeceptum, praeceptum ad praeceptum,regula ad regulam, regula ad regulam,modicum ibi, modicum ibi ",ut vadant et cadant retrorsum et conteranturet illaqueentur et capiantur.
ISA|28|14|Propter hoc audite verbum Domini,viri illusores, qui dominamini super populum meum,qui est in Ierusalem.
ISA|28|15|Dixistis enim: " Percussimus foedus cum morteet cum inferno fecimus pactum;flagellum inundans cum transierit,non veniet super nos,quia posuimus mendacium spem nostramet in fallacia absconditi sumus ".
ISA|28|16|Idcirco haec dicit Dominus Deus: Ecce ego fundamentum ponam in Sion, lapidem,lapidem probatum, angularem, pretiosum, fundatum;qui crediderit, non turbabitur.
ISA|28|17|Et ponam iudicium tamquam normamet iustitiam tamquam perpendiculum;et subvertet grando spem mendacii,et latibulum aquae inundabunt.
ISA|28|18|Et delebitur foedus vestrum cum morte,et pactum vestrum cum inferno non stabit;flagellum inundans cum transierit,eritis ei in conculcationem.
ISA|28|19|Quandocumque pertransierit, tollet vos;quoniam mane diluculo pertransibit,in die et in nocte,et erit tantummodo horrendum intellegere auditum ".
ISA|28|20|Coangustatum est enim stratum, ut quis se extendat,et pallium brevius, ut quis se operire possit.
ISA|28|21|Sicut enim in monte Pharasim stabit Dominus,sicut in valle, quae est in Gabaon, irascetur,ut faciat opus suum, novum opus suum,ut operetur operationem suam,peregrinam operationem suam.
ISA|28|22|Et nunc nolite illudere,ne forte constringantur vincula vestra;decretum enim destructionis audivia Domino, Deo exercituum,super universam terram.
ISA|28|23|Auribus percipite et audite vocem meam,attendite et audite eloquium meum.
ISA|28|24|Numquid tota die arat arans, ut serat,proscindit et sarrit humum suam?
ISA|28|25|Nonne, cum adaequaverit faciem eius,spargit nigellam et serit cuminum,ponit triticum et hordeumet far in finibus suis?
ISA|28|26|Erudit enim illum recte,Deus suus docet illum.
ISA|28|27|Non enim in serris trituratur nigella,nec rota plaustri super cuminum circuit;sed in virga excutitur nigella,et cuminum in baculo.
ISA|28|28|Numquid comminuitur triticum?Verum non in perpetuum triturans triturabit illum,neque vexabit eum rota plaustri,nec ungulis suis comminuet eum.
ISA|28|29|Et hoc a Domino, Deo exercituum, exivit;mirabile fecit consilium,magnificavit sapientiam.
ISA|29|1|Vae Ariel, Ariel, civitas,quam circumdedit David!Addite annum ad annum,sollemnitates evolvantur;
ISA|29|2|et circumvallabo Ariel,et erit maeror et maestitia,et erit mihi quasi Ariel.
ISA|29|3|Et circumdabo te quasi sphaeramet iaciam contra te aggeremet munimenta ponam in obsidionem tuam.
ISA|29|4|Humiliaberis, de terra loqueris,et de pulvere vix audietur eloquium tuum,et erit quasi pythonis de terra vox tua,et de humo eloquium tuum mussitabit.
ISA|29|5|Et erit sicut pulvis tenuis multitudo superborum tuorum,et sicut palea volans multitudo fortium.Eritque repente confestim,
ISA|29|6|a Domino exercituum visitaberisin tonitruo et commotione terrae,magno fragore, turbine et tempestateet flamma ignis devorantis.
ISA|29|7|Et erit sicut somnium visionis nocturnaemultitudo omnium gentium, quae dimicant contra Ariel,et omnes, qui pugnant contra eam et contra munimenta eius et oppressores eius;
ISA|29|8|Et sicut somniat esuriens, et ecce comedit,cum autem fuerit expergefactus, vacua est anima eius;et sicut somniat sitiens, et ecce bibitet, postquam fuerit expergefactus, lassus adhuc sitit,et anima eius vacua est,sic erit multitudo omnium gentiumdimicantium contra montem Sion.
ISA|29|9|Obstupescite et admiramini,excaecamini et caeci estote,inebriamini et non a vino,vacillate et non ab ebrietate.
ISA|29|10|Quoniam miscuit vobis Dominus spiritum soporis,clausit oculos vestroset capita vestra operuit.
ISA|29|11|Et erit vobis visio omnis sicut verba libri signati; quem cum dederint scienti litteras dicentes: " Lege istum ", respondebit: " Non possum, signatus est enim ".
ISA|29|12|Et dabitur liber nescienti litteras diceturque ei: " Lege ", et respondebit: " Nescio litteras ".
ISA|29|13|Et dixit Dominus: Eo quod appropinquat populus iste ore suoet labiis suis glorificat me,cor autem eius longe est a me,et est timor eorum erga mevelut mandatum hominum perceptum,
ISA|29|14|ideo ecce ego addam ut admirationem faciampopulo huic miraculo grandi et stupendo:peribit sapientia sapientium eius,et prudentia prudentium eius abscondetur ".
ISA|29|15|Vae, qui profunde a Dominoconsilium abscondunt,quorum sunt in tenebris opera, et dicunt: Quis videt nos, et quis novit nos? ".
ISA|29|16|Perversa cogitatio vestra!Numquid quasi lutum reputabitur figulus,ut dicat opus factori suo: Non fecisti me ";et figmentum dicat fictori suo: Non intellegis "?
ISA|29|17|Nonne adhuc in modico et in brevi convertetur Libanus in hortum,et hortus in saltum reputabitur?
ISA|29|18|Et audient in die illa surdi verba libri,et de tenebris et caligine oculi caecorum videbunt.
ISA|29|19|Et addent mites in Domino laetitiam,et pauperrimi hominum in Sancto Israel exsultabunt;
ISA|29|20|quoniam defecit, qui praevalebat,consummatus est illusor,et succisi sunt omnes, qui vigilabant super iniquitatem,
ISA|29|21|qui peccare faciebant homines in verboet arguentem in porta supplantabantet deiecerunt inanibus verbis iustum.
ISA|29|22|Propter hoc haec dicit Dominusad domum Iacob, qui redemit Abraham: Non modo confundetur Iacob,nec modo vultus eius erubescet;
ISA|29|23|sed, cum viderit opera manuum mearum,in medio sui sanctificabunt nomen meumet sanctificabunt Sanctum Iacobet Deum Israel pavebunt,
ISA|29|24|et scient errantes spiritu sapientiam,et mussitatores discent doctrinam ".
ISA|30|1|" Vae, filii desertores, dicit Dominus,eo quod facitis consilium et non ex me,et pactum statuitis et non per spiritum meum,ut addatis peccatum super peccatum!
ISA|30|2|Qui ambulatis, ut descendatis in Aegyptum,et os meum non interrogastis,sperantes auxilium in fortitudine pharaoniset habentes fiduciam in umbra Aegypti.
ISA|30|3|Et erit vobis fortitudo pharaonis in confusionem,et fiducia sub umbra Aegypti in ignominiam.
ISA|30|4|Cum fuerint enim in Tani principes tui,et nuntii tui usque ad Hanes pervenerint,
ISA|30|5|omnes confundentursuper populo, qui eis prodesse non potest;non erit in auxilium et in utilitatem sed in confusionem et opprobrium ".
ISA|30|6|Oraculum iumentorum Nageb.In terra tribulationis et angustiae,leaenae et leonis rugientis,viperae et draconis volantisportant super umeros iumentorum divitias suaset super gibbum camelorum thesauros suosad populum, qui eis prodesse non poterit.
ISA|30|7|Aegyptus enim frustra et vane auxiliabitur;ideo vocavi Rahab otiosam.
ISA|30|8|Nunc ingredere, scribe coram eis super buxumet in libro diligenter exara illud,et erit in posterumin testimonium usque in aeternum.
ISA|30|9|Populus enim rebellis est,et filii mendaces,filii nolentes audire legem Domini;
ISA|30|10|qui dicunt videntibus: " Nolite videre "et aspicientibus: " Nolite aspicere nobis ea, quae recta sunt;loquimini nobis placentia, aspicite nobis illusiones.
ISA|30|11|Recedite a via, declinate a semita,tollite a facie nostra Sanctum Israel ".
ISA|30|12|Propterea haec dicit Sanctus Israel: Pro eo quod reprobastis verbum hocet sperastis in perversitatem et in perfidiamet innixi estis super eis,
ISA|30|13|propterea erit vobis iniquitas haecsicut interruptio cadens, locus tumens in muro excelso,cuius confractio subito, dum non speratur,venit improviso;
ISA|30|14|et comminuetur, sicut conteritur lagoena figuli,contritione absque misericordia,et non invenietur de fragmentis eius testa,in qua capiatur igniculus de incendio,aut hauriatur aqua de fovea ".
ISA|30|15|Quia haec dixit Dominus Deus, Sanctus Israel: In conversione et quiete salvi eritis;in silentio et in spe erit fortitudo vestra ".Et noluistis
ISA|30|16|et dixistis: Nequaquam, sed super equis fugiemus ",ideo fugietis;et: " Super veloces ascendemus ",ideo veloces erunt, qui persequentur vos.
ISA|30|17|Mille pavebunt a facie terroris unius,et a facie terroris quinque fugietis,donec relinquaminiquasi malus in vertice montiset quasi signum super collem.
ISA|30|18|Propterea exspectat Dominus, ut misereatur vestri,et ideo exaltabitur parcens vobis,quia Deus iudicii Dominus;beati omnes, qui exspectant eum.
ISA|30|19|Nam, popule Sion, qui habitas in Ierusalem,plorans nequaquam plorabis:miserans miserebitur tui ad vocem clamoris tui;statim ut audierit, respondebit tibi.
ISA|30|20|Et dabit vobis Dominuspanem angustiae et aquam afflictionis,sed non amplius avolabit a te doctor tuus;et erunt oculi tui videntes praeceptorem tuum,
ISA|30|21|et aures tuae audient verbum post tergum monentis: Haec via, ambulate in ea ",si declinaveritis ad dexteram vel ad sinistram.
ISA|30|22|Et contaminabis laminas sculptilium argentorum tuorumet vestimentum conflatilis aurei tui;disperges ea sicut immunditiam menstruatae. Egredere " dices ei.
ISA|30|23|Et dabit pluviam semini tuo,quod seminaveris in terra,et panis frugum terrae erit uberrimus et pinguis;pascetur pecus tuum in die illo, agnus in pascuis spatiosis,
ISA|30|24|et boves tui et asini, qui operantur terram,commixtum migma comedentventilatum in pala et ventilabro.
ISA|30|25|Et erunt super omnem montem excelsumet super omnem collem elevatumrivi currentium aquarumin die interfectionis multorum,cum ceciderint turres.
ISA|30|26|Et erit lux lunae sicut lux solis,et lux solis erit septempliciter sicut lux septem dierumin die, qua alligaverit Dominus vulnus populi suiet percussuram plagae eius sanaverit.
ISA|30|27|Ecce nomen Domini venit de longinquo,ardens furor eius, et gravis eius fragor;labia eius repleta sunt indignatione,et lingua eius quasi ignis devorans.
ISA|30|28|Spiritus eius velut torrens inundans,usque ad collum pertingens,ad cribrandas gentes in cribro funesto,et frenum dolosum in maxillis populorum.
ISA|30|29|Canticum erit vobissicut nox sanctificatae sollemnitatis,et laetitia cordissicut eius, qui ad sonum tibiae pergitin montem Domini,ad petram Israel.
ISA|30|30|Et auditam faciet Dominusgloriam vocis suaeet terrorem brachii suiostendet in comminatione furoriset flamma ignis devorantis,in turbine et in imbre et in lapide grandinis.
ISA|30|31|A voce enim Domini pavebitAssyrius virga percussus.
ISA|30|32|Et erit omnis ictus baculi percutientis,quem requiescere faciet Dominussuper eum in tympanis et citharis,et in bellis agitatis expugnabit eos.
ISA|30|33|Praeparata est enim ab heri Topheth,praeparata, profunda et dilatata,in pyra eius ignis et ligna multa;flatus Domini sicut torrens sulphurissuccendit eam.
ISA|31|1|Vae, qui descendunt in Aegyptum ad auxilium,in equis speranteset habentes fiduciam super quadrigis, quia multae sunt,et super equitibus, quia praevalidi nimis,et non intendunt in Sanctum Israelet Dominum non requirunt!
ISA|31|2|Tamen et ipse sapiens adducit malumet verba sua non retractat;et consurget contra domum pessimorumet contra auxilium operantium iniquitatem.
ISA|31|3|Aegyptius homo et non Deus,et equi eorum caro et non spiritus;et Dominus inclinabit manum suam,et corruet auxiliator,et cadet, cui praestatur auxilium,simulque omnes consumentur.
ISA|31|4|Quia haec dicit Dominus ad me: Quomodo si rugit leo et catulus leonis super praedam suam,cum occurrerit ei multitudo pastorum,a voce eorum non formidabit et a multitudine eorum non pavebit,sic descendet Dominus exercituum, ut proelietur super montem Sion et super collem eius.
ISA|31|5|Sicut aves volantes,sic proteget Dominus exercituum Ierusalem,protegens et liberans,parcens et salvans ".
ISA|31|6|Convertimini ad eum, a quo penitus recesseratis,filii Israel.
ISA|31|7|In die enim illa abiciet viridola argentea sua et idola aurea sua,quae fecerunt vobis manus vestrae in peccatum;
ISA|31|8|et cadet Assyria in gladio non viri,et gladius non hominis vorabit eum,et fugiet a facie gladii,et iuvenes eius vectigales erunt.
ISA|31|9|Et fortitudo eius prae terrore transibit,et pavebunt signum principes eius,dixit Dominus, cuius ignis est in Sion,et caminus eius in Ierusalem.
ISA|32|1|Ecce in iustitia regnabit rex,et principes in iudicio praee runt.
ISA|32|2|Et erit vir sicut latibulum a ventoet refugium a tempestate,sicut rivi aquarum in sitiente terraet umbra petrae magnae in terra arida.
ISA|32|3|Non caligabunt oculi videntium,et aures audientium diligenter auscultabunt,
ISA|32|4|et cor stultorum intelleget scientiam,et lingua balborum velociter loquetur et plane.
ISA|32|5|Non vocabitur ultra is, qui insipiens est, nobilis,neque fraudulentus appellabitur maior;
ISA|32|6|stultus enim fatua loquitur,et cor eius cogitat iniquitatem,ut perficiat impietatemet loquatur contra Dominum erroreset vacuam faciat animam esurientemet potum sitienti auferat.
ISA|32|7|Fraudulenti fraudes pessimae sunt;ipse enim cogitationes concinnatad perdendos mites in sermone mendaci,etiam quando pauper iudicium vindicat.
ISA|32|8|Nobilis vero consilia nobilia datet ipse ad nobilia assurget.
ISA|32|9|Mulieres vanae, surgite, audite vocem meam;filiae confidentes, percipite auribus eloquium meum.
ISA|32|10|Post dies enim et annumvos pavebitis confidentes;consummata est enim vindemia,collectio ultra non veniet.
ISA|32|11|Obstupescite, vanae;pavete, confidentes,exuite vos et nudate vos,accingite lumbos vestros.
ISA|32|12|Super ubera plangite,super regione desiderabili,super vinea fertili.
ISA|32|13|Super humum populi meispinae et vepres ascendent,super omnes domos gaudii,super civitatem exsultantem.
ISA|32|14|Domus enim dimissa est;multitudo urbis relicta est,Ophel et Bahan erunt speluncaeusque in aeternum,gaudium onagrorum,pascua gregum,
ISA|32|15|donec effundatur super nosspiritus de excelso.Et erit desertum in hortum,et hortus in saltum reputabitur,
ISA|32|16|et habitabit in solitudine iudicium,et iustitia in horto sedebit;
ISA|32|17|et erit opus iustitiae pax,et cultus iustitiae silentium,et securitas usque in sempiternum.
ISA|32|18|Et sedebit populus meus in habitatione paciset in tabernaculis fiduciaeet in locis securis.
ISA|32|19|Et penitus cadet saltus,et profunde deprimetur civitas.
ISA|32|20|Beati, qui seminatis super omnes aquas,immittentes pedem bovis et asini.
ISA|33|1|Vae, qui praedaris, cum nemo te praedatus sit;qui devastas, cum nemo te devastaverit!Cum consummaveris depraedationem, depraedaberis;cum perfeceris devastationem, te devastabunt.
ISA|33|2|Domine, miserere nostri,te enim exspectavimus;esto brachium nostrum in maneet salus nostra in tempore tribulationis.
ISA|33|3|A voce fragoris fugerunt populi,ab exaltatione tua dispersae sunt gentes.
ISA|33|4|Et congregabuntur spolia, sicut colligitur bruchus;sicut discurrunt locustae, ad ea discurritur.
ISA|33|5|Sublimis est Dominus, quoniam habitat in excelso;implet Sion iudicio et iustitia.
ISA|33|6|Et erit firmitas in temporibus tuis;divitiae salutis sapientia et scientia:timor Domini ipse est thesaurus eius.
ISA|33|7|Ecce praecones clamabunt foris,angeli pacis amare flebunt.
ISA|33|8|Dissipatae sunt viae, cessavit transiens per semitam;irritum fecit pactum,reiecit testes,non reputavit homines.
ISA|33|9|Luget et elanguescit terra,confusus est Libanus et obsorduit,et factus est Saron sicut desertum,et exaruerunt Basan et Carmelus.
ISA|33|10|" Nunc consurgam, dicit Dominus,nunc exaltabor, nunc sublevabor.
ISA|33|11|Concipietis fenum, parietis stipulam;spiritus meus ut ignis vorabit vos.
ISA|33|12|Et erunt populi fornaces calcis:spinae congregatae igne comburentur.
ISA|33|13|Audite, qui longe estis, quae fecerim,et cognoscite, vicini, fortitudinem meam ".
ISA|33|14|Conterriti sunt in Sion peccatores,possedit tremor impios.Quis poterit habitare de vobis cum igne devorante?Quis habitabit ex vobis cum ardoribus sempiternis?
ISA|33|15|Qui ambulat in iustitiis et loquitur aequitates,qui reicit lucra ex rapiniset excutit manus suas, ne munera accipiat,qui obturat aures suas, ne audiat sanguinem,et claudit oculos suos, ne videat malum:
ISA|33|16|iste in excelsis habitabit,munimenta saxorum refugium eius;panis ei datus est, aquae eius fideles sunt.
ISA|33|17|Regem in decore suo videbunt oculi tui,cernent terram longinquam.
ISA|33|18|Cor tuum cum timore inquiret: Ubi est scriba? Ubi ponderator?Ubi computator turrium? ".
ISA|33|19|Populum impudentem non videbis,populum profundi sermonis, ininterpretabilis,linguae barbarae absque intellegentia.
ISA|33|20|Respice Sion civitatem sollemnitatum nostrarum!Oculi tui videbunt Ierusalem,habitationem securam,tabernaculum quod nequaquam transferri poterit;nec auferentur clavi eius in sempiternum,et omnes funiculi eius non rumpentur.
ISA|33|21|Quia ibi potens Dominus pro nobisloco fluviorum, rivorum late patentium;non transibit ibi navis remigum,neque navis magna transgredietur eum.
ISA|33|22|Dominus enim iudex noster, Dominus legifer noster,Dominus rex noster: ipse salvabit nos.
ISA|33|23|Laxati sunt funiculi tuinec sustinent malum suum,ut dilatare velum non queant.Tunc divident caeci praedam multam;claudi diripient rapinam.
ISA|33|24|Nec dicet incola: " Elangui ".Populus, qui habitat in ea,auferetur ab eo iniquitas.
ISA|34|1|Accedite, gentes, ad audien dum;et populi, attendite.Audiat terra et plenitudo eius,orbis et omne germen eius.
ISA|34|2|Quia indignatio Domini super omnes gentes,et furor super universam militiam eorum:ad interitum devovit eos et dedit eos in occisionem.
ISA|34|3|Interfecti eorum proicientur,et de cadaveribus eorum ascendet foetor;dissolventur montes sanguine eorum.
ISA|34|4|Et tabescet omnis militia caelorum,et complicabuntur sicut liber caeli, et omnis militia eorum defluet,sicut defluit folium de vinea et arida frons de ficu.
ISA|34|5|Quoniam inebriatus est in caelo gladius meus:ecce super Edom descendetet super populum interfectionis meae ad iudicium.
ISA|34|6|Gladius Domini repletus est sanguine,incrassatus est adipe,de sanguine agnorum et hircorum, de adipe viscerum arietum;victima enim Domini in Bosra,et interfectio magna in terra Edom.
ISA|34|7|Cadunt bubali cum eis,iuvenci cum tauris;inebriabitur terra eorum sanguine,et humus eorum adipe pinguium,
ISA|34|8|quia dies ultionis Domini,annus retributionum ad vindicandam Sion.
ISA|34|9|Et convertentur torrentes eius in picem,et humus eius in sulphur,et erit terra eius in picem ardentem.
ISA|34|10|Nocte et die non exstinguetur,in sempiternum ascendet fumus eius,a generatione in generationem desolabitur,in saecula saeculorum non erit transiens per eam.
ISA|34|11|Et possidebunt illam onocrotalus et ericius,noctua et corvus habitabunt in ea;et extendet super eam mensuram solitudiniset perpendiculum desolationis.
ISA|34|12|Nobiles eius non erunt,nec regnum proclamabunt;et omnes principes eius erunt in nihilum.
ISA|34|13|Et orientur in domibus eius spinae,urticae et paliurus in munitionibus eius;et erit cubile draconumet pascua struthionum.
ISA|34|14|Et occurrent hyaenae thoibus,et pilosus clamat ad amicum suum;ibi cubat lamiaet invenit sibi requiem.
ISA|34|15|Ibi nidificat serpens ovaque deponitet circumfodit et fovet in umbra eius;illuc congregantur milvi alter ad alterum.
ISA|34|16|Requirite in libro Domini et legite:unum ex eis non deest,alter alterum exspectare non debet;quia os Domini praecepit,et spiritus eius ipse congregavit ea.
ISA|34|17|Et ipse misit eis sortem,et manus eius divisit terram illis in mensura;usque in aeternum possidebunt eam,in generatione et generatione habitabunt in ea.
ISA|35|1|Laetentur deserta et invia,et exsultet solitudo et floreat quasi lilium.
ISA|35|2|Germinet et exsultetlaetabunda et laudans.Gloria Libani data est ei,decor Carmeli et Saron;ipsi videbunt gloriam Domini,maiestatem Dei nostri.
ISA|35|3|Confortate manus dissolutaset genua debilia roborate.
ISA|35|4|Dicite pusillanimis: Confortamini, nolite timere!Ecce Deus vester,ultio veniet, retributio Dei;ipse veniet et salvabit vos ".
ISA|35|5|Tunc aperientur oculi caecorum,et aures surdorum patebunt.
ISA|35|6|Tunc saliet sicut cervus claudus,et exsultabit lingua mutorum,quia erumpent in deserto aquae,et torrentes in solitudine.
ISA|35|7|Et terra arida erit in stagnum,et sitiens in fontes aquarum;in cubilibus, in quibus dracones habitabant,erit locus calami et iunci.
ISA|35|8|Et erit ibi semita et via;et via sancta vocabitur:non transibit per eam pollutus;et erit eis directa via,ita ut stulti non errent per eam.
ISA|35|9|Non erit ibi leo,et rapax bestia non ascendet per eamnec invenietur ibi;et ambulabunt, qui liberati fuerint,
ISA|35|10|et redempti a Domino revertentur.Et venient in Sion cum laude,et laetitia sempiterna super caput eorum:gaudium et laetitiam obtinebunt,et fugiet maeror et gemitus.
ISA|36|1|Et factum est in quarto deci mo anno regis Ezechiae, ascendit Sennacherib rex Assyriorum super omnes civitates Iudae munitas et cepit eas.
ISA|36|2|Et misit rex Assyriorum Rabsacen de Lachis in Ierusalem ad regem Ezechiam in manu gravi, et stetit in aquaeductu piscinae superioris in via agri fullonis.
ISA|36|3|Et egressus est ad eum Eliachim filius Helciae, qui erat super domum, et Sobna scriba et Ioah filius Asaph a commentariis.
ISA|36|4|Et dixit ad eos Rabsaces: " Dicite Ezechiae: Haec dicit rex magnus, rex Assyriorum: Quae est ista fiducia, qua confidis?
ISA|36|5|Dixisti: " Verbum labiorum est consilium et fortitudo ad bellum". Nunc super quem habes fiduciam, quia recessisti a me?
ISA|36|6|Ecce confidis super baculum arundineum confractum istum, super Aegyptum; cui si innixus fuerit homo, intrabit in manum eius et perforabit eam: sic pharao rex Aegypti omnibus, qui confidunt in eo.
ISA|36|7|Quod si responderis mihi: "In Domino Deo nostro confidimus"; nonne ipse est, cuius abstulit Ezechias excelsa et altaria et dixit Iudae et Ierusalem: "Coram altari isto adorabitis"?
ISA|36|8|Et nunc sponde domino meo regi Assyriorum, et dabo tibi duo milia equorum, si poteris ex te praebere ascensores eorum.
ISA|36|9|Et quomodo averteris faciem unius ex servis domini mei minoribus? Et tamen confidis in Aegypto, in quadriga et in equitibus;
ISA|36|10|et nunc, numquid sine Domino ascendi ad terram istam, ut disperderem eam? Dominus dixit ad me: "Ascende super terram istam et disperde eam" ".
ISA|36|11|Et dixit Eliachim et Sobna et Ioah ad Rabsacen: "Loquere ad servos tuos Aramaice; intellegimus enim. Ne loquaris ad nos Iudaice in auribus populi, qui est super murum ".
ISA|36|12|Et dixit Rabsaces: " Numquid ad dominum tuum et ad te misit me dominus meus, ut loquerer omnia verba ista? Et non potius ad viros, qui sedent in muro, ut comedant stercora sua et bibant urinam suam vobiscum? ".
ISA|36|13|Et stetit Rabsaces et clamavit voce magna Iudaice et dixit: " Audite verba regis magni, regis Assyriorum:
ISA|36|14|Haec dicit rex: Non seducat vos Ezechias, quia non poterit eruere vos.
ISA|36|15|Et non vobis tribuat fiduciam Ezechias super Domino dicens: "Eruens liberabit nos Dominus; non dabitur civitas ista in manu regis Assyriorum".
ISA|36|16|Nolite audire Ezechiam. Haec enim dicit rex Assyriorum: Facite mecum benedictionem et egredimini ad me; et comedite unusquisque vineam suam et unusquisque ficum suam, et bibite unusquisque aquam de cisterna sua,
ISA|36|17|donec veniam et tollam vos ad terram, quae est ut terra vestra, terram frumenti et vini, terram panis et vinearum.
ISA|36|18|Ne illudat vos Ezechias dicens: "Dominus liberabit nos". Numquid liberaverunt dii gentium unusquisque terram suam de manu regis Assyriorum?
ISA|36|19|Ubi sunt dii Emath et Arphad? Ubi sunt dii Sepharvaim? Numquid liberaverunt Samariam de manu mea?
ISA|36|20|Quinam ex omnibus diis terrarum istarum eruerunt terram suam de manu mea? Numquid eruet Dominus Ierusalem de manu mea? ".
ISA|36|21|Et siluerunt et non responderunt ei verbum; mandaverat enim rex dicens: Ne respondeatis ei ".
ISA|36|22|Et ingressus est Eliachim filius Helciae, qui erat super domum, et Sobna scriba et Ioah filius Asaph a commentariis ad Ezechiam scissis vestibus; et nuntiaverunt ei verba Rabsacis.
ISA|37|1|Et factum est cum audisset rex Ezechias, scidit vestimen ta sua et obvolutus est sacco et intravit in domum Domini;
ISA|37|2|et misit Eliachim, qui erat super domum, et Sobnam scribam et seniores de sacerdotibus opertos saccis ad Isaiam filium Amos prophetam,
ISA|37|3|et dixerunt ad eum: " Haec dicit Ezechias: Dies tribulationis et correptionis et contumeliae dies haec, quia venerunt filii usque ad partum, et virtus non est pariendi.
ISA|37|4|Forsitan audiet Dominus Deus tuus verba Rabsacis, quem misit rex Assyriorum, dominus suus, ad blasphemandum Deum viventem, et puniet sermones, quos audivit Dominus Deus tuus; leva ergo orationem pro reliquiis, quae repertae sunt ".
ISA|37|5|Et venerunt servi regis Ezechiae ad Isaiam;
ISA|37|6|et dixit ad eos Isaias: "Haec dicetis domino vestro: Haec dicit Dominus: Ne timeas a facie verborum, quae audisti, quibus blasphemaverunt pueri regis Assyriorum me.
ISA|37|7|Ecce ego dabo ei spiritum, et audiet nuntium et revertetur ad terram suam, et corruere eum faciam gladio in terra sua ".
ISA|37|8|Reversus est autem Rabsaces et invenit regem Assyriorum proeliantem adversus Lobnam; audierat enim quia profectus esset de Lachis.
ISA|37|9|Et audivit de Tharaca rege Aethiopiae dicentes: " Egressus est, ut pugnet contra te ".Quod cum audisset, misit nuntios ad Ezechiam dicens:
ISA|37|10|" Haec dicetis Ezechiae regi Iudae loquentes: Non te decipiat Deus tuus, in quo tu confidis, dicens: "Non dabitur Ierusalem in manu regis Assyriorum".
ISA|37|11|Ecce tu audisti omnia, quae fecerunt reges Assyriorum omnibus terris, quas ad interitum devoverunt, et tu poteris liberari?
ISA|37|12|Numquid eruerunt eos dii gentium, quos subverterunt patres mei, Gozan et Charran et Reseph et filios Eden, qui erant in Thelassar?
ISA|37|13|Ubi est rex Emath et rex Arphad et rex urbis Sepharvaim, Ana et Ava? ".
ISA|37|14|Et tulit Ezechias epistulam de manu nuntiorum et legit eam. Et ascendit in domum Domini et expandit eam Ezechias coram Domino.
ISA|37|15|Et oravit Ezechias ad Dominum dicens:
ISA|37|16|" Domine exercituum, Deus Israel, qui sedes super cherubim, tu es Deus solus omnium regnorum terrae, tu fecisti caelum et terram.
ISA|37|17|Inclina, Domine, aurem tuam et audi; aperi, Domine, oculos tuos et vide et audi omnia verba Sennacherib, quae misit ad blasphemandum Deum viventem.
ISA|37|18|Vere enim, Domine, dissipaverunt reges Assyriorum gentes et regiones earum
ISA|37|19|et dederunt deos earum igni: non enim erant dii, sed opera manuum hominum, lignum et lapis; et comminuerunt eos.
ISA|37|20|Et nunc, Domine Deus noster, salva nos de manu eius; et cognoscant omnia regna terrae quia tu, Domine, es solus Deus ".
ISA|37|21|Et misit Isaias filius Amos ad Ezechiam dicens: " Haec dicit Dominus, Deus Israel: Pro quibus rogasti me de Sennacherib rege Assyriorum,
ISA|37|22|hoc est verbum, quod locutus est Dominus super eum:Despexit te, subsannavit te virgo filia Sion;post te caput movit filia Ierusalem.
ISA|37|23|Cui exprobrasti et quem blasphemasti?Et super quem exaltasti vocemet levasti altitudinem oculorum tuorum?Contra Sanctum Israel!
ISA|37|24|In manu servorum tuorum exprobrasti Dominoet dixisti: "In multitudine quadrigarum mearumego ascendi altitudinem montium, iuga Libani;et succidi excelsa cedrorum eiuset electas abietes illiuset introivi altitudinem summitatis eius,silvam condensam.
ISA|37|25|Ego fodi et bibi aquam alienamet exsiccavi vestigio pedis meiomnes rivos Aegypti".
ISA|37|26|Numquid non audisti?A saeculo feci illud; a diebus antiquisego plasmavi illud et nunc adduxi,ut fiat in eradicationem,in lapides eversos civitates munitae.
ISA|37|27|Habitatores earum breviata manucontremuerunt et confusi sunt;facti sunt sicut fenum agriet gramen viride et herba tectorum, quae exaruit a facie austri.
ISA|37|28|Sessionem tuamet egressum tuum et introitum tuum cognoviet insaniam tuam contra me.
ISA|37|29|Cum fureris adversum me,et superbia tua ascenderit in aures meas,ponam circulum in naribus tuiset frenum in labiis tuiset reducam te in viam,per quam venisti.
ISA|37|30|Tibi autem hoc erit signum:Comedantur hoc anno, quae colligi poterunt,et in anno secundo, quae sponte nascuntur;in anno autem tertio seminate et metiteet plantate vineas et comedite fructum earum.
ISA|37|31|Et mittet id, quod salvatum fuerit de domo Iudae,quod reliquum est, radicem deorsumet faciet fructum sursum.
ISA|37|32|Quia de Ierusalem exibit residuum,et, quod salvum fuerit, de monte Sion.Zelus Domini exercituum faciet istud.
ISA|37|33|Propterea haec dicit Dominus de rege Assyriorum:Non introibit civitatem hancet non iaciet ibi sagittamet non opponet ei clipeumet non mittet contra eam aggerem.
ISA|37|34|In via, qua venit, per eam revertetur,et civitatem hanc non ingredietur, dicit Dominus.
ISA|37|35|Et protegam civitatem istam, ut salvem eampropter me et propter David servum meum ".
ISA|37|36|Egressus est autem angelus Domini et percussit in castris Assyriorum centum octoginta quinque milia; et surrexerunt mane, et ecce omnes illi cadavera mortuorum.
ISA|37|37|Et egressus est et abiit; et reversus est Sennacherib rex Assyriorum et habitavit in Nineve.
ISA|37|38|Et factum est, cum adoraret in templo Nesroch dei sui, Adramelech et Sarasar filii eius percusserunt eum gladio fugeruntque in terram Ararat. Et regnavit Asarhaddon filius eius pro eo.
ISA|38|1|In diebus illis aegrotavit Ezechias usque ad mortem. Et introivit ad eum Isaias filius Amos propheta et dixit ei: " Haec dicit Dominus: Dispone domui tuae, quia morieris tu et non vives".
ISA|38|2|Et convertit Ezechias faciem suam ad parietem et oravit ad Dominum
ISA|38|3|et dixit: " Obsecro, Domine; memento, quaeso, quomodo ambulaverim coram te in veritate et in corde perfecto et, quod bonum est in oculis tuis, fecerim ". Et flevit Ezechias fletu magno.
ISA|38|4|Et factum est verbum Domini ad Isaiam dicens:
ISA|38|5|" Vade et dic Ezechiae: "Haec dicit Dominus, Deus David patris tui: Audivi orationem tuam, vidi lacrimas tuas; ecce ego adiciam super dies tuos quindecim annos
ISA|38|6|et de manu regis Assyriorum eruam te et civitatem istam et protegam hanc civitatem".
ISA|38|7|Hoc autem tibi erit signum a Domino quia faciet Dominus verbum hoc, quod locutus est:
ISA|38|8|Ecce ego reverti faciam umbram graduum, per quos descenderat in horologio Achaz in sole retrorsum decem gradibus ". Et reversus est sol decem gradibus per gradus, quos descenderat.
ISA|38|9|Scriptura Ezechiae regis Iudae, cum aegrotasset et convaluisset de infirmitate sua:
ISA|38|10|" Ego dixi: In dimidio dierum meorumvadam ad portas inferi;quaesivi residuum annorum meorum.
ISA|38|11|Dixi: Non videbo Dominum Deum in terra viventium,non aspiciam hominem ultrainter habitatores orbis.
ISA|38|12|Habitaculum meum ablatum est et abductum longe a mequasi tabernaculum pastorum;convolvit sicut textor vitam meam;de stamine succidit me.De mane usque ad vesperam confecisti me.
ISA|38|13|Prostratus sum usque ad mane,quasi leo sic conterit omnia ossa mea;de mane usque ad vesperam confecisti me.
ISA|38|14|Sicut pullus hirundinis, sic mussitabo,meditabor ut columba;attenuati sunt oculi meisuspicientes in excelsum.Domine, vim patior,sponde pro me.
ISA|38|15|Quid dicam, aut quid respondebit mihi?Ipse fecit!Incedam per omnes annos meosin amaritudine animae meae.
ISA|38|16|Domine, in te sperat cor meum;vivat spiritus meus,sana me et vivifica me;
ISA|38|17|ecce in pacem versa est amaritudo mea.Tu autem eruisti animam meama fovea consumptionis,proiecisti enim post tergum tuumomnia peccata mea.
ISA|38|18|Quia non infernus confitebitur tibi,neque mors laudabit te;non exspectabunt, qui descendunt in lacum,veritatem tuam.
ISA|38|19|Vivens, vivens ipse confitebitur tibi,sicut et ego hodie;pater filiis notam faciet veritatem tuam.
ISA|38|20|Domine, salvum me fac,et ad sonum citharae cantabimuscunctis diebus vitae nostraein domo Domini ".
ISA|38|21|Et iussit Isaias, ut tollerent massam de ficis et cataplasmarent super vulnus, et sanaretur.
ISA|38|22|Et dixit Ezechias: " Quod erit signum quia ascendam in domum Domini?".
ISA|39|1|In tempore illo misit Merodachbaladan filius Baladan rex Babylonis litteras et munera ad Ezechiam; audierat enim quod aegrotasset et convaluisset.
ISA|39|2|Laetatus est autem super eis Ezechias et ostendit eis cellam thesauri sui et argentum et aurum et aromata et oleum optimum et omnes apothecas supellectilis suae et universa, quae inventa sunt in thesauris eius. Nihil fuit, quod non ostenderet eis Ezechias in domo sua et in omni potestate sua.
ISA|39|3|Introivit autem Isaias propheta ad Ezechiam regem et dixit ei: " Quid dixerunt viri isti et unde venerunt ad te? ". Et dixit Ezechias: " De terra longinqua venerunt ad me, de Babylone ".
ISA|39|4|Et dixit: "Quid viderunt in domo tua?". Et dixit Ezechias: " Omnia, quae in domo mea sunt, viderunt; non fuit res, quam non ostenderim eis in thesauris meis ".
ISA|39|5|Et dixit Isaias ad Ezechiam: " Audi verbum Domini exercituum:
ISA|39|6|Ecce dies venient, et auferentur omnia, quae in domo tua sunt, et quae thesaurizaverunt patres tui usque ad diem hanc, in Babylonem; non relinquetur quidquam, dicit Dominus.
ISA|39|7|Et de filiis tuis, qui exibunt de te, quos genueris, tollent, et erunt eunuchi in palatio regis Babylonis ".
ISA|39|8|Et dixit Ezechias ad Isaiam: " Bonum verbum Domini, quod locutus est ". Et dixit: " Dummodo fiat pax et securitas in diebus meis ".
ISA|40|1|Consolamini, consolamini populum meum,dicit Deus vester.
ISA|40|2|Loquimini ad cor Ierusalemet clamate ad eam,quoniam completa est militia eius,expiata est iniquitas illius;suscepit de manu Dominiduplicia pro omnibus peccatis suis.
ISA|40|3|Vox clamantis: In deserto parate viam Domini,rectas facite in solitudinesemitas Dei nostri.
ISA|40|4|Omnis vallis exaltetur,et omnis mons et collis humilietur;et fiant prava in directa,et aspera in plana:
ISA|40|5|et revelabitur gloria Domini,et videbit omnis caro pariterquod os Domini locutum est ".
ISA|40|6|Vox dicentis: " Clama! ".Et dixi: " Quid clamabo? ".Omnis caro fenum,et omnis gloria eius quasi flos agri;
ISA|40|7|exsiccatum est fenum, et cecidit flos,quia spiritus Domini sufflavit in eo. Vere fenum est populus.
ISA|40|8|Exsiccatum est fenum, et cecidit flos;verbum autem Dei nostri manet in aeternum.
ISA|40|9|Super montem excelsum ascende,tu, quae evangelizas Sion;exalta in fortitudine vocem tuam,quae evangelizas Ierusalem;exalta, noli timere;dic civitatibus Iudae: Ecce Deus vester,
ISA|40|10|ecce Dominus Deus in virtute venit,et brachium eius dominatur:ecce merces eius cum eo,et praemium illius coram illo.
ISA|40|11|Sicut pastor gregem suum pascit,in brachio suo congregat agnoset in sinu suo levat;fetas ipse portat ".
ISA|40|12|Quis mensus est pugillo aquaset caelos palmo disposuit,modio continuit pulverem terraeet libravit in pondere monteset colles in statera?
ISA|40|13|Quis direxit spiritum Domini?Aut quis consilium suumostendit illi?
ISA|40|14|Cum quo iniit consilium, et instruxit eumet docuit eum semitam iustitiaeet erudivit eum scientiamet viam prudentiae ostendit illi?
ISA|40|15|Ecce gentes quasi stilla situlaeet quasi momentum pulveris in statera reputantur;ecce insulae quasi pulvis exiguus.
ISA|40|16|Et Libanus non sufficiet ad succendendum,et animalia eius non sufficient ad holocaustum.
ISA|40|17|Omnes gentes, quasi non sint, coram eo;quasi nihilum et inane reputantur ab eo.
ISA|40|18|Cui ergo similem facitis Deum?Aut quam imaginem ponitis ei?
ISA|40|19|Sculptile conflat faber,et aurifex auro figurat illud,et laminis argenteis argentarius.
ISA|40|20|Nimis pauper, ut offerat lignum imputribile:exquirit sibi sapientem artificem,ut statuat simulacrum,quod non moveatur.
ISA|40|21|Numquid non scitis? Numquid non audistis?Numquid non annuntiatum est vobis ab initio?Numquid non intellexistis fundamenta terrae?
ISA|40|22|Qui sedet super gyrum terrae,et habitatores eius sunt quasi locustae;qui extendit sicut velum caeloset expandit eos sicut tabernaculum ad inhabitandum;
ISA|40|23|qui redigit in nihilum principes,iudices terrae velut inane facit.
ISA|40|24|Et quidem neque plantatus neque satusneque radicatus in terra truncus eorum;repente flavit in eos, et aruerunt,et turbo quasi stipulam aufert eos.
ISA|40|25|" Et cui assimilabitis me,quasi aequalis ei sim ego? ",dicit Sanctus.
ISA|40|26|Levate in excelsum oculos vestroset videte: Quis creavit haec?Qui educit in numero militiam eorumet omnes ex nomine vocat;prae multitudine fortitudinis et roboris virtutisque eiusneque unum deest.
ISA|40|27|Quare dicis, Iacob,et loqueris, Israel: Abscondita est via mea a Domino,et a Deo meo iudicium meum transit? ".
ISA|40|28|Numquid nescis? Aut non audisti?Deus sempiternus Dominus,qui creavit terminos terrae;non deficiet neque laborabit,nec est investigatio sapientiae eius.
ISA|40|29|Qui dat lasso virtutemet invalido robur multiplicat.
ISA|40|30|Deficient pueri et laborabunt,et iuvenes lapsu labentur;
ISA|40|31|qui autem sperant in Domino,mutabunt fortitudinem,assument pennas sicut aquilae,current et non laborabunt,ambulabunt et non deficient.
ISA|41|1|Taceant ante me insulae,et gentes renovent fortitudinem;accedant et tunc loquantur,simul ad iudicium propinquemus.
ISA|41|2|Quis suscitavit ab oriente eum,cuius gressum sequitur iustitia?Dabit in conspectu eius genteset subiciet ei reges,quos reddet quasi pulverem gladius eius,sicut stipulam vento raptam arcus eius.
ISA|41|3|Persequetur eos, transibit in pace;semita sub pedibus eius non apparebit.
ISA|41|4|Quis operatus est et fecit,vocans generationes ab exordio?Ego Dominus, primuset cum novissimis ego sum.
ISA|41|5|Viderunt insulae et timuerunt,extrema terrae obstupuerunt,appropinquaverunt et accesserunt.
ISA|41|6|Unusquisque proximo suo auxiliabituret fratri suo dicet: " Confortare ".
ISA|41|7|Confortabit faber aurificem,percutiens malleo eum, qui cudit,dicens de glutino: " Bonum est ";et roborat eum clavis,ut non moveatur.
ISA|41|8|Tu autem, Israel, serve meus,Iacob, quem elegi,semen Abraham amici mei,
ISA|41|9|quem apprehendi ab extremis terrae,et a longinquis eius vocavi teet dixi tibi: " Servus meus es tu;elegi te et non abieci te ".
ISA|41|10|Ne timeas, quia ego tecum sum;ne declines, quia ego Deus tuus:confortabo te et auxiliabor tibiet sustentabo te dextera iustitiae meae.
ISA|41|11|Ecce confundentur et erubescentomnes, qui irascuntur adversum te;erunt quasi non sintet peribunt viri, qui contradicunt tibi.
ISA|41|12|Quaeres eos et non inveniesviros, qui rixantur tecum;erunt quasi non sint et veluti nihilum,viri bellantes adversum te.
ISA|41|13|Quia ego Dominus Deus tuusapprehendens manum tuamdicensque tibi: " Ne timeas;ego auxiliabor tibi.
ISA|41|14|Noli timere, vermis Iacob,homines ex Israel.Ego auxiliabor tibi ", dicit Dominuset redemptor tuus, Sanctus Israel.
ISA|41|15|Ecce posui te quasi plaustrum triturans novum,habens rostra serrantia.Triturabis montes et comminueset colles quasi pulverem pones.
ISA|41|16|Ventilabis eos, et ventus tollet eos,et turbo disperget eos;et tu exsultabis in Domino,in Sancto Israel laetaberis.
ISA|41|17|Egeni et pauperes quaerunt aquas, et non sunt,lingua eorum siti aruit.Ego, Dominus, exaudiam eos,Deus Israel non derelinquam eos.
ISA|41|18|Aperiam in decalvatis collibus fluminaet in medio vallium fontes;ponam desertum in stagna aquarumet terram aridam in rivos aquarum.
ISA|41|19|Plantabo in deserto cedrum,acaciam et myrtum et lignum olivae;ponam in solitudine abietem,ulmum et cupressum simul,
ISA|41|20|ut videant et sciantet recogitent et intellegant pariterquia manus Domini fecit hoc,et Sanctus Israel creavit illud.
ISA|41|21|Proferte causam vestram, dicit Dominus;afferte, si quid firmum habetis, dixit Rex Iacob.
ISA|41|22|Accedant et nuntient nobis, quaecumque ventura sunt.Priora, quae fuerunt, nuntiate,ut ponamus cor nostrum et sciamus novissima eorum;et, quae ventura sunt, indicate nobis.
ISA|41|23|Annuntiate, quae ventura sunt in futurum,ut sciamus quia dii estis vos;bene quoque aut male facite,ut inspiciamus et videamus simul.
ISA|41|24|Ecce vos estis nihilum,et opus vestrum nihil valet;abominatio est, qui eligit vos.
ISA|41|25|Suscitavi ab aquilone,et venit ab ortu solis;vocavi eum nomine;et conculcabit potentes quasi lutumet velut plastes calcans humum.
ISA|41|26|Quis annuntiavit ab exordio, ut sciamus,et a principio, ut dicamus: " Iustum est "?Non est neque annuntians neque praedicensneque audiens sermones vestros.
ISA|41|27|Primus ad Sion: Ecce adsunt;et Ierusalem laeta nuntiantem do.
ISA|41|28|Et vidi, et nemo erat,ex istis nullus consiliator,ut, si eos interrogarem,responderent verbum.
ISA|41|29|Ecce omnes iniquitas,vana opera eorum;ventus et inanesimulacra eorum.
ISA|42|1|Ecce servus meus, suscipiam eum;electus meus, complacet sibi in illo anima mea;dedi spiritum meum super eum,iudicium gentibus proferet.
ISA|42|2|Non clamabit neque vociferabitur,nec audietur vox eius foris.
ISA|42|3|Calamum quassatum non conteretet linum fumigans non exstinguet;in veritatem proferet iudicium.
ISA|42|4|Non languebit nec frangetur,donec ponat in terra iudicium;et legem eius insulae exspectant.
ISA|42|5|Haec dicit Dominus Deus,creans caelos et extendens eos,firmans terram et quae germinant ex ea,dans flatum populo, qui est super eam,et spiritum calcantibus eam:
ISA|42|6|" Ego, Dominus, vocavi te in iustitiaet apprehendi manum tuam;et formavi te et dedi tein foedus populi, in lucem gentium,
ISA|42|7|ut aperires oculos caecorumet educeres de conclusione vinctum,de domo carceris sedentes in tenebris.
ISA|42|8|Ego Dominus: hoc est nomen meum;et gloriam meam alteri non daboet laudem meam sculptilibus.
ISA|42|9|Quae prima fuerunt, ecce venerunt;nova quoque ego annuntio:antequam oriantur, audita vobis faciam ".
ISA|42|10|Cantate Domino canticum novum,laus eius ab extremis terrae;qui descenditis in mare, et plenitudo eius,insulae et habitatores earum.
ISA|42|11|Exsultent desertum et civitates eius,vici, quos habitat Cedar.Iubilent habitatores Petrae,de vertice montium clament.
ISA|42|12|Ponant Domino gloriamet laudem eius in insulis nuntient.
ISA|42|13|Dominus sicut fortis egredietur,sicut vir proeliator suscitabit zelum;vociferabitur et conclamabit,super inimicos suos praevalebit.
ISA|42|14|" Tacui semper, silui, patiens fui;sicut parturiens ululabo,gemam et fremam simul.
ISA|42|15|Desertos faciam montes et colleset omne gramen eorum exsiccabo;et ponam flumina in insulaset stagna arefaciam.
ISA|42|16|Et ducam caecos in viam, quam nesciunt,et in semitis, quas ignoraverunt, ambulare eos faciam;ponam tenebras coram eis in lucemet prava in recta.Haec verba faciam eiset non dereliquam eos ".
ISA|42|17|Conversi sunt retrorsum;confundantur confusione, qui confidunt in sculptili,qui dicunt conflatili: Vos dii nostri ".
ISA|42|18|Surdi, audite;et caeci, intuemini ad videndum.
ISA|42|19|Quis caecus sicut servus meus,et surdus sicut nuntius, quem ego mittam?Quis caecus sicut qui restitutus est?Et quis caecus sicut servus Domini?
ISA|42|20|Multa vidisti, sed non servas;aures aperuisti, sed non audis.
ISA|42|21|Dominus voluit propter iustitiam suammagnificare legem et extollere.
ISA|42|22|Ipse autem populus direptus et vastatus;in foveis conclusi omnes,et in domibus carcerum absconditi sunt.Facti sunt in rapinam, nec est qui eruat;in direptionem, nec est qui dicat: " Redde! ".
ISA|42|23|Quis est in vobis, qui audiat hoc,attendat et auscultet futura?
ISA|42|24|Quis dedit in direptionem Iacobet Israel vastantibus?Nonne Dominus ipse, cui peccavimus?Et noluerunt in viis eius ambulareet non audierunt legem eius.
ISA|42|25|Et effudit super eum indignationem furoris suiet forte bellum.Et combussit eum in circuitu, et non cognovit;et succendit eum, et non intellexit.
ISA|43|1|Et nunc haec dicit Dominus,qui creavit te, Iacob, et formavit te, Israel: Noli timere, quia redemi teet vocavi te nomine tuo; meus es tu.
ISA|43|2|Cum transieris per aquas, tecum ero,et flumina non operient te;cum ambulaveris in igne, non combureris,et flamma non ardebit in te,
ISA|43|3|quia ego Dominus Deus tuus,Sanctus Israel, salvator tuus:dedi propitiationem tuam Aegyptum,Aethiopiam et Saba pro te.
ISA|43|4|Quoniam pretiosus factus es in oculis meiset gloriosus, ego diligo teet dabo homines pro teet populos pro anima tua.
ISA|43|5|Noli timere, quoniam ego tecum sum:ab oriente adducam semen tuumet ab occidente congregabo te.
ISA|43|6|Dicam aquiloni: "Da"et austro: "Noli prohibere;affer filios meos de longinquoet filias meas ab extremis terrae.
ISA|43|7|Omnem, qui vocatur nomine meo,in gloriam meam creavi eum,formavi eum et feci eum".
ISA|43|8|Educ foras populum caecum, et oculos habentem,surdos, et aures eis sunt.
ISA|43|9|Omnes gentes congregentur simul,et colligantur nationes:quis in eis annuntiabit istudet priora audire nos faciet?Dent testes suos et iustificenturet audiant et dicant: "Vere".
ISA|43|10|Vos testes mei, dicit Dominus,et servus meus, quem elegi,ut sciatis et credatis mihiet intellegatis quia ego ipse sum;ante me non est formatus Deuset post me non erit.
ISA|43|11|Ego, ego sum Dominus,et non est absque me salvator.
ISA|43|12|Ego, annuntiavi et salvavi;auditum feci, et non fuit in vobis alienus;et vos testes mei, dicit Dominus,et ego Deus,
ISA|43|13|iam ab initio ego ipse.Et non est qui de manu mea eruat; operabor, et quis avertet illud? ".
ISA|43|14|Haec dicit Dominus, redemptor vester,Sanctus Israel: Propter vos misi in Babylonemet detraxi fugitivos universoset Chaldaeos in navibus suis gloriantes.
ISA|43|15|Ego Dominus, Sanctus vester,creans Israel, rex vester ".
ISA|43|16|Haec dicit Dominus,qui dedit in mari viamet in aquis torrentibus semitam;
ISA|43|17|qui eduxit quadrigam et equum,agmen et robustum;simul iacuerunt nec resurgent,contriti sunt quasi linum et exstincti sunt.
ISA|43|18|" Ne memineritis priorumet antiqua ne intueamini:
ISA|43|19|ecce ego facio nova,et nunc orientur: nonne cognoscitis ea?Utique ponam in deserto viamet in invio flumina.
ISA|43|20|Glorificabit me bestia agri,dracones et struthiones,quia dedi in deserto aquas,flumina in invio,ut darem potum populo meo, electo meo.
ISA|43|21|Populum istum formavi mihi;laudem meam narrabunt.
ISA|43|22|Non me invocasti, Iacob;immo taedio mei affectus es, Israel.
ISA|43|23|Non obtulisti mihi agnos holocausti tuiet victimis tuis non glorificasti me;non te gravavi in oblationenec laborem tibi praebui in ture.
ISA|43|24|Non emisti mihi argento calamumet adipe victimarum tuarum non inebriasti me;verumtamen servire me fecisti in peccatis tuis,praebuisti mihi laborem in iniquitatibus tuis.
ISA|43|25|Ego, ego sum ipse, qui deleo iniquitates tuas propter meet peccatorum tuorum non recordabor.
ISA|43|26|Memorem me redde, iudicium agamus simul:narra, ut iustificeris.
ISA|43|27|Pater tuus primus peccavit,et interpretes tui praevaricati sunt in me;
ISA|43|28|et contaminavi principes sanctuarii,dedi ad internecionem Iacobet Israel in opprobrium ".
ISA|44|1|Et nunc audi, Iacob serve meus,et Israel, quem elegi.
ISA|44|2|Haec dicit Dominus, qui fecit teet formavit te ab utero,auxiliator tuus: Noli timere, serve meus Iacob,et dilecte, quem elegi.
ISA|44|3|Effundam enim aquas super terram sitientemet fluenta super aridam;effundam spiritum meum super semen tuumet benedictionem meam super stirpem tuam:
ISA|44|4|et germinabunt inter herbasquasi salices iuxta praeterfluentes aquas.
ISA|44|5|Iste dicet: "Domini ego sum",et ille vocabit se nomine Iacob;et hic scribet manu sua: "Domino", et inscribetur nomine Israel ".
ISA|44|6|Haec dicit Dominus, rex Israelet redemptor eius, Dominus exercituum: Ego primus et ego novissimus,et absque me non est Deus.
ISA|44|7|Quis similis mei? Conclamet et annuntietet exponat mihi,ex quo constitui populum antiquum;ventura et, quae futura sunt, annuntiet nobis.
ISA|44|8|Nolite timere neque conturbemini;nonne ex tunc audire te feci et annuntiavi?Vos estis testes mei.Numquid est Deus absque meaut Petra, quam ego non noverim? ".
ISA|44|9|Plastae idoli omnes nihil sunt, et pretiosa eorum non proderunt eis; testes eorum non vident neque intellegunt, ut confundantur.
ISA|44|10|Quis formavit deum et sculptile conflavit lucrum non quaerens?
ISA|44|11|Ecce omnes participes eius confundentur; fabri enim sunt ex hominibus: conveniant omnes, stent; pavebunt, confundentur simul.
ISA|44|12|Faber ferrarius securim operatur in prunis et in malleis format illam et polit eam in brachio fortitudinis suae; esurit et deficit, non bibit aquam et lassescit.
ISA|44|13|Artifex lignarius extendit normam, describit illud stilo, operatur illud scalpellis et circino describit illud quasi imaginem viri, quasi speciosum hominem, qui resideat in domo.
ISA|44|14|Succidit sibi cedros et arripit ilicem et quercum, quae steterat inter ligna saltus; plantavit pinum, quam pluvia nutrivit.
ISA|44|15|Homini facta sunt ad comburendum; sumit ex eis, ut calefaciat, et succendit et coquit panes. De reliquo autem operatur deum et adorat; facit sculptile et curvatur ante illud.
ISA|44|16|Medium eius comburit igne et medio eius carnes assat, manducat assaturam et saturatur et calefit et dicit: " Vah, calefactus sum, vidi focum ".
ISA|44|17|Reliquum autem eius deum fecit, sculptile sibi; curvatur ante illud et adorat illud et obsecrat dicens: " Libera me, quia deus meus es tu ".
ISA|44|18|Nescierunt neque intellexerunt; nam clausit oculos eorum, ne videant et ne intellegant corde suo.
ISA|44|19|Non recogitant in corde suo, scientia et intellegentia carent, ut dicant: " Medietatem eius combussi igne et coxi super carbones eius panes, coxi carnes et comedi et de reliquo eius abominationem faciam; ante truncum ligni procidam? ".
ISA|44|20|Cinere vescitur; cor insipiens decepit eum, et non liberabit animam suam neque dicet: " Nonne mendacium est in dextera mea? ".
ISA|44|21|Memento horum, Iacob,et Israel, quoniam servus meus es tu;formavi te, servus meus es tu,Israel, non decipies me.
ISA|44|22|Delevi ut nubem iniquitates tuaset quasi nebulam peccata tua;revertere ad me,quoniam redemi te.
ISA|44|23|Exsultate, caeli, quoniam hoc fecit Dominus;iubilate, fundamenta terrae,resonate, montes, laudationem,saltus et omne lignum eius,quoniam redemit Dominus Iacobet in Israel glorificabitur.
ISA|44|24|Haec dicit Dominus, redemptor tuus et formator tuus ex utero: Ego sum Dominus, qui feci omnia,extendi caelos solus,expandi terram; et quis mecum?
ISA|44|25|Qui irrita facio signa divinorumet hariolos stultos reddo;compello sapientes retrorsumet scientiam eorum vanam facio;
ISA|44|26|qui suscito verbum servi meiet consilium nuntiorum meorum compleo.Qui dico Ierusalem: "Habitaberis" et civitatibus Iudae: "Aedificabimini"et deserta eius suscitabo;
ISA|44|27|qui dico profundo: "Desolare,et flumina tua arefaciam";
ISA|44|28|qui dico de Cyro: "Pastor meus estet omnem voluntatem meam complebit";qui dico Ierusalem: "Aedificaberis",et templo: "Fundaberis" ".
ISA|45|1|Haec dicit Dominus de uncto suo Cyro: Apprehendi dexteram eius,ut subiciam ante faciem eius genteset dorsa regum vertamet aperiam coram eo ianuas;et portae non claudentur.
ISA|45|2|Ego ante te iboet montes humiliabo;portas aereas conteramet vectes ferreos confringam.
ISA|45|3|Et dabo tibi thesauros absconditoset divitias occultas,ut scias quia ego Dominus,qui vocavi te nomine tuo, Deus Israel.
ISA|45|4|Propter servum meum Iacobet Israel electum meum,et vocavi te nomine tuo;designavi te, et non cognovisti me.
ISA|45|5|Ego Dominus, et non est amplius:extra me non est Deus.Accinxi te, et non cognovisti me,
ISA|45|6|ut sciant ab ortu solis et ab occidentequoniam absque me nullus est.Ego Dominus, et non est alter,
ISA|45|7|formans lucem et creans tenebras,faciens pacem et creans malum:ego Dominus faciens omnia haec.
ISA|45|8|Rorate, caeli, desuper, et nubes pluant iustitiam;aperiatur terraet germinet salvationem;et iustitia oriatur simul:ego Dominus creavi eam ".
ISA|45|9|Vae, qui contradicit fictori suo,testa de vasis fictilibus terrae!Numquid dicet lutum figulo suo: " Quid facis? "et " Opus tuum absque manibus est "?
ISA|45|10|Vae, qui dicit patri: " Quid generas? "et mulieri: " Quid parturis? ".
ISA|45|11|Haec dicit Dominus,Sanctus Israel, plastes eius: Numquid ventura interrogatis me super filios meoset super opus manuum mearum mandatis mihi?
ISA|45|12|Ego feci terramet hominem super eam creavi ego;manus meae tetenderunt caelos,et omni militiae eorum mandavi.
ISA|45|13|Ego suscitavi eum in iustitiaet omnes vias eius dirigam;ipse aedificabit civitatem meamet captivitatem meam dimittetnon in pretio neque in muneribus ",dicit Dominus exercituum.
ISA|45|14|Haec dicit Dominus: Labor Aegypti et negotiatio Aethiopiaeet Sabaim viri sublimesad te transibunt et tui erunt;post te ambulabunt,vincti manicis pergent et te adorabuntteque deprecabuntur:Tantum in te est Deus,et non est absque te Deus!".
ISA|45|15|Vere tu es Deus absconditus,Deus Israel, salvator.
ISA|45|16|Confusi sunt et erubuerunt omnes,simul abierunt in confusionem fabricatores idolorum.
ISA|45|17|Israel salvatus est in Domino salute aeterna;non confundemini et non erubescetisusque in saeculum saeculi.
ISA|45|18|Quia haec dicit Dominus,qui creavit caelos, ipse Deus,qui formavit terram et fecit eam, ipse fundavit eam;non ut vacua esset, creavit eam,ut habitaretur, formavit eam: Ego Dominus, et non est alius.
ISA|45|19|Non in abscondito locutus sum,in loco terrae tenebroso;non dixi semini Iacob:Frustra quaerite me".Ego Dominus loquens iustitiam,annuntians recta.
ISA|45|20|Congregamini et venite et accedite simul,qui salvati estis ex gentibus.Nescierunt, qui levant lignum sculpturae suaeet rogant deum non salvantem.
ISA|45|21|Annuntiate et venite et consiliamini simul.Quis auditum fecit hoc ab initio,ex tunc praedixit illud?Numquid non ego Dominus,et non est ultra Deus absque me?Deus iustus et salvans non est praeter me.
ISA|45|22|Convertimini ad me et salvi eritis,omnes fines terrae,quia ego Deus, et non est alius.
ISA|45|23|In memetipso iuravi:Egressa est de ore meo iustitia,verbum, quod non revertetur;quia mihi curvabitur omne genu,et iurabit omnis lingua ".
ISA|45|24|" Tantum in Domino " dicent sunt iustitiae et robur! ".Ad eum venient et confundenturomnes, qui repugnant ei;
ISA|45|25|in Domino iustificabitur et laudabituromne semen Israel.
ISA|46|1|Concidit Bel, incurvavit se Nabo;fuerunt simulacra eorum bestiis et iumentis.Statuae vestrae portantur, onera lassis.
ISA|46|2|Se incurvaverunt et conciderunt simul;non potuerunt salvare onuset ipsi in captivitatem ibunt.
ISA|46|3|Audite me, domus Iacobet omne residuum domus Israel,qui portamini ab utero,qui gestamini a vulva.
ISA|46|4|Usque ad senectam ego ipseet usque ad canos ego portabo;et ego feci et ego feram,ego portabo et salvabo.
ISA|46|5|Cui assimilatis me et adaequatiset comparatis me, et erimus similes?
ISA|46|6|Qui effundunt aurum de sacculoet argentum statera ponderant,conducunt aurificem, ut faciat deum,et procidunt et adorant.
ISA|46|7|Portant illum in umeris gestanteset ponentes in loco suo;et stabit ac de loco suo non movebitur;sed et si quis clamat ad eum, non respondet;de tribulatione eius non salvabit eum.
ISA|46|8|Mementote istud et confundamini;redite, praevaricatores, ad cor.
ISA|46|9|Recordamini prioris saeculi,quoniam ego sum Deus,et non est ultra Deus,nec est similis mei.
ISA|46|10|Annuntians ab exordio novissimumet ab initio, quae necdum facta sunt,dicens: " Consilium meum stabit,et omnem voluntatem meam faciam ".
ISA|46|11|Vocans ab oriente avem rapacemet de terra longinqua virum consilii mei;et locutus sum et adducam illud,decrevi et faciam illud.
ISA|46|12|Audite me, duri corde,qui longe estis a iustitia.
ISA|46|13|Prope feci iustitiam meam, non elongabitur;et salus mea non morabitur:et dabo in Sion salutemet Israeli gloriam meam.
ISA|47|1|Descende, sede in pulvere,virgo filia Babylon;sede in terra sine solio,filia Chaldaeorum,quia ultra non vocaberismollis et tenera.
ISA|47|2|Tolle molam et mole farinam;depone velum tuum,subleva stolam, revela crura,transi flumina.
ISA|47|3|Revelabitur ignominia tua,et videbitur opprobrium tuum. Ultionem capiam,nemini parcam ",
ISA|47|4|dicit Redemptor noster, Dominus exercituum nomen illius,Sanctus Israel.
ISA|47|5|Sede tacens et intra in tenebras,filia Chaldaeorum,quia non vocaberis ultraDomina regnorum.
ISA|47|6|Iratus sum super populum meum,contaminavi hereditatem meamet dedi eos in manu tua;non posuisti eis misericordias,super senem aggravasti iugum tuum valde
ISA|47|7|et dixisti: " In sempiternum ero domina ".Non posuisti haec super cor tuumneque recordata es novissimi tui.
ISA|47|8|Et nunc audi haec, delicata,quae habitas confidenteret dicis in corde tuo: Ego, et praeter me non est altera, non sedebo vidua et orbitatem ignorabo ".
ISA|47|9|Venient tibi duo haecsubito in die una,orbitas et viduitas;repente venerunt super tepropter multitudinem maleficiorum tuorum,propter abundantiam incantationum tuarum.
ISA|47|10|Et fiduciam habuisti in malitia tuaet dixisti: " Non est qui videat me ".Sapientia tua et scientia tua,haec decepit te.Et dixisti in corde tuo: Ego, et praeter me non est altera ".
ISA|47|11|Veniet super te malum,et nescies avertere;et irruet super te calamitas,quam non poteris expiare;veniet super te repentemiseria, quam nescies.
ISA|47|12|Sta cum incantationibus tuiset cum multitudine maleficiorum tuorum,in quibus laborasti ab adulescentia tua:forte poteris iuvari, forte terrebis.
ISA|47|13|Defecisti in multitudine consiliorum tuorum;stent et salvent te, qui metiuntur caelum,qui contemplantur sideraet annuntiant singulis noviluniisventura tibi.
ISA|47|14|Ecce facti sunt quasi stipula,ignis combussit eos.Non liberabunt seipsosde manu flammae;non sunt prunae, quibus calefiant,nec focus, ut sedeant ad eum.
ISA|47|15|Sic fiunt tibi incantatores tui,in quibuscumque laborasti ab adulescentia tua;unusquisque in via sua errat,non est qui salvet te.
ISA|48|1|Audite hoc, domus Iacob,qui vocamini nomine Israelet de aquis Iudae existis,qui iuratis in nomine Dominiet Deum Israel invocatisnon in veritate neque in iustitia.
ISA|48|2|De civitate enim sancta vocati suntet super Deum Israel constabiliti sunt;Dominus exercituum nomen eius.
ISA|48|3|Priora ex tunc annuntiavi,et ex ore meo exierunt,et audita feci ea;repente operatus sum, et venerunt.
ISA|48|4|Scivi enim quia durus es tu,et nervus ferreus cervix tua,et frons tua aerea.
ISA|48|5|Praedixi tibi ex tunc;antequam venirent, indicavi tibi,ne forte diceres: "Idolum meum operatum est haec,et sculptile meum et conflatile mandaverunt ista ".
ISA|48|6|Quae audisti, vide omnia;vos autem num annuntiabitis?Audita facio tibi nova ex nuncet occulta, quae nescis.
ISA|48|7|Nunc creata sunt et non ex tunc,et ante eorum diem, et non audisti ea,ne forte diceres: "Ecce ego cognovi ea ".
ISA|48|8|Neque audisti neque cognovisti,neque ex tunc aperta est auris tua;scio enim quia praevaricans praevaricariset transgressor ex utero vocaris.
ISA|48|9|Propter nomen meum longe faciam furorem meumet propter laudem meam infrenabo me super te,ne perdam te.
ISA|48|10|Ecce excoxi te, sed non quasi argentum;probavi te in camino paupertatis.
ISA|48|11|Propter me, propter me faciam,ut non blasphemer;et gloriam meam alteri non dabo.
ISA|48|12|Audi me, Iacob,et Israel, quem ego vocavi;ego, ego primuset ego novissimus.
ISA|48|13|Manus mea fundavit terram,et dextera mea expandit caelos;ego voco eos, et stant simul.
ISA|48|14|Congregamini, omnes vos, et audite:Quis de eis annuntiavit haec?Dominus dilexit eum;faciet voluntatem suam in Babyloneet brachium suum in Chaldaeis.
ISA|48|15|Ego, ego locutus sum et vocavi eum;adduxi eum, et prospera fuit via eius.
ISA|48|16|Accedite ad me et audite hoc:Non a principio in abscondito locutus sum;ex tempore, antequam fieret, ibi eram;et nunc Dominus Deus misit me cum spiritu suo.
ISA|48|17|Haec dicit Dominus,redemptor tuus, Sanctus Israel:Ego Dominus Deus tuus docens te utilia,gubernans te in via, qua ambulas.
ISA|48|18|Utinam attendisses mandata mea!Facta fuisset sicut flumen pax tua,et iustitia tua sicut gurgites maris;
ISA|48|19|et fuisset quasi arena semen tuum,et stirps uteri tui ut lapilli eius;non interisset et non fuisset attritumnomen eius a facie mea.
ISA|48|20|Egredimini de Babylone, fugite a Chaldaeis,in voce exsultationis annuntiate;auditum facite hoc, efferte illud usque ad extrema terrae,dicite: " Redemit Dominus servum suum Iacob ".
ISA|48|21|Non sitierunt, cum per desertum duceret eos;aquam de petra produxit eiset scidit petram, et fluxerunt aquae.
ISA|48|22|Non est pax impiis, dicit Dominus.
ISA|49|1|Audite me, insulae, et attendite, populi de longe;Dominus ab utero vocavit me,de ventre matris meae recordatus est nominis mei;
ISA|49|2|et posuit os meum quasi gladium acutum,in umbra manus suae protexit meet posuit me sicut sagittam electam,in pharetra sua abscondit me
ISA|49|3|et dixit mihi: " Servus meus es tu,Israel, in quo gloriabor ".
ISA|49|4|Et ego dixi: " In vacuum laboravi,sine causa et vane fortitudinem meam consumpsi;verumtamen iudicium meum cum Domino,et merces mea cum Deo meo ".
ISA|49|5|Et nunc dicit Dominus,qui formavit me ex utero servum sibi,ut reducerem Iacob ad eum,et Israel ei congregaretur;et glorificatus sum in oculis Domini,et Deus meus factus est fortitudo mea.
ISA|49|6|Et dixit: " Parum est ut sis mihi servusad suscitandas tribus Iacobet reliquias Israel reducendas:dabo te in lucem gentium,ut sit salus mea usque ad extremum terrae ".
ISA|49|7|Haec dicit Dominus,redemptor Israel, Sanctus eius,ad contemptum in anima,ad abominatum in gente,ad servum dominorum: Reges videbunt et consurgent,principes quoque et adorabunt,propter Dominum, quia fidelis est,Sanctum Israel, qui elegit te ".
ISA|49|8|Haec dicit Dominus: In tempore beneplaciti exaudivi teet in die salutis auxiliatus sum tui;et servavi te et dedi te in foedus populi,ut suscitares terramet distribueres hereditates dissipatas;
ISA|49|9|ut diceres his, qui vincti sunt: "Exite",et his, qui in tenebris: "Revelamini".Super vias pascentur,et in omnibus collibus decalvatis pascua eorum;
ISA|49|10|non esurient neque sitient,et non percutiet eos aestus vel sol,quia miserator eorum reget eoset ad fontes aquarum adducet eos.
ISA|49|11|Et ponam omnes montes meos in viam,et semitae meae exaltabuntur.
ISA|49|12|Ecce isti de longe venient,et ecce illi ab aquilone et mari,et isti de terra Sinim ".
ISA|49|13|Laudate, caeli, et exsulta, terra;iubilate, montes, laudem,quia consolatur Dominus populum suumet pauperum suorum miseretur.
ISA|49|14|Et dixit Sion: " Dereliquit me Dominus,et Dominus oblitus est mei ".
ISA|49|15|Numquid oblivisci potest mulier infantem suum,ut non misereatur filio uteri sui?Et si illa oblita fuerit,ego tamen non obliviscar tui.
ISA|49|16|Ecce in manibus meis descripsi te;muri tui coram me semper.
ISA|49|17|Festinant structores tui;destruentes te et dissipantes a te exibunt.
ISA|49|18|Leva in circuitu oculos tuos et vide:omnes isti congregati sunt, venerunt tibi. Vivo ego, dicit Dominus,quia omnibus his velut ornamento vestieriset circumdabis tibi eos quasi sponsa ".
ISA|49|19|Quia ruinae tuae et solitudines tuaeet terra eversa:nunc angusta eris prae habitatoribus;et longe erunt, qui devorabant te.
ISA|49|20|Adhuc dicent in auribus tuisfilii orbitatis tuae: Angustus est mihi locus;fac spatium mihi, ut habitem ".
ISA|49|21|Et dices in corde tuo: Quis genuit mihi istos?Ego orbata et non pariens,transmigrata et captiva;et istos quis enutrivit?Ecce ego relicta eram sola;et isti ubi erant? ".
ISA|49|22|Haec dicit Dominus Deus: Ecce levabo ad gentes manum meamet ad populos exaltabo signum meum;et afferent filios tuos in ulnis,et filiae tuae super umeros portabuntur.
ISA|49|23|Et erunt reges nutricii tui,et reginae nutrices tuae;vultu in terram demisso adorabunt teet pulverem pedum tuorum lingent.Et scies quia ego Dominus:non confundentur, qui sperant in me ".
ISA|49|24|Numquid tolletur a forti praeda,aut, quod captum fuerit, a robusto salvari poterit?
ISA|49|25|Quia haec dicit Dominus: Equidem et captivus a forti tolletur,et, quod ablatum fuerit a robusto, salvabitur;cum his, qui contendebant tecum, ego contendamet filios tuos ego salvabo.
ISA|49|26|Et cibabo hostes tuos carnibus suis,et quasi musto sanguine suo inebriabuntur;et sciet omnis caro quia ego Dominus salvator tuus,et redemptor tuus Fortis Iacob ".
ISA|50|1|Haec dicit Dominus: Ubinam est liber repudii matris vestrae,quo dimisi eam?Aut quis est creditor meus,cui vendidi vos?Ecce in iniquitatibus vestris venditi estis,et in sceleribus vestris dimissa est mater vestra.
ISA|50|2|Cur veni, et non erat vir,vocavi, et non erat qui responderet?Numquid abbreviata est manus mea,ut non possim redimere?Aut non est in me virtus ad liberandum?Ecce in increpatione mea exsiccabo mare,ponam flumina in siccum;computrescent pisces sine aquaet morientur in siti.
ISA|50|3|Induam caelos luctuet saccum ponam operimentum eorum ".
ISA|50|4|Dominus Deus dedit mihi linguam eruditam,ut sciam sustentare eum, qui lassus est, verbo;excitat mane, mane excitat mihi aurem,ut audiam quasi discipulus.
ISA|50|5|Dominus Deus aperuit mihi aurem;ego autem non rebellavi, retrorsum non abii.
ISA|50|6|Dorsum meum dedi percutientibuset genas meas vellentibus:faciem meam non avertiab increpationibus et sputis.
ISA|50|7|Dominus Deus auxiliator meus;ideo non sum confusus,ideo posui faciem meam ut petram durissimamet scio quoniam non confundar.
ISA|50|8|Iuxta est qui iustificat me;quis contradicet mihi? Stemus simul.Quis est adversarius meus? Accedat ad me.
ISA|50|9|Ecce Dominus Deus auxiliator meus;quis est qui condemnet me?Ecce omnes quasi vestimentum conterentur,tinea comedet eos.
ISA|50|10|Quis ex vobis timet Dominum,audiens vocem servi sui?Qui ambulavit in tenebris,et non est lumen ei,speret in nomine Dominiet innitatur super Deum suum.
ISA|50|11|Ecce vos omnes, qui accenditis ignem,accincti sagittis,ambulate in lumine ignis vestriet in sagittis, quas succendistis.De manu mea factum est hoc vobis;in doloribus recumbetis.
ISA|51|1|Audite me, qui sequimini iustitiam,qui quaeritis Dominum;attendite ad petram, unde excisi estis,et ad cavernam laci, de qua praecisi estis.
ISA|51|2|Attendite ad Abraham patrem vestrumet ad Saram, quae peperit vos;quia unum vocavi eumet benedixi ei et multiplicavi eum.
ISA|51|3|Consolatur enim Dominus Sion,consolatur omnes ruinas eius;et ponit desertum eius quasi Edenet solitudinem eius quasi hortum Domini.Gaudium et laetitia invenietur in ea,gratiarum actio et vox laudis.
ISA|51|4|Attendite ad me, popule meus;et nationes, me audite,quia lex a me exiet,et iudicium meum in lucem populorum statuam.
ISA|51|5|Prope est iustitia mea,egressa est salus mea,et brachia mea populos iudicabunt;in me insulae sperabuntet ad brachium meum attendent.
ISA|51|6|Levate in caelum oculos vestroset inspicite in terram deorsum,quia caeli sicut fumus liquescent,et terra sicut vestimentum atteretur,et habitatores eius sicut haec interibunt.Salus autem mea in sempiternum erit,et iustitia mea non deficiet.
ISA|51|7|Audite me, qui scitis iustitiam,popule, in cuius corde est lex mea:nolite timere opprobrium hominumet blasphemias eorum ne metuatis.
ISA|51|8|Sicut enim vestimentum sic comedet eos vermis,et sicut lanam sic devorabit eos tinea;iustitia autem mea in sempiternum erit,et salus mea in generationes generationum.
ISA|51|9|Consurge, consurge, induere fortitudinem,brachium Domini;consurge sicut in diebus antiquis,in generationibus saeculorum.Numquid non tu percussisti Rahab,vulnerasti draconem?
ISA|51|10|Numquid non tu siccasti mare,aquam abyssi vehementis,qui posuisti profundum maris viam,ut transirent liberati?
ISA|51|11|Et redempti a Domino revertenturet venient in Sion laudantes;et laetitia sempiterna super capita eorum,gaudium et laetitiam obtinebunt;fugiet dolor et gemitus.
ISA|51|12|Ego, ego ipse consolator vester.Quis tu, ut timeas ab homine mortaliet a filio hominis, qui quasi fenum ita arescet?
ISA|51|13|Et oblitus es Domini factoris tui,qui tetendit caelos et fundavit terram;et formidasti iugiter tota diea facie furoris eius, qui te tribulabat,cum parabat ad perdendum.Ubi nunc est furor tribulantis?
ISA|51|14|Cito captivus liberabituret non morietur in fovea,nec deficiet panis eius.
ISA|51|15|Ego enim sum Dominus Deus tuus,qui conturbo mare,et intumescunt fluctus eius;Dominus exercituum nomen eius.
ISA|51|16|Posui verba mea in ore tuoet in umbra manus meae protexi te,cum extendebam caelos et fundabam terramet dicebam ad Sion: "Populus meus es tu ".
ISA|51|17|Elevare, elevare, consurge, Ierusalem,quae bibisti de manu Domini calicem irae eius;poculum soporis bibisti,epotasti.
ISA|51|18|Non est qui sustentet eamex omnibus filiis, quos genuit;et non est qui apprehendat manum eiusex omnibus filiis, quos enutrivit.
ISA|51|19|Duo sunt quae occurrerunt tibi;quis contristabitur super te?Vastitas et contritio et fames et gladius;quis consolabitur te?
ISA|51|20|Filii tui defecerunt,iacent in capite omnium viarumsicut oryx illaqueatus,pleni indignatione Domini,increpatione Dei tui.
ISA|51|21|Idcirco audi hoc, pauperculaet ebria, sed non a vino.
ISA|51|22|Haec dicit dominator tuus,Dominus et Deus tuus, qui contendit pro populo suo: Ecce tuli de manu tua calicem soporis,poculum indignationis meae;non adicies, ut bibas illum ultra.
ISA|51|23|Et ponam illum in manu eorum, qui te humiliaveruntet dixerunt tibi: "Incurvare, ut transeamus";et ponebas ut terram dorsum tuumet quasi viam transeuntibus ".
ISA|52|1|Consurge, consurge,induere fortitudine tua, Sion;induere vestimentis gloriae tuae,Ierusalem, civitas sanctitatis,quia non adiciet ultra, ut pertranseat per teincircumcisus et immundus.
ISA|52|2|Excutere de pulvere, consurge,captiva Ierusalem;solve vincula colli tui,captiva filia Sion.
ISA|52|3|Quia haec dicit Dominus: " Gratis venumdati estis et sine argento redimemini ".
ISA|52|4|Quia haec dicit Dominus Deus: " In Aegyptum descendit populus meus in principio, ut colonus esset ibi; et Assur sine causa oppressit eum.
ISA|52|5|Et nunc quid mihi est hic, dicit Dominus, quoniam ablatus est populus meus gratis? Dominatores eius ululant, dicit Dominus, et iugiter tota die nomen meum blasphematur.
ISA|52|6|Propter hoc sciet populus meus nomen meum in die illa, quia ego ipse, qui loquebar: "Ecce adsum" ".
ISA|52|7|Quam pulchri super montespedes annuntiantis, praedicantis pacem,annuntiantis bonum, praedicantis salutem,dicentis Sion: "Regnavit Deus tuus!".
ISA|52|8|Vox speculatorum tuorum: levaverunt vocem,simul exsultabunt,quia oculo ad oculum videbunt,cum redierit Dominus ad Sion.
ISA|52|9|Gaudete et exsultate simul,deserta Ierusalem,quia consolatus est Dominus populum suum,redemit Ierusalem.
ISA|52|10|Nudavit Dominus brachium sanctum suumin oculis omnium gentium;et videbunt omnes fines terraesalutare Dei nostri.
ISA|52|11|Recedite, recedite, exite inde,pollutum nolite tangere;exite de medio eius, mundamini,qui fertis vasa Domini.
ISA|52|12|Quoniam non in festinatione exibitisnec in fuga properabitis;praecedet enim vos Dominus,et colliget vos Deus Israel.
ISA|52|13|Ecce prospere aget servus meus;exaltabitur et elevabitur et sublimis erit valde.
ISA|52|14|Sicut obstupuerunt super eum multi,sic deformis erat, quasi non esset hominis species eius,filiorum hominis aspectus eius,
ISA|52|15|sic disperget gentes multas.Super ipsum continebunt reges os suum,quia, quae non sunt narrata eis, videruntet, quae non audierunt, contemplati sunt.
ISA|53|1|" Quis credidit auditui nostro,et brachium Domini cui revelatum est?
ISA|53|2|Et ascendit sicut virgultum coram eoet sicut radix de terra sitienti.Non erat species ei neque decor, ut aspiceremus eum,et non erat aspectus, ut desideraremus eum.
ISA|53|3|Despectus erat et novissimus virorum,vir dolorum et sciens infirmitatem,et quasi abscondebamus vultum coram eo;despectus, unde nec reputabamus eum.
ISA|53|4|Vere languores nostros ipse tulitet dolores nostros ipse portavit;et nos putavimus eum quasi plagatum,percussum a Deo et humiliatum.
ISA|53|5|Ipse autem vulneratus est propter iniquitates nostras,attritus est propter scelera nostra;disciplina pacis nostrae super eum,et livore eius sanati sumus.
ISA|53|6|Omnes nos quasi oves erravimus,unusquisque in viam suam declinavit;et posuit Dominus in eoiniquitatem omnium nostrum ".
ISA|53|7|Afflictus est et ipse subiecit seet non aperuit os suum;sicut agnus, qui ad occisionem ducitur,et quasi ovis, quae coram tondentibus se obmutuitet non aperuit os suum.
ISA|53|8|Angustia et iudicio sublatus est.De generatione eius quis curabit?Quia abscissus est de terra viventium;propter scelus populi mei percussus est ad mortem.
ISA|53|9|Et posuerunt sepulcrum eius cum impiis,cum divitibus tumulum eius,eo quod iniquitatem non fecerit,neque dolus fuerit in ore eius.
ISA|53|10|Et Dominus voluit conterere eum infirmitate.Si posuerit in piaculum animam suam,videbit semen longaevum,et voluntas Domini in manu eius prosperabitur.
ISA|53|11|Propter laborem animae eiusvidebit lucem, saturabitur in scientia sua.Iustificabit iustus servus meus multoset iniquitates eorum ipse portabit.
ISA|53|12|Ideo dispertiam ei multos,et cum fortibus dividet spolia,pro eo quod tradidit in mortem animam suamet cum sceleratis reputatus est;et ipse peccatum multorum tulitet pro transgressoribus rogat.
ISA|54|1|Exsulta, sterilis, quae non peperisti,laetare, gaude, quae non parturisti,quoniam multi sunt filii desertaemagis quam filii nuptae, dicit Dominus.
ISA|54|2|Dilata locum tentorii tuiet pelles tabernaculorum tuorum extende, ne parcas;longos fac funiculos tuoset clavos tuos consolida.
ISA|54|3|Ad dexteram enim et ad laevam penetrabis,et semen tuum hereditabit gentes,quae civitates desertas inhabitabunt.
ISA|54|4|Noli timere, quia non confunderis,neque erubescas, quia non te pudebit;nam confusionis adulescentiae tuae oblivisceriset opprobrii viduitatis tuae non recordaberis amplius.
ISA|54|5|Qui enim fecit te, erit sponsus tuus,Dominus exercituum nomen eius;et redemptor tuus Sanctus Israel,Deus omnis terrae vocabitur.
ISA|54|6|Quia ut mulierem derelictam et maerentem spirituvocavit te Dominus,et uxorem ab adulescentia abiectamdixit Deus tuus.
ISA|54|7|Ad punctum in modico dereliqui teet in miserationibus magnis congregabo te.
ISA|54|8|In momento indignationisabscondi faciem meam parumper a teet in misericordia sempiterna misertus sum tui,dixit redemptor tuus Dominus.
ISA|54|9|Sicut in diebus Noe istud mihi est,cui iuravi, ne inducerem aquas Noe ultra supra terram;sic iuravi, ut non irascar tibiet non increpem te.
ISA|54|10|Montes enim recedent,et colles movebuntur,misericordia autem mea non recedet a te,et foedus pacis meae non movebitur,dixit miserator tuus Dominus.
ISA|54|11|Paupercula, tempestate convulsa absque ulla consolatione,ecce ego sternam super carbunculos lapides tuoset fundabo te in sapphiris;
ISA|54|12|et ponam iaspidem propugnacula tuaet portas tuas in lapides pretiososet omnes terminos tuos in lapides desiderabiles.
ISA|54|13|Universi filii tui erunt discipuli Domini,et magna erit pax filiis tuis;
ISA|54|14|in iustitia fundaberis.Procul eris ab oppressione, quia non timebis,et a pavore, quia non appropinquabit tibi.
ISA|54|15|Ecce, si impetus fiet, non erit ex me; qui impetum fecerit in te, cadet contra te.
ISA|54|16|Ecce, ego creavi fabrumsufflantem in igne prunaset proferentem vas in opus suum;et ego creavi etiam vastatorem ad disperdendum.
ISA|54|17|Omne vas, quod fictum est contra te, frustra erit.Et omnem linguam insurgentem tibi in iudicio confutabis:haec est hereditas servorum Dominiet iustitia eorum ex me, dicit Dominus.
ISA|55|1|Heu! Omnes sitientes, venite ad aquas;et, qui non habetis argentum, properate,emite et comedite, venite, emite absque argentoet absque ulla commutatione vinum et lac.
ISA|55|2|Quare appenditis argentum non in panibuset laborem vestrum non in saturitate?Audite, audientes me, et comedite bonum,ut delectetur in crassitudine anima vestra.
ISA|55|3|Inclinate aurem vestram et venite ad me;audite, ut vivat anima vestra,et feriam vobiscum pactum sempiternum,misericordias David fideles.
ISA|55|4|Ecce testem populis dedi eum,ducem ac praeceptorem gentibus.
ISA|55|5|Ecce gentem, quam nesciebas, vocabis,et gentes, quae te non cognoverunt, ad te current,propter Dominum Deum tuumet Sanctum Israel, quia glorificavit te.
ISA|55|6|Quaerite Dominum, dum inveniri potest;invocate eum, dum prope est.
ISA|55|7|Derelinquat impius viam suam,et vir iniquus cogitationes suas;et revertatur ad Dominum, et miserebitur eius,et ad Deum nostrum, quoniam multus est ad ignoscendum.
ISA|55|8|Non enim cogitationes meae cogitationes vestrae,neque viae vestrae viae meae, dicit Dominus.
ISA|55|9|Quia sicut exaltantur caeli a terra,sic exaltatae sunt viae meae a viis vestris,et cogitationes meae a cogitationibus vestris.
ISA|55|10|Et quomodo descendit imber et nix de caeloet illuc ultra non revertitur,sed inebriat terram et infundit eamet germinare eam facitet dat semen serenti et panem comedenti,
ISA|55|11|sic erit verbum meum, quod egredietur de ore meo:non revertetur ad me vacuum,sed faciet, quaecumque volui,et prosperabitur in his, ad quae misi illud.
ISA|55|12|Quia in laetitia egredieminiet in pace deducemini;montes et colles cantabunt coram vobis laudem,et omnia ligna regionis plaudent manu.
ISA|55|13|Pro vepribus ascendet cupressus,et pro urtica crescet myrtus;et erit Domino in gloriam,in signum aeternum, quod non auferetur.
ISA|56|1|Haec dicit Dominus: Custodite iudicium et faciteiustitiam,quia iuxta est salus mea, ut veniat,et iustitia mea, ut reveletur ".
ISA|56|2|Beatus vir, qui facit hoc,et filius hominis, qui apprehendit istud,custodiens sabbatum, ne polluat illud,custodiens manum suam, ne faciat omne malum.
ISA|56|3|Et non dicat filius advenae, qui adhaeret Domino,dicens: " Separatione dividet me Dominus a populo suo ".Et non dicat eunuchus: Ecce, ego lignum aridum ".
ISA|56|4|Quia haec dicit Dominus eunuchis: Qui custodierint sabbata meaet elegerint, quae ego volui,et tenuerint foedus meum,
ISA|56|5|dabo eis in domo mea et in muris meislocum et nomen melius a filiis et filiabus:nomen sempiternum dabo eis,quod non peribit.
ISA|56|6|Et filios advenae, qui adhaerent Domino,ut colant eum,ut diligant nomen Domini,ut sint ei in servos,omnes custodientes sabbatum, ne polluant illud,et tenentes foedus meum,
ISA|56|7|adducam eos in montem sanctum meumet laetificabo eos in domo orationis meae:holocausta eorum et victimae eorumplacebunt mihi super altari meo,quia domus mea domus orationisvocabitur cunctis populis ".
ISA|56|8|Ait Dominus Deus, qui congregat dispersos Israel: Adhuc congregabo ad eum praeter congregatos eius ".
ISA|56|9|Omnes bestiae agri, venite ad devorandum,universae bestiae saltus.
ISA|56|10|Speculatores eius caeci, omnes nescierunt;universi sunt canes muti non valentes latrare,insanientes, cubantes, amantes soporem;
ISA|56|11|et canes voraces nescierunt saturitatem,ipsi pastores ignoraverunt intellegentiam:omnes in viam suam declinaverunt,unusquisque ad avaritiam suam,a summo usque ad novissimum.
ISA|56|12|" Venite, sumam vinum, et impleamur ebrietate;et cras erit sicut hodieet multo amplius ".
ISA|57|1|Iustus perit, et non est qui recogitet in corde suo;et viri misericordiae colliguntur,tamen non est qui intellegat:a facie enim malitiae collectus est iustus.
ISA|57|2|In pacem ingreditur, requiescit in cubili suo,qui ambulat in directione sua.
ISA|57|3|Vos autem accedite huc, filii auguratricis,semen adulteri et fornicariae.
ISA|57|4|Super quem luditis?Super quem dilatatis os et eicitis linguam?Numquid non vos filii scelesti, semen mendax,
ISA|57|5|qui exardescitis in terebinthissubter omne lignum frondosum,immolantes parvulos in vallibussubter scissuras petrarum?
ISA|57|6|In partibus vallis pars tua,hae sunt sors tua;et ipsis effundisti libamen, obtulisti sacrificium.Numquid super his consolabor?
ISA|57|7|Super montem excelsum et sublimem posuisti cubile tuum,et illuc ascendisti, ut immolares hostias.
ISA|57|8|Et post ostium et postem posuisti memoriale tuum;nam longe a me discooperuisti et ascendisti,dilatasti cubile tuum,et pepigisti cum eis foedus;dilexisti stratum eorum, manum respexisti.
ISA|57|9|Et ingressa es ad regem cum unguentoet multiplicasti pigmenta tua;misisti legatos tuos proculet humiliata es usque ad inferos.
ISA|57|10|In multitudine viae tuae laborasti;non dixisti: " Vanum est! ".Vitam manus tuae invenisti,propterea non aegrotasti.
ISA|57|11|Pro quo sollicita timuisti,quia mentita es et mei non es recordataneque cogitasti in corde tuo?Nonne, quia ego tacui et longo tempore,me non times?
ISA|57|12|Ego annuntiabo iustitiam tuamet opera tua, quae non proderunt tibi.
ISA|57|13|Cum clamaveris, liberent te lucra tua;et omnia illa auferet ventus, tollet aura.Qui autem fiduciam habet in me, hereditabit terramet possidebit montem sanctum meum.
ISA|57|14|Et dicent: " Sternite, sternite,parate viam, auferte offendicula de via populi mei ".
ISA|57|15|Quia haec dicit Excelsus et Sublimis,habitans aeternitatem, et sanctum nomen eius: Excelsus et sanctus habitoet cum contrito et humili spiritu,ut vivificem spiritum humiliumet vivificem cor contritorum.
ISA|57|16|Non enim in sempiternum litigaboneque usque ad finem irascar,quia spiritus a facie mea deficeret,halitus, quem ego feci.
ISA|57|17|Propter iniquitatem avaritiae eius iratus sum et percussi eum,abscondi faciem meam et indignatus sum;et abiit vagus in via cordis sui.
ISA|57|18|Vias eius vidi et sanabo eum et reducam eumet reddam consolationes ipsi et lugentibus eius.
ISA|57|19|Creo fructum labiorum pacem;pacem ei, qui longe est et qui prope, dixit Dominus,et sanabo eum ".
ISA|57|20|Impii autem quasi mare fervens,quod quiescere non potest,et redundant fluctus eius in limum et lutum.
ISA|57|21|Non est pax impiis, dicit Deus meus.
ISA|58|1|Clama fortiter, ne cesses;quasi tuba exalta vocem tuamet annuntia populo meo scelera eorumet domui Iacob peccata eorum.
ISA|58|2|Me etenim de die in diem quaerunt et scire vias meas volunt,quasi gens, quae iustitiam feceritet iudicium Dei sui non dereliquerit.Rogant me iudicia iustitiae,appropinquare Deum volunt.
ISA|58|3|" Quare ieiunavimus, et non aspexisti,humiliavimus animam nostram, et nescisti? ".Ecce, in die ieiunii vestri agitis negotiaet omnes operarios vestros opprimitis.
ISA|58|4|Ecce, ad lites et contentiones ieiunatiset percutitis pugno impie.Nolite ieiunare sicut hodie,ut audiatur in excelso clamor vester.
ISA|58|5|Numquid tale est ieiunium, quod elegi,dies, quo homo affligit animam suam?Numquid contorquere quasi iuncum caput suumet saccum et cinerem sternere?Numquid istud vocabis ieiuniumet diem acceptabilem Domino?
ISA|58|6|Nonne hoc est ieiunium, quod elegi:dissolvere vincula iniqua,solvere funes iugi,dimittere eos, qui confracti sunt, liberos,et omne iugum dirumpere?
ISA|58|7|Nonne frangere esurienti panem tuum,et egenos, vagos inducere in domum?Cum videris nudum, operi eumet carnem tuam ne despexeris.
ISA|58|8|Tunc erumpet quasi aurora lumen tuum,et sanatio tua citius orietur;et anteibit faciem tuam iustitia tua,et gloria Domini colliget te.
ISA|58|9|Tunc invocabis, et Dominus exaudiet;clamabis, et dicet: " Ecce adsum ".Si abstuleris de medio tui iugumet desieris extendere digitumet loqui iniquitatem;
ISA|58|10|si effuderis esurienti animam tuamet animam afflictam satiaveris,orietur in tenebris lux tua,et caligo tua erit sicut meridies.
ISA|58|11|Et te ducet Dominus semper,et satiabit in locis aridis animam tuamet ossa tua firmabit;et eris quasi hortus irriguuset sicut fons aquarum,cuius non deficient aquae.
ISA|58|12|Et reaedificabit gens tua ruinas antiquas;fundamenta generationis et generationis suscitabis:et vocaberis restitutor ruinarum,instaurator viarum, ut habitentur.
ISA|58|13|Si averteris a sabbato pedem tuum,facere negotia tua in die sancto meo,et vocaveris sabbatum deliciaset diem Domino sacrum gloriosum;et glorificaveris eum relinquens vias tuaset negotia tua et sermones tuos,
ISA|58|14|tunc delectaberis super Domino;et vehi te faciam super altitudines terraeet cibabo te hereditate Iacob patris tui.Os enim Domini locutum est.
ISA|59|1|Ecce non est abbreviata manus Domini,ut salvare nequeat,neque aggravata est auris eius,ut non exaudiat;
ISA|59|2|sed iniquitates vestrae diviseruntinter vos et Deum vestrum,et peccata vestra absconderunt faciem eiusa vobis, ne exaudiret.
ISA|59|3|Manus enim vestrae pollutae sunt sanguine,et digiti vestri iniquitate;labia vestra locuta sunt mendacium,et lingua vestra iniquitatem fatur.
ISA|59|4|Non est qui invocet iustitiam,neque est qui iudicet vere;confidunt in nihilo et loquuntur vanitates:conceperunt laborem et pepererunt iniquitatem.
ISA|59|5|Ova aspidum rumpuntet telas araneae texunt;qui comederit de ovis eorum, morietur,et, quod fractum est, erumpet in regulum.
ISA|59|6|Telae eorum non erunt in vestimentum,neque operientur operibus suis;opera eorum opera iniquitatis,et facinora violentiae in manibus eorum.
ISA|59|7|Pedes eorum ad malum curruntet festinant, ut effundant sanguinem innocentem;cogitationes eorum cogitationes iniquitatis,vastitas et contritio in viis eorum.
ISA|59|8|Viam pacis nescierunt,et non est iudicium in gressibus eorum;semitae eorum incurvatae sunt eis:omnis, qui calcat in eis, ignorat pacem.
ISA|59|9|Propter hoc elongatum est iudicium a nobis,et non apprehendit nos iustitia;exspectamus lucem, et ecce tenebrae,splendorem, et in caligine ambulamus.
ISA|59|10|Palpamus sicut caeci parietemet quasi absque oculis attrectamus;impegimus meridie quasi in crepusculo,inter sanos quasi mortui.
ISA|59|11|Rugimus quasi ursi omneset quasi columbae gementes gemimus;exspectamus iudicium, et non est,salutem, et elongata est a nobis.
ISA|59|12|Multiplicatae sunt enim iniquitates nostrae coram te,et peccata nostra respondent nobis;quia scelera nostra nobiscum,et iniquitates nostras cognovimus:
ISA|59|13|peccare et mentiri contra Dominumet recedere a Deo nostro,loqui violentiam et transgressionem,concipere et murmurare de corde verba mendacii.
ISA|59|14|Et conversum est retrorsum iudicium,et iustitia longe stat,quia corruit in platea veritas,et aequitas non potuit ingredi.
ISA|59|15|Et facta est veritas in oblivionem,et, qui recedit a malo, spoliatur.Et vidit Dominus, et malum apparuit in oculis eius,quia non est iudicium.
ISA|59|16|Et vidit quia non est vir,et aporiatus est, quia non est qui occurrat;et salvavit sibi brachium suum,et iustitia eius ipsa confirmavit eum.
ISA|59|17|Indutus est iustitia ut lorica,et galea salutis in capite eius;indutus est vestimentis ultioniset operuit se zelo quasi pallio.
ISA|59|18|Secundum opera sic retribuet:iram hostibus suis,retributionem inimicis suis,insulis vicem reddet.
ISA|59|19|Et timebunt, qui ab occidente, nomen Domini,et, qui ab ortu solis, gloriam eius,cum venerit quasi fluvius violentus,quem spiritus Domini cogit.
ISA|59|20|Et veniet pro Sion redemptoret eis, qui redeunt ab iniquitate in Iacob,dixit Dominus.
ISA|59|21|Hoc foedus meum cum eis,dixit Dominus: Spiritus meus, qui est super te,et verba mea, quae posui in ore tuo,non recedent de ore tuoet de ore seminis tuiet de ore seminis seminis tui,dixit Dominus, amodo et usque in sempiternum ".
ISA|60|1|Surge, illuminare, quia venit lumen tuum,et gloria Domini super te orta est.
ISA|60|2|Quia ecce tenebrae operient terramet caligo populos;super te autem orietur Dominus,et gloria eius in te videbitur.
ISA|60|3|Et ambulabunt gentes in lumine tuo,et reges in splendore ortus tui.
ISA|60|4|Leva in circuitu oculos tuos et vide:omnes isti congregati sunt, venerunt tibi;filii tui de longe veniunt,et filiae tuae in ulnis gestantur.
ISA|60|5|Tunc videbis et illuminaberis,et palpitabit et dilatabitur cor tuum,quia confluet ad te multitudo maris,fortitudo gentium veniet tibi;
ISA|60|6|inundatio camelorum operiet te,dromedarii Madian et Epha;omnes de Saba venient,aurum et tus deferenteset laudem Domini annuntiantes.
ISA|60|7|Omne pecus Cedar congregabitur tibi,arietes Nabaioth ministrabunt tibi;offerentur super placabili altari meo,et domum gloriae meae glorificabo.
ISA|60|8|Quae sunt istae, quae ut nubes volant,et quasi columbae ad fenestras suas?
ISA|60|9|Me enim insulae exspectabunt,et in principio naves Tharsis,ut adducant filios tuos de longe,argentum eorum et aurum eorum cum eis,nomini Domini Dei tui et Sancto Israel,quia glorificavit te.
ISA|60|10|Et aedificabunt filii peregrinorum muros tuos,et reges eorum ministrabunt tibi;in indignatione enim mea percussi te,sed in beneplacito meo misertus sum tui.
ISA|60|11|Et aperientur portae tuae iugiter,die ac nocte non claudentur,ut afferatur ad te fortitudo gentium,et reges earum adducantur.
ISA|60|12|Gens enim et regnum, quae non servierint tibi, peribunt,et gentes vastitate vastabuntur.
ISA|60|13|Gloria Libani ad te veniet,cupressus, ulmus et abies simul,ad ornandum locum sanctuarii mei;et locum pedum meorum glorificabo.
ISA|60|14|Et venient ad te curvi filii eorum, qui humiliaverunt te,et adorabunt vestigia pedum tuorum omnes, qui detrahebant tibi, et vocabunt te Civitatem Domini,Sion Sancti Israel.
ISA|60|15|Pro eo quod fuisti derelicta et odio habita,et non erat qui per te transiret,ponam te in superbiam saeculorum,gaudium in generationem et generationem;
ISA|60|16|et suges lac gentiumet mamilla regum lactaberiset scies quia ego Dominus salvator tuus,et redemptor tuus Fortis Iacob.
ISA|60|17|Pro aere afferam aurumet pro ferro afferam argentumet pro lignis aeset pro lapidibus ferrum;et ponam custodes tuos pacemet praepositos tuos iustitiam.
ISA|60|18|Non audietur ultra violentia in terra tua,vastitas et contritio in terminis tuis;et vocabis Salutem muros tuoset portas tuas Laudem.
ISA|60|19|Non erit tibi amplius sol ad lucendum per diem,nec splendor lunae illuminabit te,sed erit tibi Dominus in lucem sempiternam,et Deus tuus in gloriam tuam.
ISA|60|20|Non occidet ultra sol tuus,et luna tua non minuetur,quia erit tibi Dominus in lucem sempiternam,et complebuntur dies luctus tui.
ISA|60|21|Populus autem tuus omnes iusti;in perpetuum hereditabunt terram,germen plantationis meae,opus manus meae ad glorificandum.
ISA|60|22|Minimus erit in mille,et parvulus in gentem fortem.Ego Dominus in tempore eius subito faciam istud.
ISA|61|1|Spiritus Domini Dei super me,eo quod unxerit Dominus me;ad annuntiandum laeta mansuetis misit me,ut mederer contritis cordeet praedicarem captivis liberationemet clausis apertionem;
ISA|61|2|ut praedicarem annum placabilem Dominoet diem ultionis Deo nostro;ut consolarer omnes lugentes,
ISA|61|3|ut ponerem lugentibus Sionet darem eis coronam pro cinere,oleum gaudii pro luctu,pallium laudis pro spiritu maeroris.Et vocabuntur Terebinthi iustitiae,plantatio Domini ad glorificandum.
ISA|61|4|Et aedificabunt deserta a saeculoet ruinas antiquas erigentet instaurabunt civitates desertas,dissipatas in generatione et generatione.
ISA|61|5|Et stabunt alieni et pascent pecora vestra,et filii peregrinorum agricolae et vinitores vestri erunt;
ISA|61|6|vos autem Sacerdotes Domini vocabimini,Ministri Dei nostri dicetur vobis;fortitudinem gentium comedetiset in gloria earum superbietis.
ISA|61|7|Pro confusione eorum dupliciet ignominia laudabunt partem suam;propterea in terra sua duplicia possidebunt,laetitia sempiterna erit eis.
ISA|61|8|Quia ego Dominus diligens iudicium,odio habens rapinam et iniquitatem;et dabo opus eorum in veritateet foedus perpetuum feriam eis.
ISA|61|9|Et scietur in gentibus semen eorum,et germen eorum in medio populorum;omnes, qui viderint eos, cognoscent illos,quia isti sunt semen, cui benedixit Dominus.
ISA|61|10|Gaudens gaudebo in Domino,et exsultabit anima mea in Deo meo,quia induit me vestimentis salutiset indumento iustitiae circumdedit me,quasi sponsum decoratum coronaet quasi sponsam ornatam monilibus suis.
ISA|61|11|Sicut enim terra profert germen suum,et sicut hortus semen suum germinat,sic Dominus Deus germinabit iustitiamet laudem coram universis gentibus.
ISA|62|1|Propter Sion non taceboet propter Ierusalem nonquiescam,donec egrediatur ut splendor iustitia eius,et salus eius ut lampas accendatur.
ISA|62|2|Et videbunt gentes iustitiam tuam,et cuncti reges gloriam tuam;et vocaberis nomine novo,quod os Domini nominabit.
ISA|62|3|Et eris corona gloriae in manu Domini,et diadema regni in manu Dei tui.
ISA|62|4|Non vocaberis ultra Derelicta,et terra tua non vocabitur amplius Desolata;sed vocaberis Beneplacitum meum in ea,et terra tua Nupta,quia complacuit Domino in te,et terra tua erit nupta.
ISA|62|5|Nam ut iuvenis uxorem ducit virginem,ita ducent te filii tui;ut gaudet sponsus super sponsam,ita gaudebit super te Deus tuus.
ISA|62|6|Super muros tuos, Ierusalem, constitui custodes;tota die et tota nocte, in perpetuo non tacebunt.Qui commonetis Dominum, ne taceatis
ISA|62|7|et ne detis silentium ei,donec stabiliat et donec ponat Ierusalemlaudem in terra.
ISA|62|8|Iuravit Dominus in dextera suaet in brachio fortitudinis suae: Non dabo triticum tuum ultracibum inimicis tuis,neque bibent filii alienivinum tuum, in quo laborasti.
ISA|62|9|Quia, qui collegerint illud, comedentet laudabunt Dominum;et, qui vindemiam fecerint,illud bibent in atriis sanctuarii mei.
ISA|62|10|Transite, transite per portas,parate viam populo.Sternite, sternite semitam, eligite lapides,elevate signum ad populos ".
ISA|62|11|Ecce Dominus auditum fecit in extremis terrae: Dicite filiae Sion:Ecce salus tua venit,ecce merces eius cum eo,et praemium eius coram illo.
ISA|62|12|Et vocabunt eos Populus sanctus,Redempti a Domino;tu autem vocaberis Quaesita,Civitas non derelicta ".
ISA|63|1|" Quis est iste, qui venit de Edom,tinctis vestibus de Bosra?Iste formosus in stola sua,gradiens in multitudine fortitudinis suae ". Sum ego, qui loquor iustitiam,potens ad salvandum ".
ISA|63|2|" Quare ergo rubrum est indumentum tuum,et vestimenta tua sicut calcantis in torculari? ".
ISA|63|3|" Torcular calcavi solus,et de gentibus non erat vir mecum;calcavi eos in furore meoet conculcavi eos in ira mea.Et aspersus est sanguis eorum super vestimenta mea,et omnia indumenta mea inquinavi.
ISA|63|4|Dies enim ultionis in corde meo,annus redemptionis meae venit.
ISA|63|5|Circumspexi, et non erat auxiliator,miratus sum, et non fuit qui adiuvaret;et salvavit mihi brachium meum,et indignatio mea ipsa auxiliata est mihi.
ISA|63|6|Et conculcavi populos in furore meoet contrivi eos in indignatione meaet effudi in terram sanguinem eorum ".
ISA|63|7|Miserationum Domini recordabor,laudum Dominisuper omnibus, quae reddidit nobis Dominus,et super multitudinem bonorum domui Israel,quae largitus est eis secundum misericordias suaset secundum multitudinem miserationum suarum.
ISA|63|8|Et dixit: " Verumtamen populus meus est,filii, qui non deludent ";et factus est eis salvator.
ISA|63|9|In omni tribulatione eorum non legatus neque angelus,sed ipse salvavit eos.In dilectione sua et in indulgentia suaipse redemit eoset sustulit eos et portavit eoscunctis diebus saeculi.
ISA|63|10|Ipsi autem ad iracundiam provocaveruntet afflixerunt spiritum sanctitatis eius;et conversus est eis in inimicumet ipse debellavit eos.
ISA|63|11|Et recordatus est dierum antiquorum,Moysi et populi sui.Ubi est qui eduxit eos de maricum pastore gregis sui?Ubi est qui posuit in medio eiusspiritum sanctitatis suae?
ISA|63|12|Qui adduxit ad dexteram Moysibrachium maiestatis suae,qui scidit aquas ante eos,ut faceret sibi nomen sempiternum,
ISA|63|13|qui deduxit eos per abyssosquasi equum per desertum, et non impingebant?
ISA|63|14|Sicut armentum, quod descendit per vallem,spiritus Domini fecit eos quiescere;sic conduxisti populum tuum,ut faceres tibi nomen gloriae.
ISA|63|15|Attende de caelo et videde habitaculo sancto tuo et gloriae tuae;ubi est zelus tuus et fortitudo tua?Commotio viscerum tuorum et misericordiae tuaesuper me continuerunt se.
ISA|63|16|Tu enim pater noster.Abraham enim nescit nos,et Israel ignorat nos;tu, Domine, pater noster,redemptor noster: a saeculo nomen tuum.
ISA|63|17|Quare errare nos fecisti, Domine, de viis tuis,indurasti cor nostrum, ne timeremus te?Convertere propter servos tuos,tribus hereditatis tuae.
ISA|63|18|Brevi tempore hereditaverunt populum sanctum tuum,hostes nostri conculcaverunt sanctuarium tuum.
ISA|63|19|Facti sumus a saeculo,cum non dominareris nostri,neque invocaretur nomen tuum super nos.Utinam dirumperes caelos et descenderes!A facie tua montes defluerent.
ISA|64|1|Sicut ignis succendit sarmenta,aquam ebullire facit ignis,ut notum facias nomen tuum inimicis tuis,a facie tua gentes turbentur,
ISA|64|2|cum feceris mirabilia,quae non sperabamus.Descendisti, et a facie tua montes defluxerunt.
ISA|64|3|A saeculo non audierunt, neque aures perceperunt;oculus non vidit Deum, absque te,qui operaretur pro sperantibus in eum.
ISA|64|4|Occurris laetanti, facienti iustitiamet his, qui in viis tuis recordantur tui.Ecce tu iratus es, et peccavimus;in ipsis a saeculo nos salvabimur.
ISA|64|5|Et facti sumus ut immundus omnes nos,et quasi pannus inquinatus universae iustitiae nostrae;et marcuimus quasi folium universi,et iniquitates nostrae quasi ventus abstulerunt nos.
ISA|64|6|Non est qui invocet nomen tuum,qui consurgat et adhaereat tibi,quia abscondisti faciem tuam a nobiset dissolvisti nos in manu iniquitatis nostrae.
ISA|64|7|Et nunc, Domine, pater noster es tu,nos vero lutum; et fictor noster tu,et opera manuum tuarum omnes nos.
ISA|64|8|Ne irascaris, Domine, nimiset ne ultra memineris iniquitatis;ecce, respice: populus tuus omnes nos.
ISA|64|9|Urbes sanctitatis tuae factae sunt in desertum,Sion deserta facta est,Ierusalem desolata est.
ISA|64|10|Domus sanctitatis nostrae et gloriae nostrae,ubi laudaverunt te patres nostri,facta est in exustionem ignis,et omnia desiderabilia nostra versa sunt in ruinas.
ISA|64|11|Numquid super his continebis te, Domine,tacebis et affliges nos vehementer?
ISA|65|1|" Quaesitus sum ab his, qui non consulebant me,inventus sum ab his, qui non quaerebant me.Dixi: "Ecce ego, ecce ego!"ad gentem, quae non invocabat nomen meum.
ISA|65|2|Expandi manus meas tota diead populum rebellem,qui graditur in via non bonapost cogitationes suas;
ISA|65|3|populus, qui ad iracundiam provocat meante faciem meam semper,qui immolant in hortiset sacrificant super lateres,
ISA|65|4|qui morantur in sepulcriset in locis occultis pernoctant,qui comedunt carnem suillamet ius abominabile in vasis eorum,
ISA|65|5|qui dicunt: "Recede!Non appropinques mihi, quia sanctificarem te".Isti fumus sunt in naribus meis,ignis ardens tota die.
ISA|65|6|Ecce scriptum est coram me;non tacebo, sed retribuam,et retribuam in sinum eorum
ISA|65|7|iniquitates vestras et iniquitates patrum vestrorumsimul, dicit Dominus,qui sacrificaverunt super monteset super colles exprobraverunt mihi;et remetiar opus eorum primoin sinu eorum ".
ISA|65|8|Haec dicit Dominus: Quomodo si inveniatur mustum in botroet dicatur: "Ne dissipes illud,quoniam benedictio est in eo",sic faciam propter servos meos,ut non disperdam totum.
ISA|65|9|Et educam de Iacob semenet de Iuda possidentem montes meos;et hereditabunt terram electi mei,et servi mei habitabunt ibi.
ISA|65|10|Et erit Saron in pascua gregum,et vallis Achor in cubile armentorumpopulo meo, qui quaesierunt me.
ISA|65|11|Vos autem, qui derelinquitis Dominum,qui obliviscimini montem sanctum meum,qui ponitis Gad mensamet amphoram impletis Meni,
ISA|65|12|numerabo vos in gladio,et omnes in caede corruetis;pro eo quod vocavi, et non respondistis,locutus sum, et non audistis,sed fecistis malum in oculis meiset, quod displicet mihi, elegistis ".
ISA|65|13|Propter hoc haec dicit Dominus Deus: Ecce servi mei comedent,et vos esurietis;ecce servi mei bibent,et vos sitietis;ecce servi mei laetabuntur,et vos confundemini;
ISA|65|14|ecce servi mei laudabunt in exsultatione cordis,et vos clamabitis prae dolore cordiset prae contritione spiritus ululabitis.
ISA|65|15|Et relinquetis nomen vestrumin iuramentum electis meis:Interficiat te Dominus Deus";et servos suos vocabit nomine alio.
ISA|65|16|Quicumque benedicit sibi in terra,benedicet sibi in Deo Amen;et, quicumque iurat in terra,iurabit in Deo Amen;quia oblivioni tradentur angustiae priores,et quia abscondentur ab oculis meis.
ISA|65|17|Ecce enim ego creocaelos novos et terram novam,et non erunt in memoria prioraet non ascendent super cor.
ISA|65|18|Sed gaudebunt et exsultabunt usque in sempiternumin his, quae ego creo,quia ecce ego creo Ierusalem exsultationemet populum eius gaudium.
ISA|65|19|Et exsultabo in Ierusalemet gaudebo in populo meo,et non audietur in ea ultravox fletus et vox clamoris.
ISA|65|20|Non erit ibi amplius infans dierumet senex, qui non impleat dies suos.Quoniam puer erit,qui centenarius moriatur;et, qui non attingat centum annos,maledictus erit.
ISA|65|21|Et aedificabunt domos et habitabuntet plantabunt vineas et comedent fructus earum.
ISA|65|22|Non aedificabunt, ut alius habitet,non plantabunt, ut alius comedat:secundum enim dies ligni erunt dies populi mei,et operibus manuum suarum diu fruentur electi mei.
ISA|65|23|Non laborabunt frustraneque generabunt in interitum repentinum,quia semen benedictorum erunt Domini,et nepotes eorum cum eis.
ISA|65|24|Eritque: antequam clament, ego respondebo;adhuc illis loquentibus, ego exaudiam.
ISA|65|25|Lupus et agnus pascentur simul,et leo sicut bos comedet paleas,et serpenti pulvis panis eius.Non nocebunt neque occidentin omni monte sancto meo ",dicit Dominus.
ISA|66|1|Haec dicit Dominus: Caelum thronus meus,terra autem scabellum pedum meorum.Quae ista domus, quam aedificabitis mihi,et quis iste locus quietis meae?
ISA|66|2|Omnia haec manus mea fecit,et mea sunt universa ista,dicit Dominus.Ad hunc autem respiciam,ad pauperculum et contritum spirituet trementem sermones meos.
ISA|66|3|Qui immolat bovem, interficit virum;qui sacrificat ovem, excerebrat canem;qui offert oblationem, idemque sanguinem suillum;qui adolet incensum, benedicit idolo.Sicut isti elegerunt vias suas,et in abominationibus suis anima eorum delectatur,
ISA|66|4|sic ego eligam malam sortem eorumet, quae timebant, adducam eis;quia vocavi, et non erat qui responderet,locutus sum, et non audieruntfeceruntque malum in oculis meiset, quod displicet mihi, elegerunt ".
ISA|66|5|Audite verbum Domini,qui tremitis ad verbum eius.Dixerunt fratres vestri odientes voset abicientes vos propter nomen meum: Gloriam suam manifestet Dominus,ut videamus laetitiam vestram";ipsi autem confundentur.
ISA|66|6|Vox clamoris de civitate,vox de templo,vox Dominireddentis retributionem inimicis suis.
ISA|66|7|Antequam parturiret, peperit;antequam veniret partus eius, peperit masculum.
ISA|66|8|Quis audivit umquam tale?Et quis vidit huic simile?Numquid oritur terra in die una,aut parietur gens in momento?Quia parturivit, iam peperit Sion filios suos.
ISA|66|9|" Numquid aperiam uterum et parere non faciam? ",dicit Dominus. Aut ego, qui parere facio, uterum claudam? ",ait Deus tuus.
ISA|66|10|Laetamini cum Ierusalem et exsultate in ea,omnes, qui diligitis eam;gaudete cum ea gaudio,universi, qui lugebatis super eam,
ISA|66|11|ut sugatis et repleaminiab ubere consolationis eius,ut mulgeatis et deliciis affluatisex uberibus gloriae eius.
ISA|66|12|Quia haec dicit Dominus: Ecce ego dirigam ad eam quasi fluvium pacemet quasi torrentem inundantem gloriam gentium.Sugetis, in ulnis portabimini,et super genua blandientur vobis.
ISA|66|13|Quomodo si quem mater consolatur,ita ego consolabor vos;et in Ierusalem consolabimini.
ISA|66|14|Videbitis, et gaudebit cor vestrum,et ossa vestra quasi herba germinabunt,et manifestabitur manus Domini in servis eius,et indignabitur inimicis suis.
ISA|66|15|Quia ecce Dominus in igne veniet,et quasi turbo quadrigae eius,reddere in indignatione furorem suumet increpationem suam in flamma ignis;
ISA|66|16|quia in igne Dominus diiudicabitet in gladio suo omnem carnem,et multiplicabuntur interfecti a Domino.
ISA|66|17|Qui sanctificantur et purificantur, ut ingredianturin hortos post aliquem stantem in medio,qui comedunt carnem suillamet abominationem et murem,simul consumentur,dicit Dominus.
ISA|66|18|Ego autem cognoscens opera eorum et cogitationes eorum veniam, ut congregem omnes gentes et linguas; et venient et videbunt gloriam meam.
ISA|66|19|Et ponam in eis signum et mittam ex eis, qui salvati fuerint, ad gentes in Tharsis, Phut, Lud, Mosoch, Ros, Thubal et Iavan, ad insulas longinquas, ad eos, qui non audierunt de me et non viderunt gloriam meam, et annuntiabunt gloriam meam gentibus;
ISA|66|20|et adducent omnes fratres vestros de cunctis gentibus oblationem Domino, in equis et in quadrigis et in lecticis et in mulis et in dromedariis, ad montem sanctum meum Ierusalem, dicit Dominus: quomodo si inferant filii Israel oblationem in vase mundo in domum Domini.
ISA|66|21|Et assumam ex eis in sacerdotes et Levitas, dicit Dominus.
ISA|66|22|Quia sicut caeli noviet terra nova, quae ego faciam,stabunt coram me,dicit Dominus,sic stabit semen vestrum et nomen vestrum.
ISA|66|23|Et erit: unoquoque novilunioet quovis sabbatoveniet omnis caro, ut adoret coram facie mea,dicit Dominus.
ISA|66|24|Et egredientur et videbunt cadavera virorum,qui praevaricati sunt in me;nam vermis eorum non morietur,et ignis eorum non exstinguetur,et erunt abominationi omni carni ".
JER|1|1|Verba Ieremiae filii Helciae de sacerdotibus, qui fuerunt in Anathoth in terra Beniamin.
JER|1|2|Quod factum est verbum Domini ad eum in diebus Iosiae filii Amon regis Iudae, in tertio decimo anno regni eius.
JER|1|3|Et factum est in diebus Ioachim filii Iosiae regis Iudae, usque ad consummationem undecimi anni Sedeciae filii Iosiae regis Iudae, usque ad transmigrationem Ierusalem in mense quinto.
JER|1|4|Et factum est verbum Domini ad me dicens:
JER|1|5|" Priusquam te formarem in utero, novi teet, antequam exires de vulva, sanctificavi teet prophetam gentibus dedi te ".
JER|1|6|Et dixi: " Heu, Domine Deus! Ecce nescio loqui, quia puer ego sum ".
JER|1|7|Et dixit Dominus ad me: " Noli dicere: "Puer sum",quoniam, ad quoscumque mittam te, ibiset universa, quaecumque mandavero tibi, loqueris.
JER|1|8|Ne timeas a facie eorum,quia tecum ego sum, ut eruam te ",dicit Dominus.
JER|1|9|Et misit Dominus manum suam et tetigit os meum; et dixit Dominus ad me: Ecce dedi verba mea in ore tuo;
JER|1|10|ecce constitui te hodie super gentes et super regna,ut evellas et destruaset disperdas et dissipeset aedifices et plantes ".
JER|1|11|Et factum est verbum Domini ad me dicens: " Quid tu vides, Ieremia? ". Et dixi: " Virgam amygdali vigilantis ego video ".
JER|1|12|Et dixit Dominus ad me: "Bene vidisti, quia vigilo ego super verbo meo, ut faciam illud ".
JER|1|13|Et factum est verbum Domini secundo ad me dicens: " Quid tu vides? ". Et dixi: " Ollam succensam ego video; et facies eius a facie aquilonis ".
JER|1|14|Et dixit Dominus ad me: Ab aquilone pandetur malumsuper omnes habitatores terrae;
JER|1|15|quia ecce ego convocaboomnia regna aquilonis,ait Dominus,et venient et ponent unusquisque solium suumin introitu portarum Ierusalemet contra omnes muros eius in circuituet contra universas urbes Iudae;
JER|1|16|et loquar iudicia mea cum eissuper omnem malitiam eorum,qui dereliquerunt meet incensum obtulerunt diis alieniset adoraverunt opus manuum suarum.
JER|1|17|Tu ergo accinge lumbos tuoset surge et loquere ad eos omnia,quae ego praecipio tibi;ne timeas a facie eorum,alioquin timere te faciam vultum eorum.
JER|1|18|Ego quippe dedi te hodiein civitatem munitamet in columnam ferreamet in murum aereumcontra omnem terramregibus Iudae, principibus eiuset sacerdotibus et populo terrae;
JER|1|19|et bellabunt adversum te et non praevalebunt,quia tecum ego sum,ait Dominus,ut eripiam te ".
JER|2|1|Et factum est verbum Domini ad me dicens:
JER|2|2|" Vade et clama in auribus Ierusalem dicens:Haec dicit Dominus:Recordatus sum tui, caritatis adulescentiae tuaeet amoris desponsationis tuae,quando secuta es me in deserto,in terra, quae non seminatur.
JER|2|3|Sanctus Domino Israel,primitiae frugum eius;omnes, qui devorabant eum, delinquebant;mala veniebant super eos,dicit Dominus.
JER|2|4|Audite verbum Domini, domus Iacobet omnes cognationes domus Israel.
JER|2|5|Haec dicit Dominus:Quid invenerunt patres vestri in me iniquitatis,quia elongaverunt a meet ambulaverunt post vanitatemet vani facti sunt?
JER|2|6|Et non dixerunt: "Ubi est Dominus,qui ascendere nos fecit de terra Aegypti,qui traduxit nos per desertum,per terram inhabitabilem et inviam,per terram sitis et caliginis,per terram, in qua non ambulavit vir,neque habitavit homo?".
JER|2|7|Et induxi vos in terram hortorum,ut comederetis fructum eius et optima illius;et ingressi contaminastis terram meamet hereditatem meam posuistis in abominationem.
JER|2|8|Sacerdotes non dixerunt:Ubi est Dominus?".Et tractantes legem nescierunt me,et pastores praevaricati sunt in me,et prophetae prophetaverunt in Baalet, quae nihil prosunt, secuti sunt.
JER|2|9|Propterea adhuc iudicio contendam vobiscum,ait Dominus,et cum filiis filiorum vestrorum disceptabo.
JER|2|10|En transite ad insulas Cetthim et videteet in Cedar mittite et considerate vehementeret videte, si factum est huiuscemodi:
JER|2|11|si mutavit gens deos,et certe ipsi non sunt dii;populus vero meus mutavit gloriam suamin id, quod nihil prodest.
JER|2|12|Obstupescite, caeli, super hocet inhorrescite supra modum,dicit Dominus.
JER|2|13|Duo enim mala fecit populus meus:me dereliquerunt fontem aquae vivae,ut foderent sibi cisternas,cisternas dissipatas,quae continere non valent aquas.
JER|2|14|Numquid servus est Israelaut vernaculus?Quare ergo factus est in praedam?Super eum rugierunt leones
JER|2|15|et dederunt vocem suam;posuerunt terram eius in solitudinem:civitates eius exustae sunt,et non est qui habitet in eis.
JER|2|16|Filii quoque Mempheos et Taphnesdecalvabunt tibi verticem.
JER|2|17|Numquid non istud factum est tibi,quia dereliquisti Dominum Deum tuumeo tempore, quo ducebat te per viam?
JER|2|18|Et nunc quid tibi vis in via Aegypti,ut bibas aquam Nili?Et quid tibi cum via Assyriorum,ut bibas aquam Fluminis?
JER|2|19|Arguet te malitia tua,et aversio tua increpabit te;scito et vide quia malum et amarum estreliquisse te Dominum Deum tuum et non esse timorem mei apud te,dicit Dominus, Deus exercituum.
JER|2|20|A saeculo confregisti iugum tuum,rupisti vincula tuaet dixisti: "Non serviam".In omni enim colle sublimiet sub omni ligno frondosotu prosternebaris meretrix.
JER|2|21|Ego autem plantavi te vineam electam,omne semen verum;quomodo ergo conversa esin palmites vineae alienae?
JER|2|22|Si laveris te nitroet multiplicaveris tibi herbam fullonum,maculata es in iniquitate tua coram me,dicit Dominus Deus.
JER|2|23|Quomodo dicis: "Non sum polluta,post Baalim non ambulavi"?Vide viam tuam in convalle,scito quid feceris:camelus levis contorquens vias suas.
JER|2|24|Onager assuetus in solitudinein desiderio animae suae attrahit aerem;libidinem eius quis avertet?Omnes, qui quaerunt eam, non deficient,in menstruis eius invenient eam.
JER|2|25|Prohibe pedem tuum a nuditateet guttur tuum a siti.Et dixisti: "Vanum est, nequaquam;adamavi quippe alienoset post eos ambulabo".
JER|2|26|Quomodo confunditur fur, quando deprehenditur,sic confusi sunt domus Israel,ipsi et reges eorum, principeset sacerdotes et prophetae eorum
JER|2|27|dicentes ligno: "Pater meus es tu" et lapidi: "Tu me genuisti".Verterunt ad me tergum et non faciem,sed in tempore afflictionis suae dicent:Surge et libera nos!".
JER|2|28|Ubi sunt dii tui, quos fecisti tibi?Surgant et liberent te in tempore afflictionis tuae;secundum numerum quippe civitatum tuarumfacti sunt dii tui, Iuda.
JER|2|29|Quid vultis mecum iudicio contendere?Omnes praevaricati estis in me,dicit Dominus.
JER|2|30|Frustra percussi filios vestros:disciplinam non receperunt.Devoravit gladius vester prophetas vestros:quasi leo vastator.
JER|2|31|O generatio, vos videte verbum Domini:numquid solitudo factus sum Israeliaut terra tenebrarum?Quare ergo dixit populus meus: "Recessimus,non veniemus ultra ad te"?
JER|2|32|Numquid obliviscitur virgo ornamenti sui,sponsa fasciae pectoralis suae?Populus vero meus oblitus est meidiebus innumeris.
JER|2|33|Quam bene paras viam tuamad quaerendum amorem!Et insuper in malumdocuisti vias tuas,
JER|2|34|et in fimbriis tuis inventus estsanguis animarum pauperum innocentium:non effringentes invenisti eos;sed in omnibus his
JER|2|35|dixisti: "Innocens ego sum,propterea aversus est furor eius a me".Ecce ego iudicio contendam tecum, eo quod dixeris: "Non peccavi".
JER|2|36|Quam leviter mutas vias tuas!Et ab Aegypto confunderis,sicut confusa es ab Assyria.
JER|2|37|Nam et ab ista egredieris,et manus tuae erunt super caput tuum,quoniam obtrivit Dominus illos, quibus confisus es,et nihil habebis prosperum in eis.
JER|3|1|Si dimiserit vir uxorem suam,et recedens ab eoduxerit virum alterum,numquid revertetur ad eam ultra?Numquid non pollutaet contaminata est terra illa?Tu autem fornicata es cum amatoribus multiset reverteris ad me?,dicit Dominus.
JER|3|2|Leva oculos tuos ad colles et vide,ubi non prostrata sis.In viis sedebas exspectans eosquasi Arabs in solitudine;et polluisti terramin fornicationibus tuis et in malitia tua.
JER|3|3|Quam ob rem prohibitae sunt stillae pluviarum,et serotinus imber non fuit.Frons mulieris meretricis facta est tibi;noluisti erubescere.
JER|3|4|Nonne amodo vocas me: "Pater meus,dux adulescentiae meae tu es!
JER|3|5|Numquid irascetur in perpetuumaut perseverabit in finem?".Ecce locuta eset fecisti mala et praevaluisti ".
JER|3|6|Et dixit Dominus ad me in diebus Iosiae regis: " Numquid vidisti, quae fecerit aversatrix Israel? Abiit sibimet super omnem montem excelsum et sub omni ligno frondoso et fornicata est ibi.
JER|3|7|Et dixi: "Cum fecerit haec omnia, ad me revertetur"; et non est reversa. Et vidit praevaricatrix soror eius, Iuda;
JER|3|8|et vidit quia pro eo quod moechata esset aversatrix Israel, dimisissem eam et dedissem ei libellum repudii, et non timuit praevaricatrix Iuda, soror eius, sed abiit et fornicata est etiam ipsa;
JER|3|9|et facilitate fornicationis suae contaminavit terram et moechata est cum lapide et ligno.
JER|3|10|Sed in omnibus his non est reversa ad me praevaricatrix soror eius Iuda in toto corde suo sed in mendacio ", ait Dominus.
JER|3|11|Et dixit Dominus ad me: " Iustificavit animam suam aversatrix Israel comparatione praevaricatricis Iudae.
JER|3|12|Vade et clama sermones istos contra aquilonem et dices:Revertere, aversatrix Israel,ait Dominus,et non avertam faciem meam a vobis,quia pius ego sum,dicit Dominus,et non irascar in perpetuum.
JER|3|13|Verumtamen scito iniquitatem tuam,quia in Dominum Deum tuum praevaricata eset dispersisti vias tuas alienissub omni ligno frondoso;et vocem meam non audistis,ait Dominus.
JER|3|14|Convertimini, filii, qui aversi estis a me, dicit Dominus, quia ego Dominus vester sum; et assumam vos unum de civitate et duos de cognatione et introducam vos in Sion;
JER|3|15|et dabo vobis pastores iuxta cor meum, et pascent vos scientia et doctrina.
JER|3|16|Cumque multiplicati fueritis et creveritis in terra in diebus illis, ait Dominus, non dicent ultra: "Arca testamenti Domini", neque ascendet super cor, neque recordabuntur illius, nec requiretur, nec fiet ultra.
JER|3|17|In tempore illo vocabunt Ierusalem Solium Domini, et congregabuntur ad eam omnes gentes in nomine Domini in Ierusalem; et non ambulabunt ultra post pravitatem cordis sui pessimi.
JER|3|18|In diebus illis ibit domus Iudae ad domum Israel, et venient simul de terra aquilonis ad terram, quam dedi in hereditatem patribus vestris.
JER|3|19|Ego autem dixi:Quomodo ponam te in filiiset tribuam tibi terram desiderabilem,hereditatem praeclarissimam inter gentes?Et dixi: Patrem vocabitis meet post me ingredi non cessabitis.
JER|3|20|Sed, quomodo contemnit mulier amatorem suum,sic contempsistis me, domus Israel ",dicit Dominus.
JER|3|21|Vox in collibus audita est,ploratus et supplicatio filiorum Israel,quoniam iniquam fecerunt viam suam,obliti sunt Domini Dei sui.
JER|3|22|" Convertimini, filii, qui aversi estis a me,et sanabo aversiones vestras ". Ecce nos venimus ad te;tu enim es Dominus Deus noster.
JER|3|23|Vere mendaces erant colleset tumultus montium;vere in Domino Deo nostrosalus Israel.
JER|3|24|Confusio comedit laborem patrum nostrorumab adulescentia nostra,greges eorum et armenta eorum,filios eorum et filias eorum.
JER|3|25|Dormiemus in confusione nostra,et operiet nos ignominia nostra,quoniam Domino Deo nostro peccavimusnos et patres nostriab adulescentia nostra usque ad hanc diemet non audivimus vocem Domini Dei nostri ".
JER|4|1|" Si converteris, Israel,ait Dominus,ad me convertere;si abstuleris abominationes tuas a facie mea,non effugies.
JER|4|2|Et iurabis: "Vivit Dominus!"in veritate et in iudicio et in iustitia,et benedicentur in ipso genteset in ipso gloriabuntur.
JER|4|3|Haec enim dicit Dominusviro Iudae et Ierusalem:Novate vobis novaleet nolite serere super spinas.
JER|4|4|Circumcidimini Dominoet auferte praeputia cordium vestrorum,viri Iudae et habitatores Ierusalem,ne forte egrediatur ut ignis indignatio meaet succendatur, et non sit qui exstinguat,propter malitiam operum vestrorum.
JER|4|5|Annuntiate in Iudaet in Ierusalem auditum facite;et loquimini et canite tuba in terra,clamate fortiter et dicite:Congregamini, et ingrediamur civitates munitas".
JER|4|6|Levate signum in Sion,fugite, nolite stare,quia malum ego adduco ab aquiloneet contritionem magnam.
JER|4|7|Ascendit leo de cubili suo,et praedo gentium se levavit;egressus est de loco suo,ut ponat terram tuam in solitudinem:civitates tuae vastabuntur,remanentes absque habitatore.
JER|4|8|Super hoc accingite vos ciliciis,plangite et ululate,quia non est aversa ira furoris Domini a nobis.
JER|4|9|Et erit in die illa,dicit Dominus,peribit cor regiset cor principum,et obstupescent sacerdotes,et prophetae consternabuntur ".
JER|4|10|Et dixi: " Heu, Domine Deus!Ergo decepisti populum istum et Ierusalemdicens: "Pax erit vobis";et ecce pervenit gladius usque ad animam ".
JER|4|11|In tempore illo dicetur populo huic et Ierusalem: Ventus urens collium, qui sunt in deserto,invadit filiam populi meinon ad ventilandum et ad purgandum.
JER|4|12|Ventus plenior his veniet mihi,nunc et ego loquar iudicia mea cum eis ".
JER|4|13|Ecce quasi nubes ascendet,et quasi tempestas currus eius;velociores aquilis equi illius.Vae nobis, quoniam vastati sumus!
JER|4|14|Lava a malitia cor tuum,Ierusalem, ut salva fias;usquequo morabuntur in tecogitationes iniquae?
JER|4|15|Vox enim annuntiantis a Danet notam facientis calamitatem de monte Ephraim.
JER|4|16|Nuntiate gentibus. Ecce adsunt!Auditum facite hoc super Ierusalem: Custodes venerunt de terra longinquaet dederunt super civitates Iudae vocem suam;
JER|4|17|quasi custodes agrorum facti sunt super eam in gyro,quia adversus me contumax erat ",dicit Dominus.
JER|4|18|Via tua et opera tuafecerunt haec tibi;ista malitia tua, quia amara,quia tetigit cor tuum.
JER|4|19|Viscera mea, viscera mea! Doleo.Parietes cordis mei!Turbatur in me cor meum:non tacebo,quoniam vocem bucinae audivit anima mea,clamorem proelii.
JER|4|20|Contritio super contritionem vocata est,quoniam vastata est omnis terra,repente vastata sunt tabernacula mea,subito tentoria mea.
JER|4|21|Usquequo videbo vexillum,audiam vocem bucinae?
JER|4|22|" Quia stultus populus meus:me non cognoverunt;filii insipientes sunt et vecordes:sapientes sunt, ut faciant mala,bene autem facere nesciunt ".
JER|4|23|Aspexi terram, et ecce vacua erat et deserta;et caelos, et non erat lux in eis.
JER|4|24|Aspexi montes, et ecce movebantur,et omnes colles conturbati sunt.
JER|4|25|Aspexi, et ecce non erat homo,et omne volatile caeli recesserat.
JER|4|26|Aspexi, et ecce hortus desertus,et omnes urbes eius destructae sunta facie Domini et a facie irae furoris eius.
JER|4|27|Haec enim dicit Dominus: Deserta erit omnis terra,sed tamen consummationem non faciam.
JER|4|28|Super hoc lugebit terra,et maerebunt caeli desuper,eo quod locutus sum,statui et non paenitet menec avertar ab eo ".
JER|4|29|A voce equitis et mittentis sagittamfugit omnis civitas;ingressi sunt silvas condensaset ascenderunt rupes;universae urbes derelictae sunt,et non habitat in eis homo.
JER|4|30|Tu autem, vastata, quid facies?Cum vestieris te coccino,cum ornata fueris monili aureo,et pinxeris stibio oculos tuos,frustra componeris;contempserunt te amatores tui,animam tuam quaerent.
JER|4|31|Vocem enim quasi parturientis audivi,angustias ut puerperae;vox filiae Sionintermorientis expandentisque manus suas: Vae mihi, quia defecit anima meapropter interfectores! ".
JER|5|1|Circuite vias Ierusalemet aspicite et considerateet quaerite in plateis eius,an inveniatis virum,an sit qui faciat iudicium et quaerentem fidem,et propitius ero ei.
JER|5|2|Quod si etiam " Vivit Dominus! " dixerint,certe falso iurabunt.
JER|5|3|Domine, nonne oculi tui respiciunt fidem?Percussisti eos, et non doluerunt,attrivisti eos, et renuerunt accipere disciplinam:induraverunt facies suas supra petram,noluerunt reverti.
JER|5|4|Ego autem dixi: " Ecce pauperes illi stulte agunt,quia ignorant viam Domini,iudicium Dei sui.
JER|5|5|Ibo igitur ad optimateset loquar eis;ipsi enim noverunt viam Domini,iudicium Dei sui ".Ecce hi simul confregerunt iugum, ruperunt vincula.
JER|5|6|Idcirco percussit eos leo de silva,lupus deserti vastabit eos,pardus vigilans super civitates eorum:omnis, qui egressus fuerit ex eis, lacerabitur,quia multiplicatae sunt praevaricationes eorum,confortatae sunt aversiones eorum.
JER|5|7|" Super quo propitius tibi esse potero?Filii tui dereliquerunt meet iuraverunt in his, qui non sunt dii;saturavi eos, et moechati suntet in domum meretricis gregatim confluebant.
JER|5|8|Equi impinguati et admissarii facti sunt:unusquisque ad uxorem proximi sui hinniebat.
JER|5|9|Numquid super his non visitabo,dicit Dominus,et in gente tali non ulciscetur anima mea?
JER|5|10|Ascendite muros eius et dissipate,consummationem autem nolite facere;auferte propagines eius,quia non sunt Domini.
JER|5|11|Praevaricatione enim praevaricata est in medomus Israel et domus Iudae ",ait Dominus.
JER|5|12|Negaverunt Dominumet dixerunt: "Non est ipse;neque veniet super nos malum,et gladium et famem non videbimus.
JER|5|13|Prophetae erunt in ventum,et responsum non est in eis.Haec ergo evenient illis ".
JER|5|14|Propterea haec dicit Dominus, Deus exercituum: Quia locuti estis verbum istud,ecce ego do verba mea in ore tuo in ignemet populum istum in ligna,et vorabit eos.
JER|5|15|Ecce ego adducam super vos gentem de longinquo,domus Israel,ait Dominus,gentem robustam,gentem antiquam,gentem, cuius ignorabis linguamnec intelleges quid loquatur.
JER|5|16|Pharetra eius quasi sepulcrum patensuniversi fortes.
JER|5|17|Et comedet segetes tuas et panem tuum,devorabit filios tuos et filias tuas,comedet gregem tuum et armenta tua,comedet vineam tuam et ficum tuam;et conteret urbes munitas tuas,in quibus tu habes fiduciam, gladio.
JER|5|18|Verumtamen et in diebus illis,ait Dominus,non faciam in vobis consummationem ".
JER|5|19|Quod si dixeritis: " Quare fecit nobis Dominus Deus noster haec omnia?, dices ad eos: " Sicut dereliquistis me et servistis diis alienis in terra vestra, sic servietis alienis in terra non vestra ".
JER|5|20|Annuntiate hoc domui Iacobet auditum facite in Iuda dicentes:
JER|5|21|" Audi, popule stulte, qui non habes cor,qui habentes oculos non vident,et aures et non audiunt.
JER|5|22|Numquid me non timebitis,ait Dominus,et a facie mea non trepidabitis?Qui posui arenam terminum mari, praeceptum sempiternum, quod non praeteribit;et commovebuntur et non poterunt,et intumescent fluctus eius, et non transibunt illud ".
JER|5|23|Populo autem huic factum est cor contumax et rebelle;recesserunt et abierunt
JER|5|24|et non dixerunt in corde suo: Metuamus Dominum Deum nostrum,qui dat nobis pluviamtemporaneam et serotinam in tempore suo,hebdomadas statutas messiscustodientem nobis ".
JER|5|25|Iniquitates vestrae declinaverunt haec,et peccata vestra prohibuerunt bonum a vobis,
JER|5|26|quia inventi sunt in populo meo impii,insidiantes quasi incurvati aucupes,laqueos ponentes ad capiendos viros.
JER|5|27|Sicut decipula plena avibus,sic domus eorum plenae dolo;ideo magnificati sunt et ditati,
JER|5|28|incrassati sunt et impinguati:et transgressi sunt terminos mali.Causam non iudicaverunt,causam pupilli, ut ipsi prospere agant,et iudicium pauperum non iudicaverunt.
JER|5|29|Numquid super his non visitabo,dicit Dominus,aut super gentem huiuscemodinon ulciscetur anima mea?
JER|5|30|Stupor et mirabiliafacta sunt in terra:
JER|5|31|prophetae prophetabant mendacium,et sacerdotes applaudebant manibus suis,et populus meus dilexit talia.Quid igitur facietis in novissimo eius?
JER|6|1|Fugite, filii Beniamin,de medio Ierusalem;et in Thecua clangite bucinaet super Bethcharem levate vexillum,quia malum visum est ab aquiloneet contritio magna.
JER|6|2|Speciosam et delicatam silere fecifiliam Sion.
JER|6|3|Ad eam venient pastores et greges eorum,figent in ea tentoria in circuitu;pascet unusquisque partem suam.
JER|6|4|" Sanctificate super eam bellum,consurgite, et ascendamus in meridie;vae nobis, quia declinavit dies,quia longiores factae sunt umbrae vesperi!
JER|6|5|Surgite, et ascendamus in nocteet dissipemus domos eius ".
JER|6|6|Quia haec dicit Dominus exercituum: Caedite lignum eiuset fundite circa Ierusalem aggerem;haec est civitas visitationis,omnis calumnia in medio eius.
JER|6|7|Sicut effluere facit cisterna aquam suam,sic illa effluere facit malitiam suam;violentia et vastitas auditur in ea,coram me semper afflictio et plaga.
JER|6|8|Erudire, Ierusalem,ne forte recedat anima mea a te,ne forte ponam te desertam,terram inhabitabilem ".
JER|6|9|Haec dicit Dominus exercituum: Usque ad racemum colligent quasi in vineareliquias Israel.Converte manum tuamquasi vindemiator ad palmites ".
JER|6|10|Cui loquar et quem contestabor, ut audiat?Ecce incircumcisae aures eorum,et audire non possunt;ecce verbum Domini factum est eis in opprobrium,et non suscipient illud.
JER|6|11|Idcirco furore Domini plenus sum,laboravi sustinens. Effunde super parvulum foriset super concilium iuvenum simul;etiam vir cum muliere capietur,senex cum pleno dierum.
JER|6|12|Et transibunt domus eorum ad alteros,agri et uxores pariter,quia extendam manum meamsuper habitantes terram ",dicit Dominus.
JER|6|13|A minore quippe usque ad maioremomnes avaritiae student,et a propheta usque ad sacerdotemcuncti faciunt dolum.
JER|6|14|Et curant contritionem populi mei in levitatedicentes: " Pax, pax "; et non est pax.
JER|6|15|Confusi sunt, quia abominationem fecerunt;quin potius confusione non sunt confusiet erubescere nescierunt. Quam ob rem cadent inter ruentes;tempore, quo visitavero eos, corruent ",dicit Dominus.
JER|6|16|Haec dicit Dominus: State super vias et videteet interrogate de semitis antiquis,quae sit via bona, et ambulate in eaet invenietis refrigerium animabus vestris ".Et dixerunt: " Non ambulabimus! ".
JER|6|17|Et constitui super vos speculatores: Audite vocem tubae ".Et dixerunt: " Non audiemus! ".
JER|6|18|Ideo audite, gentes,et cognosce, congregatio,quanta ego faciam eis.
JER|6|19|Audi terra: " Ecce ego adducam mala super populum istum,fructum cogitationum eorum,quia verba mea non audieruntet legem meam proiecerunt.
JER|6|20|Ut quid mihi tus, quod de Saba venit,et calamus suave olens de terra longinqua?Holocautomata vestra non sunt accepta,et victimae vestrae non placent mihi ".
JER|6|21|Propterea haec dicit Dominus: Ecce ego dabo in populum istum offendicula,et offendent in eis patres et filii simul,vicinus et proximus peribunt ".
JER|6|22|Haec dicit Dominus: Ecce populus venit de terra aquilonis,et gens magna consurget a finibus terrae;
JER|6|23|arcum et acinacem arripiet,crudelis est et non miserebitur;vox eorum quasi mare sonabit,et super equos ascendent,praeparati quasi vir ad proeliumadversum te, filia Sion ".
JER|6|24|" Audivimus famam eius;dissolutae sunt manus nostrae,tribulatio apprehendit nos,dolores ut parturientem ".
JER|6|25|Nolite exire ad agroset in via ne ambuletis,quoniam gladius inimici,pavor in circuitu.
JER|6|26|Filia populi mei, accingere cilicioet volutare in cinere,luctum unigeniti fac tibi,planctum amarum,quia repente veniet vastator super nos.
JER|6|27|Probatorem dedi te in populo meo;et scies et probabis viam eorum.
JER|6|28|Omnes isti principes rebelles,ambulantes fraudulenter.Aes et ferrum,omnia isti corrumpunt.
JER|6|29|Sufflavit sufflatorium in igne,consumptum est plumbum;frustra conflavit conflator,scoriae enim non sunt separatae.
JER|6|30|Argentum reprobum vocate eos,quia Dominus proiecit illos.
JER|7|1|Verbum, quod factum est ad Ieremiam a Domino dicens:
JER|7|2|" Sta in porta domus Domini et praedica ibi verbum istud et dic: Audite verbum Domini, omnis Iuda, qui ingredimini per portas has, ut adoretis Dominum.
JER|7|3|Haec dicit Dominus exercituum, Deus Israel: Bonas facite vias vestras et opera vestra, et habitare vos faciam in loco isto.
JER|7|4|Nolite confidere in verbis mendacii dicentes: "Templum Domini, templum Domini, templum Domini est".
JER|7|5|Quoniam, si bene direxeritis vias vestras et opera vestra, si feceritis iudicium inter virum et proximum eius,
JER|7|6|advenae et pupillo et viduae non feceritis calumniam nec sanguinem innocentem effuderitis in loco hoc et post deos alienos non ambulaveritis in malum vobismetipsis,
JER|7|7|habitare vos faciam in loco isto, in terra, quam dedi patribus vestris a saeculo usque in saeculum.
JER|7|8|Ecce vos confiditis vobis in sermonibus mendacii, qui non proderunt.
JER|7|9|Quid? Furari, occidere, adulterari, iurare mendaciter, incensum offerre Baal et ire post deos alienos, quos ignoratis;
JER|7|10|et venitis et statis coram me in domo hac, super quam invocatum est nomen meum, et dicitis: "Liberati sumus", eo quod faciatis omnes abominationes istas.
JER|7|11|Numquid spelunca latronum facta est domus ista, super quam invocatum est nomen meum in oculis vestris?Ecce, etiam ego vidi, dicit Dominus.
JER|7|12|Ite ad locum meum in Silo, ubi habitavit nomen meum a principio, et videte, quae fecerim ei propter malitiam populi mei Israel.
JER|7|13|Et nunc, quia fecistis omnia opera haec, dicit Dominus, et locutus sum ad vos mane consurgens et loquens, et non audistis, et vocavi vos, et non respondistis,
JER|7|14|faciam domui huic, super quam invocatum est nomen meum, et in qua vos habetis fiduciam, et loco, quem dedi vobis et patribus vestris, sicut feci Silo;
JER|7|15|et proiciam vos a facie mea, sicut proieci omnes fratres vestros, universum semen Ephraim.
JER|7|16|Tu ergo, noli orare pro populo hoc nec assumas pro eis deprecationem et orationem et non obsistas mihi, quia non exaudiam te.
JER|7|17|Nonne vides, quid isti faciant in civitatibus Iudae et in plateis Ierusalem?
JER|7|18|Filii colligunt ligna, et patres succendunt ignem, et mulieres commiscent farinam, ut faciant placentas reginae caeli et libent diis alienis, ut me ad iracundiam provocent.
JER|7|19|Numquid me ad iracundiam provocant, dicit Dominus, nonne semetipsos in confusionem vultus sui?
JER|7|20|Ideo haec dicit Dominus Deus: Ecce furor meus et indignatio mea effunditur super locum istum, super homines et super iumenta et super lignum regionis et super fruges terrae et succendetur et non exstinguetur.
JER|7|21|Haec dicit Dominus exercituum, Deus Israel: Holocautomata vestra addite victimis vestris et comedite carnes,
JER|7|22|quia non sum locutus cum patribus vestris et non praecepi eis in die, qua eduxi eos de terra Aegypti, de verbo holocautomatum et victimarum.
JER|7|23|Sed hoc verbum praecepi eis dicens: Audite vocem meam, et ero vobis Deus, et vos eritis mihi populus; et ambulate in omni via, quam mandaverim vobis, ut bene sit vobis.
JER|7|24|Et non audierunt nec inclinaverunt aurem suam, sed abierunt in voluntatibus et in pravitate cordis sui mali factique sunt retrorsum et non in ante
JER|7|25|a die, qua egressi sunt patres eorum de terra Aegypti, usque ad diem hanc. Et misi ad vos omnes servos meos prophetas, per diem consurgens diluculo et mittens;
JER|7|26|et non audierunt me nec inclinaverunt aurem suam, sed induraverunt cervicem suam et peius operati sunt quam patres eorum.
JER|7|27|Et loqueris ad eos omnia verba haec, et non audient te; et vocabis eos, et non respondebunt tibi;
JER|7|28|et dices ad eos: Haec est gens, quae non audivit vocem Domini Dei sui nec recepit disciplinam. Periit fides et ablata est de ore eorum.
JER|7|29|Tonde capillum tuum et proiceet sume in collibus planctum,quia sprevit Dominuset proiecit generationem furoris sui.
JER|7|30|Quia fecerunt filii Iudae malum in oculis meis, dicit Dominus; posuerunt abominationes suas in domo, super quam invocatum est nomen meum, ut polluerent eam;
JER|7|31|et aedificaverunt excelsa Topheth, quae est in valle Benennom, ut incenderent filios suos et filias suas igni: quae non praecepi nec cogitavi in corde meo.
JER|7|32|Ideo ecce dies venient, dicit Dominus, et non dicetur amplius Topheth et vallis Benennom sed vallis Interfectionis; et sepelient in Topheth, eo quod non sit locus.
JER|7|33|Et erit morticinum populi huius in cibum volucribus caeli et bestiis terrae, et non erit qui abigat.
JER|7|34|Et quiescere faciam de urbibus Iudae et de plateis Ierusalem vocem gaudii et vocem laetitiae, vocem sponsi et vocem sponsae: in desolationem enim erit terra ".
JER|8|1|" In illo tempore, ait Dominus, eicient ossa regum Iudae et ossa principum eius et ossa sacerdotum et ossa prophetarum et ossa eorum, qui habitaverunt Ierusalem de sepulcris suis;
JER|8|2|et expandent ea ad solem et lunam et omnem militiam caeli, quae dilexerunt et quibus servierunt et post quae ambulaverunt et quae quaesierunt et adoraverunt; non colligentur et non sepelientur: in sterquilinium super faciem terrae erunt.
JER|8|3|Et eligent magis mortem quam vitam omnes, qui residui fuerint de cognatione hac pessima in universis locis, ad quae eiecero eos, dicit Dominus exercituum.
JER|8|4|Et dices ad eos: Haec dicit Dominus:Numquid, qui cadit, non resurget, et, qui aversus est, non revertetur?
JER|8|5|Quare ergo aversus est populus iste,Ierusalem aversione perpetua?Apprehenderunt mendaciumet noluerunt reverti.
JER|8|6|Attendi et auscultavi:nemo, quod bonum est, loquitur,nullus est, qui agat paenitentiamsuper malitia sua dicens:Quid feci?".Omnes conversi sunt ad cursum suum,quasi equus impetu vadens in proelio.
JER|8|7|Etiam ciconia in caelonovit tempus suum;turtur et hirundo et turduscustodierunt tempus adventus sui;populus autem meus non novitiudicium Domini.
JER|8|8|Quomodo dicitis: "Sapientes nos sumus,et lex Domini nobiscum est"?Vere mendacium operatus eststilus mendax scribarum.
JER|8|9|Confusi sunt sapientes,perterriti et capti sunt;verbum enim Domini proiecerunt,et sapientia nulla est in eis.
JER|8|10|Propterea dabo mulieres eorum exteris,agros eorum expugnatoribus,quia a minimo usque ad maximumomnes avaritiam sequuntur,a propheta usque ad sacerdotemcuncti faciunt mendacium.
JER|8|11|Et sanant contritionemfiliae populi mei in levitatedicentes "Pax, pax", cum non sit pax.
JER|8|12|Confusi sunt, quia abominationem fecerunt;quin immo confusione non sunt confusiet erubescere nescierunt,idcirco cadent inter corruentes,in tempore visitationis suae corruent,dicit Dominus.
JER|8|13|Congregans congregabo eos,ait Dominus;non est uva in vitibus,et non sunt ficus in ficulnea,folium defluxit,et dabo eis gradientes super eos.
JER|8|14|"Quare sedemus?Convenite, et ingrediamur civitates munitaset pereamus ibi,quia Dominus Deus noster tradidit nos in interitumet potum dedit nobis aquam fellis;peccavimus enim Domino.
JER|8|15|Exspectavimus pacem, et non est bonum,tempus medelae, et ecce formido".
JER|8|16|A Dan auditus est fremitus equorum eius,a voce hinnituum fortium equorum eiuscommota est omnis terra;et venient et devorabunt terram et plenitudinem eius,urbem et habitatores eius.
JER|8|17|Quia ecce ego mittam vobisserpentes regulos,quibus non est incantatio,et mordebunt vos ",ait Dominus.
JER|8|18|Hilaritas mea facta est dolor in me,cor meum maerens.
JER|8|19|Ecce vox clamoris filiae populi meide terra longinqua: Numquid Dominus non est in Sion?Aut rex eius non est in ea? ". Quare ergo me ad iracundiam concitaverunt in sculptilibus suiset in vanitatibus alienis? ".
JER|8|20|" Transiit messis, finita est aestas,et nos salvati non sumus ".
JER|8|21|Super contritione filiae populi meicontritus sum et contristatus;stupor obtinuit me.
JER|8|22|Numquid resina non est in Galaad?Aut medicus non est ibi?Quare enim non est obductacicatrix filiae populi mei?
JER|8|23|Quis dabit capiti meo aquamet oculis meis fontem lacrimarum,et plorabo die ac nocteinterfectos filiae populi mei?
JER|9|1|Quis dabit mihi in solitudine deversorium viatorum,et de relinquam populum meum et recedam ab eis?Quia omnes adulteri sunt,coetus praevaricatorum.
JER|9|2|" Et tenderunt linguam suam quasi arcum;mendacium, et non veritas, invaluit in terra,quia de malo ad malum egressi suntet me non cognoverunt,dicit Dominus.
JER|9|3|Unusquisque se a proximo suo custodiatet in omni fratre suo non habeat fiduciam,quia omnis frater supplantat,et omnis amicus fraudulenter incedit,
JER|9|4|et vir fratrem suum decipit,et veritatem non loquuntur;docuerunt enim linguam suam loqui mendacium,inique egerunt, noluerunt converti.
JER|9|5|Iniuria super iniuriam,dolus super dolum.Renuerunt scire me ",dicit Dominus.
JER|9|6|Propterea haec dicit Dominus exercituum: Ecce ego conflabo et probabo eos;quid enim aliud faciam filiae populi mei?
JER|9|7|Sagitta vulnerans lingua eorum;dolum locuta est in ore suo:pacem cum amico suo loquituret occulte ponit ei insidias.
JER|9|8|Numquid super his non visitabo eos,dicit Dominus,aut in gente huiusmodinon ulciscetur anima mea? ".
JER|9|9|Super montes assumam fletum ac lamentumet super pascua deserti planctum,quoniam incensa sunt,eo quod non sit vir pertransiens,et non audiunt vocem gregis;a volucre caeli usque ad pecoratransmigraverunt, recesserunt.
JER|9|10|" Et dabo Ierusalem in acervos arenaeet cubilia thoum,et civitates Iudae dabo in desolationem,eo quod non sit habitator ".
JER|9|11|Quis est vir sapiens, qui intellegat hoc,et ad quem verbum oris Domini fiat,ut annuntiet istud:Quare perierit terra,exusta sit quasi desertum,eo quod non sit qui pertranseat?
JER|9|12|Et dixit Dominus: " Quia dereliquerunt legem meam, quam dedi eis, et non audierunt vocem meam et non ambulaverunt in ea;
JER|9|13|et abierunt post pravitatem cordis sui et post Baalim, quos didicerunt a patribus suis ".
JER|9|14|Idcirco haec dicit Dominus exercituum, Deus Israel: " Ecce ego cibabo populum istum absinthio et potum dabo eis aquam fellis;
JER|9|15|et dispergam eos in gentibus, quas non noverunt ipsi et patres eorum, et mittam post eos gladium, donec consumantur.
JER|9|16|Haec dicit Dominus exercituum:Attendite et vocate lamentatrices, et veniant;et ad eas, quae sapientes sunt, mittite, et properent! ".
JER|9|17|Festinentet assumant super nos lamentum:deducant oculi nostri lacrimas,et palpebrae nostrae defluant aquis.
JER|9|18|Quia vox lamentationis audita est de Sion: Quomodo vastati sumus et confusi vehementer,quia dereliquimus terram,quoniam deiecta sunt tabernacula nostra ".
JER|9|19|Audite ergo, mulieres, verbum Domini;et assumant aures vestrae sermonem oris eius,et docete filias vestras lamentum,et unaquaeque proximam suam planctum.
JER|9|20|Quia ascendit mors per fenestras nostras,ingressa est domos nostras,disperdere parvulos deforis,iuvenes de plateis.
JER|9|21|Loquere. Haec dicit Dominus: Et cadet morticinum hominisquasi stercus super faciem regioniset quasi manipulus post tergum metentis,et non est qui colligat ".
JER|9|22|Haec dicit Dominus: Non glorietur sapiens in sapientia sua,et non glorietur fortis in fortitudine sua,et non glorietur dives in divitiis suis;
JER|9|23|sed in hoc glorietur, qui gloriatur:scire et nosse me,quia ego sum Dominus, qui facio misericordiamet iudicium et iustitiam in terra;haec enim placent mihi,ait Dominus.
JER|9|24|Ecce dies veniunt, dicit Dominus, et visitabo super omnem, qui circumcisum habet praeputium,
JER|9|25|super Aegyptum et super Iudam et super Edom et super filios Ammon et super Moab et super omnes, qui attonsi sunt in comam, habitantes in deserto, quia omnes gentes habent praeputium, omnis autem domus Israel incircumcisi sunt corde ".
JER|10|1|Audite verbum, quod locutus est Dominus super vos, domus Israel.
JER|10|2|Haec dicit Dominus: Iuxta vias gentium nolite discereet a signis caeli nolite metuere,quae timent gentes,
JER|10|3|quia leges populorum vanae sunt.Quia lignum de saltu praeciditopus manuum artificis in ascia,
JER|10|4|argento et auro decoravit illud,clavis et malleis firmavit,ut non moveatur;
JER|10|5|sicut formido in cucumerario suntet non loquentur,portantur, quia incedere non valent:nolite ergo timere ea,quia nec male possunt facere nec bene ".
JER|10|6|Non est similis tui, Domine;magnus es tu,et magnum nomen tuum in fortitudine.
JER|10|7|Quis non timebit te, o rex gentium?Te enim decet,quoniam inter cunctos sapientes gentiumet in universis regnis earum nullus est similis tui.
JER|10|8|Pariter insipientes et fatui sunt;doctrina vanitatis eorum lignum est.
JER|10|9|Argentum involutum, quod de Tharsis affertur,et aurum de Ophaz,opus artificis et manuum aurificis,hyacinthus et purpura indumentum eorum;opus artificum universa haec.
JER|10|10|Dominus autem Deus verus est,ipse Deus vivens et rex sempiternus;ab indignatione eius commovebitur terra,et non sustinebunt gentes comminationem eius.
JER|10|11|Sic ergo dicetis eis: " Dii, qui caelos et terram non fecerunt, pereant de terra et de his, quae sub caelis sunt ".
JER|10|12|Qui fecit terram in fortitudine sua,firmavit orbem in sapientia suaet prudentia sua extendit caelos.
JER|10|13|Ad vocem suam dat multitudinem aquarum in caeloet elevat nebulas ab extremitatibus terrae;fulgura in pluviam facitet educit ventum de thesauris suis.
JER|10|14|Stultus factus est omnis homo absque scientia;confusus est omnis artifex in sculptili,quoniam falsum est, quod conflavit,et non est spiritus in eis.
JER|10|15|Vana sunt et opus risu dignum;in tempore visitationis suae peribunt.
JER|10|16|Non est his similis pars Iacob:qui enim formavit omnia, ipse est,et Israel tribus hereditatis eius,Dominus exercituum nomen illi.
JER|10|17|Congrega de terra sarcinam tuam,quae habitas in obsidione,
JER|10|18|quia haec dicit Dominus: Ecce ego longe proiciam habitatores terrae in hac viceet tribulabo eos, ita ut inveniant me ".
JER|10|19|Vae mihi super contritione mea,pessima plaga mea!Ego autem dixi: Plane haec infirmitas mea est,et portabo illam ".
JER|10|20|Tabernaculum meum vastatum est, omnes funiculi mei dirupti sunt;filii mei exierunt a me et non subsistunt,non est qui extendat ultra tentorium meumet erigat pelles meas.
JER|10|21|Quia stulte egerunt pastoreset Dominum non quaesierunt;propterea non prosperati sunt,et omnis grex eorum dispersus est.
JER|10|22|Vox auditionis ecce venitet commotio magna de terra aquilonis,ut ponat civitates Iudae solitudinemet habitaculum thoum.
JER|10|23|" Scio, Domine, quia non est hominis via eius,nec viri est, ut ambulet et dirigat gressus suos.
JER|10|24|Corripe me, Domine,verumtamen in iudicio et non in furore tuo,ne forte ad nihilum redigas me ".
JER|10|25|Effunde indignationem tuam super gentes,quae non cognoverunt te,et super cognationes,quae nomen tuum non invocaverunt;quia comederunt Iacobet devoraverunt eumet consumpserunt illumet pascua eius dissipaverunt.
JER|11|1|Verbum, quod factum est ad Ieremiam a Domino dicens:
JER|11|2|" Audite verba pacti huius et loquimini ad viros Iudae et habitatores Ierusalem.
JER|11|3|Et dices ad eos: Haec dicit Dominus, Deus Israel: Maledictus vir, qui non audierit verba pacti huius,
JER|11|4|quod praecepi patribus vestris in die, qua eduxi eos de terra Aegypti, de fornace ferrea, dicens: Audite vocem meam et facite omnia, quae praecipio vobis, et eritis mihi in populum, et ego ero vobis in Deum;
JER|11|5|ut suscitem iuramentum, quod iuravi patribus vestris, daturum me eis terram fluentem lacte et melle, sicut est dies haec ". Et respondi et dixi: " Amen, Domine ".
JER|11|6|Et dixit Dominus ad me: " Vociferare omnia verba haec in civitatibus Iudae et in foris Ierusalem dicens: Audite verba pacti huius et facite illa.
JER|11|7|Quia contestans contestatus sum patres vestros in die, qua eduxi eos de terra Aegypti, usque ad diem hanc; mane consurgens contestatus sum et dixi: Audite vocem meam.
JER|11|8|Et non audierunt nec inclinaverunt aurem suam, sed abierunt unusquisque in pravitate cordis sui mali; et induxi super eos omnia verba pacti huius, quod praecepi, ut facerent, et non fecerunt ".
JER|11|9|Et dixit Dominus ad me: " Inventa est coniuratio in viris Iudae et in habitatoribus Ierusalem.
JER|11|10|Reversi sunt ad iniquitates patrum suorum priorum, qui noluerunt audire verba mea; et hi ergo abierunt post deos alienos, ut servirent eis: irritum fecerunt domus Israel et domus Iudae pactum meum, quod pepigi cum patribus eorum.
JER|11|11|Quam ob rem haec dicit Dominus: Ecce ego inducam super eos mala, de quibus exire non poterunt; et clamabunt ad me, et non exaudiam eos.
JER|11|12|Et ibunt civitates Iudae et habitatores Ierusalem et clamabunt ad deos, quibus sacrificant, et non salvabunt eos in tempore afflictionis eorum.
JER|11|13|Secundum numerum enim civitatum tuarum erant dii tui, Iuda, et secundum numerum viarum Ierusalem posuistis aras confusioni, aras ad sacrificandum Baal.
JER|11|14|Tu ergo noli orare pro populo hoc et ne assumas pro eis deprecationem et orationem, quia non exaudiam in tempore clamoris eorum ad me, in tempore afflictionis eorum.
JER|11|15|Quid est dilectae meae,ut in domo mea perficiat consilia mala?Numquid vota et carnes sanctaeauferent a te malitias tuas,in quibus glorieris? ".
JER|11|16|Olivam uberem, pulchram, fructibus speciosam,vocabit Dominus nomen tuum;ad vocem strepitus grandissuccendit ignem in ea,et combusti sunt rami eius.
JER|11|17|Et Dominus exercituum, qui plantavit te, locutus est super te malum, pro malis domus Israel et domus Iudae, quae fecerunt sibi ad irritandum me, sacrificantes Baal.
JER|11|18|Tu autem, Domine, demonstrasti mihi, et cognovi;tunc ostendisti mihi opera eorum.
JER|11|19|Et ego quasi agnus mansuetus, qui portatur ad victimam; et non cognovi quia super me cogitaverunt consilia: " Caedamus lignum in vigore eius et eradamus eum de terra viventium, et nomen eius non memoretur amplius ".
JER|11|20|Tu autem, Domine exercituum,qui iudicas iuste et probas renes et corda:videam ultionem tuam ex eis;tibi enim revelavi causam meam.
JER|11|21|Propterea haec dicit Dominus super viros Anathoth, qui quaerunt animam tuam et dicunt: " Non prophetabis in nomine Domini et non morieris in manibus nostris ".
JER|11|22|Propterea haec dicit Dominus exercituum: " Ecce ego visitabo super eos: iuvenes morientur in gladio, filii eorum et filiae eorum morientur in fame,
JER|11|23|et reliquiae non erunt eis; inducam enim malum super viros Anathoth, annum visitationis eorum ".
JER|12|1|Iustus quidem tu es, Domine, si disputem tecum;verumtamen de iudiciis loquar ad te.Quare via impiorum prosperatur?Bene est omnibus, qui praevaricantur et inique agunt.
JER|12|2|Plantasti eos, et radicem miserunt,proficiunt et faciunt fructum;prope es tu ori eorumet longe a renibus eorum.
JER|12|3|Et tu, Domine, nosti me, vidisti meet probasti cor meum tecum;segrega eos quasi gregem ad victimamet sanctifica eos in diem occisionis.
JER|12|4|Usquequo lugebit terra,et herba omnis regionis siccabiturpropter malitiam habitantium in ea?Consumptum est animal et volucre,quoniam dixerunt: "Non videbit novissima nostra".
JER|12|5|" Si cum peditibus currens laborasti,quomodo contendere poteris cum equis?Cum autem in terra pacis securus fueris,quid facies in silva condensa Iordanis?
JER|12|6|Nam et fratres tui et domus patris tui,etiam ipsi fraudulenter egerunt adversum teet clamaverunt post te plena voce;ne credas eis, cum locuti fuerint tibi bona ".
JER|12|7|" Reliqui domum meam,dimisi hereditatem meam;dedi dilectam animae meaein manu inimicorum eius.
JER|12|8|Facta est mihi hereditas meaquasi leo in silva;dedit contra me vocem, ideo odivi eam.
JER|12|9|Numquid avis discolor hereditas mea mihi?Numquid aves in circuitu contra eam?Venite, congregamini, omnes bestiae campi,properate ad devorandum.
JER|12|10|Pastores multi demoliti sunt vineam meam,conculcaverunt partem meam;dederunt portionem meam desiderabilemin desertum solitudinis.
JER|12|11|Posuerunt eam in dissipationem;lugetque coram me desolata,vastata est omnis terra,quia nullus est qui recogitet corde ".
JER|12|12|Super omnes colles in deserto venerunt vastatores,quia gladius Domini devoratab extremo terrae usque ad extremum eius;non est pax universae carni.
JER|12|13|Seminaverunt triticum et spinas messuerunt,laboraverunt, et non eis proderit;confundemini a fructibus vestrispropter iram furoris Domini.
JER|12|14|Haec dicit Dominus adversum omnes vicinos meos pessimos, qui tangunt hereditatem, quam distribui populo meo Israel: "Ecce ego evellam eos de terra sua et domum Iudae evellam de medio eorum.
JER|12|15|Et erit: cum evulsero eos, convertar et miserebor eorum et reducam eos, virum ad hereditatem suam et virum in terram suam.
JER|12|16|Et erit: si eruditi didicerint vias populi mei, ut iurent in nomine meo: "Vivit Dominus!", sicut docuerunt populum meum iurare in Baal, aedificabuntur in medio populi mei.
JER|12|17|Quod si non audierint, evellam gentem illam evulsione et perditione ", ait Dominus.
JER|13|1|Haec dixit Dominus ad me: " Vade et posside tibi lumba re lineum et pones illud super lumbos tuos et in aquam non inferes illud ".
JER|13|2|Et possedi lumbare iuxta verbum Domini et posui circa lumbos meos.
JER|13|3|Et factus est sermo Domini ad me secundo dicens:
JER|13|4|" Tolle lumbare, quod possedisti, quod est circa lumbos tuos, et surgens vade ad Euphraten et absconde ibi illud in foramine petrae ".
JER|13|5|Et abii et abscondi illud ad Euphraten, sicut praeceperat mihi Dominus.
JER|13|6|Et factum est, post dies plurimos dixit Dominus ad me: " Surge, vade ad Euphraten et tolle inde lumbare, quod praecepi tibi, ut absconderes ibi ".
JER|13|7|Et abii ad Euphraten et fodi et tuli lumbare de loco, ubi absconderam illud; et ecce, computruerat lumbare, ita ut nulli usui aptum esset.
JER|13|8|Et factum est verbum Domini ad me dicens:
JER|13|9|" Haec dicit Dominus: Sic putrescere faciam superbiam Iudae et superbiam Ierusalem multam;
JER|13|10|populus iste pessimus - qui nolunt audire verba mea et ambulant in pravitate cordis sui abieruntque post deos alienos, ut servirent eis et adorarent eos - erit sicut lumbare istud, quod nulli usui aptum est.
JER|13|11|Sicut enim adhaeret lumbare ad lumbos viri, sic agglutinavi mihi omnem domum Israel et omnem domum Iudae, dicit Dominus, ut esset mihi in populum et in nomen et in laudem et in gloriam, et non audierunt.
JER|13|12|Dices ergo ad eos sermonem istum: Haec dicit Dominus, Deus Israel: Omnis laguncula implebitur vino. Et dicent ad te: "Numquid ignoramus quia omnis laguncula implebitur vino?".
JER|13|13|Et dices ad eos: Haec dicit Dominus: Ecce ego implebo omnes habitatores terrae huius et reges, qui sedent de stirpe David super thronum eius, et sacerdotes et prophetas et omnes habitatores Ierusalem ebrietate;
JER|13|14|et collidam eos, virum in fratrem suum et patres et filios pariter, ait Dominus; non parcam et non concedam neque miserebor, ut non disperdam eos.
JER|13|15|Audite et auribus percipite; nolite elevari,quia Dominus locutus est.
JER|13|16|Date Domino Deo vestro gloriam,antequam contenebrescat,et antequam offendant pedes vestriad montes caliginosos;exspectabitis lucem,et ponet eam in umbram mortiset in caliginem.
JER|13|17|Quod si hoc non audieritis,in abscondito plorabit anima meaa facie superbiae;plorans plorabitet deducet oculus meus lacrimam,quia captus est grex Domini.
JER|13|18|" Dic regi et dominatrici:In humo sedete,quoniam descendit de capite vestrocorona gloriae vestrae.
JER|13|19|Civitates austri clausae sunt,et non est qui aperiat;translata est omnis Iudatransmigratione perfecta.
JER|13|20|Leva oculos tuos et videvenientes ab aquilone:Ubi est grex, qui datus est tibi,pecus inclitum tuum?
JER|13|21|Quid dices, cum visitaverit te?Tu enim ipsa docuisti eos adversum te,amicos in caput tuum;numquid non dolores apprehendent tequasi mulierem parturientem?
JER|13|22|Quod si dixeris in corde tuo:Quare venerunt mihi haec?".Propter multitudinem iniquitatis tuaerevelatae sunt laciniae tuae,pollutae sunt plantae tuae.
JER|13|23|Numquid mutare potest Aethiops pellem suamaut pardus varietates suas?Tunc et vos poteritis benefacere,cum didiceritis malum.
JER|13|24|Et disseminabo eos quasi stipulam,quae raptatur in vento deserti.
JER|13|25|Haec sors tua parsque mensurae tuae a me,dicit Dominus,quia oblita es meiet confisa es in mendacio.
JER|13|26|Unde et ego sublevabo lacinias tuas super faciem tuam,et apparebit ignominia tua,
JER|13|27|adulteria tua et hinnitus tuus,scelus fornicationis tuae.Super colles in agro vidi abominationes tuas.Vae tibi, Ierusalem! Non mundaberis;usquequo adhuc? ".
JER|14|1|Quod factum est verbum Domini ad Ieremiam de sic citate.
JER|14|2|Luget Iuda,et portae eius languescuntet contristatae iacent in terra,et clamor Ierusalem ascendit.
JER|14|3|Maiores eorum miserunt minores suos ad aquam:venerunt ad cisternas,non invenerunt aquam;reportaverunt vasa sua vacua,confusi sunt et afflictiet operuerunt capita sua.
JER|14|4|Propter terrae vastitatem,quia non venit pluvia in terram,confusi sunt agricolae,operuerunt capita sua.
JER|14|5|Nam et cerva in agro peperit et reliquit,quia non erat herba.
JER|14|6|Et onagri steterunt in collibus,traxerunt aerem quasi thoes;defecerunt oculi eorum,quia non erat herba.
JER|14|7|" Si iniquitates nostrae testificantur adversus nos,Domine, fac propter nomen tuum,quoniam multae sunt aversiones nostrae,tibi peccavimus.
JER|14|8|Exspectatio Israel,salvator eius in tempore tribulationis,quare quasi peregrinus es in terraet quasi viator declinans ad pernoctandum?
JER|14|9|Quare es velut vir attonitus,ut fortis, qui non potest salvare?Tu autem in medio nostri es, Domine,et nomen tuum invocatum est super nos;ne derelinquas nos ".
JER|14|10|Haec dicit Dominus populo huic: " Ita diligunt vagari, pedes suos non prohibent et Domino non placent ". Nunc recordatus est iniquitatum eorum et visitat peccata eorum.
JER|14|11|Et dixit Dominus ad me: " Noli orare pro populo isto in bonum.
JER|14|12|Cum ieiunaverint, non exaudiam preces eorum; et, si obtulerint holocautomata et oblationes, non suscipiam ea; quoniam gladio et fame et peste consumam eos ".
JER|14|13|Et dixi: " Heu, Domine Deus! Ecce prophetae dicunt eis: "Non videbitis gladium, et fames non erit in vobis, sed pacem veram dabit vobis in loco isto" ".
JER|14|14|Et dixit Dominus ad me: " Falso prophetae vaticinantur in nomine meo: non misi eos et non praecepi eis neque locutus sum ad eos; visionem mendacem et divinationem et fraudulentiam et seductionem cordis sui prophetant vobis.
JER|14|15|Idcirco haec dicit Dominus contra prophetas, qui prophetant in nomine meo, quos ego non misi, dicentes: "Gladius et fames non erit in terra hac": In gladio et fame consumentur prophetae illi;
JER|14|16|et homines, quibus prophetant, erunt proiecti in viis Ierusalem prae fame et gladio, et non erit qui sepeliat eos: ipsi et uxores eorum, filii et filiae eorum, et effundam super eos malum suum.
JER|14|17|Et dices ad eos verbum istud:Deducant oculi mei lacrimamper noctem et diem, et non taceant,quoniam contritione magna contrita estvirgo filia populi mei,plaga pessima vehementer.
JER|14|18|Si egressus fuero ad agros,ecce occisi gladio;et, si introiero in civitatem,ecce attenuati fame;propheta quoque et sacerdosabierunt per terram nescientes ".
JER|14|19|Numquid proiciens abiecisti Iudam,aut Sion abominata est anima tua?Quare ergo percussisti nos,ita ut nulla sit sanitas?Exspectavimus pacem, et non est bonum,et tempus curationis, et ecce turbatio.
JER|14|20|Cognovimus, Domine, impietates nostras,iniquitates patrum nostrorum, quia peccavimus tibi.
JER|14|21|Ne des nos in opprobrium propter nomen tuum,ne facias contumeliam solio gloriae tuae;recordare, ne irritum facias foedus tuum nobiscum.
JER|14|22|Numquid sunt in sculptilibus gentium, qui pluant,aut caeli possunt dare imbres?Nonne tu es Dominus Deus noster,quem exspectamus?Tu enim fecisti omnia haec.
JER|15|1|Et dixit Dominus ad me: " Si steterit Moyses et Samuel co ram me, non est anima mea ad populum istum; eice illos a facie mea, et egrediantur.
JER|15|2|Quod si dixerint ad te: "Quo egrediemur?", dices ad eos: Haec dicit Dominus:Qui ad mortem, ad mortem;et qui ad gladium, ad gladium;et qui ad famem, ad famem;et qui ad captivitatem, ad captivitatem.
JER|15|3|Et mandabo super eos quattuor species, dicit Dominus: gladium ad occisionem et canes ad lacerandum et volatilia caeli et bestias terrae ad devorandum et dissipandum.
JER|15|4|Et dabo eos in commotionem universis regnis terrae, propter Manassem filium Ezechiae regem Iudae, super omnibus, quae fecit in Ierusalem.
JER|15|5|Quis enim miserebitur tui, Ierusalem,aut quis contristabitur pro te,aut quis ibit ad rogandum de pace tua?
JER|15|6|Tu reppulisti me,dicit Dominus,retrorsum abiisti;et extendi manum meam super te et interfeci te:laboravi miserans.
JER|15|7|Et ventilavi eos ventilabroin portis terrae;orbavi et disperdidi populum meum:a viis suis non sunt reversi.
JER|15|8|Multiplicatae sunt mihi viduae eiussuper arenam maris,induxi eis super matremmilitem vastatorem meridie,misi super eam repenteperturbationem et terrorem.
JER|15|9|Infirmata est, quae peperit septem,exhalavit animam suam;occidit ei sol, cum adhuc esset dies,confusa est et erubuit,et residuos eorum in gladium daboin conspectu inimicorum eorum ",ait Dominus.
JER|15|10|Vae mihi, mater mea,quoniam genuisti me virum rixaeet virum discordiae in universa terra!Non feneravi, nec feneravit mihi quisquam;omnes maledicunt mihi.
JER|15|11|Amen, Domine, ministravi tibi in bonum,intercessi apud te in tempore afflictioniset in tempore tribulationis pro inimico.
JER|15|12|Numquid frangitur ferroferrum aquilonis et aes?
JER|15|13|" Divitias tuas et thesauros tuosin direptionem dabo gratis,propter omnia peccata tua,in omnibus terminis tuis.
JER|15|14|Et servire te faciam inimicis tuisin terra, quam nescis,quia ignis succensus est in furore meo:super vos ardebit ".
JER|15|15|Tu scis, Domine;recordare mei et visita meet vindica me de his, qui persequuntur me;noli in patientia tua abripere me,scito quoniam sustinui pro te opprobrium.
JER|15|16|Inventi sunt sermones tui, et comedi eos,et factum est mihi verbum tuumin gaudium et in laetitiam cordis mei,quoniam invocatum est nomen tuum super me,Domine, Deus exercituum.
JER|15|17|Non sedi in concilio ludentiumet gloriatus sum;a facie manus tuae solus sedebam,quoniam indignatione replesti me.
JER|15|18|Quare factus est dolor meus perpetuus,et plaga mea desperabilis renuit curari?Factus es mihi quasi rivus mendax,aquae infideles.
JER|15|19|Propter hoc haec dixit Dominus: Si converteris, convertam te,et ante faciem meam stabis;et si separaveris pretiosum a vili,quasi os meum eris;convertentur ipsi ad te,et tu non converteris ad eos.
JER|15|20|Et dabo te populo huicin murum aereum fortem;et bellabunt adversum teet non praevalebunt,quia ego tecum sum,ut salvem te et eruam te,dicit Dominus.
JER|15|21|Et liberabo te de manu pessimorumet redimam te de manu fortium ".
JER|16|1|Et factum est verbum Domi ni ad me dicens:
JER|16|2|" Non acci pies uxorem, et non erunt tibi filii et filiae in loco isto.
JER|16|3|Quia haec dicit Dominus super filios et filias, qui generantur in loco isto, et super matres eorum, quae genuerunt eos, et super patres eorum, de quorum stirpe sunt nati in terra hac:
JER|16|4|Mortibus aegrotationum morientur, non plangentur et non sepelientur; in sterquilinium super faciem terrae erunt et gladio et fame consumentur, et erit cadaver eorum in escam volatilibus caeli et bestiis terrae ".
JER|16|5|Haec enim dixit Dominus: "Ne ingrediaris domum convivii neque vadas ad plangendum neque lugebis eos, quia abstuli pacem meam a populo isto, dicit Dominus, misericordiam et miserationes.
JER|16|6|Et morientur grandes et parvi in terra ista, non sepelientur neque plangentur, et non se incident, neque calvitium fiet pro eis.
JER|16|7|Et non frangent lugenti panem ad consolandum super mortuo et non dabunt ei calicem ad consolandum super patre suo et matre.
JER|16|8|Et domum convivii non ingredieris, ut sedeas cum eis et comedas et bibas.
JER|16|9|Quia haec dicit Dominus exercituum, Deus Israel: Ecce ego auferam de loco isto in oculis vestris et in diebus vestris vocem gaudii et vocem laetitiae, vocem sponsi et vocem sponsae.
JER|16|10|Et cum annuntiaveris populo huic omnia verba haec, et dixerint tibi: Quare locutus est Dominus super nos omne malum grande istud? Quae iniquitas nostra et quod peccatum nostrum, quod peccavimus Domino Deo nostro?",
JER|16|11|dices ad eos: Quia dereliquerunt me patres vestri, ait Dominus, et abierunt post deos alienos et servierunt eis et adoraverunt eos et me dereliquerunt et legem meam non custodierunt.
JER|16|12|Sed et vos peius operati estis quam patres vestri: ecce enim ambulat unusquisque post pravitatem cordis sui mali, ut me non audiat.
JER|16|13|Et eiciam vos de terra hac in terram, quam ignoratis, vos et patres vestri; et servietis ibi diis alienis, die ac nocte, quia non dabo vobis gratiam.
JER|16|14|Propterea ecce dies veniunt, dicit Dominus, et non dicetur ultra: Vivit Dominus, qui eduxit filios Israel de terra Aegypti!",
JER|16|15|sed: "Vivit Dominus, qui eduxit filios Israel de terra aquilonis et de universis terris, ad quas eieci eos!". Et reducam eos in terram suam, quam dedi patribus eorum.
JER|16|16|Ecce ego mittam piscatores multos, dicit Dominus, et piscabuntur eos; et post haec mittam eis multos venatores, et venabuntur eos de omni monte et de omni colle et de cavernis petrarum.
JER|16|17|Quia oculi mei super omnes vias eorum: non sunt absconditae a facie mea, et non est occulta iniquitas eorum ab oculis meis.
JER|16|18|Et reddam primum dupliciter iniquitates et peccata eorum, quia contaminaverunt terram meam in morticinis idolorum suorum et abominationibus suis impleverunt hereditatem meam ".
JER|16|19|Domine, fortitudo mea et praesidium meumet refugium meum in die tribulationis;ad te gentes venient ab extremis terrae et dicent: Vere mendacium possederunt patres nostri,vanitatem, quae nihil prodest ".
JER|16|20|Numquid faciet sibi homo deos,et ipsi non sunt dii?
JER|16|21|" Idcirco ecce ego ostendam eis per vicem hanc,ostendam eis manum meam et virtutem meam,et scient quia nomen mihi Dominus ".
JER|17|1|Peccatum Iudae scriptum est stilo ferreo,in ungue adamantino exaratumsuper tabulam cordis eorumet in cornibus ararum eorum,
JER|17|2|ut recordarentur filii eorum ararum suarumet palorum suorum iuxta ligna frondentiain collibus excelsis,
JER|17|3|montibus in campo. Divitias tuas, omnes thesauros tuosin direptionem dabo,excelsa tua propter peccatain universis finibus tuis.
JER|17|4|Et relinques hereditatem tuam,quam dedi tibi;et servire te faciam inimicis tuisin terra, quam ignoras,quoniam ignem succendistis in naribus meis;usque in aeternum ardebit ".
JER|17|5|Haec dicit Dominus: Maledictus homo, qui confidit in homineet ponit carnem brachium suum,et a Domino recedit cor eius;
JER|17|6|erit enim quasi myricae in desertoet non videbit, cum venerit bonum,sed habitabit in siccitate in deserto,in terra salsuginis et inhabitabili.
JER|17|7|Benedictus vir, qui confidit in Domino,et erit Dominus fiducia eius;
JER|17|8|et erit quasi lignum,quod transplantatur super aquas,quod ad humorem mittit radices suaset non timebit, cum venerit aestus;et erit folium eius viride,et in anno siccitatis non erit sollicitumnec aliquando desinet facere fructum
JER|17|9|Dolosum est cor super omnia et insanabile;quis cognoscet illud?
JER|17|10|Ego Dominus scrutans cor et probans renes,qui do unicuique iuxta viam suamet iuxta fructum operum suorum.
JER|17|11|Perdix fovit, quae non peperit,ita faciens divitias sed non in iudicio.In dimidio dierum suorum derelinquet easet in novissimo suo erit insipiens ".
JER|17|12|Solium gloriae, altitudo a principio,locus sanctificationis nostrae!
JER|17|13|Exspectatio Israel, Domine,omnes, qui te derelinquunt, confundentur;recedentes a te in terra scribentur,quoniam dereliquerunt venamaquarum viventium, Dominum.
JER|17|14|Sana me, Domine, et sanabor;salvum me fac, et salvus ero,quoniam laus mea tu es.
JER|17|15|Ecce ipsi dicunt ad me: Ubi est verbum Domini? Veniat ".
JER|17|16|Et ego non institi pro malo apud teet diem calamitatis non desideravi,tu scis: quod egressum est de labiis meis,rectum in conspectu tuo fuit.
JER|17|17|Non sis mihi tu formidini;refugium meum tu in die afflictionis.
JER|17|18|Confundantur, qui me persequuntur,et non confundar ego;paveant illi, et non paveam ego;induc super eos diem afflictioniset duplici contritione contere eos.
JER|17|19|Haec dixit Dominus ad me: " Vade et sta in porta Filiorum populi, per quam ingrediuntur reges Iudae et egrediuntur, et in cunctis portis Ierusalem;
JER|17|20|et dices ad eos: Audite verbum Domini, reges Iudae et omnis Iuda cunctique habitatores Ierusalem, qui ingredimini per portas istas.
JER|17|21|Haec dicit Dominus: Custodite animas vestras et nolite portare pondera in die sabbati nec inferatis per portas Ierusalem;
JER|17|22|et nolite efferre onera de domibus vestris in die sabbati et omne opus non facietis: sanctificate diem sabbati, sicut praecepi patribus vestris.
JER|17|23|Et non audierunt nec inclinaverunt aurem suam; sed induraverunt cervicem suam, ne audirent me et ne acciperent disciplinam.
JER|17|24|Et erit: si audieritis me, dicit Dominus, ut non inferatis onera per portas civitatis huius in die sabbati, et si sanctificaveritis diem sabbati, ne faciatis in eo omne opus,
JER|17|25|ingredientur per portas civitatis huius reges et principes sedentes super solium David et ascendentes in curribus et equis, ipsi et principes eorum, viri Iudae et habitatores Ierusalem; et habitabitur civitas haec in sempiternum.
JER|17|26|Et venient de civitatibus Iudae et de circuitu Ierusalem et de terra Beniamin et de Sephela et de montuosis et a Nageb, portantes holocaustum et victimam et sacrificium et tus, et inferent oblationem laudis in domum Domini.
JER|17|27|Si autem non audieritis me, ut sanctificetis diem sabbati et ne portetis onus intrantes per portas Ierusalem in die sabbati, succendam ignem in portis eius, et devorabit domos Ierusalem et non exstinguetur ".
JER|18|1|Verbum, quod factum est ad Ieremiam a Domino dicens:
JER|18|2|" Surge et descende in domum figuli et ibi audies verba mea ".
JER|18|3|Et descendi in domum figuli, et ecce ipse faciebat opus super rotam;
JER|18|4|et dissipatum est vas, quod ipse faciebat e luto manibus suis, et rursus fecit illud vas alterum, sicut placuerat in oculis eius, ut faceret.
JER|18|5|Et factum est verbum Domini ad me dicens:
JER|18|6|" Numquid sicut figulus iste non potero vobis facere, domus Israel?, ait Dominus. Ecce, sicut lutum in manu figuli, sic vos in manu mea, domus Israel.
JER|18|7|Repente loquar adversum gentem et adversum regnum, ut eradicem et destruam et disperdam illud;
JER|18|8|si paenitentiam egerit gens illa a malo suo, propter quod locutus sum adversus eam, agam et ego paenitentiam super malo, quod cogitavi ut facerem ei.
JER|18|9|Et subito loquar de gente et de regno, ut aedificem et plantem illud;
JER|18|10|si fecerit malum in oculis meis, ut non audiat vocem meam, paenitentiam agam super bono, quod locutus sum ut facerem ei.
JER|18|11|Nunc ergo, dic viro Iudae et habitatoribus Ierusalem dicens: Haec dicit Dominus: Ecce ego fingo contra vos malum et cogito contra vos cogitationem; revertatur unusquisque a via sua mala, et dirigite vias vestras et opera vestra ".
JER|18|12|Qui dixerunt: " Vanum est; post cogitationes enim nostras ibimus et unusquisque pravitatem cordis sui mali faciemus ".
JER|18|13|Ideo haec dicit Dominus: Interrogate gentes:quis audivit talia horribilia,quae fecit nimis virgo Israel?
JER|18|14|Numquid deficiet de petra agrinix Libani,aut arescent aquae erumpentesfrigidae et defluentes?
JER|18|15|Quia oblitus est mei populus meus,vanitati sacrificanteset impingentes in viis suis,in semitis antiquis,ut ambularent per callesin itinere non trito,
JER|18|16|ut poneret terram eorum in desolationemet in sibilum sempiternum:omnis, qui praeterierit per eam, obstupescetet movebit caput suum.
JER|18|17|Sicut ventus urens dispergam eoscoram inimico;dorsum et non faciem ostendam eis in die perditionis eorum ".
JER|18|18|Et dixerunt: " Venite, et cogitemus contra Ieremiam cogitationes; non enim peribit lex a sacerdote, neque consilium a sapiente, nec sermo a propheta. Venite, et percutiamus eum lingua et non attendamus ad universos sermones eius ".
JER|18|19|Attende, Domine, ad meet audi vocem adversariorum meorum.
JER|18|20|Numquid redditur pro bono malum,quia foderunt foveam animae meae?Recordare quod steterim in conspectu tuo,ut loquerer pro eis bonumet averterem indignationem tuam ab eis.
JER|18|21|Propterea da filios eorum in famemet deduc eos in manus gladii;fiant uxores eorum absque liberis et viduae,et viri eorum interficiantur morte,iuvenes eorum confodiantur gladio in proelio.
JER|18|22|Audiatur clamor de domibus eorum;adduces enim super eos latronem repente,quia foderunt foveam, ut caperent me,et laqueos absconderunt pedibus meis.
JER|18|23|Tu autem, Domine, scis omne consilium eorumadversum me in mortem;ne propitieris iniquitati eorum,et peccatum eorum a facie tua non deleatur.Fiant corruentes in conspectu tuo;in tempore furoris tui abutere eis.
JER|19|1|Haec dicit Dominus: " Vade et eme lagunculam figuli testeam et accipe de senioribus populi et de senioribus sacerdotum
JER|19|2|et egredere ad vallem Benennom, quae est iuxta introitum portae Fictilium, et praedicabis ibi verba, quae ego loquar ad te,
JER|19|3|et dices: Audite verbum Domini, reges Iudae et habitatores Ierusalem: Haec dicit Dominus exercituum, Deus Israel: Ecce ego inducam afflictionem super locum istum, ita ut omnis, qui audierit illam, tinniant aures eius,
JER|19|4|eo quod dereliquerint me et alienum fecerint locum istum et sacrificaverint in eo diis alienis, quos nescierunt ipsi et patres eorum et reges Iudae; et repleverunt locum istum sanguine innocentium;
JER|19|5|et aedificaverunt excelsa Baal ad comburendos filios suos igne in holocaustum Baal: quae non praecepi nec locutus sum, nec ascenderunt in cor meum.
JER|19|6|Propterea ecce dies veniunt, dicit Dominus, et non vocabitur amplius locus iste Topheth et vallis Benennom sed vallis Occisionis.
JER|19|7|Et dissipabo consilium Iudae et Ierusalem in loco isto; et subvertam eos gladio in conspectu inimicorum suorum et in manu quaerentium animas eorum et dabo cadavera eorum escam volatilibus caeli et bestiis terrae.
JER|19|8|Et ponam civitatem hanc in stuporem et in sibilum; omnis, qui praeterierit per eam, obstupescet et sibilabit super universa plaga eius.
JER|19|9|Et cibabo eos carnibus filiorum suorum et carnibus filiarum suarum; et unusquisque carnem amici sui comedet in obsidione et in angustia, in qua concludent eos inimici eorum et qui quaerunt animas eorum.
JER|19|10|Et conteres lagunculam in oculis virorum, qui ibunt tecum,
JER|19|11|et dices ad eos: Haec dicit Dominus exercituum: Sic conteram populum istum et civitatem istam, sicut conteritur vas figuli, quod non potest ultra instaurari; et in Topheth sepelientur, eo quod non sit alius locus ad sepeliendum.
JER|19|12|Sic faciam loco huic, ait Dominus, et habitatoribus eius, ut ponam civitatem istam sicut Topheth;
JER|19|13|et erunt domus Ierusalem et domus regum Iudae sicut locus Topheth, immundae: omnes domus, in quarum domatibus sacrificaverunt omni militiae caeli et libaverunt libamina diis alienis ".
JER|19|14|Venit autem Ieremias de Topheth, quo miserat eum Dominus ad prophetandum, et stetit in atrio domus Domini et dixit ad omnem populum:
JER|19|15|" Haec dicit Dominus exercituum, Deus Israel: Ecce ego inducam super civitatem hanc et super omnes urbes eius universa mala, quae locutus sum adversum eam, quoniam induraverunt cervicem suam, ut non audirent sermones meos ".
JER|20|1|Et audivit Phassur filius Em mer sacerdos, qui constitutus erat princeps in domo Domini, Ieremiam prophetantem sermones istos;
JER|20|2|et percussit Phassur Ieremiam prophetam et misit eum in nervum, quod erat in porta Beniamin superiore in domo Domini.
JER|20|3|Cumque illuxisset in crastinum, eduxit Phassur Ieremiam de nervo; et dixit ad eum Ieremias: " Non Phassur vocavit Dominus nomen tuum sed Pavorem undique.
JER|20|4|Quia haec dicit Dominus: Ecce ego dabo te in pavorem, te et omnes amicos tuos, et corruent gladio inimicorum suorum, et oculi tui videbunt; et omnem Iudam dabo in manu regis Babylonis, et traducet eos in Babylonem et percutiet eos gladio.
JER|20|5|Et dabo universam substantiam civitatis huius et omnem laborem eius omneque pretium et cunctos thesauros regum Iudae dabo in manu inimicorum eorum; et diripient eos et tollent et ducent in Babylonem.
JER|20|6|Tu autem, Phassur et omnes habitatores domus tuae, ibitis in captivitatem; et in Babylonem venies et ibi morieris ibique sepelieris, tu et omnes amici tui, quibus prophetasti mendacium ".
JER|20|7|Seduxisti me, Domine, et seductus sum;fortior me fuisti et invaluisti.Factus sum in derisum tota die,omnes subsannant me.
JER|20|8|Quia quotiescumque loquor, vociferor,iniquitatem et vastitatem clamito;et factus est mihi sermo Dominiin opprobrium et in derisum tota die.
JER|20|9|Et dixi: " Non recordabor eiusneque loquar ultra in nomine illius ".Et factus est in corde meo quasi ignis exaestuansclaususque in ossibus meis:et defeci, ferre non sustinens.
JER|20|10|Audivi enim contumelias multorumet terrorem in circuitu: Denuntiate, et denuntiemus eum ".Omnes pacifici mei observabant lapsum meum: Forte decipietur, et praevalebimus adversus eumet consequemur ultionem ex eo ".
JER|20|11|Dominus autem mecum est quasi bellator fortis;idcirco, qui persequuntur me,cadent et infirmi erunt.Confundentur vehementer, quia non prosperati sunt;opprobrium sempiternum, quod numquam delebitur.
JER|20|12|Et tu, Domine exercituum,probator iusti, qui vides renes et cor,videam, quaeso, ultionem tuam ex eis;tibi enim revelavi causam meam.
JER|20|13|Cantate Domino, laudate Dominum,quia liberavit animam pauperisde manu malorum.
JER|20|14|Maledicta dies, in qua natus sum;dies, in qua peperit me mater mea,non sit benedicta.
JER|20|15|Maledictus vir, qui annuntiavit patri meodicens: " Natus est tibi puer masculus "et gaudio laetificavit eum;
JER|20|16|sit homo ille, ut sunt civitates,quas subvertit Dominuset non paenituit eum:audiat clamorem maneet ululatum in tempore meridiano,
JER|20|17|qui non me interfecit a vulva,ut fieret mihi mater mea sepulcrum,et vulva eius conceptus aeternus.
JER|20|18|Quare de vulva egressus sum,ut viderem laborem et dolorem,et consumerentur in confusione dies mei?
JER|21|1|Verbum, quod factum est ad Ieremiam a Domino, quando misit ad eum rex Sedecias Phassur filium Melchiae et Sophoniam filium Maasiae sacerdotem dicens:
JER|21|2|" Interroga pro nobis Dominum, quia Nabuchodonosor rex Babylonis proeliatur adversum nos; si forte faciat Dominus nobiscum secundum omnia mirabilia sua, et recedat a nobis ".
JER|21|3|Et dixit Ieremias ad eos: " Sic dicetis Sedeciae:
JER|21|4|Haec dicit Dominus, Deus Israel: Ecce ego convertam vasa belli, quae in manibus vestris sunt et quibus vos pugnatis adversum regem Babylonis et Chaldaeos, qui obsident vos in circuitu murorum; et congregabo eos in medio civitatis huius.
JER|21|5|Et debellabo ego vos in manu extenta et in brachio forti et in furore et in indignatione et in ira grandi
JER|21|6|et percutiam habitatores civitatis huius, homines et bestias: pestilentia magna morientur.
JER|21|7|Et post haec, ait Dominus, dabo Sedeciam regem Iudae et servos eius et populum eius, qui derelicti sunt in civitate hac a peste et gladio et fame, in manu Nabuchodonosor regis Babylonis et in manu inimicorum eorum et in manu quaerentium animam eorum; et percutiet eos in ore gladii et non flectetur neque parcet nec miserebitur.
JER|21|8|Et ad populum hunc dices: Haec dicit Dominus: Ecce ego do coram vobis viam vitae et viam mortis:
JER|21|9|qui habitaverit in urbe hac, morietur gladio et fame et peste; qui autem egressus fuerit et transfugerit ad Chaldaeos, qui obsident vos, vivet, et erit ei anima sua quasi spolium.
JER|21|10|Posui enim faciem meam super civitatem hanc in malum et non in bonum, ait Dominus: in manu regis Babylonis dabitur, et exuret eam igni.
JER|21|11|Et domui regis Iudae:Audite verbum Domini,
JER|21|12|domus David. Haec dicit Dominus:Iudicate mane iudiciumet eruite vi oppressum de manu expoliantis,ne forte egrediatur ut ignis indignatio meaet succendatur, et non sit qui exstinguat,propter malitiam operum vestrorum.
JER|21|13|Ecce ego ad te, habitatricem vallis,petram in planitie,ait Dominus;qui dicitis: "Quis invadet nos?Et quis ingredietur domos nostras?".
JER|21|14|Et visitabo super vos iuxta fructum operum vestrorum,dicit Dominus;et succendam ignem in saltu eius,et devorabit omnia in circuitu eius ".
JER|22|1|Haec dicit Dominus: " Descende in domum regis Iudae et loqueris ibi verbum hoc
JER|22|2|et dices: Audi verbum Domini, rex Iudae, qui sedes super solium David, tu et servi tui et populus tuus, qui ingredimini per portas istas.
JER|22|3|Haec dicit Dominus: Facite iudicium et iustitiam et liberate vi oppressum de manu expoliantis et advenam et pupillum et viduam nolite affligere neque opprimatis inique et sanguinem innocentem ne effundatis in loco isto.
JER|22|4|Si enim facientes feceritis verbum istud, ingredientur per portas domus huius reges, sedentes de genere David super thronum eius et ascendentes currus et equos, ipsi et servi et populus eorum.
JER|22|5|Quod si non audieritis verba haec, in memetipso iuravi, dicit Dominus, quia in solitudinem erit domus haec.
JER|22|6|Quia haec dicit Dominus super domum regis Iudae:Galaad tu mihi,caput Libani,verumtamen ponam te solitudinem,urbes inhabitabiles,
JER|22|7|et sanctificabo super teinterficientem virum et arma eius,et succident electas cedros tuaset praecipitabunt in ignem.
JER|22|8|Et pertransibunt gentes multae per civitatem hanc, et dicet unusquisque proximo suo: "Quare fecit Dominus sic civitati huic grandi?".
JER|22|9|Et respondebunt: "Eo quod dereliquerint pactum Domini Dei sui et adoraverint deos alienos et servierint eis" ".
JER|22|10|Nolite flere mortuumneque lugeatis super eum fletu;plangite eum, qui egreditur,quia non revertetur ultranec videbit terram nativitatis suae.
JER|22|11|Quia haec dicit Dominus ad Sellum filium Iosiae regem Iudae, qui regnavit pro Iosia patre suo: " Qui egressus est de loco isto, non revertetur huc amplius,
JER|22|12|sed in loco, ad quem transtulerunt eum, ibi morietur et terram istam non videbit amplius ".
JER|22|13|Vae, qui aedificat domum suam in iniustitiaet cenacula sua non in iudicio,proximum suum servire facit gratiset mercedem eius non reddet ei;
JER|22|14|qui dicit: " Aedificabo mihi domum latamet cenacula spatiosa ";qui aperit sibi fenestraset facit laquearia cedrinapingitque sinopide!
JER|22|15|Numquid regnabis,quoniam gloriaris in cedris?Pater tuus numquid non comedit et bibit?Sed fecit iudicium et iustitiam,tunc bene erat ei.
JER|22|16|Iudicavit causam pauperis et egeni,tunc bene. Numquid non hoc est nosse me? ",dicit Dominus.
JER|22|17|Tui vero oculi et cor tuum nonnisi ad avaritiamet ad sanguinem innocentem fundendumet ad calumniam et ad oppressionem faciendam.
JER|22|18|Propterea haec dicit Dominus ad Ioachim filium Iosiae regem Iudae: Non plangent eum:Vae, frater meus!" et "Vae, soror!".Non concrepabunt ei:Vae, domine!" et "Vae, inclite!".
JER|22|19|Sepultura asini sepelietur,tractus et proiectus longeextra portas Ierusalem ".
JER|22|20|Ascende Libanum et clamaet in Basan da vocem tuamet clama de Abarim,quia contriti sunt omnes amatores tui.
JER|22|21|Locutus sum ad te in securitate tua,et dixisti: " Non audiam! ".Haec est via tua ab adulescentia tua,quia non audisti vocem meam.
JER|22|22|Omnes pastores tuos pascet ventus,et amatores tui in captivitatem ibunt,quia tunc confunderis et erubescesab omni malitia tua.
JER|22|23|Quae sedes in Libanoet nidificas in cedris,quomodo congemisces,cum venerint tibi doloresquasi dolores parturientis!
JER|22|24|" Vivo ego, dicit Dominus, quia si fuerit Iechonias, filius Ioachim rex Iudae, anulus in manu dextera mea, inde evellam eum
JER|22|25|et dabo te in manu quaerentium animam tuam et in manu, quorum tu formidas faciem, in manu Nabuchodonosor, regis Babylonis, et in manu Chaldaeorum;
JER|22|26|et mittam te et matrem tuam, quae genuit te, in terram alienam, in qua nati non estis, ibique moriemini;
JER|22|27|et in terram, ad quam ipsi levant animam suam, ut revertantur, illuc non revertentur ".
JER|22|28|Numquid vas despectum et contritum, vir iste Iechonias? Numquid vas absque omni voluptate? Quare abiecti sunt, ipse et semen eius, et proiecti in terram, quam ignoraverunt?
JER|22|29|Terra, terra, terra, audi sermonem Domini!
JER|22|30|Haec dicit Dominus: " Scribite virum istum sterilem, virum, qui in diebus suis non prosperabitur; nec enim erit de semine eius vir, qui sedeat super solium David et potestatem habeat ultra in Iuda ".
JER|23|1|"Vae pastoribus, qui disper dunt et dissipant gregem pascuae meae!, dicit Dominus.
JER|23|2|Ideo haec dicit Dominus, Deus Israel, ad pastores, qui pascunt populum meum: Vos dissipastis gregem meum et eiecistis eos et non visitastis eos; ecce ego visitabo super vos malitiam operum vestrorum, ait Dominus.
JER|23|3|Et ego congregabo reliquias gregis mei de omnibus terris, ad quas eiecero eos, et convertam eos ad rura sua, et crescent et multiplicabuntur.
JER|23|4|Et suscitabo super eos pastores, et pascent eos; non formidabunt ultra et non pavebunt, et nullus quaeretur ex numero, dicit Dominus.
JER|23|5|Ecce dies veniunt,dicit Dominus,et suscitabo David germen iustum;et regnabit rex et sapiens eritet faciet iudicium et iustitiam in terra.
JER|23|6|In diebus illis salvabitur Iuda,et Israel habitabit confidenter;et hoc est nomen, quod vocabunt eum:Dominus iustitia nostra.
JER|23|7|Propter hoc ecce dies veniunt, dicit Dominus, et non dicent ultra: Vivit Dominus, qui eduxit filios Israel de terra Aegypti!",
JER|23|8|sed: "Vivit Dominus, qui eduxit et adduxit semen domus Israel de terra aquilonis et de cunctis terris!", ad quas eieceram eos; et habitabunt in terra sua ".
JER|23|9|Ad prophetas.Contritum est cor meum in medio mei,contremuerunt omnia ossa mea;factus sum quasi vir ebriuset quasi homo madidus a vino,a facie Dominiet a facie verborum sanctorum eius;
JER|23|10|quia adulteris repleta est terra,quia a facie maledictionis luxit terra,arefacta sunt arva deserti,factus est cursus eorum malus,et fortitudo eorum iniustitia.
JER|23|11|" Propheta namque et sacerdos polluti sunt,et in domo mea inveni malum eorum,ait Dominus.
JER|23|12|Idcirco via eorum erit quasi lubricum;in tenebras proicientur et cadent in eis;afferam enim super eos mala,annum visitationis eorum,ait Dominus.
JER|23|13|Et in prophetis Samariae vidi fatuitatem:prophetabant in Baalet decipiebant populum meum Israel.
JER|23|14|Et in prophetis Ierusalem vidi horribilia:adulterium faciunt et in mendacio ambulant;et confortaverunt manus pessimorum,ut non converteretur unusquisque a malitia sua:facti sunt mihi omnes ut Sodoma,et habitatores eius quasi Gomorra ".
JER|23|15|Propterea haec dicit Dominus exercituum ad prophetas: Ecce ego cibabo eos absinthioet potabo eos felle;a prophetis enim Ierusalemegressa est pollutio super omnem terram.
JER|23|16|Haec dicit Dominus exercituum: Nolite audire verba prophetarum, qui prophetant vobis et decipiunt vos; visionem cordis sui loquuntur, non de ore Domini.
JER|23|17|Dicunt his, qui despiciunt me:Locutus est Dominus: Pax erit vobis";et omni, qui ambulat in pravitate cordis sui,dixerunt: "Non veniet super vos malum".
JER|23|18|Quis enim affuit in consilio Domini et vidit et audivit sermonem eius? Quis consideravit verbum illius et audivit?
JER|23|19|Ecce turbo Domini, indignatio egressa est,et tempestas erumpens super caput impiorum irruet.
JER|23|20|Non cessabit furor Domini, usque dum faciatet usque dum compleat cogitationes cordis sui;in novissimis diebus intellegetis consilium eius.
JER|23|21|Non mittebam prophetas,et ipsi currebant;non loquebar ad eos,et ipsi prophetabant.
JER|23|22|Si stetissent in consilio meo,nota fecissent verba mea populo meoet avertissent utique eos a via sua malaet ab operibus suis pessimis.
JER|23|23|Putasne Deus e vicino ego sum,dicit Dominus,et non Deus de longe?
JER|23|24|Si occultabitur vir in absconditis,ego non videbo eum?,dicit Dominus.Numquid non caelum et terram ego impleo?,dicit Dominus.
JER|23|25|Audivi, quae dixerunt prophetae prophetantes in nomine meo mendacium atque dicentes: "Somniavi, somniavi".
JER|23|26|Usquequo istud est in corde prophetarum vaticinantium mendacium et prophetantium seductionem cordis sui?
JER|23|27|Qui volunt facere, ut obliviscatur populus meus nominis mei, propter somnia eorum, quae narrat unusquisque ad proximum suum, sicut obliti sunt patres eorum nominis mei propter Baal.
JER|23|28|Propheta, qui habet somnium, narret somnium et, qui habet sermonem meum, loquatur sermonem meum vere.Quid paleis ad triticum?,dicit Dominus.
JER|23|29|Numquid non verba mea sunt quasi ignis,dicit Dominus,et quasi malleus conterens petram?
JER|23|30|Propterea ecce ego ad prophetas, ait Dominus, qui furantur verba mea unusquisque a proximo suo.
JER|23|31|Ecce ego ad prophetas, ait Dominus, qui assumunt linguas suas et aiunt: Dicit Dominus".
JER|23|32|Ecce ego ad prophetantes somnia mendacii, ait Dominus, qui narraverunt ea et seduxerunt populum meum in mendaciis suis et in iactantia sua, cum ego non misissem eos nec mandassem eis; qui nihil profuerunt populo huic, dicit Dominus.
JER|23|33|Si interrogaverit te populus iste vel propheta aut sacerdos dicens: Quod est onus Domini", dices ad eos: Vos estis onus; proiciam quippe vos, dicit Dominus.
JER|23|34|Et propheta et sacerdos et populus, qui dicit: "Onus Domini", visitabo super virum illum et super domum eius.
JER|23|35|Haec dicetis unusquisque ad proximum et ad fratrem suum: "Quid respondit Dominus?" et "Quid locutus est Dominus?".
JER|23|36|Sed "Onus Domini" ultra non memorabitis, quia onus erit unicuique sermo suus, et pervertitis verba Dei viventis, Domini exercituum, Dei nostri.
JER|23|37|Haec dices ad prophetam: "Quid respondit tibi Dominus?" et "Quid locutus est Dominus?".
JER|23|38|Si autem "Onus Domini" dixeritis, propter hoc haec dicit Dominus: Quia dixistis sermonem istum: "Onus Domini", et misi ad vos dicens: Nolite dicere: "Onus Domini";
JER|23|39|propterea, ecce ego tollam vos portans et proiciam vos et civitatem, quam dedi vobis et patribus vestris, a facie mea;
JER|23|40|et dabo vos in opprobrium sempiternum et in ignominiam aeternam, quae numquam oblivione delebitur ".
JER|24|1|Ostendit mihi Dominus, et ecce duo calathi pleni ficis positi ante templum Domini, postquam transtulit Nabuchodonosor rex Babylonis Iechoniam filium Ioachim regem Iudae et principes eius et fabrum et inclusorem de Ierusalem et adduxit eos in Babylonem.
JER|24|2|Calathus unus ficus bonas habebat nimis, ut solent ficus esse primi temporis; et calathus unus ficus habebat malas nimis, quae comedi non poterant, eo quod essent malae.
JER|24|3|Et dixit Dominus ad me: " Quid tu vides, Ieremia? ". Et dixi: " Ficus, ficus bonas, bonas valde, et malas, malas valde, quae comedi non possunt, eo quod sint malae ".
JER|24|4|Et factum est verbum Domini ad me dicens:
JER|24|5|" Haec dicit Dominus, Deus Israel: Sicut ficus hae bonae, sic cognoscam transmigrationem Iudae, quam emisi de loco isto in terram Chaldaeorum, in bonum.
JER|24|6|Et ponam oculos meos super eos ad placandum et reducam eos in terram hanc et aedificabo eos et non destruam et plantabo eos et non evellam.
JER|24|7|Et dabo eis cor, ut sciant me quia ego sum Dominus; et erunt mihi in populum, et ego ero eis in Deum, quia revertentur ad me in toto corde suo.
JER|24|8|Et sicut ficus pessimae, quae comedi non possunt, eo quod sint malae, haec dicit Dominus, sic dabo Sedeciam regem Iudae et principes eius et reliquos de Ierusalem, qui remanserunt in terra hac et qui habitant in terra Aegypti.
JER|24|9|Et dabo eos in vexationem afflictionemque omnibus regnis terrae, in opprobrium et in proverbium et in derisum et in maledictionem in universis locis, ad quae eieci eos.
JER|24|10|Et mittam in eis gladium et famem et pestem, donec consumantur de terra, quam dedi eis et patribus eorum ".
JER|25|1|Verbum, quod factum est ad Ieremiam de omni populo Iudae in anno quarto Ioachim filii Iosiae regis Iudae - ipse est annus primus Nabuchodonosor regis Babylonis -
JER|25|2|quod locutus est Ieremias propheta ad omnem populum Iudae et ad universos habitatores Ierusalem dicens:
JER|25|3|" A tertio decimo anno Iosiae filii Amon regis Iudae usque ad diem hanc, iste tertius et vicesimus est annus, factum est verbum Domini ad me, et locutus sum ad vos de nocte consurgens et loquens, et non audistis.
JER|25|4|Et misit Dominus ad vos omnes servos suos prophetas, consurgens diluculo mittensque; et non audistis neque inclinastis aures vestras, ut audiretis,
JER|25|5|cum diceret: "Revertimini unusquisque a via sua mala et a pessimis cogitationibus vestris, et habitabitis in terra, quam dedit Dominus vobis et patribus vestris, a saeculo et usque in saeculum;
JER|25|6|et nolite ire post deos alienos, ut serviatis eis adoretisque eos, neque me ad iracundiam provocetis in operibus manuum vestrarum, et non affligam vos.
JER|25|7|Et non audistis me, dicit Dominus, ut me ad iracundiam provocaretis in operibus manuum vestrarum, in malum vestrum".
JER|25|8|Propterea haec dicit Dominus exercituum: Pro eo quod non audistis verba mea,
JER|25|9|ecce ego mittam et assumam universas cognationes aquilonis, ait Dominus, et Nabuchodonosor regem Babylonis, servum meum, et adducam eos super terram istam et super habitatores eius et super omnes nationes, quae in circuitu illius sunt; et interficiam eos et ponam eos in stuporem et in sibilum et in ruinas sempiternas.
JER|25|10|Perdamque ex eis vocem gaudii et vocem laetitiae, vocem sponsi et vocem sponsae, vocem molae et lumen lucernae,
JER|25|11|et erit universa terra haec in solitudinem et in stuporem, et servient omnes gentes istae regi Babylonis septuaginta annis.
JER|25|12|Cumque impleti fuerint septuaginta anni, visitabo super regem Babylonis et super gentem illam, dicit Dominus, iniquitatem eorum et super terram Chaldaeorum; et ponam illam in solitudines sempiternas.
JER|25|13|Et adducam super terram illam omnia verba mea, quae locutus sum contra eam, omne, quod scriptum est in libro isto, quaecumque prophetavit Ieremias adversum omnes gentes.
JER|25|14|Quia servient eis etiam illi, gentes multae et reges magni, et reddam eis secundum opera eorum et secundum facta manuum suarum ".
JER|25|15|Quia sic dicit Dominus, Deus Israel, ad me: " Sume calicem vini furoris huius de manu mea et propinabis de illo cunctis gentibus, ad quas ego mittam te;
JER|25|16|et bibent et turbabuntur et insanient a facie gladii, quem ego mittam inter eos ".
JER|25|17|Et accepi calicem de manu Domini et propinavi cunctis gentibus, ad quas misit me Dominus,
JER|25|18|Ierusalem et civitatibus Iudae et regibus eius et principibus eius, ut darem eos in solitudinem et in stuporem, in sibilum et in maledictionem, sicut est dies ista;
JER|25|19|pharaoni regi Aegypti et servis eius et principibus eius et omni populo eius;
JER|25|20|et omni vulgo promiscuo et cunctis regibus terrae Us et cunctis regibus terrae Philisthim et Ascaloni et Gazae et Accaroni et reliquiis Azoti,
JER|25|21|Edom et Moab et filiis Ammon;
JER|25|22|et cunctis regibus Tyri et universis regibus Sidonis et regibus terrae insularum, qui sunt trans mare;
JER|25|23|et Dedan et Thema et Buz et universis, qui attonsi sunt in comam;
JER|25|24|et cunctis regibus Arabiae et cunctis regibus vulgi promiscui, qui habitant in deserto,
JER|25|25|et cunctis regibus Zimri et cunctis regibus Elam et cunctis regibus Medorum,
JER|25|26|cunctis quoque regibus aquilonis de prope et de longe, unicuique post fratrem suum et omnibus regnis terrae, quae super faciem eius sunt; et rex Sesach bibet post eos.
JER|25|27|" Et dices ad eos: Haec dicit Dominus exercituum, Deus Israel: Bibite et inebriamini et vomite; et cadite neque surgatis a facie gladii, quem ego mittam inter vos.
JER|25|28|Cumque noluerint accipere calicem de manu tua, ut bibant, dices ad eos: Haec dicit Dominus exercituum: Bibentes bibetis;
JER|25|29|quia ecce in civitate, super quam invocatum est nomen meum, ego incipio affligere, et vos immunes eritis? Non eritis immunes; gladium enim ego voco super omnes habitatores terrae, dicit Dominus exercituum.
JER|25|30|Et tu prophetabis ad eos omnia verba haec et dices ad illos:Dominus de excelso rugietet de habitaculo sancto suo dabit vocem suam;rugiens rugiet super pascua sua,celeuma quasi calcantium concineturadversus omnes habitatores terrae.
JER|25|31|Pervenit sonitus usque ad extrema terrae,quia iudicium Domino cum gentibus;in iudicium venit ipse cum omni carne;impios tradidit gladio,dicit Dominus.
JER|25|32|Haec dicit Dominus exercituum:Ecce afflictio egreditur de gente in gentem,et turbo magnus surgit a summitatibus terrae ".
JER|25|33|Et erunt interfecti Domini in die illa a summo terrae usque ad summum eius; non plangentur et non colligentur neque sepelientur: in sterquilinium super faciem terrae erunt.
JER|25|34|Ululate, pastores, et clamate;et volutamini vos in pulvere, optimates gregis,quia completi sunt dies vestri ad occisionemet ad dispersionem vestram,et cadetis quasi vasa pretiosa.
JER|25|35|Et peribit fuga a pastoribus,et salvatio ab optimatibus gregis.
JER|25|36|Vox clamoris pastorumet ululatus optimatium gregis,quia vastavit Dominus pascua eorum.
JER|25|37|Et conticuerunt arva pacisa facie irae furoris Domini.
JER|25|38|Dereliquit quasi leo umbraculum suum,quia facta est terra eorum in desolationem,a facie irae violentaeet a facie irae furoris Domini.
JER|26|1|In principio regni Ioachim filii Iosiae regis Iudae factum est verbum istud a Domino dicens:
JER|26|2|" Haec dicit Dominus: Sta in atrio domus Domini et loqueris ad omnes civitates Iudae, de quibus veniunt, ut adorent in domo Domini, universos sermones, quos ego mandavi tibi, ut loquaris ad eos: noli subtrahere verbum,
JER|26|3|si forte audiant et convertantur unusquisque a via sua mala, et paeniteat me mali, quod cogito facere eis propter malitiam operum eorum.
JER|26|4|Et dices ad eos: Haec dicit Dominus: Si non audieritis me, ut ambuletis in lege mea, quam dedi vobis,
JER|26|5|ut audiatis sermones servorum meorum prophetarum, quos ego misi ad vos de nocte consurgens et dirigens, et non audistis,
JER|26|6|dabo domum istam sicut Silo et urbem hanc dabo in maledictionem cunctis gentibus terrae ".
JER|26|7|Et audierunt sacerdotes et prophetae et omnis populus Ieremiam loquentem verba haec in domo Domini.
JER|26|8|Cumque complesset Ieremias loquens omnia, quae praeceperat ei Dominus, ut loqueretur ad universum populum, apprehenderunt eum sacerdotes et prophetae et omnis populus dicens: " Morte moriaris!
JER|26|9|Quare prophetasti in nomine Domini dicens: "Sicut Silo erit domus haec, et urbs ista desolabitur, eo quod non sit habitator"? ".Et congregatus est omnis populus adversus Ieremiam in domo Domini.
JER|26|10|Et audierunt principes Iudae verba haec et ascenderunt de domo regis in domum Domini et sederunt in introitu portae domus Domini Novae.
JER|26|11|Et locuti sunt sacerdotes et prophetae ad principes et ad omnem populum dicentes: " Iudicium mortis est viro huic, quia prophetavit adversus civitatem istam, sicut audistis auribus vestris ".
JER|26|12|Et ait Ieremias ad omnes principes et ad universum populum dicens: " Dominus misit me, ut prophetarem ad domum istam et ad civitatem hanc omnia verba, quae audistis.
JER|26|13|Nunc ergo bonas facite vias vestras et opera vestra et audite vocem Domini Dei vestri, et paenitebit Dominum mali, quod locutus est adversum vos.
JER|26|14|Ego autem ecce in manibus vestris sum; facite mihi, quod bonum et rectum est in oculis vestris.
JER|26|15|Verumtamen scitote et cognoscite quod si occideritis me, sanguinem innocentem tradetis contra vosmetipsos et contra civitatem istam et habitatores eius; in veritate enim misit me Dominus ad vos, ut loquerer in auribus vestris omnia verba haec ".
JER|26|16|Et dixerunt principes et omnis populus ad sacerdotes et prophetas: " Non est viro huic iudicium mortis, quia in nomine Domini Dei nostri locutus est ad nos ".
JER|26|17|Surrexerunt ergo viri de senioribus terrae et dixerunt ad omnem coetum populi loquentes:
JER|26|18|" Michaeas Morasthites fuit propheta in diebus Ezechiae regis Iudae et ait ad omnem populum Iudae dicens: "Haec dicit Dominus exercituum:Sion quasi ager arabitur,et Ierusalem in acervum lapidum erit,et mons domus in excelsa silvarum".
JER|26|19|Numquid morte condemnavit eum Ezechias rex Iudae et omnis Iuda? Numquid non timuerunt Dominum et deprecati sunt faciem Domini, et paenituit Dominum mali, quod locutus fuerat adversum eos? Et nos facimus malum grande contra animas nostras! ".
JER|26|20|Fuit quoque vir prophetans in nomine Domini Urias filius Semei de Cariathiarim et prophetavit adversus civitatem istam et adversus terram hanc iuxta omnia verba Ieremiae.
JER|26|21|Et audivit rex Ioachim et omnes potentes et principes eius verba haec, et quaesivit rex interficere eum; et audivit Urias et timuit fugitque et ingressus est Aegyptum.
JER|26|22|Et misit rex Ioachim viros in Aegyptum, Elnathan filium Achobor et viros cum eo in Aegyptum;
JER|26|23|et eduxerunt Uriam de Aegypto et adduxerunt eum ad regem Ioachim, et percussit eum gladio et proiecit cadaver eius in sepulcris filiorum vulgi.
JER|26|24|Igitur manus Ahicam filii Saphan fuit cum Ieremia, ut non traderetur in manus populi, et interficerent eum.
JER|27|1|In principio regni Sedeciae filii Iosiae regis Iudae factum est verbum istud ad Ieremiam a Domino dicens:
JER|27|2|" Haec dicit Dominus ad me: Fac tibi vincula et iuga et pones ea in collo tuo
JER|27|3|et mittes ea ad regem Edom et ad regem Moab et ad regem filiorum Ammon et ad regem Tyri et ad regem Sidonis in manu nuntiorum, qui venerunt Ierusalem ad Sedeciam regem Iudae;
JER|27|4|et praecipies eis, ut ad dominos suos loquantur: Haec dicit Dominus exercituum, Deus Israel: Haec dicetis ad dominos vestros:
JER|27|5|Ego feci terram et hominem et iumenta, quae sunt super faciem terrae, in fortitudine mea magna et in brachio meo extento et dedi eam ei, qui placuit in oculis meis.
JER|27|6|Et nunc itaque ego dedi omnes terras istas in manu Nabuchodonosor regis Babylonis servi mei, insuper et bestias agri dedi ei, ut serviant illi;
JER|27|7|et servient ei omnes gentes et filio eius et filio filii eius, donec veniat tempus terrae eius etiam ipsius; et servient ei gentes multae et reges magni.
JER|27|8|Gens autem et regnum, quod non servierit Nabuchodonosor regi Babylonis, et quicumque non curvaverit collum suum sub iugo regis Babylonis, in gladio et in fame et in peste visitabo super gentem illam, ait Dominus, donec consumam eos in manu eius.
JER|27|9|Vos ergo nolite audire prophetas vestros et divinos et somniatores et augures et maleficos, qui dicunt vobis: "Non servietis regi Babylonis",
JER|27|10|quia mendacium prophetant vobis, ut longe vos faciant de terra vestra, et eiciam vos, et pereatis.
JER|27|11|Porro gens, quae subiecerit cervicem suam sub iugo regis Babylonis et servierit ei, dimittam eam in terra sua, dicit Dominus, et colet eam et habitabit in ea ".
JER|27|12|Et ad Sedeciam regem Iudae locutus sum secundum omnia verba haec dicens: " Subicite colla vestra sub iugo regis Babylonis et servite ei et populo eius, et vivetis.
JER|27|13|Quare moriemini tu et populus tuus gladio, fame et peste, sicut locutus est Dominus ad gentem, quae servire noluerit regi Babylonis?
JER|27|14|Nolite audire verba prophetarum dicentium vobis: "Non servietis regi Babylonis", quia mendacium ipsi loquuntur vobis.
JER|27|15|Quia non misi eos, ait Dominus, et ipsi prophetant in nomine meo mendaciter, ut eiciam vos et pereatis, tam vos quam prophetae, qui vaticinantur vobis ".
JER|27|16|Et ad sacerdotes et ad populum istum locutus sum dicens: " Haec dicit Dominus: Nolite audire verba prophetarum vestrorum, qui prophetant vobis dicentes: "Ecce vasa domus Domini revertentur de Babylone nunc cito". Mendacium enim prophetant vobis.
JER|27|17|Nolite ergo audire eos, sed servite regi Babylonis, ut vivatis. Quare datur haec civitas in solitudinem?
JER|27|18|Et si prophetae sunt, et est verbum Domini in eis, occurrant Domino exercituum, ut non veniant vasa, quae derelicta fuerant in domo Domini et in domo regis Iudae et in Ierusalem, in Babylonem ".
JER|27|19|Quia haec dicit Dominus exercituum ad columnas et ad mare et ad bases et ad reliqua vasorum, quae remanserunt in civitate hac,
JER|27|20|quae non tulit Nabuchodonosor rex Babylonis, cum transferret Iechoniam filium Ioachim regem Iudae de Ierusalem in Babylonem et omnes optimates Iudae et Ierusalem;
JER|27|21|quia haec dicit Dominus exercituum, Deus Israel, ad vasa, quae derelicta sunt in domo Domini et in domo regis Iudae et Ierusalem:
JER|27|22|"In Babylonem transferentur et ibi erunt usque ad diem visitationis eorum, dicit Dominus; et afferri faciam ea et restitui in loco isto ".
JER|28|1|Et factum est in anno illo, in principio regni Sedeciae regis Iudae, in anno quarto in mense quinto, dixit ad me Hananias filius Azur propheta de Gabaon in domo Domini coram sacerdotibus et omni populo dicens:
JER|28|2|" Haec dicit Domi nus exercituum, Deus Israel: Contrivi iugum regis Babylonis.
JER|28|3|Adhuc duo anni dierum, et ego referri faciam ad locum istum omnia vasa domus Domini, quae tulit Nabuchodonosor rex Babylonis de loco isto et transtulit ea in Babylonem.
JER|28|4|Et Iechoniam filium Ioachim regem Iudae et omnem transmigrationem Iudae, qui ingressi sunt in Babylonem, ego convertam ad locum istum, ait Dominus; conteram enim iugum regis Babylonis ".
JER|28|5|Et dixit Ieremias propheta ad Hananiam prophetam in oculis sacerdotum et in oculis omnis populi, qui stabat in domo Domini,
JER|28|6|et ait Ieremias propheta: " Amen, sic faciat Dominus! Suscitet Dominus verba tua, quae prophetasti, ut referantur vasa in domum Domini et omnis transmigratio de Babylone ad locum istum.
JER|28|7|Verumtamen audi verbum hoc, quod ego loquor in auribus tuis et in auribus universi populi:
JER|28|8|Prophetae, qui fuerunt ante me et ante te ab initio et prophetaverunt super terras multas et super regna magna de proelio et de afflictione et de peste;
JER|28|9|propheta, qui vaticinatur pacem, cum venerit verbum eius, scietur propheta, quem misit Dominus in veritate ".
JER|28|10|Et tulit Hananias propheta iugum de collo Ieremiae prophetae et confregit illud;
JER|28|11|et ait Hananias in conspectu omnis populi dicens: " Haec dicit Dominus: Sic confringam iugum Nabuchodonosor regis Babylonis post duos annos dierum de collo omnium gentium ". Et abiit Ieremias propheta in viam suam.
JER|28|12|Et factum est verbum Domini ad Ieremiam, postquam confregit Hananias propheta iugum de collo Ieremiae prophetae, dicens:
JER|28|13|"Vade et dices Hananiae: Haec dicit Dominus: Iuga lignea contrivisti et facies pro eis iuga ferrea.
JER|28|14|Quia haec dicit Dominus exercituum, Deus Israel: Iugum ferreum posui super collum cunctarum gentium istarum, ut serviant Nabuchodonosor regi Babylonis, et servient ei; insuper et bestias terrae dedi ei ".
JER|28|15|Et dixit Ieremias propheta ad Hananiam prophetam: "Audi, Hanania! Non misit te Dominus, et tu confidere fecisti populum istum in mendacio.
JER|28|16|Idcirco haec dicit Dominus: Ecce emittam te a facie terrae; hoc anno morieris, adversum enim Dominum praevaricationem locutus es ".
JER|28|17|Et mortuus est Hananias propheta in anno illo, mense septimo.
JER|29|1|Et haec sunt verba epistulae, quam misit Ieremias propheta de Ierusalem ad reliquias seniorum transmigrationis et ad sacerdotes et ad prophetas et ad omnem populum, quem traduxerat Nabuchodonosor de Ierusalem in Babylonem,
JER|29|2|postquam egressus est Iechonias rex et domina et eunuchi et principes Iudae et Ierusalem et faber et inclusor de Ierusalem,
JER|29|3|in manu Elasa filii Saphan et Gamariae filii Helciae, quos misit Sedecias rex Iudae ad Nabuchodonosor regem Babylonis in Babylonem dicens:
JER|29|4|" Haec dicit Dominus exercituum, Deus Israel, omni transmigrationi, quam transtuli de Ierusalem in Babylonem:
JER|29|5|Aedificate domos et habitate et plantate hortos et comedite fructum eorum,
JER|29|6|accipite uxores et generate filios et filias et date filiis vestris uxores et filias vestras date viris, et pariant filios et filias, et multiplicamini ibi et nolite esse pauci numero.
JER|29|7|Et quaerite pacem civitatis, ad quam transmigrare vos feci, et orate pro ea ad Dominum, quia in pace illius erit pax vobis.
JER|29|8|Haec enim dicit Dominus exercituum, Deus Israel: Non vos seducant prophetae vestri, qui sunt in medio vestrum, et divini vestri, et ne attendatis ad somnia vestra, quae vos somniatis,
JER|29|9|quia falso ipsi prophetant vobis in nomine meo, et non misi eos, dicit Dominus.
JER|29|10|Quia haec dicit Dominus: Cum impleti fuerint in Babylone septuaginta anni, visitabo vos et suscitabo super vos verbum meum bonum, ut reducam vos ad locum istum.
JER|29|11|Ego enim scio cogitationes, quas ego cogito super vos, ait Dominus, cogitationes pacis et non afflictionis, ut dem vobis posteritatem et spem.
JER|29|12|Et invocabitis me et ibitis; et orabitis me, et ego exaudiam vos.
JER|29|13|Quaeretis me et invenietis, cum quaesieritis me in toto corde vestro.
JER|29|14|Et inveniar a vobis, ait Dominus, et reducam captivitatem vestram et congregabo vos de universis gentibus et de cunctis locis, ad quae expuli vos, dicit Dominus; et reverti vos faciam ad locum, de quo transmigrare vos feci.
JER|29|15|Quia dixistis: "Suscitavit nobis Dominus prophetas in Babylone".
JER|29|16|Quia haec dicit Dominus ad regem, qui sedet super solium David, et ad omnem populum habitatorem urbis huius, ad fratres vestros, qui non sunt egressi vobiscum in transmigrationem,
JER|29|17|haec dicit Dominus exercituum: Ecce mittam in eis gladium et famem et pestem et ponam eos quasi ficus malas, quae comedi non possunt, eo quod pessimae sint;
JER|29|18|et persequar eos in gladio et in fame et in pestilentia et dabo eos in vexationem universis regnis terrae, in maledictionem et in stuporem et in sibilum et in opprobrium cunctis gentibus, ad quas ego eieci eos,
JER|29|19|eo quod non audierint verba mea, dicit Dominus, quae misi ad eos per servos meos prophetas, de nocte consurgens et mittens, et non audistis, dicit Dominus.
JER|29|20|Vos ergo audite verbum Domini, omnis transmigratio, quam emisi de Ierusalem in Babylonem.
JER|29|21|Haec dicit Dominus exercituum, Deus Israel, ad Achab filium Colaiae et ad Sedeciam filium Maasiae, qui prophetant vobis in nomine meo mendaciter: Ecce ego tradam eos in manu Nabuchodonosor regis Babylonis, et percutiet eos in oculis vestris;
JER|29|22|et assumetur ex eis maledictio omni transmigrationi Iudae, quae est in Babylone, dicentium: "Ponat te Dominus sicut Sedeciam et sicut Achab, quos frixit rex Babylonis in igne!";
JER|29|23|pro eo quod fecerint stultitiam in Israel et moechati sunt in uxores amicorum suorum et locuti sunt verbum in nomine meo mendaciter, quod non mandavi eis. Ego enim scio et sum testis, dicit Dominus.
JER|29|24|Et ad Semeiam Nehelamiten dices:
JER|29|25|Haec dicit Dominus exercituum, Deus Israel, pro eo quod misisti in nomine tuo epistulas ad omnem populum, qui est in Ierusalem, et ad Sophoniam filium Maasiae sacerdotem et ad universos sacerdotes dicens:
JER|29|26|"Dominus dedit te sacerdotem pro Ioiada sacerdote, ut sis praefectus in domo Domini super omnem virum arrepticium et prophetantem, ut mittas eum in nervum et in vincula.
JER|29|27|Et nunc quare non increpasti Ieremiam Anathothiten, qui prophetat vobis?
JER|29|28|Quia super hoc misit ad nos in Babylonem dicens: Longum est; aedificate domos et habitate et plantate hortos et comedite fructum eorum" ".
JER|29|29|Legit ergo Sophonias sacerdos epistulam istam in auribus Ieremiae prophetae.
JER|29|30|Et factum est verbum Domini ad Ieremiam dicens:
JER|29|31|" Mitte ad omnem transmigrationem dicens: Haec dicit Dominus ad Semeiam Nehelamiten: Pro eo quod prophetavit vobis Semeias, et ego non misi eum, et fecit vos confidere in mendacio,
JER|29|32|idcirco haec dicit Dominus: Ecce ego visitabo super Semeiam Nehelamiten et super semen eius; non erit ei vir sedens in medio populi huius, et non videbit bonum, quod ego faciam populo meo, ait Dominus, quia praevaricationem locutus est adversus Dominum ".
JER|30|1|Verbum, quod factum est ad Ieremiam a Domino dicens:
JER|30|2|" Haec dicit Dominus, Deus Israel, dicens: Scribe tibi omnia verba, quae locutus sum ad te, in libro;
JER|30|3|ecce enim dies veniunt, dicit Dominus, et convertam sortem populi mei Israel et Iudae, ait Dominus, et convertam eos ad terram, quam dedi patribus eorum, et possidebunt eam ".
JER|30|4|Et haec verba, quae locutus est Dominus ad Israel et ad Iudam:
JER|30|5|" Quoniam haec dicit Dominus:Vocem terroris audivimus,formido et non est pax.
JER|30|6|Interrogate et videte, si generat masculus;quare ergo vidi omnis viri manumsuper lumbum suum quasi parturientis,et conversae sunt universae facies in auruginem?
JER|30|7|Vae, quia magna dies illa,nec est similis eius,tempusque tribulationis est Iacob,et ex ipso salvabitur.
JER|30|8|Et erit: in die illa, ait Dominus exercituum, conteram iugum eius de collo tuo et vincula tua dirumpam; et non dominabuntur ei amplius alieni,
JER|30|9|sed servient Domino Deo suo et David regi suo, quem suscitabo eis.
JER|30|10|Tu ergo ne timeas, serve meus Iacob,ait Dominus,neque paveas, Israel,quia ecce ego salvabo te de terra longinquaet semen tuum de terra captivitatis eorum;et revertetur Iacob et quiescetet securus erit, et non erit quem formidet;
JER|30|11|quoniam tecum ego sum,ait Dominus,ut salvem te.Faciam enim consummationem in cunctis gentibus,in quibus dispersi te;te autem non faciam in consummationem,sed castigabo te in iudicionec quasi innocenti parcam tibi.
JER|30|12|Quia haec dicit Dominus:Insanabilis fractura tua,pessima plaga tua;
JER|30|13|non est qui iudicet iudicium tuum;sunt ulceri medicamina,tibi vero cicatrix non obducitur.
JER|30|14|Omnes amatores tui obliti sunt tui,te non quaerunt;plaga enim inimici percussi tecastigatione crudeli:propter multitudinem iniquitatis tuaedura facta sunt peccata tua.
JER|30|15|Quid clamas super contritione tua?Insanabilis est dolor tuus.Propter multitudinem iniquitatis tuaeet propter dura peccata tua feci haec tibi.
JER|30|16|Propterea omnes, qui comedunt te, devorabuntur,et universi hostes tui in captivitatem ducentur,et, qui te vastant, vastabuntur,cunctosque praedatores tuos dabo in praedam.
JER|30|17|Obducam enim cicatricem tibiet a vulneribus tuis sanabo te,dicit Dominus,quia Eiectam vocaverunt te,Sion haec, quae non habebat requirentem.
JER|30|18|Haec dicit Dominus:Ecce ego convertam sortem tabernaculorum Iacobet tectis eius miserebor,et aedificabitur civitas in ruinis suis,et arx in loco suo fundabitur;
JER|30|19|et egredietur de eis laus voxque ludentium.Et multiplicabo eos, et non imminuentur,et glorificabo eos, et non attenuabuntur.
JER|30|20|Et erunt filii eius sicut a principio,et coetus eius coram me permanebit,et visitabo adversum omnes, qui tribulant eum.
JER|30|21|Et erit dux eius ex eo,et princeps de medio eius procedet; et applicabo eum, et accedet ad me.Quis enim iste est, qui pignori dabit cor suum,ut appropinquet mihi?,ait Dominus.
JER|30|22|Et eritis mihi in populum,et ego ero vobis in Deum.
JER|30|23|Ecce turbo Domini, furor egrediens,procella ruens;in capite impiorum conquiescet.
JER|30|24|Non cessabit ab ira indignationis Dominus,donec faciat et compleatcogitationes cordis sui;in novissimo dierum intellegetis ea.
JER|31|1|In tempore illo,dicit Dominus,ero Deus universis cognationibus Israel,et ipsi erunt mihi in populum.
JER|31|2|Haec dicit Dominus:Invenit gratiam in desertopopulus, qui remanserat a gladio;vadet ad requiem suam Israel ".
JER|31|3|De longe Dominus apparuit mihi: In caritate perpetua dilexi te;ideo attraxi te in misericordia.
JER|31|4|Rursumque aedificabo te, et aedificaberis,virgo Israel;adhuc ornaberis tympanis tuiset egredieris in choro ludentium.
JER|31|5|Adhuc plantabis vineas in montibus Samariae;plantabunt plantanteset vindemiabunt.
JER|31|6|Quia erit dies, in qua clamabunt custodesin monte Ephraim:Surgite, et ascendamus in Sionad Dominum Deum nostrum".
JER|31|7|Quia haec dicit Dominus:Exsultate in laetitia propter Iacobet hinnite capiti gentium;personate, canite et dicite:Salva, Domine, populum tuum,reliquias Israel".
JER|31|8|Ecce ego adducam eos de terra aquiloniset congregabo eos ab extremis terrae;inter quos erunt caecus et claudus, praegnans et pariens simul:coetus magnus revertentium huc.
JER|31|9|In fletu venient,et in deprecatione reducam eoset adducam eos per torrentes aquarumin via recta, et non impingent in ea, quia factus sum Israeli pater,et Ephraim primogenitus meus est ".
JER|31|10|Audite verbum Domini, gentes,et annuntiate in insulis, quae procul sunt, et dicite: Qui dispersit Israel, congregabit eumet custodiet eum sicut pastor gregem suum ".
JER|31|11|Redemit enim Dominus Iacobet liberavit eum de manu potentioris.
JER|31|12|Et venient et laudabunt in monte Sionet confluent ad bona Dominisuper frumento et vino et oleoet fetu pecorum et armentorum;eritque anima eorum quasi hortus irriguus,et ultra non esurient.
JER|31|13|Tunc laetabitur virgo in choro,iuvenes et senes simul. Et convertam luctum eorum in gaudiumet consolabor eos et laetificabo a dolore suo.
JER|31|14|Et inebriabo animam sacerdotum pinguedine,et populus meus bonis meis adimplebitur ",ait Dominus.
JER|31|15|Haec dicit Dominus: Vox in Rama audita estlamentationis, luctus et fletusRachel plorantis filios suoset nolentis consolari super eis, quia non sunt ".
JER|31|16|Haec dicit Dominus: Quiescat vox tua a ploratu,et oculi tui a lacrimis,quia est merces operi tuo,ait Dominus,et revertentur de terra inimici.
JER|31|17|Et est spes novissimis tuis,ait Dominus,et revertentur filii ad terminos suos.
JER|31|18|Audiens audivi Ephraim transmigrantem:Castigasti me, et eruditus sumquasi iuvenculus indomitus;converte me, et convertar,quia tu Dominus Deus meus.
JER|31|19|Postquam enim convertisti me,egi paenitentiam;et postquam ostendisti mihi,percussi femur meum;confusus sum et erubui,quoniam sustinui opprobrium adulescentiae meae".
JER|31|20|Estne filius honorabilis mihi Ephraimaut puer delectabilis,quia ex quo locutus sum de eo,adhuc recordabor eius?Idcirco conturbata sunt viscera mea super eum:miserans miserebor eius ",ait Dominus.
JER|31|21|Statue tibi lapides,pone tibi signa,dirige cor tuum in iter,viam, in qua ambulasti;revertere, virgo Israel,revertere ad civitates tuas istas.
JER|31|22|Usquequo vagaberis,filia rebellis?Quia creavit Dominus novum super terram:femina circumdabit virum.
JER|31|23|Haec dicit Dominus exercituum, Deus Israel: " Adhuc dicent verbum istud in terra Iudae et in urbibus eius, cum convertero sortem eorum: "Benedicat tibi Dominus, habitaculum iustitiae, mons sanctus".
JER|31|24|Et habitabunt in eo Iudas et omnes civitates eius simul, agricolae et minantes greges.
JER|31|25|Quia inebriavi animam lassam et omnem animam esurientem saturavi ".
JER|31|26|Ideo quasi de somno suscitatus sum et vidi, et somnus meus dulcis mihi.
JER|31|27|" Ecce dies veniunt, dicit Dominus, et seminabo domum Israel et domum Iudae semine hominum et semine iumentorum.
JER|31|28|Et sicut vigilavi super eos, ut evellerem et demolirer et dissiparem et disperderem et affligerem, sic vigilabo super eos, ut aedificem et plantem, ait Dominus.
JER|31|29|In diebus illis non dicent ultra:Patres comederunt uvam acerbam, et dentes filiorum obstupuerunt",
JER|31|30|sed unusquisque in iniquitate sua morietur; omnis homo, qui comederit uvam acerbam, obstupescent dentes eius.
JER|31|31|Ecce dies veniunt, dicit Dominus, et feriam domui Israel et domui Iudae pactum novum;
JER|31|32|non secundum pactum, quod pepigi cum patribus eorum in die qua apprehendi manum eorum, ut educerem eos de terra Aegypti, pactum, quod irritum fecerunt, et ego dominatus sum eorum, dicit Dominus.
JER|31|33|Sed hoc erit pactum, quod feriam cum domo Israel post dies illos, dicit Dominus: Dabo legem meam in visceribus eorum et in corde eorum scribam eam; et ero eis in Deum, et ipsi erunt mihi in populum.
JER|31|34|Et non docebit ultra vir proximum suum, et vir fratrem suum dicens: Cognosce Dominum"; omnes enim cognoscent me, a minimo eorum usque ad maximum, ait Dominus, quia propitiabor iniquitati eorum et peccati eorum non memorabor amplius ".
JER|31|35|Haec dicit Dominus,qui dat solem in lumine diei,ordinem lunae et stellarum in lumine noctis,qui turbat mare, et fremunt fluctus eius,Dominus exercituum nomen illi:
JER|31|36|" Si defecerint leges istae coram me,dicit Dominus,tunc et semen Israel deficiet,ut non sit gens coram me cunctis diebus ".
JER|31|37|Haec dicit Dominus: Si mensurari potuerint caeli sursum,et investigari fundamenta terrae deorsum,et ego abiciam universum semen Israelpropter omnia, quae fecerunt,dicit Dominus.
JER|31|38|Ecce dies veniunt, dicit Dominus, et aedificabitur civitas Domino a turre Hananeel usque ad portam Anguli,
JER|31|39|et exibit ultra norma mensurae in conspectu eius super collem Gareb et vertetur in Goa,
JER|31|40|et omnis vallis cadaverum et cineris et universa regio usque ad torrentem Cedron et usque ad angulum portae Equorum orientalis sanctum Domini; non evelletur et non destruetur ultra in perpetuum ".
JER|32|1|Verbum, quod factum est ad Ieremiam a Domino in anno decimo Sedeciae regis Iudae; ipse est annus decimus octavus Nabuchodonosor.
JER|32|2|Tunc exercitus regis Babylonis obsidebat Ierusalem, et Ieremias propheta erat clausus in atrio custodiae, qui erat in domo regis Iudae.
JER|32|3|Clauserat enim eum Sedecias rex Iudae dicens: " Quare vaticinaris dicens: "Haec dicit Dominus: Ecce ego dabo civitatem istam in manu regis Babylonis, et capiet eam;
JER|32|4|et Sedecias rex Iudae non effugiet de manu Chaldaeorum, sed tradetur in manus regis Babylonis, et loquetur os eius cum ore illius, et oculi eius oculos illius videbunt;
JER|32|5|et in Babylonem ducet Sedeciam, et ibi erit, donec visitem eum, ait Dominus; si autem dimicaveritis adversum Chaldaeos, nihil prosperum habebitis"? ".
JER|32|6|Et dixit Ieremias: " Factum est verbum Domini ad me dicens:
JER|32|7|Ecce Hanameel filius Sellum patruelis tuus veniet ad te dicens: "Eme tibi agrum meum, qui est in Anathoth; tibi enim competit ex propinquitate, ut emas".
JER|32|8|Et venit ad me Hanameel filius patrui mei secundum verbum Domini ad vestibulum custodiae et ait ad me: "Posside agrum meum, qui est in Anathoth in terra Beniamin, quia tibi competit hereditas, et tu propinquus es, ut possideas". Intellexi autem quod verbum Domini esset
JER|32|9|et emi agrum ab Hanameel filio patrui mei, qui est in Anathoth, et appendi ei argentum: septem et decem siclos argenteos.
JER|32|10|Et scripsi in libro et signavi et adhibui testes et appendi argentum in statera.
JER|32|11|Et accepi librum possessionis signatum, continentem stipulationes et rata, et apertum;
JER|32|12|et dedi librum possessionis Baruch filio Neriae filii Maasiae in oculis Hanameel patruelis mei et in oculis testium, qui obsignaverant in libro emptionis, et in oculis omnium Iudaeorum, qui sedebant in atrio custodiae.
JER|32|13|Et praecepi Baruch coram eis dicens:
JER|32|14|Haec dicit Dominus exercituum, Deus Israel: Sume libros istos, librum emptionis hunc signatum et librum hunc, qui apertus est; et pones illos in vase fictili, ut permanere possint diebus multis.
JER|32|15|Haec enim dicit Dominus exercituum, Deus Israel: Adhuc possidebuntur domus et agri et vineae in terra ista.
JER|32|16|Et oravi ad Dominum, postquam tradidi librum possessionis Baruch filio Neriae, dicens:
JER|32|17|Heu, Domine Deus, ecce tu fecisti caelum et terram in fortitudine tua magna et in brachio tuo extento; non erit tibi difficile omne verbum,
JER|32|18|qui facis misericordiam in milibus et reddis iniquitatem patrum in sinum filiorum eorum post eos; Deus magne, potens, Dominus exercituum nomen eius:
JER|32|19|magnus consilio et potens in operibus, cuius oculi aperti sunt super omnes vias filiorum Adam, ut reddas unicuique secundum vias suas et secundum fructum operum eius.
JER|32|20|Qui posuisti signa et portenta in terra Aegypti usque ad diem hanc et in Israel et in hominibus; et fecisti tibi nomen, sicut est dies haec.
JER|32|21|Et eduxisti populum tuum Israel de terra Aegypti in signis et in portentis et in manu robusta et in brachio extento et in terrore magno.
JER|32|22|Et dedisti eis terram hanc, quam iurasti patribus eorum, ut dares eis, terram fluentem lacte et melle.
JER|32|23|Et ingressi sunt et possederunt eam; et non oboedierunt voci tuae et in lege tua non ambulaverunt: omnia, quae mandasti eis, ut facerent, non fecerunt; et occurrere fecisti eis omnia mala haec.
JER|32|24|Ecce munitiones exstructae sunt adversum civitatem, ut capiatur, et urbs data est in manu Chaldaeorum, qui proeliantur adversus eam, in gladio et fame et pestilentia; et quaecumque locutus es, acciderunt, ut tu ipse cernis.
JER|32|25|Et tu dicis mihi, Domine Deus: Eme agrum argento et adhibe testes, cum urbs data sit in manu Chaldaeorum ".
JER|32|26|Et factum est verbum Domini ad Ieremiam dicens:
JER|32|27|" Ecce ego Dominus, Deus universae carnis; numquid mihi difficile erit omne verbum?
JER|32|28|Propterea haec dicit Dominus: Ecce ego tradam civitatem istam in manus Chaldaeorum et in manus regis Babylonis, et capiet eam.
JER|32|29|Et venient Chaldaei proeliantes adversum urbem hanc et succendent eam igni et comburent eam et domos, in quarum domatibus sacrificabant Baal et libabant diis alienis libamina ad irritandum me.
JER|32|30|Erant enim filii Israel et filii Iudae iugiter facientes malum in oculis meis ab adulescentia sua, filii Israel, qui usque nunc exacerbant me in opere manuum suarum, dicit Dominus.
JER|32|31|Quia in furorem et in indignationem meam facta est mihi civitas haec a die, qua aedificaverunt eam, usque ad diem istam, qua auferetur de conspectu meo
JER|32|32|propter omnem malitiam filiorum Israel et filiorum Iudae, quam fecerunt, ad iracundiam me provocantes, ipsi et reges eorum, principes eorum et sacerdotes eorum et prophetae eorum, viri Iudae et habitatores Ierusalem.
JER|32|33|Et verterunt ad me terga et non facies, cum docerem eos diluculo consurgens et erudiens, et nollent audire, ut acciperent disciplinam.
JER|32|34|Et posuerunt idola sua in domo, super quam invocatum est nomen meum, ut polluerent eam;
JER|32|35|et aedificaverunt excelsa Baal, quae sunt in valle Benennom, ut initiarent filios suos et filias suas Moloch; quod non mandavi eis, nec ascendit in cor meum, ut facerent abominationem hanc et in peccatum deducerent Iudam ".
JER|32|36|Et nunc propter ista, haec dicit Dominus, Deus Israel, ad civitatem hanc, de qua vos dicitis quod tradatur in manus regis Babylonis in gladio et in fame et in peste:
JER|32|37|" Ecce ego congregabo eos de universis terris, ad quas eieci eos in furore meo et in ira mea et in indignatione grandi; et reducam eos ad locum istum et habitare eos faciam confidenter.
JER|32|38|Et erunt mihi in populum, et ego ero eis in Deum.
JER|32|39|Et dabo eis cor unum et viam unam, ut timeant me universis diebus, et bene sit eis et filiis eorum post eos.
JER|32|40|Et feriam eis pactum sempiternum et non desinam eis benefacere et timorem meum dabo in corde eorum, ut non recedant a me.
JER|32|41|Et laetabor super eis, cum bene eis fecero, et plantabo eos in terra ista in veritate, in toto corde meo et in tota anima mea.
JER|32|42|Quia haec dicit Dominus: Sicut adduxi super populum istum omne malum hoc grande, sic adducam super eos omne bonum, quod ego loquor ad eos,
JER|32|43|et possidebuntur agri in terra ista, de qua vos dicitis quod deserta sit, eo quod non remanserit homo et iumentum, et data sit in manu Chaldaeorum.
JER|32|44|Agri ementur pecunia et scribentur in libro, et imprimetur signum, et testes adhibebuntur in terra Beniamin et in circuitu Ierusalem, in civitatibus Iudae et in civitatibus montanis et in civitatibus Sephelae et in civitatibus, quae ad austrum sunt, quia convertam sortem eorum ", ait Dominus.
JER|33|1|Et factum est verbum Domi ni ad Ieremiam secundo, cum adhuc clausus esset in atrio custodiae, dicens:
JER|33|2|" Haec dicit Dominus, qui facturus est id, Dominus, qui formaturus est illud et paraturus, Dominus nomen eius:
JER|33|3|Clama ad me, et exaudiam te et annuntiabo tibi grandia et inaccessibilia, quae nescis.
JER|33|4|Quia haec dicit Dominus, Deus Israel, super domos urbis huius et ad domos regis Iudae, quae destructae sunt, pro munitionibus et pro gladio
JER|33|5|venientium, ut dimicent cum Chaldaeis et impleant eas cadaveribus hominum, quos percussi in furore meo et in indignatione mea, abscondens faciem meam a civitate hac propter omnem malitiam eorum.
JER|33|6|Ecce ego obducam ei cicatricem et sanitatem et curabo eos et revelabo illis abundantiam pacis et veritatis
JER|33|7|et convertam sortem Iudae et sortem Israel et aedificabo eos sicut a principio.
JER|33|8|Et emundabo illos ab omni iniquitate sua, in qua peccaverunt mihi, et propitius ero cunctis iniquitatibus eorum, in quibus deliquerunt mihi et spreverunt me;
JER|33|9|et erit mihi in nomen et in gaudium et in laudem et in exsultationem cunctis gentibus terrae, quae audierint omnia bona, quae ego facturus sum eis; et pavebunt et turbabuntur in universis bonis et in omni pace, quam ego faciam eis.
JER|33|10|Haec dicit Dominus: Adhuc audietur in loco isto, quem vos dicitis esse desertum, eo quod non sit homo et iumentum in civitatibus Iudae et foris Ierusalem, quae desolatae sunt absque homine et absque habitatore et absque pecore,
JER|33|11|vox gaudii et vox laetitiae, vox sponsi et vox sponsae, vox dicentium:Confitemini Domino exercituum, quoniam bonus Dominus,quoniam in aeternum misericordia eius";et portantium vota in domum Domini; reducam enim sortem terrae sicut a principio, dicit Dominus.
JER|33|12|Haec dicit Dominus exercituum: Adhuc erit in loco isto deserto, absque homine et absque iumento, et in cunctis civitatibus eius habitaculum pastorum accubantium gregum.
JER|33|13|In civitatibus montuosis et in civitatibus Sephelae et in civitatibus, quae ad austrum sunt, et in terra Beniamin et in circuitu Ierusalem et in civitatibus Iudae adhuc transibunt greges ad manum numerantis, ait Dominus.
JER|33|14|Ecce dies veniunt, dicit Dominus, et suscitabo verbum bonum, quod locutus sum ad domum Israel et ad domum Iudae.
JER|33|15|In diebus illis et in tempore illo germinare faciam David germen iustitiae, et faciet iudicium et iustitiam in terra.
JER|33|16|In diebus illis salvabitur Iuda, et Ierusalem habitabit confidenter; et hoc est nomen, quod vocabit eam: Dominus iustitia nostra.
JER|33|17|Quia haec dicit Dominus: Non interibit de David vir, qui sedeat super thronum domus Israel;
JER|33|18|et de sacerdotibus Levitis non interibit vir a facie mea, qui offerat holocautomata et incendat sacrificium et caedat victimas omnibus diebus ".
JER|33|19|Et factum est verbum Domini ad Ieremiam dicens:
JER|33|20|" Haec dicit Dominus: Si irritum potest fieri pactum meum cum die et pactum meum cum nocte, ut non sit dies et nox in tempore suo,
JER|33|21|et pactum meum irritum esse poterit cum David servo meo, ut non sit ex eo filius, qui regnet in throno eius, et cum Levitis sacerdotibus ministris meis.
JER|33|22|Sicuti enumerari non possunt stellae caeli et metiri arena maris, sic multiplicabo semen David servi mei et Levitas ministros meos ".
JER|33|23|Et factum est verbum Domini ad Ieremiam dicens:
JER|33|24|" Numquid non vidisti quid populus hic locutus sit dicens: "Duae cognationes, quas elegerat Dominus, abiectae sunt", et populum meum despexerunt, eo quod non sit ultra gens coram eis?
JER|33|25|Haec dicit Dominus: Si pactum meum inter diem et noctem et leges caelo et terrae non posui,
JER|33|26|equidem et semen Iacob et David servi mei proiciam, ut non assumam de semine eius principes seminis Abraham et Isaac et Iacob; reducam enim sortem eorum et miserebor eis ".
JER|34|1|Verbum, quod factum est ad Ieremiam a Domino, quando Nabuchodonosor rex Babylonis et omnis exercitus eius universaque regna terrae, quae erant sub potestate manus eius, et omnes populi bellabant contra Ierusalem et contra omnes urbes eius, dicens:
JER|34|2|" Haec dicit Dominus, Deus Israel: Vade et loquere ad Sedeciam regem Iudae et dices ad eum: Haec dicit Dominus: Ecce ego tradam civitatem hanc in manus regis Babylonis, et succendet eam igni;
JER|34|3|et tu non effugies de manu eius, sed comprehensione capieris et in manu eius traderis, et oculi tui oculos regis Babylonis videbunt, et os eius cum ore tuo loquetur, et Babylonem introibis.
JER|34|4|Attamen audi verbum Domini, Sedecia rex Iudae. Haec dicit Dominus ad te: Non morieris in gladio,
JER|34|5|sed in pace morieris et secundum combustiones patrum tuorum regum priorum, qui fuerunt ante te, sic comburent tibi et "Vae, domine!" plangent te, quia verbum ego locutus sum ", dicit Dominus.
JER|34|6|Et locutus est Ieremias propheta ad Sedeciam regem Iudae universa verba haec in Ierusalem;
JER|34|7|et exercitus regis Babylonis pugnabat contra Ierusalem et contra omnes civitates Iudae, quae reliquae erant, contra Lachis et contra Azeca: hae enim supererant de civitatibus Iudae urbes munitae.
JER|34|8|Verbum, quod factum est ad Ieremiam a Domino, postquam percussit rex Sedecias foedus cum omni populo in Ierusalem praedicans eis libertatem,
JER|34|9|ut dimitteret unusquisque servum suum et unusquisque ancillam suam, Hebraeum et Hebraeam, liberos et nequaquam dominarentur eis, id est in Iudaeo et fratre suo.
JER|34|10|Audierunt ergo omnes principes et universus populus, qui inierant pactum, ut dimitteret unusquisque servum suum et unusquisque ancillam suam liberos et ultra non dominarentur eis; audierunt igitur et dimiserunt.
JER|34|11|Et conversi sunt deinceps et retraxerunt servos et ancillas suas, quos dimiserant liberos, et subiugaverunt in famulos et in famulas.
JER|34|12|Et factum est verbum Domini ad Ieremiam a Domino dicens:
JER|34|13|" Haec dicit Dominus, Deus Israel: Ego percussi foedus cum patribus vestris in die, qua eduxi eos de terra Aegypti de domo servitutis, dicens:
JER|34|14|Cum completi fuerint septem anni, dimittat unusquisque fratrem suum Hebraeum, qui venditus est ei, et serviet tibi sex annis, et dimittes eum a te liberum, et non audierunt patres vestri me nec inclinaverunt aurem suam.
JER|34|15|Et conversi estis vos hodie et fecistis, quod rectum est in oculis meis, ut praedicaretis libertatem unusquisque ad proximum suum; et inistis pactum in conspectu meo in domo, super quam invocatum est nomen meum.
JER|34|16|Et reversi estis et commaculastis nomen meum et reduxistis unusquisque servum suum et unusquisque ancillam suam, quos dimiseratis, ut essent liberi et suae potestatis, et subiugastis eos, ut sint vobis servi et ancillae.
JER|34|17|Propterea haec dicit Dominus: Vos non audistis me, ut praedicaretis libertatem unusquisque fratri suo et unusquisque amico suo; ecce ego praedico vobis libertatem, ait Dominus, ad gladium et pestem et famem et dabo vos in commotionem cunctis regnis terrae.
JER|34|18|Et dabo viros, qui praevaricantur foedus meum et non observaverunt verba foederis, quibus assensi sunt in conspectu meo, sicut vitulum, quem conciderunt in duas partes et transierunt inter divisiones eius,
JER|34|19|principes Iudae et principes Ierusalem, eunuchi et sacerdotes et omnis populus terrae, qui transierunt inter divisiones vituli;
JER|34|20|et dabo eos in manu inimicorum suorum et in manu quaerentium animam eorum, et erit morticinum eorum in escam volatilibus caeli et bestiis terrae.
JER|34|21|Et Sedeciam regem Iudae et principes eius dabo in manus inimicorum suorum et in manus quaerentium animas eorum et in manus exercituum regis Babylonis, qui recesserunt a vobis.
JER|34|22|Ecce ego praecipio, dicit Dominus, et reducam eos in civitatem hanc; et proeliabuntur adversus eam et capient eam et incendent igni; et civitates Iudae dabo in solitudinem, eo quod non sit habitator ".
JER|35|1|Verbum, quod factum est ad Ieremiam a Domino in die bus Ioachim filii Iosiae regis Iudae dicens:
JER|35|2|" Vade ad domum Rechabitarum et loquere eis; et introduces eos in domum Domini in unam exedram et dabis eis bibere vinum ".
JER|35|3|Et assumpsi Iezoniam filium Ieremiae filii Habsaniae et fratres eius et omnes filios eius et universam domum Rechabitarum;
JER|35|4|et introduxi eos in domum Domini ad exedram filiorum Hanan filii Iegdaliae hominis Dei, quod erat iuxta exedram principum super exedram Maasiae filii Sellum, qui erat custos vestibuli.
JER|35|5|Et posui coram filiis domus Rechabitarum scyphos plenos vino et calices et dixi ad eos: " Bibite vinum ".
JER|35|6|Qui responderunt: " Non bibemus vinum, quia Ionadab filius Rechab pater noster praecepit nobis dicens: "Non bibetis vinum, vos et filii vestri, usque in sempiternum
JER|35|7|et domum non aedificabitis et sementem non seretis et vineas non plantabitis, nec habebitis, sed in tabernaculis habitabitis cunctis diebus vestris, ut vivatis diebus multis super faciem terrae, in qua vos peregrinamini".
JER|35|8|Oboedivimus ergo voci Ionadab filii Rechab patris nostri in omnibus, quae praecepit nobis, ita ut non biberemus vinum cunctis diebus nostris, nos et mulieres nostrae, filii et filiae nostrae,
JER|35|9|et non aedificaremus domos ad habitandum et vineam et agrum et sementem non habuimus,
JER|35|10|sed habitavimus in tabernaculis; et oboedientes fecimus iuxta omnia, quae praecepit nobis Ionadab pater noster.
JER|35|11|Cum autem ascendisset Nabuchodonosor rex Babylonis ad terram, diximus: Venite, et ingrediamur Ierusalem a facie exercitus Chaldaeorum et a facie exercitus Syriae. Et mansimus in Ierusalem ".
JER|35|12|Et factum est verbum Domini ad Ieremiam dicens:
JER|35|13|" Haec dicit Dominus exercituum, Deus Israel: Vade et dic viris Iudae et habitatoribus Ierusalem: Numquid non recipietis disciplinam, ut oboediatis verbis meis?, dicit Dominus.
JER|35|14|Praevaluerunt sermones Ionadab filii Rechab, quos praecepit filiis suis, ut non biberent vinum, et non biberunt usque ad diem hanc, quia oboedierunt praecepto patris sui; ego autem locutus sum ad vos de mane consurgens et loquens, et non oboedistis mihi.
JER|35|15|Misique ad vos omnes servos meos prophetas, consurgens diluculo mittensque et dicens: Convertimini unusquisque a via sua pessima et bona facite opera vestra et nolite sequi deos alienos neque colatis eos, et habitabitis in terra, quam dedi vobis et patribus vestris, et non inclinastis aurem vestram neque audistis me.
JER|35|16|Firmaverunt igitur filii Ionadab filii Rechab praeceptum patris sui, quod praeceperat eis; populus autem iste non oboedivit mihi.
JER|35|17|Idcirco haec dicit Dominus exercituum, Deus Israel: Ecce ego adducam super Iudam et super omnes habitatores Ierusalem universam afflictionem, quam locutus sum adversum illos, eo quod locutus sum ad illos, et non audierunt, vocavi illos, et non responderunt mihi ".
JER|35|18|Domui autem Rechabitarum dixit Ieremias: " Haec dicit Dominus exercituum, Deus Israel: Pro eo quod oboedistis praecepto Ionadab patris vestri et custodistis omnia mandata eius et fecistis universa, quae praecepit vobis,
JER|35|19|propterea haec dicit Dominus exercituum, Deus Israel: Non deficiet vir de stirpe Ionadab filii Rechab stans in conspectu meo cunctis diebus ".
JER|36|1|Et factum est in anno quarto Ioachim filii Iosiae regis Iudae, factum est verbum hoc ad Ieremiam a Domino dicens:
JER|36|2|" Tolle volumen libri et scribes in eo omnia verba, quae locutus sum tibi adversum Israel et Iudam et adversum omnes gentes a die qua locutus sum ad te ex diebus Iosiae usque ad diem hanc,
JER|36|3|si forte, audiente domo Iudae universa mala, quae ego cogito facere eis, revertatur unusquisque a via sua pessima, et propitius ero iniquitati et peccato eorum ".
JER|36|4|Vocavit ergo Ieremias Baruch filium Neriae; et scripsit Baruch ex ore Ieremiae omnes sermones Domini, quos locutus est ad eum, in volumine libri.
JER|36|5|Et praecepit Ieremias Baruch dicens: " Ego impeditus sum nec valeo ingredi domum Domini.
JER|36|6|Ingredere ergo tu et lege de volumine, in quo scripsisti ex ore meo verba Domini, audiente populo in domo Domini, in die ieiunii; insuper et audiente universo Iuda, qui veniunt de civitatibus suis, leges eis,
JER|36|7|si forte cadat oratio eorum in conspectu Domini, et revertatur unusquisque a via sua pessima, quoniam magnus furor et indignatio est, quam locutus est Dominus adversus populum hunc ".
JER|36|8|Et fecit Baruch filius Neriae iuxta omnia, quae praeceperat ei Ieremias propheta, legens ex volumine sermones Domini in domo Domini.
JER|36|9|Factum est autem in anno quinto Ioachim filii Iosiae regis Iudae, in mense nono, praedicaverunt ieiunium in conspectu Domini omni populo in Ierusalem et universae multitudini, quae confluxerat de civitatibus Iudae in Ierusalem.
JER|36|10|Legitque Baruch ex volumine sermones Ieremiae in domo Domini, in exedra Gamariae filii Saphan scribae in vestibulo superiore, in introitu portae Novae domus Domini, audiente omni populo.
JER|36|11|Cumque audisset Michaeas filius Gamariae filii Saphan omnes sermones Domini ex libro,
JER|36|12|descendit in domum regis ad exedram scribae; et ecce ibi omnes principes sedebant: Elisama scriba et Dalaias filius Semiae et Elnathan filius Achobor et Gamarias filius Saphan et Sedecias filius Hananiae et universi principes.
JER|36|13|Et nuntiavit eis Michaeas omnia verba, quae audivit, legente Baruch ex volumine in auribus populi.
JER|36|14|Miserunt itaque omnes principes ad Baruch Iudi filium Nathaniae filii Selemiae filii Chusi dicentes: " Volumen, ex quo legisti audiente populo, sume in manu tua et veni ". Tulit ergo Baruch filius Neriae volumen in manu sua et venit ad eos.
JER|36|15|Et dixerunt ad eum: " Sede et lege haec in auribus nostris "; et legit Baruch in auribus eorum.
JER|36|16|Igitur cum audissent omnia verba, obstupuerunt unusquisque ad proximum suum; et dixerunt ad Baruch: "Nuntiare debemus regi omnes sermones istos".
JER|36|17|Et interrogaverunt Baruch dicentes: " Indica nobis, quomodo scripsisti omnes sermones istos ex ore eius ".
JER|36|18|Dixit autem eis Baruch: " Ex ore suo loquebatur ad me omnes sermones istos, et ego scribebam in volumine atramento ".
JER|36|19|Et dixerunt principes ad Baruch: " Vade et abscondere, tu et Ieremias, et nemo sciat, ubi sitis ".
JER|36|20|Et ingressi sunt ad regem in atrium, porro volumen deposuerunt in exedra Elisamae scribae; et nuntiaverunt audiente rege omnes sermones.
JER|36|21|Misitque rex Iudi, ut sumeret volumen; qui, tollens illud de exedra Elisamae scribae, legit audiente rege et universis principibus, qui stabant circa regem.
JER|36|22|Rex autem sedebat in domo hiemali in mense nono, et posita erat arula coram eo plena prunis;
JER|36|23|cumque legisset Iudi tres pagellas vel quattuor, scidit eas scalpello scribae et proiecit in ignem, qui erat super arulam, donec consumeretur omne volumen igni, qui erat in arula.
JER|36|24|Et non timuerunt neque sciderunt vestimenta sua rex et omnes servi eius, qui audierunt universos sermones istos.
JER|36|25|Verumtamen Elnathan et Dalaias et Gamarias instanter rogaverunt regem, ne combureret librum, et non audivit eos.
JER|36|26|Et praecepit rex Ierameel filio regis et Saraiae filio Azriel et Selemiae filio Abdeel, ut comprehenderent Baruch scribam et Ieremiam prophetam; abscondit autem eos Dominus.
JER|36|27|Et factum est verbum Domini ad Ieremiam, postquam combusserat rex volumen et sermones, quos scripserat Baruch ex ore Ieremiae, dicens:
JER|36|28|"Rursum tolle volumen aliud et scribe in eo omnes sermones priores, qui erant in primo volumine, quod combussit Ioachim rex Iudae.
JER|36|29|Et super Ioachim regem Iudae dices: Haec dicit Dominus: Tu combussisti volumen illud dicens: "Quare scripsisti in eo annuntians: Certe veniet rex Babylonis et vastabit terram hanc et cessare faciet ex illa hominem et iumentum?".
JER|36|30|Propterea haec dicit Dominus contra Ioachim regem Iudae: Non erit ex eo, qui sedeat super solium David, et cadaver eius proicietur ad aestum per diem et ad gelu per noctem;
JER|36|31|et visitabo contra eum et contra semen eius et contra servos eius iniquitates suas; et adducam super eos et super habitatores Ierusalem et super viros Iudae omne malum, quod locutus sum ad eos, et non audierunt ".
JER|36|32|Ieremias autem tulit volumen aliud et dedit illud Baruch filio Neriae scribae; qui scripsit in eo ex ore Ieremiae omnes sermones libri, quem combusserat Ioachim rex Iudae igni; et insuper additi sunt multi sermones similes illis.
JER|37|1|Et regnavit rex Sedecias filius Iosiae pro Iechonia filio Ioachim; quem constituit regem Nabuchodonosor rex Babylonis in terra Iudae.
JER|37|2|Et non oboedivit, ipse et servi eius et populus terrae, verbis Domini, quae locutus est in manu Ieremiae prophetae.
JER|37|3|Et misit rex Sedecias Iuchal filium Selemiae et Sophoniam filium Maasiae sacerdotem ad Ieremiam prophetam dicens: " Ora pro nobis Dominum Deum nostrum ".
JER|37|4|Ieremias autem libere ambulabat in medio populi; non enim miserant eum in custodiam carceris.
JER|37|5|Igitur exercitus pharaonis egressus est de Aegypto, et audientes Chaldaei, qui obsidebant Ierusalem, huiuscemodi nuntium recesserunt ab Ierusalem.
JER|37|6|Et factum est verbum Domini ad Ieremiam prophetam dicens:
JER|37|7|" Haec dicit Dominus, Deus Israel: Sic dicetis regi Iudae, qui misit vos ad me interrogandum: Ecce exercitus pharaonis, qui egressus est vobis in auxilium, revertetur in terram suam in Aegyptum;
JER|37|8|et redient Chaldaei et bellabunt contra civitatem hanc et capient eam et succendent eam igni.
JER|37|9|Haec dicit Dominus: Nolite decipere animas vestras dicentes: "Euntes abibunt et recedent a nobis Chaldaei", quia non abibunt.
JER|37|10|Sed et si percusseritis omnem exercitum Chaldaeorum, qui proeliantur adversum vos, et derelicti fuerint ex eis aliqui vulnerati, singuli de tentorio suo consurgent et incendent civitatem hanc igni ".
JER|37|11|Ergo cum recessisset exercitus Chaldaeorum ab Ierusalem propter exercitum pharaonis,
JER|37|12|egressus est Ieremias de Ierusalem, ut iret in terram Beniamin et divideret ibi possessionem in conspectu populi.
JER|37|13|Cumque pervenisset ad portam Beniamin, erat ibi custos portae nomine Ierias filius Selemiae filii Hananiae; et apprehendit Ieremiam prophetam dicens: " Ad Chaldaeos profugis ".
JER|37|14|Et respondit Ieremias: " Falsum est! Non fugio ad Chaldaeos ". Et non audivit eum; sed comprehendit Ierias Ieremiam et adduxit eum ad principes.
JER|37|15|Et irati sunt principes contra Ieremiam, quem caesum miserunt in carcerem, qui erat in domo Ionathan scribae; eam enim in carcerem fecerant.
JER|37|16|Itaque ingressus est Ieremias in domum laci fornice tectam; et sedit ibi Ieremias diebus multis.
JER|37|17|Mittens autem Sedecias rex tulit eum et interrogavit eum in domo sua abscondite et dixit: " Putasne est sermo a Domino? ". Et dixit Ieremias: " Est "; et ait: "In manus regis Babylonis traderis ".
JER|37|18|Et dixit Ieremias ad regem Sedeciam: " Quid peccavi tibi et servis tuis et populo isti, quia misistis me in domum carceris?
JER|37|19|Ubi sunt prophetae vestri, qui prophetabant vobis et dicebant: "Non veniet rex Babylonis super vos et super terram hanc"?
JER|37|20|Nunc ergo audi, obsecro, domine mi rex; valeat deprecatio mea in conspectu tuo, et ne me remittas in domum Ionathan scribae, ne moriar ibi.
JER|37|21|Praecepit ergo rex Sedecias, ut traderetur Ieremias in vestibulo custodiae, et daretur ei torta panis cotidie ex vico Pistorum, donec consumerentur omnes panes de civitate. Et mansit Ieremias in vestibulo custodiae.
JER|38|1|Audivit autem Saphatias fi lius Matthan et Godolias fi lius Phassur et Iuchal filius Selemiae et Phassur filius Melchiae sermones, quos Ieremias loquebatur ad omnem populum dicens:
JER|38|2|" Haec dicit Dominus: Quicumque manserit in civitate hac, morietur gladio et fame et peste; qui autem profugerit ad Chaldaeos, vivet, et erit anima eius quasi spolium et vivet.
JER|38|3|Haec dicit Dominus: Certe tradetur civitas haec in manu exercitus regis Babylonis, et capiet eam ".
JER|38|4|Et dixerunt principes regi: " Rogamus, ut occidatur homo iste; de industria enim dissolvit manus virorum bellantium, qui remanserunt in civitate hac, et manus universi populi loquens ad eos iuxta verba haec; siquidem homo iste non quaerit pacem populo huic sed malum ".
JER|38|5|Et dixit rex Sedecias: " Ecce ipse in manibus vestris est; nequit enim rex vobis quidquam negare ".
JER|38|6|Tulerunt ergo Ieremiam et proiecerunt eum in lacum Melchiae filii regis, qui erat in vestibulo custodiae. Et submiserunt Ieremiam funibus. Et in lacu non erat aqua sed lutum; descendit itaque Ieremias in caenum.
JER|38|7|Audivit autem Abdemelech Aethiops, vir eunuchus, qui erat in domo regis, quod misissent Ieremiam in lacum; porro rex sedebat in porta Beniamin.
JER|38|8|Et egressus est Abdemelech de domo regis et locutus est ad regem dicens:
JER|38|9|" Domine mi rex, malefecerunt viri isti omnia, quaecumque perpetrarunt contra Ieremiam prophetam, mittentes eum in lacum, ut moriatur ibi fame; non sunt enim panes ultra in civitate ".
JER|38|10|Praecepit itaque rex Abdemelech Aethiopi dicens: " Tolle tecum hinc triginta viros et leva Ieremiam prophetam de lacu, antequam moriatur ".
JER|38|11|Assumptis ergo Abdemelech secum viris, ingressus est domum regis, in conclave, quod erat sub thesauro, et tulit inde pannos ex vestibus veteribus et scissis et submisit eos ad Ieremiam in lacum per funiculos.
JER|38|12|Dixitque Abdemelech Aethiops ad Ieremiam: " Pone veteres pannos et haec scissa sub scapuli et postea funes ". Fecit ergo Ieremias sic;
JER|38|13|et extraxerunt Ieremiam funibus et eduxerunt eum de lacu. Mansit autem Ieremias in vestibulo custodiae.
JER|38|14|Et misit rex Sedecias et tulit ad se Ieremiam prophetam ad ostium tertium, quod erat in domo Domini; et dixit rex ad Ieremiam: "Interrogo ego te sermonem, ne abscondas a me aliquid ".
JER|38|15|Dixit autem Ieremias ad Sedeciam: " Si annuntiavero tibi, numquid non interficies me? Et si consilium dedero tibi, non me audies ".
JER|38|16|Iuravit ergo rex Sedecias Ieremiae clam dicens: " Vivit Dominus, qui fecit nobis animam hanc, non occidam te et non tradam te in manu virorum istorum, qui quaerunt animam tuam ".
JER|38|17|Et dixit Ieremias ad Sedeciam: " Haec dicit Dominus exercituum, Deus Israel: Si profectus exieris ad principes regis Babylonis, vivet anima tua, et civitas haec non succendetur igni, et salvus eris tu et domus tua;
JER|38|18|si autem non exieris ad principes regis Babylonis, tradetur civitas haec in manu Chaldaeorum, et succendent eam igni, et tu non effugies de manu eorum ".
JER|38|19|Et dixit rex Sedecias ad Ieremiam: " Sollicitus sum propter Iudaeos, qui transfugerunt ad Chaldaeos, ne forte tradar in manus eorum, et illudant mihi ".
JER|38|20|Respondit autem Ieremias: " Non te tradent; audi, quaeso, vocem Domini, quam ego loquor ad te, et bene tibi erit, et vivet anima tua.
JER|38|21|Quod si nolueris egredi, iste est sermo, quem ostendit mihi Dominus:
JER|38|22|Ecce omnes mulieres, quae remanserunt in domo regis Iudae, educentur ad principes regis Babylonis et ipsae dicent:Seduxerunt te et praevaluerunt adversum teviri pacifici tui;demersi sunt in caeno pedes tui,illi autem recesserunt a te".
JER|38|23|Et omnes uxores tuae et filii tui educentur ad Chaldaeos, et non effugies manus eorum, sed in manu regis Babylonis capieris; et civitatem hanc comburet igni ".
JER|38|24|Dixit ergo Sedecias ad Ieremiam: " Nullus sciat verba haec, et non morieris.
JER|38|25|Si autem audierint principes quia locutus sum tecum, et venerint ad te et dixerint tibi: "Indica nobis, quid locutus sis cum rege, ne celes nos, et non te interficiemus, et quid locutus est tecum rex",
JER|38|26|dices ad eos: "Prostravi ego preces meas coram rege, ne me reduci iuberet in domum Ionathan, et ibi morerer" ".
JER|38|27|Venerunt ergo omnes principes ad Ieremiam et interrogaverunt eum, et locutus est eis iuxta omnia verba, quae praeceperat ei rex; et cessaverunt ab eo: nihil enim fuerat auditum.
JER|38|28|Mansit vero Ieremias in vestibulo custodiae usque ad diem, quo capta est Ierusalem.Et factum est ut caperetur Ierusalem.
JER|39|1|Anno nono Sedeciae regis Iudae, mense decimo, venit Nabuchodonosor rex Babylonis et omnis exercitus eius ad Ierusalem et obsidebant eam.
JER|39|2|Undecimo autem anno Sedeciae, mense quarto, nona mensis, aperta est civitas;
JER|39|3|et ingressi sunt omnes principes regis Babylonis et sederunt in porta Media: Nergelsereser Samegarnabu, Sarsachim princeps eunuchorum, Nergelsereser princeps magorum et omnes reliqui principes regis Babylonis.
JER|39|4|Cumque vidisset eos Sedecias rex Iudae et omnes viri bellatores, fugerunt et egressi sunt nocte de civitate per viam horti regis et per portam, quae erat inter duos muros, et egressi sunt ad viam Arabae.
JER|39|5|Persecutus est autem eos exercitus Chaldaeorum; et comprehenderunt Sedeciam in campestribus Iericho et captum adduxerunt ad Nabuchodonosor regem Babylonis in Rebla, quae est in terra Emath; et locutus est ad eum iudicia.
JER|39|6|Et occidit rex Babylonis filios Sedeciae in Rebla in oculis eius, et omnes nobiles Iudae occidit rex Babylonis;
JER|39|7|oculos quoque Sedeciae eruit et vinxit eum compedibus, ut duceretur in Babylonem.
JER|39|8|Domum quoque regis et domum vulgi succenderunt Chaldaei igni; et murum Ierusalem subverterunt.
JER|39|9|Et reliquias populi, quae remanserant in civitate, et perfugas, qui transfugerant ad eum, et superfluos artificum, qui remanserant, transtulit Nabuzardan magister satellitum in Babylonem.
JER|39|10|Et de plebe pauperum, qui nihil penitus habebant, dimisit Nabuzardan magister satellitum in terra Iudae; et dedit eis vineas et agros in die illa.
JER|39|11|Praeceperat autem Nabuchodonosor rex Babylonis de Ieremia Nabuzardan magistro satellitum dicens:
JER|39|12|" Tolle illum et pone super eum oculos tuos nihilque ei mali facias, sed, ut voluerit, sic facies ei ".
JER|39|13|Misit ergo Nabuzardan princeps satellitum et Nabusezban princeps eunuchorum et Nergelsereser princeps magorum et omnes optimates regis Babylonis
JER|39|14|miserunt et tulerunt Ieremiam de vestibulo custodiae et tradiderunt eum Godoliae filio Ahicam filii Saphan, ut duceret domum. Et habitavit in populo.
JER|39|15|Ad Ieremiam autem factus fuerat sermo Domini, cum clausus esset in vestibulo custodiae, dicens:
JER|39|16|" Vade et dic Abdemelech Aethiopi dicens: Haec dicit Dominus exercituum, Deus Israel: Ecce ego inducam sermones meos super civitatem hanc in malum et non in bonum; et erunt in conspectu tuo in die illa.
JER|39|17|Et liberabo te in die illa, ait Dominus, et non traderis in manus virorum, quos tu formidas;
JER|39|18|sed eruens liberabo te, et gladio non cades, sed erit tibi anima tua quasi spolium, quia in me habuisti fiduciam ", ait Dominus.
JER|40|1|Sermo, qui factus est ad Ieremiam a Domino, postquam dimissus est a Nabuzardan magistro satellitum de Rama, quando tulit eum vinctum catenis in medio omnium, qui migrabant de Ierusalem et Iuda et ducebantur in Babylonem.
JER|40|2|Tollens ergo princeps satellitum Ieremiam, dixit ad eum: " Dominus Deus tuus locutus est malum hoc super locum istum
JER|40|3|et adduxit; et fecit Dominus, sicut locutus est, quia peccastis Domino et non audistis vocem eius, et factus est vobis sermo hic.
JER|40|4|Nunc ergo ecce solvi te hodie de catenis, quae sunt in manibus tuis. Si placet tibi, ut venias mecum in Babylonem, veni, et ponam oculos meos super te; si autem displicet tibi venire mecum in Babylonem, reside; ecce omnis terra in conspectu tuo est: quod elegeris et quo placuerit tibi ut vadas, illuc perge ".
JER|40|5|Cum nondum reverteretur, dixit: " Revertere ad Godoliam filium Ahicam filii Saphan, quem praeposuit rex Babylonis civitatibus Iudae; habita ergo cum eo in medio populi vel quocumque placuerit tibi ut vadas, vade ". Dedit quoque ei magister satellitum cibaria et munuscula et dimisit eum.
JER|40|6|Venit autem Ieremias ad Godoliam filium Ahicam in Maspha et habitavit cum eo in medio populi, qui relictus fuerat in terra.
JER|40|7|Cumque audissent omnes principes exercitus, qui dispersi fuerant per regiones, ipsi et viri eorum, quod praefecisset rex Babylonis Godoliam filium Ahicam terrae et quod commendasset ei viros et mulieres et parvulos et de pauperibus terrae, qui non fuerant translati in Babylonem,
JER|40|8|venerunt ad Godoliam in Maspha; Ismael, inquam, filius Nathaniae et Iohanan et Ionathan filii Caree et Saraia filius Thanehumeth et filii Ophi, qui erant de Netopha, et Iezonias filius Maachathi, ipsi et viri eorum.
JER|40|9|Et iuravit eis Godolias filius Ahicam filii Saphan et comitibus eorum dicens: "Nolite timere servire Chaldaeis; habitate in terra et servite regi Babylonis, et bene erit vobis.
JER|40|10|Ecce ego habito in Maspha, ut stem coram Chaldaeis, qui veniunt ad nos; vos autem colligite vindemiam et messem et oleum et condite in vasis vestris et manete in urbibus vestris, quas tenetis ".
JER|40|11|Sed et omnes Iudaei, qui erant in Moab et in filiis Ammon et in Edom et in universis regionibus, audito quod dedisset rex Babylonis reliquias in Iudaea et quod praeposuisset super eos Godoliam filium Ahicam filii Saphan,
JER|40|12|reversi sunt, inquam, omnes Iudaei de universis locis, ad quae profugerant, et venerunt in terram Iudae ad Godoliam in Maspha et collegerunt vinum et messem multam nimis.
JER|40|13|Iohanan autem filius Caree et omnes principes exercitus, qui dispersi fuerant in regionibus, venerunt ad Godoliam in Maspha
JER|40|14|et dixerunt ei: " Scito quod Baalis rex filiorum Ammon misit Ismael filium Nathaniae percutere animam tuam "; et non credidit eis Godolias filius Ahicam.
JER|40|15|Iohanan vero filius Caree dixit ad Godoliam seorsum in Maspha loquens: Ibo et percutiam Ismael filium Nathaniae, nullo sciente, ne interficiat animam tuam, et dissipentur omnes Iudaei, qui congregati sunt ad te, et peribunt reliquiae Iudae ".
JER|40|16|Et ait Godolias filius Ahicam ad Iohanan filium Caree: " Noli facere verbum hoc; falsum enim tu loqueris de Ismael ".
JER|41|1|Et factum est in mense septi mo, venit Ismael filius Nathaniae filii Elisama de semine regali et optimates regis et decem viri cum eo ad Godoliam filium Ahicam in Maspha; et comederunt ibi panes simul in Maspha.
JER|41|2|Surrexit autem Ismael filius Nathaniae et decem viri, qui cum eo erant, et percusserunt Godoliam filium Ahicam filii Saphan gladio; et interfecerunt eum, quem praefecerat rex Babylonis terrae.
JER|41|3|Omnes quoque Iudaeos, qui erant cum Godolia in Maspha, et Chaldaeos, qui reperti sunt ibi, et viros bellatores percussit Ismael.
JER|41|4|Secundo autem die postquam occiderat Godoliam, nullo adhuc sciente,
JER|41|5|venerunt viri de Sichem et de Silo et de Samaria, octoginta viri, rasi barba et scissis vestibus et incisi in cute, et munera et tus habebant in manu, ut offerrent in domo Domini.
JER|41|6|Egressus ergo Ismael filius Nathaniae in occursum eorum de Maspha, incedens et plorans ibat. Cum autem occurrisset eis, dixit ad eos: " Venite ad Godoliam filium Ahicam ".
JER|41|7|Qui cum venissent ad medium civitatis, interfecit eos Ismael filius Nathaniae et proiecit in medium laci, ipse et viri, qui erant cum eo.
JER|41|8|Decem autem viri reperti sunt inter eos, qui dixerunt ad Ismael: " Noli occidere nos, quia habemus thesauros in agro, frumenti et hordei et olei et mellis "; et cessavit et non interfecit eos cum fratribus suis.
JER|41|9|Lacus autem, in quem proiecerat Ismael omnia cadavera virorum, quos percussit, est lacus magnus, quem fecit rex Asa propter Baasa regem Israel; ipsum replevit Ismael filius Nathaniae occisis.
JER|41|10|Et captivas duxit Ismael omnes reliquias populi, qui erant in Maspha, filias regis et universum populum, qui remanserat in Maspha, quos commendaverat Nabuzardan princeps satellitum Godoliae filio Ahicam; et cepit eos Ismael filius Nathaniae et abiit, ut transiret ad filios Ammon.
JER|41|11|Audivit autem Iohanan filius Caree et omnes principes bellatorum, qui erant cum eo, omne malum, quod fecerat Ismael filius Nathaniae,
JER|41|12|et, assumptis universis viris, profecti sunt, ut bellarent adversum Ismael filium Nathaniae; et invenerunt eum ad aquas multas, quae sunt in Gabaon.
JER|41|13|Cumque vidisset omnis populus, qui erat cum Ismael, Iohanan filium Caree et universos principes bellatorum, qui erant cum eo, laetati sunt.
JER|41|14|Et omnis populus, quem ceperat Ismael in Maspha, reversus est et abiit ad Iohanan filium Caree;
JER|41|15|Ismael autem filius Nathaniae fugit cum octo viris a facie Iohanan et abiit ad filios Ammon.
JER|41|16|Tulit ergo Iohanan filius Caree et omnes principes bellatorum, qui erant cum eo, universas reliquias vulgi, quas reduxerat ab Ismael filio Nathaniae venientes de Maspha, postquam percussit Godoliam filium Ahicam, viros fortes ad proelium et mulieres et pueros et eunuchos, quos reduxerat de Gabaon.
JER|41|17|Et abierunt et sederunt in Gherutchamaam, quae est iuxta Bethlehem, ut pergerent et introirent Aegyptum
JER|41|18|a facie Chaldaeorum; timebant enim eos, quia percusserat Ismael filius Nathaniae Godoliam filium Ahicam, quem praeposuerat rex Babylonis in regione.
JER|42|1|Et accesserunt omnes princi pes bellatorum, scilicet Iohanan filius Caree et Iezonias filius Osaiae et universum vulgus, a parvo usque ad magnum,
JER|42|2|dixeruntque ad Ieremiam prophetam: " Cadat oratio nostra in conspectu tuo, et ora pro nobis ad Dominum Deum tuum pro universis reliquiis istis, quia derelicti sumus pauci de pluribus, sicut oculi tui nos intuentur;
JER|42|3|et annuntiet nobis Dominus Deus tuus viam, per quam pergamus, et verbum, quod faciamus ".
JER|42|4|Dixit autem ad eos Ieremias propheta: " Audivi. Ecce ego oro ad Dominum Deum vestrum secundum verba vestra; omne verbum, quodcumque responderit pro vobis, indicabo vobis nec celabo vos quidquam ".
JER|42|5|Et illi dixerunt ad Ieremiam: " Sit Dominus inter nos testis verax et fidelis, si non iuxta omne verbum, in quo miserit te Dominus Deus tuus ad nos, sic faciemus.
JER|42|6|Sive bonum est sive malum, voci Domini Dei nostri, ad quem mittimus te, oboediemus, ut bene sit nobis, cum audierimus vocem Domini Dei nostri ".
JER|42|7|Cum autem completi essent decem dies, factum est verbum Domini ad Ieremiam;
JER|42|8|vocavitque Iohanan filium Caree et omnes principes bellatorum, qui erant cum eo, et universum populum a minimo usque ad magnum
JER|42|9|et dixit ad eos: " Haec dicit Dominus, Deus Israel, ad quem misistis me, ut prosternerem preces vestras in conspectu eius:
JER|42|10|Si quiescentes manseritis in terra hac, aedificabo vos et non destruam, plantabo et non evellam; iam enim placatus sum super malo, quod feci vobis.
JER|42|11|Nolite timere a facie regis Babylonis, quem vos pavidi formidatis; nolite metuere eum, dicit Dominus, quia vobiscum sum ego, ut salvos vos faciam et eruam de manu eius;
JER|42|12|et dabo vobis, ut misericordiam inveniatis, et ipse miserebitur vestri et habitare vos faciet in terra vestra.
JER|42|13|Si autem dixeritis vos: "Non habitabimus in terra ista", nec audieritis vocem Domini Dei vestri
JER|42|14|dicentes: "Nequaquam, sed ad terram Aegypti pergemus, ubi non videbimus bellum et clangorem tubae non audiemus et famem non sustinebimus et ibi habitabimus",
JER|42|15|propter hoc nunc audite verbum Domini, reliquiae Iudae: Haec dicit Dominus exercituum, Deus Israel: Si posueritis faciem vestram, ut ingrediamini Aegyptum, et intraveritis, ut ibi peregrinemini,
JER|42|16|gladius, quem vos formidatis, ibi comprehendet vos in terra Aegypti, et fames, pro qua estis solliciti, adhaerebit vobis in Aegypto, et ibi moriemini.
JER|42|17|Omnesque viri, qui posuerunt faciem suam, ut ingrediantur Aegyptum et peregrinentur ibi, morientur gladio et fame et peste: nullus de eis remanebit nec effugiet a facie mali, quod ego afferam super eos.
JER|42|18|Quia haec dicit Dominus exercituum, Deus Israel: Sicut effusus est furor meus et indignatio mea super habitatores Ierusalem, sic effundetur indignatio mea super vos, cum ingressi fueritis Aegyptum, et eritis in exsecrationem et in stuporem et in maledictum et in opprobrium et nequaquam ultra videbitis locum istum ".
JER|42|19|Verbum Domini super vos, reliquiae Iudae: " Nolite intrare Aegyptum; scientes scietis quia obtestatus sum vos hodie,
JER|42|20|quia decepistis animas vestras. Vos enim misistis me ad Dominum Deum nostrum dicentes: "Ora pro nobis ad Dominum Deum nostrum et iuxta omnia, quaecumque dixerit tibi Dominus Deus noster, sic annuntia nobis, et faciemus".
JER|42|21|Et annuntiavi vobis hodie, et non audistis vocem Domini Dei vestri super universis, pro quibus misit me ad vos.
JER|42|22|Nunc ergo scientes scietis quia gladio et fame et peste moriemini in loco, ad quem voluistis intrare et ibi peregrinari ".
JER|43|1|Factum est autem, cum complesset Ieremias loquens ad populum universos sermones Domini Dei eorum, pro quibus miserat eum Dominus Deus eorum ad illos omnia verba haec,
JER|43|2|dixit Azarias filius Osaiae et Iohanan filius Caree et omnes viri superbi dicentes ad Ieremiam: " Mendacium tu loqueris; non misit te Dominus Deus noster dicens: "Ne ingrediamini Aegyptum, ut illic peregrinemini",
JER|43|3|sed Baruch filius Neriae incitat te adversum nos, ut tradat nos in manu Chaldaeorum, ut interficiant nos et traducant in Babylonem ".
JER|43|4|Et non audivit Iohanan filius Caree et omnes principes bellatorum et universus populus vocem Domini, ut manerent in terra Iudae.
JER|43|5|Sed tollens Iohanan filius Caree et universi principes bellatorum universos reliquiarum Iudae, qui reversi fuerant de cunctis gentibus, ad quas fuerant ante dispersi, ut peregrinarentur in terra Iudae,
JER|43|6|viros et mulieres et parvulos et filias regis et omnem animam, quam reliquerat Nabuzardan princeps satellitum cum Godolia filio Ahicam filii Saphan, et Ieremiam prophetam et Baruch filium Neriae,
JER|43|7|et ingressi sunt terram Aegypti, quia non oboedierunt voci Domini; et venerunt usque ad Taphnas.
JER|43|8|Et factus est sermo Domini ad Ieremiam in Taphnis dicens:
JER|43|9|" Sume lapides grandes in manu tua et absconde eos in caemento, sub pavimento, quod est ad portam domus pharaonis in Taphnis, cernentibus viris Iudaeis;
JER|43|10|et dices ad eos: Haec dicit Dominus exercituum, Deus Israel: Ecce ego mittam et assumam Nabuchodonosor regem Babylonis servum meum et ponam thronum eius super lapides istos, quos abscondi, et statuet solium suum super eos;
JER|43|11|veniensque percutiet terram Aegypti, quos in mortem, in mortem et, quos in captivitatem, in captivitatem et, quos in gladium, in gladium;
JER|43|12|et succendet ignem in delubris deorum Aegypti et comburet ea et captivos ducet illos et excutiet terram Aegypti, sicut pastor pediculis excutit pallium suum, et egredietur inde in pace;
JER|43|13|et conteret statuas domus Solis, quae sunt in terra Aegypti, et delubra deorum Aegypti comburet igni ".
JER|44|1|Verbum, quod factum est per Ieremiam ad omnes Iudaeos, qui habitabant in terra Aegypti, habitantes in Magdolo et in Taphnis et in Memphi et in terra Phatures, dicens:
JER|44|2|" Haec dicit Dominus exercituum, Deus Israel: Vos vidistis omne malum istud, quod adduxi super Ierusalem et super omnes urbes Iudae; et ecce desertae sunt hodie, et non est in eis habitator
JER|44|3|propter malitiam, quam fecerunt, ut me ad iracundiam provocarent et irent, ut sacrificarent et colerent deos alienos, quos nesciebant et illi et vos et patres vestri.
JER|44|4|Et misi ad vos omnes servos meos prophetas, de nocte consurgens mittensque et dicens: Nolite facere verbum abominationis huiuscemodi, quam odivi.
JER|44|5|Et non audierunt nec inclinaverunt aurem suam, ut converterentur a malis suis et non sacrificarent diis alienis;
JER|44|6|et effusa est indignatio mea et furor meus et succensa est in civitatibus Iudae et in plateis Ierusalem, et versae sunt in solitudinem et vastitatem secundum diem hanc.
JER|44|7|Et nunc haec dicit Dominus exercituum, Deus Israel: Quare vos facitis malum grande contra animas vestras, ut intereat ex vobis vir et mulier, parvulus et lactans de medio Iudae, nec relinquatur vobis quidquam residuum,
JER|44|8|provocantes me in operibus manuum vestrarum, sacrificando diis alienis in terra Aegypti, in quam ingressi estis, ut ibi peregrinemini, et dissipet vos, et sitis in maledictionem et in opprobrium cunctis gentibus terrae?
JER|44|9|Numquid obliti estis mala patrum vestrorum et mala regum Iudae et mala uxorum eius et mala vestra et mala uxorum vestrarum, quae fecerunt in terra Iudae et in plateis Ierusalem?
JER|44|10|Non sunt contriti usque ad diem hanc et non timuerunt et non ambulaverunt in lege mea et in praeceptis meis, quae dedi coram vobis et coram patribus vestris.
JER|44|11|Ideo haec dicit Dominus exercituum, Deus Israel: Ecce ego ponam faciem meam in vobis in malum et disperdam omnem Iudam.
JER|44|12|Et assumam reliquias Iudae, qui posuerunt facies suas, ut ingrederentur terram Aegypti et peregrinarentur ibi, et consumentur omnes in terra Aegypti: cadent in gladio et in fame et consumentur a minimo usque ad maximum, in gladio et in fame morientur; et erunt in exsecrationem et in stuporem et in maledictionem et in opprobrium.
JER|44|13|Et visitabo super habitatores terrae Aegypti, sicut visitavi super Ierusalem, in gladio et in fame et in peste:
JER|44|14|et non erit qui effugiat et sit residuus de reliquiis Iudaeorum, qui venerunt, ut peregrinarentur in terra Aegypti et reverterentur in terram Iudae, ad quam ipsi elevant animas suas, ut revertantur et habitent ibi; non revertentur, nisi qui fugerint ".
JER|44|15|Responderunt autem Ieremiae omnes viri, scientes quod sacrificarent uxores eorum diis alienis, et universae mulieres, quarum stabat multitudo grandis, et omnis populus habitantium in terra Aegypti in Phatures, dicentes:
JER|44|16|" Sermonem, quem locutus es ad nos in nomine Domini, non audiemus ex te,
JER|44|17|sed facientes faciemus omne verbum, quod egressum est de ore nostro, ut sacrificemus reginae caeli et libemus ei libamina, sicut fecimus nos et patres nostri, reges nostri et principes nostri in urbibus Iudae et in plateis Ierusalem, et saturati sumus panibus et bene nobis erat malumque non vidimus.
JER|44|18|Ex eo autem tempore, quo cessavimus sacrificare reginae caeli et libare ei libamina, indigemus omnibus et gladio et fame consumpti sumus.
JER|44|19|Quod si nos sacrificamus reginae caeli et libamus ei libamina, numquid sine viris nostris fecimus ei placentas ad effingendum eam et libandum ei libamina? ".
JER|44|20|Et dixit Ieremias ad omnem populum, adversum viros et adversum mulieres et adversum universam plebem, qui responderant ei verbum, dicens:
JER|44|21|" Numquid non sacrificium, quod sacrificastis in civitatibus Iudae et in plateis Ierusalem, vos et patres vestri, reges vestri et principes vestri et populus terrae, horum recordatus est Dominus, et ascendit super cor eius?
JER|44|22|Et non poterat Dominus ultra portare propter malitiam operum vestrorum et propter abominationes, quas fecistis; et facta est terra vestra in desolationem et in stuporem et in maledictum, eo quod non sit habitator, sicut est dies haec.
JER|44|23|Propterea quod sacrificaveritis et peccaveritis Domino et non audieritis vocem Domini et in lege et in praeceptis et in testimoniis eius non ambulaveritis, idcirco evenerunt vobis mala haec, sicut est dies haec.
JER|44|24|Dixit autem Ieremias ad omnem populum et ad universas mulieres: " Audite verbum Domini, omnis Iuda, qui estis in terra Aegypti.
JER|44|25|Haec dicit Dominus exercituum, Deus Israel, dicens: Vos et uxores vestrae locuti estis ore vestro et manibus vestris implestis dicentes: Faciamus vota nostra, quae vovimus, ut sacrificemus reginae caeli et libemus ei libamina". Implete vota vestra et opere perpetrate ea.
JER|44|26|Ideo audite verbum Domini, omnis Iuda, qui habitatis in terra Aegypti: Ecce ego iuravi in nomine meo magno, ait Dominus, quia nequaquam ultra vocabitur nomen meum ex ore omnis viri Iudae dicentis: "Vivit Dominus Deus", in omni terra Aegypti.
JER|44|27|Ecce ego vigilabo super eos in malum et non in bonum, et consumentur omnes viri Iudae, qui sunt in terra Aegypti, gladio et fame, donec penitus consumantur.
JER|44|28|Et, qui fugerint gladium, revertentur de terra Aegypti in terram Iudae, viri pauci, et scient omnes reliquiae Iudae, quae ingressae sunt terram Aegypti, ut peregrinarentur ibi, cuius sermo compleatur, meus an illorum.
JER|44|29|Et hoc vobis signum, ait Dominus, quod visitem ego super vos in loco isto, ut sciatis quia vere complebuntur sermones mei contra vos in malum.
JER|44|30|Haec dicit Dominus: Ecce ego tradam pharaonem Ophree, regem Aegypti, in manu inimicorum eius et in manu quaerentium animam illius, sicut tradidi Sedeciam regem Iudae in manu Nabuchodonosor regis Babylonis inimici sui et quaerentis animam eius ".
JER|45|1|Verbum, quod locutus est Ieremias propheta ad Baruch filium Neriae, cum scriberet verba haec in libro ex ore Ieremiae, anno quarto Ioachim filii Iosiae regis Iudae, dicens:
JER|45|2|" Haec dicit Dominus, Deus Israel, super te, Baruch.
JER|45|3|Dixisti: "Vae misero mihi, quoniam addidit Dominus dolorem maerori meo; laboravi in gemitu meo et requiem non inveni".
JER|45|4|Haec dices ad eum: Sic dicit Dominus: Ecce, quod aedificavi, ego destruo et, quod plantavi, ego evello, universam terram hanc;
JER|45|5|et tu quaeris tibi grandia? Noli quaerere, quia ecce ego adducam malum super omnem carnem, ait Dominus, et dabo tibi animam tuam quasi spolium in omnibus locis, ad quaecumque perrexeris ".
JER|46|1|Quod factum est verbum Domini ad Ieremiam prophetam contra gentes.
JER|46|2|Ad Aegyptum.Adversum exercitum pharaonis Nechao regis Aegypti, qui erat iuxta fluvium Euphraten in Charchamis, quem percussit Nabuchodonosor rex Babylonis in quarto anno Ioachim filii Iosiae regis Iudae.
JER|46|3|" Praeparate scutum et clipeumet procedite ad bellum.
JER|46|4|Iungite equos et ascendite, equites;state in galeis, polite lanceas, induite vos loricis.
JER|46|5|Quid igitur? Vidi ipsos pavidos et terga vertentes,fortes eorum caesos;fugerunt conciti nec respexerunt:terror undique,ait Dominus.
JER|46|6|Non fugiat velox,nec salvari se putet fortis;ad aquilonem iuxta flumen Euphratenvicti sunt et ruerunt.
JER|46|7|Quis est iste, qui quasi Nilus ascendit,et veluti fluviorum intumescunt gurgites eius?
JER|46|8|Aegyptus Nili instar ascendit,et velut flumina moventur fluctus eius,et dixit: "Ascendens operiam terram,perdam civitatem et habitatores eius".
JER|46|9|Ascendite, equi, et irruite, currus;et procedant fortes,Aethiopia et Phut tenentes scutum et Ludii arripientes et iacientes sagittas.
JER|46|10|Dies autem ille Domini, Dei exercituum, dies ultionis,ut sumat vindictam de inimicis suis: devorat gladius, et saturatur,et inebriatur sanguine eorum;victima enim Domini, Dei exercituum,in terra aquilonis iuxta flumen Euphraten.
JER|46|11|Ascende in Galaad et tolle resinam,virgo filia Aegypti;frustra multiplicas medicamina,tibi vero cicatrix non obducitur.
JER|46|12|Audierunt gentes ignominiam tuam, et ululatus tuus replevit terram,quia fortis impegit in fortem,et ambo pariter conciderunt ".
JER|46|13|Verbum, quod locutus est Dominus ad Ieremiam prophetam super eo quod veniret Nabuchodonosor rex Babylonis percussurus terram Aegypti.
JER|46|14|" Annuntiate Aegyptoet auditum facite in Magdolo,et resonet in Memphi et in Taphnis,dicite: "Sta et praepara te,quia devoravit gladius ea,quae per circuitum tuum sunt".
JER|46|15|Quare deiectus est fortis tuus?Non stetit, quoniam Dominus subvertit eum.
JER|46|16|Multiplicavit ruentes,ceciditque vir ad proximum suum, et dixerunt: "Surge,et revertamur ad populum nostrumet ad terram nativitatis nostrae,a facie gladii saevientis".
JER|46|17|Vocate nomen pharaonis regis Aegypti:Tumultum, qui praetermisit tempus opportunum.
JER|46|18|Vivo ego, inquit rex,Dominus exercituum nomen eius,quoniam sicut Thabor in montibuset sicut Carmelus ad mare veniet.
JER|46|19|Vasa transmigrationis fac tibi,habitatrix filia Aegypti,quia Memphis in solitudinem eritet destruetur et inhabitabilis erit.
JER|46|20|Vitula elegans atque formosa Aegyptus,stimulus ab aquilone venit ei.
JER|46|21|Mercennarii quoque eius,qui versabantur in medio eius quasi vituli saginati,versi sunt et fugerunt simulnec stare potuerunt,quia dies interfectionis eorum venit super eos,tempus visitationis eorum.
JER|46|22|Vox eius quasi serpentis sibilantis,quoniam cum exercitu properabunt et cum securibus venient ei,quasi caedentes ligna.
JER|46|23|Succiderunt saltum eius,ait Dominus,qui supputari non potest;multiplicati sunt enim super locustas,et non est eis numerus.
JER|46|24|Confusa est filia Aegyptiet tradita in manu populi aquilonis ".
JER|46|25|Dixit Dominus exercituum, Deus Israel: " Ecce ego visitabo super Amon de No et super pharaonem et super Aegyptum et super deos eius et super reges eius et super pharaonem et super eos, qui confidunt in eo;
JER|46|26|et dabo eos in manu quaerentium animam eorum et in manu Nabuchodonosor regis Babylonis et in manu servorum eius; et post haec habitabitur sicut diebus pristinis, ait Dominus.
JER|46|27|Et tu ne timeas, serve meus Iacob,et ne paveas, Israel,quia ecce ego salvum te faciam de longinquoet semen tuum de terra captivitatis eorum;et revertetur Iacob et requiescet,securus erit, et non erit qui exterreat eum.
JER|46|28|Et tu noli timere, serve meus Iacob,ait Dominus,quia tecum ego sum,quia ego consumam cunctas gentes, ad quas eieci te;te vero non consumam,sed castigabo te in iudicionec quasi innocenti parcam tibi ".
JER|47|1|Quod factum est verbum Domini ad Ieremiam prophe tam contra Philisthim, antequam percuteret pharao Gazam.
JER|47|2|Haec dicit Dominus: Ecce, aquae ascendunt ab aquiloneet erunt quasi torrens inundanset operient terram et plenitudinem eius,urbem et habitatores eius.Clamabunt homines,et ululabunt omnes habitatores terrae
JER|47|3|a strepitu ungularum fortium equorum eius,a commotione quadrigarum eiuset tumultu rotarum illius;non respexerunt patres filios, manibus dissolutis,
JER|47|4|pro adventu diei, in quo vastabuntur omnes Philisthim,et dissipabitur Tyro et Sidoni omnis superstes auxiliator:depopulatus est enim Dominus Philisthim,reliquias insulae Caphtor.
JER|47|5|Venit calvitium super Gazam,conticuit Ascalon;reliquiae Enacim,usquequo incidetis vos?
JER|47|6|O mucro Domini,usquequo non quiesces?Ingredere in vaginam tuam,refrigerare et sile.
JER|47|7|Quomodo quiescet,cum Dominus praeceperit ei adversus Ascalonemet adversus maritimas regionesibique condixerit illi? ".
JER|48|1|Ad Moab.Haec dicit Dominus exercituum, Deus Israel: Vae super Nabo, quoniam vastata est et confusa!Capta est Cariathaim, confusa est arx et tremuit.
JER|48|2|Non est ultra exsultatio in Moab;in Hesebon cogitaverunt malum contra eam:Venite et disperdamus eam de gente".Tu quoque, Madmen, conticesces, sequeturque te gladius.
JER|48|3|Vox clamoris de Oronaim:Vastitas et contritio magna".
JER|48|4|Contrita est Moab,auditum fecerunt clamorem usque ad Segor.
JER|48|5|Per ascensum enim Luithplorans ascendit in fletu,quoniam in descensu Oronaimhostes ululatum contritionis audierunt:
JER|48|6|"Fugite, salvate animas vestraset eritis quasi myricae in deserto".
JER|48|7|Pro eo enim quod habuisti fiduciamin operibus tuis et in thesauris tuis,tu quoque capieris;et ibit Chamos in transmigrationem,sacerdotes eius et principes eius simul.
JER|48|8|Et veniet praedo ad omnem urbem, et urbs nulla salvabitur;et peribit vallis, et dissipabuntur campestria,quoniam dixit Dominus.
JER|48|9|Date pennas ad volandum;et civitates eius desertae erunt et inhabitabiles.
JER|48|10|Maledictus, qui facit opus Domini neglegenter,et maledictus, qui prohibet gladium suum a sanguine.
JER|48|11|Securus fuit Moab ab adulescentia suaet requievit in faecibus suisnec transfusus est de vase in vaset in transmigrationem non abiit;idcirco permansit gustus eius in eo,et odor eius non est immutatus.
JER|48|12|Propterea, ecce, dies veniunt,dicit Dominus,et mittam ei stratores laguncularum;et sternent eumet vasa eius exhaurientet lagunculas eorum collident.
JER|48|13|Et confundetur Moab a Chamos, sicut confusa est domus Israel a Bethel, in qua habebat fiduciam.
JER|48|14|Quomodo dicitis: "Fortes sumuset viri robusti ad proeliandum"?
JER|48|15|Vastata est Moab,et ascenderunt civitates illius,et electi iuvenes eius descenderunt in occisionem,ait rex, Dominus exercituum nomen eius.
JER|48|16|Prope est interitus Moab ut veniat,et malum eius velociter accurret nimis.
JER|48|17|Lugete super eum,omnes, qui estis in circuitu eius;et universi, qui scitis nomen eius,dicite: "Quomodo confracta est virga fortis,baculus gloriosus?".
JER|48|18|Descende de gloria et sede in siti,habitatrix filia Dibon,quoniam vastator Moab ascendit ad te,dissipavit munitiones tuas.
JER|48|19|Ad viam sta et prospice,habitatrix Aroer;interroga fugientemet eam, quae evasit.Dic: "Quid accidit?".
JER|48|20|Confusus est Moab, quoniam victus est.Ululate et clamate;annuntiate in Arnon,quoniam vastatus est Moab.
JER|48|21|Et iudicium venit ad terram campestrem super Helon et super Iasa et super Mephaath
JER|48|22|et super Dibon et super Nabo et super Bethdeblathaim,
JER|48|23|et super Cariathaim et super Bethgamul et super Bethmaon
JER|48|24|et super Carioth et super Bosra et super omnes civitates terrae Moab, quae longe et quae prope sunt.
JER|48|25|Abscissum est cornu Moab,et brachium eius contritum est,ait Dominus.
JER|48|26|Inebriate eum, quoniam contra Dominum erectus est; et allidet manum Moab in vomitu suo, et erit in derisum etiam ipse.
JER|48|27|Nonne in derisum tibi fuit Israel? Num inter fures repertus est? Quotiescumque enim adversum illum loquebaris, caput movebas.
JER|48|28|Relinquite civitates et habitate in petra,habitatores Moab,et estote quasi columba nidificansin parietibus apertae voraginis.
JER|48|29|Audivimus superbiam Moab,superbus est valde;sublimitatem eius et arrogantiamet superbiam et altitudinem cordis eius.
JER|48|30|Ego scio, ait Dominus, iactantiam eius, et quod non sint rectae fabulationes, nec recta fecerint.
JER|48|31|Ideo super Moab eiulabo et super Moab universam clamabo, super viros Cirhareseth plorabitur.
JER|48|32|Plus quam in planctu Iazer plorabo tibi,vinea Sabama;propagines tuae transierunt mare,usque ad Iazer pervenerunt.Super messem tuam et vindemiam tuampraedo irruit.
JER|48|33|Ablata est laetitia et exsultatiode horto et de terra Moab,et vinum de torcularibus sustuli;nequaquam calcator uvaesolitum celeuma cantabit.
JER|48|34|De clamore Hesebon usque Eleale et Iasa dederunt vocem suam, a Segor usque ad Oronaim, ad Eglatselisiam; aquae quoque Nemrim pessimae erunt.
JER|48|35|Et auferam de Moab, ait Dominus, offerentem in excelsis et sacrificantem diis eius.
JER|48|36|Propterea cor meum ad Moab quasi tibia resonabit, et cor meum ad viros Cirhareseth dabit sonitum tibiarum; quia depositum, quod acquisierunt, periit.
JER|48|37|Omne enim caput calvitium et omnis barba rasa erit, in cunctis manibus incisiones et super lumbos cilicium.
JER|48|38|Super omnia tecta Moab et in plateis eius omnis planctus, quoniam contrivi Moab sicut vas, quod nemini placet, ait Dominus.
JER|48|39|Quomodo victa est, et ululaverunt? Quomodo vertit dorsum Moab et confusus est? Eritque Moab in derisum et in terrorem omnibus in circuitu suo.
JER|48|40|Haec dicit Dominus:Ecce quasi aquila volabitet extendet alas suas ad Moab.
JER|48|41|Capta sunt oppida,et munitiones comprehensae sunt,et erit cor fortium Moab in die illasicut cor mulieris parturientis.
JER|48|42|Et cessabit Moab esse populus,quoniam contra Dominum gloriatus est.
JER|48|43|Pavor et fovea et laqueus super te,o habitator Moab,dicit Dominus.
JER|48|44|Qui fugerit a facie pavoris, cadet in foveam,et, qui conscenderit de fovea, capietur laqueo;adducam enim super Moabannum visitationis eorum,ait Dominus.
JER|48|45|In umbra Hesebon steterunt sine viribus fugientes,sed ignis egressus est de Hesebon,et flamma de medio Sehon,et devoravit tempora Moabet verticem filiorum tumultus.
JER|48|46|Vae tibi, Moab!Periit populus Chamos,quia comprehensi sunt filii tuiet filiae tuae in captivitatem.
JER|48|47|Et convertam sortem Moab in novissimis diebus ",ait Dominus.Hucusque iudicia Moab.
JER|49|1|Ad filios Ammon.Haec dicit Dominus: Numquid filii non sunt Israel,aut heres non est ei?Cur igitur hereditate possedit Melchom Gad,et populus eius in urbibus eius habitavit?
JER|49|2|Ideo ecce dies veniunt,dicit Dominus,et auditum faciam super Rabba filiorum Ammonfremitum proelii;et erit in tumulum dissipata,filiaeque eius igni succendentur,et possidebit Israel possessores suos, ait Dominus.
JER|49|3|Ulula, Hesebon, quoniam vastata es, ut sis in acervum lapidum;clamate, filiae Rabba,accingite vos ciliciis, plangiteet circuite per muros,quoniam Melchom in transmigrationem ducetur,sacerdotes eius et principes eius simul.
JER|49|4|Quid gloriaris in vallibus?Copiose fluxit vallis tua, filia rebellis,quae confidebas in thesauris tuiset dicebas: "Quis veniet ad me?".
JER|49|5|Ecce ego inducam super te terrorem,ait Dominus, Deus exercituum,ab omnibus, qui sunt in circuitu tuo;et dispergemini singuli in viam suam,nec erit qui congreget fugientes.
JER|49|6|Et post haec convertamsortem filiorum Ammon ",ait Dominus.
JER|49|7|Ad Edom.Haec dicit Dominus exercituum: Numquid non ultra est sapientia in Theman?Periit consilium a prudentibus,inutilis facta est sapientia eorum.
JER|49|8|Fugite, terga vertite, descendite in voraginem,habitatores Dedan,quoniam perditionem Esau adduxi super eum,tempore quo visitavi eum.
JER|49|9|Si vindemiatores veniunt super te,non relinquent racemum;si fures in nocte,diripiunt, quod placet sibi.
JER|49|10|Ego vero discooperui Esau,revelavi abscondita eius,et celari non poterit;vastatum est semen eiuset fratres eius et vicini eius, et non erit.
JER|49|11|Relinque pupillos tuos, ego faciam eos vivere;et viduae tuae in me sperabunt.
JER|49|12|Quia haec dicit Dominus: Ecce quibus non erat iudicium, ut biberent calicem, bibentes bibent; et tu quasi innocens relinqueris? Non eris innocens, sed bibens bibes.
JER|49|13|Quia per memetipsum iuravi, dicit Dominus, quod in solitudinem et in opprobrium et in desertum et in maledictionem erit Bosra; et omnes civitates eius erunt in solitudines sempiternas ".
JER|49|14|Auditum audivi a Domino,et legatus ad gentes missus est: Congregamini et venite contra eamet consurgite in proelium ".
JER|49|15|" Ecce enim parvulum dedi te in gentibus,contemptibilem inter homines.
JER|49|16|Arrogantia tua decepit te,et superbia cordis tui,qui habitas in cavernis petraeet tenes altitudinem collis;cum exaltaveris quasi aquila nidum tuum,inde detraham te,dicit Dominus.
JER|49|17|Et erit Edom in desolationem: omnis, qui transibit per eam, stupebit et sibilabit super omnes plagas eius.
JER|49|18|Sicut subversa est Sodoma et Gomorra et vicinae eius, ait Dominus, non habitabit ibi vir, et non peregrinabitur in ea filius hominis.
JER|49|19|Ecce quasi leo ascendet de silva condensa Iordanis ad prata semper virentia, quia subito currere faciam eos ex illa; et, qui erit electus, illum praeponam ei. Quis enim similis mei? Et quis vocabit me in iudicium? Et quis est iste pastor, qui resistat vultui meo?
JER|49|20|Propterea audite consilium Domini, quod iniit de Edom, et cogitationes eius, quas cogitavit de habitatoribus Theman:Certe abstrahent parvulos gregis,certe desolabuntur super eos pascua eorum.
JER|49|21|A voce ruinae eorum commota est terra,clamor in mari Rubro auditus est ocis eius.
JER|49|22|Ecce quasi aquila ascendet et volabitet expandet alas suas super Bosram;et erit cor fortium Edom in die illaquasi cor mulieris parturientis ".
JER|49|23|Ad Damascum. Confusa est Emath et Arphad,quia auditum pessimum audierunt;turbati sunt in mari sollicitudinis,quod quiescere non potuit.
JER|49|24|Dissoluta est Damascus, versa in fugam;tremor apprehendit eam,angustia et dolores tenuerunt eamquasi parturientem.
JER|49|25|Quomodo non erit derelicta civitas laudabilis,urbs laetitiae?
JER|49|26|Ideo cadent iuvenes eius in plateis eius,et omnes viri proelii conticescent in die illa,ait Dominus exercituum.
JER|49|27|Et succendam ignem in muro Damasci,et devorabit moenia Benadad ".
JER|49|28|Ad Cedar et ad regna Asor, quae percussit Nabuchodonosor rex Babylonis.Haec dicit Dominus: Surgite, ascendite ad Cedaret vastate filios orientis.
JER|49|29|Tabernacula eorum et greges eorum capient;tentoria eorum et omnia vasa eorumet camelos eorum tollent sibi;et vocabunt super eos formidinem in circuitu.
JER|49|30|Fugite, abite vehementer,in voraginibus sedete,qui habitatis Asor,ait Dominus;iniit enim contra vosNabuchodonosor rex Babylonis consiliumet cogitavit adversum vos cogitationes.
JER|49|31|Consurgite, et ascenditead gentem quietam et habitantem confidenter,ait Dominus;non ostia nec vectes eis:soli habitant.
JER|49|32|Et erunt cameli eorum in direptionem,et multitudo iumentorum in praedam;et dispergam eos in omnem ventum, qui sunt attonsi in comam,et ex omni confinio eorumadducam interitum super eos,ait Dominus.
JER|49|33|Et erit Asor in habitaculum thoum,deserta usque in aeternum;non manebit ibi vir,nec peregrinabitur in ea filius hominis ".
JER|49|34|Quod factum est verbum Domini ad Ieremiam prophetam super Elam, in principio regni Sedeciae regis Iudae, dicens:
JER|49|35|" Haec dicit Dominus exercituum:Ecce ego confringam arcum Elam, summam fortitudinem eorum;
JER|49|36|et inducam super Elamquattuor ventos a quattuor plagis caeli,et ventilabo eos in omnes ventos istos,et non erit gens,ad quam non perveniant profugi Elam.
JER|49|37|Et pavere faciam Elam coram inimicis suiset in conspectu quaerentium animam eorum;et adducam super eos malumiram furoris mei,dicit Dominus,et mittam post eos gladium,donec consumam eos.
JER|49|38|Et ponam solium meum in Elamet perdam inde regem et principes, ait Dominus.
JER|49|39|In novissimis autem diebusconvertam sortem Elam ",dicit Dominus.
JER|50|1|Verbum, quod locutus est Dominus de Babylone et de terra Chaldaeorum in manu Ieremiae prophetae:
JER|50|2|" Annuntiate in gentibus et auditum facite,levate signum;praedicate et nolite celare, dicite:Capta est Babylon,confusus est Bel,victus est Merodach.Confusa sunt sculptilia eius,superata sunt idola eorum".
JER|50|3|Quoniam ascendit contra eam gens ab aquilone, quae ponet terram eius in solitudinem, et non erit qui habitet in ea ab homine usque ad pecus: et moti sunt et abierunt.
JER|50|4|In diebus illis et in tempore illo, ait Dominus, venient filii Israel ipsi et filii Iudae simul; ambulantes et flentes properabunt et Dominum Deum suum quaerent.
JER|50|5|De Sion interrogabunt, ad cuius viam facies eorum: "Venite, et apponamur ad Dominum foedere sempiterno, quod nulla oblivione delebitur".
JER|50|6|Grex perditus factus est populus meus, pastores eorum seduxerunt eos feceruntque vagari in montibus; de monte in collem transierunt, obliti sunt cubilis sui.
JER|50|7|Omnes, qui invenerunt, comederunt eos, et hostes eorum dixerunt: "Non delinquimus, pro eo quod peccaverunt Domino, habitaculo iustitiae et exspectationi patrum eorum Domino".
JER|50|8|Recedite de medio Babyloniset de terra Chaldaeorum egredimini;et estote quasi haedi ante gregem.
JER|50|9|Quoniam ecce ego suscito et adducam in Babylonemcongregationem gentium magnarumde terra aquilonis;et praeparabuntur adversus eam,et inde capietur:sagitta eorum quasi bellatoris electinon revertetur vacua.
JER|50|10|Et erit Chaldaea in praedam;omnes vastantes eam replebuntur ",ait Dominus.
JER|50|11|Dum exsultatis et magna loquiminidiripientes hereditatem meamdum effusi estis sicut vituli super herbamet hinnitis sicut equi fortes,
JER|50|12|confusa est mater vestra nimis,et in opprobrium facta est, quae genuit vos;ecce novissima erit in gentibus,deserta, invia et arens.
JER|50|13|Ab ira Domini non habitabitur,sed redigetur tota in solitudinem;omnis, qui transibit per Babylonem, stupebitet sibilabit super universis plagis eius.
JER|50|14|Praeparamini contra Babylonem per circuitumomnes, qui tenditis arcum;debellate eam, non parcatis iaculis,quia Domino peccavit.
JER|50|15|Clamate adversus eam;ubique dedit manum,ceciderunt fundamenta eius,destructi sunt muri eius,quoniam ultio Domini est;ultionem accipite de ea:sicut fecit, facite ei.
JER|50|16|Disperdite satorem de Babyloneet tenentem falcem in tempore messis;a facie gladii saevientisunusquisque ad populum suum convertetur,et singuli ad terram suam fugient.
JER|50|17|Ovis dispersa Israel;leones eiecerunt eum.Primus comedit eum rex Assyriae;iste novissimus exossavit eumNabuchodonosor rex Babylonis.
JER|50|18|Propterea haec dicit Dominus exercituum, Deus Israel: " Ecce ego visitabo regem Babylonis et terram eius, sicut visitavi regem Assyriae;
JER|50|19|et reducam Israel ad pascua sua, et pascetur Carmelum et Basan, et in monte Ephraim et Galaad saturabitur anima eius.
JER|50|20|In diebus illis et in tempore illo, ait Dominus, quaeretur iniquitas Israel et non erit, et peccatum Iudae et non invenietur, quoniam propitius ero eis, quos reliquero.
JER|50|21|Super terram Merataim ascendeet super habitatores Phacud.Dissipa et interfice persequens eos,ait Dominus,et fac iuxta omnia, quae praecepi tibi ".
JER|50|22|Vox belli in terraet contritio magna.
JER|50|23|Quomodo confractus est et contritusmalleus universae terrae?Quomodo versa est in desolationem Babylon in gentibus?
JER|50|24|Illaqueavi te, et capta es, Babylon,et nesciebas;inventa es et apprehensa,quoniam Dominum provocasti.
JER|50|25|Aperuit Dominus thesaurum suumet protulit vasa irae suae,quoniam opus est Domino Deo exercituumin terra Chaldaeorum.
JER|50|26|Venite ad eam ab extremis finibus,aperite horrea eius;redigite eam in acervos lapidum quasi manipuloset interficite eam,nec sit quidquam reliquum.
JER|50|27|Dissipate universos tauros eius,descendant in occisionem.Vae eis, quia venit dies eorum,tempus visitationis eorum!
JER|50|28|Vox fugientiumet eorum, qui evaserunt de terra Babylonis,ut annuntient in Sionultionem Domini Dei nostri,ultionem templi eius.
JER|50|29|Convocate in Babylonem sagittarios,omnes, qui tendunt arcum;consistite adversus eam per gyrum, et nullus evadat:reddite ei secundum opus suum,iuxta omnia, quae fecit, facite illi,quia contra Dominum erecta est,adversum Sanctum Israel.
JER|50|30|" Idcirco cadent iuvenes eius in plateis eius,et omnes viri bellatores eius conticescent in die illa,ait Dominus.
JER|50|31|Ecce ego ad te, Superbia,dicit Dominus, Deus exercituum,quia venit dies tuus,tempus visitationis tuae.
JER|50|32|Et cadet Superbia et corruet,et non erit qui suscitet eam;et succendam ignem in urbibus eius,et devorabit omnia in circuitu eius ".
JER|50|33|Haec dicit Dominus exercituum: " Calumniam sustinent filii Israel et filii Iudae simul; omnes, qui ceperunt eos, tenent, nolunt dimittere eos.
JER|50|34|Redemptor eorum fortis, Dominus exercituum nomen eius, iudicio defendet causam eorum, ut quietem det terrae et conturbet habitatores Babylonis.
JER|50|35|Gladius ad Chaldaeos,ait Dominus,et ad habitatores Babyloniset ad principes et ad sapientes eius!
JER|50|36|Gladius ad divinos eius, qui stulti erunt!Gladius ad fortes illius, qui timebunt!
JER|50|37|Gladius ad equos eius et ad currus eiuset ad omne vulgus, quod est in medio eius;et erunt quasi mulieres!Gladius ad thesauros eius, qui diripientur!
JER|50|38|Siccitas super aquas eius erit, et arescent,quia terra sculptilium est,et in portentis insaniunt.
JER|50|39|Propterea habitabunt dracones cum thoibus, et habitabunt in ea struthiones; et non inhabitabitur ultra usque in sempiternum nec exstruetur usque ad generationem et generationem.
JER|50|40|Sicut subvertit Deus Sodomam et Gomorram et vicinas eius, ait Dominus, non habitabit ibi vir, et non peregrinabitur in ea filius hominis.
JER|50|41|Ecce populus venit ab aquilone, et gens magna et reges multi consurgent a finibus terrae.
JER|50|42|Arcum et acinacem apprehendent, crudeles sunt et immisericordes; vox eorum quasi mare sonabit, et super equos ascendent sicut vir paratus ad proelium contra te, filia Babylon.
JER|50|43|Audivit rex Babylonis famam eorum, et dissolutae sunt manus eius; angustia apprehendit eum, dolor quasi parturientem.
JER|50|44|Ecce quasi leo ascendet de silva condensa Iordanis ad prata semper virentia, quia subito currere faciam eos ex illa et, qui erit electus, illum praeponam ei. Quis enim similis mei? Et quis vocabit me in iudicium? Et quis est iste pastor, qui resistat vultui meo? ".
JER|50|45|Propterea audite consilium Domini, quod mente concepit adversum Babylonem, et cogitationes eius, quas cogitavit super terram Chaldaeorum: certe abstrahent parvulos gregis, certe desolabuntur super eos pascua eorum.
JER|50|46|A voce captivitatis Babylonis commota est terra, et clamor inter gentes auditus est.
JER|51|1|Haec dicit Dominus: Ecce ego suscitabo super Babylonemet super habitatores Chaldaeaequasi ventum pestilentem;
JER|51|2|et mittam in Babylonem ventilatores,et ventilabunt eamet demolientur terram eius,quoniam venerunt super eam undiquein die afflictionis.
JER|51|3|Non tendat, qui tendit arcum suum,et non ascendat loricatus;nolite parcere iuvenibus eius,interficite omnem militiam eius ".
JER|51|4|Et cadent interfecti in terra Chaldaeorumet vulnerati in plateis eius,
JER|51|5|quoniam non est viduatus Israel et Iudaa Deo suo, Domino exercituum;terra autem eorum repleta est delictoin conspectu Sancti Israel.
JER|51|6|Fugite de medio Babylonis,et salvet unusquisque animam suam;nolite perire in poena eius,quoniam tempus ultionis est Domino:vicissitudinem ipse retribuet ei.
JER|51|7|Calix aureus Babylon in manu Dominiinebrians omnem terram;de vino eius biberunt genteset ideo insaniunt.
JER|51|8|Subito cecidit Babylon et contrita est.Ululate super eam;tollite resinam ad dolorem eius,si forte sanetur.
JER|51|9|" Curavimus Babylonem,et non est sanata.Derelinquite eam,et eamus unusquisque in terram suam,quoniam pervenit usque ad caelos iudicium eiuset elevatum est usque ad nubes.
JER|51|10|Protulit Dominus iustitias nostras;venite, et narremus in Sionopus Domini Dei nostri ".
JER|51|11|Acuite sagittas, implete pharetras;suscitavit Dominus spiritum regum Medorum,et contra Babylonem mens eius est, ut perdat eam,quoniam ultio Dominiest ultio templi sui.
JER|51|12|Super muros Babylonis levate signum,augete custodiam,ponite custodes, praeparate insidias,quia cogitavit Dominus,et facit quaecumque locutus estcontra habitatores Babylonis.
JER|51|13|Quae habitas super aquas multas,locuples in thesauris,venit finis tuus,pedalis praecisionis tuae.
JER|51|14|Iuravit Dominus exercituum per animam suam: Quoniam, etsi replevero te hominibus quasi brucho,super te celeuma cantabitur ".
JER|51|15|Qui fecit terram in fortitudine sua,praeparavit orbem in sapientia sua et prudentia sua extendit caelos;
JER|51|16|dante eo vocem, multiplicantur aquae in caelo;qui levat nubes ab extremo terrae,fulgura in pluviam facitet producit ventum de thesauris suis.
JER|51|17|Stultus factus est omnis homo, absque scientia;confusus est omnis conflator in sculptili,quia mendax conflatio eius,nec est spiritus in eis.
JER|51|18|Vana sunt opera et risu digna,in tempore visitationis suae peribunt.
JER|51|19|Non sicut haec pars Iacob,quia, qui fecit omnia, ipse est,et Israel tribus hereditatis eius:Dominus exercituum nomen eius.
JER|51|20|" Malleus tu mihi, vas belli:et ego collisi in te genteset dispersi in te regna
JER|51|21|et collisi in te equum et equitem eiuset collisi in te currum et ascensorem eius
JER|51|22|et collisi in te virum et mulieremet collisi in te senem et puerumet collisi in te iuvenem et virginem
JER|51|23|et collisi in te pastorem et gregem eiuset collisi in te agricolam et iugales eiuset collisi in te duces et magistratus.
JER|51|24|Et reddam Babyloni et cunctis habitatoribus Chaldaeae omne malum suum, quod fecerunt in Sion in oculis vestris, ait Dominus.
JER|51|25|Ecce ego ad te, mons pestifer,ait Dominus,qui corrumpis universam terram;et extendam manum meam super teet evolvam te de petriset dabo te in montem combustionis.
JER|51|26|Et non tollent de te lapidem in angulumet lapidem in fundamenta,sed perditus in aeternum eris ",ait Dominus.
JER|51|27|Levate signum in terra,clangite bucina in gentibus,sanctificate super eam gentes,vocate contra illam regnaArarat, Menni et Aschenez.Constituite super eam scribas,adducite equos quasi bruchum aculeatum.
JER|51|28|Sanctificate contra eam gentes, reges Mediae, duces eius et universos magistratus eius cunctamque terram potestatis eius.
JER|51|29|Et commovebitur terra et conturbabitur,quia impletur contra Babylonem cogitatio Domini,ut ponat terram Babylonisdesertam et inhabitabilem.
JER|51|30|Cessaverunt fortes Babylonis a proelio,habitaverunt in praesidiis;devoratum est robur eorum,et facti sunt quasi mulieres;incensa sunt tabernacula eius,contriti sunt vectes eius.
JER|51|31|Currens obviam currenti veniet,et nuntius obvius nuntianti,ut annuntiet regi Babylonisquia capta est civitas eiusa summo usque ad summum.
JER|51|32|Et vada praeoccupata sunt,et paludes incensae sunt igni;et viri bellatores conturbati sunt.
JER|51|33|Quia haec dicit Dominus exercituum, Deus Israel: Filia Babylonis quasi area tempore triturae eius;adhuc modicum, et veniet tempus messionis eius ".
JER|51|34|" Comedit me, devoravit me Nabuchodonosor;rex Babylonis reddidit me quasi vas inane,absorbuit me quasi draco,replevit ventrem suum deliciis meis et eiecit me ".
JER|51|35|" Iniquitas adversum me et caro mea super Babylonem! ",dicit habitatio Sion. Et sanguis meus super habitatores Chaldaeae! ",dicit Ierusalem.
JER|51|36|Propterea haec dicit Dominus: Ecce ego iudicabo causam tuamet ulciscar ultionem tuamet desertum faciam mare eiuset siccabo venam eius;
JER|51|37|et erit Babylon in tumulos,habitatio thoum,stupor et sibilus,eo quod non sit habitator.
JER|51|38|Simul ut leones rugient,frement veluti catuli leonum.
JER|51|39|In calore eorum ponam potus eorumet inebriabo eos, ut sopianturet dormiant somnum sempiternum et non consurgant,dicit Dominus.
JER|51|40|Deducam eos quasi agnos ad victimam,quasi arietes cum haedis ".
JER|51|41|Quomodo capta est Babel,et comprehensa est gloria universae terrae?Quomodo facta est in stuporemBabylon inter gentes?
JER|51|42|Ascendit super Babylonem mare,multitudine fluctuum eius operta est.
JER|51|43|Factae sunt civitates eius in stuporem,terra inhabitabilis et deserta,terra, in qua nullus habitet,nec transeat per eam filius hominis.
JER|51|44|" Et visitabo super Bel in Babyloneet eiciam, quod absorbuerat, de ore eius;et non confluent ad eum ultra gentes,siquidem et murus Babylonis corruet.
JER|51|45|Egredimini de medio eius, populus meus,ut salvet unusquisque animam suamab ira furoris Domini.
JER|51|46|Et ne forte mollescat cor vestrum, et timeatis auditum, qui audietur in terra; et veniet in anno auditio, et post hunc annum auditio, et iniquitas in terra, et dominator super dominatorem.
JER|51|47|Propterea ecce dies veniunt, et visitabo super sculptilia Babylonis, et omnis terra eius confundetur, et universi interfecti eius cadent in medio eius.
JER|51|48|Et laudabunt super Babylonem caeli et terra et omnia, quae in eis sunt, quia ab aquilone venient ei praedones, ait Dominus.
JER|51|49|Et Babylon cadet, occisi in Israel, sicut pro Babylone ceciderunt occisi universae terrae.
JER|51|50|Qui fugistis gladium, ite, nolite stare; recordamini procul Domini, et Ierusalem ascendat super cor vestrum.
JER|51|51|"Confusi sumus, quoniam audivimus opprobrium; operuit ignominia facies nostras, quia venerunt alieni super sanctificationem domus Domini".
JER|51|52|Propterea ecce dies veniunt, ait Dominus, et visitabo super sculptilia eius, et in omni terra eius gemet vulneratus.
JER|51|53|Si ascenderit Babylon in caelum et firmaverit in excelso robur suum, a me venient vastatores eius ", ait Dominus.
JER|51|54|Vox clamoris de Babylone et contritio magna de terra Chaldaeorum,
JER|51|55|quoniam vastavit Dominus Babylonem et perdidit ex ea vocem magnam; et sonabunt fluctus eorum quasi aquae multae, dedit sonitum vox eorum.
JER|51|56|Quia venit super eam, id est super Babylonem, praedo; et apprehensi sunt fortes eius, et fractus est arcus eorum, quia Deus ultor Dominus reddens retribuet.
JER|51|57|" Et inebriabo principes eius et sapientes eius et duces eius et magistratus eius et fortes eius; et dormient somnum sempiternum et non expergiscentur ", ait rex, Dominus exercituum nomen eius.
JER|51|58|Haec dicit Dominus exercituum: Murus Babylonis ille latissimus funditus suffodietur,et portae eius excelsae igni comburentur;et laboraverunt populi pro nihilo,et gentes pro igni lassatae sunt ".
JER|51|59|Verbum, quod praecepit Ieremias propheta Saraiae filio Neriae filii Maasiae, cum pergeret cum Sedecia rege Iudae in Babylonem in anno quarto regni eius; Saraias autem erat princeps, qui mansionibus praeerat.
JER|51|60|Et scripsit Ieremias omne malum, quod venturum erat super Babylonem, in libro uno, omnia verba haec, quae scripta sunt contra Babylonem.
JER|51|61|Et dixit Ieremias ad Saraiam: " Cum veneris in Babylonem et videris et legeris omnia verba haec,
JER|51|62|dices: "Domine, tu locutus es contra locum istum, ut disperderes eum, ne sit qui in eo habitet ab homine usque ad pecus, et ut sit perpetua solitudo".
JER|51|63|Cumque compleveris legere librum istum, ligabis ad eum lapidem et proicies illum in medium Euphraten
JER|51|64|et dices: "Sic submergetur Babylon et non consurget a facie afflictionis, quam ego adduco super eam, et dissolvetur" ".Hucusque verba Ieremiae.
JER|52|1|Filius viginti et unius anni erat Sedecias, cum regnare coepisset, et undecim annis regnavit in Ierusalem; et nomen matris eius Amital filia Ieremiae de Lobna.
JER|52|2|Et fecit malum in oculis Domini iuxta omnia, quae fecerat Ioachim,
JER|52|3|quoniam furor Domini erat in Ierusalem et in Iuda, usquequo proiceret eos a facie sua.Et recessit Sedecias a rege Babylonis.
JER|52|4|Factum est autem in anno nono regni eius, in mense decimo decima mensis, venit Nabuchodonosor rex Babylonis, ipse et omnis exercitus eius, adversus Ierusalem; et obsederunt eam et aedificaverunt contra eam munitiones in circuitu.
JER|52|5|Et fuit civitas obsessa usque ad undecimum annum regis Sedeciae.
JER|52|6|Mense autem quarto, nona mensis, obtinuit fames in civitate, et non erant alimenta populo terrae.
JER|52|7|Et dirupta est civitas, et omnes viri bellatores fugerunt exieruntque de civitate nocte per viam portae, quae est inter duos muros et ducit ad hortum regis, Chaldaeis obsidentibus urbem in gyro, et abierunt per viam, quae ducit in Arabam.
JER|52|8|Persecutus est autem Chaldaeorum exercitus regem, et apprehenderunt Sedeciam in campestribus Iericho, et omnis comitatus eius diffugit ab eo.
JER|52|9|Cumque comprehendissent regem, adduxerunt eum ad regem Babylonis in Rebla, quae est in terra Emath; et locutus est ad eum iudicia.
JER|52|10|Et iugulavit rex Babylonis filios Sedeciae in oculis eius, sed et omnes principes Iudae occidit in Rebla;
JER|52|11|et oculos Sedeciae eruit et vinxit eum compedibus et adduxit eum rex Babylonis in Babylonem et posuit eum in domo carceris usque ad diem mortis eius.
JER|52|12|In mense autem quinto, decima mensis, ipse est annus nonus decimus Nabuchodonosor regis Babylonis, venit Nabuzardan princeps satellitum, qui stabat coram rege Babylonis, in Ierusalem.
JER|52|13|Et incendit domum Domini et domum regis; et omnes domos Ierusalem et omnem domum magnam igni combussit;
JER|52|14|et totum murum Ierusalem per circuitum destruxit cunctus exercitus Chaldaeorum, qui erat cum magistro satellitum.
JER|52|15|De pauperibus autem populi et de reliquo vulgo, quod remanserat in civitate, et de perfugis, qui transfugerant ad regem Babylonis, et superfluos artificum transtulit Nabuzardan princeps satellitum.
JER|52|16|De pauperibus vero terrae reliquit Nabuzardan princeps satellitum in vinitores et in agricolas.
JER|52|17|Columnas quoque aereas, quae erant in domo Domini, et bases et mare aereum, quod erat in domo Domini, confregerunt Chaldaei et tulerunt omne aes eorum in Babylonem.
JER|52|18|Et lebetes et vatilla et cultros et phialas et mortariola et omnia vasa aerea, quae in ministerio fuerant, tulerunt;
JER|52|19|et pelves et thymiamateria et phialas et lebetes et candelabra et mortaria et cyathos, quotquot aurea aurea, et quotquot argentea argentea, tulit magister satellitum;
JER|52|20|columnas duas et mare unum et vitulos duodecim aereos, qui erant subtus basi, quam fecerat rex Salomon domui Domini. Non erat pondus aeris omnium horum vasorum.
JER|52|21|De columnis autem, decem et octo cubiti altitudinis erant in columna una, et funiculus duodecim cubitorum circuibat eam; porro grossitudo eius quattuor digitorum, et intrinsecus cava erat.
JER|52|22|Et capitella super utramque aerea: altitudo capitelli unius quinque cubitorum, et retiacula et malogranata super capitellum in circuitu omnia aerea; similiter columnae secundae.
JER|52|23|Et malogranata nonaginta sex dependentia; omnia malogranata centum super retiacula in circuitu.
JER|52|24|Et tulit magister satellitum Saraiam sacerdotem primum et Sophoniam sacerdotem secundum et tres custodes vestibuli.
JER|52|25|Et de civitate tulit eunuchum unum, qui erat praepositus super viros bellatores, et septem viros de his, qui videbant faciem regis, qui inventi sunt in civitate, et scribam principis militum, qui ex populo terrae probabat tirones, et sexaginta viros de populo terrae, qui inventi sunt in medio civitatis.
JER|52|26|Tulit autem eos Nabuzardan magister satellitum et duxit eos ad regem Babylonis in Rebla;
JER|52|27|et percussit eos rex Babylonis et interfecit eos in Rebla in terra Emath. Et translatus est Iuda de terra sua.
JER|52|28|Iste est populus, quem transtulit Nabuchodonosor: in anno septimo, Iudaeos tria millia et viginti tres;
JER|52|29|in anno octavo decimo Nabuchodonosor de Ierusalem animas octingentas triginta duas;
JER|52|30|in anno vicesimo tertio Nabuchodonosor transtulit Nabuzardan magister satellitum animas Iudaeorum septingentas quadraginta quinque; omnes ergo animae quattuor milia sescentae.
JER|52|31|Et factum est in tricesimo septimo anno transmigrationis Ioachin regis Iudae, duodecimo mense vicesima quinta mensis, elevavit Evilmerodach rex Babylonis, ipso anno regni sui, caput Ioachin regis Iudae; et eduxit eum de domo carceris.
JER|52|32|Et locutus est cum eo bona et posuit thronum eius super thronos regum, qui erant secum in Babylone.
JER|52|33|Et mutavit vestimenta carceris eius, et comedebat panem coram eo semper cunctis diebus vitae suae.
JER|52|34|Et cibaria eius, cibaria perpetua dabantur ei a rege Babylonis statuta per singulos dies, usque ad diem mortis suae, cunctis diebus vitae eius.
LAM|1|1|ALEPH. Quomodo sedet solacivitas plena populo!Facta est quasi viduadomina gentium;princeps provinciarumfacta est sub tributo.
LAM|1|2|BETH. Plorans plorat in nocte,et lacrimae eius in maxillis eius;non est qui consoletur eamex omnibus caris eius:omnes amici eius spreverunt eamet facti sunt ei inimici.
LAM|1|3|GHIMEL. Migravit Iudas prae afflictioneet multitudine servitutis;habitat inter gentesnec invenit requiem:omnes persecutores eius apprehenderunt eaminter angustias.
LAM|1|4|DALETH. Viae Sion lugent,eo quod non sint qui veniant ad sollemnitatem;omnes portae eius destructae,sacerdotes eius gementes,virgines eius afflictae,et ipsa oppressa amaritudine.
LAM|1|5|HE. Facti sunt hostes eius in caput,inimici eius in securitate,quia Dominus afflixit eampropter multitudinem iniquitatum eius;parvuli eius ducti sunt captiviante faciem tribulantis.
LAM|1|6|VAU. Et egressus est a filia Sionomnis decor eius;facti sunt principes eius velut cervinon invenientes pascuaet abierunt absque fortitudineante faciem persequentis.
LAM|1|7|ZAIN. Recordata est Ierusalemdierum afflictionis suae et peregrinationis,omnium desiderabilium suorum,quae habuerat a diebus antiquis,cum caderet populus eius in manu hostili,et non esset auxiliator;viderunt eam hosteset deriserunt interitum eius.
LAM|1|8|HETH. Peccatum peccavit Ierusalem,propterea abominabilis facta est;omnes, qui glorificabant eam, spreverunt illam,quia viderunt ignominiam eius:ipsa autem gemensconversa est retrorsum.
LAM|1|9|TETH. Sordes eius in fimbriis eius,nec recordata est finis sui;deposita est vehementer,non habens consolatorem. Vide, Domine, afflictionem meam, quoniam erectus est inimicus! ".
LAM|1|10|IOD. Manum suam misit hostisad omnia desiderabilia eius,quia vidit gentesingressas sanctuarium suum,de quibus praeceperas,ne intrarent in ecclesiam tuam.
LAM|1|11|CAPH. Omnis populus eius gemenset quaerens panem;dederunt pretiosa quaeque pro ciboad refocillandam animam. Vide, Domine, et considera,quoniam facta sum vilis!
LAM|1|12|LAMED. O vos omnes, qui transitis per viam,attendite et videte,si est dolor sicut dolor meus,quem paravit mihi,quo afflixit me Dominusin die irae furoris sui.
LAM|1|13|MEM. De excelso misit ignem,in ossa mea immisit eum;expandit rete pedibus meis,convertit me retrorsum:posuit me desolatam,tota die maerore confectam.
LAM|1|14|NUN. Vigilavit super iniquitates meas,in manu eius convolutae suntet impositae collo meo;debilitavit virtutem meam:dedit me Dominus in manu,de qua non potero surgere.
LAM|1|15|SAMECH. Sprevit omnes fortes meosDominus in medio mei;vocavit adversum me conventum,ut contereret iuvenes meos:torcular calcavit Dominusvirgini filiae Iudae.
LAM|1|16|AIN. Idcirco ego plorans,et oculus meus deducens aquas,quia longe factus est a me consolatorreficiens animam meam;facti sunt filii mei desolati,quoniam invaluit inimicus ".
LAM|1|17|PHE. Expandit Sion manus suas,non est qui consoletur eam;mandavit Dominus adversum Iacobin circuitu eius hostes eius:facta est Ierusalemquasi polluta menstruis inter eos.
LAM|1|18|SADE. " Iustus est Dominus,quia contra os eius rebellis fui.Audite, obsecro, universi populi,et videte dolorem meum:virgines meae et iuvenes meiabierunt in captivitatem.
LAM|1|19|COPH. Vocavi amicos meos,et ipsi deceperunt me;sacerdotes mei et senes meiin urbe consumpti sunt,quia quaesierunt cibum sibi,ut refocillarent animam suam.
LAM|1|20|RES. Vide, Domine, quoniam tribulor;efferbuerunt viscera mea,subversum est cor meum in memetipsa,quoniam valde rebellis fui;foris orbavit me gladiuset domi mors.
LAM|1|21|SIN. Audi, quia ingemisco ego,et non est qui consoletur me;omnes inimici mei audierunt malum meum,laetati sunt quoniam tu fecisti.Adduc diem, quem proclamasti,et fient similes mei.
LAM|1|22|THAU. Ingrediatur omne malum eorum coram te,et fac eis,sicut fecisti mihipropter omnes iniquitates meas;multi enim gemitus mei,et cor meum maerens ".
LAM|2|1|ALEPH. Quomodo obtexit caligine in furore suoDominus filiam Sion!Proiecit de caelo in terramgloriam Israelet non est recordatus scabelli pedum suorumin die furoris sui.
LAM|2|2|BETH. Praecipitavit Dominusnec pepercit omnia pascua Iacob;destruxit in furore suomunitiones filiae Iudae;deiecit in terram, polluitregnum et principes eius.
LAM|2|3|GHIMEL. Confregit in ira furoris suiomne cornu Israel;avertit retrorsum dexteram suama facie inimiciet succendit in Iacob quasi ignem flammaedevorantis in gyro.
LAM|2|4|DALETH. Tetendit arcum suum quasi inimicus,firmavit dexteram suam quasi hostiset occidit omne,quod pulchrum erat visu,in tabernaculo filiae Sion;effudit quasi ignem indignationem suam.
LAM|2|5|HE. Factus est Dominus velut inimicus,deglutivit Israel,deglutivit omnia moenia eius,dissipavit munitiones eiuset multiplicavit in filia Iudaemaerorem et maestitiam.
LAM|2|6|VAU. Et dissipavit quasi hortum saepem suam,demolitus est tabernaculum suum; oblivioni tradidit Dominus in Sion festivitatem et sabbatumet despexit in indignatione furoris suiregem et sacerdotem.
LAM|2|7|ZAIN. Reppulit Dominus altare suum,maledixit sanctuario suo;tradidit in manu inimicimuros domorum eius:vocem dederunt in domo Dominisicut in die sollemni.
LAM|2|8|HETH. Cogitavit Dominus dissiparemurum filiae Sion;tetendit funiculum,non avertit manum suam a perditione;et in luctum redegit antemurale et murum:pariter elanguerunt.
LAM|2|9|TETH. Defixae sunt in terra portae eius;perdidit et contrivit vectes eius.Rex eius et principes eius in gentibus;non est lex,et prophetae eius non inveneruntvisionem a Domino.
LAM|2|10|IOD. Sederunt in terra,conticuerunt senes filiae Sion,consperserunt cinere capita sua,accincti sunt ciliciis;abiecerunt in terram capita suavirgines Ierusalem.
LAM|2|11|CAPH. Defecerunt prae lacrimis oculi mei,efferbuerunt viscera mea;effusum est in terra iecur meumsuper contritione filiae populi mei,cum deficeret parvulus et lactansin plateis oppidi.
LAM|2|12|LAMED. Matribus suis dixerunt: Ubi est triticum et vinum? ",cum deficerent quasi vulneratiin plateis civitatis,cum exhalarent animas suasin sinu matrum suarum.
LAM|2|13|MEM. Cui comparabo te vel cui assimilabo te,filia Ierusalem?Cui exaequabo te et consolabor te, virgo filia Sion?Magna est enim velut mare contritio tua;quis medebitur tui?
LAM|2|14|NUN. Prophetae tui viderunt tibi falsa et stultanec aperiebant iniquitatem tuam,ut converterent sortem tuam;viderunt autem tibi oraculamendacii et seductionis.
LAM|2|15|SAMECH. Plauserunt super te manibusomnes transeuntes per viam;sibilaverunt et moverunt caput suumsuper filiam Ierusalem: Haeccine est urbs, quam vocabant perfectum decorem,gaudium universae terrae? ".
LAM|2|16|PHE. Aperuerunt super te os suumomnes inimici tui;sibilaverunt et fremuerunt dentibuset dixerunt: " Devoravimus;en ista est dies, quam exspectabamus:invenimus, vidimus ".
LAM|2|17|AIN. Fecit Dominus, quae cogitavit;complevit sermonem suum,quem praeceperat a diebus antiquis:destruxit et non pepercit.Et laetificavit super te inimicumet exaltavit cornu hostium tuorum.
LAM|2|18|SADE. Clamet cor tuum ad Dominumsuper muros filiae Sion;deduc quasi torrentem lacrimasper diem et noctem.Non des requiem tibi,neque taceat pupilla oculi tui.
LAM|2|19|COPH. Consurge, lamentare in noctein principio vigiliarum,effunde sicut aquam cor tuumante conspectum Domini;leva ad eum manus tuaspro anima parvulorum tuorum,qui defecerunt in famein capite omnium compitorum.
LAM|2|20|RES. " Vide, Domine, et considera,cui feceris ita;ergone comedent mulieres fructum suum,parvulos diligenter fovendos?Num occidetur in sanctuario Dominisacerdos et propheta?
LAM|2|21|SIN. Iacuerunt in terra forispuer et senex;virgines meae et iuvenes meiceciderunt in gladio:interfecisti in die furoris tui,percussisti nec misertus es.
LAM|2|22|THAU. Vocasti quasi ad diem sollemnem,qui terrerent me de circuitu,et non fuit in die furoris Domini,qui effugeret et relinqueretur:quos fovi et enutrivi,inimicus meus consumpsit eos ".
LAM|3|1|ALEPH. Ego vir videns paupertatem meamin virga indignationis eius.
LAM|3|2|ALEPH. Me minavit et adduxitin tenebras et non in lucem.
LAM|3|3|ALEPH. Tantum in me vertit et convertitmanum suam tota die.
LAM|3|4|BETH. Consumpsit pellem meam et carnem meam,contrivit ossa mea.
LAM|3|5|BETH. Aedificavit in gyro meoet circumdedit me felle et labore.
LAM|3|6|BETH. In tenebrosis collocavit mequasi mortuos sempiternos.
LAM|3|7|GHIMEL. Circumaedificavit adversum me, ut non egrediar,aggravavit compedem meum.
LAM|3|8|GHIMEL. Sed et cum clamavero et rogavero,exclusit orationem meam.
LAM|3|9|GHIMEL. Conclusit vias meas lapidibus quadris,semitas meas subvertit.
LAM|3|10|DALETH. Ursus insidians factus est mihi,leo in absconditis.
LAM|3|11|DALETH. Semitas meas subvertit et confregit me,posuit me desolatam.
LAM|3|12|DALETH. Tetendit arcum suum et posuit mequasi signum ad sagittam.
LAM|3|13|HE. Misit in renibus meisfilias pharetrae suae.
LAM|3|14|HE. Factus sum in derisum omni populo meo,canticum eorum tota die.
LAM|3|15|HE. Replevit me amaritudinibus,inebriavit me absinthio.
LAM|3|16|VAU. Et fregit in glarea dentes meos,depressit me cinere.
LAM|3|17|VAU. Et repulsa est a pace anima mea,oblitus sum bonorum.
LAM|3|18|VAU. Et dixi: " Periit splendor meus et spes mea a Domino ".
LAM|3|19|ZAIN. Recordare paupertatis et peregrinationis meae,absinthii et fellis.
LAM|3|20|ZAIN. Memoria memor estet tabescit in me anima mea.
LAM|3|21|ZAIN. Haec recolam in corde meo,ideo sperabo.
LAM|3|22|HETH. Misericordiae Domini, quia non sumus consumpti,quia non defecerunt miserationes eius.
LAM|3|23|HETH. Novae sunt omni mane,magna est fides tua.
LAM|3|24|HETH. " Pars mea Dominus, dixit anima mea;propterea exspectabo eum ".
LAM|3|25|TETH. Bonus est Dominus sperantibus in eum,animae quaerenti illum.
LAM|3|26|TETH. Bonum est praestolari cum silentiosalutare Domini.
LAM|3|27|TETH. Bonum est viro, cum portaveritiugum ab adulescentia sua.
LAM|3|28|IOD. Sedebit solitarius et tacebit,cum istud imponitur ei.
LAM|3|29|IOD. Ponet in pulvere os suum,si forte sit spes.
LAM|3|30|IOD. Dabit percutienti se maxillam,saturabitur opprobriis.
LAM|3|31|CAPH. Quia non repellet in sempiternumDominus.
LAM|3|32|CAPH. Quia si afflixit, et miserebitursecundum multitudinem misericordiarum suarum.
LAM|3|33|CAPH. Non enim humiliat ex corde suoet affligit filios hominum.
LAM|3|34|LAMED. Conterere sub pedibus suisomnes vinctos terrae.
LAM|3|35|LAMED. Declinare iudicium viriin conspectu vultus Altissimi.
LAM|3|36|LAMED. Pervertere hominem in iudicio suo,num Dominus haec ignorat?
LAM|3|37|MEM. Quis est iste, qui dixit, et factum est?Dominus non iussit?
LAM|3|38|MEM. Ex ore Altissimi nonne egrediunturet mala et bona?
LAM|3|39|MEM. Quid murmurabit homo vivens,vir pro peccatis suis?
LAM|3|40|NUN. " Scrutemur vias nostras et quaeramuset revertamur ad Dominum.
LAM|3|41|NUN. Levemus corda nostra cum manibusad Dominum in caelos.
LAM|3|42|NUN. Nos inique egimus et rebelles fuimus;idcirco tu inexorabilis fuisti.
LAM|3|43|SAMECH. Operuisti in furore et percussisti nos;occidisti nec pepercisti.
LAM|3|44|SAMECH. Opposuisti nubem tibi,ne transeat oratio.
LAM|3|45|SAMECH. In eradicationem et abiectionem posuisti nosin medio populorum.
LAM|3|46|PHE. Aperuerunt super nos os suumomnes inimici nostri.
LAM|3|47|PHE. Formido et fovea facta est nobis,vastatio et contritio ".
LAM|3|48|PHE. Rivos aquarum deducit oculus meusin contritione filiae populi mei.
LAM|3|49|AIN. Oculus meus lacrimas effundit nec tacet,eo quod non sit requies.
LAM|3|50|AIN. Donec respiciat et videatDominus de caelis.
LAM|3|51|AIN. Oculus meus affligit animam meamprae cunctis filiabus urbis meae.
LAM|3|52|SADE. Venatione venati sunt me quasi aveminimici mei gratis.
LAM|3|53|SADE. Perdiderunt in lacu vitam meamet iecerunt lapides super me.
LAM|3|54|SADE. Inundaverunt aquae super caput meum,dixi: " Perii ".
LAM|3|55|COPH. Invocavi nomen tuum, Domine,de profunditate lacus.
LAM|3|56|COPH. Vocem meam audisti: " Ne avertasaurem tuam a singultu meo et clamoribus ".
LAM|3|57|COPH. Appropinquasti in die, quando invocavi te,dixisti: " Ne timeas ".
LAM|3|58|RES. Iudicasti, Domine, causam animae meae,redemisti vitam meam.
LAM|3|59|RES. Vidisti, Domine, afflictionem meam;iudica iudicium meum.
LAM|3|60|RES. Vidisti omnem furorem eorum, universas cogitationes eorum adversum me.
LAM|3|61|SIN. Audisti opprobrium eorum, Domine,omnes cogitationes eorum adversum me.
LAM|3|62|SIN. Labia insurgentium mihi et meditationes eorumadversum me tota die.
LAM|3|63|SIN. Sessionem eorum et resurrectionem eorum vide;ego sum psalmus eorum.
LAM|3|64|THAU. Reddes eis vicem, Domine,iuxta opera manuum suarum.
LAM|3|65|THAU. Dabis eis duritiam cordis,exsecrationem tuam.
LAM|3|66|THAU. Persequeris in furore et conteres eossub caelis tuis, Domine.
LAM|4|1|ALEPH. Quomodo obscuratum est aurum,mutatum est obryzum optimum!Dispersi sunt lapides sanctiin capite omnium platearum.
LAM|4|2|BETH. Filii Sion inclitiet ponderati auro primo,quomodo reputati sunt in vasa testea,opus manuum figuli!
LAM|4|3|GHIMEL. Sed et thoes nudaverunt mammam,lactaverunt catulos suos;filia populi mei crudelisquasi struthio in deserto.
LAM|4|4|DALETH. Adhaesit lingua lactantisad palatum eius in siti;parvuli petierunt panem,et non erat qui frangeret eis.
LAM|4|5|HE. Qui vescebantur voluptuose,interierunt in viis;qui nutriebantur in coccinis,amplexati sunt stercora.
LAM|4|6|VAU. Et maior effecta est iniquitas filiae populi meipeccato Sodomae,quae subversa est in momento,et non laborabant in ea manus.
LAM|4|7|ZAIN. Candidiores nazaraei eius nive,nitidiores lacte,rubicundiores in corpore coralliis,sapphirus aspectus eorum.
LAM|4|8|HETH. Denigrata est super carbones facies eorum,et non sunt cogniti in plateis:adhaesit cutis eorum ossibus,aruit et facta est quasi lignum.
LAM|4|9|TETH. Melius fuit occisis gladioquam interfectis fame,quoniam isti extabuerunt consumptia sterilitate terrae.
LAM|4|10|IOD. Manus mulierum misericordiumcoxerunt filios suos:facti sunt cibus earumin contritione filiae populi mei.
LAM|4|11|CAPH. Complevit Dominus furorem suum,effudit iram indignationis suae;et succendit ignem in Sion,qui devoravit fundamenta eius.
LAM|4|12|LAMED. Non crediderunt reges terraeet universi habitatores orbis,quoniam ingrederetur hostis et inimicusper portas Ierusalem.
LAM|4|13|MEM. Propter peccata prophetarum eiuset iniquitates sacerdotum eius,qui effuderunt in medio eiussanguinem iustorum.
LAM|4|14|NUN. Erraverunt caeci in plateis,polluti sunt in sanguine,ita ut nemo posset attingerelacinias eorum.
LAM|4|15|SAMECH. " Recedite! Pollutus est ", clamaverunt eis; Recedite, abite, nolite tangere! ".Cum fugerent et errarent, dixerunt inter gentes: Non addent ultra ut incolant ".
LAM|4|16|PHE. Facies Domini dispersit eos,non addet ut respiciat eos;facies sacerdotum non respexeruntneque senum miserti sunt.
LAM|4|17|AIN. Adhuc deficiunt oculi nostriad auxilium nostrum vanum?In specula nostra respeximusad gentem, quae salvare non potest.
LAM|4|18|SADE. Insidiati sunt vestigiis nostris,ne iremus per plateas nostras. Appropinquavit finis noster, completi sunt dies nostri,quia venit finis noster ".
LAM|4|19|COPH. Velociores fuerunt persecutores nostriaquilis caeli;super montes persecuti sunt nos,in deserto insidiati sunt nobis.
LAM|4|20|RES. Spiritus oris nostri, unctus Domini,captus est in foveis eorum,de quo dicebamus: " Sub umbra suavivemus in gentibus ".
LAM|4|21|SIN. Gaude et laetare, filia Edom,quae habitas in terra Us;ad te quoque perveniet calix,inebriaberis atque nudaberis.
LAM|4|22|THAU. Completa est iniquitas tua, filia Sion,non addet ultra ut transmigret te;visitavit iniquitatem tuam, filia Edom,discooperuit peccata tua.
LAM|5|1|Recordare, Domine, quid acci derit nobis;intuere et respice opprobrium nostrum.
LAM|5|2|Hereditas nostra versa est ad alienos,domus nostrae ad extraneos.
LAM|5|3|Pupilli facti sumus absque patre,matres nostrae quasi viduae.
LAM|5|4|Aquam nostram pecunia bibimus,ligna nostra pretio comparamus.
LAM|5|5|Iugum in cervicibus nostris minamur;lassis non datur requies.
LAM|5|6|Aegyptiis dedimus manum et Assyriis,ut saturaremur pane.
LAM|5|7|Patres nostri peccaverunt et non sunt,et nos iniquitates eorum portamus.
LAM|5|8|Servi dominantur nostri;non est qui redimat de manu eorum.
LAM|5|9|Vitae nostrae periculo afferimus panem nobisa facie gladii in deserto.
LAM|5|10|Pellis nostra quasi clibanus exusta estpropter aestum famis.
LAM|5|11|Mulieres in Sion humiliaveruntet virgines in civitatibus Iudae.
LAM|5|12|Principes manu eorum suspensi sunt;facies senum honorem non habuerunt.
LAM|5|13|Adulescentes molam portaverunt,et pueri sub lignis corruerunt.
LAM|5|14|Senes deficiunt de portis,iuvenes de choro psallentium.
LAM|5|15|Defecit gaudium cordis nostri;versus est in luctum chorus noster.
LAM|5|16|Cecidit corona capitis nostri;vae nobis, quia peccavimus!
LAM|5|17|Propterea maestum factum est cor nostrum,ideo contenebrati sunt oculi nostri,
LAM|5|18|propter montem Sion, quia desolatus est:vulpes ambulant in eo.
LAM|5|19|Tu autem, Domine, in aeternum permanebis,solium tuum in generationem et generationem.
LAM|5|20|Quare in perpetuum oblivisceris nostri,derelinques nos in longitudinem dierum?
LAM|5|21|Converte nos, Domine, ad te, et convertemur;innova dies nostros sicut a principio.
LAM|5|22|Ergone proiciens reppulisti nos,iratus es contra nos vehementer?
EZEK|1|1|Et factum est in tricesimo anno, in quarto mense, in quinta men sis, cum essem in medio captivorum iuxta fluvium Chobar, aperti sunt caeli, et vidi visiones Dei.
EZEK|1|2|In quinta mensis, ipse est annus quintus transmigrationis regis Ioachin,
EZEK|1|3|factum est verbum Domini ad Ezechielem filium Buzi, sacerdotem, in terra Chaldaeorum secus flumen Chobar, et facta est super eum ibi manus Domini.
EZEK|1|4|Et vidi: et ecce ventus turbinis veniebat ab aquilone et nubes magna et ignis conglobatus, et splendor in circuitu eius, et de medio eius quasi species electri, id est de medio ignis;
EZEK|1|5|et ex medio eius similitudo quattuor animalium, et hic aspectus eorum: similitudo hominis erat eis.
EZEK|1|6|Quattuor facies uni et quattuor pennae uni;
EZEK|1|7|pedes eorum pedes recti, et planta pedis eorum quasi planta pedis vituli, et scintillabant quasi aspectus aeris candentis.
EZEK|1|8|Et manus hominis erant sub pennis eorum in quattuor partibus. Facies autem et pennae illorum quattuor:
EZEK|1|9|iunctae erant pennae eorum altera ad alteram; non revertebantur, cum incederent, sed unumquodque ante faciem suam gradiebatur.
EZEK|1|10|Similitudo autem vultus eorum: facies hominis et facies leonis a dextris ipsorum quattuor, facies autem bovis a sinistris ipsorum quattuor et facies aquilae ipsorum quattuor.
EZEK|1|11|Et pennae eorum extentae desuper; duae pennae singulorum iungebantur, et duae tegebant corpora eorum.
EZEK|1|12|Et unumquodque coram facie sua ambulabat: ubi erat impetus spiritus, illuc gradiebantur nec revertebantur, cum ambularent.
EZEK|1|13|Et in medio animalium, aspectus quasi carbonum ignis ardentium, quasi aspectus lampadarum discurrentium in medio animalium; et splendor erat ignis, et de igne fulgur egrediens.
EZEK|1|14|Et animalia ibant et revertebantur in similitudinem fulguris coruscantis.
EZEK|1|15|Cumque aspicerem animalia, apparuit rota una super terram iuxta singula animalia.
EZEK|1|16|Et aspectus rotarum et opus earum quasi species chrysolithi, et una similitudo ipsarum quattuor; et aspectus earum et opera, quasi sit rota in medio rotae.
EZEK|1|17|Per quattuor partes earum euntes ibant et non revertebantur, cum ambularent.
EZEK|1|18|Canthis autem earum erat altitudo et horribilis aspectus; et canthi earum erant oculis pleni in circuitu ipsarum quattuor.
EZEK|1|19|Cumque ambularent animalia, ambulabant pariter et rotae iuxta ea; et cum elevarentur animalia de terra, elevabantur simul et rotae.
EZEK|1|20|Quocumque impellebat spiritus ut irent, ibant, et rotae pariter levabantur sequentes eum; spiritus enim animalium erat in rotis.
EZEK|1|21|Cum euntibus ibant et cum stantibus stabant; et cum elevatis a terra pariter elevabantur, et rotae sequentes ea, quia spiritus animalium erat in rotis.
EZEK|1|22|Et similitudo super capita animalium firmamenti quasi aspectus crystalli horribilis et extenti super capita eorum desuper.
EZEK|1|23|Sub firmamento autem pennae eorum rectae altera ad alteram; unumquodque duabus alis velabat corpus suum.
EZEK|1|24|Et audiebam sonum alarum quasi sonum aquarum multarum, quasi sonum Omnipotentis: cum ambularent, erat strepitus vehemens ut sonus castrorum; cumque starent, demittebantur pennae eorum.
EZEK|1|25|Nam cum fieret vox supra firmamentum, quod erat super caput eorum, stabant et submittebant alas suas.
EZEK|1|26|Et super firmamentum, quod erat imminens capiti eorum, quasi aspectus lapidis sapphiri similitudo throni; et super similitudinem throni similitudo quasi aspectus hominis desuper.
EZEK|1|27|Et vidi quasi speciem electri, velut aspectum ignis per circuitum ab aspectu lumborum eius et desuper; et ab aspectu lumborum eius usque deorsum vidi quasi speciem ignis splendentis in circuitu.
EZEK|1|28|Velut aspectus arcus, cum fuerit in nube in die pluviae: sic erat aspectus splendoris per gyrum. Haec visio similitudinis gloriae Domini. Et vidi et cecidi in faciem meam et audivi vocem loquentis.
EZEK|2|1|Et dixit ad me: " Fili hominis, sta super pedes tuos, et loquar tecum ".
EZEK|2|2|Et ingressus est in me spiritus, postquam locutus est mihi et statuit me supra pedes meos, et audivi loquentem ad me
EZEK|2|3|et dicentem: " Fili hominis, mitto ego te ad filios Israel, ad gentes apostatrices, quae recesserunt a me; ipsi et patres eorum praevaricati sunt in me usque ad diem hanc.
EZEK|2|4|Et filii dura facie et obstinato corde sunt, ad quos ego mitto te; et dices ad eos: Haec dicit Dominus Deus.
EZEK|2|5|Ipsi sive audiant, sive contemnant - quoniam domus exasperans est - sciant tamen quia propheta fuerit in medio eorum.
EZEK|2|6|Tu ergo, fili hominis, ne timeas eos neque sermones eorum metuas, etsi cardui et spinae te circumdant, et cum scorpionibus habitas. Verba eorum ne timeas et vultus eorum ne formides, quia domus exasperans est.
EZEK|2|7|Loqueris ergo verba mea ad eos, sive audiant, sive contemnant, quoniam exasperantes sunt.
EZEK|2|8|Tu autem, fili hominis, audi, quaecumque loquor ad te, et noli esse exasperans, sicut domus exasperatrix est; aperi os tuum et comede, quaecumque ego do tibi ".
EZEK|2|9|Et vidi: et ecce manus missa ad me, in qua erat involutus liber; et expandit illum coram me, qui erat scriptus intus et foris, et scriptae erant in eo lamentationes et gemitus et vae.
EZEK|3|1|Et dixit ad me: " Fili hominis, quodcumque inveneris, comede; comede volumen istud et vadens loquere ad filios Israel ".
EZEK|3|2|Et aperui os meum, et cibavit me volumine illo
EZEK|3|3|et dixit ad me: " Fili hominis, venter tuus comedet, et viscera tua complebuntur volumine isto, quod ego do tibi ". Et comedi illud, et factum est in ore meo sicut mel dulce.
EZEK|3|4|Et dixit ad me: " Fili hominis, vade ad domum Israel et loqueris verba mea ad eos.
EZEK|3|5|Non enim ad populum profundi sermonis et ignotae linguae tu mitteris, ad domum Israel;
EZEK|3|6|neque ad populos multos profundi sermonis et ignotae linguae, quorum non possis audire sermones; et si ad illos mittereris, ipsi audirent te.
EZEK|3|7|Domus autem Israel nolunt audire te, quia nolunt audire me; omnis quippe domus Israel dura fronte est et obstinato corde.
EZEK|3|8|Ecce dedi faciem tuam valentiorem faciebus eorum et frontem tuam duriorem frontibus eorum;
EZEK|3|9|ut adamantem et duriorem silice dedi faciem tuam: ne timeas eos neque metuas a facie eorum, quia domus exasperans est ".
EZEK|3|10|Et dixit ad me: " Fili hominis, omnes sermones meos, quos loquor ad te, assume in corde tuo et auribus tuis audi.
EZEK|3|11|Et vade, ingredere ad transmigrationem, ad filios populi tui, et loqueris ad eos et dices eis: Haec dicit Dominus Deus; sive audiant, sive contemnant ".
EZEK|3|12|Et assumpsit me spiritus, et audivi post me vocem commotionis magnae, cum elevaretur gloria Domini de loco suo;
EZEK|3|13|et vocem alarum animalium percutientium alteram ad alteram et vocem rotarum sequentium animalia et vocem commotionis magnae.
EZEK|3|14|Spiritus quoque levavit me et assumpsit me; et abii amarus in indignatione spiritus mei: manus enim Domini erat super me gravis.
EZEK|3|15|Et veni ad transmigrationem, ad Telabib, ad eos, qui habitabant iuxta flumen Chobar; et sedi, ubi illi sedebant, et mansi ibi septem diebus obstupefactus in medio eorum.
EZEK|3|16|Cum autem pertransissent septem dies, factum est verbum Domini ad me dicens:
EZEK|3|17|" Fili hominis, speculatorem dedi te domui Israel; et audies de ore meo verbum et commonebis eos ex me.
EZEK|3|18|Si, dicente me ad impium: Morte morieris, non commonueris eum neque locutus fueris ei, ut avertatur a via sua impia et vivat, ipse impius in iniquitate sua morietur, sanguinem autem eius de manu tua requiram.
EZEK|3|19|Si autem tu commonueris impium, et ille non fuerit conversus ab impietate sua et a via sua impia, ipse quidem in iniquitate sua morietur, tu autem animam tuam liberasti.
EZEK|3|20|Sed et si conversus iustus a iustitia sua, fecerit iniquitatem, ponam offendiculum coram eo; ipse morietur, quia non commonuisti eum: in peccato suo morietur, et non erunt in memoria iustitiae eius, quas fecit; sanguinem vero eius de manu tua requiram.
EZEK|3|21|Si autem tu commonueris iustum, ut non peccet iustus, et ille non peccaverit, vivens vivet, quia commonuisti eum et tu animam tuam liberasti.
EZEK|3|22|Et facta est super me manus Domini, et dixit ad me: " Surgens egredere in campum, et ibi loquar tecum ".
EZEK|3|23|Et surgens egressus sum in campum, et ecce ibi gloria Domini stabat quasi gloria, quam vidi iuxta fluvium Chobar, et cecidi in faciem meam.
EZEK|3|24|Et ingressus est in me spiritus et statuit me super pedes meos et locutus est mihi et dixit ad me: " Ingredere et includere in medio domus tuae.
EZEK|3|25|Et tu, fili hominis, ecce data sunt super te vincula, et ligabunt te in eis, et non egredieris in medio eorum;
EZEK|3|26|et linguam tuam adhaerere faciam palato tuo, et eris mutus nec quasi vir obiurgans, quia domus exasperans est.
EZEK|3|27|Cum autem locutus fuero tibi, aperiam os tuum, et dices ad eos: Haec dicit Dominus Deus. Qui audit, audiat; et, qui contemnit, contemnat, quia domus exasperans est ".
EZEK|4|1|" Et tu, fili hominis, sume tibi laterem et pones eum coram te et describes in eo civitatem Ierusalem.
EZEK|4|2|Et ordinabis adversus eam obsidionem et aedificabis munitiones et comportabis aggerem et dabis contra eam castra et pones arietes in gyro.
EZEK|4|3|Et tu sume tibi sartaginem ferream et pones eam in murum ferreum inter te et inter civitatem; et obfirmabis faciem tuam ad eam, et erit in obsidionem, et circumdabis eam: signum est domui Israel.
EZEK|4|4|Et tu recumbes super latus tuum sinistrum et pones iniquitates domus Israel super eo; numero dierum, quibus recumbes super illud, assumes iniquitatem eorum.
EZEK|4|5|Ego autem dedi tibi annos iniquitatis eorum numero dierum trecentos et nonaginta dies, et portabis iniquitatem domus Israel.
EZEK|4|6|Et cum compleveris haec, recumbes super latus tuum dextrum secundo et assumes iniquitatem domus Iudae quadraginta diebus; diem pro anno, diem, inquam, pro anno dedi tibi.
EZEK|4|7|Et ad obsidionem Ierusalem convertes faciem tuam, et brachium tuum erit exsertum, et prophetabis adversus eam.
EZEK|4|8|Ecce circumdedi te vinculis, et non te convertes a latere tuo in latus aliud, donec compleas dies obsidionis tuae.
EZEK|4|9|Et tu sume tibi frumentum et hordeum et fabam et lentem et milium et far et mittes ea in vas unum et facies tibi panes numero dierum, quibus recumbes super latus tuum: trecentis et nonaginta diebus comedes illud.
EZEK|4|10|Cibus autem tuus, quo vesceris, erit in pondere viginti stateres in die; a tempore usque ad tempus comedes illud.
EZEK|4|11|Et aquam in mensura bibes, sextam partem hin; a tempore usque ad tempus bibes illud.
EZEK|4|12|Et quasi subcinericium hordeaceum comedes illud; et stercore, quod egreditur de homine, coques illud in oculis eorum".
EZEK|4|13|Et dixit Dominus: " Sic comedent filii Israel panem suum pollutum inter gentes, ad quas eiciam eos ".
EZEK|4|14|Et dixi: " Heu, Domine Deus, ecce anima mea non est polluta, et morticinum et laceratum a bestiis non comedi ab infantia mea usque nunc, et non est ingressa in os meum caro immunda ".
EZEK|4|15|Et dixit ad me: " Ecce dedi tibi fimum boum pro stercoribus humanis, et facies panem tuum in eo ".
EZEK|4|16|Et dixit ad me: " Fili hominis, ecce ego conteram baculum panis in Ierusalem, et comedent panem in pondere et in sollicitudine et aquam in mensura et in desolatione bibent,
EZEK|4|17|ut, deficientibus pane et aqua, desoletur unusquisque cum fratre suo, et contabescant in iniquitatibus suis.
EZEK|5|1|Et tu, fili hominis, sume tibi gladium acutum radentem pilos et assumes eum et duces per caput tuum et per barbam tuam et assumes tibi stateram ponderis et divides eos.
EZEK|5|2|Tertiam partem igne combures in medio civitatis, post completionem dierum obsidionis; et assumens tertiam partem, concides gladio in circuitu eius; tertiam vero aliam disperges in ventum, et gladium nudabo post eos.
EZEK|5|3|Et sumes inde parvum numerum et ligabis eos in summitate pallii tui;
EZEK|5|4|et ex eis rursum tolles et proicies eos in medio ignis et combures eos igne; ex eo egredietur ignis. Et dices ad omnem domum Israel:
EZEK|5|5|Haec dicit Dominus Deus: Ista est Ierusalem! In medio gentium posui eam et in circuitu eius terras.
EZEK|5|6|Et contempsit iudicia mea, ut plus esset impia quam gentes, et praecepta mea ultra quam terrae, quae in circuitu eius sunt: iudicia enim mea proiecerunt et in praeceptis meis non ambulaverunt.
EZEK|5|7|Idcirco haec dicit Dominus Deus: Quia tumultuati estis magis quam gentes, quae in circuitu vestro sunt, et in praeceptis meis non ambulastis et iudicia mea non fecistis et iuxta iudicia gentium, quae in circuitu vestro sunt, non estis operati,
EZEK|5|8|ideo haec dicit Dominus Deus: Ecce ego ad te et ipse ego faciam in medio tui iudicia in oculis gentium
EZEK|5|9|et faciam in te, quae non feci et quibus similia ultra non faciam, propter omnes abominationes tuas.
EZEK|5|10|Ideo patres comedent filios in medio tui, et filii comedent patres suos, et faciam in te iudicia et ventilabo universas reliquias tuas in omnem ventum.
EZEK|5|11|Idcirco vivo ego, dicit Dominus Deus, vere pro eo quod sanctum meum violasti in omnibus offensionibus tuis et in omnibus abominationibus tuis, ego quoque radam, et non parcet oculus meus, et non miserebor.
EZEK|5|12|Tertia tui pars peste morietur et fame consumetur in medio tui, et tertia tui pars in gladio cadet in circuitu tuo, tertiam vero partem tuam in omnem ventum dispergam et gladium evaginabo post eos.
EZEK|5|13|Et complebo furorem meum et requiescere faciam indignationem meam in eis et consolabor; et scient quia ego Dominus locutus sum in zelo meo, cum implevero indignationem meam in eis.
EZEK|5|14|Et dabo te in desertum et in opprobrium in gentibus, quae in circuitu tuo sunt, in conspectu omnis praetereuntis;
EZEK|5|15|et eris opprobrium et blasphemia, exemplum et stupor in gentibus, quae in circuitu tuo sunt, cum fecero in te iudicia in furore et in indignatione et in castigationibus irae.
EZEK|5|16|Ego Dominus locutus sum. Quando misero sagittas famis pessimas in vos, quae erunt mortiferae, et quas mittam, ut destruam vos, et famem congregabo super vos et conteram vobis baculum panis;
EZEK|5|17|et immittam in vos famem et bestias pessimas, et absque liberis facient te, et pestilentia et sanguis transibunt per te, et gladium inducam super te. Ego Dominus locutus sum ".
EZEK|6|1|Et factus est sermo Domini ad me dicens:
EZEK|6|2|" Fili hominis, pone faciem tuam ad montes Israel et prophetabis ad eos
EZEK|6|3|et dices: Montes Israel, audite verbum Domini Dei. Haec dicit Dominus Deus montibus et collibus, voraginibus et vallibus: Ecce ego inducam super vos gladium et destruam excelsa vestra;
EZEK|6|4|et demoliar aras vestras, et confringentur delubra vestra, et deiciam interfectos vestros ante idola vestra.
EZEK|6|5|Et dabo cadavera filiorum Israel ante faciem simulacrorum vestrorum et dispergam ossa vestra circum aras vestras;
EZEK|6|6|in omnibus habitationibus vestris urbes desertae erunt, et excelsa demolientur, ut dissipentur et intereant arae vestrae, et confringantur et cessent idola vestra, et conterantur delubra vestra, et deleantur opera vestra.
EZEK|6|7|Et cadet interfectus in medio vestri, et scietis quia ego Dominus.
EZEK|6|8|Et relinquam in vobis eos, qui fugerint gladium in gentibus, cum dispersero vos in terris;
EZEK|6|9|et recordabuntur mei liberati vestri in gentibus, ad quas captivi ducti sunt, quia contrivi cor eorum fornicans et recedens a me, et oculos eorum fornicantes post idola sua; et displicebunt sibimet super malis, quae fecerunt in universis abominationibus suis,
EZEK|6|10|et scient quia ego Dominus non frustra locutus sum, ut facerem eis malum hoc.
EZEK|6|11|Haec dicit Dominus Deus: Plaude manu tua et percute pede tuo et dic: Heu ad omnes abominationes malas domus Israel, quia gladio, fame et peste ruituri sunt!
EZEK|6|12|Qui longe est, peste morietur; qui autem prope, gladio corruet; et, qui relictus fuerit et obsessus, fame morietur, et complebo indignationem meam in eis.
EZEK|6|13|Et scietis quia ego Dominus, cum fuerint interfecti eorum in medio idolorum suorum, in circuitu ararum suarum, in omni colle excelso, in cunctis summitatibus montium et subtus omne lignum nemorosum et subtus universam quercum frondosam, locum ubi obtulerunt tura redolentia universis idolis suis.
EZEK|6|14|Et extendam manum meam super eos et faciam terram desolatam et destitutam a deserto usque Rebla in omnibus habitationibus eorum, et scient quia ego Dominus ".
EZEK|7|1|Et factus est sermo Domini ad me dicens:
EZEK|7|2|" Et tu, fili hominis, loquere. Haec dicit Dominus Deus terrae Israel: Finis venit, finis super quattuor plagas terrae;
EZEK|7|3|nunc finis super te, et immittam furorem meum in te et iudicabo te iuxta vias tuas et ponam super te omnes abominationes tuas.
EZEK|7|4|Et non parcet oculus meus super te, et non miserebor, sed vias tuas ponam super te, et abominationes tuae in medio tui erunt, et scietis quia ego Dominus.
EZEK|7|5|Haec dicit Dominus Deus: Afflictio super afflictionem ecce venit.
EZEK|7|6|Finis venit, venit finis; evigilavit adversum te, ecce venit.
EZEK|7|7|Venit contractio super te, qui habitas in terra; venit tempus, prope est dies turbationis et non iubilationis in montibus.
EZEK|7|8|Nunc de propinquo effundam iram meam super te et complebo furorem meum in te et iudicabo te iuxta vias tuas et imponam tibi omnia scelera tua;
EZEK|7|9|et non parcet oculus meus, nec miserebor, sed vias tuas imponam tibi, et abominationes tuae in medio tui erunt, et scietis quia ego sum Dominus percutiens.
EZEK|7|10|Ecce dies, ecce venit; egressa est contractio, floruit iniustitia, germinavit superbia;
EZEK|7|11|violentia surrexit, ut esset virga impietatis: non ex eis et non ex pompa eorum neque ex sonitu eorum; et non erit requies in eis.
EZEK|7|12|Venit tempus, appropinquavit dies: qui emit, non laetetur; et, qui vendit, non lugeat, quia ira super omnem pompam eius.
EZEK|7|13|Quia, qui vendit, ad id quod vendidit non revertetur, cum adhuc sit in viventibus vita eorum. Visio enim ad omnem pompam eius non regredietur, et unusquisque in iniquitate sua vitam suam non confortabit.
EZEK|7|14|Canite tuba, praeparentur omnia, sed non est qui vadat ad proelium; ira enim mea super universam pompam eius.
EZEK|7|15|Gladius foris, pestis et fames intrinsecus. Qui in agro est, gladio morietur; et, qui in civitate, fame et pestilentia devorabuntur.
EZEK|7|16|Et salvabuntur, qui fugerint ex eis, et erunt in montibus quasi columbae convallium omnes gementes, unusquisque in iniquitate sua.
EZEK|7|17|Omnes manus dissolventur, et omnia genua fluent aquis.
EZEK|7|18|Et accingent se ciliciis, et operiet eos formido; et in omni facie confusio, et in universis capitibus eorum calvitium.
EZEK|7|19|Argentum suum foras proicient, et aurum eorum in immunditiam erit; argentum eorum et aurum eorum non valebit liberare eos in die furoris Domini; animam suam non saturabunt, et ventres eorum non implebuntur, quia scandalum iniquitatis eorum factum est,
EZEK|7|20|et ornamentum monilium suorum in superbiam posuerunt et imagines abominationum suarum et simulacrorum fecerunt ex eo; propter hoc dedi eis illud in immunditiam.
EZEK|7|21|Et dabo illud in manus alienorum ad diripiendum et impiis terrae in praedam, et contaminabunt illud.
EZEK|7|22|Et avertam faciem meam ab eis, et violabunt thesaurum meum absconditum; et introibunt in illud praedones et contaminabunt illud
EZEK|7|23|et facient ex illo catenas; quoniam terra plena est iudicio sanguinum, et civitas plena iniquitate.
EZEK|7|24|Et adducam pessimos de gentibus, et possidebunt domos eorum; et quiescere faciam superbiam potentium, et possidebunt sanctuaria eorum.
EZEK|7|25|Angustia superveniente, requirent pacem, et non erit.
EZEK|7|26|Calamitas super calamitatem veniet, et auditus super auditum; et quaerent visionem de propheta, et lex peribit a sacerdote, et consilium a senioribus.
EZEK|7|27|Rex lugebit, et princeps induetur horrore, et manus populi terrae conturbabuntur. Secundum viam eorum faciam eis et secundum iudicia eorum iudicabo eos, et scient quia ego Dominus ".
EZEK|8|1|Et factum est in anno sexto, in sexto mense, in quinta mensis, ego sedebam in domo mea, et senes Iudae sedebant coram me, et cecidit super me ibi manus Domini Dei,
EZEK|8|2|et vidi: et ecce similitudo quasi aspectus viri, ab aspectu lumborum eius et deorsum ignis, et a lumbis eius et sursum quasi aspectus splendoris ut visio electri.
EZEK|8|3|Emisit similitudinem manus et apprehendit me in cincinno capitis mei; et elevavit me spiritus inter terram et caelum et adduxit in Ierusalem, in visionibus Dei, iuxta ostium interius, quod respiciebat aquilonem, ubi erat statutum idolum zeli ad provocandam aemulationem.
EZEK|8|4|Et ecce ibi gloria Dei Israel secundum visionem, quam videram in campo;
EZEK|8|5|et dixit ad me: " Fili hominis, leva oculos tuos ad viam aquilonis ". Et levavi oculos meos ad viam aquilonis, et ecce ab aquilone portae altaris hoc idolum zeli in introitu.
EZEK|8|6|Et dixit ad me: " Fili hominis, putasne vides tu, quid isti faciunt, abominationes magnas, quas domus Israel facit hic, ut procul recedam a sanctuario meo? Et adhuc conversus videbis abominationes maiores ".
EZEK|8|7|Et duxit me ad ostium atrii, et vidi: et ecce foramen unum in pariete.
EZEK|8|8|Et dixit ad me: "Fili hominis, fode parietem"; et cum perfodissem parietem, apparuit ostium unum.
EZEK|8|9|Et dixit ad me: " Ingredere et vide abominationes pessimas, quas isti faciunt hic ".
EZEK|8|10|Et ingressus vidi: et ecce omnis similitudo reptilium et animalium abominatio et universa idola domus Israel depicta erant in pariete in circuitu per totum;
EZEK|8|11|et septuaginta viri de senioribus domus Israel, et Iezonias filius Saphan stabat in medio eorum stantium ante picturas, et unusquisque habebat turibulum in manu sua, et vapor nebulae de ture consurgebat.
EZEK|8|12|Et dixit ad me: " Certe vides, fili hominis, quae seniores domus Israel faciunt in tenebris, unusquisque in cubiculo simulacri sui; dicunt enim: Non videt Dominus nos, dereliquit Dominus terram"".
EZEK|8|13|Et dixit ad me: " Adhuc videbis abominationes maiores, quas isti faciunt ".
EZEK|8|14|Et duxit me ad ostium portae domus Domini, quod respiciebat ad aquilonem, et ecce ibi mulieres sedebant plangentes Thammuz.
EZEK|8|15|Et dixit ad me: "Certe vidisti, fili hominis; adhuc videbis abominationes maiores his ".
EZEK|8|16|Et introduxit me in atrium domus Domini interius, et ecce in ostio templi Domini, inter vestibulum et altare, quasi viginti quinque viri dorsa habentes contra templum Domini et facies ad orientem, et adorabant ad ortum solis.
EZEK|8|17|Et dixit ad me: " Certe vidisti, fili hominis; numquid parum est hoc domui Iudae, ut facerent abominationes istas, quas fecerunt hic, quia replentes terram iniquitate iterum irritaverunt me et ecce applicant ramum ad nares suas.
EZEK|8|18|Ergo et ego faciam in furore: non parcet oculus meus, nec miserebor et, cum clamaverint ad aures meas voce magna, non exaudiam eos ".
EZEK|9|1|Et clamavit in auribus meis voce magna dicens: " Appro pinquaverunt visitationes urbis, et unusquisque vas interfectionis habet in manu sua ".
EZEK|9|2|Et ecce sex viri veniebant de via portae superioris, quae respicit ad aquilonem, et uniuscuiusque vas interitus in manu eius; vir quoque unus in medio eorum vestitus lineis, et atramentarium scriptoris ad renes eius; et ingressi sunt et steterunt iuxta altare aereum.
EZEK|9|3|Et gloria Dei Israel elevata est de cherub, super quem erat, ad limen domus; et vocavit virum, qui indutus erat lineis et atramentarium scriptoris habebat in lumbis suis.
EZEK|9|4|Et dixit Dominus ad eum: " Transi per mediam civitatem in medio Ierusalem et signa thau super frontes virorum gementium et dolentium super cunctis abominationibus, quae fiunt in medio eius ".
EZEK|9|5|Et illis dixit, audiente me: " Transite per civitatem sequentes eum et percutite; non parcat oculus vester, neque misereamini:
EZEK|9|6|senem, adulescentulum et virginem et parvulum et mulieres interficite usque ad internecionem; omnem autem, super quem videritis thau, ne occidatis, et a sanctuario meo incipite ". Coeperunt ergo a viris senioribus, qui erant ante faciem domus.
EZEK|9|7|Et dixit ad eos: "Contaminate domum et implete atria interfectis. Egredimini ". Et egressi sunt et percutiebant eos, qui erant in civitate.
EZEK|9|8|Et caede completa, remansi ego ruique super faciem meam et clamans aio: Heu, Domine Deus! Ergone disperdes omnes reliquias Israel, effundens furorem tuum super Ierusalem? ".
EZEK|9|9|Et dixit ad me: " Iniquitas domus Israel et Iudae magna est nimis valde; et repleta est terra sanguinibus, et civitas repleta est iniustitia. Dixerunt enim: "Dereliquit Dominus terram, et Dominus non videt";
EZEK|9|10|igitur et meus non parcet oculus, neque miserebor: viam eorum super caput eorum reddam ".
EZEK|9|11|Et ecce vir, qui indutus erat lineis, qui habebat atramentarium in lumbis suis, respondit verbum dicens: " Feci, sicut praecepisti mihi ".
EZEK|10|1|Et vidi: et ecce super fir mamentum, quod erat super caput cherubim, quasi lapis sapphirus, quasi species similitudinis solii apparuit super ea.
EZEK|10|2|Et dixit ad virum, qui indutus erat lineis, et ait: " Ingredere in medio rotarum, quae sunt subtus cherub, et imple manus tuas prunis ignis, quae sunt inter cherubim, et effunde super civitatem ". Ingressusque est in conspectu meo.
EZEK|10|3|Cherubim autem stabant a dextris domus, cum ingrederetur vir, et nubes implevit atrium interius.
EZEK|10|4|Et elevata est gloria Domini desuper cherub ad limen domus, et repleta est domus nube, et atrium repletum est splendore gloriae Domini.
EZEK|10|5|Et sonitus alarum cherubim audiebatur usque ad atrium exterius, quasi vox Dei omnipotentis loquentis.
EZEK|10|6|Cumque praecepisset viro, qui indutus erat lineis, dicens: " Sume ignem de medio rotarum, de medio cherubim ", ingressus ille stetit iuxta rotam;
EZEK|10|7|et extendit cherub manum de medio cherubim ad ignem, qui erat inter cherubim, et sumpsit et dedit in manus eius, qui indutus erat lineis; qui accipiens egressus est.
EZEK|10|8|Et apparuit in cherubim similitudo manus hominis subtus pennas eorum,
EZEK|10|9|et vidi: et ecce quattuor rotae iuxta cherubim; rota una iuxta cherub unum, et rota alia iuxta cherub unum, species autem rotarum erat quasi species lapidis chrysolithi,
EZEK|10|10|et aspectus earum similitudo una illis quattuor, quasi sit rota in medio rotae.
EZEK|10|11|Cumque ambularent in quattuor partes, gradiebantur et non convertebantur ambulantes, sed ad locum, ad quem ire declinabat quae prima erat, sequebantur et ceterae nec convertebantur, cum ambularent.
EZEK|10|12|Et omne corpus eorum et terga et manus et pennae et rotae plena erant oculis in circuitu illis quattuor;
EZEK|10|13|et rotae istae vocatae sunt Volubiles, audiente me.
EZEK|10|14|Quattuor autem facies habebat unumquodque: facies prima facies cherub, et facies secunda facies hominis, et tertia facies leonis, et quarta facies aquilae.
EZEK|10|15|Et elevati sunt cherubim: ipsum est animal, quod videram iuxta fluvium Chobar.
EZEK|10|16|Cumque ambularent, cherubim ibant pariter, et rotae iuxta ea; et cum elevarent cherubim alas suas, ut exaltarentur de terra, non convertebantur rotae, sed et ipsae iuxta erant.
EZEK|10|17|Stantibus illis, stabant et cum elevatis elevabantur; spiritus enim animalium erat in eis.
EZEK|10|18|Et egressa est gloria Domini a limine templi et stetit super cherubim;
EZEK|10|19|et elevantes cherubim alas suas exaltata sunt a terra coram me, et, illis egredientibus, rotae quoque subsecutae sunt; et stetit in introitu portae domus Domini orientalis, et gloria Dei Israel erat super eos.
EZEK|10|20|Ipsum est animal, quod vidi subter Deum Israel iuxta fluvium Chobar, et intellexi quia cherubim essent.
EZEK|10|21|Quattuor per quattuor vultus unicuique, et quattuor alae unicuique, et similitudo manus hominis sub alis eorum;
EZEK|10|22|et similitudo vultuum eorum, ipsi vultus quorum aspectum videram iuxta fluvium Chobar. Et singuli ante faciem suam gradiebantur.
EZEK|11|1|Et elevavit me spiritus et duxit me ad portam domus Domini orientalem, quae respicit solis ortum; et ecce in introitu portae viginti quinque viri, et vidi in medio eorum Iezoniam filium Azur et Pheltiam filium Banaiae, principes populi.
EZEK|11|2|Dixitque ad me: " Fili hominis, hi sunt viri, qui cogitant iniquitatem et tractant consilium pessimum in urbe ista
EZEK|11|3|dicentes: "Nonne dudum aedificatae sunt domus? Haec est lebes, nos autem carnes".
EZEK|11|4|Idcirco vaticinare de eis; vaticinare, fili hominis ".
EZEK|11|5|Et irruit in me spiritus Domini et dixit ad me: " Loquere. Haec dicit Dominus: Sic locuti estis, domus Israel, et cogitationes cordis vestri ego novi.
EZEK|11|6|Plurimos occidistis in urbe hac et implestis vias eius interfectis.
EZEK|11|7|Propterea haec dicit Dominus Deus: Interfecti vestri, quos posuistis in medio eius, hi sunt carnes, et haec est lebes, et educam vos de medio eius.
EZEK|11|8|Gladium metuitis, et gladium inducam super vos, ait Dominus Deus.
EZEK|11|9|Et eiciam vos de medio eius daboque vos in manu hostium et faciam in vobis iudicia.
EZEK|11|10|Gladio cadetis, in finibus Israel iudicabo vos, et scietis quia ego Dominus.
EZEK|11|11|Haec non erit vobis in lebetem, et vos non eritis in medio eius in carnes: in finibus Israel iudicabo vos;
EZEK|11|12|et scietis quia ego Dominus, qui in praeceptis meis non ambulastis et iudicia mea non fecistis, sed iuxta iudicia gentium, quae in circuitu vestro sunt, estis operati ".
EZEK|11|13|Et factum est cum prophetarem, Pheltias filius Banaiae mortuus est; et cecidi in faciem meam, clamans voce magna, et dixi: " Heu, Domine Deus, consummationem tu facis reliquiarum Israel! ".
EZEK|11|14|Et factum est verbum Domini ad me dicens:
EZEK|11|15|" Fili hominis, fratres tui, fratres tui, viri propinqui tui et omnis domus Israel, universi, quibus dixerunt habitatores Ierusalem: "Longe sunt a Domino; nobis data est terra in possessionem".
EZEK|11|16|Propterea haec dicit Dominus Deus: Quia longe feci eos in gentibus et quia dispersi eos in terris, ero eis in sanctificationem modicam in terris, ad quas venerunt.
EZEK|11|17|Propterea loquere: Haec dicit Dominus Deus: Congregabo vos de populis et adunabo de terris, in quibus dispersi estis, daboque vobis humum Israel.
EZEK|11|18|Et ingredientur illuc et auferent omnes offensiones cunctasque abominationes eius de illa.
EZEK|11|19|Et dabo eis cor aliud et spiritum novum tribuam in visceribus eorum; et auferam cor lapideum de carne eorum et dabo eis cor carneum,
EZEK|11|20|ut in praeceptis meis ambulent et iudicia mea custodiant faciantque ea et sint mihi in populum, et ego sim eis in Deum.
EZEK|11|21|Quorum cor post offendicula et abominationes suas ambulat, horum viam in capite suo ponam ", dicit Dominus Deus.
EZEK|11|22|Et elevaverunt cherubim alas suas, et rotae cum eis, et gloria Dei Israel erat super eos;
EZEK|11|23|et ascendit gloria Domini de medio civitatis stetitque super montem, qui est ad orientem urbis.
EZEK|11|24|Et spiritus levavit me adduxitque in Chaldaeam ad transmigrationem in visione in spiritu Dei; et sublata est a me visio, quam videram.
EZEK|11|25|Et locutus sum ad transmigrationem omnia verba Domini, quae ostenderat mihi.
EZEK|12|1|Et factus est sermo Domini ad me dicens:
EZEK|12|2|" Fili hominis, in medio domus exasperantis tu habitas, qui oculos habent ad videndum et non vident, et aures ad audiendum et non audiunt, quia domus exasperans est.
EZEK|12|3|Tu ergo, fili hominis, fac tibi vasa transmigrationis et transmigrabis per diem coram eis; transmigrabis autem de loco tuo ad locum alterum in conspectu eorum, si forte aspiciant, quia domus exasperans est.
EZEK|12|4|Et efferes foras vasa tua quasi vasa transmigrantis per diem in conspectu eorum; tu autem egredieris vespere coram eis, sicut egreditur migrans.
EZEK|12|5|Ante oculos eorum perfode tibi parietem et efferes per eum;
EZEK|12|6|in conspectu eorum in umeris portabis, in caligine efferes: faciem tuam velabis et non videbis terram, quia portentum dedi te domui Israel ".
EZEK|12|7|Feci ergo, sicut praeceperat mihi Dominus: vasa mea protuli quasi vasa transmigrantis per diem et vespere perfodi mihi parietem manu; et in caligine extuli in umeris portans in conspectu eorum.
EZEK|12|8|Et factus est sermo Domini ad me mane dicens:
EZEK|12|9|" Fili hominis, numquid non dixerunt ad te domus Israel, domus exasperans: "Quid tu facis?".
EZEK|12|10|Dic ad eos: Haec dicit Dominus Deus: Super ducem onus istud, qui est in Ierusalem, et super omnem domum Israel, quae est in medio eius.
EZEK|12|11|Dic: Ego portentum vestrum. Quomodo feci, sic fiet illis: in transmigrationem et in captivitatem ibunt.
EZEK|12|12|Et dux, qui est in medio eorum, in umeris portabit, in caligine, et egredietur; parietem perfodient, ut transitus fiat per eum; faciem suam operiet, ut non videat oculo terram.
EZEK|12|13|Et extendam rete meum super illum, et capietur in tendicula mea; et adducam eum in Babylonem in terram Chaldaeorum, et ipsam non videbit ibique morietur.
EZEK|12|14|Et omnes, qui circa eum sunt, praesidium eius et agmina eius, dispergam in omnem ventum; et gladium evaginabo post eos.
EZEK|12|15|Et scient quia ego Dominus, quando dispersero illos in gentibus et disseminavero eos in terris.
EZEK|12|16|Et relinquam ex eis viros paucos a gladio et fame et pestilentia, ut narrent omnia scelera eorum in gentibus, ad quas ingredientur, et scient quia ego Dominus ".
EZEK|12|17|Et factus est sermo Domini ad me dicens:
EZEK|12|18|" Fili hominis, panem tuum in conturbatione comede; sed et aquam tuam in trepidatione et sollicitudine bibe.
EZEK|12|19|Et dices ad populum terrae: Haec dicit Dominus Deus ad eos, qui habitant in Ierusalem in terra Israel: Panem suum in sollicitudine comedent et aquam suam in desolatione bibent, quia desolabitur terra a plenitudine sua propter violentiam omnium, qui habitant in ea;
EZEK|12|20|et civitates, quae nunc habitantur, desolatae erunt, terraque deserta, et scietis quia ego Dominus ".
EZEK|12|21|Et factus est sermo Domini ad me dicens:
EZEK|12|22|" Fili hominis, quod est proverbium istud vobis in terra Israel dicentibus: "In longum differentur dies, et peribit omnis visio"?
EZEK|12|23|Ideo dic ad eos: Haec dicit Dominus Deus: Quiescere faciam proverbium istud, neque vulgo dicetur ultra in Israel; et loquere ad eos quod appropinquaverint dies et sermo omnis visionis.
EZEK|12|24|Non enim erit ultra omnis visio vana neque divinatio ambigua in medio filiorum Israel,
EZEK|12|25|quia ego Dominus loquar; quodcumque locutus fuero verbum, et fiet: non prolongabitur amplius, sed in diebus vestris, domus exasperans, loquar verbum et faciam illud ", dicit Dominus Deus.
EZEK|12|26|Et factus est sermo Domini ad me dicens:
EZEK|12|27|" Fili hominis, ecce domus Israel dicentium: "Visio, quam hic videt, in dies multos et in tempora longa iste prophetat";
EZEK|12|28|propterea dic ad eos: Haec dicit Dominus Deus: Non differetur ultra omnis sermo meus; verbum, quod locutus fuero, complebitur ", dicit Dominus Deus.
EZEK|13|1|Et factus est sermo Domini ad me dicens:
EZEK|13|2|" Fili hominis, vaticinare ad prophetas Israel, qui prophetant; et dices prophetantibus de corde suo: Audite verbum Domini.
EZEK|13|3|Haec dicit Dominus Deus: Vae prophetis insipientibus, qui sequuntur spiritum suum et nihil vident!
EZEK|13|4|Quasi vulpes in ruinis prophetae tui, Israel, facti sunt.
EZEK|13|5|Non ascendistis confractiones neque opposuistis murum pro domo Israel, ut staretis in proelio in die Domini.
EZEK|13|6|Vident vana et divinant mendacium dicentes: "Ait Dominus", cum Dominus non miserit eos; et exspectant, ut confirmet sermonem.
EZEK|13|7|Numquid non visionem cassam vidistis et divinationem mendacem locuti estis, et dicitis: "Ait Dominus", cum ego non sim locutus?
EZEK|13|8|Propterea haec dicit Dominus Deus: Quia locuti estis vana et vidistis mendacium, ideo ecce ego ad vos, ait Dominus Deus;
EZEK|13|9|et erit manus mea super prophetas, qui vident vana et divinant mendacium: in consilio populi mei non erunt et in scriptura domus Israel non scribentur nec in terram Israel ingredientur, et scietis quia ego Dominus Deus.
EZEK|13|10|Eo quod deceperint populum meum dicentes: "Pax", et non est pax; et ipse aedificabat parietem, illi autem liniebant eum calce.
EZEK|13|11|Dic ad eos, qui liniunt calce, quod casurus sit; erit enim imber inundans, et dabo lapides grandinis desuper irruentes et ventum procellae dissipantem.
EZEK|13|12|Siquidem ecce cecidit paries; numquid non dicetur vobis: "Ubi est litura, quam levistis?".
EZEK|13|13|Propterea haec dicit Dominus Deus: Et erumpere faciam spiritum tempestatum in indignatione mea, et imber inundans in furore meo erit, et lapides grandinis in ira in consumptionem;
EZEK|13|14|et destruam parietem, quem levistis calce, et adaequabo eum terrae, et revelabitur fundamentum eius, et cadet, et consumemini in medio eius et scietis quia ego sum Dominus.
EZEK|13|15|Et complebo indignationem meam in pariete et in his, qui leverunt eum calce, dicamque vobis: Non est paries, et non sunt qui leverunt eum;
EZEK|13|16|prophetae Israel, qui prophetant ad Ierusalem et vident ei visionem pacis, et non est pax, ait Dominus Deus.
EZEK|13|17|Et tu, fili hominis, pone faciem tuam contra filias populi tui, quae prophetant de corde suo, et vaticinare super eas
EZEK|13|18|et dic: Haec dicit Dominus Deus: Vae, quae consuunt fascias pro omni articulo manus et faciunt velamina pro capite omnis staturae ad capiendas animas! Numquid capietis animas de populo meo et vivificabitis animas vobis?
EZEK|13|19|Et violastis me ad populum meum pro pugillo hordei et fragmento panis, ut interficeretis animas, quae mori non deberent, et vivificastis animas, quae non deberent vivere, mentientes populo meo credenti mendaciis.
EZEK|13|20|Propter hoc haec dicit Dominus Deus: Ecce ego ad fascias vestras, quibus vos capitis animas quasi volatilia, et disrumpam eas de brachiis vestris; et dimittam animas, quas vos cepistis, animas quasi volatilia,
EZEK|13|21|et disrumpam velamina vestra et liberabo populum meum de manu vestra, neque erunt ultra in manibus vestris ad praedandum, et scietis quia ego Dominus.
EZEK|13|22|Pro eo quod maerere fecistis cor iusti mendaciter, quem ego non contristavi, et confortastis manus impii, ut non reverteretur a via sua mala et viveret,
EZEK|13|23|propterea vana non videbitis et divinationes non divinabitis amplius, et eruam populum meum de manu vestra, et scietis quia ego Dominus ".
EZEK|14|1|Et venerunt ad me viri seniorum Israel et sederunt coram me.
EZEK|14|2|Et factus est sermo Domini ad me dicens:
EZEK|14|3|" Fili hominis, viri isti posuerunt idola sua in cordibus suis et scandalum iniquitatis suae statuerunt contra faciem suam; numquid interrogatus respondebo eis?
EZEK|14|4|Propter hoc loquere eis et dices ad eos: Haec dicit Dominus Deus: Omnis homo de domo Israel, qui posuerit idola sua in corde suo et scandalum iniquitatis suae statuerit contra faciem suam et venerit ad prophetam interrogans per eum me, ego Dominus respondebo ei per me pro multitudine idolorum suorum,
EZEK|14|5|ut capiam domum Israel in corde suo, quo recesserunt a me in cunctis idolis suis.
EZEK|14|6|Propterea dic ad domum Israel: Haec dicit Dominus Deus: Convertimini et recedite ab idolis vestris et ab universis contaminationibus vestris avertite facies vestras.
EZEK|14|7|Quia omnis homo de domo Israel et de advenis, quicumque advena fuerit in Israel, si alienatus fuerit a me et posuerit idola sua in corde suo et scandalum iniquitatis suae statuerit contra faciem suam et venerit ad prophetam, ut interroget per eum me, ego Dominus respondebo ei per me;
EZEK|14|8|et ponam faciem meam contra hominem illum et faciam eum in exemplum et in proberbium et disperdam eum de medio populi mei, et scietis quia ego Dominus.
EZEK|14|9|Et propheta cum erraverit et locutus fuerit verbum, ego Dominus decepi prophetam illum et extendam manum meam contra eum et delebo eum de medio populi mei Israel.
EZEK|14|10|Et portabunt iniquitatem suam: sicut iniquitas interrogantis, sic et iniquitas prophetae erit,
EZEK|14|11|ut non erret ultra domus Israel a me neque polluatur in universis praevaricationibus suis, sed sit mihi in populum, et ego sim eis in Deum, ait Dominus Deus.
EZEK|14|12|Et factus est sermo Domini ad me dicens:
EZEK|14|13|" Fili hominis, terra cum peccaverit mihi, ut praevaricetur praevaricans, extendam manum meam super eam et conteram virgam panis eius et immittam in eam famem et interficiam de ea hominem et iumentum;
EZEK|14|14|et si fuerint tres viri isti in medio eius, Noe, Danel et Iob, ipsi iustitia sua liberabunt animas suas, ait Dominus Deus.
EZEK|14|15|Quod si et bestias pessimas induxero super terram, ut absque liberis faciant eam, et fuerit deserta, in qua nullus pertranseat propter bestias,
EZEK|14|16|tres viri isti si fuerint in ea, vivo ego, dicit Dominus Deus, quia nec filios nec filias liberabunt, sed ipsi soli liberabuntur, terra autem desolabitur.
EZEK|14|17|Vel si gladium induxero super terram illam et dixero gladio: Transi per terram, et interfecero de ea hominem et iumentum,
EZEK|14|18|et tres viri isti fuerint in medio eius, vivo ego, dicit Dominus Deus, non liberabunt filios neque filias, sed ipsi soli liberabuntur.
EZEK|14|19|Vel si pestilentiam immisero super terram illam et effudero indignationem meam super eam in sanguine, ut auferam ex ea hominem et iumentum,
EZEK|14|20|et Noe et Danel et Iob fuerint in medio eius, vivo ego, dicit Dominus Deus, quia filium et filiam non liberabunt, sed ipsi iustitia sua liberabunt animas suas.
EZEK|14|21|Quoniam haec dicit Dominus Deus: Quod si et quattuor iudicia mea pessima, gladium et famem et bestias malas et pestilentiam misero in Ierusalem, ut interficiam de ea hominem et pecus,
EZEK|14|22|tamen relinquetur in ea salvatio educentium filios et filias: ecce ipsi egredientur ad vos, et videbitis viam eorum et opera eorum et consolabimini super malo, quod induxi in Ierusalem in omnibus, quae importavi super eam.
EZEK|14|23|Et consolabuntur vos, cum videritis viam eorum et opera eorum, et cognoscetis quod non frustra fecerim omnia, quae feci in ea ", ait Dominus Deus.
EZEK|15|1|Et factus est sermo Domini ad me dicens:
EZEK|15|2|" Fili hominis, quid habet lignum vitisprae omnibus lignis sarmentorum,quae sunt inter ligna silvarum?
EZEK|15|3|Numquid tolletur de ea lignum,ut fiat opus,aut fabricabitur de ea paxillus,ut dependeat in eo quodcumque vas?
EZEK|15|4|Ecce igni datum est in escam,utramque partem eius consumpsit ignis,et medietas eius adusta est;numquid utile erit ad opus?
EZEK|15|5|Etiam cum esset integrum,non erat aptum ad opus;quanto magis cum ignis illud devoraverit et combusserit,nihil ex eo fiet operis.
EZEK|15|6|Propterea haec dicit Dominus Deus:Quomodo lignum vitis inter ligna silvarum,quod dedi igni ad devorandum,sic tradam habitatores Ierusalem.
EZEK|15|7|Et ponam faciem meam in eos:de igne egressi sunt,et ignis consumet eos.Et scietis quia ego Dominus,cum posuero faciem meam in eos
EZEK|15|8|et dedero terram inviam et desolatam,eo quod praevaricatores exstiterint ",dicit Dominus Deus.
EZEK|16|1|Et factus est sermo Domini ad me dicens:
EZEK|16|2|" Fili hominis, notas fac Ierusalem abominationes suas
EZEK|16|3|et dices: Haec dicit Dominus Deus ad Ierusalem: Radix tua et generatio tua de terra Chanaan, pater tuus Amorraeus et mater tua Hetthaea.
EZEK|16|4|Et quando nata es, in die ortus tui non est praecisus umbilicus tuus, et in aqua non es lota in emundationem nec sale salita nec involuta pannis.
EZEK|16|5|Non pepercit super te oculus, ut faceret tibi unum de his, miseratus tui, sed proiecta es super faciem terrae in abiectione animae tuae in die, qua nata es.
EZEK|16|6|Praeteriens autem te, vidi te palpitare in sanguine tuo et dixi tibi, cum esses in sanguine tuo: Vive. Dixi, inquam, tibi: In sanguine tuo vive.
EZEK|16|7|Crescentem quasi germen agri dedi te, et crevisti et grandis effecta es et pervenisti ad mundum muliebrem: ubera tua intumuerunt, et pilus tuus germinavit; sed eras nuda et confusione plena.
EZEK|16|8|Et transivi per te et vidi te; et ecce tempus tuum, tempus amantium. Et expandi amictum meum super te et operui ignominiam tuam; et iuravi tibi et ingressus sum pactum tecum, ait Dominus Deus, et facta es mea.
EZEK|16|9|Et lavi te aqua et emundavi sanguinem tuum ex te et unxi te oleo;
EZEK|16|10|et vestivi te discoloribus et calceavi te calceis corii delphini et cinxi te bysso et indui te serico.
EZEK|16|11|Et ornavi te ornamento et dedi armillas in manibus tuis et torquem circa collum tuum;
EZEK|16|12|et dedi inaurem super os tuum et circulos auribus tuis et coronam decoris in capite tuo.
EZEK|16|13|Et ornata es auro et argento et vestita es bysso et serico et multicoloribus. Similam et mel et oleum comedisti et decora facta es vehementer nimis et apta ad regnum.
EZEK|16|14|Et egressum est nomen tuum in gentes propter speciem tuam, quia perfecta eras in decore meo, quem posueram super te, dicit Dominus Deus.
EZEK|16|15|Et habens fiduciam in pulchritudine tua fornicata es in nomine tuo et exposuisti fornicationem tuam omni transeunti, quisquis fuerit.
EZEK|16|16|Et sumens de vestimentis tuis fecisti tibi excelsa variegata et fornicata es super eis, sicut non est factum neque futurum est.
EZEK|16|17|Et tulisti vasa decoris tui de auro meo atque argento meo, quae dedi tibi, et fecisti tibi imagines masculinas et fornicata es in eis.
EZEK|16|18|Et sumpsisti vestimenta tua multicoloria et operuisti illas et oleum meum et thymiama meum posuisti coram eis.
EZEK|16|19|Et panem meum, quem dedi tibi, similam et oleum et mel, quibus enutrivi te, posuisti in conspectu eorum in odorem suavitatis, et factum est, ait Dominus Deus.
EZEK|16|20|Et tulisti filios tuos et filias tuas, quas generasti mihi, et immolasti eis ad devorandum. Numquid parva est fornicatio tua?
EZEK|16|21|Immolasti filios meos et dedisti illos consecrans eis.
EZEK|16|22|Et post omnes abominationes tuas et fornicationes non es recordata dierum adulescentiae tuae, quando eras nuda et confusione plena, palpitans in sanguine tuo.
EZEK|16|23|Et accidit post omnem malitiam tuam - vae, vae tibi!, ait Dominus Deus
EZEK|16|24|et aedificasti tibi fornicem et fecisti tibi excelsum in cunctis plateis;
EZEK|16|25|ad omne caput viae aedificasti locum elevatum tuum et abominabilem fecisti decorem tuum et divisisti pedes tuos omni transeunti et multiplicasti fornicationes tuas.
EZEK|16|26|Et fornicata es cum filiis Aegypti vicinis tuis magnorum membrorum et multiplicasti fornicationem tuam ad irritandum me.
EZEK|16|27|Ecce ego extendi manum meam super te et imminui portionem tuam et dedi te in animam odientium te, filiarum Palaestinarum, quae erubescunt in via tua scelerata.
EZEK|16|28|Et fornicata es in filiis Assyriorum, eo quod necdum fueris expleta; et, postquam fornicata es, nec sic es satiata.
EZEK|16|29|Et multiplicasti fornicationem tuam usque ad terram mercatorum Chaldaeam, et nec sic satiata es.
EZEK|16|30|In quo mundabo cor tuum, ait Dominus Deus, cum faceres omnia haec opera mulieris meretricis et procacis?
EZEK|16|31|Quia fabricasti fornicem tuum in capite omnis viae et excelsum tuum fecisti in omni platea; nec facta es quasi meretrix, quia sprevisti pretium.
EZEK|16|32|Mulier adultera loco viri sui accipit alienos.
EZEK|16|33|Omnibus meretricibus dantur mercedes, tu autem dedisti mercedes cunctis amatoribus tuis et donabas eis, ut intrarent ad te undique ad fornicandum tecum.
EZEK|16|34|Factumque in te est contra consuetudinem mulierum in fornicationibus tuis, et post te non sunt fornicati; in eo enim quod dedisti mercedes et mercedes non accepisti, factum est in te contrarium.
EZEK|16|35|Propterea, meretrix, audi verbum Domini.
EZEK|16|36|Haec dicit Dominus Deus: Quia effusum est aes tuum, et revelata est ignominia tua in fornicationibus tuis ad amatores tuos et ad omnia idola abominabilia tua, in sanguine filiorum tuorum, quos dedisti eis,
EZEK|16|37|ideo ecce ego congregabo omnes amatores tuos, quibus iucunda fuisti, et omnes, quos dilexisti, cum universis, quos oderas; et congregabo eos super te undique et nudabo ignominiam tuam coram eis, et videbunt omnem turpitudinem tuam.
EZEK|16|38|Et iudicabo te iudiciis adulterarum et effundentium sanguinem et dabo te in sanguinem furoris et zeli.
EZEK|16|39|Et dabo te in manus eorum, et destruent fornicem tuum et demolientur excelsa tua et denudabunt te vestimentis tuis et auferent vasa decoris tui et derelinquent te nudam plenamque ignominia.
EZEK|16|40|Et convocabunt contra te congregationem et lapidabunt te lapidibus et trucidabunt te gladiis suis.
EZEK|16|41|Et comburent domos tuas igni et facient in te iudicia in oculis mulierum plurimarum; et faciam ut desinas fornicari, et mercedes ultra non dabis.
EZEK|16|42|Et satiabo indignationem meam in te, et auferetur zelus meus a te; et quiescam nec irascar amplius.
EZEK|16|43|Eo quod non fueris recordata dierum adulescentiae tuae et provocasti me in omnibus his, propterea et ego vias tuas in capite tuo dabo, ait Dominus Deus, et non feci iuxta scelera tua in omnibus abominationibus tuis.
EZEK|16|44|Ecce omnis, qui dicit vulgo proverbium in te, assumet illud dicens: Sicut mater, ita et filia eius".
EZEK|16|45|Filia matris tuae es tu, quae sprevit virum suum et filios suos; et soror sororum tuarum es tu, quae spreverunt viros suos et filios suos. Mater vestra Hetthaea, et pater vester Amorraeus.
EZEK|16|46|Et soror tua maior Samaria, ipsa et filiae eius, quae habitat ad sinistram tuam; soror autem tua minor te, quae habitat a dextris tuis, Sodoma et filiae eius.
EZEK|16|47|Sed nec in viis earum ambulasti neque secundum scelera earum fecisti; quasi parum fuisset, sceleratiora fecisti illis in omnibus viis tuis.
EZEK|16|48|Vivo ego, dicit Dominus Deus, non fecit Sodoma soror tua, ipsa et filiae eius, sicut fecisti tu et filiae tuae.
EZEK|16|49|Ecce haec fuit iniquitas Sodomae, sororis tuae: superbia, saturitas panis et securum otium erat ei et filiabus eius, et manum egeni et pauperis non sustentabant;
EZEK|16|50|et elevatae sunt et fecerunt abominationes coram me, et abstuli eas, sicut vidisti.
EZEK|16|51|Et Samaria dimidium peccatorum tuorum non peccavit, sed vicisti eas sceleribus tuis et iustificasti sorores tuas in omnibus abominationibus tuis, quas operata es.
EZEK|16|52|Ergo et tu porta confusionem tuam, quae absolvisti sorores tuas peccatis tuis, sceleratius agens quam illae; iustificatae sunt enim a te. Ergo et tu confundere et porta ignominiam tuam, quae iustificasti sorores tuas.
EZEK|16|53|Et convertam sortem earum, sortem Sodomorum cum filiabus suis et sortem Samariae et filiarum eius; et convertam sortem tuam in medio earum,
EZEK|16|54|ut portes ignominiam tuam et confundaris in omnibus, quae fecisti consolans eas.
EZEK|16|55|Et soror tua Sodoma et filiae eius revertentur ad pristinum statum suum, et Samaria et filiae eius revertentur ad pristinum statum suum, et tu et filiae tuae revertimini ad pristinum statum vestrum.
EZEK|16|56|Nonne fuit Sodoma, soror tua, in fabulam in ore tuo in die superbiae tuae,
EZEK|16|57|antequam revelaretur malitia tua, sicut hoc tempore tu es in opprobrium filiarum Syriae et cunctarum in circuitu tuo filiarum Palaestinarum, quae ambiunt te per gyrum?
EZEK|16|58|Scelus tuum et ignominiam tuam tu portabis, ait Dominus.
EZEK|16|59|Quia haec dicit Dominus Deus: Et faciam tibi, sicut fecisti, qui despexisti iuramentum, ut irritum faceres pactum.
EZEK|16|60|Et recordabor ego pacti mei tecum in diebus adulescentiae tuae et suscitabo tibi pactum sempiternum.
EZEK|16|61|Et recordaberis viarum tuarum et confunderis, cum receperis sorores tuas te maiores cum minoribus tuis, et dabo eas tibi in filias sed non ex pacto tuo.
EZEK|16|62|Et suscitabo ego pactum meum tecum, et scies quia ego Dominus,
EZEK|16|63|ut recorderis et confundaris, et non sit tibi ultra aperire os prae confusione tua, cum placatus fuero tibi in omnibus, quae fecisti ", ait Dominus Deus.
EZEK|17|1|Et factum est verbum Do mini ad me dicens:
EZEK|17|2|"Fili ho minis, propone aenigma et narra parabolam ad domum Israel
EZEK|17|3|et dices:Haec dicit Dominus Deus:Aquila grandismagnarum alarum,longo pennarum ductu,plena plumis et varietate,venit ad Libanumet tulit cacumen cedri;
EZEK|17|4|summitatem frondium eius avellitet transportavit eam in terram Chanaan,in urbem negotiatorum posuit illam.
EZEK|17|5|Et tulit de semine terraeet posuit illud in terra pro semine,super aquas multas,quasi salicem posuit illud,
EZEK|17|6|ut germinaret et cresceret in vineam latioremhumili statura,respicientibus ramis eius ad illam,et radices eius sub illa essent.Facta est ergo vineaet fructificavit in palmiteset emisit propagines.
EZEK|17|7|Et fuit aquila altera grandis,magnis alismultisque plumis;et ecce vinea ista,quasi mittens radices suas ad eam,palmites suos extendit ad illam,ut irrigaret eam abundantiusquam areolae, in quibus erat plantata.
EZEK|17|8|In terra bonasuper aquas multasplantata est,ut faciat frondeset portet fructumet sit in vineam grandem.
EZEK|17|9|Dic: Haec dicit Dominus Deus:Ergone prosperabitur?Nonne radices eius evelletet fructum eius distringet,et marcescent omnia recentia germina eius, et arescet?Et non opus erit brachio grandi neque populo multo,ut evellat eam radicitus.
EZEK|17|10|Ecce plantata est; ergone prosperabitur?Nonne, cum tetigerit eam ventus urens,siccabituret in areis, in quibus germinaverat, arescet? ".
EZEK|17|11|Et factum est verbum Domini ad me dicens:
EZEK|17|12|" Dic ad domum exasperantem: Nescitis quid ista significent? Dic: Ecce venit rex Babylonis Ierusalem et assumpsit regem et principes eius et adduxit eos ad semetipsum in Babylonem;
EZEK|17|13|et tulit de semine regni pepigitque cum eo foedus et accepit ab eo iusiurandum, sed et fortes terrae sustulit,
EZEK|17|14|ut esset regnum humile et non elevaretur, sed custodiret pactum eius et servaret illud.
EZEK|17|15|Qui recedens ab eo, misit nuntios ad Aegyptum, ut daret sibi equos et populum multum. Numquid prosperabitur vel consequetur salutem, qui fecit haec? Et, qui dissolvit pactum, numquid effugiet?
EZEK|17|16|Vivo ego, dicit Dominus Deus, quoniam in loco regis, qui constituit eum regem, cuius fecit irritum iuramentum et solvit pactum, quod habebat cum eo, in medio Babylonis morietur.
EZEK|17|17|Et non in exercitu grandi neque in populo multo adiuvabit eum pharao in proelio, in iactu aggeris et in exstructione munitionum, ut interficiat animas multas.
EZEK|17|18|Spreverat enim iuramentum, ut solveret foedus, et ecce dedit manum suam et, cum omnia haec fecerit, non effugiet.
EZEK|17|19|Propterea haec dicit Dominus Deus: Vivo ego, quoniam iuramentum meum, quod sprevit, et foedus meum, quod praevaricatus est, ponam in caput eius
EZEK|17|20|et expandam super eum rete meum, et comprehendetur tendicula mea, et adducam eum in Babylonem et iudicabo illum ibi in praevaricatione, qua praevaricatus est in me.
EZEK|17|21|Et omnes electi eius in universo agmine suo gladio cadent; residui autem in omnem ventum dispergentur, et scietis quia ego Dominus locutus sum.
EZEK|17|22|Haec dicit Dominus Deus:Et sumam ego de cacumine cedri sublimis et ponam;de vertice ramorum eius tenerum distringamet plantabo super montem excelsum et eminentem.
EZEK|17|23|In monte sublimi Israel plantabo illud;et erumpet in germen et faciet fructumet erit in cedrum magnam;et habitabunt sub ea omnes volucres,et universum volatile sub umbra frondium eius nidificabit.
EZEK|17|24|Et scient omnia ligna regionisquia ego Dominushumiliavi lignum sublimeet exaltavi lignum humileet siccavi lignum virideet frondere feci lignum aridum.Ego Dominus locutus sum et feci ".
EZEK|18|1|Et factus est sermo Domini ad me dicens:
EZEK|18|2|"Quid est vo bis quod vulgo dicitis proverbium istud in terra Israel dicentes:Patres comederunt uvam acerbam,et dentes filiorum obstupescunt"?
EZEK|18|3|Vivo ego, dicit Dominus Deus, non dicetis ultra hoc proverbium in Israel.
EZEK|18|4|Ecce omnes animae meae sunt: ut anima patris, ita et anima filii mea est; anima, quae peccaverit, ipsa morietur.
EZEK|18|5|Et vir, si fuerit iustus et fecerit iudicium et iustitiam,
EZEK|18|6|in montibus non comederit et oculos suos non levaverit ad idola domus Israel et uxorem proximi sui non violaverit et ad mulierem menstruatam non accesserit
EZEK|18|7|et hominem non afflixerit, pignus debitori reddiderit, per vim nihil rapuerit, panem suum esurienti dederit et nudum operuerit vestimento,
EZEK|18|8|ad usuram non commodaverit et fenus non acceperit, ab iniquitate averterit manum suam, iudicium verum fecerit inter virum et virum,
EZEK|18|9|in praeceptis meis ambulaverit et iudicia mea custodierit, ut faciat veritatem, hic iustus est, vita vivet, ait Dominus Deus.
EZEK|18|10|Quod si genuerit filium latronem, effundentem sanguinem et facientem unum de istis,
EZEK|18|11|cum ipse haec omnia non fecerit, et etiam in montibus comedentem et uxorem proximi sui polluentem,
EZEK|18|12|egenum et pauperem affligentem, rapientem rapinas, pignus non reddentem et ad idola levantem oculos suos, abominationem facientem,
EZEK|18|13|ad usuram dantem et fenus accipientem, numquid vivet? Non vivet. Cum universa detestanda haec fecerit, morte morietur; sanguis eius in ipso erit.
EZEK|18|14|Quod si genuerit filium, qui videns omnia peccata patris sui, quae fecit, timuerit et non fecerit simile eis:
EZEK|18|15|super montes non comederit et oculos suos non levaverit ad idola domus Israel et uxorem proximi sui non violaverit
EZEK|18|16|et virum non afflixerit, pignus non retinuerit et rapinam non rapuerit, panem suum esurienti dederit et nudum operuerit vestimento,
EZEK|18|17|ab iniuria averterit manum suam, usuram et fenus non acceperit, iudicia mea fecerit, in praeceptis meis ambulaverit, hic non morietur in iniquitate patris sui, sed vita vivet.
EZEK|18|18|Pater eius, quia calumniatus est et fecit rapinas nec bonum operatus est in medio populi sui, ecce mortuus est in iniquitate sua.
EZEK|18|19|Et dicitis: "Quare non portavit filius iniquitatem patris?". Videlicet, quia filius iudicium et iustitiam operatus est, omnia praecepta mea custodivit et fecit illa, vivet vita.
EZEK|18|20|Anima, quae peccaverit, ipsa morietur; filius non portabit iniquitatem patris, et pater non portabit iniquitatem filii. Iustitia iusti super eum erit, et impietas impii erit super eum.
EZEK|18|21|Si autem impius egerit paenitentiam ab omnibus peccatis suis, quae operatus est, et custodierit universa praecepta mea et fecerit iudicium et iustitiam, vita vivet, non morietur.
EZEK|18|22|Omnes iniquitates eius, quas operatus est, non memorabuntur ei; in iustitia sua, quam operatus est, vivet.
EZEK|18|23|Numquid voluntatis meae est mors impii, dicit Dominus Deus, et non ut convertatur a viis suis et vivat?
EZEK|18|24|Si autem averterit se iustus a iustitia sua et fecerit iniquitatem secundum omnes abominationes, quas operari solet impius, numquid vivet? Omnes iustitiae eius, quas fecerat, non recordabuntur; in praevaricatione, qua praevaricatus est, et in peccato suo, quod peccavit, in ipsis morietur.
EZEK|18|25|Et dixistis: "Non est aequa via Domini". Audite ergo, domus Israel: Numquid via mea non est aequa, et non magis viae vestrae pravae sunt?
EZEK|18|26|Cum enim averterit se iustus a iustitia sua et fecerit iniquitatem, morietur; in iniustitia, quam operatus est, morietur.
EZEK|18|27|Et cum averterit se impius ab impietate sua, quam operatus est, et fecerit iudicium et iustitiam, ipse animam suam vivificabit;
EZEK|18|28|considerans enim et avertens se ab omnibus iniquitatibus suis, quas operatus est, vita vivet, non morietur.
EZEK|18|29|Et dicunt domus Israel: "Non est aequa via Domini". Numquid viae meae non sunt aequae, domus Israel, et non magis viae vestrae pravae?
EZEK|18|30|Idcirco unumquemque iuxta vias suas iudicabo, domus Israel, ait Dominus Deus. Convertimini et agite paenitentiam ab omnibus iniquitatibus vestris, et non erit vobis in scandalum iniquitatis.
EZEK|18|31|Proicite a vobis omnes praevaricationes vestras, in quibus praevaricati estis, et facite vobis cor novum et spiritum novum. Et quare moriemini, domus Israel?
EZEK|18|32|Quia nolo mortem morientis, dicit Dominus Deus. Revertimini et vivite.
EZEK|19|1|Et tu, assume planctum super principes Israel
EZEK|19|2|et dices:Qualis erat mater tua leaenainter leones!Cubavit in medio leunculorum,enutrivit catulos suos.
EZEK|19|3|Et educavit unum de leunculis suis;leo factus estet didicit capere praedam,homines devoravit.
EZEK|19|4|Et convocaverunt contra eum gentes,in fovea earum captus est;et adduxerunt eum in circulisin terram Aegypti.
EZEK|19|5|Quae cum vidisset quoniam exspectaverat,et perierat spes eius,tulit alium de leunculis suis,leonem constituit eum.
EZEK|19|6|Qui incedebat inter leones,factus est leoet didicit praedam capere,homines devoravit;
EZEK|19|7|et fregit arces eorumet civitates eorum vastavit.Et obstupuit terra et plenitudo eiusa voce rugitus illius.
EZEK|19|8|Et convenerunt adversum eum gentesundique de provinciiset expanderunt super eum rete suum,in fovea earum captus est.
EZEK|19|9|Et miserunt eum in caveam in circuliset adduxerunt eum ad regem Babylonis;qui misit eum in carcerem,ne audiretur vox eius ultrasuper montes Israel.
EZEK|19|10|Mater tua vineae assimilabatursuper aquam plantata.Fructus eius et frondes eius creveruntex aquis multis;
EZEK|19|11|et factae sunt ei virgae solidaein sceptra dominantium,et exaltata est statura eiususque in nubes,et apparuit in altitudine sua,in multitudine palmitum suorum.
EZEK|19|12|Et evulsa est in irain terramque proiecta,et ventus urens siccavit fructum eius;abrepta et arefacta est virga roboris eius,ignis comedit eam.
EZEK|19|13|Et nunc transplantata est in desertum,in terra invia et sitienti.
EZEK|19|14|Et egressus est ignis de virga ramorum eius,qui fructum eius comedit;et non fuit in ea virga fortis,sceptrum regni ".Planctus est, et erit in planctum.
EZEK|20|1|Et factum est in anno sep timo, in quinto mense, in de cima mensis, venerunt viri de senioribus Israel, ut interrogarent Dominum, et sederunt coram me.
EZEK|20|2|Et factus est sermo Domini ad me dicens:
EZEK|20|3|" Fili hominis, loquere senioribus Israel et dices ad eos: Haec dicit Dominus Deus: Num ad interrogandum me vos venistis? Vivo ego, quia non respondebo vobis, ait Dominus Deus.
EZEK|20|4|Numquid iudicabis eos, numquid iudicabis, fili hominis? Abominationes patrum eorum ostende eis.
EZEK|20|5|Et dices ad eos: Haec dicit Dominus Deus: In die qua elegi Israel et levavi manum meam pro stirpe domus Iacob et apparui eis in terra Aegypti et levavi manum meam pro eis dicens: Ego Dominus Deus vester;
EZEK|20|6|in die illa levavi manum meam pro eis, ut educerem eos de terra Aegypti in terram, quam provideram eis fluentem lacte et melle, quae est egregia inter omnes terras.
EZEK|20|7|Et dixi ad eos: Unusquisque abominationes oculorum suorum abiciat, et in idolis Aegypti nolite pollui: ego Dominus Deus vester.
EZEK|20|8|Et irritaverunt me nolueruntque me audire; unusquisque abominationes oculorum suorum non proiecit, nec idola Aegypti reliquerunt. Et dixi, ut effunderem indignationem meam super eos et consummarem iram meam in eis in medio terrae Aegypti.
EZEK|20|9|Et feci propter nomen meum, ut non violaretur coram gentibus, in quarum medio erant, et inter quas apparui eis, ut educerem eos de terra Aegypti.
EZEK|20|10|Eduxi ergo eos de terra Aegypti et duxi in desertum.
EZEK|20|11|Et dedi eis praecepta mea et iudicia mea ostendi eis, quae faciat homo et vivat in eis.
EZEK|20|12|Insuper et sabbata mea dedi eis, ut essent signum inter me et eos, et scirent quia ego Dominus sanctificans eos.
EZEK|20|13|Et irritaverunt me domus Israel in deserto: in praeceptis meis non ambulaverunt et iudicia mea proiecerunt, quae faciens homo vivet in eis, et sabbata mea violaverunt vehementer. Dixi ergo, ut effunderem furorem meum super eos in deserto et consumerem eos.
EZEK|20|14|Et feci propter nomen meum, ne violaretur coram gentibus, de quibus eduxi eos in conspectu earum.
EZEK|20|15|Attamen ego levavi quoque manum meam super eos in deserto, ne inducerem eos in terram, quam dedi eis fluentem lacte et melle, praecipuam terrarum omnium;
EZEK|20|16|quia iudicia mea proiecerunt et in praeceptis meis non ambulaverunt et sabbata mea violaverunt, post idola enim sua cor eorum gradiebatur.
EZEK|20|17|Et pepercit oculus meus super eos, ut non interficerem eos; nec consumpsi eos in deserto.
EZEK|20|18|Dixi autem ad filios eorum in solitudine: In praeceptis patrum vestrorum nolite incedere nec iudicia eorum custodiatis nec in idolis eorum polluamini.
EZEK|20|19|Ego Dominus Deus vester. In praeceptis meis ambulate et iudicia mea custodite et facite ea
EZEK|20|20|et sabbata mea sanctificate, ut sint signum inter me et vos, et sciatur quia ego Dominus Deus vester.
EZEK|20|21|Et exacerbaverunt me filii; in praeceptis meis non ambulaverunt et iudicia mea non custodierunt, ut facerent ea, quae cum fecerit homo, vivet in eis, et sabbata mea violaverunt. Et comminatus sum, ut effunderem furorem meum super eos et consummarem iram meam in eis in deserto.
EZEK|20|22|Averti autem manum meam et feci propter nomen meum, ut non violaretur coram gentibus, de quibus eduxi eos in oculis earum.
EZEK|20|23|Iterum levavi manum meam in eos in solitudine, ut dispergerem illos in nationes et ventilarem in terras,
EZEK|20|24|eo quod iudicia mea non fecissent et praecepta mea reprobassent et sabbata mea violassent et post idola patrum suorum fuissent oculi eorum.
EZEK|20|25|Ergo et ego dedi eis praecepta non bona et iudicia, in quibus non vivent;
EZEK|20|26|et pollui eos in muneribus suis, cum offerrent omne, quod aperit vulvam, ut horrorem eis incuterem, et sciant quia ego Dominus.
EZEK|20|27|Quam ob rem loquere ad domum Israel, fili hominis, et dices ad eos: Haec dicit Dominus Deus: Adhuc et in hoc blasphemaverunt me patres vestri, cum sprevissent me contemnentes,
EZEK|20|28|et induxissem eos in terram, super quam levavi manum meam, ut darem eis. Viderunt omnem collem excelsum et omne lignum nemorosum et immolaverunt ibi victimas suas et dederunt ibi irritationem oblationis suae et posuerunt ibi odorem suavitatis suae et libaverunt libationes suas.
EZEK|20|29|Et dixi ad eos: Quid est excelsum, ad quod vos ingredimini? Et vocatum est nomen eius Excelsum usque ad hanc diem.
EZEK|20|30|Propterea dic ad domum Israel: Haec dicit Dominus Deus: Certe in via patrum vestrorum vos polluimini et post offendicula eorum vos fornicamini
EZEK|20|31|et in oblatione donorum vestrorum, cum traducitis filios vestros per ignem; vos polluimini in omnibus idolis vestris usque hodie, et ego respondebo vobis, domus Israel? Vivo ego, dicit Dominus Deus, quia non respondebo vobis.
EZEK|20|32|Neque cogitatio mentis vestrae fiet dicentium: "Erimus sicut gentes et sicut cognationes terrarum, ut colamus ligna et lapides".
EZEK|20|33|Vivo ego, dicit Dominus Deus, quoniam in manu forti et brachio extento et in furore effuso regnabo super vos.
EZEK|20|34|Et educam vos de populis et congregabo vos de terris, in quibus dispersi estis; in manu valida et brachio extento et in furore effuso.
EZEK|20|35|Et adducam vos in desertum populorum et iudicio contendam vobiscum ibi facie ad faciem.
EZEK|20|36|Sicut iudicio contendi adversum patres vestros in deserto terrae Aegypti, sic iudicio contendam vobiscum, dicit Dominus Deus,
EZEK|20|37|et transire vos faciam sub baculo meo et inducam vos in vinculis foederis.
EZEK|20|38|Et segregabo de vobis transgressores et impios et de terra incolatus eorum educam eos, et terram Israel non ingredientur, et scietis quia ego Dominus.
EZEK|20|39|Et vos, domus Israel, haec dicit Dominus Deus: Singuli post idola vestra ambulate et servite eis. Sed postea nonne audietis me et nomen meum sanctum non polluetis ultra in muneribus vestris et in idolis vestris?
EZEK|20|40|In monte enim sancto meo, in monte excelso Israel, ait Dominus Deus, ibi serviet mihi omnis domus Israel: omnes, inquam, in terra, in qua placebunt mihi; et ibi quaeram donaria vestra et primitias oblationum vestrarum in omnibus sanctificationibus vestris.
EZEK|20|41|In odorem suavitatis suscipiam vos, cum eduxero vos de populis et congregavero vos de terris, in quas dispersi estis, et sanctificabor in vobis in oculis nationum.
EZEK|20|42|Et scietis quia ego Dominus, cum induxero vos ad terram Israel, in terram, pro qua levavi manum meam, ut darem eam patribus vestris.
EZEK|20|43|Et recordabimini ibi viarum vestrarum et omnium scelerum vestrorum, quibus polluti estis, et displicebitis vobis in conspectu vestro in omnibus malitiis vestris, quas fecistis.
EZEK|20|44|Et scietis quia ego Dominus, cum benefecero vobis propter nomen meum, non secundum vias vestras malas neque secundum scelera vestra pessima, domus Israel ", ait Dominus Deus.
EZEK|21|1|Et factus est sermo Domini ad me dicens:
EZEK|21|2|" Fili hominis, pone faciem tuam contra meridiem et stilla ad austrum et propheta ad saltum agri Nageb.
EZEK|21|3|Et dices saltui Nageb: Audi verbum Domini. Haec dicit Dominus Deus: Ecce ego succendam in te ignem, et comburet in te omne lignum viride et omne lignum aridum; non exstinguetur flamma succensionis, et comburetur in ea omnis facies ab austro usque ad aquilonem.
EZEK|21|4|Et videbit universa caro quia ego Domínus succendi eam, nec exstinguetur.
EZEK|21|5|Et dixi: " Heu, Domine Deus! Ipsi dicunt de me: "Numquid non per parabolas loquitur iste?" ".
EZEK|21|6|Et factus est sermo Domini ad me dicens:
EZEK|21|7|" Fili hominis, pone faciem tuam ad Ierusalem et stilla ad sanctuaria et propheta contra humum Israel.
EZEK|21|8|Et dices terrae Israel: Haec dicit Dominus Deus: Ecce ego ad te, et eiciam gladium meum de vagina sua et occidam in te iustum et impium.
EZEK|21|9|Pro eo autem quod occidi in te iustum et impium, idcirco egredietur gladius meus de vagina sua ad omnem carnem, ab austro ad aquilonem,
EZEK|21|10|ut sciat omnis caro quia ego Dominus eduxi gladium meum de vagina sua irrevocabilem.
EZEK|21|11|Et tu, fili hominis, ingemisce in contritione lumborum et in amaritudinibus ingemisce coram eis.
EZEK|21|12|Cumque dixerint ad te: "Quare tu gemis?", dices: Pro auditu quia venit et tabescet omne cor, et dissolventur universae manus, et infirmabitur omnis spiritus, et per cuncta genua fluent aquae; ecce venit et fiet ", ait Dominus Deus.
EZEK|21|13|Et factus est sermo Domini ad me dicens:
EZEK|21|14|" Fili hominis, propheta et dices: Haec dicit Dominus Deus: Loquere:Gladius, gladius exacutus estet etiam limatus;
EZEK|21|15|ut caedat victimas exacutus est,ut splendeat limatus est.
EZEK|21|16|Et datus est ad levigandum,ut teneatur manu.Iste exacutus est gladius et iste limatus,ut sit in manu interficientis.
EZEK|21|17|Clama et ulula, fili hominis,quia hic directus est in populum meum,hic in cunctos duces Israel,qui gladio traditi sunt cum populo meo.
EZEK|21|18|Idcirco plaude super femur,quia probatio est,dicit Dominus Deus.
EZEK|21|19|Tu ergo, fili hominis,propheta et percute manu ad manum.Et duplicetur gladius,ac triplicetur gladius interfectorum: hic est gladius occisionis magnae,qui eos circumdat,
EZEK|21|20|ut cor tabescat,et multiplicentur corruentes.In omnibus portis eorumdedi occisionem gladii:eheu, facti acuti et limati ad fulgendum,politi ad caedem!
EZEK|21|21|"Exacuere, vade ad dexteram sive ad sinistram,quocumque acies tuae sunt destinatae".
EZEK|21|22|Quin et ego plaudam manu ad manumet saturabo indignationem meam,ego Dominus locutus sum ".
EZEK|21|23|Et factus est sermo Domini ad me dicens:
EZEK|21|24|"Et tu, fili hominis, pone tibi duas vias, ut veniat gladius regis Babylonis: de terra una egrediantur ambae; et indicem statue, in capite viae civitatis statue.
EZEK|21|25|Viam pones, quo veniat gladius, ad Rabba filiorum Ammon et ad Iudam in Ierusalem munitissimam.
EZEK|21|26|Stat enim rex Babylonis in bivio in capite duarum viarum, divinationem quaerens, commiscens sagittas; interrogat teraphim, iecur consulit.
EZEK|21|27|Ad dexteram eius facta est divinatio super Ierusalem, ut ponat arietes, ut aperiat os ad caedem, ut elevet vocem in ululatu, ut ponat arietes contra portas, ut comportet aggerem, ut aedificet munitiones.
EZEK|21|28|Eritque quasi consulens frustra oraculum in oculis eorum, et iuramenta sanctissima sunt eis; ipse autem in memoriam revocabit iniquitatem ad capiendum.
EZEK|21|29|Idcirco haec dicit Dominus Deus: Pro eo quod in memoriam revocastis iniquitatem vestram, et revelatae sunt praevaricationes vestrae, et apparuerunt peccata vestra in omnibus operibus vestris; pro eo, inquam, quod in memoriam revocati estis, manu capiemini.
EZEK|21|30|Tu autem, profane, impie dux Israel, cuius venit dies in tempore iniquitatis finitae -
EZEK|21|31|haec dicit Dominus Deus - auferatur cidaris, tollatur corona; hoc non erit amplius. Humile sublevetur, et sublime humilietur.
EZEK|21|32|Ruinam, ruinam, ruinam ponam illud; et hoc non fiet, donec veniat, cuius est iudicium, et tradam ei.
EZEK|21|33|Et tu, fili hominis, propheta et dic: Haec dicit Dominus Deus ad filios Ammon et ad opprobrium eorum; et dices: Gladius, gladius est evaginatus ad occidendum, limatus ad consumendum, ut fulgeat,
EZEK|21|34|cum tibi videntur vana, et divinantur mendacia, ut ponatur gladius ad colla profanorum impiorum, quorum venit dies in tempore iniquitatis finitae.
EZEK|21|35|Revertatur ad vaginam suam. In loco, in quo creatus es, in terra nativitatis tuae iudicabo te.
EZEK|21|36|Et effundam super te indignationem meam, in igne furoris mei sufflabo in te; daboque te in manus hominum insipientium et fabricantium interitum.
EZEK|21|37|Igni eris cibus, sanguis tuus erit in medio terrae; oblivioni traderis, quia ego Dominus locutus sum ".
EZEK|22|1|Et factum est verbum Do mini ad me dicens:
EZEK|22|2|" Et tu, fili hominis, num iudicas, num iudicas civitatem sanguinum?
EZEK|22|3|Et ostendes ei omnes abominationes suas et dices: Haec dicit Dominus Deus: Civitas effundens sanguinem in medio sui, ut veniat tempus eius et, quae fecit idola contra semetipsam, ut pollueretur.
EZEK|22|4|In sanguine tuo, qui a te effusus est, deliquisti; et in idolis tuis, quae fecisti, polluta es; et appropinquare fecisti dies tuos et adduxisti tempus annorum tuorum. Propterea dedi te opprobrium gentibus et irrisionem universis terris.
EZEK|22|5|Quae iuxta sunt et quae procul a te, triumphabunt de te, sordibus famosa, grandis tumultu.
EZEK|22|6|Ecce principes Israel singuli pro brachio suo fuerunt in te ad effundendum sanguinem.
EZEK|22|7|Pater et mater contempti sunt in te, advena oppressus est in medio tui, pupillum et viduam afflixerunt apud te.
EZEK|22|8|Sanctuaria mea sprevisti et sabbata mea profanasti.
EZEK|22|9|Viri detractores fuerunt in te ad effundendum sanguinem et super montes comederunt in te; scelus operati sunt in medio tui.
EZEK|22|10|Verecundiora patris discooperuerunt in te, immunditiam menstruatae humiliaverunt in te;
EZEK|22|11|et unus in uxorem proximi sui operatus est abominationem, et alter nurum suam polluit nefarie; frater sororem suam, filiam patris sui, oppressit in te.
EZEK|22|12|Munera acceperunt apud te ad effundendum sanguinem, usuram et fenus accepisti et avare proximos tuos calumniabaris meique oblita es, ait Dominus Deus.
EZEK|22|13|Ecce complosi manus meas super lucrum tuum, quod fecisti, et super sanguinem, qui effusus est in medio tui.
EZEK|22|14|Numquid sustinebit cor tuum, aut praevalebunt manus tuae in diebus, quos ego faciam tibi? Ego Dominus locutus sum et faciam;
EZEK|22|15|et dispergam te in nationes et ventilabo te in terras et deficere faciam immunditiam tuam a te:
EZEK|22|16|et profanabo me in te in conspectu gentium, et scies quia ego Dominus.
EZEK|22|17|Et factum est verbum Domini ad me dicens:
EZEK|22|18|" Fili hominis, versa est mihi domus Israel in scoriam; omnes isti argentum et aes et stannum et ferrum et plumbum in medio fornacis, scoria facti sunt.
EZEK|22|19|Propterea haec dicit Dominus Deus: Eo quod versi estis omnes in scoriam, propterea ecce ego congregabo vos in medio Ierusalem
EZEK|22|20|congregatione argenti et aeris et ferri et plumbi et stanni in medio fornacis, ut succendatur in ea ignis ad conflandum: sic congregabo in furore meo et in ira mea et ponam et conflabo vos
EZEK|22|21|et congregabo vos et succendam vos in igne furoris mei, et conflabimini in medio eius.
EZEK|22|22|Ut conflatur argentum in medio fornacis, sic conflabimini in medio eius; et scietis quia ego Dominus effuderim indignationem meam super vos.
EZEK|22|23|Et factum est verbum Domini ad me dicens:
EZEK|22|24|" Fili hominis, dic ei: Tu es terra, super quam non cecidit pluvia neque imber in die furoris,
EZEK|22|25|cuius duces in medio eius sicut leo rugiens capiensque praedam: animas devoraverunt, opes et pretium acceperunt, viduas eius multiplicaverunt in medio illius.
EZEK|22|26|Sacerdotes eius contempserunt legem meam et polluerunt sanctuaria mea, inter sanctum et profanum non habuerunt distantiam et inter pollutum et mundum non docuerunt distinguere et a sabbatis meis averterunt oculos suos, et coinquinabar in medio eorum.
EZEK|22|27|Principes eius in medio illius quasi lupi rapientes praedam ad effundendum sanguinem et perdendas animas et avare sectanda lucra.
EZEK|22|28|Prophetae autem eius liniebant eis omnia calce, videntes vana et divinantes eis mendacium, dicentes: "Haec dicit Dominus Deus", cum Dominus non sit locutus.
EZEK|22|29|Populus terrae calumniabatur calumniam et rapiebat violenter; egenum et pauperem affligebant et advenam opprimebant absque iudicio.
EZEK|22|30|Et quaesivi de eis virum, qui interponeret saepem et staret in confractione contra me pro terra, ne dissiparem eam, et non inveni.
EZEK|22|31|Et effudi super eos indignationem meam, in igne irae meae consumpsi eos, viam eorum in caput eorum reddidi ", ait Dominus Deus.
EZEK|23|1|Et factus est sermo Domini ad me dicens:
EZEK|23|2|" Fili hominis, duae mulieres filiae matris unius fuerunt
EZEK|23|3|et fornicatae sunt in Aegypto, in adulescentia sua fornicatae sunt; ibi subacta sunt ubera earum, et tactae sunt mammae virginitatis earum.
EZEK|23|4|Nomina autem earum Oolla maior et Ooliba soror eius; et habui eas, et pepererunt filios et filias: porro earum nomina Samaria Oolla et Ierusalem Ooliba.
EZEK|23|5|Fornicata est igitur Oolla discedens a me; et insanivit in amatores suos, in Assyrios: bellatores
EZEK|23|6|vestitos hyacintho, principes et magistratus, iuvenes desiderabiles universi, equites ascensores equorum.
EZEK|23|7|Et dedit fornicationes suas ad eos electos filiorum Assyriae universos; et apud omnes, in quos insanivit, in omnibus idolis eorum polluta est.
EZEK|23|8|Insuper et fornicationes suas, quas habuerat in Aegypto, non reliquit; nam et illi dormierunt cum ea in adulescentia eius, et illi tetigerant ubera virginitatis eius et effuderant fornicationem suam super eam.
EZEK|23|9|Propterea tradidi eam in manus amatorum suorum, in manus filiorum Assyriae, in quos insanivit;
EZEK|23|10|ipsi discooperuerunt ignominiam eius, filios et filias illius tulerunt et ipsam occiderunt gladio; et facta est famosa mulieribus, et iudicia perpetrarunt in ea.
EZEK|23|11|Quod cum vidisset soror eius Ooliba, plus quam illa insanivit libidine et fornicatione sua super fornicationem sororis suae.
EZEK|23|12|In filios Assyriorum amore exarsit: duces et magistratus, bellatores indutos veste pretiosa, equites, qui vectabantur equis, adulescentes cuncti desiderabiles.
EZEK|23|13|Et vidi quod polluta esset: via una ambarum;
EZEK|23|14|et auxit fornicationes suas. Cumque vidisset viros depictos in pariete, imagines Chaldaeorum expressas sinopide,
EZEK|23|15|et accinctos balteis renes, et tiaras defluentes in capitibus eorum; aspectus essedariorum omnibus, similitudo filiorum Babylonis, quorum patria Chaldaea.
EZEK|23|16|Et insanivit super eos concupiscentia oculorum suorum et misit nuntios ad eos in Chaldaeam.
EZEK|23|17|Cumque venissent ad eam filii Babylonis ad cubile amoris, polluerunt eam stupris suis; et, cum polluta esset ab eis, recessit anima eius ab illis.
EZEK|23|18|Cum manifestasset fornicationes suas et discooperuisset ignominiam suam, recessit anima mea ab ea, sicut recesserat anima mea a sorore eius.
EZEK|23|19|Multiplicavit autem fornicationes suas, recordans dies adulescentiae suae, quibus fornicata est in terra Aegypti;
EZEK|23|20|et insanivit libidine in amatores suos, quorum membra sunt ut membra asinorum, et sicut fluxus equorum fluxus eorum.
EZEK|23|21|Et desiderasti scelus adulescentiae tuae, quando subacta sunt in Aegypto ubera tua, et tactae mammae pubertatis tuae.
EZEK|23|22|Propterea, Ooliba, haec dicit Dominus Deus: Ecce ego suscitabo amatores tuos contra te, de quibus recessit anima tua; et congregabo eos adversum te in circuitu,
EZEK|23|23|filios Babylonis et universos Chaldaeos, Phacud et Sue et Cue, omnes filios Assyriorum cum eis, iuvenes desiderabiles, duces et magistratus universos, essedarios et nominatos, ascensores equorum omnes.
EZEK|23|24|Et venient super te instructi curru et rota, cum multitudine populorum; scuto et clipeo et galea armabuntur contra te undique, et dabo coram eis iudicium, et iudicabunt te iudiciis suis.
EZEK|23|25|Et ponam zelum meum in te, quem exercent tecum in furore: nasum tuum et aures tuas praecident et, quae remanserint de te, gladio concident; ipsi filios tuos et filias tuas capient, et novissimum tuum devorabitur igni.
EZEK|23|26|Et denudabunt te vestimentis tuis et tollent vasa gloriae tuae;
EZEK|23|27|et cessare faciam scelus tuum de te et fornicationem tuam de terra Aegypti, nec levabis oculos tuos ad eos et Aegypti non recordaberis amplius.
EZEK|23|28|Quia haec dicit Dominus Deus: Ecce ego tradam te in manu eorum, quos odisti, in manu, de quibus recessit anima tua;
EZEK|23|29|et agent tecum in odio et tollent omnes labores tuos et dimittent te nudam et ignominia plenam, et revelabitur ignominia fornicationum tuarum, scelus tuum et fornicationes tuae.
EZEK|23|30|Fecerunt haec tibi, quia fornicata es post gentes, inter quas polluta es in idolis earum.
EZEK|23|31|In via sororis tuae ambulasti, et dabo calicem eius in manu tua.
EZEK|23|32|Haec dicit Dominus Deus:Calicem sororis tuae bibesprofundum et latumC eris in derisum et in subsannationem C:est capacissimus.
EZEK|23|33|Ebrietate et dolore repleberis,calice stuporis et horroris,calice sororis tuae Samariae,
EZEK|23|34|et bibes illum et epotabis usque ad faeces;et fragmenta eius rodeset ubera tua lacerabis,quia ego locutus sum ",ait Dominus Deus.
EZEK|23|35|Propterea haec dicit Dominus Deus: " Quia oblita es mei et proiecisti me post tergum tuum, tu quoque porta scelus tuum et fornicationes tuas ".
EZEK|23|36|Et ait Dominus ad me: " Fili hominis, numquid iudicas Oollam et Oolibam? Annuntia ergo eis scelera earum.
EZEK|23|37|Quia adulteratae sunt, et sanguis in manibus earum, et cum idolis suis fornicatae sunt; insuper et filios suos, quos genuerunt mihi, obtulerunt eis ad devorandum.
EZEK|23|38|Sed et hoc fecerunt mihi: polluerunt sanctuarium meum in die illa et sabbata mea profanaverunt.
EZEK|23|39|Cumque immolarent filios suos idolis suis et ingrederentur sanctuarium meum in die illa, ut polluerent illud, ecce haec fecerunt in medio domus meae.
EZEK|23|40|Quin et miserunt ad viros venientes de longe, ad quos nuntius missus erat; itaque ecce venerunt. Quibus te lavisti et circumlevisti stibio oculos tuos et ornata es mundo muliebri;
EZEK|23|41|sedisti in lecto pulcherrimo, et mensa ornata est ante te, thymiama meum et unguentum meum posuisti super eam.
EZEK|23|42|Et vox multitudinis exsultantis erat apud eam et apud viros multitudo hominum, qui adducebantur de deserto; et posuerunt armillas in manibus earum et coronas speciosas in capitibus earum.
EZEK|23|43|Et dixi de ea, quae attrita est in adulteriis: Nunc fornicabitur in fornicatione sua etiam haec.
EZEK|23|44|Et ingressi sunt ad eam quasi ad mulierem meretricem; sic ingrediebantur ad Oollam et ad Oolibam, mulieres nefarias.
EZEK|23|45|Viri ergo iusti sunt; hi iudicabunt eas iudicio adulterarum et iudicio effundentium sanguinem, quia adulterae sunt, et sanguis in manibus earum.
EZEK|23|46|Haec enim dicit Dominus Deus: " Adduc ad eas congregationem et trade eas in terrorem et in rapinam;
EZEK|23|47|et lapidentur lapidibus congregationis et confodiantur gladiis eorum; filios et filias earum interficiant et domos earum igne succendant.
EZEK|23|48|Et auferam scelus de terra, et discent omnes mulieres, ne faciant secundum scelus vestrum;
EZEK|23|49|et dabunt scelus vestrum super vos, et peccata idolorum vestrorum portabitis et scietis quia ego Dominus Deus ".
EZEK|24|1|Et factum est verbum Do mini ad me in anno nono, in mense decimo, decima mensis, dicens:
EZEK|24|2|"Fili hominis, scribe tibi nomen diei huius, in qua aggressus est rex Babylonis adversum Ierusalem hodie.
EZEK|24|3|Et dices per proverbium ad domum irritatricem parabolam et loqueris ad eos: Haec dicit Dominus Deus:Pone ollam; pone, inquam,et mitte in ea aquam.
EZEK|24|4|Congere frusta eius in ea,omnem partem bonam, femur et armum,electis ossibus imple eam,
EZEK|24|5|pinguissimum pecus assume.Compone quoque struem lignorum sub ea;effervescant frusta eius,et coque ossa illius in medio eius.
EZEK|24|6|Propterea haec dicit Dominus Deus:Vae civitati sanguinum,ollae, cuius rubigo in ea est,et rubigo eius non exivit de ea!Per partes et per partes suas eice ex ea,neque cadat super eam sors.
EZEK|24|7|Sanguis enim eius in medio eius est,super limpidissimam petram effudit illum;non effudit illum super terram,ut possit operiri pulvere;
EZEK|24|8|ut superducerem indignationem meamet vindicta ulciscerer,dedi sanguinem eiussuper petram limpidissimam, ne operiretur.
EZEK|24|9|Propterea haec dicit Dominus Deus:Vae civitati sanguinum,cuius ego grandem faciam pyram!
EZEK|24|10|Congere ligna, succende ignem,coque carnes usque ad consumptionemet effunde ius,et ossa comburentur.
EZEK|24|11|Relinque quoque eam super prunas vacuam,ut incalescat, et ardescat aes eius,et confletur in medio eius inquinamentum eius,et consumatur rubigo eius.
EZEK|24|12|Multo labore sudatum est,et non exibit de ea nimia rubigo eius,neque per ignem.
EZEK|24|13|Immunditia tua execrabilis, quia mundare te volui, et non es mundata a sordibus tuis; sed nec mundaberis prius, donec quiescere faciam indignationem meam in te.
EZEK|24|14|Ego Dominus locutus sum; veniet et faciam: non indulgebo nec parcam nec placabor. Iuxta vias tuas et iuxta opera tua iudicabo te ", dicit Dominus.
EZEK|24|15|Et factum est verbum Domini ad me dicens:
EZEK|24|16|" Fili hominis, ecce ego tollo a te delicias oculorum tuorum in plaga, et non planges neque plorabis, neque fluent lacrimae tuae.
EZEK|24|17|Ingemisce tacens, mortuorum luctum non facies, corona tua circumligata sit tibi, et calceamenta tua pones in pedibus tuis nec amictu ora velabis nec cibos lugentium comedes ".
EZEK|24|18|Locutus sum ergo ad populum mane, et mortua est uxor mea vespere; fecique mane, sicut praeceperat mihi.
EZEK|24|19|Et dixit ad me populus: " Quare non indicas nobis, quid ista significent, quae tu facis? ".
EZEK|24|20|Et dixi ad eos: " Sermo Domini factus est ad me dicens:
EZEK|24|21|Loquere domui Israel: Haec dicit Dominus Deus: Ecce ego polluam sanctuarium meum, superbiam roboris vestri et delicias oculorum vestrorum et sollicitudinem animae vestrae. Filii vestri et filiae, quas reliquistis, gladio cadent.
EZEK|24|22|Et facietis, sicut feci: ora amictu non velabitis et cibos lugentium non comedetis,
EZEK|24|23|coronas habebitis in capitibus vestris et calceamenta in pedibus, non plangetis neque flebitis, sed tabescetis in iniquitatibus vestris, et unusquisque gemet ad fratrem suum.
EZEK|24|24|Eritque Ezechiel vobis in portentum: iuxta omnia, quae fecit, facietis, cum venerit istud, et scietis quia ego Dominus Deus.
EZEK|24|25|Et tu, fili hominis, ecce in die, quo tollam ab eis fortitudinem eorum et gaudium magnificentiae et delicias oculorum eorum et desiderium animae eorum, filios et filias eorum;
EZEK|24|26|in die illa, cum venerit fugiens ad te, ut annuntiet tibi,
EZEK|24|27|in die, inquam, illa aperietur os tuum cum eo, qui fugit; et loqueris et non silebis ultra erisque eis in portentum, et scient quia ego Dominus.
EZEK|25|1|Et factus est sermo Domini ad me dicens:
EZEK|25|2|" Fili hominis, pone faciem tuam contra filios Ammon et propheta de eis
EZEK|25|3|et dices filiis Ammon: Audite verbum Domini Dei.Haec dicit Dominus Deus: Pro eo quod dixisti: "Euge!" super sanctuarium meum, quia pollutum est, et super terram Israel, quoniam desolata est, et super domum Iudae, quoniam ducti sunt in captivitatem,
EZEK|25|4|idcirco ego tradam te filiis orientalibus in hereditatem, et collocabunt castra sua in te et ponent in te tentoria sua; ipsi comedent fruges tuas, et ipsi bibent lac tuum.
EZEK|25|5|Daboque Rabba in pascua camelorum et filios Ammon in cubile pecorum, et scietis quia ego Dominus.
EZEK|25|6|Quia haec dicit Dominus Deus: Pro eo quod plausisti manu et percussisti pede et gavisa es ex toto affectu super terram Israel,
EZEK|25|7|idcirco ecce ego extendam manum meam super te et tradam te in direptionem gentium et interficiam te de populis et perdam de terris et conteram, et scies quia ego Dominus.
EZEK|25|8|Haec dicit Dominus Deus: Pro eo quod dixerunt Moab et Seir: "Ecce sicut omnes gentes domus Iudae!",
EZEK|25|9|idcirco ecce ego aperiam latus Moab privans eam civitatibus, civitatibus, inquam, eius, a finibus eius, decore terrae: Bethiesimoth et Baalmeon et Cariathaim;
EZEK|25|10|filiis orientis cum filiis Ammon dabo eam in hereditatem, ut non sit memoria ultra filiorum Ammon in gentibus.
EZEK|25|11|Et in Moab faciam iudicia, et scient quia ego Dominus.
EZEK|25|12|Haec dicit Dominus Deus: Pro eo quod fecit Idumaea ultionem, ut se vindicaret de domo Iudae, peccavitque delinquens et vindictam expetivit de eis,
EZEK|25|13|idcirco haec dicit Dominus Deus: Extendam manum meam super Idumaeam et auferam de ea hominem et iumentum et faciam eam desertum; de Theman et usque Dedan gladio cadent.
EZEK|25|14|Et dabo ultionem meam super Idumaeam per manum populi mei Israel, et facient in Edom iuxta iram meam et furorem meum, et scient vindictam meam, dicit Dominus Deus.
EZEK|25|15|Haec dicit Dominus Deus: Pro eo quod fecerunt Palaestini in vindicta et ulti se sunt toto animo interficientes et implentes inimicitias sempiternas,
EZEK|25|16|propterea haec dicit Dominus Deus: Ecce ego extendam manum meam super Palaestinos et interficiam Cherethaeos et perdam reliquias maritimae regionis;
EZEK|25|17|faciamque in eis ultiones magnas, arguens in furore, et scient quia ego Dominus, cum dedero vindictam meam super eos ".
EZEK|26|1|Et factum est in undecimo anno, prima mensis, factus est sermo Domini ad me dicens:
EZEK|26|2|"Fili hominis, pro eo quod dixit Tyrus de Ierusalem:Euge, confracta estporta populorum!Conversa est ad me;quae erat plena, deserta est",
EZEK|26|3|propterea haec dicit Dominus Deus:Ecce ego super te, Tyre,et ascendere faciam ad te gentes multas,sicut ascendit mare fluctuans;
EZEK|26|4|et dissipabunt muros Tyriet destruent turres eius,et radam pulverem eius de ea,et dabo eam in limpidissimam petram.
EZEK|26|5|Siccatio sagenarumerit in medio maris,quia ego locutus sum,ait Dominus Deus;et erit in direptionem gentibus.
EZEK|26|6|Filiae quoque eius, quae sunt in agro,gladio interficientur,et scient quia ego Dominus.
EZEK|26|7|Quia haec dicit Dominus Deus:Ecce ego adducam ad TyrumNabuchodonosor, regem Babylonis,ab aquilone, regem regum,cum equis et curribus et equitibuset coetu populoque magno.
EZEK|26|8|Filias tuas, quae sunt in agro,gladio interficiet,et circumdabit te munitionibuset comportabit aggerem in gyroet levabit contra te clipeum
EZEK|26|9|et vineas et arietes temperabit in muros tuoset turres tuas destruet in armatura sua.
EZEK|26|10|Inundatione equorum eiusoperiet te pulvis eorum,a sonitu equitumet rotarum et curruummovebuntur muri tui,dum ingressus fuerit portas tuasquasi per introitus urbis dissipatae.
EZEK|26|11|Ungulis equorum suorumconculcabit omnes plateas tuas,populum tuum gladio caedet,et columnae tuae fortissimaein terram corruent.
EZEK|26|12|Vastabunt opes tuas,diripient negotiationes tuaset destruent muros tuoset domos tuas praeclaras subvertentet lapides tuos et ligna tua et pulverem tuumin medio aquarum ponent.
EZEK|26|13|Et quiescere faciam tumultum canticorum tuorum,et sonitus cithararum tuarum non audietur amplius,
EZEK|26|14|et dabo te in limpidissimam petram;siccatio sagenarum eris,nec aedificaberis ultra,quia ego locutus sum,dicit Dominus Deus.
EZEK|26|15|Haec dicit Dominus Deus Tyro: Numquid non a sonitu ruinae tuae et gemitu interfectorum tuorum, cum occisi fuerint in medio tui, commovebuntur insulae?
EZEK|26|16|Et descendent de sedibus suis omnes principes maris et auferent pallia sua et vestimenta sua varia abicient; et induentur stupore, in terra sedebunt et attoniti et tremefacti stupebunt super te.
EZEK|26|17|Et assumentes super te lamentum dicent tibi:Quomodo peristi, quae habitas in mari,urbs inclita,quae fuisti fortis in maricum habitatoribus tuis,quos formidabant universi!
EZEK|26|18|Nunc stupebunt navesin die ruinae tuae,et turbabuntur insulae in mariob exitum tuum".
EZEK|26|19|Quia haec dicit Dominus Deus: Cum dedero te urbem desolatam sicut civitates, quae non habitantur, et adduxero super te abyssum, et operuerint te aquae multae,
EZEK|26|20|detraham te cum his, qui descendunt in lacum, ad populum pristinum et collocabo te in profundis terrae sicut ruinas a saeculo cum his, qui descendunt in lacum, ut non habiteris et consistas in terra viventium;
EZEK|26|21|in nihilum redigam te, et non eris et requisita non invenieris ultra in sempiternum ", dicit Dominus Deus.
EZEK|27|1|Et factum est verbum Do mini ad me dicens:
EZEK|27|2|"Tu er go, fili hominis, assume super Tyrum lamentum
EZEK|27|3|et dices Tyro, quae habitat in introitu maris, negotiatrici populorum ad insulas multas: Haec dicit Dominus Deus:O Tyre, tu dixisti: "Perfecti decoris ego sum!".
EZEK|27|4|In corde maris fines tui;qui te aedificaverunt, impleverunt decorem tuum.
EZEK|27|5|Abietibus de Sanir exstruxerunttibi omnia tabulata;cedrum de libano tulerunt,ut facerent tibi malum;
EZEK|27|6|quercus de Basandolaverunt in remos tuoset transtra tua fecerunt ex eboreet cupressis de insulis Cetthim.
EZEK|27|7|Byssus varia texta de Aegyptoerat tibi in velum,ut poneretur in malo,hyacinthus et purpura de insulis Elisafacta sunt operimentum tuum.
EZEK|27|8|Habitatores Sidonis et Aradiifuerunt remiges tui;sapientes tui, Tyre,facti sunt nautae tui.
EZEK|27|9|Senes Gibli et prudentes eius fuerunt in te,ut sarcirent rimas tuas.Omnes naves maris et nautae earumfuerunt in te, ut mercarentur merces tuas.
EZEK|27|10|Persae et Lud et Phuterant in exercitu tuo,viri bellatores tui.Clipeum et galeam suspenderunt in te;ipsi dederunt tibi splendorem.
EZEK|27|11|Filii Aradii cum exercitu tuo erant super muros tuos in circuitu, et Gammadii erant in turribus tuis. Clipeos suos suspenderunt in muris tuis per gyrum; ipsi compleverunt pulchritudinem tuam.
EZEK|27|12|Tharsis negotiatrix tua propter multitudinem cunctarum divitiarum; argentum, ferrum, stannum plumbumque dederunt pro mercibus tuis.
EZEK|27|13|Iavan, Thubal et Mosoch ipsi institores tui; mancipia et vasa aerea adduxerunt tibi in commutationem populo tuo.
EZEK|27|14|De domo Thogorma equos et equites et mulos adduxerunt pro mercibus tuis ad forum tuum;
EZEK|27|15|filii Rhodi negotiatores tui; insulae multae negotiatio manus tuae: dentes eburneos et ebenina reddiderunt tibi ut tributum.
EZEK|27|16|Edom negotiator tuus propter multitudinem operum tuorum; carbunculum, purpuram et scutulata et byssum et corallia et rubinum attulerunt pro mercibus tuis.
EZEK|27|17|Iuda et terra Israel ipsi institores tui; frumentum primum, balsamum et mel et oleum et resinam attulerunt tibi in commutationem.
EZEK|27|18|Damascenus negotiator tuus propter multitudinem operum tuorum, propter multitudinem diversarum opum; vinum de Helbon et lanam de Sahar
EZEK|27|19|et vinum de Uzal pro mercibus tuis dederunt; ferrum fabrefactum, cassia et calamus in commutatione tua erat.
EZEK|27|20|Dedan institores tui in tapetibus ad equitandum.
EZEK|27|21|Arabia et universi principes Cedar ipsi negotiatores manus tuae; cum agnis et arietibus et haedis, cum quibus erant negotiatores tui.
EZEK|27|22|Venditores Saba et Regma, ipsi negotiatores tui, universa prima aromata et omnem lapidem pretiosum et aurum dederunt pro mercibus tuis.
EZEK|27|23|Charran et Chenne et Eden negotiatores tui; Saba, Assyria et Chelmad venditores tui.
EZEK|27|24|Ipsi negotiatores tui cum vestibus splendidis, involucris hyacinthinis et polymitis texturisque discoloribus, funibus obvolutis et cedris in negotiationibus tuis.
EZEK|27|25|Naves Tharsis, principes tuiin negotiatione tua;et repleta es et glorificata nimisin corde maris.
EZEK|27|26|In aquis multis adduxerunt teremiges tui;ventus auster contrivit tein corde maris.
EZEK|27|27|Divitiae tuae et thesauri tui et multiplices merces tuae,nautae tui et gubernatores tui,resarcientes rimas tuas et commutantes merces tuas,omnes quoque viri bellatores tui,qui sunt in te,cum universa multitudine tua,quae est in medio tui,cadent in corde marisin die ruinae tuae.
EZEK|27|28|A sonitu clamoris gubernatorum tuorumconturbabuntur litora.
EZEK|27|29|Et descendent de navibus suisomnes, qui tenebant remum;nautae et universi gubernatores marisin terra stabunt.
EZEK|27|30|Et eiulabunt super te voce magnaet clamabunt amare;et superiacient pulverem capitibus suis,in cinere volutabuntur.
EZEK|27|31|Et radent super te calvitiumet accingentur ciliciiset plorabunt te in amaritudine animaeploratu amarissimo;
EZEK|27|32|et assument super te congementes carmen lugubreet plangent te:Quae est ut Tyrus, quae obmutuitin medio maris?
EZEK|27|33|Cum venissent merces tuae de mari, satiasti populos multos;in multitudine divitiarum tuarum et mercium tuarumditasti reges terrae.
EZEK|27|34|Nunc contrita es a mariin profundis aquarum.Opes tuae et omnis multitudo tua,quae erat in medio tui,ceciderunt.
EZEK|27|35|Universi habitatores insularumobstupuerunt super te,et reges earum horrore formidarunt vultu conturbato;
EZEK|27|36|negotiatores in populis sibilaverunt super te.In horrorem facta eset non eris usque in perpetuum" ".
EZEK|28|1|Et factus est sermo Domini ad me dicens:
EZEK|28|2|" Fili hominis, dic principi Tyri: Haec dicit Dominus Deus:Eo quod elevatum est cor tuum,et dixisti: "Deus ego sumet in cathedra deorum sedeoin corde maris!",cum sis homo et non Deus,et dedisti cor tuum quasi cor Dei.
EZEK|28|3|Ecce sapientior es tu Danel,omne secretum non est absconditum a te,
EZEK|28|4|in sapientia et prudentia tuafecisti tibi opeset acquisisti aurum et argentumin thesauris tuis;
EZEK|28|5|in multitudine sapientiae tuae et in negotiatione tuamultiplicasti tibi opes,et elevatum est cor tuum in opibus tuis.
EZEK|28|6|Propterea haec dicit Dominus Deus: Eo quod fecisti cor tuum quasi cor Dei,
EZEK|28|7|idcirco ecce ego adducam super tealienos violentissimos gentium;et nudabunt gladios suos super pulchritudinem sapientiae tuaeet polluent splendorem tuum.
EZEK|28|8|In fossam detrahent te, et morierisinteritu occisorum in corde maris.
EZEK|28|9|Numquid dicens loqueris: "Deus ego sum!"coram interficientibus te,cum sis homo et non Deusin manu occidentium te?
EZEK|28|10|Morte incircumcisorum morierisin manu alienorum,quia ego locutus sum ",ait Dominus Deus.
EZEK|28|11|Et factus est sermo Domini ad me dicens: " Fili hominis, leva planctum super regem Tyri
EZEK|28|12|et dices ei: Haec dicit Dominus Deus:Tu signaculum perfectum,plenus sapientia et perfectus decore;
EZEK|28|13|in deliciis paradisi Dei fuisti,omnis lapis pretiosus operimentum tuum:sardius, topazius et iaspis,chrysolithus et onyx et beryllus,sapphirus et carbunculus et smaragdus,aurum opus caelaturae in te;in die, qua conditus es, praeparata sunt.
EZEK|28|14|Cum cherub extento et protegente te posui te,in monte sancto Dei fuisti,in medio lapidum ignitorum ambulasti,
EZEK|28|15|perfectus in viis tuisa die conditionis tuae,donec inventa est iniquitas in te.
EZEK|28|16|In multitudine negotiationis tuae repleta sunt interiora tuainiquitate, et peccasti.Et eieci te de monte Dei,et perdidit te cherub protegensde medio lapidum ignitorum.
EZEK|28|17|Elevatum est cor tuum in decore tuo;perdidisti sapientiam tuam propter splendorem tuum:in terram proieci te,ante faciem regum dedi te, ut cernerent te.
EZEK|28|18|In multitudine iniquitatum tuarumet iniquitate negotiationis tuaepolluisti sanctuaria tua;producam ergo ignem de medio tui,qui comedat te,et dabo te in cinerem super terramin conspectu omnium videntium te.
EZEK|28|19|Omnes, qui viderint te, in gentibusobstupescent super te;in horrorem factus eset non eris in perpetuum ".
EZEK|28|20|Et factus est sermo Domini ad me dicens:
EZEK|28|21|" Fili hominis, pone faciem tuam contra Sidonem et propheta de ea
EZEK|28|22|et dices: Haec dicit Dominus Deus:Ecce ego ad te, Sidon,et glorificabor in medio tui,et scient quia ego Dominus,cum fecero in ea iudiciaet sanctificatus fuero in ea.
EZEK|28|23|Et immittam ei pestilentiamet sanguinem in plateis eius,et corruent interfecti in medio eius gladio per circuitum,et scient quia ego Dominus.
EZEK|28|24|Et non erit ultra domui Israel stimulus amaritudinis et spina dolorem inferens undique per circuitum eorum, qui adversantur eis, et scient quia ego Dominus Deus.
EZEK|28|25|Haec dicit Dominus Deus: Quando congregavero domum Israel de populis, in quibus dispersi sunt, sanctificabor in eis coram gentibus, et habitabunt in terra sua, quam dedi servo meo Iacob;
EZEK|28|26|et habitabunt in ea securi et aedificabunt domos plantabuntque vineas et habitabunt confidenter, cum fecero iudicia in omnibus, qui adversantur eis per circuitum, et scient quia ego Dominus Deus eorum ".
EZEK|29|1|In anno decimo, in decimo mense, duodecima mensis, factum est verbum Domini ad me dicens:
EZEK|29|2|" Fili hominis, pone faciem tuam contra pharaonem, regem Aegypti, et prophetabis de eo et de Aegypto universa.
EZEK|29|3|Loquere et dices: Haec dicit Dominus Deus:Ecce ego ad te, pharao,rex Aegypti,draco magne, qui cubasin medio fluminum tuorumet dicis: "Meus est fluvius,et ego feci memetipsum!".
EZEK|29|4|Et ponam uncos in maxillis tuiset agglutinabo pisces fluminum tuorum squamis tuiset extraham te de medio fluminum tuorum,et universi pisces tui squamis tuis adhaerebunt.
EZEK|29|5|Et proiciam te in desertumet omnes pisces fluminum tuorum.Super faciem terrae cades;non colligeris neque congregaberis.Bestiis terrae et volatilibus caelidedi te ad devorandum.
EZEK|29|6|Et scient omnes habitatores Aegyptiquia ego Dominus,pro eo quod fuisti baculus arundineusdomui Israel:
EZEK|29|7|quando apprehenderunt te manu,confractus es et lacerasti omnem umerum eorumet, innitentibus eis super te,comminutus eset dissolvisti omnes lumbos eorum.
EZEK|29|8|Propterea haec dicit Dominus Deus: Ecce ego adducam super te gladium et interficiam de te hominem et iumentum;
EZEK|29|9|et erit terra Aegypti in desertum et solitudinem, et scient quia ego Dominus. Pro eo quod dixeris: "Fluvius meus est, et ego feci!",
EZEK|29|10|idcirco ecce ego ad te et ad flumina tua, daboque terram Aegypti in solitudines, gladio dissipatam a Magdolo ad Syenen et usque ad terminos Chus.
EZEK|29|11|Non pertransibit eam pes hominis, neque pes iumenti gradietur in ea, et non habitabitur quadraginta annis;
EZEK|29|12|daboque terram Aegypti desertam in medio terrarum desertarum, et civitates eius in medio urbium subversarum erunt desolatae quadraginta annis, et dispergam Aegyptios in nationes et ventilabo eos in terras.
EZEK|29|13|Quia haec dicit Dominus Deus: Post finem quadraginta annorum congregabo Aegyptios de populis, in quibus dispersi fuerunt,
EZEK|29|14|et convertam sortem Aegypti et collocabo eos in terra Phatures, in terra nativitatis suae; et erunt ibi in regnum humile.
EZEK|29|15|Inter regna cetera erit humillima et non elevabitur ultra super nationes, et imminuam eos, ne imperent gentibus.
EZEK|29|16|Neque erunt ultra domui Israel in confidentiam, in memoriam revocans iniquitatem, cum sequerentur eos, et scient quia ego Dominus Deus ".
EZEK|29|17|Et factum est in vicesimo et septimo anno, in primo, in una mensis, factum est verbum Domini ad me dicens:
EZEK|29|18|" Fili hominis, Nabuchodonosor, rex Babylonis, servire fecit exercitum suum servitute magna adversus Tyrum; omne caput decalvatum et omnis umerus attritus est, et merces non est reddita ei neque exercitui eius de Tyro pro servitute, qua servivit adversum eam.
EZEK|29|19|Propterea haec dicit Dominus Deus: Ecce ego dabo Nabuchodonosor, regi Babylonis, terram Aegypti, et accipiet opes eius et depraedabitur manubias eius et diripiet spolia eius, et erit merces exercitui illius,
EZEK|29|20|ut stipendium eius, pro quo servivit adversum eam. Dedi ei terram Aegypti pro eo quod laboraverunt mihi, ait Dominus Deus.
EZEK|29|21|In die illo germinare faciam cornu domui Israel, et tibi dabo apertum os in medio eorum, et scient quoniam ego Dominus ".
EZEK|30|1|Et factum est verbum Do mini ad me dicens:
EZEK|30|2|" Fili ho minis, propheta et dic: Haec dicit Dominus Deus:Ululate, vae diei,
EZEK|30|3|quia iuxta est dies,et appropinquat dies Domini,dies nubis; tempus gentium erit.
EZEK|30|4|Et veniet gladius in Aegyptum,et erit pavor in Chus,cum ceciderint vulnerati in Aegypto,et ablatae fuerint opes illius,et destructa fundamenta eius.
EZEK|30|5|Chus et Phut et Lud et omne vulgus promiscuumet Chub et filii terrae foederiscum eis gladio cadent.
EZEK|30|6|Haec dicit Dominus Deus:Et corruent fulcientes Aegyptum,et destruetur superbia potentiae eius;a Magdolo usque ad Syenen gladio cadent in ea,ait Dominus Deus.
EZEK|30|7|Et dissipabuntur in medio terrarum desolatarum, et urbes eius in medio civitatum desertarum erunt;
EZEK|30|8|et scient quia ego Dominus, cum dedero ignem in Aegyptum, et attriti fuerint omnes auxiliatores eius.
EZEK|30|9|In die illa egredientur nuntii a facie mea in navibus ad conterendam confidentiam Chus, et erit pavor in eis in die Aegypti, quia veniet.
EZEK|30|10|Haec dicit Dominus Deus: Cessare faciam pompam Aegypti in manu Nabuchodonosor, regis Babylonis.
EZEK|30|11|Ipse et populus eius cum eo violentissimi gentium adducentur ad disperdendam terram; et evaginabunt gladios suos super Aegyptum et implebunt terram interfectis.
EZEK|30|12|Et faciam alveos fluminum aridos et tradam terram in manu pessimorum et dissipabo terram et plenitudinem eius in manu alienorum. Ego Dominus locutus sum.
EZEK|30|13|Haec dicit Dominus Deus:Et disperdam simulacraet cessare faciam idola de Memphi,et dux de terra Aegyptinon erit amplius,et dabo terrorem in terra Aegypti.
EZEK|30|14|Et disperdam terram Phatureset dabo ignem in Taniet faciam iudicia in No.
EZEK|30|15|Et effundam indignationem meam super Sin, robur Aegypti, et interficiam multitudinem No.
EZEK|30|16|Et dabo ignem in Aegypto; quasi parturiens dolebit Sin, et in No scissura erit, et contra Memphin hostes plena die.
EZEK|30|17|Iuvenes Heliopoleos et Bubasti gladio cadent, et ipsae captivae ducentur.
EZEK|30|18|Et in Taphnis nigrescet dies, cum contrivero ibi sceptra Aegypti, et defecerit in ea superbia potentiae eius; ipsam nubes operiet, filiae autem eius in captivitatem ducentur.
EZEK|30|19|Et faciam iudicia in Aegypto, et scient quia ego Dominus ".
EZEK|30|20|Et factum est in undecimo anno, in primo, in septima mensis, factum est verbum Domini ad me dicens:
EZEK|30|21|" Fili hominis, brachium pharaonis, regis Aegypti, confregi, et ecce non est obvolutum, ut restitueretur ei sanitas, ut ligaretur pannis et farciretur linteolis, ut recepto robore posset tenere gladium.
EZEK|30|22|Propterea haec dicit Dominus Deus: Ecce ego ad pharaonem, regem Aegypti, et comminuam brachium eius forte sed confractum et deiciam gladium de manu eius
EZEK|30|23|et dispergam Aegyptum in gentibus et ventilabo eos in terris.
EZEK|30|24|Et confortabo brachia regis Babylonis daboque gladium meum in manu eius; et confringam brachia pharaonis, et gemet gemitibus sicut transfixus coram facie eius.
EZEK|30|25|Et confortabo brachia regis Babylonis, et brachia pharaonis concident; et scient quia ego Dominus, cum dedero gladium meum in manu regis Babylonis, et extenderit eum super terram Aegypti.
EZEK|30|26|Et dispergam Aegyptum in nationes et ventilabo eos in terras, et scient quia ego Dominus ".
EZEK|31|1|Et factum est in anno unde cimo, in tertio, una mensis, factum est verbum Domini ad me dicens:
EZEK|31|2|" Fili hominis, dic pharaoni, regi Aegypti, et pompae eius:Cui similis factus es in magnitudine tua?
EZEK|31|3|Ecce abies, quasi cedrus in Libano,pulcher ramis et frondibus nemorosusexcelsusque altitudine,et inter nubes elevatum est cacumen eius;
EZEK|31|4|aquae nutrierunt illum,abyssus exaltavit eum,flumina eius manabantin circuitu radicum eius,et rivos suos emisitad universa ligna campi.
EZEK|31|5|Propterea elevata est altitudo eiussuper omnia ligna campi,et multiplicata sunt arbusta eius,et elevati sunt rami eiuspropter aquas multas.
EZEK|31|6|Cumque extendisset umbram suam,in ramis eius fecerunt nidosomnia volatilia caeli,et sub frondibus eius genueruntomnes bestiae campi,et sub umbra illius habitabatuniversa multitudo gentium;
EZEK|31|7|eratque pulcherrimus in magnitudine suaet in dilatatione arbustorum suorum,erat enim radix illiusiuxta aquas multas.
EZEK|31|8|Cedri non fuerunt pares illiin paradiso Dei;abietes non adaequaveruntramos eius,et platani non fueruntaequae frondibus illius;omne lignum paradisi Deinon est assimilatum illi et pulchritudini eius,
EZEK|31|9|quoniam speciosum feci eumet multis condensisque frondibus:et aemulata sunt eum omnia ligna Eden,quae erant in paradiso Dei.
EZEK|31|10|Propterea haec dicit Dominus Deus: Pro eo quod sublimatus est in altitudine et dedit summitatem suam usque in nubes, et elevatum est cor eius in altitudine sua,
EZEK|31|11|tradam eum in manu potentis principis gentium; faciens faciet ei: iuxta impietatem eius eieci eum.
EZEK|31|12|Et succident illum alieni, violentissimi nationum; et proicient eum super montes, et in cunctis convallibus corruent rami eius, et confringentur arbusta eius in universis voraginibus terrae, et recedent de umbra eius omnes populi terrae et relinquent eum.
EZEK|31|13|Super ruinam eius habitabuntomnia volatilia caeli,et in ramis eius eruntuniversae bestiae campi,
EZEK|31|14|ne eleventur in altitudine suaomnia ligna aquarum neque ponantsublimitatem suam inter nubes necstent apud eas in sublimitate suaomnia, quae irrigantur aquis, quiaomnes traditi sunt in mortemad inferiora terrae,in medio filiorum hominum,ad eos, qui descendunt in lacum.
EZEK|31|15|Haec dicit Dominus Deus: In die, quando descendit ad inferos, induxi luctum, operui propter eum abyssum et prohibui flumina eius et coercui aquas multas; obscuravi super eum Libanum, et omnia ligna agri concussa sunt.
EZEK|31|16|A sonitu ruinae eius commovi gentes, cum deducerem eum ad infernum cum his, qui descendebant in lacum; et consolata sunt in inferioribus terrae omnia ligna Eden, egregia atque praeclara in Libano, universa, quae irrigabantur aquis.
EZEK|31|17|Nam et ipsi cum eo descenderunt ad infernum ad interfectos gladio et auxiliatores eius, qui sederant sub umbra eius in medio nationum.
EZEK|31|18|Cui assimilatus es, o inclite atque sublimis inter ligna Eden? Et ecce deductus es cum lignis Eden ad inferiora terrae; in medio incircumcisorum dormies cum his, qui interfecti sunt gladio. Ipse est pharao et omnis pompa eius ", dicit Dominus Deus.
EZEK|32|1|Et factum est duodecimo anno, in mense duodecimo, in una mensis, factum est verbum Domini ad me dicens:
EZEK|32|2|" Fili hominis, assume lamentum super pharaonem, regem Aegypti, et dices ad eum:Leo gentium peristi,et eras sicut draco in mari;et bulliebas in fluminibus tuiset conturbabas aquas pedibus tuiset turbida faciebas flumina earum.
EZEK|32|3|Haec dicit Dominus Deus:Expandam super te rete meumin coetu populorum multorum,et extrahent te in sagena mea;
EZEK|32|4|et proiciam te in terram,super faciem agri abiciam teet habitare faciam super te omnia volatilia caeliet saturabo de te bestias universae terrae;
EZEK|32|5|et dabo carnes tuas super monteset implebo valles sanie tua.
EZEK|32|6|Et irrigabo terram paedoresanguinis tui super montes,et voragines implebuntur ex te;
EZEK|32|7|et operiam, cum exstinctus fueris, caelumet nigrescere faciam stellas eius:solem nube tegam,et luna non dabit lumen suum;
EZEK|32|8|omnia luminaria caelimaerere faciam super teet dabo tenebras super terram tuam,dicit Dominus Deus.
EZEK|32|9|Et commovebo cor populorum multorum, cum induxero contritionem tuam in gentibus super terras, quas nescis.
EZEK|32|10|Et stupescere faciam super te populos multos, et reges eorum horrore nimio formidabunt super te, cum volare coeperit gladius meus coram facie eorum, et obstupescet tremefactus unusquisque pro anima sua in die ruinae tuae.
EZEK|32|11|Quia haec dicit Dominus Deus: Gladius regis Babylonis veniet tibi,
EZEK|32|12|in gladiis fortium deiciam multitudinem tuam;violentissimae gentium omnium haeet vastabunt superbiam Aegypti,et dissipabitur omnis pompa eius.
EZEK|32|13|Et perdam omnia iumenta eius,quae erant super aquas plurimas,et non conturbabit eas pes hominis ultra,neque ungula iumentorum turbabit eas;
EZEK|32|14|tunc purissimas reddam aquas eorumet flumina eorum quasi oleum adducam,ait Dominus Deus.
EZEK|32|15|Cum dedero terram Aegypti desolatam,deseretur autem terra a plenitudine sua, quando percussero omnes habitatores eius,scient quia ego Dominus.
EZEK|32|16|Planctus est, et plangent eum; filiae gentium plangent eum, super Aegyptum et super omnem pompam eius plangent eum ", ait Dominus Deus.
EZEK|32|17|Et factum est in duodecimo anno, in quinta decima mensis, factum est verbum Domini ad me dicens:
EZEK|32|18|" Fili hominis, cane lugubre super pompam Aegypti et detrahe eam, ipsam et filias gentium robustarum ad inferiora terrae cum his, qui descendunt in lacum.
EZEK|32|19|Quo pulchrior es?Descende et dormi cum incircumcisis.
EZEK|32|20|In medio interfectorum gladio cadent; gladius datus est, attraxerunt eam et omnes populos eius.
EZEK|32|21|Loquentur ei potentissimi robustorum de medio inferni, cum auxiliatoribus eius descenderunt:Tacent incircumcisi interfecti gladio!".
EZEK|32|22|Ibi Assyria et omnis multitudo eius, in circuitu illius sepulcra eius, omnes interfecti, qui ceciderunt gladio;
EZEK|32|23|quorum data sunt sepulcra in profundissimis laci, et facta est multitudo eius per gyrum sepulcri eius; universi interfecti, cadentes gladio, qui dederant quondam formidinem in terra viventium.
EZEK|32|24|Ibi Elam et omnis pompa eius per gyrum sepulcri sui; omnes hi interfecti ruentesque gladio, qui descenderunt incircumcisi ad inferiora terrae, qui dederant quondam formidinem suam in terra viventium et sustulerunt ignominiam suam cum his, qui descendunt in lacum.
EZEK|32|25|In medio interfectorum posuerunt cubile eius, in omni pompa eius, in circuitu eius sepulcra illius, omnes hi incircumcisi interfectique gladio; dederant enim terrorem suum in terra viventium et sustulerunt ignominiam suam cum his, qui descendunt in lacum, in medio interfectorum positi sunt.
EZEK|32|26|Ibi Mosoch, Thubal et omnis pompa eius, in circuitu illius sepulcra eius, omnes hi incircumcisi interfectique gladio, quia dederunt formidinem suam in terra viventium;
EZEK|32|27|et non dormient cum fortibus, qui ceciderunt a saeculo et descenderunt ad infernum cum armis suis et posuerunt gladios suos sub capitibus suis, et fuerunt scuta eorum super ossa eorum, quia terror fortium erat in terra viventium.
EZEK|32|28|Et tu ergo in medio incircumcisorum contereris et dormies cum interfectis gladio.
EZEK|32|29|Ibi Idumaea, reges eius et omnes duces eius, qui dati sunt in robore suo cum interfectis gladio et qui cum incircumcisis dormiunt et cum his, qui descenderunt in lacum.
EZEK|32|30|Ibi principes aquilonis omnes et universi Sidonii, qui deducti sunt cum interfectis in terrore suo, in sua fortitudine confusi; qui dormiunt incircumcisi cum interfectis gladio et sustulerunt confusionem suam cum his, qui descendunt in lacum.
EZEK|32|31|Videbit eos pharao et consolabitur super universa pompa sua. Interfecti sunt gladio pharaonis et omnis exercitus eius, ait Dominus Deus,
EZEK|32|32|quia dedi terrorem meum in terra viventium; et prostratus est in medio incircumcisorum cum interfectis gladio pharaonis et omnis pompa eius ", ait Dominus Deus.
EZEK|33|1|Et factum est verbum Do mini ad me dicens:
EZEK|33|2|" Fili ho minis, loquere ad filios populi tui et dices ad eos: Terra, cum induxero super eam gladium, et tulerit populus terrae virum unum de finibus suis et constituerit eum sibi speculatorem,
EZEK|33|3|et ille viderit gladium venientem super terram et cecinerit bucina et annuntiaverit populo;
EZEK|33|4|audiens autem quisquis ille est sonum bucinae, non se observaverit, veneritque gladius et tulerit eum: sanguis ipsius super caput eius erit;
EZEK|33|5|sonum bucinae audivit et non se observavit, sanguis eius in ipso erit. Si autem se custodierit, animam suam salvavit.
EZEK|33|6|Quod si speculator viderit gladium venientem et non insonuerit bucina, et populus non se custodierit; veneritque gladius et tulerit de eis animam: ille quidem in iniquitate sua captus est, sanguinem autem eius de manu speculatoris requiram.
EZEK|33|7|Te autem, fili hominis, speculatorem dedi domui Israel. Audiens ergo ex ore meo sermonem, commonebis eos ex me.
EZEK|33|8|Si, me dicente ad impium: Impie, morte morieris, non fueris locutus, ut se custodiat impius a via sua, ipse impius in iniquitate sua morietur, sanguinem autem eius de manu tua requiram.
EZEK|33|9|Si autem commonueris impium, ut a viis suis convertatur, et ille non fuerit conversus a via sua, ipse in iniquitate sua morietur, porro tu animam tuam liberasti.
EZEK|33|10|Tu ergo, fili hominis, dic ad domum Israel: Sic locuti estis, dicentes: Iniquitates nostrae et peccata nostra super nos sunt, et in ipsis nos tabescimus; quomodo ergo vivere poterimus?".
EZEK|33|11|Dic ad eos: Vivo ego, dicit Dominus Deus; nolo mortem impii, sed ut revertatur impius a via sua et vivat. Convertimini, convertimini a viis vestris pessimis; et quare moriemini, domus Israel?
EZEK|33|12|Tu itaque, fili hominis, dic ad filios populi tui: Iustitia iusti non liberabit eum in quacumque die praevaricatus fuerit; et impietas impii non nocebit ei in quacumque die conversus fuerit ab impietate sua; et iustus non poterit vivere in iustitia sua in quacumque die peccaverit.
EZEK|33|13|Etiamsi dixero iusto quod vita vivat, et, confisus in iustitia sua, fecerit iniquitatem, omnes iustitiae eius oblivioni tradentur, et in iniquitate sua, quam operatus est, in ipsa morietur.
EZEK|33|14|Sin autem dixero impio: Morte morieris, et egerit paenitentiam a peccato suo feceritque iudicium et iustitiam,
EZEK|33|15|pignus restituerit ille impius rapinamque reddiderit, in mandatis vitae ambulaverit nec fecerit quidquam iniustum, vita vivet et non morietur;
EZEK|33|16|omnia peccata eius, quae peccavit, non imputabuntur ei: iudicium et iustitiam fecit, vita vivet.
EZEK|33|17|Et dicunt filii populi tui: "Non est aequa via Domini"; et ipsorum via iniqua est.
EZEK|33|18|Cum enim recesserit iustus a iustitia sua feceritque iniquitates, morietur in eis;
EZEK|33|19|et cum recesserit impius ab impietate sua feceritque iudicium et iustitiam, vivet in eis.
EZEK|33|20|Et dicitis: "Non est recta via Domini". Unumquemque iuxta vias suas iudicabo de vobis, domus Israel ".
EZEK|33|21|Et factum est in duodecimo anno, in decimo, in quinta mensis transmigrationis nostrae, venit ad me, qui fugerat de Ierusalem, dicens: " Vastata est civitas ".
EZEK|33|22|Manus autem Domini facta fuerat ad me vespere, antequam veniret qui fugerat; aperuitque os meum, donec veniret ad me mane, et, aperto ore meo, non silui amplius.
EZEK|33|23|Et factum est verbum Domini ad me dicens:
EZEK|33|24|" Fili hominis, qui habitant in ruinosis his super humum Israel, loquentes aiunt: "Unus erat Abraham et hereditate possedit terram; nos autem multi, nobis data est terra in possessionem".
EZEK|33|25|Idcirco dices ad eos: Haec dicit Dominus Deus: Qui in sanguine comeditis et oculos vestros levatis ad idola vestra et sanguinem funditis, numquid terram hereditate possidebitis?
EZEK|33|26|Stetistis in gladiis vestris, fecistis abominationes, et unusquisque uxorem proximi sui polluit, et terram hereditate possidebitis?
EZEK|33|27|Haec dices ad eos: Sic dicit Dominus Deus: Vivo ego, qui in ruinosis habitant, gladio cadent; et, qui in agro est, bestiis tradetur ad devorandum; qui autem in praesidiis et in speluncis sunt, peste morientur.
EZEK|33|28|Et dabo terram in solitudinem et desertum, et deficiet superba fortitudo eius, et desolabuntur montes Israel, ita ut nullus sit qui per eos transeat;
EZEK|33|29|et scient quia ego Dominus, cum dedero terram desolatam et desertam propter universas abominationes suas, quas operati sunt.
EZEK|33|30|Et tu, fili hominis, filii populi tui, qui loquuntur de te iuxta parietes et in ostiis domorum et dicunt unus ad alterum, vir ad fratrem suum, loquentes: "Venite et audite, qui sit sermo egrediens a Domino".
EZEK|33|31|Et veniunt ad te quasi si conveniat populus, et sedent coram te populus meus; et audiunt sermones tuos et non faciunt eos, quia quasi amatores loquuntur, et avaritiam suam sequitur cor eorum.
EZEK|33|32|Et es eis quasi carmen amatorum, quod suavi voce et cum dulci chordarum sono canitur, et audiunt verba tua et non faciunt ea.
EZEK|33|33|Et cum venerit, quod praedictum est - ecce enim venit - tunc scient quod prophetes fuerit inter eos ".
EZEK|34|1|Et factum est verbum Do mini ad me dicens:
EZEK|34|2|" Fili ho minis, propheta de pastoribus Israel, propheta et dices pastoribus: Haec dicit Dominus Deus: Vae pastoribus Israel, qui pascebant semetipsos! Nonne greges pascuntur a pastoribus?
EZEK|34|3|Lac comedebatis et lana operiebamini et, quod crassum erat, occidebatis, gregem autem non pascebatis;
EZEK|34|4|quod infirmum fuit, non consolidastis et, quod aegrotum, non sanastis; quod fractum est, non alligastis et, quod eiectum est, non reduxistis et, quod perierat, non quaesistis et super forte imperabatis cum violentia.
EZEK|34|5|Et dispersae sunt oves meae, eo quod non esset pastor; et factae sunt in devorationem omnium bestiarum agri et dispersae sunt.
EZEK|34|6|Erraverunt greges mei in cunctis montibus et in universo colle excelso, et super omnem faciem terrae dispersi sunt greges mei; et non erat qui requireret, non erat qui requireret.
EZEK|34|7|Propterea, pastores, audite verbum Domini:
EZEK|34|8|Vivo ego, dicit Dominus Deus, pro eo quod factus est grex meus in rapinam et oves meae in devorationem omnium bestiarum agri, eo quod non esset pastor, neque enim quaesierunt pastores mei gregem meum, sed pascebant pastores semetipsos et gregem meum non pascebant,
EZEK|34|9|propterea, pastores, audite verbum Domini.
EZEK|34|10|Haec dicit Dominus Deus: Ecce ego ipse super pastores requiram gregem meum de manu eorum et cessare eos faciam, ut ultra non pascant gregem nec pascant amplius pastores semetipsos; et liberabo gregem meum de ore eorum, et non erit ultra eis in escam.
EZEK|34|11|Quia haec dicit Dominus Deus: Ecce ego ipse requiram oves meas et visitabo eas.
EZEK|34|12|Sicut visitat pastor gregem suum in die, quando fuerit in medio ovium suarum dissipatarum, sic visitabo oves meas et liberabo eas de omnibus locis, in quibus dispersae fuerant in die nubis et caliginis.
EZEK|34|13|Et educam eas de populis et congregabo eas de terris et inducam eas in terram suam et pascam eas in montibus Israel, in rivis et in cunctis sedibus terrae.
EZEK|34|14|In pascuis uberrimis pascam eas, et in montibus excelsis Israel erunt pascua earum; ibi requiescent in herbis virentibus et in pascuis pinguibus pascentur super montes Israel.
EZEK|34|15|Ego pascam oves meas et ego eas accubare faciam, dicit Dominus Deus.
EZEK|34|16|Quod perierat, requiram et, quod eiectum erat, reducam et, quod confractum fuerat, alligabo et, quod infirmum erat, consolidabo et, quod pingue et forte, custodiam et pascam illas in iudicio.
EZEK|34|17|Vos autem, grex meus, haec dicit Dominus Deus: Ecce ego iudico inter pecus et pecus, inter arietes et hircos.
EZEK|34|18|Nonne satis vobis erat pascuam bonam depasci? Insuper et reliquias pascuarum vestrarum conculcastis pedibus vestris et, cum purissimam aquam biberetis, reliquam pedibus vestris turbabatis;
EZEK|34|19|et oves meae his, quae conculcata pedibus vestris fuerant, pascebantur et, quae pedes vestri turbaverant, haec bibebant.
EZEK|34|20|Propterea haec dicit Dominus Deus ad eos: Ecce ego ipse iudico inter pecus pingue et macilentum;
EZEK|34|21|pro eo quod lateribus et umeris impingebatis et cornibus vestris ventilabatis omnia infirma pecora, donec dispergerentur foras,
EZEK|34|22|salvabo gregem meum, et non erit ultra in rapinam, et iudicabo inter pecus et pecus.
EZEK|34|23|Et suscitabo super eas pastorem unum, qui pascat eas, servum meum David; ipse pascet eas et ipse erit eis in pastorem.
EZEK|34|24|Ego autem Dominus ero eis in Deum, et servus meus David princeps in medio eorum. Ego Dominus locutus sum.
EZEK|34|25|Et faciam cum eis pactum pacis et cessare faciam bestias pessimas de terra, et habitabunt in deserto securi et dormient in saltibus;
EZEK|34|26|et ponam eos et, quae sunt in circuitu collis mei, benedictionem et deducam imbrem in tempore suo: pluviae benedictionis erunt.
EZEK|34|27|Et dabit lignum agri fructum suum, et terra dabit germen suum, et erunt in terra sua absque timore et scient quia ego Dominus, cum contrivero vectes iugi eorum et eruero eos de manu imperantium sibi.
EZEK|34|28|Et non erunt ultra in rapinam gentibus, neque bestiae terrae devorabunt eos, sed habitabunt confidenter absque ullo terrore.
EZEK|34|29|Et suscitabo eis germen nominatum, et non erunt ultra imminuti fame in terra neque portabunt ultra opprobrium gentium;
EZEK|34|30|et scient quia ego Dominus Deus eorum cum eis, et ipsi populus meus domus Israel, ait Dominus Deus.
EZEK|34|31|Vos autem grex meus, grex pascuae meae vos, et ego Dominus Deus vester, dicit Dominus Deus.
EZEK|35|1|Et factus est sermo Domini ad me dicens:
EZEK|35|2|" Fili hominis, pone faciem tuam adversum montem Seir et propheta de eo et dices illi:
EZEK|35|3|Haec dicit Dominus Deus:Ecce ego ad te, mons Seir;et extendam manum meam super teet dabo te desolatum atque desertum.
EZEK|35|4|Urbes tuas demoliar,et tu desertus eriset scies quia ego Dominus.
EZEK|35|5|Eo quod fueris inimicus sempiternus et concluseris filios Israel in manus gladii in tempore afflictionis eorum, in tempore poenae extremae;
EZEK|35|6|propterea, vivo ego, dicit Dominus Deus, sanguini tradam te, et sanguis te persequetur et, cum sanguinem non oderis, sanguis persequetur te.
EZEK|35|7|Et dabo montem Seir desolatum atque desertum et auferam de eo euntem et redeuntem
EZEK|35|8|et implebo montes eius occisorum suorum, in collibus tuis et in vallibus tuis, atque in omnibus torrentibus tuis interfecti gladio cadent.
EZEK|35|9|In solitudines sempiternas tradam te, et civitates tuae non habitabuntur, et scietis quoniam ego Dominus.
EZEK|35|10|Eo quod dixeris: "Duae gentes et duae terrae meae erunt, et hereditate possidebo eas!", cum Dominus esset ibi;
EZEK|35|11|propterea, vivo ego, dicit Dominus Deus, faciam iuxta iram tuam et secundum zelum tuum, quem fecisti odio habens eos, et notus efficiar in eis, cum te iudicavero.
EZEK|35|12|Et scies quia ego Dominus audivi universa opprobria tua, quae locutus es de montibus Israel dicens: "Deserti nobis ad devorandum dati sunt!".
EZEK|35|13|Et insurrexistis super me ore vestro et vociferati estis vobis adversum me verba vestra; ego audivi.
EZEK|35|14|Haec dicit Dominus Deus: Laetante universa terra, in solitudinem te redigam;
EZEK|35|15|sicuti gavisus es super hereditatem domus Israel, eo quod fuerit dissipata, sic faciam tibi: dissipatus eris, mons Seir, et Idumaea omnis, et scient quia ego Dominus.
EZEK|36|1|Tu autem, fili hominis, pro pheta super montes Israel et dices: Montes Israel, audite verbum Domini.
EZEK|36|2|Haec dicit Dominus Deus: Eo quod dixerit inimicus de vobis: "Euge, altitudines sempiternae in hereditatem datae sunt nobis";
EZEK|36|3|propterea vaticinare et dic: Haec dicit Dominus Deus: Pro eo quod desolati estis, et inhiaverunt vobis per circuitum, ut fieretis in hereditatem reliquis gentibus, et ascendistis super labium linguae et opprobrium populi;
EZEK|36|4|propterea, montes Israel, audite verbum Domini Dei: Haec dicit Dominus Deus montibus et collibus, torrentibus vallibusque et desertis dissipatis et urbibus derelictis, quae depopulatae sunt et subsannatae a reliquis gentibus per circuitum;
EZEK|36|5|propterea haec dicit Dominus Deus: In igne zeli mei locutus sum de reliquis gentibus et de Idumaea universa, quae dederunt terram meam sibi in hereditatem cum gaudio et toto corde et ex animo maligno, ut pascua eius depraedarentur.
EZEK|36|6|Idcirco vaticinare super humum Israel et dices montibus et collibus, torrentibus et vallibus: Haec dicit Dominus Deus: Ecce ego in zelo meo et in furore meo locutus sum, eo quod confusionem gentium sustinueritis;
EZEK|36|7|idcirco haec dicit Dominus Deus: Ego levavi manum meam: gentes, quae in circuitu vestro sunt, ipsae confusionem suam portabunt;
EZEK|36|8|vos autem, montes Israel, ramos vestros germinabitis et fructum vestrum afferetis populo meo Israel, prope est enim ut veniat.
EZEK|36|9|Quia ecce ego ad vos et convertar ad vos, et arabimini et accipietis sementem;
EZEK|36|10|et multiplicabo in vobis homines, omnem domum Israel, et habitabuntur civitates, et ruinosa instaurabuntur.
EZEK|36|11|Et replebo vos hominibus et iumentis, et multiplicabuntur et crescent; et habitari vos faciam, sicut a principio bonisque donabo maioribus quam habuistis ab initio, et scietis quia ego Dominus.
EZEK|36|12|Et adducam super vos homines, populum meum Israel, et hereditate possidebunt te, et eris eis in hereditatem et non addes ultra ut eos facias absque liberis.
EZEK|36|13|Haec dicit Dominus Deus: Pro eo quod dicunt de vobis: "Devoratrix hominum es et faciens gentem tuam absque liberis";
EZEK|36|14|propterea homines non comedes amplius et gentem tuam non facies ultra absque liberis, ait Dominus Deus.
EZEK|36|15|Nec auditam faciam in te amplius ignominiam gentium, et opprobrium populorum nequaquam portabis ultra et gentem tuam non facies amplius absque liberis ", ait Dominus Deus.
EZEK|36|16|Et factum est verbum Domini ad me dicens:
EZEK|36|17|" Fili hominis, domus Israel habitaverunt in humo sua et polluerunt eam in viis suis et in operibus suis; iuxta immunditiam menstruatae facta est via eorum coram me.
EZEK|36|18|Et effudi indignationem meam super eos pro sanguine, quem fuderunt super terram, et in idolis suis polluerunt eam.
EZEK|36|19|Et dispersi eos in gentes, et ventilati sunt in terras; iuxta vias eorum et iuxta opera eorum iudicavi eos.
EZEK|36|20|Et ingressi sunt ad gentes, ad quas introierunt, et polluerunt nomen sanctum meum, cum diceretur de eis: "Populus Domini iste est, et de terra eius egressi sunt".
EZEK|36|21|Et peperci nomini meo sancto, quod polluerat domus Israel in gentibus, ad quas ingressi sunt.
EZEK|36|22|Idcirco dices domui Israel: Haec dicit Domihus Deus: Non propter vos ego faciam, domus Israel, sed propter nomen sanctum meum, quod polluistis in gentibus, ad quas intrastis;
EZEK|36|23|et sanctificabo nomen meum magnum, quod pollutum est inter gentes, quod polluistis in medio earum, ut sciant gentes quia ego Dominus, ait Dominus Deus, cum sanctificatus fuero in vobis coram eis.
EZEK|36|24|Tollam quippe vos de gentibus et congregabo vos de universis terris et adducam vos in terram vestram;
EZEK|36|25|et effundam super vos aquam mundam, et mundabimini ab omnibus inquinamentis vestris, et ab universis idolis vestris mundabo vos.
EZEK|36|26|Et dabo vobis cor novum et spiritum novum ponam in medio vestri et auferam cor lapideum de carne vestra et dabo vobis cor carneum;
EZEK|36|27|et spiritum meum ponam in medio vestri et faciam, ut in praeceptis meis ambuletis et iudicia mea custodiatis et operemini.
EZEK|36|28|Et habitabitis in terra, quam dedi patribus vestris, et eritis mihi in populum, et ego ero vobis in Deum.
EZEK|36|29|Et salvabo vos ex universis inquinamentis vestris et vocabo frumentum et multiplicabo illud et non imponam vobis famem.
EZEK|36|30|Et multiplicabo fructum ligni et genimina agri, ut non portetis ultra opprobrium famis in gentibus.
EZEK|36|31|Et recordabimini viarum vestrarum pessimarum operumque non bonorum, et displicebunt vobis iniquitates vestrae et scelera vestra.
EZEK|36|32|Non propter vos ego faciam, ait Dominus Deus, notum sit vobis; confundimini et erubescite super viis vestris, domus Israel.
EZEK|36|33|Haec dicit Dominus Deus: In die, qua mundavero vos ex omnibus iniquitatibus vestris et inhabitari fecero urbes et instauravero ruinosa,
EZEK|36|34|et terra deserta fuerit exculta, quae quondam erat desolata in oculis omnis viatoris,
EZEK|36|35|dicent: "Terra illa inculta facta est ut hortus Eden, et civitates desertae et destitutae atque destructae munitae inhabitantur".
EZEK|36|36|Et scient gentes, quaecumque derelictae fuerint in circuitu vestro, quia ego Dominus aedificavi dissipata plantavique inculta; ego Dominus locutus sum et facio.
EZEK|36|37|Haec dicit Dominus Deus: Adhuc in hoc exorabor a domo Israel, ut faciam eis: multiplicabo eos sicut gregem hominum,
EZEK|36|38|ut gregem sanctum, ut gregem Ierusalem in sollemnitatibus eius; sic erunt civitates desertae plenae gregibus hominum, et scient quia ego Dominus ".
EZEK|37|1|Facta est super me manus Domini et eduxit me in spiri tu Domini et posuit me in medio campi, qui erat plenus ossibus,
EZEK|37|2|et circumduxit me per ea in gyro: erant autem multa valde super faciem campi siccaque vehementer.
EZEK|37|3|Et dixit ad me: " Fili hominis, putasne vivent ossa ista? ". Et dixi: " Domine, tu nosti ".
EZEK|37|4|Et dixit ad me: " Vaticinare super ossa ista et dices eis: Ossa arida, audite verbum Domini.
EZEK|37|5|Haec dicit Dominus Deus ossibus his: Ecce ego intromittam in vos spiritum, et vivetis,
EZEK|37|6|et dabo super vos nervos et succrescere faciam super vos carnes et superextendam in vobis cutem et dabo vobis spiritum, et vivetis et scietis quia ego Dominus ".
EZEK|37|7|Et prophetavi, sicut praeceperat mihi. Factus est autem sonitus, prophetante me, et ecce commotio; et accesserunt ossa ad ossa, unumquodque ad iuncturam suam.
EZEK|37|8|Et vidi: et ecce super ea nervi et carnes ascenderunt, et extenta est in eis cutis desuper, sed spiritum non habebant.
EZEK|37|9|Et dixit ad me: " Vaticinare ad spiritum; vaticinare, fili hominis, et dices ad spiritum: Haec dicit Dominus Deus: A quattuor ventis veni, spiritus, et insuffla super interfectos istos, ut reviviscant ".
EZEK|37|10|Et prophetavi, sicut praeceperat mihi, et ingressus est in ea spiritus; et vixerunt steteruntque super pedes suos, exercitus grandis nimis valde.
EZEK|37|11|Et dixit ad me: " Fili hominis, ossa haec universa domus Israel est. Ipsi dicunt: "Aruerunt ossa nostra, et periit spes nostra, et abscissi sumus".
EZEK|37|12|Propterea vaticinare et dices ad eos: Haec dicit Dominus Deus: Ecce ego aperiam tumulos vestros et educam vos de sepulcris vestris, populus meus, et inducam vos in terram Israel;
EZEK|37|13|et scietis quia ego Dominus, cum aperuero sepulcra vestra et eduxero vos de tumulis vestris, populus meus.
EZEK|37|14|Et dabo spiritum meum in vobis, et vivetis, et collocabo vos super humum vestram, et scietis quia ego Dominus. Locutus sum et facio ", ait Dominus Deus.
EZEK|37|15|Et factus est sermo Domini ad me dicens:
EZEK|37|16|" Et tu, fili hominis, sume tibi lignum unum et scribe super illud: Iudae et filiis Israel sociis eius. Et tolle lignum alterum et scribe super illud: Ioseph, lignum Ephraim, et cunctae domui Israel sociis eius.
EZEK|37|17|Et adiunge illa unum ad alterum tibi in lignum unum; et erunt in unionem in manu tua.
EZEK|37|18|Cum autem dixerint ad te filii populi tui loquentes: "Nonne indicas nobis, quid in his tibi velis?",
EZEK|37|19|loqueris ad eos: Haec dicit Dominus Deus: Ecce ego assumam lignum Ioseph, quod est in manu Ephraim, et tribus Israel, quae iunctae sunt ei, et dabo eas pariter cum ligno Iudae et faciam eas in lignum unum, et erunt unum in manu mea.
EZEK|37|20|Erunt autem ligna, super quae scripseris, in manu tua in oculis eorum,
EZEK|37|21|et dices ad eos: Haec dicit Dominus Deus: Ecce ego assumam filios Israel de medio nationum, ad quas abierunt, et congregabo eos undique et adducam eos ad humum suam
EZEK|37|22|et faciam eos in gentem unam in terra, in montibus Israel; et rex unus erit omnibus imperans, et non erunt ultra duae gentes nec dividentur amplius in duo regna.
EZEK|37|23|Neque polluentur ultra in idolis suis et abominationibus suis et in cunctis iniquitatibus suis, et salvos eos faciam de universis aversionibus suis, quibus peccaverunt, et mundabo eos, et erunt mihi populus, et ego ero eis Deus.
EZEK|37|24|Et servus meus David rex super eos, et pastor unus erit omnium eorum; in iudiciis meis ambulabunt et mandata mea custodient et facient ea.
EZEK|37|25|Et habitabunt super terram, quam dedi servo meo Iacob, in qua habitaverunt patres vestri; et habitabunt super eam, ipsi et filii eorum et filii filiorum eorum usque in sempiternum, et David servus meus princeps eorum in perpetuum.
EZEK|37|26|Et percutiam illis foedus pacis, pactum sempiternum erit eis, et fundabo eos et multiplicabo; et dabo sanctuarium meum in medio eorum in perpetuum,
EZEK|37|27|et erit habitaculum meum in eis, et ero eis Deus, et ipsi erunt mihi populus;
EZEK|37|28|et scient gentes quia ego Dominus sanctificator Israel, cum fuerit sanctuarium meum in medio eorum in perpetuum ".
EZEK|38|1|Et factus est sermo Domini ad me dicens:
EZEK|38|2|" Fili hominis, pone faciem tuam contra Gog, in terra Magog, principem summum Mosoch et Thubal, et vaticinare de eo
EZEK|38|3|et dices: Haec dicit Dominus Deus: Ecce ego ad te, Gog, principem summum Mosoch et Thubal,
EZEK|38|4|et circumagam te et ponam uncos in maxillis tuis et educam te et omnem exercitum tuum, equos et equites vestitos perfecte universos, multitudinem magnam cum scuto et clipeo arripientes gladium.
EZEK|38|5|Persae, Chus et Phut cum eis, omnes scutati et galeati;
EZEK|38|6|Gomer et universa agmina eius, domus Thogorma de extremo aquilone et totum robur eius, populi multi tecum.
EZEK|38|7|Praepara et instrue te et omnem multitudinem tuam, quae coacervata est ad te, et esto mihi in custodiam.
EZEK|38|8|Post dies multos evocaberis; in novissimo annorum venies ad terram, quae reversa est a gladio, congregata est de populis multis ad montes Israel, qui fuerunt deserti iugiter: haec de populis educta est, et habitant in ea confidenter universi.
EZEK|38|9|Ascendens autem quasi tempestas venies, quasi nubes, ut operias terram, tu et omnia agmina tua et populi multi tecum.
EZEK|38|10|Haec dicit Dominus Deus: In die illa ascendent sermones super cor tuum, et cogitabis cogitationem pessimam
EZEK|38|11|et dices: "Ascendam ad terram absque muro, veniam ad quiescentes habitantesque secure; hi omnes habitant sine muro, vectes et portae non sunt eis";
EZEK|38|12|ut diripias spolia et capias praedam, ut inferas manum tuam super deserta iterum inhabitata et super populum, qui est congregatus ex gentibus, qui acquisivit pecora et substantiam et habitat in umbilico terrae.
EZEK|38|13|Saba et Dedan et negotiatores Tharsis et omnes principes eius dicent tibi: "Numquid ad sumenda spolia tu venis? Numquid ad diripiendam praedam congregasti multitudinem tuam, ut tollas argentum et aurum, auferas pecora atque substantiam et diripias manubias infinitas?".
EZEK|38|14|Propterea vaticinare, fili hominis, et dices ad Gog: Haec dicit Dominus Deus: Numquid non in die illo, cum habitaverit populus meus Israel confidenter, consurges?
EZEK|38|15|Et venies de loco tuo ab extremo aquilone, tu et populi multi tecum, ascensores equorum universi, coetus magnus et exercitus vehemens.
EZEK|38|16|Et ascendes super populum meum Israel quasi nubes, ut operias terram. In novissimis diebus erit, et adducam te super terram meam, ut sciant gentes me, cum sanctificatus fuero in te in oculis eorum, o Gog.
EZEK|38|17|Haec dicit Dominus Deus: Tu ergo ille es, de quo locutus sum in diebus antiquis in manu servorum meorum prophetarum Israel, qui prophetaverunt in diebus illis per annos, ut adducerem te super eos.
EZEK|38|18|Et erit in die illa, in die adventus Gog super terram Israel, ait Dominus Deus, ascendet indignatio mea in furore meo.
EZEK|38|19|Et in zelo meo, in igne irae meae locutus sum: In die illa erit commotio magna super terram Israel,
EZEK|38|20|et commovebuntur a facie mea pisces maris et volucres caeli et bestiae agri et omne reptile, quod movetur super humum, cunctique homines, qui sunt super faciem terrae; et subvertentur montes, et cadent rupes, et omnis murus in terram corruet.
EZEK|38|21|Et convocabo adversus eum in cunctis montibus meis gladium, ait Dominus Deus; gladius uniuscuiusque in fratrem suum dirigetur.
EZEK|38|22|Et iudicabo eum peste et sanguine et imbre vehementi et lapidibus grandinis; ignem et sulphur pluam super eum et super exercitum eius et super populos multos, qui sunt cum eo,
EZEK|38|23|et magnificabor et sanctificabor et notus ero in oculis multarum gentium, et scient quia ego Dominus.
EZEK|39|1|Tu autem, fili hominis, va ticinare adversum Gog et dices: Haec dicit Dominus Deus: Ecce ego super te, Gog, principem summum Mosoch e Thubal;
EZEK|39|2|et circumagam te et seducam te et ascendere faciam de extremo aquilone et adducam te super montes Israel.
EZEK|39|3|Et percutiam arcum tuum in manu sinistra tua et sagittas tuas de manu dextera tua deiciam.
EZEK|39|4|Super montes Israel cades, tu et omnia agmina tua et populi, qui sunt tecum; feris avibus, omni volatili et bestiis terrae dedi te devorandum:
EZEK|39|5|super faciem agri cades, quia ego locutus sum, ait Dominus Deus.
EZEK|39|6|Et emittam ignem in Magog et in his, qui habitant in insulis confidenter, et scient quia ego Dominus.
EZEK|39|7|Et nomen sanctum meum notum faciam in medio populi mei Israel et non polluam nomen sanctum meum amplius, et scient gentes quia ego Dominus, sanctus in Israel.
EZEK|39|8|Ecce venit et fit, ait Dominus Deus; haec est dies, de qua locutus sum.
EZEK|39|9|Et egredientur habitatores de civitatibus Israel et succendent et comburent arma, clipeum et scutum, arcum et sagittas et baculos, manus et contos, et succendent ea igne septem annis.
EZEK|39|10|Et non portabunt ligna de campis neque succident de saltibus, quoniam arma succendent igne et depraedabuntur eos, quibus praedae fuerant, et diripient vastatores suos, ait Dominus Deus.
EZEK|39|11|Et erit, in die illa dabo Gog locum nominatum sepulcrum in Israel, vallem viatorum ad orientem maris, quae oppilat viam praetereuntibus; et sepelient ibi Gog et omnem multitudinem eius, et vocabitur vallis Multitudinis Gog.
EZEK|39|12|Et sepelient eos domus Israel, ut mundent terram septem mensibus;
EZEK|39|13|sepeliet autem eum omnis populus terrae, et erit eis nominata dies, in qua glorificatus sum, ait Dominus Deus.
EZEK|39|14|Et viros iugiter constituent lustrantes terram, qui sepeliant eos, qui remanserant super faciem terrae, ut emundent eam; post menses autem septem quaerere incipient
EZEK|39|15|et circuibunt peragrantes terram; cumque viderint os hominis, statuent iuxta illud titulum, donec sepeliant illud pollinctores in valle Multitudinis Gog.
EZEK|39|16|Nomen quoque civitatis Amona, et mundabunt terram.
EZEK|39|17|Tu ergo, fili hominis, haec dicit Dominus Deus, dic volucri, universis avibus cunctisque bestiis agri: Convenite, properate, concurrite undique ad victimam meam, quam ego immolo vobis, victimam grandem super montes Israel, ut comedatis carnes et bibatis sanguinem.
EZEK|39|18|Carnes fortium comedetis et sanguinem principum terrae bibetis: arietes, agni et hirci taurique saginati de Basan sunt omnes;
EZEK|39|19|et comedetis adipem in saturitatem et bibetis sanguinem in ebrietatem de victima, quam ego immolabo vobis.
EZEK|39|20|Et saturabimini super mensam meam de equo et de iugali currus, de forti et de universis viris bellatoribus, ait Dominus Deus.
EZEK|39|21|Et ponam gloriam meam in gentibus, et videbunt omnes gentes iudicium meum, quod fecerim, et manum meam, quam posuerim super eos;
EZEK|39|22|et scient domus Israel quia ego Dominus Deus eorum a die illa et deinceps,
EZEK|39|23|et scient gentes quoniam in iniquitate sua capta sit domus Israel, eo quod reliquerint me, et absconderim faciem meam ab eis et tradiderim eos in manus hostium suorum, et ceciderint in gladio universi.
EZEK|39|24|Iuxta immunditiam eorum et scelera eorum feci eis et abscondi faciem meam ab illis.
EZEK|39|25|Propterea haec dicit Dominus Deus: Nunc restituam Iacob et miserebor omnis domus Israel et assumam zelum pro nomine sancto meo.
EZEK|39|26|Et portabunt confusionem suam et omnem praevaricationem, quam praevaricati sunt in me, cum habitaverint in terra sua confidenter; et nemo erit qui exterreat.
EZEK|39|27|Et reduxero eos de populis et congregavero de terris inimicorum suorum et sanctificatus fuero in eis in oculis gentium plurimarum,
EZEK|39|28|et scient quia ego Dominus Deus eorum, eo quod transtulerim eos in nationes et congregaverim eos super terram suam et non dereliquerim quemquam ex eis ibi.
EZEK|39|29|Et non abscondam ultra faciem meam ab eis, eo quod effuderim spiritum meum super domum Israel ", ait Dominus Deus.
EZEK|40|1|In vicesimo et quinto anno transmigrationis nostrae, in exordio anni, decima mensis, quarto decimo anno, postquam percussa est civitas, in ipsa hac die facta est super me manus Domini et adduxit me illuc.
EZEK|40|2|In visionibus Dei adduxit me in terram Israel et posuit me super montem excelsum nimis, super quem erat quasi aedificium civitatis ad austrum.
EZEK|40|3|Et introduxit me illuc; et ecce vir, cuius erat species quasi species aeris, et funiculus lineus in manu eius, et calamus mensurae in manu eius, stabat autem in porta.
EZEK|40|4|Et locutus est ad me idem vir: " Fili hominis, vide oculis tuis et auribus tuis audi et pone cor tuum in omnia, quae ego ostendam tibi, quia ut ostendantur tibi, adductus es huc; annuntia omnia, quae tu vides, domui Israel ".
EZEK|40|5|Et ecce murus forinsecus in circuitu domus undique, et in manu viri calamus mensurae sex cubitorum, qui habebant cubitum et palmum; et mensus est latitudinem aedificii calamo uno, altitudinem quoque calamo uno.
EZEK|40|6|Et venit ad portam, quae respiciebat viam orientalem, et ascendit per gradus eius et mensus est limen portae calamo uno latitudinem
EZEK|40|7|et cubiculum uno calamo in longum et uno calamo in latum et inter cubicula quinque cubitos et limen portae iuxta vestibulum portae intrinsecus calamo uno.
EZEK|40|8|Et mensus est vestibulum portae
EZEK|40|9|octo cubitorum et postem eius duobus cubitis; vestibulum autem portae erat intrinsecus.
EZEK|40|10|Porro cubicula portae ad viam orientalem, tria hinc et tria inde, mensura una trium et mensura una postium ex utraque parte.
EZEK|40|11|Et mensus est latitudinem ostii portae decem cubitorum et longitudinem portae tredecim cubitorum,
EZEK|40|12|et saeptum ante cubicula cubiti unius utrimque; cubicula autem sex cubitorum erant hinc et inde.
EZEK|40|13|Et mensus est portam a tecto cubiculi usque ad tectum eius a contra, latitudinem viginti et quinque cubitorum, ostium contra ostium,
EZEK|40|14|()
EZEK|40|15|et a facie ingressus portae usque ad faciem vestibuli portae intrinsecus, quinquaginta cubitos.
EZEK|40|16|Et erant fenestrae marginatae in cubiculis et in postibus intra portam undique per circuitum; similiter autem erant et in vestibulo fenestrae per gyrum intrinsecus, et ante postes pictura palmarum.
EZEK|40|17|Et eduxit me ad atrium exterius, et ecce exedrae et pavimentum stratum lapide in atrio per circuitum, triginta exedrae in circuitu pavimenti;
EZEK|40|18|et pavimentum ad latus portarum secundum longitudinem portarum; hoc erat pavimentum inferius.
EZEK|40|19|Et mensus est latitudinem a facie portae inferioris usque ad frontem portae interioris extrinsecus, centum cubitos. Sic oriens. Et sic aquilo.
EZEK|40|20|Portam quoque, quae respiciebat viam aquilonis atrii exterioris, mensus est, tam in longitudine quam in latitudine;
EZEK|40|21|et cubicula eius, tria hinc et tria inde, et postes eius et vestibulum eius secundum mensuram portae prioris; quinquaginta cubitorum longitudo eius et latitudo viginti quinque cubitorum.
EZEK|40|22|Et fenestrae vestibuli eius et sculpturae palmarum secundum mensuram portae, quae respiciebat ad orientem; et septem graduum erat ascensus eius, et vestibulum intrinsecus.
EZEK|40|23|Et porta atrii interioris contra portam aquilonis sicut in porta orientali; et mensus est a porta usque ad portam centum cubitos.
EZEK|40|24|Et duxit me ad viam australem, et ecce porta, quae respiciebat ad austrum; et mensus est postes eius et vestibulum eius iuxta mensuras superiores.
EZEK|40|25|Et fenestrae eius et vestibuli in circuitu sicut fenestrae ceterae; quinquaginta cubitorum longitudo erat et latitudo viginti quinque cubitorum.
EZEK|40|26|Et in gradibus septem ascendebatur ad eam, et vestibulum erat intrinsecus, et caelatae palmae erant, una hinc et altera inde, in postibus eius.
EZEK|40|27|Et porta erat atrio interiori in via australi, et mensus est a porta usque ad portam in via australi centum cubitos.
EZEK|40|28|Et introduxit me in atrium interius per portam australem et mensus est portam iuxta mensuras superiores;
EZEK|40|29|cubicula eius et postes eius, et vestibulum eius eisdem mensuris; et fenestrae erant ei et vestibulo eius in circuitu. Quinquaginta cubitorum longitudo erat et latitudo viginti quinque cubitorum.
EZEK|40|30|()
EZEK|40|31|Et vestibulum eius respiciebat ad atrium exterius, et palmae in postibus eius, et octo gradus erant, quibus ascendebatur ad eam.
EZEK|40|32|Et introduxit me in atrium interius per viam orientalem et mensus est portam secundum mensuras superiores;
EZEK|40|33|cubicula eius et postes eius et vestibulum eius sicut supra; et fenestrae erant ei et vestibulo eius in circuitu. Longitudo erat quinquaginta cubitorum et latitudo viginti quinque cubitorum.
EZEK|40|34|Et vestibulum eius respiciebat ad atrium exterius, et palmae caelatae in postibus eius hinc et inde et in octo gradibus ascensus eius.
EZEK|40|35|Et introduxit me ad portam, quae respiciebat ad aquilonem, et mensus est secundum mensuras superiores
EZEK|40|36|cubicula eius et postes eius et vestibulum eius; et fenestrae ei erant per circuitum. Longitudo quinquaginta cubitorum erat et latitudo viginti quinque cubitorum.
EZEK|40|37|Et vestibulum eius respiciebat ad atrium exterius, et caelatura palmarum in postibus illius hinc et inde et in octo gradibus ascensus eius.
EZEK|40|38|Et erat exedra, cuius ostium in vestibulo portae; ibi lavabunt holocaustum.
EZEK|40|39|Et in vestibulo portae duae mensae hinc et duae mensae inde, ut mactetur super eas holocaustum et pro peccato et pro delicto.
EZEK|40|40|Et ad latus extra vestibulum ad ostium portae, quae respicit ad aquilonem, duae mensae; et ad la tus alterum vestibuli portae duae mensae.
EZEK|40|41|Quattuor mensae hinc et quattuor mensae inde ad latus portae: octo mensae erant, super quas mactabunt.
EZEK|40|42|Quattuor autem mensae ad holocaustum de lapidibus quadris exstructae longitudine cubiti unius et dimidii et latitudine cubiti unius et dimidii et altitudine cubiti unius, super ista ponant vasa, quibus mactetur holocaustum et victima,
EZEK|40|43|et labia palmi unius reflexa intrinsecus per circuitum; super mensas autem carnes oblationis.
EZEK|40|44|Et extra portam interiorem exedrae duae, in atrio interiori; una erat in latere portae respicientis ad aquilonem, et facies eius contra viam australem, et una ex latere portae australis, quae respiciebat ad viam aquilonis.
EZEK|40|45|Et dixit ad me: " Haec est exedra, quae respicit viam meridianam; sacerdotum erit, qui excubant in custodiis templi.
EZEK|40|46|Porro exedra, quae respicit ad viam aquilonis, sacerdotum erit, qui excubant ad ministerium altaris: isti sunt filii Sadoc, qui accedunt de filiis Levi ad Dominum, ut ministrent ei ".
EZEK|40|47|Et mensus est atrium longitudine centum cubitorum et latitudine centum cubitorum per quadrum. Altare autem erat ante faciem templi.
EZEK|40|48|Et introduxit me in vestibulum templi; et mensus est postes vestibuli quinque cubitis hinc et quinque cubitis inde et latitudinem portae quattuordecim cubitorum et latera portae trium cubitorum hinc et trium cubitorum inde;
EZEK|40|49|longitudinem autem vestibuli viginti cubitorum et latitudinem duodecim cubitorum, et decem gradibus ascendebatur ad illud, et columnae erant in postibus, una hinc et altera inde.
EZEK|41|1|Et introduxit me in templum et mensus est postes: sex cu bitos latitudinis hinc et sex cubitos latitudinis inde.
EZEK|41|2|Et latitudo portae decem cubitorum erat, et latera portae quinque cubitis hinc et quinque cubitis inde; et mensus est longitudinem eius quadraginta cubitorum et latitudinem viginti cubitorum.
EZEK|41|3|Et introgressus intrinsecus, mensus est in poste portae duos cubitos et portam sex cubitorum et latitudinem laterum portae septem cubitorum hinc et septem cubitorum inde.
EZEK|41|4|Et mensus est longitudinem eius viginti cubitorum et latitudinem viginti cubitorum versus faciem templi. Et dixit ad me: " Hoc est Sanctum sanctorum ".
EZEK|41|5|Et mensus est parietem domus sex cubitorum et latitudinem aedificii adiacentis quattuor cubitorum undique per circuitum domus;
EZEK|41|6|cubicula autem adiacentia, cubiculum super cubiculum, in tribus tabulatis. Et erant margines eminentes in pariete domus pro cubiculis adiacentibus per circuitum, ut essent fulcra, neque essent fulcra intra parietem domus,
EZEK|41|7|et latitudo ambitus sursum ascendens iuxta cubicula adiacentia, quia circumdata erat domus usque sursum circa domum; idcirco amplificata erat domus usque sursum, et de inferiore tabulato ascendebatur ad superius per medium.
EZEK|41|8|Et vidi in domo altitudinem per circuitum, fundamenta aedificii adiacentis mensura calami pleni, id est sex cubitorum, in altitudine.
EZEK|41|9|Et latitudo parietis aedificii adiacentis forinsecus erat quinque cubitorum. Et area vacua inter cubicula domui adiacentia,
EZEK|41|10|et inter exedras habebat latitudinem viginti cubitorum in circuitu domus undique.
EZEK|41|11|Et ostia aedificii adiacentis ad aream vacuam, ostium unum ad viam aquilonis et ostium unum ad viam australem; et latitudo muri areae vacuae quinque cubitorum in circuitu.
EZEK|41|12|Et aedificium, quod erat ex adverso areae separatae versumque ad viam respicientem ad mare, latitudinis septuaginta cubitorum; paries autem aedificii quinque cubitorum latitudinis per circuitum et longitudo eius nonaginta cubitorum.
EZEK|41|13|Et mensus est domus longitudinem centum cubitorum et areae separatae et aedificii et parietum eius longitudinem centum cubitorum;
EZEK|41|14|latitudinem autem faciei domus et areae separatae contra orientem centum cubitorum.
EZEK|41|15|Et mensus est longitudinem aedificii ex adverso areae separatae ad dorsum et parietum eius ex utraque parte centum cubitorum. Et templum interius et vestibulum exterius
EZEK|41|16|strata erant ligno, et fenestrae marginatae et margines in circuitu triplices contra limen erant strato ligno per gyrum in circuitu, et a terra usque ad fenestras - et fenestrae poterant claudi - usque ad superiora ostii;
EZEK|41|17|et usque ad domum interiorem et forinsecus et per omnem parietem in circuitu, intrinsecus et forinsecus, ad mensuram
EZEK|41|18|fabrefacti cherubim et palmae, et palma inter cherub et cherub; duasque facies habebat cherub,
EZEK|41|19|faciem hominis versam ad palmam ex hac parte et faciem leonis versam ad palmam ex alia parte: expressi per omnem domum in circuitu.
EZEK|41|20|De terra usque ad superiora portae cherubim et palmae caelatae erant. In pariete templi
EZEK|41|21|postes portae quadruplices, et coram sanctuario aspectus quasi aspectus
EZEK|41|22|altaris lignei trium cubitorum altitudo, et longitudo eius duorum cubitorum, et anguli eius et bases eius et parietes eius lignei. Et locutus est ad me: " Haec est mensa coram Domino ".
EZEK|41|23|Et duo ostia erant templo et sanctuario
EZEK|41|24|duo ostia. Ostiis erant duae valvae versatiles usque ad parietem, valvae duae ostio uni et valvae duae ostio alteri.
EZEK|41|25|Et caelati erant in ipsis ostiis templi cherubim et sculpturae palmarum, sicut in parietibus quoque expressi erant; et tectum ligneum erat in vestibuli fronte forinsecus.
EZEK|41|26|Et fenestrae marginatae et similitudo palmarum hinc atque inde in lateribus vestibuli et in cubiculis adiacentibus domus.
EZEK|42|1|Et eduxit me in atrium ex terius per viam ducentem ad aquilonem; et duxit me ad exedram, quae erat contra aream separatam, et contra aedem ad aquilonem.
EZEK|42|2|Longitudo erat centum cubitorum in latere aquilonis et latitudo quinquaginta cubitorum.
EZEK|42|3|Contra viginti cubitos atrii interioris et contra pavimentum stratum lapide atrii exterioris elevabatur pars iuxta partem in tribus gradibus.
EZEK|42|4|Et ante exedras deambulatio decem cubitorum latitudinis, ad interiora respiciens, longitudinis centum cubitorum; et ostia eorum ad aquilonem.
EZEK|42|5|Exedrae superiores angustiores erant, quia gradus auferebant eis spatium, prae inferioribus et mediis aedificii.
EZEK|42|6|Tristega enim erant et non habebant columnas, sicut erant columnae exteriorum; sic ergo in gradibus de inferioribus, et de mediis a terra surgebat aedificium.
EZEK|42|7|Et murus exterior secundum exedras erat in via atrii exterioris ante exedras, longitudo eius quinquaginta cubitorum,
EZEK|42|8|quia longitudo erat exedrarum atrii exterioris quinquaginta cubitorum, quae erant ante faciem illarum, totum erat centum cubitorum.
EZEK|42|9|Et erat subter exedras has introitus ab oriente ingredientibus in ea de atrio exteriori
EZEK|42|10|in capite muri atrii. Contra viam meridianam in facie areae separatae, et erant exedrae ante aedificium,
EZEK|42|11|et via ante faciem earum iuxta similitudinem exedrarum, quae erant in via aquilonis; secundum longitudinem earum et latitudinem earum, sic et omnes exitus earum et dispositiones et ostia earum.
EZEK|42|12|Et ad ostia exedrarum, quae erant in via respiciente ad notum, ostium in capite viae, quae via erat ante murum protegentem per viam orientalem ingredientibus.
EZEK|42|13|Et dixit ad me: "Exedrae aquilonis et exedrae austri, quae sunt ante aream separatam, hae sunt exedrae sanctae, in quibus vescuntur sacerdotes, qui appropinquant ad Dominum sancta sanctorum: ibi ponent sancta sanctorum et oblationem et pro peccato et pro delicto, locus enim sanctus est.
EZEK|42|14|Cum autem ingressi fuerint sacerdotes, non egredientur de sanctis in atrium exterius, sed ibi reponent vestimenta sua, in quibus ministrant, quia sancta sunt; vestienturque vestimentis aliis et sic procedent ad locum populi ".
EZEK|42|15|Cumque complesset mensuras interioris areae domus, eduxit me per viam portae, quae respiciebat ad viam orientalem, et mensus est ibi undique per circuitum.
EZEK|42|16|Mensus est autem contra ventum orientalem calamo mensurae quingentos calamos in calamo mensurae per circuitum.
EZEK|42|17|Et mensus est contra ventum aquilonis quingentos calamos in calamo mensurae per gyrum.
EZEK|42|18|Et ad ventum australem mensus est quingentos calamos in calamo mensurae per circuitum.
EZEK|42|19|Et conversus ad ventum occidentalem mensus est quingentos calamos in calamo mensurae.
EZEK|42|20|Per quattuor ventos mensus est illud; murus ei erat undique per circuitum longitudine quingentorum cubitorum et latitudine quingentorum cubitorum, dividens inter sanctuarium et locum profanum.
EZEK|43|1|Et duxit me ad portam, quae respiciebat ad viam orientalem,
EZEK|43|2|et ecce gloria Dei Israel ingrediebatur per viam orientalem, et vox erat ei quasi vox aquarum multarum, et terra splendebat a maiestate eius.
EZEK|43|3|Et vidi visionem secundum speciem, quam videram, quando venit, ut disperderet civitatem, et species secundum aspectum, quem videram iuxta fluvium Chobar; et cecidi super faciem meam.
EZEK|43|4|Et maiestas Domini ingressa est templum per viam portae, quae respiciebat ad orientem.
EZEK|43|5|Et levavit me spiritus et introduxit me in atrium interius; et ecce repleta erat gloria Domini domus.
EZEK|43|6|Et audivi loquentem ad me de domo, cum vir staret iuxta me,
EZEK|43|7|et dixit ad me: " Fili hominis, locus solii mei et locus vestigiorum pedum meorum, ubi habitabo in medio filiorum Israel in aeternum; et non polluent ultra domus Israel nomen sanctum meum, ipsi et reges eorum, in fornicationibus suis et in cadaveribus regum suorum in morte eorum,
EZEK|43|8|qui fabricati sunt limen suum iuxta limen meum et postes suos iuxta postes meos, et paries erat inter me et eos, et polluerunt nomen sanctum meum in abominationibus, quas fecerunt; propter quod consumpsi eos in ira mea.
EZEK|43|9|Nunc ergo repellant procul fornicationem suam et cadavera regum suorum a me, et habitabo in medio eorum semper.
EZEK|43|10|Tu autem, fili hominis, ostende domui Israel templum, et confundantur ab iniquitatibus suis et metiantur fabricam.
EZEK|43|11|Et si erubuerint ex omnibus, quae fecerunt, describe domum et supellectilem eius, exitus et introitus, et omnem figuram eius et universa praecepta eius et omnes leges eius ostende eis et scribes oculis eorum, ut custodiant omnem figuram eius et omnia praecepta illius et faciant ea.
EZEK|43|12|Ista est lex domus in summitate montis: omnes fines eius in circuitu sanctum sanctorum sunt; haec est ergo lex domus ".
EZEK|43|13|Istae autem mensurae altaris in cubitis, cubitus habebat cubitum et palmum; fossae in circuitu eius erat cubitus in altitudine et cubitus in latitudine; et saepto eius ad marginem eius in circuitu palmus unus. Haec autem erat altitudo altaris:
EZEK|43|14|de fossa terrae usque ad crepidinem inferiorem duo cubiti, et latitudo cubiti unius; et a crepidine minore usque ad crepidinem maiorem quattuor cubiti, et latitudo unius cubiti.
EZEK|43|15|Ipse autem focus quattuor cubitorum, et a foco usque sursum cornua quattuor.
EZEK|43|16|Et focus duodecim cubitorum in longitudine per duodecim cubitos latitudinis, quadrangulatum aequis lateribus.
EZEK|43|17|Et crepido quattuordecim cubitorum longitudinis per quattuordecim cubitos latitudinis in quattuor angulis eius; et saeptum in circuitu eius dimidii cubiti, et fossa eius unius cubiti per circuitum; gradus autem eius versi ad orientem.
EZEK|43|18|Et dixit ad me: " Fili hominis, haec dicit Dominus Deus: Hi sunt ritus altaris: in qua die fuerit fabricatum, ut offeratur super illud holocaustum, et effundatur sanguis,
EZEK|43|19|dabis sacerdotibus levitis, qui sunt de semine Sadoc, qui accedunt ad me, ait Dominus Deus, ut ministrent mihi, vitulum de armento pro peccato.
EZEK|43|20|Et assumens de sanguine eius, pones super quattuor cornua eius et super quattuor angulos crepidinis et super saeptum in circuitu et mundabis illud et expiabis.
EZEK|43|21|Et tolles vitulum, qui oblatus fuerit pro peccato, et combures illum in destinato loco domus extra sanctuarium.
EZEK|43|22|Et in die secunda offeres hircum caprarum immaculatum pro peccato, et expiabunt altare, sicut expiaverunt in vitulo.
EZEK|43|23|Cumque compleveris expians illud, offeres vitulum de armento immaculatum et arietem de grege immaculatum;
EZEK|43|24|et offeres eos in conspectu Domini, et mittent sacerdotes super eos sal et offerent eos holocaustum Domino.
EZEK|43|25|Septem diebus facies hircum pro peccato cotidie, et vitulum de armento et arietem de pecoribus immaculatos offerent.
EZEK|43|26|Septem diebus expiabunt altare et mundabunt illud et consecrabunt illud.
EZEK|43|27|Expletis autem diebus, in die octava et ultra facient sacerdotes super altare holocausta vestra et pacifica, et placatus ero vobis ", ait Dominus Deus.
EZEK|44|1|Et convertit me ad viam portae sanctuarii exterioris, quae respiciebat ad orientem, et erat clausa;
EZEK|44|2|et dixit Dominus ad me: " Porta haec clausa erit; non aperietur, et vir non transibit per eam, quoniam Dominus, Deus Israel, ingressus est per eam, eritque clausa.
EZEK|44|3|Princeps, ut princeps ipse sedebit in ea, ut comedat panem coram Domino; per viam vestibuli portae ingredietur et per eandem viam egredietur ".
EZEK|44|4|Et adduxit me per viam portae aquilonis in conspectum domus; et vidi: et ecce implevit gloria Domini domum Domini, et cecidi in faciem meam.
EZEK|44|5|Et dixit ad me Dominus: " Fili hominis, pone cor tuum et vide oculis tuis et auribus tuis audi omnia, quae ego loquor ad te de universis caeremoniis domus Domini et de cunctis legibus eius; et pones cor tuum in introitu templi et in omni exitu sanctuarii
EZEK|44|6|et dices ad exasperantem me domum Israel: Haec dicit Dominus Deus: Sufficiant vobis omnes abominationes vestrae, domus Israel,
EZEK|44|7|eo quod induxistis alienigenas incircumcisos corde et incircumcisos carne, ut essent in sanctuario meo et polluerent domum meam, cum offertis panem meum, adipem et sanguinem; et dissolvistis pactum meum in omnibus abominationibus vestris
EZEK|44|8|et non explevistis ministerium sanctorum meorum et posuistis illos ministrantes mihi in sanctuario meo. Propterea
EZEK|44|9|haec dicit Dominus Deus: Omnis alienigena incircumcisus corde et incircumcisus carne non ingredietur sanctuarium meum, omnis alienigena, qui est in medio filiorum Israel.
EZEK|44|10|Sed Levitae, qui longe recesserint a me in errore filiorum Israel, qui erraverunt a me post idola sua, portabunt iniquitatem suam
EZEK|44|11|et erunt in sanctuario meo aeditui et ianitores portarum domus et ministri domus: ipsi mactabunt holocausta et victimas populo et ipsi stabunt in conspectu eorum, ut ministrent eis.
EZEK|44|12|Pro eo quod ministraverunt illis in conspectu idolorum suorum et facti sunt domui Israel in offendiculum iniquitatis, idcirco levavi manum meam super eos, dicit Dominus Deus; portabunt iniquitatem suam.
EZEK|44|13|Et non appropinquabunt ad me, ut sacerdotio fungantur mihi, neque accedent ad omnia sancta mea, ad sanctissima, sed portabunt confusionem suam et abominationes suas, quas fecerunt.
EZEK|44|14|Et faciam eos ministros in omni ministerio domus et in universis, quae facienda sunt in ea.
EZEK|44|15|Sacerdotes autem levitae filii Sadoc, qui custodierunt caeremonias sanctuarii mei, cum errarent filii Israel a me, ipsi accedent ad me, ut ministrent mihi, et stabunt in conspectu meo, ut offerant mihi adipem et sanguinem, ait Dominus Deus.
EZEK|44|16|Ipsi ingredientur sanctuarium meum et ipsi accedent ad mensam meam, ut serviant mihi et custodiant ministerium meum.
EZEK|44|17|Cumque ingredientur portas atrii interioris, vestibus lineis induentur, nec ascendet super eos quidquam laneum, quando ministrant in portis atrii interioris et in domo.
EZEK|44|18|Vittae lineae erunt in capitibus eorum, et feminalia linea erunt in lumbis eorum, et non accingentur in sudore.
EZEK|44|19|Cumque egredientur atrium exterius ad populum, exuent se vestimenta sua, in quibus ministraverunt, et reponent ea in exedris sanctis et vestient se vestimentis aliis et non sanctificabunt populum in vestibus suis.
EZEK|44|20|Caput autem suum non radent neque comam nutrient, sed tondentes attondent capita sua.
EZEK|44|21|Et vinum non bibet omnis sacerdos, quando ingressurus est atrium interius.
EZEK|44|22|Et viduam et repudiatam non accipient sibi uxores sed virgines de semine domus Israel; sed et viduam, quae fuerit vidua a sacerdote, accipient.
EZEK|44|23|Et populum meum docebunt quid sit inter sanctum et profanum et inter mundum et immundum ostendent eis.
EZEK|44|24|Et cum fuerit controversia, stabunt ad iudicandum et in iudiciis meis iudicabunt; leges meas et praecepta mea in omnibus sollemnitatibus meis custodient et sabbata mea sanctificabunt.
EZEK|44|25|Et ad mortuum hominem non ingredientur, ne polluantur, nisi ad patrem et matrem et filium et filiam et fratrem et sororem, quae virum non habuit: in quibus contaminabuntur.
EZEK|44|26|Et postquam fuerit emundatus, septem dies numerabuntur ei,
EZEK|44|27|et in die introitus sui in sanctuarium ad atrium interius, ut ministret mihi in sanctuario, offeret pro peccato suo, ait Dominus Deus.
EZEK|44|28|Et erit eis in hereditatem: ego hereditas eorum; et possessionem non dabitis eis in Israel: ego enim possessio eorum.
EZEK|44|29|Oblationem et pro peccato et pro delicto ipsi comedent, et omne anathema in Israel ipsorum erit;
EZEK|44|30|et primitiva omnium primogenitorum et omnia libamenta ex omnibus, quae offertis, sacerdotum erunt; et primitiva farinae vestrae dabitis sacerdoti, ut reponat benedictionem domui tuae.
EZEK|44|31|Omne morticinum et captum a bestia de avibus et de pecoribus non comedent sacerdotes.
EZEK|45|1|Cumque coeperitis terram dividere sortito, separate oblationem Domino sanctificatum de terra, longitudine viginti quinque milia et latitudine viginti milia: sanctificatum erit in omni termino suo per circuitum;
EZEK|45|2|ex quo sanctuarium obtinebit quingentos per quingentos, quadrifariam per circuitum, et quinquaginta cubitos pascua eius per gyrum.
EZEK|45|3|Et a mensura ista mensurabis longitudinem viginti quinque milium et latitudinem decem milium, et in ipso erit templum, Sanctum sanctorum.
EZEK|45|4|Sanctificatum de terra erit sacerdotibus ministris sanctuarii, qui accedunt ad ministerium Domini; et erit eis locus in domos et in pascua pecoribus.
EZEK|45|5|Viginti quinque autem milia longitudinis et decem milia latitudinis erunt Levitis, qui ministrant domui; ipsis in possessionem, civitates ad habitandum.
EZEK|45|6|Et possessionem civitatis dabitis quinque milia latitudinis et longitudinis viginti quinque milia, iuxta oblationem sacram; omni domui Israel erit.
EZEK|45|7|Principi quoque ex utraque parte oblationis sacrae et possessionis civitatis, secundum oblationem sacram et possessionem urbis, a latere maris usque ad mare et a latere orientis versus orientem, longitudinem autem iuxta unamquamque partium, a termino occidentali usque ad terminum orientalem.
EZEK|45|8|Haec terra erit ei possessio in Israel, et non depopulabuntur ultra principes mei populum meum; sed terram dabunt domui Israel secundum tribus eorum.
EZEK|45|9|Haec dicit Dominus Deus: Sufficiat vobis, principes Israel; violentiam et rapinas omittite et iudicium et iustitiam facite; auferte exactiones vestras a populo meo, ait Dominus Deus.
EZEK|45|10|Statera iusta et ephi iustum et batus iustus sit vobis;
EZEK|45|11|ephi et batus aequalia et unius mensurae sint, ut capiat decimam partem homer batus, et decimam partem homer ephi: iuxta mensuram homer sit aequa libratio eorum.
EZEK|45|12|Siclus autem viginti gera habeat; quinque sicli sint quinque, et decem sicli sint decem, et quinquaginta sint vobis mina.
EZEK|45|13|Haec est oblatio, quam offeratis: sextam partem ephi de gomor frumenti et sextam partem ephi de gomor hordei.
EZEK|45|14|Praeceptum quoque de oleo - batus est mensura olei C: decimam partem bati offeratis de choro - decem bati homer faciunt, quia decem bati implent chorum C.
EZEK|45|15|Et pecus unum de grege ducentorum, de pascuis irriguis Israel, in oblationem et in holocaustum et in pacifica ad expiandum pro eis, ait Dominus Deus.
EZEK|45|16|Omnis populus terrae tenebitur ad hanc oblationem principi in Israel;
EZEK|45|17|et super principem erunt holocausta et oblationes et libamina in diebus festis et in calendis et in sabbatis et in universis sollemnitatibus domus Israel; ipse faciet pro peccato et oblationem et holocaustum et pacifica ad expiandum pro domo Israel.
EZEK|45|18|Haec dicit Dominus Deus: In primo mense, una mensis, sumes vitulum de armento immaculatum et expiabis sanctuarium.
EZEK|45|19|Et tollet sacerdos de sanguine hostiae pro peccato et ponet in postibus domus et in quattuor angulis crepidinis altaris et in postibus portae atrii interioris.
EZEK|45|20|Et sic facies in septima mensis pro unoquoque, qui ignoravit et errore deceptus est, et expiabitis pro domo.
EZEK|45|21|In primo mense, quarta decima die mensis, erit vobis Paschae sollemnitas; septem diebus azyma comedentur.
EZEK|45|22|Et faciet princeps in die illa pro se et pro universo populo terrae vitulum pro peccato;
EZEK|45|23|et in septem dierum sollemnitate faciet holocaustum Domino septem vitulos et septem arietes immaculatos cotidie septem diebus et pro peccato hircum caprarum cotidie;
EZEK|45|24|et oblationem ephi per vitulum et ephi per arietem faciet et olei hin per singula ephi.
EZEK|45|25|Septimo mense, quinta decima die mensis, in sollemnitate faciet, sicut supra dicta sunt, per septem dies, tam pro peccato quam pro holocausto et in oblatione et in oleo.
EZEK|46|1|Haec dixit Dominus Deus: Porta atrii interioris, quae respicit ad orientem, erit clausa sex diebus, in quibus opus fit; die autem sabbati aperietur, sed et in die calendarum aperietur,
EZEK|46|2|et intrabit princeps per viam vestibuli portae deforis et stabit in poste portae, et facient sacerdotes holocaustum eius et pacifica eius, et adorabit super limen portae et egredietur; porta autem non claudetur usque ad vesperam.
EZEK|46|3|Et adorabit populus terrae ad ostium portae illius in sabbatis et in calendis coram Domino.
EZEK|46|4|Holocaustum autem hoc offeret princeps Domino: in die sabbati sex agnos immaculatos et arietem immaculatum
EZEK|46|5|et oblationem ephi per arietem, per agnos autem oblationem, quantum dederit manus eius, et olei hin per singula ephi;
EZEK|46|6|in die autem calendarum vitulum de armento immaculatum et sex agni et aries immaculati erunt
EZEK|46|7|et ephi per vitulum, ephi quoque per arietem faciet oblationem, per agnos autem sicut invenerit manus eius, et olei hin per singula ephi.
EZEK|46|8|Cumque ingressurus est princeps, per viam vestibuli portae ingrediatur et per eandem viam exeat.
EZEK|46|9|Et cum intrabit populus terrae in conspectu Domini in sollemnitatibus, qui ingreditur per portam aquilonis, ut adoret, egrediatur per viam portae meridianae; porro qui ingreditur per viam portae meridianae, egrediatur per viam portae aquilonis: non revertetur per viam portae, per quam ingressus est, sed e regione illius egredietur.
EZEK|46|10|Princeps autem in medio eorum cum ingredientibus ingredietur et cum egredientibus egredietur.
EZEK|46|11|Et in diebus festis et in sollemnitatibus erit oblatio ephi per vitulum et ephi per arietem, per agnos autem erit oblatio, quantum invenerit manus eius, et olei hin per singula ephi.
EZEK|46|12|Cum autem fecerit princeps spontaneum holocaustum aut pacifica voluntaria Domino, aperietur ei porta, quae respicit ad orientem, et faciet holocaustum suum et pacifica sua, sicut facere solet in die sabbati, et egredietur, claudeturque porta, postquam exierit.
EZEK|46|13|Et agnum anniculum immaculatum facies holocaustum cotidie Domino; semper mane facies illud.
EZEK|46|14|Et oblationem facies super eo mane mane sextam partem ephi, et de oleo tertiam partem hin, ut conspergatur simila; oblatio Domino, legitimum iuge atque perpetuum.
EZEK|46|15|Facient agnum et oblationem et oleum mane mane, holocaustum sempiternum.
EZEK|46|16|Haec dixit Dominus Deus: Si dederit princeps donum alicui de filiis suis de hereditate sua, filiorum suorum erit; possidebunt illud hereditarie.
EZEK|46|17|Si autem dederit legatum de hereditate sua uni servorum suorum, erit illius usque ad annum remissionis et revertetur ad principem; sola hereditas filiorum eius illorum erit.
EZEK|46|18|Et non accipiet princeps de hereditate populi, ut expellat eos de possessione eorum, sed de possessione sua hereditatem dabit filiis suis, ut non dispergatur populus meus unusquisque a possessione sua ".
EZEK|46|19|Et introduxit me per ingressum, qui erat ex latere portae, in exedras sacras sacerdotum, quae respiciebant ad aquilonem, et erat ibi locus in extrema parte vergens ad occidentem;
EZEK|46|20|et dixit ad me: " Iste est locus, ubi coquent sacerdotes pro delicto et pro peccato, ubi coquent oblationem, ut non efferant in atrium exterius, et sanctificetur populus ".
EZEK|46|21|Et eduxit me in atrium exterius et circumduxit me per quattuor angulos atrii, et ecce atriola singula per angulos atrii.
EZEK|46|22|In quattuor angulis atrii atriola inclusa quadraginta cubitorum per longum et triginta per latum: mensurae unius quattuor erant.
EZEK|46|23|Et paries per circuitum ambiens quattuor atriola, et culinae fabricatae erant subter parietes per gyrum.
EZEK|46|24|Et dixit ad me: "Hae sunt domus culinarum, in quibus coquent ministri domus Domini victimas populi ".
EZEK|47|1|Et convertit me ad portam domus, et ecce aquae egre diebantur subter limen domus ad orientem; facies enim domus respiciebat ad orientem, aquae autem descendebant a latere templi dextro a meridie altaris.
EZEK|47|2|Et eduxit me per viam portae aquilonis et convertit me ad viam foras ad portam exteriorem, quae respiciebat ad orientem; et ecce aquae exeuntes a latere dextro.
EZEK|47|3|Cum egrederetur vir ad orientem, qui habebat funiculum in manu sua, mensus est mille cubitos et traduxit me per aquam usque ad talos.
EZEK|47|4|Rursumque mensus est mille et traduxit me per aquam usque ad genua.
EZEK|47|5|Et mensus est mille et traduxit me per aquam usque ad renes. Et mensus est mille; torrens, quem non potui pertransire, quoniam intumuerant aquae, aquae ad natandum; torrens, qui non poterat transvadari.
EZEK|47|6|Et dixit ad me: " Certe vidisti, fili hominis "; et duxit me et convertit ad ripam torrentis.
EZEK|47|7|Cumque me convertissem, ecce in ripa torrentis ligna multa nimis ex utraque parte;
EZEK|47|8|et ait ad me: " Aquae istae, quae egrediuntur ad regionem orientalem et descendunt ad Arabam, intrabunt mare, aquas salsas, et sanabuntur aquae:
EZEK|47|9|et omnis anima vivens, quae movetur, quocumque venerit torrens, vivet, et erunt pisces multi satis, postquam venerint illuc aquae istae, et sanabuntur et vivent omnia, ad quae venerit torrens.
EZEK|47|10|Et stabunt super mare piscatores; ab Engaddi usque ad Engallim siccatio sagenarum erit; plurimae species erunt piscium eius, sicut pisces maris Magni, multitudinis nimiae.
EZEK|47|11|Palustria autem eius et stagna non sanabuntur, quia in salinas dabuntur.
EZEK|47|12|Et super torrentem orietur in ripis eius ex utraque parte omne lignum pomiferum; non defluet folium ex eo, et non deficiet fructus eius: per singulos menses afferet primitiva, quia aquae eius de sanctuario egredientur, et erunt fructus eius in cibum, et folia eius ad medicinam.
EZEK|47|13|Haec dicit Dominus Deus: Hic est terminus, in quo possidebitis terram in duodecim tribubus Israel, quia Ioseph duplicem funiculum habet;
EZEK|47|14|possidebitis autem eam, singuli aeque ut frater suus, super quam levavi manum meam, ut darem patribus vestris; et cadet terra haec vobis in possessionem.
EZEK|47|15|Hic est autem terminus terrae: ad plagam septentrionalem a mari Magno via Hethalon ad introitum Emath,
EZEK|47|16|Sedada, Berotha, Sabarim, quae est inter terminum Damasci et confinium Emath, usque ad Asarenon, quae est iuxta terminum Auran;
EZEK|47|17|erit ergo terminus a mari usque ad Asarenon, cum fines Damasci et fines Emath sint in aquilone; haec est plaga septentrionalis.
EZEK|47|18|Porro plaga orientalis de loco inter Auran et inter Damascum et in medio inter Galaad et terram Israel, Iordanis disterminans usque ad mare orientale, usque Thamar; haec est plaga orientalis.
EZEK|47|19|Plaga autem australis meridiana a Thamar usque ad aquas Meribathcades et torrentem usque ad mare Magnum; haec est plaga ad meridiem australis.
EZEK|47|20|Et plaga maris, mare Magnum a confinio per directum, donec venias Emath; haec est plaga maris.
EZEK|47|21|Et dividetis terram istam vobis per tribus Israel
EZEK|47|22|et mittetis eam in hereditatem, vobis et advenis, qui accesserint ad vos, qui genuerint filios in medio vestrum, et erunt vobis sicut indigenae inter filios Israel: vobiscum divident possessionem in medio tribuum Israel;
EZEK|47|23|in tribu autem quacumque fuerit advena, ibi dabitis possessionem illi, ait Dominus Deus.
EZEK|48|1|Et haec nomina tribuum: in finibus aquilonis iuxta viam Hethalon ad introitum Emath, Asarenon - fines Damasci ad aquilonem iuxta Emath - erit a plaga orientali usque ad mare, Dan pars una.
EZEK|48|2|Et iuxta terminum Dan a plaga orientali usque ad plagam maris, Aser una.
EZEK|48|3|Et iuxta terminum Aser a plaga orientali usque ad plagam maris, Nephthali una.
EZEK|48|4|Et iuxta terminum Nephthali a plaga orientali usque ad plagam maris, Manasse una.
EZEK|48|5|Et iuxta terminum Manasse a plaga orientali usque ad plagam maris, Ephraim una.
EZEK|48|6|Et iuxta terminum Ephraim a plaga orientali usque ad plagam maris, Ruben una.
EZEK|48|7|Et iuxta terminum Ruben a plaga orientali usque ad plagam maris, Iudae una.
EZEK|48|8|Et iuxta terminum Iudae a plaga orientali usque ad plagam maris oblatio, quam separabitis viginti quinque milibus latitudinis et longitudinis, sicuti singulae partes a plaga orientali usque ad plagam maris; et erit sanctuarium in medio eius.
EZEK|48|9|Oblatio, quam separabitis Domino, longitudo viginti quinque milibus et latitudo viginti milibus.
EZEK|48|10|His autem est oblatio sacra: sacerdotibus, ad aquilonem viginti quinque milia et ad mare latitudinis decem milia et ad orientem latitudinis decem milia et ad meridiem longitudinis viginti quinque milia; et erit sanctuarium Domini in medio eius.
EZEK|48|11|Sacerdotibus consecratis erit, filiis Sadoc, qui custodierunt caeremonias meas et non erraverunt, cum errarent filii Israel, sicut erraverunt Levitae.
EZEK|48|12|Et erit eis oblatio de oblatione terrae sanctum sanctorum iuxta terminum Levitarum;
EZEK|48|13|sed et Levitis similiter secundum fines sacerdotum, viginti quinque milia longitudinis et latitudinis decem milia, totum in longitudine viginti et quinque milia et in latitudine viginti milia;
EZEK|48|14|et non venumdabunt ex eo neque mutabunt, neque transferetur oblatio terrae, quia sanctificata est Domino.
EZEK|48|15|Quinque milia autem, quae supersunt in latitudine per viginti quinque milia, profana erunt urbi in habitaculum et in pascua, et erit civitas in medio eius.
EZEK|48|16|Et hae mensurae eius: ad plagam septentrionalem quingenti et quattuor milia et ad plagam meridianam quingenti et quattuor milia et ad plagam orientalem quingenti et quattuor milia et ad plagam occidentalem quingenti et quattuor milia.
EZEK|48|17|Erunt autem pascua civitatis ad aquilonem ducenti quinquaginta et ad meridiem ducenti quinquaginta et ad orientem ducenti quinquaginta et ad mare ducenti quinquaginta.
EZEK|48|18|Quod autem reliquum fuerit in longitudine iuxta oblationem sacram, decem milia ad orientem et decem milia ad occidentem, erunt iuxta oblationem sacram, et erunt fruges eius in panem his, qui serviunt civitati.
EZEK|48|19|Servientes autem civitati operabuntur ex omnibus tribubus Israel.
EZEK|48|20|Tota oblatio viginti quinque milium, per viginti quinque milia: in quadrum; separabitis oblationem sacram una cum possessione civitatis.
EZEK|48|21|Quod autem reliquum fuerit, principis erit, ex utraque parte oblationis sacrae et possessionis civitatis, e regione viginti quinque milium oblationis usque ad terminum orientalem, sed et ad mare e regione viginti quinque milium usque ad terminum maris secundum partes tribuum, principis erit. Et erit oblatio sacra et sanctuarium templi in medio eius,
EZEK|48|22|segregata a possessione Levitarum et a possessione civitatis in medio partium principis: inter terminum Iudae et inter terminum Beniamin erit possessio principis.
EZEK|48|23|Et reliquis tribubus: a plaga orientali usque ad plagam occidentalem, Beniamin una.
EZEK|48|24|Et iuxta terminum Beniamin a plaga orientali usque ad plagam occidentalem, Simeon una.
EZEK|48|25|Et iuxta terminum Simeonis a plaga orientali usque ad plagam occidentalem, Issachar una.
EZEK|48|26|Et iuxta terminum Issachar a plaga orientali usque ad plagam occidentalem, Zabulon una.
EZEK|48|27|Et iuxta terminum Zabulon a plaga orientali usque ad plagam maris, Gad una.
EZEK|48|28|Et iuxta terminum Gad ad plagam austri in meridiem, erit finis de Thamar usque ad aquas Meribathcades, ad torrentem usque ad mare Magnum.
EZEK|48|29|Haec est terra, quam mittetis in sortem tribubus Israel, et hae partitiones earum, ait Dominus Deus.
EZEK|48|30|Et hi egressus civitatis: a plaga septentrionali, cuius mensura quingenti et quattuor milia,
EZEK|48|31|portae civitatis in nominibus tribuum Israel: portae tres a septentrione, porta Ruben una, porta Iudae una, porta Levi una.
EZEK|48|32|Et ad plagam orientalem quingentorum et quattuor milium, portae tres: porta Ioseph una, porta Beniamin una, porta Dan una.
EZEK|48|33|Et ad plagam meridianam, cuius mensura quingenti et quattuor milia, portae tres: porta Simeonis una, porta Issachar una, porta Zabulon una.
EZEK|48|34|Et ad plagam occidentalem quingentorum et quattuor milium, portae tres: porta Gad una, porta Aser una, porta Nephthali una.
EZEK|48|35|Per circuitum decem et octo milia, et nomen civitatis ex illa die: Dominus ibidem ".
DAN|1|1|Anno tertio regni Ioachim regis Iudae venit Nabuchodonosor rex Babylonis Ierusalem et obsedit eam;
DAN|1|2|et tradidit Dominus in manu eius Ioachim regem Iudae et partem vasorum domus Dei, et asportavit ea in terram Sennaar in domum deorum suorum et vasa intulit in domum thesauri deorum suorum.
DAN|1|3|Et ait rex Asfanaz praeposito eunuchorum suorum, ut introduceret de filiis Israel et de semine regio et tyrannorum
DAN|1|4|pueros, in quibus nulla esset macula, decoros forma et eruditos omni sapientia, cautos scientia et doctos disciplina, et qui possent stare in palatio regis, et ut docerent eos litteras et linguam Chaldaeorum.
DAN|1|5|Et constituit eis rex annonam per singulos dies de cibis suis et de vino, unde bibebat ipse, ut enutriti tribus annis postea starent in conspectu regis.
DAN|1|6|Fuerunt ergo inter eos de filiis Iudae Daniel, Ananias, Misael et Azarias.
DAN|1|7|Et imposuit eis praepositus eunuchorum nomina: Danieli Baltassar et Ananiae Sedrac, Misaeli Misac et Azariae Abdenago.
DAN|1|8|Proposuit autem Daniel in corde suo, ne pollueretur de mensa regis neque de vino potus eius, et rogavit eunuchorum praepositum, ne contaminaretur.
DAN|1|9|Dedit autem Deus Danieli gratiam et misericordiam in conspectu principis eunuchorum;
DAN|1|10|et ait princeps eunuchorum ad Daniel: " Timeo ego dominum meum regem, qui constituit vobis cibum et potum; qui si viderit vultus vestros macilentiores prae ceteris adulescentibus coaevis vestris, condemnabitis caput meum regi ".
DAN|1|11|Et dixit Daniel ad custodem, quem constituerat princeps eunuchorum super Daniel, Ananiam, Misael et Azariam:
DAN|1|12|" Tenta nos, obsecro, servos tuos diebus decem, et dentur nobis legumina ad vescendum et aqua ad bibendum;
DAN|1|13|et videantur in conspectu tuo vultus nostri et vultus puerorum, qui vescuntur cibo regio, et, sicut videris, facies cum servis tuis ".
DAN|1|14|Qui, audito sermone huiuscemodi, tentavit eos diebus decem.
DAN|1|15|Post dies autem decem apparuerunt vultus eorum meliores et corpulentiores prae omnibus pueris, qui vescebantur cibo regio.
DAN|1|16|Porro custos tollebat cibaria et vinum potus eorum dabatque eis legumina.
DAN|1|17|Quattuor autem pueris his dedit Deus scientiam et disciplinam in omni scriptura et sapientia, Danieli autem intellegentiam omnium visionum et somniorum.
DAN|1|18|Completis itaque diebus, post quos dixerat rex, ut introducerentur, introduxit eos praepositus eunuchorum in conspectu Nabuchodonosor.
DAN|1|19|Cumque locutus eis fuisset rex, non sunt inventi de universis tales ut Daniel, Ananias, Misael et Azarias; et steterunt in conspectu regis.
DAN|1|20|Et omne verbum sapientiae et intellectus, quod sciscitatus est ab eis, rex invenit in eis decuplum super cunctos hariolos et magos, qui erant in universo regno eius.
DAN|1|21|Fuit autem Daniel usque ad annum primum Cyri regis.
DAN|2|1|In anno secundo regni Nabu chodonosor vidit Nabuchodo nosor somnium, et conterritus est spiritus eius, et somnus eius fugit ab eo.
DAN|2|2|Praecepit autem rex, ut convocarentur harioli et magi et malefici et Chaldaei et indicarent regi somnia sua; qui cum venissent, steterunt coram rege.
DAN|2|3|Et dixit ad eos rex: " Vidi somnium, et spiritus meus conterritus est, ut intellegat somnium ".
DAN|2|4|Responderuntque Chaldaei regi Aramaice: " Rex, in sempiternum vive! Dic somnium servis tuis, et interpretationem eius indicabimus ".
DAN|2|5|Et respondens rex ait Chaldaeis: " Sermo recessit a me. Nisi indicaveritis mihi somnium et coniecturam eius, in frusta concidemini, et domus vestrae in sterquilinium ponentur;
DAN|2|6|si autem somnium et coniecturam eius narraveritis, praemia et dona et honorem multum accipietis a me. Somnium igitur et interpretationem eius indicate mihi ".
DAN|2|7|Responderunt secundo atque dixerunt: " Rex somnium dicat servis suis, et interpretationem illius indicabimus ".
DAN|2|8|Respondit rex et ait: " Certe novi quia tempus redimitis, scientes quod recesserit a me sermo.
DAN|2|9|Si ergo somnium non indicaveritis mihi, una est de vobis sententia. Et verbum fallax et deceptione plenum composuistis, ut loquamini mihi, donec tempus pertranseat; somnium itaque dicite mihi, ut sciam quod interpretationem eius loquamini mihi ".
DAN|2|10|Respondentes ergo Chaldaei coram rege dixerunt: " Non est homo super terram qui sermonem regis possit indicare; quapropter neque regum quisquam magnus et potens verbum huiuscemodi sciscitatur ab omni hariolo et mago et Chaldaeo.
DAN|2|11|Sermo enim, quem tu quaeris, rex, gravis est, nec reperietur quisquam qui indicet illum in conspectu regis, exceptis diis, quorum non est cum hominibus conversatio ".
DAN|2|12|Quo audito, rex in furore et in ira magna praecepit, ut perirent omnes sapientes Babylonis.
DAN|2|13|Et egressa sententia, ut sapientes interficerentur, quaerebantur Daniel et socii eius, ut perirent.
DAN|2|14|Tunc Daniel interrogavit cum consilio et prudentia Arioch, principem militiae regis, qui egressus fuerat ad interficiendos sapientes Babylonis;
DAN|2|15|respondens dixit ad Arioch, qui a rege potestatem acceperat, quam ob causam tam crudelis sententia a facie esset regis egressa. Cum ergo rem indicasset Arioch Danieli,
DAN|2|16|Daniel ingressus rogavit regem, ut tempus daret sibi ad solutionem indicandam regi;
DAN|2|17|et ingressus est domum suam Ananiaeque, Misaeli et Azariae sociis suis indicavit negotium,
DAN|2|18|ut quaererent misericordiam a facie Dei caeli super sacramento isto et non perirent Daniel et socii eius cum ceteris sapientibus Babylonis.
DAN|2|19|Tunc Danieli per visionem nocte mysterium revelatum est, et benedixit Daniel Deo caeli
DAN|2|20|et locutus Daniel ait: Sit nomen Dei benedictuma saeculo et usque in saeculum,quia sapientia et fortitudo eius sunt;
DAN|2|21|et ipse mutat tempora et aetates,transfert atque constituit reges,dat sapientiam sapientibuset scientiam intellegentibus disciplinam:
DAN|2|22|ipse revelat profunda et absconditaet novit in tenebris constituta,et lux cum eo inhabitat,
DAN|2|23|Tibi, Deus patrum meorum, confiteor teque laudo,quia sapientiam et fortitudinem dedisti mihiet nunc ostendisti mihi, quae rogavimus te,quia sermonem regis aperuisti nobis ".
DAN|2|24|Propterea Daniel, ingressus ad Arioch, quem constituerat rex, ut perderet sapientes Babylonis, sic ei locutus est: " Sapientes Babylonis ne perdas; introduc me in conspectu regis et solutionem regi enarrabo ".
DAN|2|25|Tunc Arioch festinus introduxit Danielem ad regem et dixit ei: " Inveni hominem de filiis transmigrationis Iudae, qui solutionem regi annuntiet ".
DAN|2|26|Respondit rex et dixit Danieli, cuius nomen erat Baltassar: " Putasne vere potes mihi indicare somnium, quod vidi, et interpretationem eius?".
DAN|2|27|Et respondens Daniel coram rege ait: " Mysterium, quod rex interrogat, sapientes, magi et harioli et haruspices non queunt indicare regi;
DAN|2|28|sed est Deus in caelo revelans mysteria, qui indicavit tibi, rex Nabuchodonosor, quae ventura sunt in novissimis temporibus. Somnium tuum et visiones capitis tui in cubili tuo huiuscemodi sunt:
DAN|2|29|Tu, rex, cogitare coepisti in strato tuo quid esset futurum post haec; et, qui revelat mysteria, ostendit tibi, quae ventura sunt.
DAN|2|30|Mihi quoque non in sapientia, quae est in me plus quam in cunctis viventibus, sacramentum hoc revelatum est, sed ut interpretatio regi manifesta fieret, et cogitationes mentis tuae scires.
DAN|2|31|Tu, rex, videbas, et ecce statua una grandis: statua illa magna et statura sublimis stabat contra te, et intuitus eius erat terribilis.
DAN|2|32|Huius statuae caput ex auro optimo erat, pectus autem et brachia de argento, porro venter et femora ex aere,
DAN|2|33|tibiae autem ferreae, pedum quaedam pars erat ferrea, quaedam autem fictilis.
DAN|2|34|Videbas ita, donec abscissus est lapis sine manibus et percussit statuam in pedibus eius ferreis et fictilibus et comminuit eos;
DAN|2|35|tunc contrita sunt pariter ferrum, testa, aes, argentum et aurum, et fuerunt quasi folliculus ex areis aestivis, et rapuit ea ventus, nullusque locus inventus est eis; lapis autem, qui percusserat statuam, factus est mons magnus et implevit universam terram.
DAN|2|36|Hoc est somnium; interpretationem quoque eius dicemus coram te, rex.
DAN|2|37|Tu rex regum es, et Deus caeli regnum et fortitudinem et imperium et gloriam dedit tibi;
DAN|2|38|et omnia, in quibus habitant filii hominum et bestiae agri volucresque caeli, dedit in manu tua et te dominum universorum constituit: tu es caput aureum.
DAN|2|39|Et post te consurget regnum aliud minus te et regnum tertium aliud aereum, quod imperabit universae terrae.
DAN|2|40|Et regnum quartum erit robustum velut ferrum; quomodo ferrum comminuit et domat omnia, et sicut ferrum comminuens conteret et comminuet omnia haec.
DAN|2|41|Porro quia vidisti pedum et digitorum partem testae figuli et partem ferream, regnum divisum erit; et robur ferri erit ei, secundum quod vidisti ferrum mixtum testae ex luto.
DAN|2|42|Et digitos pedum ex parte ferreos et ex parte fictiles, ex parte regnum erit solidum et ex parte contritum.
DAN|2|43|Quod autem vidisti ferrum mixtum testae ex luto, commiscebuntur quidem humano semine, sed non adhaerebunt sibi, sicuti ferrum misceri non potest testae.
DAN|2|44|In diebus autem regnorum illorum suscitabit Deus caeli regnum, quod in aeternum non dissipabitur, et regnum populo alteri non tradetur: comminuet et consumet universa regna haec, et ipsum stabit in aeternum.
DAN|2|45|Secundum quod vidisti quod de monte abscisus est lapis sine manibus et comminuit testam et ferrum et aes et argentum et aurum, Deus magnus ostendit regi, quae ventura sunt postea; et verum est somnium et fidelis interpretatio eius ".
DAN|2|46|Tunc rex Nabuchodonosor cecidit in faciem suam et Danielem adoravit et hostias et incensum praecepit, ut sacrificarent ei.
DAN|2|47|Loquens ergo rex ait Danieli: " Vere Deus vester Deus deorum est et Dominus regum et revelans mysteria, quoniam potuisti aperire sacramentum hoc ".
DAN|2|48|Tunc rex Danielem in sublime extulit et munera multa et magna dedit ei et constituit eum principem super omnes provincias Babylonis et principem praefectorum super cunctos sapientes Babylonis.
DAN|2|49|Daniel autem postulavit a rege et constituit super opera provinciae Babylonis Sedrac, Misac et Abdenago; ipse autem Daniel erat in foribus regis.
DAN|3|1|Nabuchodonosor rex fecit sta tuam auream altitudine cubito rum sexaginta, latitudine cubitorum sex; et statuit eam in campo Dura in provincia Babylonis.
DAN|3|2|Itaque Nabuchodonosor rex misit ad congregandos satrapas, magistratus et iudices, duces et tyrannos et praefectos omnesque principes provinciarum, ut convenirent ad dedicationem statuae, quam erexerat Nabuchodonosor rex.
DAN|3|3|Tunc congregati sunt satrapae, magistratus et iudices, duces et tyranni et optimates, qui erant in potestatibus constituti, et universi principes provinciarum ad dedicationem statuae, quam erexerat Nabuchodonosor rex. Stabant autem in conspectu statuae, quam posuerat Nabuchodonosor,
DAN|3|4|et praeco clamabat valenter: " Vobis dicitur, populi, tribus et linguae:
DAN|3|5|in hora, qua audieritis sonitum tubae et fistulae et citharae, sambucae et psalterii et symphoniae et universi generis musicorum, cadentes adorate statuam auream, quam constituit Nabuchodonosor rex.
DAN|3|6|Si quis autem non prostratus adoraverit, eadem hora mittetur in fornacem ignis ardentis ".
DAN|3|7|Post haec igitur, statim ut audierunt omnes populi sonitum tubae, fistulae et citharae, sambucae et psalterii et symphoniae et omnis generis musicorum, cadentes omnes populi tribus et linguae adoraverunt statuam auream, quam constituerat Nabuchodonosor rex.
DAN|3|8|Statimque et in ipso tempore accedentes viri Chaldaei accusaverunt Iudaeos
DAN|3|9|dixeruntque Nabuchodonosor regi: " Rex, in aeternum vive!
DAN|3|10|Tu, rex, posuisti decretum, ut omnis homo, qui audierit sonitum tubae, fistulae et citharae, sambucae et psalterii et symphoniae et universi generis musicorum, prosternat se et adoret statuam auream;
DAN|3|11|si quis autem non procidens adoraverit, mittetur in fornacem ignis ardentis.
DAN|3|12|Sunt ergo viri Iudaei, quos constituisti super opera provinciae Babylonis, Sedrac, Misac et Abdenago; viri isti te, rex, non honorant: deos tuos non colunt et statuam auream, quam erexisti, non adorant ".
DAN|3|13|Tunc Nabuchodonosor in furore et in ira praecepit, ut adducerentur Sedrac, Misac et Abdenago; tunc viri illi adducti sunt in conspectu regis.
DAN|3|14|Pronuntiansque Nabuchodonosor rex ait eis: " Verene, Sedrac, Misac et Abdenago, deos meos non colitis et statuam auream, quam constitui, non adoratis?
DAN|3|15|Numquid estis nunc parati, quacumque hora audieritis sonitum tubae, fistulae, citharae, sambucae, psalterii et symphoniae omnisque generis musicorum, prosternere vos et adorare statuam, quam feci? Quod si non adoraveritis, eadem hora mittemini in fornacem ignis ardentis; et quis est deus, qui eripiat vos de manu mea? ".
DAN|3|16|Respondentes Sedrac, Misac et Abdenago dixerunt regi Nabuchodonosor: " Non oportet nos de hac re respondere tibi:
DAN|3|17|Si enim Deus noster, quem colimus, potest eripere nos de camino ignis ardentis, et de manu tua, rex, liberabit.
DAN|3|18|Quod si noluerit, notum sit tibi, rex, quia deos tuos non colimus et statuam auream, quam erexisti, non adoramus ".
DAN|3|19|Tunc Nabuchodonosor repletus est furore, et aspectus faciei illius immutatus est super Sedrac, Misac et Abdenago; et respondens praecepit, ut succenderetur fornax septuplum quam succendi consueverat;
DAN|3|20|et viris fortissimis de exercitu suo iussit, ut ligarent Sedrac, Misac et Abdenago et mitterent eos in fornacem ignis ardentis;
DAN|3|21|et confestim viri illi vincti, cum bracis suis et tiaris et calceamentis et vestibus missi sunt in medium fornacis ignis ardentis;
DAN|3|22|itaque, quia iussio regis urgebat, et fornax succensa erat nimis, viros illos, qui miserant Sedrac, Misac et Abdenago, interfecit flamma ignis.
DAN|3|23|Viri autem tres, Sedrac, Misac et Abdenago, ceciderunt in medio camino ignis ardentis colligati.Quae sequuntur in Hebraeis voluminibus non repperi).
DAN|3|24|Et ambulabant in medio flammae laudantes Deum et benedicentes Domino.
DAN|3|25|Stans autem Azarias oravit sic aperiensque os suum in medio ignis ait:
DAN|3|26|" Benedictus es, Domine, Deus patrum nostrorum,et laudabilis et gloriosum nomen tuum in saecula,
DAN|3|27|quia iustus es in omnibus, quae fecisti nobis,et universa opera tua vera, et viae tuae rectae,et omnia iudicia tua veritas.
DAN|3|28|Iudicia enim vera fecistiiuxta omnia, quae induxisti super noset super civitatem sanctam patrum nostrorum Ierusalem,quia in veritate et in iudicio induxisti omnia haecpropter peccata nostra.
DAN|3|29|Peccavimus enim et inique egimus recedentes a teet deliquimus in omnibus;
DAN|3|30|et praecepta tua non audivimusnec observavimusnec fecimus, sicut praeceperas nobis,ut bene nobis esset.
DAN|3|31|Omnia ergo, quae induxisti super nos,et universa, quae fecisti nobis,vero iudicio fecisti;
DAN|3|32|et tradidisti nos in manibus inimicorum nostroruminiquorum et pessimorum praevaricatorumqueet regi iniusto et pessimo ultra omnem terram.
DAN|3|33|Et nunc non possumus aperire os;confusio et opprobrium facta suntservis tuis et his, qui colunt te.
DAN|3|34|Ne, quaesumus, tradas nos in perpetuumpropter nomen tuumet ne dissipes testamentum tuum
DAN|3|35|neque auferas misericordiam tuam a nobispropter Abraham dilectum tuumet Isaac servum tuumet Israel sanctum tuum,
DAN|3|36|quibus dixistiquod multiplicares semen eorum sicut stellas caeliet sicut arenam, quae est in litore maris;
DAN|3|37|quia, Domine,imminuti sumus plus quam omnes gentessumusque humiles in universa terrahodie propter peccata nostra;
DAN|3|38|et non est in tempore hocprinceps et propheta et duxneque holocaustum neque sacrificiumneque oblatio neque incensumneque locus primitiarum coram te,ut possimus invenire misericordiam;
DAN|3|39|sed in anima contrita et spiritu humilitatis suscipiamursicut in holocausto arietum et taurorum
DAN|3|40|et sicut in milibus agnorum pinguium;sic fiat sacrificium nostrum in conspectu tuo hodie,et perfice subsequentes te,quoniam non est confusio confidentibus in te.
DAN|3|41|Et nunc sequimur te in toto cordeet timemus te et quaerimus faciem tuam;
DAN|3|42|ne confundas nos,sed fac nobiscum iuxta mansuetudinem tuamet secundum multitudinem misericordiae tuae
DAN|3|43|et erue nos in mirabilibus tuiset da gloriam nomini tuo, Domine.
DAN|3|44|Et confundantur omnes, qui ostendunt servis tuis mala;confundantur absque ulla potentia,et robur eorum conteratur.
DAN|3|45|Sciant quia tu es Dominus,Deus solus et gloriosus super orbem terrarum ".
DAN|3|46|Et non cessabant, qui immiserant eos, ministri regis succendere fornacem naphta et stuppa et pice et malleolis,
DAN|3|47|et effundebatur flamma super fornacem cubitis quadraginta novem
DAN|3|48|et erupit et incendit, quos repperit iuxta fornacem de Chaldaeis.
DAN|3|49|Angelus autem Domini descendit cum Azaria et sociis eius in fornacem et excussit flammam ignis de fornace
DAN|3|50|et fecit medium fornacis quasi ventum roris flantem; et non tetigit eos omnino ignis neque contristavit nec quidquam molestiae intulit.
DAN|3|51|Tunc hi tres, quasi ex uno ore, laudabant et glorificabant et benedicebant Deo in fornace dicentes:
DAN|3|52|" Benedictus es, Domine, Deus patrum nostrorum,et laudabilis et superexaltatus in saecula;et benedictum nomen gloriae tuae sanctumet superlaudabile et superexaltatum in saecula.
DAN|3|53|Benedictus es in templo sanctae gloriae tuaeet superlaudabilis et supergloriosus in saecula.
DAN|3|54|Benedictus es in throno regni tuiet superlaudabilis et superexaltatus in saecula.
DAN|3|55|Benedictus es, qui intueris abyssos sedens super cherubim,et laudabilis et superexaltatus in saecula.
DAN|3|56|Benedictus es in firmamento caeliet laudabilis et gloriosus in saecula.
DAN|3|57|Benedicite, omnia opera Domini, Domino,laudate et superexaltate eum in saecula.
DAN|3|58|Benedicite, caeli, Domino,laudate et superexaltate eum in saecula.
DAN|3|59|Benedicite, angeli Domini, Domino,laudate et superexaltate eum in saecula.
DAN|3|60|Benedicite, aquae omnes, quae super caelos sunt, Domino,laudate et superexaltate eum in saecula.
DAN|3|61|Benedicat omnis virtus Domino,laudate et superexaltate eum in saecula.
DAN|3|62|Benedicite, sol et luna, Domino,laudate et superexaltate eum in saecula.
DAN|3|63|Benedicite, stellae caeli, Domino,laudate et superexaltate eum in saecula.
DAN|3|64|Benedicite, omnis imber et ros, Domino,laudate et superexaltate eum in saecula.
DAN|3|65|Benedicite, omnes venti, Domino,laudate et superexaltate eum in saecula.
DAN|3|66|Benedicite, ignis et aestus, Domino,laudate et superexaltate eum in saecula.
DAN|3|67|Benedicite, frigus et aestus, Domino,laudate et superexaltate eum in saecula.
DAN|3|68|Benedicite, rores et pruina, Domino,laudate et superexaltate eum in saecula.
DAN|3|69|Benedicite, gelu et frigus, Domino,laudate et superexaltate eum in saecula.
DAN|3|70|Benedicite, glacies et nives, Domino,laudate et superexaltate eum in saecula.
DAN|3|71|Benedicite, noctes et dies, Domino,laudate et superexaltate eum in saecula.
DAN|3|72|Benedicite, lux et tenebrae, Domino,laudate et superexaltate eum in saecula.
DAN|3|73|Benedicite, fulgura et nubes, Domino,laudate et superexaltate eum in saecula.
DAN|3|74|Benedicat terra Dominum,laudet et superexaltet eum in saecula.
DAN|3|75|Benedicite, montes et colles, Domino,laudate et superexaltate eum in saecula.
DAN|3|76|Benedicite, universa germinantia in terra, Domino,laudate et superexaltate eum in saecula.
DAN|3|77|Benedicite, maria et flumina, Domino,laudate et superexaltate eum in saecula.
DAN|3|78|Benedicite, fontes, Domino,laudate et superexaltate eum in saecula.
DAN|3|79|Benedicite, cete et omnia quae moventur in aquis, Domino,laudate et superexaltate eum in saecula.
DAN|3|80|Benedicite, omnes volucres caeli, Domino,laudate et superexaltate eum in saecula.
DAN|3|81|Benedicite, omnes bestiae et pecora, Domino,laudate et superexaltate eum in saecula.
DAN|3|82|Benedicite, filii hominum, Domino,laudate et superexaltate eum in saecula.
DAN|3|83|Benedic, Israel, Domino,laudate et superexaltate eum in saecula.
DAN|3|84|Benedicite, sacerdotes Domini, Domino,laudate et superexaltate eum in saecula.
DAN|3|85|Benedicite, servi Domini, Domino,laudate et superexaltate eum in saecula.
DAN|3|86|Benedicite, spiritus et animae iustorum, Domino,laudate et superexaltate eum in saecula.
DAN|3|87|Benedicite, sancti et humiles corde, Domino,laudate et superexaltate eum in saecula.
DAN|3|88|Benedicite, Anania, Azaria, Misael, Domino,laudate et superexaltate eum in saecula;quia eruit nos de inferno et salvos fecit de manu mortiset liberavit nos de medio fornacis ardentis flammaeet de medio ignis eruit nos.
DAN|3|89|Confitemini Domino, quoniam bonus,quoniam in saeculum misericordia eius.
DAN|3|90|Benedicite, omnes, qui timetis Dominum, Deo deorum;laudate et confitemini ei, quia in saecula misericordia eius ".Hucusque non habetur in Hebraeo et, quae posuimus, de Theodotionis editione translata sunt).
DAN|3|91|24 Tunc Nabuchodonosor rex obstupuit et surrexit propere; respondens ait optimatibus suis: " Nonne tres viros misimus in medium ignis compeditos?". Qui respondentes dixerunt regi: " Vere, rex ".
DAN|3|92|25 Respondit et ait: " Ecce ego video viros quattuor solutos et ambulantes in medio ignis, et nihil corruptionis in eis est, et species quarti similis filio deorum ".
DAN|3|93|26 Tunc accessit Nabuchodonosor ad ostium fornacis ignis ardentis et ait: " Sedrac, Misac et Abdenago, servi Dei excelsi, egredimini et venite. Statimque egressi sunt Sedrac, Misac et Abdenago de medio ignis.
DAN|3|94|27 Et congregati satrapae, magistratus et iudices et potentes regis contemplabantur viros illos, quoniam nihil potestatis habuisset ignis in corporibus eorum, et capillus capitis eorum non esset adustus, et sarabara eorum non fuissent immutata, et odor ignis non transisset per eos.
DAN|3|95|28 Et erumpens Nabuchodonosor ait: " Benedictus Deus eorum, Sedrac, Misac et Abdenago, qui misit angelum suum et eruit servos suos, qui crediderunt in eo, et verbum regis immutaverunt et tradiderunt corpora sua, ne servirent et ne adorarent omnem deum, excepto Deo suo.
DAN|3|96|29 A me ergo positum est decretum, ut omnis populus, tribus et lingua quaecumque locuta fuerit blasphemiam contra Deum Sedrac, Misac et Abdenago, in frusta concidatur, et domus eius in sterquilinium fiat, eo quod non est Deus alius, qui possit ita salvare ".
DAN|3|97|30 Tunc rex promovit Sedrac, Misac et Abdenago in provincia Babylonis.
DAN|3|98|31 Nabuchodonosor rex omnibus populis, gentibus et linguis, quae habitant in universa terra: " Pax vobis multiplicetur.
DAN|3|99|32 Signa et mirabilia, quae fecit apud me Deus excelsus, placuit mihi praedicare:
DAN|3|100|33 Signa eius quam magna sunt,et mirabilia eius quam fortia!Et regnum eius regnum sempiternum,et potestas eius in generationem et generationem ".
DAN|4|1|Ego Nabuchodonosor quietus eram in domo mea et florens in palatio meo;
DAN|4|2|somnium vidi, quod perterruit me, et cogitationes in stratu meo et visiones capitis mei conturbaverunt me.
DAN|4|3|Et per me propositum est decretum, ut introducerentur in conspectu meo cuncti sapientes Babylonis, ut solutionem somnii indicarent mihi.
DAN|4|4|Tunc ingrediebantur harioli, magi, Chaldaei et haruspices; et somnium narravi in conspectu eorum, et solutionem eius non indicaverunt mihi;
DAN|4|5|donec denique ingressus est in conspectu meo Daniel, cui nomen Baltassar secundum nomen dei mei et qui habet spiritum deorum sanctorum in semetipso. Et somnium coram ipso locutus sum:
DAN|4|6|Baltassar, princeps hariolorum, quem ego scio quod spiritum deorum sanctorum habeas in te, et omne sacramentum non est impossibile tibi, visiones somnii mei, quas vidi, et solutionem eius narra.
DAN|4|7|Visio capitis mei in cubili meo:Videbam, et ecce arbor in medio terrae,et altitudo eius nimia.
DAN|4|8|Magna arbor et fortis,et proceritas eius contingens caelum;aspectus illius erat usque ad terminos universae terrae.
DAN|4|9|Folia eius pulcherrima,et fructus eius nimius,et esca universorum in ea.Subter eam habitabant bestiae agri,et in ramis eius conversabantur volucres caeli,et ex ea vescebatur omnis caro.
DAN|4|10|Videbam in visione capitis mei super stratum meum,et ecce vigil et sanctus de caelo descendit.
DAN|4|11|Clamavit fortiter et sic ait:Succidite arborem et praecidite ramos eius,excutite folia eius et dispergite fructus eius.Fugiant bestiae de sub ea,et volucres de ramis eius.
DAN|4|12|Verumtamen germen radicum eius in terra siniteet in vinculo ferreo et aereo in herbis agri,et rore caeli tingatur,et cum feris pars eius in herba terrae.
DAN|4|13|Cor eius ab humano commutetur,et cor ferae detur ei,et septem tempora mutentur super eum.
DAN|4|14|In sententia vigilum decretum est,et sermo sanctorum petitio,ut cognoscant viventesquoniam dominatur Excelsus in regno hominumet, cuicumque voluerit, dabit illudet humillimum hominem constituet super eo".
DAN|4|15|Hoc somnium vidi ego rex Nabuchodonosor. Tu ergo, Baltassar, interpretationem narra, quia omnes sapientes regni mei non queunt solutionem edicere mihi; tu autem potes, quia spiritus deorum sanctorum in te est ".
DAN|4|16|Tunc Daniel, cuius nomen Baltassar, obstupuit quasi una hora, et cogitationes eius conturbabant eum. Respondens autem rex ait: " Baltassar, somnium et interpretatio eius non conturbent te ". Respondit Baltassar et dixit: " Domine mi, somnium his, qui te oderunt, et interpretatio eius hostibus tuis sit.
DAN|4|17|Arborem, quam vidisti sublimem atque robustam, cuius altitudo pertingit ad caelum, et aspectus illius in omnem terram,
DAN|4|18|et rami eius pulcherrimi, et fructus eius nimius, et esca omnium in ea, subter eam habitantes bestiae agri, et in ramis eius commorantes aves caeli,
DAN|4|19|tu es, rex, qui magnificatus es et invaluisti, et magnitudo tua crevit et pervenit usque ad caelum, et potestas tua in terminos terrae.
DAN|4|20|Quod autem vidit rex vigilem et sanctum descendere de caelo et dicere: Succidite arborem et dissipate illam; attamen germen radicum eius in terra dimittite, et vinculo ferreo et aereo in herbis agri, et rore caeli conspergatur, et cum feris sit pars eius, donec septem tempora mutentur super eum",
DAN|4|21|haec est interpretatio, rex, et sententia Altissimi, quae pervenit super dominum meum regem:
DAN|4|22|et eicient te ab hominibus, et cum bestiis feris erit habitatio tua, et fenum ut boves comedes et rore caeli infunderis; septem quoque tempora mutabuntur super te, donec scias quod dominetur Excelsus super regnum hominum et, cuicumque voluerit, det illud.
DAN|4|23|Quod autem praeceperunt, ut relinqueretur germen radicum eius, id est arboris, regnum tuum tibi manebit, postquam cognoveris potestatem caeli.
DAN|4|24|Quam ob rem, rex, consilium meum placeat tibi, et peccata tua eleemosynis redime et iniquitates tuas misericordiis pauperum; sic longitudo erit prosperitati tuae ".
DAN|4|25|Omnia haec venerunt super Nabuchodonosor regem.
DAN|4|26|Post finem mensium duodecim in palatio regni Babylonis deambulabat;
DAN|4|27|responditque rex et ait: " Nonne haec est Babylon magna, quam ego aedificavi in domum regni, in robore fortitudinis meae et in gloria decoris mei? ".
DAN|4|28|Cum adhuc sermo esset in ore regis, vox de caelo ruit: " Tibi dicitur, Nabuchodonosor rex: Regnum tuum transiit a te,
DAN|4|29|et ab hominibus te eicient, et cum bestiis feris erit habitatio tua: fenum quasi boves comedes; et septem tempora mutabuntur super te, donec scias quod dominetur Excelsus in regno hominum et, cuicumque voluerit, det illud ".
DAN|4|30|Eadem hora sermo completus est super Nabuchodonosor, et ex hominibus abiectus est et fenum ut boves comedit, et rore caeli corpus eius infectum est, donec capilli eius in similitudinem aquilarum crescerent, et ungues eius quasi avium.
DAN|4|31|" Igitur post finem dierum ego Nabuchodonosor oculos meos ad caelum levavi, et sensus meus redditus est mihi, et Altissimo benedixi et Viventem in sempiternum laudavi et glorificavi,quia potestas eius potestas sempiterna,et regnum eius in generationem et generationem;
DAN|4|32|et omnes habitatores terrae apud eum in nihilum reputati sunt:iuxta voluntatem enim suam facittam in virtutibus caeli quam in habitatoribus terrae,et non est qui resistat manui eiuset dicat ei: "Quid facis?".
DAN|4|33|In ipso tempore sensus meus reversus est ad me, et ad honorem regni mei maiestas mea et splendor meus reversa sunt ad me; et optimates mei et magistratus mei requisierunt me, et in regno meo constitutus sum, et magnificentia amplior addita est mihi.
DAN|4|34|Nunc igitur ego Nabuchodonosor laudo et magnifico et glorifico Regem caeli, quia omnia opera eius veritas, et viae eius iudicium, et gradientes in superbia potest humiliare ".
DAN|5|1|Balthasar rex fecit grande con vivium optimatibus suis mille et coram his milibus vinum bibebat.
DAN|5|2|Balthasar ergo praecepit iam temulentus, ut afferrentur vasa aurea et argentea, quae asportaverat Nabuchodonosor pater eius de templo, quod fuit in Ierusalem, ut biberent in eis rex et optimates eius uxoresque eius et concubinae.
DAN|5|3|Tunc allata sunt vasa aurea, quae asportaverat de templo, quod fuerat in Ierusalem; et biberunt in eis rex et optimates eius, uxores et concubinae illius:
DAN|5|4|bibebant vinum et laudabant deos suos aureos et argenteos, aereos, ferreos ligneosque et lapideos.
DAN|5|5|In eadem hora apparuerunt digiti manus hominis et scripserunt contra candelabrum in superficie parietis palatii regis; et rex aspiciebat articulos manus scribentis.
DAN|5|6|Tunc regis facies commutata est, et cogitationes eius conturbabant eum, et compages renum eius solvebantur, et genua eius ad se invicem collidebantur.
DAN|5|7|Exclamavit itaque rex fortiter, ut introducerent magos, Chaldaeos et haruspices; et proloquens rex ait sapientibus Babylonis: " Quicumque legerit scripturam hanc et interpretationem eius manifestam mihi fecerit, purpura vestietur et torquem auream habebit in collo et tertius in regno meo dominabitur ".
DAN|5|8|Tunc ingressi sunt omnes sapientes regis et non potuerunt nec scripturam legere nec interpretationem indicare regi;
DAN|5|9|unde rex Balthasar satis conturbatus est, et vultus illius immutatus est super eum, sed et optimates eius turbabantur.
DAN|5|10|Regina autem, sermonum regis optimatiumque eius causa, domum convivii ingressa est; et regina proloquens ait: " Rex, in aeternum vive! Non te conturbent cogitationes tuae, neque facies tua immutetur.
DAN|5|11|Est vir in regno tuo, qui spiritum deorum sanctorum habet in se, et in diebus patris tui scientia et intellegentia et sapientia quasi sapientia deorum inventae sunt in eo; nam et rex Nabuchodonosor pater tuus principem magorum, incantatorum, Chaldaeorum et haruspicum constituit eum; pater tuus, o rex,
DAN|5|12|quia spiritus amplior et prudentia intellegentiaque et interpretatio somniorum et ostensio secretorum ac solutio ligatorum inventae sunt in eo, in Daniele, cui rex posuit nomen Baltassar. Nunc itaque Daniel vocetur et interpretationem narrabit ".
DAN|5|13|Igitur introductus est Daniel coram rege; ad quem praefatus rex ait: " Tu es Daniel de filiis captivitatis Iudae, quem adduxit rex pater meus de Iuda?
DAN|5|14|Audivi de te quoniam spiritum deorum habeas, et scientia intellegentiaque ac sapientia ampliores inventae sint in te.
DAN|5|15|Et nunc introgressi sunt in conspectu meo sapientes, magi, ut scripturam hanc legerent et interpretationem eius indicarent mihi et nequiverunt sensum huius sermonis edicere.
DAN|5|16|Porro ego audivi de te quod possis obscura interpretari et ligata dissolvere; si ergo vales scripturam legere et interpretationem eius indicare mihi, purpura vestieris et torquem auream circa collum tuum habebis et tertius in regno meo princeps eris ".
DAN|5|17|Tunc respondens Daniel ait coram rege: " Munera tua sint tibi, et dona tua alteri da; scripturam autem legam tibi, rex, et interpretationem eius ostendam tibi.
DAN|5|18|O rex, Deus altissimus regnum et magnificentiam et gloriam et honorem dedit Nabuchodonosor patri tuo.
DAN|5|19|Et propter magnificentiam, quam dederat ei, universi populi, tribus et linguae tremebant et metuebant eum; quos volebat, interficiebat et, quos volebat, percutiebat et, quos volebat, exaltabat et, quos volebat, humiliabat.
DAN|5|20|Quando autem elevatum est cor eius, et spiritus illius obfirmatus est ad superbiam, depositus est de solio regni sui, et gloria eius ablata est ab eo;
DAN|5|21|et a filiis hominum eiectus est, sed et cor eius cum bestiis positum est, et cum onagris erat habitatio eius, fenum quoque ut boves comedebat, et rore caeli corpus eius infectum est, donec cognosceret quod potestatem haberet Deus altissimus in regno hominum et, quemcumque voluerit, suscitabit super illud.
DAN|5|22|Tu quoque filius eius, Balthasar, non humiliasti cor tuum, cum scires haec omnia,
DAN|5|23|sed adversum Dominum caeli elevatus es, et vasa domus eius allata sunt coram te, et tu et optimates tui et uxores tuae et concubinae tuae vinum bibistis in eis; deos quoque argenteos et aureos et aereos, ferreos ligneosque et lapideos, qui non vident neque audiunt neque sentiunt, laudasti, porro Deum, qui habet flatum tuum in manu sua et omnes vias tuas, non glorificasti.
DAN|5|24|Idcirco ab eo missi sunt articuli manus, et scriptura haec exarata est.
DAN|5|25|Haec est autem scriptura, quae digesta est: mane, thecel, upharsin.
DAN|5|26|Et haec est interpretatio sermonis: mane, numeravit Deus regnum tuum et complevit illud;
DAN|5|27|thecel, appensus es in statera et inventus es minus habens;
DAN|5|28|phares, divisum est regnum tuum et datum est Medis et Persis ".
DAN|5|29|Tunc, iubente Balthasar, indutus est Daniel purpura, et circumdata est torques aurea collo eius, et praedicatum est de eo quod haberet potestatem tertius in regno suo.
DAN|5|30|Eadem nocte interfectus est Balthasar rex Chaldaeorum.
DAN|6|1|Et Darius Medus successit in regnum annos natus sexaginta duos.
DAN|6|2|Placuit Dario et constituit super regnum satrapas centum viginti, ut essent in toto regno suo,
DAN|6|3|et super eos principes tres, ex quibus Daniel unus erat, ut satrapae illis redderent rationem, et rex non sustineret molestiam.
DAN|6|4|Igitur ille Daniel superabat omnes principes et satrapas, quia spiritus Dei amplior erat in eo. Porro rex cogitabat constituere eum super omne regnum;
DAN|6|5|unde principes et satrapae quaerebant, ut invenirent occasionem Danieli ex latere regni, nullamque causam et suspicionem reperire potuerunt, eo quod fidelis esset, et omnis culpa et suspicio non inveniretur in eo.
DAN|6|6|Dixerunt ergo viri illi: " Non inveniemus Danieli huic aliquam occasionem, nisi forte inveniamus adversus eum in lege Dei sui ".
DAN|6|7|Tunc principes et satrapae illi concurrerunt ad regem et sic locuti sunt ei: " Darie rex, in aeternum vive!
DAN|6|8|Consilium inierunt cuncti principes regni, magistratus et satrapae, optimates et iudices, ut decretum regis promulget et edictum confirmet, ut omnis, qui petierit aliquam petitionem a quocumque deo et homine usque ad dies triginta, nisi a te, rex, mittatur in lacum leonum.
DAN|6|9|Nunc itaque, rex, confirma sententiam et signa decretum, ut non immutetur iuxta legem Medorum et Persarum, quam praevaricari non licet ".
DAN|6|10|Porro rex Darius signavit edictum et decretum.
DAN|6|11|Daniel autem, cum comperisset decretum signatum esse, ingressus est domum suam et, fenestris apertis in cenaculo suo contra Ierusalem, tribus temporibus in die flectebat genua sua et adorabat confitebaturque coram Deo suo, sicut et ante facere consueverat.
DAN|6|12|Viri ergo illi accesserunt et invenerunt Danielem orantem et obsecrantem Deum suum.
DAN|6|13|Tunc accesserunt et locuti sunt coram rege super edicto: " Rex, numquid non signasti decretum, ut omnis homo, qui rogaret quemquam de diis et hominibus usque ad dies triginta, nisi a te, rex, mitteretur in lacum leonum? ". Respondens rex ait: " Verus est sermo iuxta decretum Medorum atque Persarum, quod praevaricari non licet ".
DAN|6|14|Tunc respondentes dixerunt coram rege: " Daniel de filiis captivitatis Iudae non curavit de te, rex, et de edicto, quod constituisti, sed tribus temporibus per diem orat obsecratione sua".
DAN|6|15|Quod verbum cum audisset, rex satis contristatus est; et pro Daniele posuit cor, ut liberaret eum, et usque ad occasum solis laborabat, ut erueret illum.
DAN|6|16|Viri autem illi accesserunt ad regem et dixerunt ei: " Scito, rex, quia lex Medorum est atque Persarum, ut omne decretum et edictum, quod constituit rex, non liceat immutari ".
DAN|6|17|Tunc rex praecepit, et adduxerunt Danielem et miserunt eum in lacum leonum. Dixitque rex Danieli: " Deus tuus, quem colis semper, ipse liberet te ".
DAN|6|18|Allatusque est lapis unus et positus est super os laci; quem obsignavit rex anulo suo et anulo optimatum suorum, ne quid fieret contra Danielem.
DAN|6|19|Et abiit rex in domum suam et dormivit incenatus, cibique non sunt illati coram eo; insuper et somnus recessit ab eo.
DAN|6|20|Tunc rex primo diluculo consurgens festinus ad lacum leonum perrexit;
DAN|6|21|appropinquansque lacui Danielem voce lacrimabili inclamavit et affatus est Danielem: " Daniel, serve Dei viventis, Deus tuus, cui tu servis semper, putasne valuit liberare te a leonibus?".
DAN|6|22|Et Daniel regi respondens ait: " Rex, in aeternum vive!
DAN|6|23|Deus meus misit angelum suum et conclusit ora leonum, et non nocuerunt mihi, quia coram eo iustitia inventa est in me; sed et coram te, rex, delictum non feci ".
DAN|6|24|Tunc rex vehementer gavisus est super eo et Danielem praecepit educi de lacu; eductusque est Daniel de lacu, et nulla laesio inventa est in eo, quia credidit Deo suo.
DAN|6|25|Dixit autem rex, et adducti sunt viri illi, qui accusaverant Danielem, et in lacum leonum missi sunt, ipsi et filii eorum et uxores eorum, et non pervenerunt usque ad pavimentum laci, donec potirentur eis leones, et omnia ossa eorum comminuerunt.
DAN|6|26|Tunc Darius rex scripsit universis populis, tribubus et linguis, habitantibus in universa terra: "Pax vobis multiplicetur!
DAN|6|27|A me constitutum est decretum, ut in universo imperio regni mei tremescant et paveant Deum Danielis:ipse est enim Deus vivenset permanens in saecula,et regnum eius non dissipabitur,et potestas eius usque in aeternum;
DAN|6|28|ipse liberator atque salvatoret faciens signa et mirabiliain caelo et in terra.Liberavit autem Danielemde manu leonum ".
DAN|6|29|Porro Daniel prosperatus est in regno Darii et in regno Cyri Persae.
DAN|7|1|Anno primo Balthasar regis Babylonis Daniel somnium vidit et visionem capitis eius in cubili suo; tunc et somnium scripsit. Caput verborum, quae locutus est.
DAN|7|2|Respondit Daniel et dixit: " Videbam in visione mea nocte: et ecce quattuor venti caeli conturbabant mare Magnum,
DAN|7|3|et quattuor bestiae grandes ascendebant de mari diversae inter se.
DAN|7|4|Prima quasi leaena et alas habebat aquilae; aspiciebam, donec evulsae sunt alae eius; et sublata est de terra et super pedes quasi homo stetit, et cor hominis datum est ei.
DAN|7|5|Et ecce bestia alia, secunda, similis urso in parte stetit, et tres costae erant in ore eius et in dentibus eius; et sic dicebant ei: "Surge, comede carnes plurimas".
DAN|7|6|Post hoc aspiciebam, et ecce alia quasi pardus et alas habebat avis quattuor super se, et quattuor capita erant in bestia; et potestas data est ei.
DAN|7|7|Post hoc aspiciebam in visione noctis, et ecce bestia quarta terribilis atque mirabilis et fortis nimis; dentes ferreos habebat magnos, comedens atque comminuens et reliqua pedibus suis conculcans; dissimilis autem erat ceteris bestiis, quas videram ante eam, et habebat cornua decem.
DAN|7|8|Considerabam cornua, et ecce cornu aliud parvulum ortum est de medio eorum, et tria de cornibus primis evulsa sunt a facie eius; et ecce oculi quasi oculi hominis erant in cornu isto, et os loquens ingentia.
DAN|7|9|Aspiciebam,donec throni positi sunt,et Antiquus dierum sedit.Vestimentum eius quasi nix candidum,et capilli capitis eius quasi lana munda;thronus eius flammae ignis,rotae eius ignis accensus.
DAN|7|10|Fluvius igneus effluebatet egrediebatur a facie eius;milia milium ministrabant ei,et decies milies centena milia assistebant ei:iudicium sedit,et libri aperti sunt.
DAN|7|11|Aspiciebam tunc propter vocem sermonum grandium, quos cornu illud loquebatur; et vidi quoniam interfecta esset bestia, et perisset corpus eius, et tradita esset ad comburendum igni;
DAN|7|12|aliarum quoque bestiarum ablata esset potestas, et tempora vitae constituta essent eis usque ad tempus et tempus.
DAN|7|13|Aspiciebam ergo in visione noctis:et ecce cum nubibus caeliquasi Filius hominis veniebatet usque ad Antiquum dierum pervenit,et in conspectu eius obtulerunt eum;
DAN|7|14|et data sunt ei potestas et honor et regnum;et omnes populi, tribus et linguaeipsi servierunt:potestas eius potestas aeterna,quae non auferetur,et regnum eius, quod non corrumpetur.
DAN|7|15|Horruit spiritus meus: ego Daniel territus sum in his, et visiones capitis mei conturbaverunt me.
DAN|7|16|Accessi ad unum de assistentibus et veritatem quaerebam ab eo de omnibus his; qui dixit mihi et interpretationem sermonum edocuit me:
DAN|7|17|"Hae bestiae magnae quattuor, quattuor regna consurgent de terra;
DAN|7|18|suscipient autem regnum sancti Dei altissimi et obtinebunt regnum usque in saeculum et saeculum saeculorum".
DAN|7|19|Post hoc volui diligenter discere de bestia quarta, quae erat dissimilis valde ab omnibus his et terribilis nimis, dentes ferrei et ungues eius aerei, comedens et comminuens et reliquias pedibus suis conculcans,
DAN|7|20|et de cornibus decem, quae habebat in capite, et de alio, quod ortum fuerat ante, et ceciderant tria cornua, de cornu illo, quod habebat oculos et os loquens grandia et maius erat ceteris.
DAN|7|21|Aspiciebam, et ecce cornu illud faciebat bellum adversus sanctos et praevalebat eis,
DAN|7|22|donec venit Antiquus dierum et iudicium dedit sanctis Excelsi, et tempus advenit, et regnum obtinuerunt sancti.
DAN|7|23|Et sic ait: "Bestia quarta regnum quartum erit in terra, quod maius erit omnibus regnis et devorabit universam terram et conculcabit et comminuet eam.
DAN|7|24|Porro cornua decem regni decem reges erunt; et alius consurget post eos et ipse potentior erit prioribus et tres reges humiliabit
DAN|7|25|et sermones contra Excelsum loquetur et sanctos Altissimi conteret et putabit quod possit mutare tempora et legem, et tradentur in manu eius usque ad tempus et tempora et dimidium temporis;
DAN|7|26|et iudicium sedebit, et potentiam eius auferent, ut conteratur et dispereat usque in finem;
DAN|7|27|regnum autem et potestas et magnitudo regnorum, quae sunt subter omne caelum, detur populo sanctorum Altissimi, cuius regnum regnum sempiternum est, et omnes reges servient ei et oboedient" ".
DAN|7|28|Hucusque finis verbi. Ego Daniel multum cogitationibus meis conturbabar, et facies mea mutata est in me; verbum autem in corde meo conservavi.
DAN|8|1|Anno tertio regni Balthasar regis visio apparuit mihi, ego Daniel, post id quod mihi apparuerat in principio.
DAN|8|2|Vidi in visione, et factum est, dum viderem, eram in Susis castro, quod est in Elam provincia; vidi autem in visione esse me super rivum Ulai.
DAN|8|3|Et levavi oculos meos et vidi: et ecce aries unus stabat ante rivum habens cornua et cornua excelsa et unum excelsius altero, et excelsius crescebat in postero.
DAN|8|4|Vidi arietem cornibus ventilantem contra occidentem et contra aquilonem et contra meridiem, et omnes bestiae non poterant resistere ei neque liberari de manu eius; fecitque secundum voluntatem suam et magnificatus est.
DAN|8|5|Et ego intellegebam: ecce autem hircus caprarum veniebat ab occidente super faciem totius terrae et non tangebat terram; porro hircus habebat cornu insigne inter oculos suos.
DAN|8|6|Et venit usque ad arietem illum cornutum, quem videram stantem ante rivum, et cucurrit ad eum in impetu fortitudinis suae.
DAN|8|7|Vidi eum appropinquantem prope arietem, et efferatus est in eum et percussit arietem et comminuit duo cornua eius, et non poterat aries resistere ei; cumque eum misisset in terram, conculcavit, et nemo quibat liberare arietem de manu eius.
DAN|8|8|Hircus autem caprarum magnus factus est nimis; cumque crevisset, fractum est cornu magnum, et orta sunt quattuor cornua loco illius per quattuor ventos caeli.
DAN|8|9|De uno autem ex eis egressum est cornu unum modicum et factum est grande contra meridiem et contra orientem et contra fortitudinem
DAN|8|10|et magnificatum est usque ad fortitudinem caeli et deiecit de fortitudine et de stellis et conculcavit eas;
DAN|8|11|et usque ad principem fortitudinis magnificatum est et ab eo tulit iuge sacrificium et deiecit locum sanctificationis eius.
DAN|8|12|Militia autem data est contra iuge sacrificium propter peccata, et prostrata est veritas in terra; cornu autem fecit et prosperatum est.
DAN|8|13|Et audivi unum de sanctis loquentem, et dixit unus sanctus alteri, nescio cui, loquenti: " Usquequo visio et iuge sacrificium et peccatum desolationis, quae facta est, et sanctuarium et fortitudo conculcabitur?.
DAN|8|14|Et dixit ei: " Usque ad vesperam et mane, dies duo milia trecenti; et mundabitur sanctuarium ".
DAN|8|15|Factum est autem cum viderem ego Daniel visionem et quaererem intellegentiam, ecce stetit in conspectu meo quasi species viri;
DAN|8|16|et audivi vocem viri inter Ulai, et clamavit et ait: " Gabriel, fac intellegere istum visionem ".
DAN|8|17|Et venit et stetit iuxta, ubi ego stabam; cumque venisset, pavens corrui in faciem meam, et ait ad me: "Intellege, fili hominis, quoniam in tempore finis complebitur visio ".
DAN|8|18|Cumque loqueretur ad me, collapsus sum pronus in terram, et tetigit me et statuit me in gradu meo
DAN|8|19|dixitque: " Ecce ego ostendam tibi, quae futura sint in novissimo maledictionis, quoniam in tempore erit finis.
DAN|8|20|Aries, quem vidisti habere cornua, reges Medorum est atque Persarum;
DAN|8|21|porro hircus caprarum rex Graecorum est, et cornu grande, quod erat inter oculos eius, ipse est rex primus.
DAN|8|22|Quod autem, fracto illo, surrexerunt quattuor pro eo, quattuor regna de gente eius consurgent sed non in fortitudine eius.
DAN|8|23|Et post regnum eorum, cum creverint iniquitate, consurget rex impudens facie et intellegens propositiones;
DAN|8|24|et roborabitur fortitudo eius sed non in viribus suis, et supra quam credi potest universa vastabit et prosperabitur et faciet et interficiet robustos et populum sanctorum,
DAN|8|25|et secundum sapientiam suam prosperabitur dolus in manu eius, et in corde suo magnificabitur et in tranquillitate occidet plurimos et contra principem principum consurget et sine manu conteretur.
DAN|8|26|Et visio vespere et mane, quae dicta est, vera est; tu ergo signa visionem, quia post dies multos erit ".
DAN|8|27|Et ego Daniel langui et aegrotavi per dies; cumque surrexissem, faciebam opera regis et stupebam ad visionem, et non erat qui intellegeret.
DAN|9|1|In anno primo Darii filii Asueri de semine Medorum, qui impe ravit super regnum Chaldaeorum,
DAN|9|2|anno uno regni eius, ego Daniel intellexi in libris numerum annorum, de quo factus est sermo Domini ad Ieremiam prophetam, ut complerentur desolationes Ierusalem, septuaginta anni;
DAN|9|3|et posui faciem meam ad Dominum Deum meum, ut quaererem rogationem et deprecationem in ieiuniis, sacco et cinere.
DAN|9|4|Et oravi Dominum Deum et confessus sum et dixi: Obsecro, Domine, Deus magne et terribilis, custodiens pactum et misericordiam diligentibus eum et custodientibus mandata eius;
DAN|9|5|peccavimus, inique fecimus, impie egimus et recessimus et declinavimus a mandatis tuis ac iudiciis tuis;
DAN|9|6|non oboedivimus servis tuis prophetis, qui locuti sunt in nomine tuo regibus nostris, principibus nostris, patribus nostris omnique populo terrae.
DAN|9|7|Tibi, Domine, iustitia; nobis autem confusio faciei, sicut est hodie viro Iudae et habitatoribus Ierusalem et omni Israel, his qui prope sunt et his qui procul in universis terris, ad quas eiecisti eos propter iniquitates eorum, in quibus peccaverunt in te.
DAN|9|8|Domine, nobis confusio faciei, regibus nostris, principibus nostris et patribus nostris, quia peccavimus tibi;
DAN|9|9|Domino autem, Deo nostro, misericordia et propitiatio, quia recessimus a te.
DAN|9|10|Et non audivimus vocem Domini Dei nostri, ut ambularemus in lege eius, quam posuit nobis per servos suos prophetas;
DAN|9|11|et omnis Israel praevaricati sunt legem tuam et declinaverunt, ne audirent vocem tuam, et stillavit super nos maledictio et detestatio, quae scripta est in libro Moysis servi Dei, quia peccavimus ei.
DAN|9|12|Et statuit sermones suos, quos locutus est super nos et super iudices nostros, qui iudicaverunt nos, ut superducerent in nos magnum malum, quale numquam fuit sub omni caelo, secundum quod factum est in Ierusalem.
DAN|9|13|Sicut scriptum est in lege Moysis, omne malum hoc venit super nos, et non rogavimus faciem Domini Dei nostri, ut reverteremur ab iniquitatibus nostris et cogitaremus veritatem tuam.
DAN|9|14|Et vigilavit Dominus super malitiam et adduxit eam super nos, quia iustus Dominus Deus noster in omnibus operibus suis, quae fecit; non enim audivimus vocem eius.
DAN|9|15|Et nunc, Domine Deus noster, qui eduxisti populum tuum de terra Aegypti in manu forti et fecisti tibi nomen secundum diem hanc, peccavimus, iniquitatem fecimus,
DAN|9|16|Domine, in omnem iustitiam tuam; avertatur, obsecro, ira tua et furor tuus a civitate tua Ierusalem et monte sancto tuo; propter peccata enim nostra et iniquitates patrum nostrorum Ierusalem et populus tuus in opprobrium sunt omnibus per circuitum nostrum.
DAN|9|17|Nunc ergo exaudi, Deus noster, orationem servi tui et preces eius et ostende faciem tuam super sanctuarium tuum, quod desertum est, propter temetipsum.
DAN|9|18|Inclina, Deus meus, aurem tuam et audi; aperi oculos tuos et vide desolationem nostram et civitatem, super quam invocatum est nomen tuum; neque enim in iustificationibus nostris prosternimus preces ante faciem tuam sed in miserationibus tuis multis.
DAN|9|19|Exaudi, Domine! Placare, Domine! Attende et fac! Ne moreris propter temetipsum, Deus meus, quia nomen tuum invocatum est super civitatem et super populum tuum ".
DAN|9|20|Cumque adhuc loquerer et orarem et confiterer peccata mea et peccata populi mei Israel et prosternerem preces meas in conspectu Dei mei pro monte sancto Dei mei,
DAN|9|21|adhuc me loquente in oratione, ecce vir Gabriel, quem videram in visione principio, cito volans tetigit me in tempore sacrificii vespertini;
DAN|9|22|et docuit me et locutus est mihi dixitque: "Daniel, nunc egressus sum, ut docerem te, et intellegeres.
DAN|9|23|Ab exordio precum tuarum egressus est sermo; ego autem veni, ut indicarem, quia vir desideriorum es tu; ergo animadverte sermonem et intellege visionem.
DAN|9|24|Septuaginta hebdomades decretae suntsuper populum tuum et super urbem sanctam tuam,ut consummetur praevaricatio,et finem accipiat peccatum,et deleatur iniquitas,et adducatur iustitia sempiterna,et impleatur visio et prophetes,et ungatur Sanctus sanctorum.
DAN|9|25|Scito ergo et animadverte:ab exitu sermonisut iterum aedificetur Ierusalemusque ad christum ducem,hebdomades septem.Et hebdomades sexaginta duae erunt;et rursum aedificabitur platea et muriin angustia temporum.
DAN|9|26|Et post hebdomades sexaginta duasoccidetur christus;et nihil erit ei.Et civitatem et sanctuarium dissipabitpopulus ducis venturi,et finis eius vastitas,et usque ad finem bellistatuta desolatio.
DAN|9|27|Confirmabit autem pactum multishebdomade una;et in dimidio hebdomadideficiet hostia et sacrificium,et erit super alam abominationis vastator,et usquedum consummatio et decretumeffundantur super vastatorem ".
DAN|10|1|Anno tertio Cyri regis Per sarum verbum revelatum est Danieli cognomento Baltassar, et verum verbum et acies magna; intellexitque sermonem, intellegentia enim fuit ei in visione.
DAN|10|2|In diebus illis ego Daniel lugebam tribus hebdomadis dierum,
DAN|10|3|panem desiderabilem non comedi, et caro et vinum non introierunt in os meum, sed neque unguento unctus sum, donec complerentur tres hebdomades dierum.
DAN|10|4|Die autem vicesima et quarta mensis primi eram iuxta fluvium magnum, qui est Tigris,
DAN|10|5|et levavi oculos meos et vidi: et ecce vir unus vestitus lineis, et renes eius accincti auro obryzo;
DAN|10|6|et corpus eius quasi chrysolithus, et facies eius velut species fulgoris, et oculi eius ut lampas ardens, et brachia eius et, quae deorsum sunt usque ad pedes, quasi species aeris candentis, et vox sermonum eius ut vox multitudinis.
DAN|10|7|Vidi autem ego Daniel solus visionem; porro viri, qui erant mecum, visionem non viderunt, sed terror nimius irruit super eos, et fugerunt in absconditum.
DAN|10|8|Ego autem relictus solus vidi visionem grandem hanc, et non remansit in me fortitudo, sed et species mea immutata est in me usque ad dissipationem, nec habui quidquam virium.
DAN|10|9|Et audivi vocem sermonum eius; et audiens vocem sermonum eius iacebam consternatus super faciem meam, et vultus meus haerebat terrae.
DAN|10|10|Et ecce manus tetigit me et erexit me super genua mea et super palmas manuum mearum,
DAN|10|11|et dixit ad me: " Daniel, vir desideriorum, intellege verba, quae ego loquor ad te, et sta in gradu tuo; nunc enim sum missus ad te ". Cumque dixisset mihi sermonem istum, steti tremens.
DAN|10|12|Et ait ad me: " Noli metuere, Daniel, quia ex die primo, quo posuisti cor tuum ad intellegendum et ad humiliandum te in conspectu Dei tui, exaudita sunt verba tua; et ego veni propter sermones tuos.
DAN|10|13|Princeps autem regni Persarum restitit mihi viginti et uno diebus; et ecce Michael, unus de principibus primis, venit in adiutorium meum; et ego remansi ibi iuxta regem Persarum.
DAN|10|14|Veni autem, ut docerem te, quae ventura sunt populo tuo in novissimis diebus, quoniam adhuc visio in dies ".
DAN|10|15|Cumque loqueretur mihi huiuscemodi verbis, deieci vultum meum ad terram et tacui.
DAN|10|16|Et ecce quasi similitudo filiorum hominis tetigit labia mea; et aperiens os meum locutus sum et dixi ad eum, qui stabat contra me: " Domine mi, in visione angustiae venerunt super me, et nihil in me remansit virium.
DAN|10|17|Et quomodo poterit servus domini mei loqui cum hoc domino meo? Nihil enim in me remansit virium, et halitus meus non remansit in me ".
DAN|10|18|Rursum ergo tetigit me quasi visio hominis et confortavit me
DAN|10|19|et dixit: "Noli timere, vir desideriorum; pax tibi, confortare et esto robustus ". Cumque loqueretur mecum, convalui et dixi: " Loquere, domine mi, quia confortasti me ".
DAN|10|20|Et ait: " Numquid scis, quare venerim ad te? Et nunc revertar, ut proelier adversum principem Persarum. Et ego egrediar, et ecce princeps Graecorum veniens.
DAN|10|21|Verumtamen annuntiabo tibi, quod expressum est in scriptura veritatis; et nemo est adiutor meus adversus hos, nisi Michael princeps vester.
DAN|11|1|Ego autem ab anno primo Darii Medi astabam ei, ut confortaretur et roboraretur.
DAN|11|2|Et nunc veritatem annuntiabo tibi: Ecce adhuc tres reges stabunt pro Perside, et quartus ditabitur opibus nimis super omnes et, cum invaluerit divitiis suis, concitabit omnia adversum regnum Graeciae.
DAN|11|3|Surget vero rex fortis et dominabitur dominatione multa et faciet, quod placuerit ei;
DAN|11|4|et cum steterit, conteretur regnum eius et dividetur in quattuor ventos caeli, sed non in posteros eius neque secundum potentiam illius, qua dominatus est; lacerabitur enim regnum eius etiam ad alios, exceptis his.
DAN|11|5|Et confortabitur rex austri, et unus de principibus eius praevalebit super eum et dominabitur dominatione super dominationem eius.
DAN|11|6|Et post finem annorum foederabuntur; filiaque regis austri veniet ad regem aquilonis facere amicitiam. Et non obtinebit fortitudinem brachii, nec stabit brachium eius; et tradetur ipsa, et qui adduxerunt eam, et adulescens eius, et qui confortabat eam in temporibus.
DAN|11|7|Et stabit de germine radicum eius plantatio loco eius et veniet ad exercitum et ingredietur oppidum regis aquilonis; et faciet adversus eos et confortabitur.
DAN|11|8|Insuper et deos eorum cum sculptilibus eorum et vasis pretiosis argenti et auri captivos ducet in Aegyptum: ipse per aliquot annos praevalebit adversus regem aquilonis.
DAN|11|9|Et intrabit in regnum regis austri et revertetur ad terram suam.
DAN|11|10|Filii autem eius provocabuntur et congregabunt multitudinem exercituum plurimorum; et veniet properans et inundans et revertetur et concitabitur et congredietur usque ad oppidum eius.
DAN|11|11|Et provocabitur rex austri et egredietur et pugnabit adversus eum, adversus regem aquilonis; et praeparabit multitudinem nimiam, et dabitur multitudo in manu eius.
DAN|11|12|Et tolletur multitudo, et exaltabitur cor eius, et deiciet multa milia, sed non praevalebit.
DAN|11|13|Revertetur enim rex aquilonis et praeparabit multitudinem maiorem quam prius; et in fine temporum annorumque veniet properans cum exercitu magno et opibus nimis.
DAN|11|14|Et in temporibus illis multi consurgent adversus regem austri, filii quoque praevaricatorum populi tui extollentur, ut impleant visionem, et corruent.
DAN|11|15|Et veniet rex aquilonis et comportabit aggerem et capiet urbem munitissimam; et brachia austri non sustinebunt, et populo electorum eius non erit fortitudo ad resistendum.
DAN|11|16|Et faciet veniens super eum iuxta placitum suum, et non erit qui stet contra faciem eius; et stabit in terra inclita, et consumptio in manu eius.
DAN|11|17|Et ponet faciem suam, ut veniat ad tenendum universum regnum eius, et recta faciet cum eo et filiam feminarum dabit ei, ut evertat illud; et non stabit nec illius erit.
DAN|11|18|Et convertet faciem suam ad insulas et capiet multas, et cessare faciet princeps opprobrium eius, et opprobrium eius convertetur in eum.
DAN|11|19|Et convertet faciem suam ad oppida terrae suae et impinget et corruet, et non invenietur.
DAN|11|20|Et stabit in loco eius, qui mittat exactorem in decus regni; et in paucis diebus conteretur, non in furore nec in proelio.
DAN|11|21|Et stabit in loco eius despectus, et non tribuetur ei honor regius; et veniet clam et obtinebit regnum in fraudulentia.
DAN|11|22|Et brachia pugnantis expugnabuntur a facie eius et conterentur; insuper et dux foederis.
DAN|11|23|Et post amicitias, cum eo faciet dolum et ascendet et superabit in modico populo.
DAN|11|24|In prosperitate uberes urbes ingredietur et faciet, quae non fecerunt patres eius et patres patrum eius: rapinas et praedam et divitias eorum dissipabit et contra oppida cogitationes inibit, et hoc usque ad tempus.
DAN|11|25|Et concitabitur fortitudo eius et cor eius adversum regem austri in exercitu magno; et rex austri provocabitur ad bellum multis auxiliis et fortibus nimis, et non stabit, quia inibunt adversus eum consilia.
DAN|11|26|Et comedentes panem cum eo conterent illum; exercitusque eius opprimetur, et cadent interfecti plurimi.
DAN|11|27|Duorum quoque regum cor erit, ut malefaciant et ad mensam unam mendacium loquentur et non proficient, quia adhuc finis in aliud tempus.
DAN|11|28|Et revertetur in terram suam cum opibus multis, et cor eius adversum testamentum sanctum; et faciet et revertetur in terram suam.
DAN|11|29|Statuto tempore revertetur et veniet ad austrum, et non erit priori simile novissimum.
DAN|11|30|Et venient super eum trieres, Romani; et percutietur et revertetur et indignabitur contra testamentum sanctum et faciet reverteturque et cogitabit adversum eos, qui dereliquerunt testamentum sanctum.
DAN|11|31|Et brachia ex eo stabunt et polluent sanctuarium fortitudinis et auferent iuge sacrificium et dabunt abominationem vastatoris.
DAN|11|32|Et impios in testamentum errare faciet fraudulenter; populus autem scientium Deum suum obtinebit et faciet.
DAN|11|33|Et docti in populo docebunt plurimos; et ruent in gladio et in flamma et in captivitate et in rapina per dies.
DAN|11|34|Cumque corruerint, sublevabuntur auxilio parvulo, et applicabuntur eis plurimi fraudulenter.
DAN|11|35|Et de eruditis ruent, ut aliqui eorum conflentur et purgentur et dealbentur usque ad tempus praefinitum, quia adhuc aliud tempus erit.
DAN|11|36|Et faciet iuxta voluntatem suam rex et elevabitur et magnificabitur adversus omnem deum et adversus Deum deorum loquetur magnifica et prosperabitur, donec compleatur iracundia; perpetrata quippe est definitio.
DAN|11|37|Et deos patrum suorum non reputabit neque concupiscentiam feminarum nec quemquam deorum curabit, quia super universa magnificabit se;
DAN|11|38|deum autem oppidorum in loco suo venerabitur et deum, quem ignoraverunt patres eius, colet auro et argento et lapide pretioso rebusque pretiosis
DAN|11|39|et faciet adversus oppida munita cum deo alieno; qui cognoverit eum, multiplicabit gloriam eius et dabit eis potestatem in multis et terram dividet pretio.
DAN|11|40|Et in tempore praefinito proeliabitur adversus eum rex austri, et quasi tempestas veniet contra illum rex aquilonis in curribus et in equitibus et in classe magna, et ingredietur terras et conteret et pertransiet.
DAN|11|41|Et introibit in terram gloriosam, et multae corruent; hae autem solae salvabuntur de manu eius: Edom et Moab et principium filiorum Ammon.
DAN|11|42|Et mittet manum suam in terras, et terra Aegypti non effugiet;
DAN|11|43|et dominabitur thesaurorum auri et argenti et in omnibus pretiosis Aegypti, et Libyes et Aethiopes in vestigia eius transibunt.
DAN|11|44|Et fama turbabit eum ab oriente et ab aquilone; et veniet in ira magna, ut conterat et interficiat plurimos,
DAN|11|45|et figet tabernacula palatii sui inter maria super montem sanctum decoris; et veniet usque ad summitatem eius, et nemo auxiliabitur ei.
DAN|12|1|In tempore autem illo con surget Michael, princeps magnus, qui stat pro filiis populi tui, et erit tempus angustiae, quale non fuit ab eo, quo gentes esse coeperunt, usque ad tempus illud. Et in tempore illo salvabitur populus tuus, omnis, qui inventus fuerit scriptus in libro.
DAN|12|2|Et multi de his, qui dormiunt in terra pulveris, evigilabunt: alii in vitam aeternam, et alii in opprobrium sempiternum.
DAN|12|3|Qui autem docti fuerint, fulgebunt quasi splendor firmamenti; et, qui ad iustitiam erudierint multos, quasi stellae in perpetuas aeternitates.
DAN|12|4|Tu autem, Daniel, claude sermones et signa librum usque ad tempus finis; pertransibunt plurimi, et multiplex erit scientia ".
DAN|12|5|Et vidi ego Daniel: et ecce duo alii stabant, unus hinc super ripam fluminis, et alius inde ex altera ripa fluminis.
DAN|12|6|Et dixit viro, qui indutus erat lineis, qui stabat super aquas fluminis: Usquequo finis horum mirabilium? ".
DAN|12|7|Et audivi virum, qui indutus erat lineis, qui stabat super aquas fluminis, cum levasset dexteram et sinistram suam in caelum et iurasset per Viventem in aeternum: " Quia in tempus, tempora et dimidium temporis; et cum completa fuerit dispersio manus populi sancti, complebuntur universa haec ".
DAN|12|8|Et ego audivi et non intellexi et dixi: " Domine mi, quid erit finis horum? ".
DAN|12|9|Et ait: " Vade, Daniel, quia clausi sunt signatique sermones usque ad tempus praefinitum.
DAN|12|10|Purificabuntur et dealbabuntur et probabuntur multi, et impie agent impii, neque intellegent omnes impii; porro docti intellegent.
DAN|12|11|Et a tempore, cum ablatum fuerit iuge sacrificium, et posita fuerit abominatio vastatoris, dies mille ducenti nonaginta.
DAN|12|12|Beatus, qui exspectat et pervenit usque ad dies mille trecentos triginta quinque.
DAN|12|13|Tu autem vade ad finem et requiesce; et stabis in sorte tua in fine dierum ".Hucusque Daniel in Hebraeo volumine legimus. Cetera, quae sequuntur usque ad finem libri, de Theodotionis editione translata sunt).
DAN|13|1|Et erat vir habitans in Ba bylone, et nomen eius Ioa chim;
DAN|13|2|et accepit uxorem nomine Susannam, filiam Helciae, pulchram nimis et timentem Dominum;
DAN|13|3|parentes enim illius, cum essent iusti, erudierunt filiam suam secundum legem Moysis.
DAN|13|4|Erat autem Ioachim dives valde, et erat ei pomerium vicinum domui suae; et ad ipsum confluebant Iudaei, eo quod esset honorabilior omnium.
DAN|13|5|Et constituti sunt de populo duo senes iudices in anno illo, de quibus locutus est Dominus quia egressa est iniquitas de Babylone a senibus iudicibus, qui videbantur regere populum.
DAN|13|6|Isti frequentabant domum Ioachim, et veniebant ad eos omnes, qui habebant iudicia.
DAN|13|7|Cum autem populus revertisset per meridiem, ingrediebatur Susanna et deambulabat in pomerio viri sui.
DAN|13|8|Et videbant eam duo senes cotidie ingredientem et deambulantem et facti sunt in concupiscentia eius
DAN|13|9|et everterunt sensum suum et declinaverunt oculos suos, ut non viderent caelum neque recordarentur iudiciorum iustorum.
DAN|13|10|Erant ergo ambo vulnerati amore eius nec indicaverunt sibi vicissim dolorem suum;
DAN|13|11|erubescebant enim indicare concupiscentiam suam, volentes concumbere cum ea.
DAN|13|12|Et observabant cotidie sollicitius videre eam. Dixitque alter ad alterum:
DAN|13|13|" Eamus domum, quia prandi hora est ". Et egressi recesserunt a se.
DAN|13|14|Cumque revertissent, venerunt in unum et, sciscitantes ab invicem causam, confessi sunt concupiscentiam suam; et tunc in commune statuerunt tempus, quando eam possent invenire solam.
DAN|13|15|Factum est autem, cum observarent diem aptum, ingressa est aliquando sicut heri et nudiustertius cum duabus solis puellis voluitque lavari in pomerio, aestus quippe erat.
DAN|13|16|Et non erat ibi quisquam, praeter duos senes absconditos et contemplantes eam.
DAN|13|17|Dixit ergo puellis: " Afferte mihi oleum et smegmata et ostia pomerii claudite, ut laver ".
DAN|13|18|Et fecerunt, sicut praeceperat; clauseruntque ostia pomerii et egressae sunt per posticium, ut afferrent, quae iusserat; nesciebantque senes intus esse absconditos.
DAN|13|19|Cum autem egressae essent puellae, surrexerunt duo senes et accurrerunt ad eam et dixerunt:
DAN|13|20|" Ecce ostia pomerii clausa sunt, et nemo nos videt, et in concupiscentia tui sumus; quam ob rem assentire nobis et commiscere nobiscum.
DAN|13|21|Quod si nolueris, dicemus testimonium contra te, quod fuerit tecum iuvenis et ob hanc causam emiseris puellas a te ".
DAN|13|22|Ingemuit Susanna et ait: " Angustiae sunt mihi undique: si enim hoc egero, mors mihi est; si autem non egero, non effugiam manus vestras;
DAN|13|23|sed melius mihi est absque opere incidere in manus vestras quam peccare in conspectu Domini ".
DAN|13|24|Et exclamavit voce magna Susanna; exclamaverunt autem et senes adversus eam,
DAN|13|25|et, cum cucurrisset unus, aperuit ostia pomerii.
DAN|13|26|Cum ergo audissent clamorem in pomerio famuli domus, irruerunt per posticam, ut viderent quidnam esset ei.
DAN|13|27|Postquam autem senes locuti sunt sermones suos, erubuerunt servi vehementer, quia numquam dictus fuerat sermo huiuscemodi de Susanna. Et factum est die crastina,
DAN|13|28|cum venisset populus ad virum eius Ioachim, venerunt et duo presbyteri pleni iniqua cogitatione adversum Susannam, ut interficerent eam;
DAN|13|29|et dixerunt coram populo: " Mittite ad Susannam, filiam Helciae, quae est uxor Ioachim "; et miserunt.
DAN|13|30|Et venit cum parentibus et filiis et universis cognatis suis.
DAN|13|31|Porro Susanna erat delicata nimis et pulchra specie.
DAN|13|32|At iniqui illi iusserunt, ut discooperiretur - erat enim cooperta - ut satiarentur decore eius.
DAN|13|33|Flebant igitur sui et omnes, qui videbant eam.
DAN|13|34|Consurgentes autem duo presbyteri in medio populi, posuerunt manus super caput eius;
DAN|13|35|quae flens suspexit ad caelum: erat enim cor eius fiduciam habens in Domino.
DAN|13|36|Et dixerunt presbyteri: " Cum deambularemus in pomerio soli, ingressa est haec cum duabus puellis et clausit ostia pomerii et dimisit puellas;
DAN|13|37|venitque ad eam adulescens, qui erat absconditus, et concubuit cum ea.
DAN|13|38|Porro nos cum essemus in angulo pomerii, videntes iniquitatem cucurrimus ad eos et vidimus eos commisceri.
DAN|13|39|Et illum quidem non quivimus comprehendere, quia fortior nobis erat et, apertis ostiis, exilivit.
DAN|13|40|Hanc autem cum apprehendissemus, interrogavimus, quisnam esset adulescens, et noluit indicare nobis. Huius rei testes sumus ".
DAN|13|41|Credidit eis multitudo quasi senibus populi et iudicibus, et condemnaverunt eam ad mortem.
DAN|13|42|Exclamavit autem voce magna Susanna et dixit: " Deus aeterne, qui absconditorum es cognitor, qui nosti omnia antequam fiant,
DAN|13|43|tu scis quoniam falsum contra me tulerunt testimonium; et ecce morior, cum nihil horum fecerim, quae isti malitiose composuerunt adversum me ".
DAN|13|44|Exaudivit autem Dominus vocem eius.
DAN|13|45|Cumque duceretur ad mortem, suscitavit Deus spiritum sanctum pueri iunioris, cuius nomen Daniel;
DAN|13|46|et exclamavit voce magna: " Innocens ego sum a sanguine huius ".
DAN|13|47|Et conversus omnis populus ad eum dixit: " Quis est iste sermo, quem tu locutus es? ".
DAN|13|48|Qui cum staret in medio eorum, ait: " Sic fatui, filii Israel? Non iudicantes neque, quod verum est, cognoscentes, condemnastis filiam Israel!
DAN|13|49|Revertimini ad iudicium, quia falsum testimonium locuti sunt adversum eam ".
DAN|13|50|Reversus est ergo omnis populus cum festinatione, et dixerunt ei senes: Veni et sede in medio nostrum et indica nobis, quia tibi dedit Deus honorem senectutis ".
DAN|13|51|Et dixit ad eos Daniel: " Separate illos ab invicem procul, et diiudicabo eos ".
DAN|13|52|Cum ergo divisi essent alter ab altero, vocavit unum de eis et dixit ad eum: " Inveterate dierum malorum, nunc venerunt peccata tua, quae operabaris prius,
DAN|13|53|iudicans iudicia iniusta, innocentes opprimens et dimittens noxios, dicente Domino: "Innocentem et iustum non interficies".
DAN|13|54|Nunc ergo, si vidisti eam, dic sub qua arbore videris eos loquentes sibi ". Qui ait: " Sub schino ".
DAN|13|55|Dixit autem Daniel: " Recte mentitus es in caput tuum; ecce enim angelus Dei, accepta sententia a Deo, scindet te medium ".
DAN|13|56|Et amoto eo, iussit adduci alium et dixit ei: " Semen Chanaan et non Iudae, species decepit te, et concupiscentia subvertit cor tuum.
DAN|13|57|Sic faciebatis filiabus Israel, et illae timentes loquebantur vobis, sed non filia Iudae sustinuit iniquitatem vestram.
DAN|13|58|Nunc ergo dic mihi sub qua arbore comprehenderis eos colloquentes sibi.Qui ait: " Sub prino ".
DAN|13|59|Dixit autem ei Daniel: " Recte mentitus es et tu in caput tuum; manet enim angelus Dei, gladium habens, ut secet te medium et interficiat vos ".
DAN|13|60|Exclamavit itaque omnis coetus voce magna et benedixerunt Deo, qui salvat sperantes in se.
DAN|13|61|Et consurrexerunt adversum duos presbyteros - convicerat enim eos Daniel ex ore suo falsum dixisse testimonium - feceruntque eis, sicut male egerant adversum proximum,
DAN|13|62|ut facerent secundum legem Moysis; et interfecerunt eos, et salvatus est sanguis innoxius in die illa.
DAN|13|63|Helcias autem et uxor eius laudaverunt Deum pro filia sua Susanna, cum Ioachim marito eius et cognatis omnibus, quia non esset inventa in ea res turpis.
DAN|13|64|Daniel autem factus est magnus in conspectu populi a die illa et deinceps.
DAN|14|1|Et rex Astyages appositus est ad patres suos, et suscepit Cyrus Perses regnum eius.
DAN|14|2|Erat autem Daniel conviva regis et honoratus super omnes amicos eius.
DAN|14|3|Erat quoque idolum nomine Bel apud Babylonios, ct impendebantur in eo per dies singulos similae artabae duodecim et oves quadraginta vinique metretae sex.
DAN|14|4|Rex quoque colebat eum et ibat per singulos dies adorare eum; porro Daniel adorabat Deum suum. Dixitque ei rex: " Quare non adoras Bel? ".
DAN|14|5|Qui respondens ait ei: " Quia non colo idola manufacta sed viventem Deum, qui creavit caelum et terram et habet potestatem omnis carnis ".
DAN|14|6|Et dixit ad eum rex: "Non tibi videtur esse Bel vivens deus? An non vides, quanta comedat et bibat cotidie? ".
DAN|14|7|Et ait Daniel arridens: " Ne erres, rex; iste enim intrinsecus luteus est et forinsecus aereus, neque comedit neque bibit aliquando ".
DAN|14|8|Et iratus rex vocavit sacerdotes eius et ait eis: " Nisi dixeritis mihi, quis est qui comedat impensas has, moriemini;
DAN|14|9|si autem ostenderitis quoniam Bel comedat haec, morietur Daniel, quia blasphemavit in Bel ". Et dixit Daniel regi: " Fiat iuxta verbum tuum ".
DAN|14|10|Erant autem sacerdotes Bel septuaginta, exceptis uxoribus et parvulis et filiis. Et venit rex cum Daniele in templum Belis.
DAN|14|11|Et dixerunt sacerdotes Belis: " Ecce nos egredimur foras; et tu, rex, affer escas et vinum miscens pone et claude ostium et signa anulo tuo;
DAN|14|12|et, cum ingressus fueris mane, nisi inveneris omnia comesta a Bel, morte moriemur, vel Daniel, qui mentitus est adversum nos ".
DAN|14|13|Contemnebant autem, quia fecerant sub mensa absconditum introitum et per illum ingrediebantur semper et devorabant ea.
DAN|14|14|Factum est igitur, postquam egressi sunt illi, et rex posuit cibos ante Bel; et praecepit Daniel pueris suis, et attulerunt cinerem et cribraverunt per totum templum coram rege solo et egressi clauserunt ostium et signantes anulo regis abierunt.
DAN|14|15|Sacerdotes autem ingressi sunt nocte iuxta consuetudinem suam et uxores et filii eorum et comederunt omnia et biberunt.
DAN|14|16|Surrexit autem rex primo diluculo, et Daniel cum eo;
DAN|14|17|et ait rex: " Salvane sunt signa, Daniel? ". Qui respondit: " Salva, rex ".
DAN|14|18|Statimque cum aperuisset ostium, intuitus rex mensam, exclamavit voce magna: " Magnus es, Bel, et non est apud te dolus quisquam ".
DAN|14|19|Et risit Daniel et tenuit regem, ne ingrederetur intro, et dixit: " Ecce pavimentum; animadverte, cuius vestigia sunt haec ".
DAN|14|20|Et dixit rex: " Video vestigia virorum et mulierum et infantium ". Et iratus est rex.
DAN|14|21|Tunc apprehendit sacerdotes et uxores et filios eorum, et ostenderunt ei abscondita ostiola, per quae ingrediebantur et consumebant, quae erant super mensam.
DAN|14|22|Occidit ergo illos rex et tradidit Bel in potestate Danieli, qui subvertit eum et templum eius.
DAN|14|23|Et erat draco magnus, et colebant eum Babylonii.
DAN|14|24|Et dixit rex Danieli: " Non potes dicere quia iste non sit deus vivens; adora ergo eum ".
DAN|14|25|Dixitque Daniel: " Dominum Deum meum adoro, quia ipse est Deus vivens.
DAN|14|26|Tu autem, rex, da mihi potestatem, et interficiam draconem absque gladio et fuste ". Et ait rex: " Do tibi ".
DAN|14|27|Tulit ergo Daniel picem et adipem et pilos et coxit pariter; fecitque massas et dedit in os draconis et, cum comedisset, diruptus est draco. Et dixit: " Ecce quae colebatis ".
DAN|14|28|Cum audissent Babylonii, indignati sunt vehementer et congregati adversum regem dixerunt: "Iudaeus factus est rex; Bel destruxit, draconem interfecit et sacerdotes occidit ".
DAN|14|29|Et dixerunt, cum venissent ad regem: " Trade nobis Danielem; alioquin interficiemus te et domum tuam ".
DAN|14|30|Vidit ergo rex quod irruerent in eum vehementer et, necessitate compulsus, tradidit eis Danielem.
DAN|14|31|Qui miserunt eum in lacum leonum, et erat ibi diebus sex.
DAN|14|32|Porro in lacu erant septem leones, et dabantur eis cotidie duo corpora et duae oves; et tunc non data sunt eis, ut devorarent Danielem.
DAN|14|33|Erat autem Abacuc propheta in Iudaea et ipse coxerat pulmentum et intriverat panes in alveolo et ibat in campum, ut ferret messoribus.
DAN|14|34|Dixitque angelus Domini ad Abacuc: " Fer prandium, quod habes, in Babylonem Danieli, qui est in lacu leonum ".
DAN|14|35|Et dixit Abacuc: " Domine, Babylonem non vidi et lacum nescio ".
DAN|14|36|Et apprehendit eum angelus Domini in vertice eius et portavit eum capillo capitis sui posuitque eum in Babylone supra lacum in impetu spiritus sui.
DAN|14|37|Et clamavit Abacuc dicens: " Daniel, Daniel, tolle prandium, quod misit tibi Deus ".
DAN|14|38|Et ait Daniel: "Recordatus es enim mei, Deus, et non dereliquisti diligentes te ".
DAN|14|39|Surgensque Daniel comedit. Porro angelus Dei restituit Abacuc confestim in loco suo.
DAN|14|40|Venit ergo rex die septima, ut lugeret Danielem; et venit ad lacum et introspexit, et ecce Daniel sedens.
DAN|14|41|Et exclamavit rex voce magna dicens: "Magnus es, Domine, Deus Danielis, et non est alius praeter te ".
DAN|14|42|Porro illos, qui perditionis eius causa fuerant, intromisit in lacum; et devorati sunt in momento coram eo.
HOS|1|1|Verbum Domini, quod factum est ad Osee filium Beeri in die bus Oziae, Ioatham, Achaz, Ezechiae regum Iudae, et in diebus Ieroboam filii Ioas regis Israel.
HOS|1|2|Principium verbi Domini per Osee. Dixit Dominus ad Osee: Vade, sume tibi mulierem fornicationumet filios fornicationum,quia fornicans fornicatur terra a Domino ".
HOS|1|3|Et abiit et accepit Gomer filiam Debelaim, quae concepit et peperit ei filium.
HOS|1|4|Et dixit Dominus ad eum: " Voca nomen eius 'Iezrahel', quoniam adhuc modicum et visitabo sanguinem Iezrahel super domum Iehu et cessare faciam regnum domus Israel;
HOS|1|5|et in illa die conteram arcum Israel in valle Iezrahel ".
HOS|1|6|Et concepit adhuc et peperit filiam; et dixit ei: " Voca nomen eius Absque misericordia", quia non addam ultra misereri domui Israel, ut ignoscam eis.
HOS|1|7|Et domui Iudae miserebor et salvabo eos in Domino Deo suo et non salvabo eos in arcu et gladio et in bello et in equis et in equitibus ".
HOS|1|8|Et ablactavit eam, quae erat 'Absque misericordia', et concepit et peperit filium.
HOS|1|9|Et dixit: " Voca nomen eius 'Non populus meus', quia vos non populus meus, et ego 'Non sum' vobis.
HOS|2|1|Et erit numerus filiorum Israelquasi arena maris,quae sine mensura est et non numerabitur.Et erit: in loco, ubi dicebatur eis:Non populus meus vos",dicetur eis: "Filii Dei viventis".
HOS|2|2|Et congregabuntur filii Iudaeet filii Israel pariteret ponent sibimet caput unumet ascendent de terra,quia magnus dies Iezrahel.
HOS|2|3|Dicite fratribus vestris: "Populus meus"et sororibus vestris: "Misericordiam consecuta".
HOS|2|4|Contendite adversum matrem vestram; contendite,quoniam ipsa non uxor mea,et ego non vir eius;auferat fornicationes suas a facie suaet adulteria sua de medio uberum suorum,
HOS|2|5|ne forte exspoliem eam nudamet statuam eam secundum diem nativitatis suaeet ponam eam quasi solitudinemet statuam eam velut terram aridamet interficiam eam siti.
HOS|2|6|Et filiorum illius non miserebor,quoniam filii fornicationum sunt,
HOS|2|7|quia fornicata est mater eorum,turpiter egit, quae concepit eos;quia dixit: "Vadam post amatores meos,qui dant panes mihi et aquas meas,lanam meam et linum meum,oleum meum et potum meum".
HOS|2|8|Propter hoc ecce ego saepiamviam tuam spiniset saepiam eam maceria,et semitas suas non inveniet;
HOS|2|9|et sequetur amatores suoset non apprehendet eos;et quaeret eos et non invenietet dicet: "Vadam et revertarad virum meum priorem,quia bene mihi erat tunc magis quam nunc".
HOS|2|10|Et haec nescivit quia egodedi ei frumentum et vinum et oleumet argentum multiplicavi eiet aurum, quae fecerunt Baal.
HOS|2|11|Idcirco convertar et sumamfrumentum meum in tempore suoet vinum meum in tempore suo;et auferam lanam meam et linum meum,quae operiebant pudenda eius,
HOS|2|12|et nunc revelabo ignominiam eiusin oculis amatorum eius,et nullus est qui eruat eam de manu mea.
HOS|2|13|Et cessare faciam omne gaudium eius,sollemnitatem eius, neomeniam eius,sabbatum eius et omnia festa tempora eius;
HOS|2|14|et corrumpam vineam eius et ficum eius,de quibus dixit: "Mercedes hae meae sunt,quas dederunt mihi amatores mei".Et ponam eas in saltum,et comedet illas bestia agri.
HOS|2|15|Et visitabo super eam dies Baalim,quibus accendebat incensumet ornabatur inaure sua et monili suoet ibat post amatores suos,sed mei obliviscebatur,dicit Dominus.
HOS|2|16|Propter hoc ecce ego lactabo eamet ducam eam in solitudinemet loquar ad cor eius;
HOS|2|17|et dabo ei vineas eius ex eodem locoet vallem Achor, portam spei,et respondebit ibiiuxta dies iuventutis suaeet iuxta dies ascensionis suae de terra Aegypti.
HOS|2|18|Et erit: in die illa,ait Dominus,vocabis me: "Vir meus"et non vocabis me ultra: "Baal meus".
HOS|2|19|Et auferam nomina Baalim de ore eius,et non recordabitur ultra nominis eorum.
HOS|2|20|Et percutiam eis foedus in die illacum bestia agri et cum volucre caeli et cum reptili terrae;et arcum et gladium et bellumconteram de terraet cubare eos faciam confidenter.
HOS|2|21|Et sponsabo te mihi in sempiternum;et sponsabo te mihi in iustitia et iudicioet in misericordia et miserationibus.
HOS|2|22|Et sponsabo te mihi in fide,et cognosces Dominum.
HOS|2|23|Et erit: in illa die exaudiam,dicit Dominus,exaudiam caelos,et illi exaudient terram;
HOS|2|24|et terra exaudiettriticum et vinum et oleum,et haec exaudient Iezrahel.
HOS|2|25|Et seminabo eam mihi in terramet miserebor eius, quae fuit "Absque misericordia";
HOS|2|26|et dicam "Non populo meo": "Populus meus tu";et ipse dicet: "Deus meus es tu" ".
HOS|3|1|Et dixit Dominus ad me: " Adhuc vade, dilige mulierem dilectam amico et adulteram, sicut diligit Dominus filios Israel, et ipsi respectant ad deos alienos et diligunt placentas uvarum ".
HOS|3|2|Et emi eam mihi quindecim argenteis et choro hordei et dimidio choro hordei.
HOS|3|3|Et dixi ad eam: " Dies multos exspectabis me; non fornicaberis et non eris viro, neque ibo ego ad te ".
HOS|3|4|Quia dies multos sedebunt filii Israel sine rege et sine principe et sine sacrificio et sine lapide et sine ephod et sine theraphim.
HOS|3|5|Et post haec revertentur filii Israel et quaerent Dominum Deum suum et David regem suum et pavebunt ad Dominum et ad bonum eius in fine dierum.
HOS|4|1|" Audite verbum Domini,filii Israel,quia iudicium Dominocum habitatoribus terrae:non est enim veritas, et non est benignitas,et non est scientia Dei in terra;
HOS|4|2|maledictum et mendaciumet homicidium et furtum et adulterium inundaverunt,et sanguis sanguinem tetigit.
HOS|4|3|Propter hoc lugebit terra,et infirmabitur omnis, qui habitat in ea,cum bestia agri et volucre caeli,sed et pisces maris auferentur.
HOS|4|4|Verumtamen non sit qui contendatnec qui arguat,sed tecum iudicium meum, sacerdos.
HOS|4|5|Et corrues plena die,et corruet etiam propheta tecum nocte;et perdam matrem tuam.
HOS|4|6|Perit populus meus,eo quod non habuerit scientiam.Quia tu scientiam reppulisti,repellam te, ne sacerdotio fungaris mihi;et quia oblitus es legis Dei tui,obliviscar filiorum tuorum et ego.
HOS|4|7|Secundum multitudinem eorum, sic peccaverunt mihi;gloriam eorum in ignominiam commutabo.
HOS|4|8|Peccatum populi mei comeduntet ad iniquitatem eorum sublevabunt animas eorum.
HOS|4|9|Et erit sicut populus sic sacerdos;et visitabo super eum vias eiuset opera eius reddam ei.
HOS|4|10|Et comedent et non saturabuntur;fornicabuntur et non multiplicabuntur,quoniam Dominum reliqueruntin non custodiendo.
HOS|4|11|Fornicatio et vinum et ebrietas auferunt cor.
HOS|4|12|Populus meus in ligno suo interrogat,et baculus eius annuntiat ei;spiritus enim fornicationum decepit eos,et fornicantur a Deo suo.
HOS|4|13|Super capita montium sacrificantet super colles accendunt thymiama,subtus quercum et populum et terebinthum,quia bona est umbra eius;ideo fornicantur filiae vestrae,et sponsae vestrae adulterae sunt.
HOS|4|14|Non visitabo super filias vestras,cum fuerint fornicatae,et super sponsas vestras,cum adulteraverint,quoniam hi ipsi cum meretricibus seceduntet cum prostibulis delubrorum sacrificant,et populus non intellegens corruet.
HOS|4|15|Si fornicaris tu, Israel,non delinquat saltem Iuda;et nolite ingredi in Galgalaet ne ascenderitis in Bethavenneque iuraveritis: "Vivit Dominus".
HOS|4|16|Quoniam sicut vacca lasciviensIsrael contumax est;nunc pascet eos Dominusquasi agnum in latitudine?
HOS|4|17|Particeps idolorum Ephraim,dimitte eum.
HOS|4|18|Transiit convivium eorum,fornicatione fornicati sunt,diligunt vehementerignominiam impudicitiae.
HOS|4|19|Ligabit spiritus eos in alis suis,et confundentur a sacrificiis suis.
HOS|5|1|Audite hoc, sacerdotes,et attendite, domus Israel;et domus regis, auscultate,quia vobis iudicium est;quoniam laqueus facti estis pro Masphaet rete expansum super Thabor.
HOS|5|2|Et foveam Settim profundam fecerunt;ego autem castigabo vos omnes.
HOS|5|3|Ego scio Ephraim,et Israel non est absconditus a me;quia nunc fornicatus es, Ephraim,contaminatus est Israel.
HOS|5|4|Non dabunt opera sua,ut revertantur ad Deum suum,quia spiritus fornicationis in medio eorum,et Dominum non cognoverunt.
HOS|5|5|Et testatur arrogantia Israel in faciem suam,et Israel et Ephraim ruent in iniquitate sua:ruet etiam Iudas cum eis.
HOS|5|6|In gregibus suis et in armentis suisvadent ad quaerendum Dominumet non invenient;subtraxit se ab eis.
HOS|5|7|In Dominum praevaricati sunt,quia filios alienos genuerunt;nunc devorabit eos uno mense cum partibus suis.
HOS|5|8|Clangite bucina in Gabaa,tuba in Rama,conclamate in Bethaven,exterrete Beniamin.
HOS|5|9|Ephraim vastabitur in die correptionis;in tribubus Israel annuntio rem certam.
HOS|5|10|Facti sunt principes Iudaequasi transferentes terminos;super eos effundamquasi aquam iram meam.
HOS|5|11|Oppressus est Ephraim,fractum est ius,quoniam voluit abire post sordem.
HOS|5|12|Et ego quasi sanies Ephraim,et quasi putredo domui Iudae.
HOS|5|13|Et vidit Ephraim languorem suum,et Iuda ulcus suum;et abiit Ephraim ad Assyriamet misit ad regem magnum;sed et ipse non poterit sanare vosnec solvere poterit vos ab ulcere.
HOS|5|14|Quoniam ego quasi leaena Ephraimet quasi catulus leonis domui Iudae;ego, ego capiam et vadam,tollam, et non est qui eruat.
HOS|5|15|Vadens revertar ad locum meum,donec poenas solvantet quaerant faciem meam,in tribulatione sua me desiderent.
HOS|6|1|"Venite, et revertamur ad Do minum,quia ipse laceravit et sanabit nos,percussit et curabit nos.
HOS|6|2|Vivificabit nos post duos dies,in die tertia suscitabit nos,et vivemus in conspectu eius.
HOS|6|3|Sciamus sequamurque,ut cognoscamus Dominum.Quasi diluculum praeparatus est egressus eius,et veniet quasi imber nobis temporaneus,quasi imber serotinus irrigans terram".
HOS|6|4|Quid faciam tibi, Ephraim?Quid faciam tibi, Iuda?Caritas vestra quasi nubes matutinaet quasi ros mane pertransiens.
HOS|6|5|Propter hoc dolavi per prophetas,occidi eos in verbis oris mei,sed ius meum quasi lux egredietur;
HOS|6|6|quia caritatem volo et non sacrificium,et scientiam Dei plus quam holocausta.
HOS|6|7|Ipsi autem in Adam transgressi sunt pactum;ibi praevaricati sunt in me.
HOS|6|8|Galaad civitas operantium iniquitatemmaculata sanguine.
HOS|6|9|Et quasi insidiantes virum latronescaterva sacerdotum;in via interficiunt pergentes Sichem,vere scelus operantur.
HOS|6|10|In domo Israel vidi horrendum:ibi fornicationes Ephraim,contaminatus est Israel.
HOS|6|11|Sed et tibi, Iuda, parata est messis,cum convertero sortem populi mei.
HOS|7|1|Cum sanare vellem Israel,revelata est iniquitas Ephraimet malitia Samariae,quia operati sunt mendacium;et fur ingressus est,foris autem spoliat turma latronum.
HOS|7|2|Et non dicunt in cordibus suisomnem malitiam eorum me recordari.Nunc circumdederunt eos opera sua,coram facie mea facta sunt.
HOS|7|3|In malitia sua laetificaverunt regem et in mendaciis suis principes.
HOS|7|4|Omnes adulterantes;quasi clibanus succensus illi,pistor cessat excitare ignema commixtione fermenti, donec fermentetur totum.
HOS|7|5|Die regis nostriinfirmi facti sunt principes ardore vini,quod apprehendit protervos.
HOS|7|6|Quia applicuerunt quasi clibanum cor suumin insidiando;tota nocte dormivit ira eorum,mane ipsa ardet quasi ignis flammae.
HOS|7|7|Omnes calefacti sunt quasi clibanuset devorant iudices suos.Omnes reges eorum ceciderunt;non est qui clamet in eis ad me.
HOS|7|8|Ephraim in populis ipse commiscebatur;Ephraim factus est subcinericius panis, qui non reversatur.
HOS|7|9|Comederunt alieni robur eius,et ipse nescit;sed et cani effusi sunt in eo,et ipse ignorat.
HOS|7|10|Et testatur superbia Israel in faciem suam,nec reversi sunt ad Dominum Deum suumet non quaesierunt eum in omnibus his.
HOS|7|11|Et factus est Ephraim quasi columbainsipiens non habens sensum:Aegyptum invocabant,ad Assyrios abierunt.
HOS|7|12|Et cum profecti fuerint,expandam super eos rete meum;quasi volucrem caeli detraham eos, corripiam eos secundum auditionem coetus eorum.
HOS|7|13|Vae eis, quoniam recesserunt a me!Vastabuntur, quia praevaricati sunt in me.Et ego redimam eos,cum ipsi locuti sint contra me mendacia?
HOS|7|14|Et non clamaverunt ad me in corde suo,sed ululabant in cubilibus suis;super triticum et vinum se incidebant,contumaces sunt adversum me.
HOS|7|15|Et ego erudivi eos et confortavi brachia eorum,et in me cogitaverunt malitiam.
HOS|7|16|Convertuntur ad eum, qui non prodest,facti sunt quasi arcus dolosus;cadent in gladio principes eorumpropter execrationem linguae suae: ista subsannatio eorum in terra Aegypti.
HOS|8|1|In gutture tuo sit tuba!Quasi aquila super domum Do minipro eo quod transgressi sunt foedus meumet legem meam praevaricati sunt.
HOS|8|2|Me invocant: "Deus meus";cognovimus te, Israel.
HOS|8|3|Proiecit Israel bonum;inimicus persequetur eum.
HOS|8|4|Ipsi constituerunt reges, et non ex me;principes constituerunt, et non cognovi:argentum suum et aurum suumfecerunt sibi idola,ut interirent.
HOS|8|5|Proiectus est vitulus tuus, Samaria;iratus est furor meus in eos.Usquequo non poterunt emundari?
HOS|8|6|Quia ex Israel et ipse est:artifex fecit illum,et non est Deus;quoniam in scintillas eritvitulus Samariae.
HOS|8|7|Quia ventum seminabuntet turbinem metent;cum culmus non sit in eo,germen non faciet farinam:quod et si fecerit,alieni comedent eam.
HOS|8|8|Devoratus est Israel,nunc factus est in nationibusquasi vas immundum.
HOS|8|9|Quia ipsi ascenderunt ad Assyriam, onager est solitarius sibi;Ephraim autem munera dederunt amatoribus.
HOS|8|10|Sed et cum mercede conduxerint nationes,nunc compellam eos,et trement paulisper sub onere regis principum.
HOS|8|11|Cum multiplicaret Ephraim altaria pro peccato,factae sunt ei arae in peccatum.
HOS|8|12|Scribebam ei multiplices leges meas;velut alienae computatae sunt.
HOS|8|13|Hostias amant,immolant carnes et comedunt;sed Dominus non suscipiet eas.Nunc recordabitur iniquitatis eorumet visitabit peccata eorum:ipsi in Aegyptum convertentur.
HOS|8|14|Et oblitus est Israel factoris suiet aedificavit delubra;et Iudas multiplicavit urbes munitas.Et mittam ignem in civitates eius,et devorabit aedes illius.
HOS|9|1|Noli laetari, Israel;noli exsultare sicut populi,quia fornicatus es a Deo tuo,dilexisti mercedem super omnes areas tritici.
HOS|9|2|Area et torcular non pascet eos,et vinum mentietur eis.
HOS|9|3|Non manebunt in terra Domini:revertetur Ephraim in Aegyptum,et in Assyria pollutum comedent.
HOS|9|4|Non libabunt Domino vinum,et non placebunt ei sacrificia eorum;quasi panis lugentium erunt eis:omnes, qui comedent eum, contaminabuntur,quia panis eorum erit tantummodo pro vita ipsorum;non intrabit in domum Domini.
HOS|9|5|Quid facietis in die sollemni,in die festivitatis Domini?
HOS|9|6|Ecce enim profecti sunt a vastitate;Aegyptus congregabit eos,Memphis sepeliet eos:desiderabile argentum eorumurtica hereditabit,spina in tabernaculis eorum.
HOS|9|7|Venerunt dies visitationis,venerunt dies retributionis:sciat Israel!Stultus - clamet - est propheta;insanus vir spiritalis".Secundum multitudinem iniquitatis tuaemultae sunt inimicitiae tuae.
HOS|9|8|Speculatur Ephraim, populus Dei mei, prophetam;laqueus aucupis super omnes vias eius,inimicitiae in ipsa domo Dei eius.
HOS|9|9|Profunde peccaveruntsicut in diebus Gabaa;recordabitur iniquitatis eorumet visitabit peccata eorum.
HOS|9|10|Quasi uvas in desertoinveni Israel,quasi prima poma ficulneae in initio eiusvidi patres vestros;ipsi autem intraverunt ad Baalphegoret se consecraverunt Confusioniet facti sunt abominabilessicut id, quod dilexerunt.
HOS|9|11|Ephraim quasi avis avolabit gloria eorum,a partu et ab utero et a conceptu.
HOS|9|12|Quod si et enutrierint filios suos,absque liberis eos faciam, absque hominibus;sed et vae eis,cum recessero ab eis!
HOS|9|13|Ephraim, ut vidi, in venationem posuit sibi filios suos,et Ephraim educit ad interfectorem filios suos.
HOS|9|14|"Da eis, Domine! Quid dabis eis?Da eis vulvam sine liberis et ubera arentia!".
HOS|9|15|Omnes nequitiae eorum in Galgala,profecto ibi exosos habui eos.Propter malitiam operum eorumde domo mea eiciam eos.Non addam ut diligam eos;omnes principes eorum rebelles.
HOS|9|16|Percussus est Ephraim,radix eorum exsiccata est,fructum nequaquam facient;quod si et genuerint,interficiam amantissima uteri eorum ".
HOS|9|17|Abiciet eos Deus meus,quia non audierunt eum;et erunt vagi in nationibus.
HOS|10|1|Vitis frondosa Israel,fructum producens sibi;secundum multitudinem fructus sui multiplicavit altaria,iuxta ubertatem terrae suaedecoravit simulacra.
HOS|10|2|Divisum est cor eorum,nunc poenas solvent;ipse confringet aras eorum,depopulabitur simulacra eorum.
HOS|10|3|Profecto nunc dicent: Non est rex nobis;non enim timemus Dominum,et rex quid faciet nobis? ".
HOS|10|4|Loqui verba, iurare in vanum,ferire foedus;et germinabit quasi venenum iussuper sulcos agri.
HOS|10|5|De vitulo Bethaventrement habitatores Samariae;quia luget super eum populus eius;dum sacerdotes eius super eumexsultant in gloria eius;vere migrabit ab eo.
HOS|10|6|Siquidem et ipse in Assyriam delatus est,munus regi magno;confusio Ephraim capiet,et confundetur Israel in consilio suo.
HOS|10|7|Perit Samaria,rex eius quasi festuca super faciem aquae.
HOS|10|8|Et disperdentur excelsa impietatis,peccatum Israel;spina et tribulus ascendetsuper aras eorum,et dicent montibus: " Operite nos! "et collibus: " Cadite super nos! ".
HOS|10|9|Ex diebus Gabaa peccavit Israel;ibi perstiterunt.Non comprehendet eos in Gabaaproelium super filios iniquitatis?
HOS|10|10|" Iuxta desiderium meum corripiam eos;congregabuntur super eos populi,cum corripientur propter duas iniquitates suas.
HOS|10|11|Ephraim vitula docta,diligens trituram.Et ego transivi super pulchritudinem colli eius;iunxi Ephraim aratro,arabit Iudas,sarriet sibi Iacob.
HOS|10|12|Seminate vobis in iustitia,metite secundum caritatem;innovate vobis novale.Tempus est requirendi Dominum,donec veniat, ut pluat vobis iustitiam.
HOS|10|13|Arastis impietatem,iniquitatem messuistis,comedistis frugem mendacii,quia confisus es in curribus tuis,in multitudine fortium tuorum.
HOS|10|14|Consurget tumultus in populo tuo,et omnes munitiones tuae vastabuntur,sicut vastavit Salman Betharbeelin die proelii,matre super filios allisa.
HOS|10|15|Sic faciet vobis Bethelpropter maximam nequitiam vestram.Mane interibit rex Israel.
HOS|11|1|Cum puer esset Israel, dilexi eumet ex Aegypto vocavi filium meum.
HOS|11|2|Quanto magis vocabam eos,tanto recesserunt a facie mea;ipsi Baalim immolabantet simulacris sacrificabant.
HOS|11|3|Et ego dirigebam gressus Ephraim,portabam eos in brachiis meis,et nescierunt quod curarem eos.
HOS|11|4|In funiculis humanitatis trahebam eos,in vinculis caritatis;et fui eis, quasi qui elevant infantem ad maxillas suas,et declinavi ad eum, ut vesceretur.
HOS|11|5|Revertetur in terram Aegypti,et Assur ipse rex eius,quoniam noluerunt converti.
HOS|11|6|Saeviet gladius in civitatibus eiuset consumet garrulos eiuset comedet eos propter consilia eorum.
HOS|11|7|Populus meus pendet ad praevaricandum contra me;vocant eum ad altum, sed simul non erigunt eum.
HOS|11|8|Quomodo dabo te, Ephraim,tradam te, Israel?Quomodo dabo te sicut Adama,ponam te ut Seboim?Convertitur in me cor meum,simul exardescit miseratio mea.
HOS|11|9|Non faciam furorem irae meae,non convertar, ut disperdam Ephraim,quoniam Deus egoet non homo,in medio tui Sanctuset non veniam in terrore.
HOS|11|10|Post Dominum ambulabunt;quasi leo rugiet,quia ipse rugiet,et in tremore accurrent filii ab occidente.
HOS|11|11|Et avolabunt quasi avis ex Aegyptoet quasi columba de terra Assyriae;et collocabo eos in domibus suis,dicit Dominus.
HOS|12|1|Circumdedit me in fraude Ephraim,et in dolo domus Israel;C Iudas autem, dum adhuc vagatur, est cum Deoet cum Sancto fidelis " C.
HOS|12|2|Ephraim pascit ventumet sequitur aestum;tota die mendacium et violentiam multiplicatet foedus cum Assyriis initet oleum in Aegyptum fert.
HOS|12|3|Iudicium ergo Domini cum Iuda,et visitatio super Iacob;iuxta vias eius et iuxta opera eius reddet ei.
HOS|12|4|In utero supplantavit fratrem suumet in robore suo luctatus est cum Deo.
HOS|12|5|Et luctatus est cum angelo et praevaluit;flevit et deprecatus est eum.In Bethel invenit eumet ibi locutus est nobiscum
HOS|12|6|Dominus, Deus exercituum:Dominus memoriale eius.
HOS|12|7|" Et tu ad Deum tuum converteris;caritatem et iudicium custodiet spera in Deo tuo semper ".
HOS|12|8|Chanaan, in manu eius statera dolosa,fraudem diligit.
HOS|12|9|Et dixit Ephraim: " Verumtamen dives effectus sum,inveni opes mihi,omnes labores mei non invenient mihiiniquitatem, quam peccavi ".
HOS|12|10|" Ego autem Dominus, Deus tuusex terra Aegypti;adhuc sedere te faciam in tabernaculis,sicut in diebus conventus.
HOS|12|11|Et loquar ad prophetaset ego visionem multiplicaboet in manu prophetarum proponam similitudines ".
HOS|12|12|Si Galaad iniquitas fuerat,prorsus inanes facti sunt;in Galgala bobus immolantes,etiam altaria eorum erunt quasi acervisuper sulcos agri.
HOS|12|13|Fugit Iacob in regionem Aram;et servivit Israel pro uxoreet pro uxore custos fuit.
HOS|12|14|Per prophetam autem eduxit DominusIsrael de Aegypto,et per prophetam custoditus est.
HOS|12|15|Ad iracundiam provocavit Ephraim amarissime,sed sanguinem eius super eum relinquetet opprobrium eius retribuet ei Dominus suus.
HOS|13|1|Loquente Ephraim, horror factus est;dux erat in Israel.Et deliquit in Baalet mortuus est.
HOS|13|2|Et nunc addunt ad peccandumfaciuntque sibi conflatile de argento suo,secundum intellegentiam suam simulacra;factura artificum totum est. His - ipsi dicunt - immolate! ".Homines vitulos osculantur.
HOS|13|3|Idcirco erunt quasi nubes matutinaet sicut ros matutinus praeteriens,sicut palea turbine rapta ex areaet sicut fumus de fumario.
HOS|13|4|" Ego autem Dominus, Deus tuusex terra Aegypti;et Deum absque me nescies,et salvator non est praeter me.
HOS|13|5|Ego pavi te in deserto,in terra ardenti solitudinis.
HOS|13|6|Iuxta pascua sua saturati suntet saturati elevaverunt cor suum,propterea obliti sunt mei.
HOS|13|7|Et ego ero eis quasi leaena,sicut pardus iuxta viam insidiabor.
HOS|13|8|Occurram eis quasi ursa, raptis catulis,et dirumpam claustrum cordis eorum:et consumam eos ibi quasi leo;bestia agri scindet eos.
HOS|13|9|Perdo te, Israel;quis est auxiliator tuus?
HOS|13|10|Ubinam est rex tuus,ut salvet te in omnibus urbibus tuis,et iudices tui, de quibus dixisti:Da mihi regem et principes"?
HOS|13|11|Do tibi regem in furore meoet aufero in indignatione mea.
HOS|13|12|Colligata est iniquitas Ephraim,absconditum peccatum eius.
HOS|13|13|Dolores parturientis venient ei;erit filius non sapiens:suo enim tempore non stabitin ore vulvae.
HOS|13|14|De manu inferni liberabo eos,de morte redimam eos?Ubi pestilentiae tuae, o mors?Ubi pestis tua, inferne?Consolatio abscondita est ab oculis meis ".
HOS|13|15|Dum ipse inter fratres fructificat,veniet ventus urens, ventus Dominide deserto ascendens,et siccabit venas eiuset desolabit fontem eius.Ipse diripiet thesaurum,omne vas desiderabile.
HOS|14|1|Poenas solvet Samaria,quoniam rebellavit contra Deum suum:in gladio peribunt,parvuli eorum elidentur,et praegnantes discindentur.
HOS|14|2|Convertere, Israel, ad Dominum Deum tuum,quoniam corruisti in iniquitate tua.
HOS|14|3|Tollite vobiscum verbaet convertimini ad Dominum;dicite ei: " Omnem aufer iniquitatemet accipe bonum,et reddemus fructum labiorum nostrorum.
HOS|14|4|Assyria non salvabit nos;super equum non ascendemusnec vocabimus ultra: "Deos nostros!"opera manuum nostrarum,quia in te misericordiam consequetur pupillus ".
HOS|14|5|" Sanabo praevaricationem eorum,diligam eos spontanee,quia aversus est furor meus ab eis.
HOS|14|6|Ero quasi ros pro Israel;germinabit quasi liliumet mittet radices suas ut Libanus.
HOS|14|7|Expandentur rami eius;et erit quasi oliva gloria eius,et odor eius ut Libani.
HOS|14|8|Convertentur sedentes in umbra mea,colent triticumet germinabunt quasi vinea;memoriale eius sicut vinum Libani.
HOS|14|9|Ephraim, quid ei ultra idola?Ego exaudio et respicio in eum.Ego ut abies virens:ex me fructus tuus invenitur ".
HOS|14|10|Qui sapiens est, intellegat ista;intellegens sciat haec!Quia rectae viae Domini,et iusti ambulabunt in eis;praevaricatores vero corruent in eis.
JOEL|1|1|Verbum Domini, quod factum est ad loel filium Phatuel.
JOEL|1|2|Audite hoc, senes,et auribus percipite, omnes habitatores terrae,si factum est istud in diebus vestrisaut in diebus patrum vestrorum.
JOEL|1|3|Super hoc filiis vestris narrate,et filii vestri filiis suis,et filii eorum generationi alterae.
JOEL|1|4|Residuum erucae comedit locusta,et residuum locustae comedit bruchus,et residuum bruchi comedit gryllus.
JOEL|1|5|Expergiscimini, ebrii, et flete,et ululate, omnes, qui bibitis vinum,propter mustum,quoniam periit ab ore vestro.
JOEL|1|6|Gens enim ascendit super terram meamfortis et innumerabilis;dentes eius ut dentes leonis,et molares leaenae sunt ei.
JOEL|1|7|Posuit vineam meam in desertumet ficum meam in lignum confractum;nudans spoliavit eam et proiecit,albi facti sunt rami eius.
JOEL|1|8|Plange, quasi virgo accincta saccosuper virum pubertatis suae.
JOEL|1|9|Periit oblatio et libatiode domo Domini;luxerunt sacerdotesministri Domini.
JOEL|1|10|Depopulata est regio;luxit humus,quoniam devastatum est triticum,defecit mustum,elanguit oleum.
JOEL|1|11|Confundemini, agricolae,ululate, vinitores,super frumento et hordeo,quia periit messis agri.
JOEL|1|12|Vinea exaruit,et ficus elanguit,malogranatum et palma et malumet omnia ligna agri aruerunt,quia evanuit gaudiuma filiis hominum.
JOEL|1|13|Accingite vos et plangite, sacerdotes;ululate, ministri altaris.Ingredimini, cubate in sacco,ministri Dei mei,quoniam interiit de domo Dei vestrioblatio et libatio.
JOEL|1|14|Sanctificate ieiunium,vocate coetum,congregate senes,omnes habitatores terraein domum Dei vestri,et clamate ad Dominum:
JOEL|1|15|" Heu diei!Quia prope est dies Domini,et quasi vastitas a potente veniet.
JOEL|1|16|Numquid non coram oculis vestrisalimenta perierunt,de domo Dei nostrilaetitia et exsultatio?".
JOEL|1|17|Computruerunt seminasubtus glebas suas,demolita sunt horrea,dissipatae sunt apothecae,eo quod exaruit triticum.
JOEL|1|18|Quid ingemuit animal,perterrita sunt armenta boum,quia non est pascua eis?Sed et greges pecorum disperierunt.
JOEL|1|19|Ad te, Domine, clamo,quia ignis comeditpascua deserti,et flamma succenditomnia ligna agri.
JOEL|1|20|Sed et bestiae agrisuspirant ad te,quoniam exsiccati sunt fontes aquarum,et ignis devoravitpascua deserti.
JOEL|2|1|Canite tuba in Sion,ululate in monte sancto meo;conturbentur omnes habitatores terrae,quia venit dies Domini,quia prope est.
JOEL|2|2|Dies tenebrarum et caliginis,dies nubis et turbinis;quasi aurora expansa super montespopulus multus et fortis:similis ei non fuit a principio,et post eum non eritusque in annos generationis et generationis.
JOEL|2|3|Ante faciem eius ignis vorat,et post eum exurit flamma.Quasi hortus Eden terra coram eo,et post eum solitudo deserti;neque est quod effugiat eum.
JOEL|2|4|Quasi aspectus equorum aspectus eorum,et quasi equites sic current.
JOEL|2|5|Sicut sonitus quadrigarumsuper capita montium exsiliunt,sicut sonitus flammae ignisdevorantis stipulam,velut populus fortispraeparatus ad proelium.
JOEL|2|6|A facie eius cruciabuntur populi,omnes vultus candentes.
JOEL|2|7|Sicut fortes currunt,quasi viri bellatores ascendunt murum;unusquisque in viis suis graditur,et non declinant a semitis suis.
JOEL|2|8|Unusquisque fratrem suum non coarctat,singuli in calle suo ambulant,per media tela prorumpuntsine intermissione.
JOEL|2|9|Urbem ingrediuntur,in murum discurrunt,domos conscendunt,per fenestras intrant quasi fur.
JOEL|2|10|A facie eius contremuit terra,moti sunt caeli,sol et luna obtenebrati sunt,et stellae retraxerunt splendorem suum.
JOEL|2|11|Et Dominus dedit vocem suam ante faciem exercitus sui,quia multa sunt nimis castra eius,quia fortia et facientia verbum eius;magnus enim dies Dominiet terribilis valde, et quis sustinebit eum?
JOEL|2|12|" Nunc ergo,dicit Dominus,convertimini ad me in toto corde vestro,in ieiunio et in fletu et in planctu;
JOEL|2|13|et scindite corda vestra et non vestimenta vestra,et convertimini ad Dominum Deum vestrum,quia benignus et misericors est,patiens et multae misericordiaeet placabilis super malitia ".
JOEL|2|14|Quis scit, si convertatur et ignoscatet relinquat post se benedictionem,oblationem et libationemDomino Deo vestro?
JOEL|2|15|Canite tuba in Sion,sanctificate ieiunium, vocate coetum;congregate populum, sanctificate conventum,coadunate senes,
JOEL|2|16|congregate parvulos et sugentes ubera,egrediatur sponsus de cubili suo,et sponsa de thalamo suo.
JOEL|2|17|Inter vestibulum et altare plorentsacerdotes ministri Dominiet dicant: "Parce, Domine, populo tuoet ne des hereditatem tuam in opprobrium,ut dominentur eis nationes ".Quare dicent in populis: Ubi est Deus eorum "?
JOEL|2|18|Zelatus est Dominus terram suamet pepercit populo suo.
JOEL|2|19|Et respondit Dominus et dixit populo suo: Ecce ego mittam vobisfrumentum et vinum et oleum,et replebimini eis;et non dabo vos ultraopprobrium in gentibus.
JOEL|2|20|Et eum, qui ab aquilone est,procul faciam a vobiset expellam eum in terraminviam et desertam:facies eius contra mare orientale,et extremum eius ad mare occidentale;et ascendet foetor eius,et ascendet putredo eius,quia magna operatus est.
JOEL|2|21|Noli timere, terra;exsulta et laetare,quoniam magna Dominus operatus est.
JOEL|2|22|Nolite timere, animalia regionis,quia germinaverunt pascua deserti,quia lignum attulit fructum suum,ficus et vinea dederunt divitias suas.
JOEL|2|23|Et, filii Sion, exsultateet laetamini in Domino Deo vestro,quia dedit vobispluviam iustitiaeet descendere fecit ad vosimbrem matutinum et serotinum sicut prius.
JOEL|2|24|Et implebuntur areae frumento,et redundabunt torculariavino et oleo;
JOEL|2|25|et reddam vobis annos,quos comedit locusta, bruchuset gryllus et eruca,exercitus meus magnus,quem misi in vos.
JOEL|2|26|Et comedetis vescentes et saturabiminiet laudabitis nomen Domini Dei vestri,qui mirabilia fecit vobiscum;et non confundetur populus meus in sempiternum.
JOEL|2|27|Et scietis quia in medio Israel ego sum,et ego Dominus Deus vester,et non est amplius;et non confundetur populus meus in aeternum ".
JOEL|3|1|Et erit post haec:effundam spiritum meum super omnem carnem,et prophetabunt filii vestri et filiae vestrae,senes vestri somnia somniabunt,et iuvenes vestri visiones videbunt;
JOEL|3|2|sed et super servos meos et ancillasin diebus illis effundam spiritum meum.
JOEL|3|3|Et dabo prodigia in caelo et in terra,sanguinem et ignem et columnas fumi;
JOEL|3|4|sol convertetur in tenebras,et luna in sanguinem,antequam veniat dies Dominimagnus et horribilis.
JOEL|3|5|Et erit:omnis, qui invocaverit nomen Domini, salvus erit,quia in monte Sion et in Ierusalemerit salvatio, sicut dixit Dominus,et in residuis, quos Dominus vocaverit.
JOEL|4|1|Quia ecce in diebus illiset in tempore illo,cum convertero sortemIudae et Ierusalem,
JOEL|4|2|congregabo omnes genteset deducam eas in vallem Iosaphatet disceptabo cum eis ibisuper populo meo et hereditate mea Israel,quos disperserunt in nationibus,et terram meam diviserunt.
JOEL|4|3|Et super populum meum miserunt sortem;et dederunt puerum pro meretriceet puellam vendiderunt pro vino, ut biberent.
JOEL|4|4|Verum quid vobis et mihi, Tyrus et Sidon et omnes termini Philisthaeae? Numquid ultionem vos reddetis mihi? Et si ulciscimini vos contra me, cito velociter reddam ultionem vestram super caput vestrum.
JOEL|4|5|Argentum enim meum et aurum tulistis et pretiosa bona mea intulistis in delubra vestra.
JOEL|4|6|Et filios Iudae et filios Ierusalem vendidistis filiis Graecorum, ut longe faceretis eos de finibus suis.
JOEL|4|7|Ecce ego suscitabo eos de loco, in quo vendidistis eos, et reddam ultionem vestram in caput vestrum.
JOEL|4|8|Et vendam filios vestros et filias vestras in manibus filiorum Iudae; et venumdabunt eos Sabaeis, genti longinquae, quia Dominus locutus est.
JOEL|4|9|Clamate hoc in gentibus,sanctificate bellum,suscitate robustos;accedant, ascendantomnes viri bellatores.
JOEL|4|10|Concidite vomeres vestros in gladioset falces vestras in lanceas;infirmus dicat: Fortis ego sum ".
JOEL|4|11|Erumpite et venite,omnes gentes de circuitu,et congregamini ibi!Deduc, Domine, robustos tuos!
JOEL|4|12|Consurgant et ascendant gentesin vallem Iosaphat,quia ibi sedebo, ut iudicemomnes gentes in circuitu.
JOEL|4|13|Mittite falces,quoniam maturavit messis;venite et premite,quia plenum est torcular:exuberant torcularia,quia magna est malitia eorum.
JOEL|4|14|Populi, populiin valle Decisionis,quia iuxta est dies Dominiin valle Decisionis.
JOEL|4|15|Sol et luna obtenebrati sunt,et stellae retraxerunt splendorem suum.
JOEL|4|16|Et Dominus de Sion rugietet de Ierusalem dabit vocem suam;et movebuntur caeli et terra,et Dominus refugium populo suoet fortitudo filiis Israel.
JOEL|4|17|Et scietis quia ego Dominus Deus vesterhabitans in Sion monte sancto meo;et erit Ierusalem locus sanctus,et alieni non transibunt per eam amplius.
JOEL|4|18|Et erit in die illa:stillabunt montes mustum,et colles fluent lacte;et per omnes rivos Iudae ibunt aquae,et fons de domo Domini egredieturet irrigabit torrentem Settim.
JOEL|4|19|Aegyptus in desolationem erit,et Idumaea in desertum desolationis,pro eo quod inique egerint in filios Iudaeet effuderint sanguinem innocentem in terra eorum.
JOEL|4|20|Et Iuda in aeternum habitabitur,et Ierusalem in generationem et generationem;
JOEL|4|21|et vindicabo sanguinem eorum, quem non relinquam impunitum;et Dominus commoratur in Sion.
AMOS|1|1|Verba Amos, qui fuit in pastori bus de Thecua; quae vidit super Israel in diebus Oziae regis Iudae et in diebus Ieroboam filii Ioas regis Israel, duobus annis ante terraemotum.
AMOS|1|2|Et dixit: Dominus de Sion rugitet de Ierusalem dat vocem suam;et lugent pascua pastorum,et exsiccatur vertex Carmeli ".
AMOS|1|3|Haec dicit Dominus: Super tribus sceleribus Damasciet super quattuor verbum non revocabo:eo quod trituraverint in plaustris ferreis Galaad,
AMOS|1|4|mittam ignem in domum Hazael,et devorabit aedes Benadad;
AMOS|1|5|conteram vectem Damasciet disperdam habitatorem de Biceatavenet tenentem sceptrum de Betheden;et transferetur populus Syriae Cir ",dicit Dominus.
AMOS|1|6|Haec dicit Dominus: Super tribus sceleribus Gazaeet super quattuor verbum non revocabo:eo quod transtulerint captivitatem perfectam,ut traderent eam in Edom,
AMOS|1|7|mittam ignem in murum Gazae,et devorabit aedes eius;
AMOS|1|8|disperdam habitatorem de Azotoet tenentem sceptrum de Ascalone;convertam manum meam super Accaron,et peribunt reliqui Philisthinorum ",dicit Dominus Deus.
AMOS|1|9|Haec dicit Dominus: Super tribus sceleribus Tyriet super quattuor verbum non revocabo:eo quod tradiderint captivitatem perfectam in Edomet non sint recordati foederis fratrum,
AMOS|1|10|mittam ignem in murum Tyri,et devorabit aedes eius ".
AMOS|1|11|Haec dicit Dominus: Super tribus sceleribus Edomet super quattuor verbum non revocabo:eo quod persecutus sit in gladio fratrem suumet violaverit misericordiam eiuset tenuerit ultra furorem suumet indignationem suam servaverit usque in finem,
AMOS|1|12|mittam ignem in Theman,et devorabit aedes Bosrae ".
AMOS|1|13|Haec dicit Dominus: Super tribus sceleribus filiorum Ammonet super quattuor verbum non revocabo:eo quod dissecuerint praegnantes Galaadad dilatandum terminum suum,
AMOS|1|14|succendam ignem in muro Rabba,et devorabit aedes eius in ululatu in die belliet in turbine in die procellae;
AMOS|1|15|et ibit rex eorum in captivitatem,ipse et principes eius simul ",dicit Dominus.
AMOS|2|1|Haec dicit Dominus: Super tribus sceleribus Moabet super quattuor verbum non revocabo:eo quod incenderit ossa regis Edomusque ad cinerem,
AMOS|2|2|mittam ignem in Moab,et devorabit aedes Carioth,et morietur in tumultu Moab,in clamore et voce tubae;
AMOS|2|3|disperdam iudicem de medio eiuset omnes principes eius interficiam cum eo ",dicit Dominus.
AMOS|2|4|Haec dicit Dominus: Super tribus sceleribus Iudaeet super quattuor verbum non revocabo:eo quod abiecerint legem Dominiet mandata eius non custodierintC deceperunt enim eos idola sua,post quae abierant patres eorum C
AMOS|2|5|mittam ignem in Iudam,et devorabit aedes Ierusalem ".
AMOS|2|6|Haec dicit Dominus: Super tribus sceleribus Israelet super quattuor verbum non revocabo:eo quod vendiderint pro argento iustumet pauperem pro calceamentis;
AMOS|2|7|qui contriverint super pulverem terrae capita pauperumet viam humilium declinaverint,et filius ac pater eius iverint ad puellam,ut violarent nomen sanctum meum;
AMOS|2|8|et super vestimentis pignoratis accubuerintiuxta omne altareet vinum damnatorum biberintin domo Dei sui.
AMOS|2|9|Ego autem exterminaveramAmorraeum a facie eorum,cuius altitudo sicut altitudo cedrorum,et fortitudo quasi quercuum;exterminaveram fructum eius desuperet radices eius subter.
AMOS|2|10|Ego ascendere vos fecide terra Aegyptiet duxi vos in desertoquadraginta annis,ut possideretis terram Amorraei;
AMOS|2|11|et suscitavi de filiis vestris prophetas et de iuvenibus vestris nazaraeos.Numquid non ita est, filii Israel?,dicit Dominus.
AMOS|2|12|Et propinastis nazaraeis vinumet prophetis mandastis dicentes:Ne prophetetis".
AMOS|2|13|Ecce ego comprimam vos ad solum,sicut comprimit plaustrumonustum feno;
AMOS|2|14|deerit fuga a veloce,et fortis non firmabit virtutem suam,et robustus non salvabit animam suam;
AMOS|2|15|tenens arcum non stabit,et velox pedibus suis non salvabitur;ascensor equi non salvabit animam suam,
AMOS|2|16|et fortissimus corde inter robustosnudus fugiet in illa die ",dicit Dominus.
AMOS|3|1|Audite verbum hoc, quod locutus est Dominus super vos, filii Israel, super omnem cognationem, quam eduxi de terra Aegypti, dicens:
AMOS|3|2|" Tantummodo vos cognoviex omnibus cognationibus terrae;idcirco visitabo super vosomnes iniquitates vestras.
AMOS|3|3|Numquid ambulabunt duo pariter, nisi convenerint?
AMOS|3|4|Numquid rugiet leo in saltu,nisi habuerit praedam?Numquid dabit catulus leonis vocem de cubili suo,nisi aliquid apprehenderit?
AMOS|3|5|Numquid cadet avis super terramabsque laqueo?Numquid laxatur laqueus de terra, antequam quid ceperit?
AMOS|3|6|Si clanget tuba in civitate,populus non expavescet?Si erit malum in civitate,nonne Dominus fecit?
AMOS|3|7|Nihil enim faciet Dominus Deus,nisi revelaverit secretum suumad servos suos prophetas.
AMOS|3|8|Leo rugit,quis non timebit?Dominus Deus locutus est,quis non prophetabit?
AMOS|3|9|Auditum facite in aedibus Assyriaeet in aedibus terrae Aegyptiet dicite: "Congregamini super montes Samariae";et videte insanias multas in medio eiuset oppressos in sinu eius.
AMOS|3|10|Et nescierunt facere rectum,dicit Dominus,thesaurizantes violentiam et rapinasin aedibus suis ".
AMOS|3|11|Propterea haec dicit Dominus Deus: Inimicus circumdabit terram,et detrahetur ex te fortitudo tua,et diripientur aedes tuae ".
AMOS|3|12|Haec dicit Dominus: Quomodo si eruat pastor de ore leonisduo crura aut extremum auriculae, sic eruentur filii Israel,qui habitant in Samaria,in margine lectuliet in Damasci grabato.
AMOS|3|13|Audite et contestamini in domo Iacob,dicit Dominus, Deus exercituum:
AMOS|3|14|In die cum visitavero praevaricationes Israel,super eum visitabo et super altaria Bethel,et amputabuntur cornua altariset cadent in terram;
AMOS|3|15|et percutiam domum hiemalemcum domo aestiva,et peribunt domus eburneae,et dissipabuntur aedes magnae ",dicit Dominus.
AMOS|4|1|Audite verbum hoc,vaccae Basan,quae estis in monte Samariae,quae opprimitis egenoset vexatis pauperes,quae dicitis dominis vestris: Affer, ut bibamus ".
AMOS|4|2|Iuravit Dominus Deusin sanctitate sua: Ecce dies venient super vos,et levabunt vos in contiset posteros vestros in hamis piscatoriis;
AMOS|4|3|et per aperturas exibitis altera contra alteramet proiciemini in Armon ",dicit Dominus.
AMOS|4|4|" Venite in Bethel et impie agite,ad Galgalam et multiplicate praevaricationem;et offerte mane victimas vestras,tribus diebus decimas vestras,
AMOS|4|5|et sacrificate de fermentato laudemet vocate voluntarias oblationes et annuntiate;sic enim diligitis, filii Israel ",dicit Dominus Deus.
AMOS|4|6|" Unde et ego dedi vobisvacuitatem dentium in cunctis urbibus vestriset indigentiam panis in omnibus locis vestris;et non estis reversi ad me ",dicit Dominus.
AMOS|4|7|" Ego quoque prohibui a vobis imbrem,cum adhuc tres menses superessent usque ad messem;et plui super unam civitatemet super alteram civitatem non plui: pars una compluta est,et pars, super quam non plui, aruit.
AMOS|4|8|Tunc fugiebant duae, tres civitatesad unam civitatem, ut biberent aquam,et non satiabantur;sed non redistis ad me ",dicit Dominus.
AMOS|4|9|" Percussi vos in vento urente et in aurugine;multitudinem hortorum vestrorum et vinearum vestrarum,ficeta vestra et oliveta vestracomedit eruca;sed non redistis ad me ",dicit Dominus.
AMOS|4|10|" Misi in vos pestemsicut pestem Aegypti,percussi in gladio iuvenes vestros,captis equis vestris;et ascendere feci putredinemcastrorum vestrorum in nares vestras;sed non redistis ad me ",dicit Dominus.
AMOS|4|11|" Subverti vos,sicut subvertit Deus Sodomam et Gomorram,et facti estis quasi torrisraptus ab incendio;sed non redistis ad me ",dicit Dominus.
AMOS|4|12|Quapropter haec faciam tibi, Israel,et quia haec faciam tibi,praeparare in occursum Dei tui, Israel;
AMOS|4|13|quia ecce formans montes et creans ventumet annuntians homini cogitationem eius,faciens auroram et tenebraset gradiens super excelsa terrae;Dominus, Deus exercituum, nomen eius.
AMOS|5|1|Audite verbum istud,quod ego levo super vos,planctum, domus Israel:
AMOS|5|2|Cecidit, non adiciet ut resurgatvirgo Israel;proiecta est in terram suam,non est qui suscitet eam.
AMOS|5|3|Quia haec dicit Dominus Deus: Urbs, de qua egrediebantur mille,relinquentur in ea centum;et de qua egrediebantur centum,relinquentur in ea decempro domo Israel ".
AMOS|5|4|Quia haec dicit Dominus domui Israel: Quaerite me et vivetis;
AMOS|5|5|et nolite quaerere Bethelet in Galgalam nolite intrareet in Bersabee nolite transire,quia Galgala captiva ducetur,et Bethel erit iniquitas ".
AMOS|5|6|Quaerite Dominum et vivite;ne forte invadat sicut ignisdomum Ioseph,et devoret, et non sitqui exstinguat Bethel.
AMOS|5|7|Qui convertunt in absinthium iudiciumet iustitiam in terram deiciunt.
AMOS|5|8|Qui facit stellas Pliadis et Orionemet convertit in mane tenebraset diem in noctem obscurat;qui vocat aquas mariset effundit eas super faciem terrae;Dominus nomen eius.
AMOS|5|9|Qui micare facit vastitatem super robustumet vastitatem super arcem affert.
AMOS|5|10|Odio habuerunt corripientem in portaet loquentem perfecte abominati sunt.
AMOS|5|11|Idcirco, pro eo quod conculcastis pauperemet portionem frumenti abstulistis ab eo,domos quadro lapide aedificastiset non habitabitis in eis,vineas plantastis amantissimaset non bibetis vinum earum.
AMOS|5|12|Quia cognovi multa scelera vestraet fortia peccata vestra,opprimentes iustum, accipientes munuset pauperes deprimentes in porta.
AMOS|5|13|Ideo prudens in tempore illo tacet,quia tempus malum est.
AMOS|5|14|Quaerite bonum et non malum,ut vivatis,ita ut sit Dominus, Deus exercituum,vobiscum, sicut dixistis.
AMOS|5|15|Odite malum et diligite bonumet constituite in porta iudicium,si forte misereatur Dominus, Deus exercituum,reliquiis Ioseph.
AMOS|5|16|Propterea haec dicit Dominus,Deus exercituum, dominator: In omnibus plateis planctus,et in cunctis viis dicetur: "Vae, vae!";et vocabunt agricolam ad luctumet ad planctum eos, qui sciunt lamentationem.
AMOS|5|17|Et in omnibus vineis erit luctus,quia pertransibo in medio tui ",dicit Dominus.
AMOS|5|18|Vae desiderantibus diem Domini!Ad quid vobis dies Domini?Tenebrae et non lux.
AMOS|5|19|Quomodo si fugiat vir a facie leonis,et occurrat ei ursus;et ingrediatur domumet innitatur manu sua super parietem,et mordeat eum coluber.
AMOS|5|20|Numquid non tenebrae dies Domini et non lux?Et caligo sine splendore in ea?
AMOS|5|21|" Odi, proieci festivitates vestraset non delector coetibus vestris.
AMOS|5|22|Quod si obtuleritis mihi holocautomata,oblationes vestras non suscipiamet sacrificia pinguium vestrorum non respiciam.
AMOS|5|23|Aufer a me tumultum carminum tuorum,et canticum lyrarum tuarum non audiam.
AMOS|5|24|Et affluat quasi aqua iudicium,et iustitia quasi torrens perennis.
AMOS|5|25|Numquid hostias et oblationes obtulistis mihi in desertoquadraginta annis, domus Israel?
AMOS|5|26|Et portastis Saccut regem vestrum,et Caivan, imagines vestras,sidus deorum vestrorum, quae fecistis vobis.
AMOS|5|27|Et migrare vos faciam trans Damascum ",dicit Dominus; Deus exercituum nomen eius.
AMOS|6|1|Vae, qui tranquilli sunt in Sionet confidunt in monte Samariae;designati primitiae populorum,ad quos venit domus Israel!
AMOS|6|2|Transite in Chalanne et videte;et ite inde in Emath magnamet descendite in Geth Palaestinorum.Numquid meliores regnis istis vos,aut latior terminus eorum termino vestro est?
AMOS|6|3|Qui removetis diem malumet appropinquare facitis solium violentiae.
AMOS|6|4|Qui dormiunt in lectis eburneis,recumbentes in stratis suis,comedentes agnos de gregeet vitulos de medio armenti;
AMOS|6|5|canentes ad vocem psalterii,sicut David excogitant sibi vasa cantici;
AMOS|6|6|bibentes vinum in phialis,optimis unguentis delibuti,et non sunt contristati super ruina Ioseph.
AMOS|6|7|Quapropter nunc migrabunt in capite transmigrantium,et auferetur factio lascivientium.
AMOS|6|8|Iuravit Dominus Deus in anima sua,dicit Dominus, Deus exercituum: Detestor ego superbiam Iacobet domos eius odiet tradam civitatem et plenitudinem eius ".
AMOS|6|9|Quod si reliqui fuerintdecem viri in domo una,et ipsi morientur;
AMOS|6|10|et tollet eum propinquus suuset comburet eum, ut efferat ossa de domo,et dicet ei, qui in penetralibus domus est: Numquid adhuc est penes te? ".Et respondebit: "Non est";et dicet ei: "Tace!";non est qui recordetur nominis Domini.
AMOS|6|11|Quia ecce Dominus mandatet percutiet domum maiorem ruiniset domum minorem scissionibus.
AMOS|6|12|Numquid currunt in petris equi,aut aratur mare in bobus,quoniam convertistis in venenum iudiciumet fructum iustitiae in absinthium?
AMOS|6|13|Qui laetantur pro Lodabar,qui dicunt: " Numquid non in fortitudine nostracepimus nobis Carnaim? ".
AMOS|6|14|" Ecce enim suscitabo super vos, domus Israel,dicit Dominus, Deus exercituum, gentem;et oppriment vos ab introitu Emathusque ad torrentem Arabae ".
AMOS|7|1|Haec ostendit mihi Dominus Deus: et ecce, ipse formabat lo custas in principio, cum germinarent serotinae fruges; et ecce fruges serotinae post fruges demessas regis.
AMOS|7|2|Et factum est, cum consummasset comedere herbam terrae, dixi: "Domine Deus, propitius esto, obsecro; quomodo stabit Iacob, quia parvulus est? ".
AMOS|7|3|Misertus est Dominus super hoc. " Non erit ", dixit Dominus Deus.
AMOS|7|4|Haec ostendit mihi Dominus Deus: et ecce, vocabat ad iudicium per ignem Dominus Deus, et devoravit abyssum magnam et comedit simul partem.
AMOS|7|5|Et dixi: " Domine Deus, quiesce, obsecro; quomodo stabit Iacob, quia parvulus est? ".
AMOS|7|6|Misertus est Dominus super hoc. " Sed et istud non erit ", dicit Dominus Deus.
AMOS|7|7|Haec ostendit mihi Dominus Deus: ecce vir stans super murum litum, et in manu eius trulla caementarii.
AMOS|7|8|Et dixit Dominus ad me: " Quid tu vides, Amos? ". Et dixi: " Trullam caementarii ". Et dixit Dominus: "Ecce ego ponam trullam in medio populi mei Israel; non adiciam ultra ignoscere ei.
AMOS|7|9|Et demolientur excelsa Isaac, et sanctuaria Israel desolabuntur, et consurgam super domum Ieroboam in gladio ".
AMOS|7|10|Et misit Amasias sacerdos Bethel ad Ieroboam regem Israel dicens: " Conspiravit contra te Amos in medio domus Israel; non poterit terra sustinere universos sermones eius.
AMOS|7|11|Haec enim dicit Amos: "In gladio morietur Ieroboam, et Israel captivus migrabit de terra sua" ".
AMOS|7|12|Et dixit Amasias ad Amos: " Qui vides, gradere. Fuge in terram Iudae et comede ibi panem et prophetabis ibi;
AMOS|7|13|et in Bethel non adicies ultra ut prophetes, quia sanctuarium regis est, et domus regni est ".
AMOS|7|14|Responditque Amos et dixit ad Amasiam: Non sum prophetaet non sum filius prophetae;sed armentarius ego sum, vellicans sycomoros.
AMOS|7|15|Et tulit me Dominus,cum sequerer gregem,et dixit Dominus ad me:Vade, propheta ad populum meum Israel".
AMOS|7|16|Et nunc audi verbum Domini. Tu dicis: "Non prophetabis super Israel et non stillabis verba super domum Isaac".
AMOS|7|17|Propter hoc haec dicit Dominus: "Uxor tua in civitate fornicabitur, et filii tui et filiae tuae in gladio cadent, et humus tua funiculo metietur; et tu in terra polluta morieris, et Israel captivus migrabit de terra sua".
AMOS|8|1|Haec ostendit mihi Dominus Deus:et ecce canistrum pomorum.
AMOS|8|2|Et dixit: " Quid tu vides, Amos? ".Et dixi: " Canistrum pomorum ".Et dixit Dominus ad me: Venit finis super populum meum Israel;non adiciam ultra ignoscere ei.
AMOS|8|3|Et lugent cantatrices palatii in die illa,dicit Dominus Deus;multa erunt cadavera,in omni loco proicientur: silentium.
AMOS|8|4|Audite hoc, qui conteritis pauperemet deficere facitis egenos terrae,
AMOS|8|5|dicentes: "Quando transibit neomenia,et venumdabimus merces?Et sabbatum, et aperiemus frumentum,ut imminuamus mensuram et augeamus siclumet supponamus stateras dolosas,
AMOS|8|6|ut possideamus in argento egenoset pauperem pro calceamentiset quisquilias frumenti vendamus?"".
AMOS|8|7|Iuravit Dominus in superbia Iacob: Non obliviscar in perpetuum omnia opera eorum.
AMOS|8|8|Numquid super isto non commovebitur terra,et lugebit omnis habitator eius,et ascendet quasi fluvius universa,fervebit et decrescet quasi flumen Aegypti?
AMOS|8|9|Et erit: in die illa,dicit Dominus Deus,occidere faciam solem in meridieet tenebrescere faciam terram in die luminis
AMOS|8|10|et convertam festivitates vestras in luctumet omnia cantica vestra in planctum;et inducam super omnes lumbos saccumet super omne caput calvitium;et ponam eam quasi luctum unigenitiet novissima eius quasi diem amarum.
AMOS|8|11|Ecce dies veniunt,dicit Dominus,et mittam famem in terram;non famem panis neque sitim aquae,sed audiendi verbum Domini ".
AMOS|8|12|Et fugient a mari usque ad mare;et ab aquilone usque ad orientem circuibunt,quaerentes verbum Domini,et non invenient.
AMOS|8|13|In die illa deficient virgines pulchraeet adulescentes in siti.
AMOS|8|14|Qui iurant in delicto Samariaeet dicunt: " Vivit Deus tuus, Dan! "et " Vivit via, Bersabee! ",et cadent et non resurgent ultra.
AMOS|9|1|Vidi Dominumstantem super altare,et dixit: "Percute capitellum,et commoveantur superliminaria;frange eos in capite omnes,et novissimum eorum in gladio interficiam;non fugiet ex eis fugitivus,et non salvabitur superstes eis.
AMOS|9|2|Si descenderint usque ad infernum,inde manus mea educet eos;et si ascenderint usque in caelum,inde detraham eos.
AMOS|9|3|Et si absconditi fuerint in vertice Carmeli,inde quaeram et auferam eos;et si celaverint se ab oculis meisin profundo maris,ibi mandabo serpenti, et mordebit eos;
AMOS|9|4|et si abierint in captivitatemcoram inimicis suis,ibi mandabo gladio, et occidet eos,et ponam oculos meos super eosin malum et non in bonum ".
AMOS|9|5|Et Dominus, Deus exercituum,qui tangit terram, et tabescet.Et lugebunt omnes habitantes in ea;et ascendet sicut fluvius ea omniset decrescet sicut flumen Aegypti.
AMOS|9|6|Qui aedificat in caelo ascensus suoset cameram suam super terram fundat,qui vocat aquas mariset effundit eas super faciem terrae;Dominus nomen eius.
AMOS|9|7|" Numquid non ut filii Aethiopumvos estis mihi, filii Israel?,ait Dominus.Numquid non Israel ascendere fecide terra Aegyptiet Philisthim de Caphtoret Syros de Cir?
AMOS|9|8|Ecce oculi Domini Deisuper regnum peccans,et conteram illuda facie terrae;verumtamen conterens non conteramdomum Iacob,dicit Dominus.
AMOS|9|9|Ecce enim mandabo egoet concutiam in omnibus gentibus domum Israel,sicut concutitur triticum in cribro,et non cadet lapillus super terram.
AMOS|9|10|In gladio morientur omnes peccatores populi mei,qui dicunt: "Non appropinquabit et non venietsuper nos malum".
AMOS|9|11|In die illa suscitabotabernaculum David, quod cecidit,et reaedificabo rupturas eius;et ea, quae corruerant, instauraboet reaedificabo illud sicut diebus antiquis,
AMOS|9|12|ut possideantreliquias Edomet omnes nationes,super quas invocatum est nomen meum,dicit Dominus, qui faciet haec.
AMOS|9|13|Ecce dies veniunt,dicit Dominus,et comprehendet arator messorem,et calcator uvae mittentem semen; et stillabunt montes mustum,et omnes colles liquefient.
AMOS|9|14|Et convertam captivitatem populi mei Israel;et aedificabunt civitates vastatas et inhabitabuntet plantabunt vineas et bibent vinum earumet facient hortos et comedent fructus eorum.
AMOS|9|15|Et plantabo eos super humum suam,et non evellentur ultrade terra sua, quam dedi eis ",dicit Dominus Deus tuus.
OBAD|1|1|Visio Abdiae.Haec dicit Dominus Deus ad Edom.Auditum audivimus a Domino,et legatus ad gentes missus est: Surgite, et consurgamusadversus eum in proelium! ".
OBAD|1|2|" Ecce parvulum te dabo in gentibus,contemptibilis tu es valde.
OBAD|1|3|Superbia cordis tui decepit tehabitantem in scissuris petrae,exaltantem solium suum;qui dicit in corde suo:Quis detrahet me in terram?".
OBAD|1|4|Si exaltatus fueris ut aquilaet si inter sidera posueris nidum tuum,inde detraham te ",dicit Dominus.
OBAD|1|5|Si fures introissent ad te,si latrones per noctem,quomodo periisses!Nonne furati essent sufficientia sibi?Si vindemiatores introissent ad te,nonne racemos tantum reliquissent?
OBAD|1|6|Quomodo scrutati sunt Esau?Investigaverunt abscondita eius.
OBAD|1|7|Usque ad terminum eiecerunt te,omnes viri foederis tui deceperunt te,invaluerunt adversum te viri pacis tuae;qui comedunt tecum, ponent insidias subter te.Non est prudentia in eo.
OBAD|1|8|" Numquid non in die illa,dicit Dominus,perdam sapientes de Edomet prudentiam de monte Esau?
OBAD|1|9|Et timebunt fortes tui Theman,ut intereat omnis vir de monte Esau.
OBAD|1|10|Propter interfectionemet propter iniquitatemin fratrem tuum Iacoboperiet te confusio,et peribis in aeternum.
OBAD|1|11|In die cum stares ex adverso,quando capiebant alieni exercitum eius,et extranei ingrediebantur portas eiuset super Ierusalem mittebant sortem,tu quoque eras quasi unus ex eis ".
OBAD|1|12|Et non respicies diem fratris tui,diem calamitatis eius;et non laetaberis super filios Iudaein die perditionis eorum;et non magnificabis os tuumin die angustiae.
OBAD|1|13|Neque ingredieris portam populi meiin die ruinae eorum;neque respicies et tu malum eiusin die vastitatis illiuset non mittes manum in opes eiusin die vastitatis illius;
OBAD|1|14|neque stabis in exitibus,ut interficias eos, qui fugerint,et non trades reliquos eiusin die tribulationis.
OBAD|1|15|Quoniam iuxta est dies Dominisuper omnes gentes:sicut fecisti, fiet tibi,retributio tua convertetur in caput tuum.
OBAD|1|16|Quomodo enim bibistis super montem sanctum meum,bibent omnes gentes iugiter;et bibent et absorbebuntet erunt quasi non fuerint.
OBAD|1|17|Et in monte Sion erit salvatio,et erit sanctum;et possidebit domus Iacobeos, qui se possederant.
OBAD|1|18|Et erit domus Iacob ignis,et domus Ioseph flamma,et domus Esau stipula;et succendentur in eis, et devorabunt eos,et non erunt reliquiae domus Esau,quia Dominus locutus est.
OBAD|1|19|Et hereditabunt austrum,montem Esau,et Sephelam Philisthim;et possidebunt regionem Ephraimet regionem Samariae,et Beniamin possidebit Galaad;
OBAD|1|20|et transmigratio prima filiorum Israelpossidebit terram Chananaeorum usque ad Sareptam;et transmigratio Ierusalem, quae in Sapharad est,possidebit civitates austri.
OBAD|1|21|Et ascendent salvatores in montem Sioniudicare montem Esau,et erit Domino regnum.
JONAH|1|1|Et factum est verbum Domini ad Ionam filium Amathi dicens:
JONAH|1|2|" Surge et vade in Nineven civitatem grandem et praedica in ea, quia ascendit malitia eius coram me ".
JONAH|1|3|Et surrexit Ionas, ut fugeret in Tharsis a facie Domini; et descendit Ioppen et invenit navem euntem in Tharsis et dedit naulum eius et descendit in eam, ut iret cum eis in Tharsis a facie Domini.
JONAH|1|4|Dominus autem misit ventum magnum in mare, et facta est tempestas magna in mari, et navis periclitabatur conteri.
JONAH|1|5|Et timuerunt nautae et clamaverunt unusquisque ad deum suum et miserunt vasa, quae erant in navi, in mare, ut alleviaretur ab eis. Ionas autem descenderat ad interiora navis et, cum recubuisset, dormiebat sopore gravi.
JONAH|1|6|Et accessit ad eum gubernator et dixit ei: " Quid? Tu sopore deprimeris? Surge, invoca Deum tuum, si forte recogitet Deus de nobis, et non pereamus.
JONAH|1|7|Et dixit unusquisque ad collegam suum: " Venite, et mittamus sortes, ut sciamus quare hoc malum sit nobis ". Et miserunt sortes, et cecidit sors super Ionam.
JONAH|1|8|Et dixerunt ad eum: " Indica nobis cuius causa malum istud sit nobis. Quod est opus tuum, et unde venis? Quae terra tua, et ex quo populo es tu?.
JONAH|1|9|Et dixit ad eos: " Hebraeus ego sum et Dominum, Deum caeli, ego timeo, qui fecit mare et aridam ".
JONAH|1|10|Et timuerunt viri timore magno et dixerunt ad eum: " Quid hoc fecisti?. Cognoverant enim viri quod a facie Domini fugeret, quia indicaverat eis.
JONAH|1|11|Et dixerunt ad eum: " Quid faciemus tibi, ut conticescat mare a nobis?. Mare enim magis ac magis intumescebat.
JONAH|1|12|Et dixit ad eos: " Tollite me et mittite in mare, et cessabit mare a vobis; scio enim ego quoniam propter me tempestas haec grandis super vos.
JONAH|1|13|Et remigabant viri, ut reverterentur ad aridam; et non valebant, quia mare magis intumescebat super eos.
JONAH|1|14|Et clamaverunt ad Dominum et dixerunt: " Quaesumus, Domine, ne pereamus in anima viri istius, et ne des super nos sanguinem innocentem; quia tu, Domine, sicut voluisti, fecisti ".
JONAH|1|15|Et tulerunt Ionam et miserunt in mare; et stetit mare a fervore suo.
JONAH|1|16|Et timuerunt viri timore magno Dominum et immolaverunt hostias Domino et voverunt vota.
JONAH|2|1|Et praeparavit Dominus piscem grandem, ut deglutiret Ionam; et erat Ionas in ventre piscis tribus diebus et tribus noctibus.
JONAH|2|2|Et oravit Ionas ad Dominum Deum suum de ventre piscis
JONAH|2|3|et dixit: " Clamavi de tribulatione mea ad Dominum,et respondit mihi;de ventre inferi clamavi,et exaudisti vocem meam.
JONAH|2|4|Et proiecisti me in profundum in corde maris,et flumen circumdedit me;omnes gurgites tui et fluctus tuisuper me transierunt.
JONAH|2|5|Et ego dixi: "Abiectus suma conspectu oculorum tuorum;verumtamen rursus videbotemplum sanctum tuum".
JONAH|2|6|Circumdederunt me aquae usque ad guttur,abyssus vallavit me,iuncus alligatus est capiti meo.
JONAH|2|7|Ad extrema montium descendi,terrae vectes concluserunt me in aeternum,sed eduxisti de fovea vitam meam,Domine Deus meus.
JONAH|2|8|Cum angustiaretur in me anima mea,Domini recordatus sum,et venit ad te oratio mea,ad templum sanctum tuum.
JONAH|2|9|Qui colunt idola vana,pietatem suam derelinquunt;
JONAH|2|10|ego autem in voce laudisimmolabo tibi,quaecumque vovi, reddam;salus Domini est ".
JONAH|2|11|Et dixit Dominus pisci, et evomuit Ionam in aridam.
JONAH|3|1|Et factum est verbum Domini ad Ionam secundo dicens:
JONAH|3|2|" Surge, vade in Nineven civitatem magnam et praedica in ea praedicationem, quam ego loquor ad te ".
JONAH|3|3|Et surrexit Ionas et abiit in Nineven iuxta verbum Domini.Et Nineve erat civitas magna coram Deo, itinere trium dierum.
JONAH|3|4|Et coepit Ionas introire in civitatem itinere diei unius; et clamavit et dixit: " Adhuc quadraginta dies, et Nineve subvertetur ".
JONAH|3|5|Et crediderunt viri Ninevitae in Deo; et praedicaverunt ieiunium et vestiti sunt saccis a maiore usque ad minorem.
JONAH|3|6|Et pervenit verbum ad regem Nineve; et surrexit de solio suo et abiecit pallium suum a se et indutus est sacco et sedit in cinere.
JONAH|3|7|Et clamavit et dixit in Nineve decreto regis et principum eius dicens: " Homines et iumenta et boves et pecora non gustent quidquam nec pascantur et aquam non bibant;
JONAH|3|8|et operiantur saccis homines et iumenta et clament ad Deum in fortitudine, et convertatur vir a via sua mala et a violentia, quae est in manibus eorum.
JONAH|3|9|Quis scit si convertatur et ignoscat Deus et revertatur a furore irae suae, et non peribimus? ".
JONAH|3|10|Et vidit Deus opera eorum, quia conversi sunt de via sua mala; et misertus est Deus super malum, quod lo cutus fuerat ut faceret eis, etnon fecit.
JONAH|4|1|Et afflictus est Ionas afflictione magna et iratus est;
JONAH|4|2|et oravit ad Dominum et dixit: " Obsecro, Domine, numquid non hoc est verbum meum, cum adhuc essem in terra mea? Propter hoc praeoccupavi ut fugerem in Tharsis. Sciebam enim quia tu Deus clemens et misericors es, longanimis et multae miserationis et ignoscens super malitia.
JONAH|4|3|Et nunc, Domine, tolle, quaeso, animam meam a me, quia melior est mihi mors quam vita".
JONAH|4|4|Et dixit Dominus: " Putasne bene irasceris tu? ".
JONAH|4|5|Et egressus est Ionas de civitate et sedit contra orientem civitatis et fecit sibimet umbraculum ibi et sedebat subter illud in umbra, donec videret quid accideret in civitate.
JONAH|4|6|Et praeparavit Dominus Deus hederam, et ascendit super Ionam, ut esset umbra super caput eius et protegeret eum ab afflictione sua. Et laetatus est Ionas super hedera laetitia magna.
JONAH|4|7|Et paravit Deus vermem, cum surgeret aurora in crastinum, et percussit hederam, quae exaruit.
JONAH|4|8|Et, cum ortus fuisset sol, praecepit Deus vento orientali calido; et percussit sol super caput Ionae, et elanguit; et petivit animae suae, ut moreretur, et dixit: " Melius est mihi mori quam vivere "
JONAH|4|9|Et dixit Deus ad Ionam: " Putasne bene irasceris tu super hedera? ". Et dixit: " Bene irascor ego usque ad mortem ".
JONAH|4|10|Et dixit Dominus: " Tu doles super hederam, in qua non laborasti neque fecisti, ut cresceret, quae sub una nocte nata est et sub una nocte periit.
JONAH|4|11|Et ego non parcam Nineve civitati magnae, in qua sunt plus quam centum viginti milia hominum, qui nesciunt quid sit inter dexteram et sinistram suam, et iumenta multa? ".
MIC|1|1|Verbum Domini, quod factum est ad Michaeam Morasthiten in diebus Ioatham, Achaz, Ezechiae regum Iudae, quod vidit super Samariam et Ierusalem.
MIC|1|2|Audite, populi omnes,et attendat terra et plenitudo eius;et sit Dominus Deus vobis in testem,Dominus de templo sancto suo.
MIC|1|3|Quia ecce Dominus egreditur de loco suoet descendet et calcabitsuper excelsa terrae;
MIC|1|4|et liquescent montes subtus eum,et valles scindentursicut cera a facie ignis,sicut aquae, quae decurrunt in praeceps.
MIC|1|5|In scelere Iacob omne istudet in peccatis domus Israel.Quod scelus Iacob?Nonne Samaria?Et quae excelsa Iudae?Nonne Ierusalem?
MIC|1|6|Et ponam Samariam in acervum lapidum,in agrum, ubi plantatur vinea;et detraham in vallem lapides eiuset fundamenta eius revelabo.
MIC|1|7|Et omnia sculptilia eius concidentur,et omnes mercedes eius comburentur igne,et omnia idola eius ponam in perditionem,quia de mercedibus meretricis congregata suntet usque ad mercedem meretricis revertentur.
MIC|1|8|Super hoc plangam et ululabo;vadam spoliatus et nudus,faciam planctum velut thoumet luctum quasi struthionum,
MIC|1|9|quia desperata est plaga eius,quia venit usque ad Iudam,tetigit portam populi meiusque ad Ierusalem.
MIC|1|10|In Geth nolite annuntiare,lacrimis ne ploretis,in Bethleaphra in pulvere volutamini.
MIC|1|11|Et transite vobis, habitatores Saphir,confusi ignominia;non sunt egressi habitatores Saanan.Planctus Betheselauferet a vobis mansionem suam.
MIC|1|12|Profecto trement de bonohabitatores Maroth,quia descendit malum a Dominoin portam Ierusalem.
MIC|1|13|Iungite quadrigae equos, habitatores Lachis;principium peccati est filiae Sion,quia in te inventa sunt scelera Israel.
MIC|1|14|Propterea dabis dimissionemsuper Moresethgeth.Domus Achzib in deceptionemregibus Israel.
MIC|1|15|Adhuc expugnatorem adducam tibi,quae habitas in Maresa;usque Odollam venietgloria Israel.
MIC|1|16|Decalvare et tonderesuper filios deliciarum tuarum;dilata calvitium tuum sicut aquila, quoniam captivi ducti sunt ex te.
MIC|2|1|Vae, qui cogitant iniquitatemet operantur malum in cubilibus suis!In luce matutina faciunt illud,quoniam est in potestate manus eorum.
MIC|2|2|Concupiscunt agros, et violenter tollunt,domos, et rapiunt.Et opprimunt virum et domum eius,hominem et hereditatem eius.
MIC|2|3|Idcirco haec dicit Dominus: Ecce ego cogitosuper familiam istam malum,unde non auferetiscolla vestra;et non ambulabitis erecti,quoniam tempus pessimum est.
MIC|2|4|In die illasumetur super vos parabola,et assumetur lamentum dicentium: "Depopulatione vastati sumus;pars populi mei commutatur,quam nemo ei restituet;infideli regiones nostrae dividuntur".
MIC|2|5|Propter hoc non erit tibimittens funiculum sortisin coetu Domini ".
MIC|2|6|" Ne vaticinemini! ". " Vaticinentur,non vaticinentur de his,non cedet confusio! ".
MIC|2|7|Numquid maledicta est domus Iacob?Numquid abbreviatus est spiritus Domini,aut tales sunt actiones eius?Nonne verba eius bona suntcum eo, qui recte graditur?
MIC|2|8|Vos autem contra populum meumut adversarium consurgitis.Desuper tunica pallium tollitis ei;qui transibant fiducialiter,fiunt quasi bello capti.
MIC|2|9|Mulieres populi mei eicitisde domo deliciarum suarum;a parvulis earum aufertisdecorem meum in perpetuum.
MIC|2|10|" Surgite et ite,quia non habetis hic requiem! ".Propter immunditiam peribitisperditione pessima.
MIC|2|11|Si esset vir vento excitatuset mendacium loqueretur: Vaticinabor tibi de vino et sicera ",hic esset vates populi istius.
MIC|2|12|Congregatione congregabo, Iacob, totum te;in unum conducam reliquias Israel,pariter ponam illum quasi gregem in ovili,quasi pecus in medio pascuae;et tumultuabuntur a multitudine hominum.
MIC|2|13|Ascendet enim pandens iter ante eos;erumpent et transibunt portam, egredientur per eam.Et transibit rex eorum coram eis,et Dominus in capite eorum.
MIC|3|1|Et dixi: Audite, principes Iacobet duces domus Israel:Numquid non vestrum est scire iudicium? ".
MIC|3|2|Sed odio habetis bonum et diligitis malum.Violenter tollitis pelles eorum desuper eoset carnem eorum desuper ossibus eorum.
MIC|3|3|Qui comedunt carnem populi meiet pellem eorum desuper excoriant; et ossa eorum confringuntet secant sicut carnem assam in lebeteet quasi carnem in medio ollae.
MIC|3|4|Tunc clamabunt ad Dominum,et non exaudiet eoset abscondet faciem suam ab eisin tempore illo,sicut pessima fecerunt opera sua.
MIC|3|5|Haec dicit Dominus super prophetas,qui seducunt populum meum,qui cum habent, quid mordeant dentibus suis,praedicant pacem;et, si quis non dederit in ore eorum quippiam,sanctificant super eum proelium.
MIC|3|6|Propterea nox vobis sine visione erit,et tenebrae vobis sine divinatione; et occumbet sol super prophetas,et obtenebrabitur super eos dies.
MIC|3|7|Et confundentur videntes,et confundentur divini,et operient labia sua omnes,quia non est responsum Dei.
MIC|3|8|Verumtamen ego repletus sumfortitudine spiritus Domini,iudicio et virtute,ut annuntiem Iacob scelus suumet Israel peccatum suum.
MIC|3|9|Audite hoc, principes domus Iacobet iudices domus Israel,qui abominamini iudiciumet omnia recta pervertitis,
MIC|3|10|qui aedificatis Sion in sanguinibuset Ierusalem in iniquitate.
MIC|3|11|Principes eius in muneribus iudicant,et sacerdotes eius in mercede docent,et prophetae eius in pecunia divinant;et super Dominum requiescunt dicentes: Numquid non Dominus in medio nostrum?Non venient super nos mala ".
MIC|3|12|Propter hoc causa vestriSion quasi ager arabitur,et Ierusalem quasi acervus lapidum erit,et mons templi in excelsa silvarum.
MIC|4|1|Et erit in novissimis diebus:Erit mons domus Dominipraeparatus in vertice montiumet sublimis super colles;et fluent ad eum populi.
MIC|4|2|Et properabunt gentes multae et dicent: Venite, ascendamus ad montem Dominiet ad domum Dei Iacob,et docebit nos de viis suis,et ibimus in semitis eius ";quia de Sion egredietur lex,et verbum Domini de Ierusalem.
MIC|4|3|Et iudicabit inter populos multoset decernet gentibus fortibus usque in longinquum;et concident gladios suos in vomereset hastas suas in falces;non sumet gens adversus gentem gladium,et non discent ultra belligerare.
MIC|4|4|Et sedebit unusquisque subtus vitem suamet subtus ficum suam,et non erit qui deterreat;quia os Domini exercituum locutum est.
MIC|4|5|Quia omnes populi ambulabuntunusquisque in nomine dei sui;nos autem ambulabimus in nomine DominiDei nostri in aeternum et ultra.
MIC|4|6|" In die illa, dicit Dominus,congregabo claudicantem,et eam, quam eieceram, colligamet quam afflixeram;
MIC|4|7|et ponam claudicantem in reliquiaset eam, quae laboraverat, in gentem robustam ".Et regnabit Dominus super eos in monte Sionex hoc nunc et usque in aeternum.
MIC|4|8|Et tu, turris gregis,collis filiae Sion,usque ad te veniet et pervenietpotestas prima,regnum filiae Ierusalem.
MIC|4|9|Nunc quare clamas clamore magno?Numquid rex non est in te,aut consiliarius tuus periit,quia comprehendit te dolor sicut parturientem?
MIC|4|10|Dole et satage,filia Sion, quasi parturiens;quia nunc egredieris de civitateet habitabis in campoet venies usque ad Babylonem;ibi liberaberis,ibi redimet te Dominusde manu inimicorum tuorum.
MIC|4|11|Nunc autem congregatae sunt super tegentes multae,quae dicunt: "Profanetur,et aspiciat in Sion oculus noster ".
MIC|4|12|Ipsi autem non cognoveruntcogitationes Dominiet non intellexerunt consilium eius,quia congregavit eos quasi manipulos in area.
MIC|4|13|Surge et tritura, filia Sion,quia cornu tuum ponam ferreumet ungulas tuas ponam aereas,et comminues populos multoset vovebis Domino rapinas eorumet divitias eorum Domino universae terrae.
MIC|4|14|Nunc incide te, filia incisionis!Obsidionem posuerunt super nos;in virga percutiuntmaxillam iudicis Israel.
MIC|5|1|Sed tu, Bethlehem Ephratha,parvulus in milibus Iudae,ex te mihi egredietur,qui sit dominator in Israel;et egressus eius a temporibus antiquis,a diebus aeternitatis.
MIC|5|2|Propter hoc dabit eosusque ad tempus, in quo parturiens pariet;et reliquiae fratrum eiusconvertentur ad filios Israel.
MIC|5|3|Et stabit et pascet in fortitudine Domini,in sublimitate nominis Domini Dei sui;et habitabunt secure, quia nunc magnus eritusque ad terminos terrae,
MIC|5|4|et erit iste pax.Assyrius cum venerit in terram nostramet quando calcaverit in domibus nostris,suscitabimus super eum septem pastoreset octo primates hominum.
MIC|5|5|Et pascent terram Assyriae in gladio et terram Nemrod in lanceis;et liberabit ab Assyrio,cum venerit in terram nostramet cum calcaverit in finibus nostris.
MIC|5|6|Et erunt reliquiae Iacobin medio populorum multorumquasi ros a Dominoet quasi imbres super herbam,quae non exspectat virumet non praestolatur filios homi num.
MIC|5|7|Et erunt reliquiae Iacob in gentibus,in medio populorum multorum,quasi leo in iumentis silvarumet quasi catulus leonis in gregibus pecorum;qui cum transierit et conculcaverit et ceperit,non est qui eruat.
MIC|5|8|Exaltabitur manus tua super hostes tuos,et omnes inimici tui interibunt.
MIC|5|9|"Et erit in die illa,dicit Dominus,auferam equos tuos de medio tuiet disperdam quadrigas tuas
MIC|5|10|et perdam civitates terrae tuaeet destruam omnes munitiones tuas.
MIC|5|11|Et auferam veneficia de manu tua,et divini non erunt in te.
MIC|5|12|Et perire faciam sculptilia tuaet lapides tuos de medio tui,et non adorabis ultraopera manuum tuarum;
MIC|5|13|et evellam palos tuos de medio tuiet conteram idola tua.
MIC|5|14|Et faciam in furoreet in indignatione ultionemin omnibus gentibus,quae non audierunt ".
MIC|6|1|Audite, quae Dominus loqui tur: Surge, contende iudicio coram montibus,et audiant colles vocem tuam ".
MIC|6|2|Audite, montes, iudicium Domini,et auscultate, fundamenta terrae;quia iudicium Domini cum populo suo,et cum Israel iudicio contendit.
MIC|6|3|" Popule meus, quid feci tibiet quid molestus fui tibi?Responde mihi.
MIC|6|4|Ego eduxi te de terra Aegyptiet de domo servientium liberavi teet misi ante faciem tuam Moysenet Aaron et Mariam.
MIC|6|5|Popule meus, memento, quaeso,quid cogitaverit Balac rex Moab,et quid responderit ei Balaam filius Beor,de Settim usque ad Galgalam,ut cognoscas iustitias Domini ".
MIC|6|6|" Quid dignum offeram Domino,dum curvo genu Deo excelso?Numquid offeram ei holocautomataet vitulos anniculos?
MIC|6|7|Numquid placebunt Domino milia arietum,multa milia torrentium olei?Numquid dabo primogenitum meum pro scelere meo,fructum ventris mei pro peccato animae meae?".
MIC|6|8|Indicatum est tibi, o homo, quid sit bonum,et quid Dominus quaerat a te:utique facere iudicium et diligere caritatemet sollicitum ambulare cum Deo tuo.
MIC|6|9|Vox Domini ad civitatem clamat et sapientia est timere nomen tuum -: Audite, tribus et coetus civitatis!
MIC|6|10|Numquid tolerabo batum iniquumet ephi minus maledictum?
MIC|6|11|Numquid iustificabo stateram impiamet saccelli pondera dolosa?
MIC|6|12|Quia divites eius repleti sunt iniquitate,et habitantes in ea loquebantur mendacium,et lingua eorum fraudulenta in ore eorum.
MIC|6|13|Ego ergo coepi percutere teperditione super peccatis tuis.
MIC|6|14|Tu comedes et non saturaberis,et sordes tuae in medio tui.Tu removebis et non salvabis;et, quos salvaveris, in gladium dabo.
MIC|6|15|Tu seminabis et non metes,tu calcabis olivam et non ungeris oleo,mustum et non bibes vinum.
MIC|6|16|Custodisti praecepta Amriet omne opus domus Achab;et ambulasti in voluntatibus eorum,ut darem te in perditionemet habitantes tuos in sibilum:et opprobrium populorum portabitis ".
MIC|7|1|Vae mihi, quia factum est mihisicut congregata messe,sicut collecta vindemia!Non est botrus ad comedendum,nec praecoqua ficus, quam desideravit anima mea.
MIC|7|2|Periit pius de terra,et rectus in hominibus non est;omnes in sanguine insidiantur,vir fratrem suum rete venatur.
MIC|7|3|Ad malum manus eorum paratae sunt;princeps postulat,et iudex est pro mercede,et magnus manifestat desiderium animae suae;vae eis, qui pervertunt illud!
MIC|7|4|Qui optimus in eis, est quasi paliurus,et, qui rectus, quasi spina de saepe; dies speculatorum tuorum, visitatio tua venit:nunc erit confusio eorum.
MIC|7|5|Nolite credere amico,nolite confidere in proximo;ab ea, quae dormit in sinu tuo,custodi claustra oris tui;
MIC|7|6|quia filius contumeliam facit patri,filia consurgit adversus matrem suam,nurus adversus socrum suam:inimici hominis domestici eius.
MIC|7|7|Ego autem ad Dominum aspiciam,exspectabo Deum salvatorem meum; audiet me Deus meus.
MIC|7|8|Ne laeteris, inimica mea, super mequia cecidi: consurgam;cum sedeo in tenebris,Dominus lux mea est.
MIC|7|9|Iram Domini porto,quoniam peccavi ei,donec iudicet causam meamet faciat iudicium meum;educet me in lucem,videbo iustitiam eius.
MIC|7|10|Et aspiciet inimica meaet operietur confusione,quae dicit ad me: Ubi est Dominus Deus tuus? ".Oculi mei videbunt in eam;nunc erit in conculcationemut lutum platearum.
MIC|7|11|Dies veniet ut aedificentur maceriae tuae;in die illa dilatabuntur fines tui.
MIC|7|12|In die illa usque ad te venienthabitantes ab Assyria usque ad Aegyptumet ab Aegypto usque ad flumenet a mari usque ad mareet a monte usque ad montem.
MIC|7|13|Terra autem erit in desolationempropter habitatores suoset propter fructum operum eorum.
MIC|7|14|Pasce populum tuum in virga tua,gregem hereditatis tuae,habitantes solos in saltu,in medio hortorum;pascantur Basan et Galaadiuxta dies antiquos.
MIC|7|15|Secundum dies egressionis tuae de terra Aegyptiostende nobis mirabilia.
MIC|7|16|Videbunt gentes et confundentursuper omni fortitudine sua,ponent manum super os,aures eorum surdae erunt;
MIC|7|17|lingent pulverem sicut serpens,velut reptilia terrae.Trementes exibunt de aedibus suis " ad Dominum Deum nostrum "formidabunt et timebunt te.
MIC|7|18|Quis Deus similis tui,qui aufers iniquitatemet transis peccatumreliquiarum hereditatis tuae?Non servat in aeternum furorem suum,quoniam volens misericordiam est.
MIC|7|19|Revertetur et miserebitur nostri,calcabit iniquitates nostraset proiciet in profundum marisomnia peccata nostra.
MIC|7|20|Dabis veritatem Iacob,misericordiam Abraham,quae iurasti patribus nostrisa diebus antiquis.
NAH|1|1|Oraculum Nineve. Liber visio nis Nahum Elcesaei.
NAH|1|2|Deus aemulator et ulciscens Dominus,ulciscens Dominus et habens furorem,ulciscens Dominus in hostes suoset servans iram inimicis suis.
NAH|1|3|Dominus patiens et magnus fortitudine,nullumque impunitum derelinquet Dominus.In tempestate et turbine via eius,et nubes pulvis pedum eius.
NAH|1|4|Increpans mare et exsiccans illudet omnia flumina ad desertum deducens.Elanguit Basan et Carmelus,et flos Libani elanguit.
NAH|1|5|Montes commoti sunt ab eo,et colles conturbati;et contremuit terra a facie eiuset orbis et omnes habitantes in eo.
NAH|1|6|Ante faciem indignationis eius quis stabit,et quis resistet in aestu furoris eius? Indignatio eius effusa est ut ignis,et petrae dissolutae sunt ab eo.
NAH|1|7|Bonus Dominus,refugium in die tribulationiset sciens sperantes in se
NAH|1|8|et in diluvio transeunte;consummationem faciet adversariorum suorum,et inimicos eius persequentur tenebrae.
NAH|1|9|Quid cogitatis contra Dominum?Consummationem ipse faciet;non consurget duplex tribulatio.
NAH|1|10|Sicut spinae condensae se invicem complectenteset sicut potatores inebriaticonsumentur quasi stipula omnino arida.
NAH|1|11|Ex te exivit cogitans contra Dominum malitiam,mente pertractans praevaricationem.
NAH|1|12|Haec dicit Dominus: Et si incolumes fuerint et numerosi,sic quoque attondentur et pertransibunt;afflixi te et non affligam te ultra.
NAH|1|13|Et nunc conteram virgam eius de dorso tuoet vincula tua disrumpam ".
NAH|1|14|Et praecipiet super te Dominus: Non seminabitur ex nomine tuo amplius.De domo dei tui disperdam sculptile et conflatile;ponam sepulcrum tuum,quia inhonoratus es ".
NAH|2|1|Ecce super montes pedes evan gelizantiset annuntiantis pacem.Celebra, Iuda, festivitates tuaset redde vota tua,quia non adiciet ultra ut pertranseat in te Belial:totus interiit.
NAH|2|2|Ascendit, qui dispergat, contra te. Custodi munitionem,contemplare viam, conforta lumbos, robora virtutem valde ".
NAH|2|3|Quia restituet Dominus magnificentiam Iacobsicut magnificentiam Israel,quia praedones praedati sunt eoset propagines eorum corruperunt.
NAH|2|4|Clipeus fortium eius ruber,viri exercitus in coccineis;ignitae laminae ferreae curruum,quando praeparat bellum,et equites agitantur.
NAH|2|5|In viis furibundae currunt quadrigae,invicem colliduntur in plateis;aspectus eorum quasi lampades,quasi fulgura discurrentia.
NAH|2|6|Recordatur fortium suorum,ruunt in itineribus suis;currunt ad murum,et praeparatur umbraculum.
NAH|2|7|Portae fluviorum apertae sunt,palatium tremit.
NAH|2|8|Et speciosa denudatur, tollitur,et ancillae eius gemunt ut columbae et percutiunt corda sua.
NAH|2|9|Et Nineve quasi piscina aquarum,cuius aquae fugiunt. State, state! ";sed non est qui revertatur.
NAH|2|10|" Diripite argentum, diripite aurum! ".Et non est finis divitiarum;thesaurus ex omnibus vasis desiderabilibus.
NAH|2|11|Dissipata et vastata et dilacerata,et cor tabescens,et dissolutio geniculorum;et tremor in cunctis renibus,et facies omnium eorum candentes.
NAH|2|12|Ubi est habitaculum leonum,et spelunca catulorum leonum,ad quam ivit leo, ut duceret illuc catulum leonis,et non erat qui exterreret?
NAH|2|13|Leo cepit sufficienter catulis suiset necavit leaenis suis;et implevit praeda speluncas suaset cubile suum rapina.
NAH|2|14|" Ecce ego ad te,dicit Dominus exercituum,et succendam usque ad fumum quadrigas tuas;et leunculos tuos comedet gladius,et exterminabo de terra praedam tuam,et non audietur ultra vox nuntiorum tuorum ".
NAH|3|1|Vae, civitas sanguinum,universa mendaciipraeda plena!Non recedet a te rapina.
NAH|3|2|Vox flagellorum et vox strepitus rotarum,equi frementes et quadrigae ferventes,equites irruentes
NAH|3|3|et gladii micantes et hastae fulguranteset multitudo interfectorum et acervi mortuorum;nec est finis cadaverum,et corruunt super corpora.
NAH|3|4|Hoc propter multitudinem fornicationum meretricisspeciosae et gratae et habentis maleficia,quae vendidit gentes fornicationibus suiset nationes maleficiis suis.
NAH|3|5|" Ecce ego ad te,dicit Dominus exercituum;et levabo vestimentum tuum in faciem tuamet ostendam gentibus nuditatem tuamet regnis ignominiam tuam.
NAH|3|6|Et proiciam super te abominationeset contumeliis te afficiam;et ponam te in exemplum.
NAH|3|7|Et erit: omnis, qui viderit te,resiliet a te et dicet:Vastata est Nineve!Quis dolebit super eam?Unde quaeram consolatorem tibi?".
NAH|3|8|Numquid melior es quam Noamon,quae habitabat in fluminibus?Aquae in circuitu eius:cuius vallum mare,aquae muri eius.
NAH|3|9|Chus fuit fortitudo eiuset Aegyptus, cuius non est finis;Phut et Libyes fuerunt in auxilio eius.
NAH|3|10|Sed et ipsa in transmigrationem ducta est,ivit in captivitatem.Parvuli eius elisi suntin capite omnium viarum;et super inclitos eius miserunt sortem,et omnes optimates eius constricti sunt in compedibus.
NAH|3|11|Et tu ergo inebriaberis,eris despecta;et tu quaeresrefugium ab inimico.
NAH|3|12|Omnes munitiones tuae sicut ficuscum ficis praecocibus:si concussae fuerint,cadent in os comedentis.
NAH|3|13|Ecce populus tuus,mulieres in medio tui;inimicis tuis late patebuntportae terrae tuae;devorabit ignis vectes tuos.
NAH|3|14|Aquam propter obsidionem hauri tibi,firma munitiones tuas;intra in lutum et calca argillam,tene typum laterum.
NAH|3|15|Ibi comedet te ignis,peribis gladio,devorabit te ut bruchus.Augere ut bruchus,multiplicare ut locusta.
NAH|3|16|Plures fecisti negotiatores tuosquam stellae sint caeli;bruchus exuit pellemet avolavit.
NAH|3|17|Custodes tui quasi locustae,et scribae tui quasi agmen locustarum,quae considunt in saepibusin die frigoris;sol ortus est,et avolaverunt,non est cognitus locus earum,ubi fuerint.
NAH|3|18|Dormiunt pastores tui, rex Assyriae,requiescunt principes tui;dispersus est populus tuus in montibus,et non est qui congreget.
NAH|3|19|Non est remedium fracturae tuae,insanabilis est plaga tua;omnes, qui audierint auditionem tuam,plaudent manibus super te,quia super quem non transiitmalitia tua semper? ".
HAB|1|1|Oraculum, quod vidit Habacuc propheta.
HAB|1|2|Usquequo, Domine, clamabo,et non exaudis?Vociferabor ad te: " Violentia! ",et non salvas?
HAB|1|3|Quare ostendisti mihi iniquitatemet malitiam vides?Et vastitas et violentia est coram me,et facta est contentio, et iurgium exoritur.
HAB|1|4|Propter hoc languet lex,et non pervenit usque ad finem iudicium.Quia impius praevalet adversus iustum,propterea egreditur iudicium perversum.
HAB|1|5|" Aspicite in gentibus et videte,admiramini et obstupescite,quia opus facio in diebus vestris,quod nemo credet, cum narrabitur.
HAB|1|6|Quia ecce ego suscitabo Chaldaeos,gentem amaram et velocem,ambulantem super latitudinem terrae,ut possideat tabernacula non sua.
HAB|1|7|Horribilis et terribilis est,ex semetipsa iudicium eiuset maiestas eius egredietur.
HAB|1|8|Leviores pardis equi eiuset saeviores lupis deserti;et accurrunt equites eius:equites namque eius de longe venient,volabunt quasi aquilafestinans ad comedendum.
HAB|1|9|Omnes, ut violentiam faciant, venient,omnes facies eorum ventus urens;et congregabunt quasi arenam captivos.
HAB|1|10|Et ipsa reges subsannabit,tyrannis illudet;ipsa super omnem munitionem ridebitet comportabit aggerem et capiet eam.
HAB|1|11|Tunc ultra progrediens quasi ventus pertransibitet constituet fortitudinem suam deum suum ".
HAB|1|12|Numquid non tu a principio, Domine,Deus meus, sanctus meus,qui non morieris?Domine, ad iudicium posuisti eam; petra mea, ad corripiendum fundasti eam.
HAB|1|13|Mundi sunt oculi tui, ne videas malum;et respicere ad iniquitatem non poteris.Quare respicis super inique agentes et taces, devorante impio iustiorem se?
HAB|1|14|Fecisti homines quasi pisces maris,quasi reptile non habens principem super se.
HAB|1|15|Omnes in hamo sublevat,trahit eos in sagena suaet congregat in rete suo;super hoc laetatur et exsultat.
HAB|1|16|Propterea immolat sagenae suaeet sacrificat reti suo,quia in ipsis incrassata est portio eius,et cibus eius pinguis.
HAB|1|17|Propter hoc ergo evaginabit gladium suum semper,ut interficiat gentes sine misericordia?
HAB|2|1|Super custodiam meam staboet consistam super speculamet contemplabor, ut videam quid dicat mihiet quid respondeat ad querelam meam.
HAB|2|2|Et respondit mihi Dominus et dixit: Scribe visumet explana eum super tabulas,ut percurrat, qui legerit eum.
HAB|2|3|Quia adhuc visus ad tempus constitutum,sed anhelat in finem et non mentietur;si moram fecerit, exspecta illum,quia veniens veniet et non tardabit.
HAB|2|4|Ecce languidus, in quo non est anima recta;iustus autem in fide sua vivet ".
HAB|2|5|Et profecto divitiae decipiunt virum superbum,et non perveniet ad finem;qui dilatat quasi infernus fauces suaset ipse quasi mors et non adimpletur:et congregat ad se omnes genteset coacervat ad se omnes populos.
HAB|2|6|Numquid non omnes isti super eum parabolam sumentet loquelam aenigmatum dicentes: Vae ei, qui multiplicat non sua - usquequo? Cet aggravat pignora super se! ".
HAB|2|7|Numquid non repente consurgent, qui mordeant te,et evigilabunt agitantes te,et eris in rapinam eis?
HAB|2|8|Quia tu spoliasti gentes multas,spoliabunt te omnes, qui reliqui fuerint de populis;propter sanguinem hominum et oppressionem terrae,civitatum et omnium habitantium in eis.
HAB|2|9|Vae, qui congregat lucrum iniustum in malum domui suae,ut ponat in excelso nidum suumet salvet se de manu mali!
HAB|2|10|Consilium cepisti in confusionem domui tuaeconcidendi populos multoset peccasti in animam tuam.
HAB|2|11|Quia lapis de pariete clamabit,et trabes de contignatione respondebit ei.
HAB|2|12|Vae, qui aedificat civitatem in sanguinibuset condit urbem in iniquitate!
HAB|2|13|Numquid non haec a Domino sunt exercituum,ut laborent populi pro igne,et gentes in vacuum fatigentur?
HAB|2|14|Quia replebitur terra cognitione gloriae Domini,sicut aquae operiunt mare.
HAB|2|15|Vae, qui potum dat amico suomittens venenum suum et inebrians eum,ut aspiciat nuditatem eius!
HAB|2|16|Repleris ignominia pro gloria;bibe tu quoque et denudare!Transibit ad te calix dexterae Domini,et veniet ignominia super gloriam tuam.
HAB|2|17|Quia vastitas Libani operiet te,et miseria animalium deterrebit tepropter sanguinem hominum et oppressionem terrae,civitatum et omnium habitantium in eis.
HAB|2|18|Quid prodest sculptile,quia sculpsit illud fictor suus;conflatile et oraculum mendax,quia speravit in figmento fictor eius, ut faceret simulacra muta?
HAB|2|19|Vae, qui dicit ligno: " Expergiscere! ", " Surge! " lapidi tacenti!Numquid ipse docere poterit?Ecce iste coopertus est auro et argento,et omnis spiritus non est in visceribus eius.
HAB|2|20|Dominus autem in templo sancto suo; sileat a facie eius omnis terra.
HAB|3|1|Oratio Habacuc prophetae.Secundum melodiam lamentationum.
HAB|3|2|Domine, audivi auditionem tuamet timui, Domine, opus tuum.In medio annorum vivifica illud,in medio annorum notum facies.Cum iratus fueris, misericordiae recordaberis.
HAB|3|3|Deus a Theman veniet,et Sanctus de monte Pharan. - Selah.Operit caelos gloria eius,et laudis eius plena est terra.
HAB|3|4|Splendor eius ut lux erit,radii ex manibus eius:ibi abscondita est fortitudo eius.
HAB|3|5|Ante faciem eius ibit mors,et egredietur pestis post pedes eius.
HAB|3|6|Stetit et concussit terram,aspexit et dissolvit gentes.Et contriti sunt montes saeculi,incurvati sunt colles antiquiab itineribus aeternitatis eius.
HAB|3|7|In afflictione vidi tentoria Chusan;turbantur pelles terrae Madian.
HAB|3|8|Numquid in fluminibus iratus es, Domine,aut in fluminibus furor tuusvel in mari indignatio tua?Quia ascendes super equos tuos,quadrigas tuas victrices.
HAB|3|9|Suscitans suscitabis arcum tuum,sagittis replevisti pharetram tuam. - Selah.In fluvios scindes terram,
HAB|3|10|viderunt te et doluerunt montes.Effuderunt aquas nubes,dedit abyssus vocem suam,in altum levavit manus suas.
HAB|3|11|Sol et luna steterunt in habitaculo suo,prae luce sagittarum tuarum discedunt,prae splendore fulgurantis hastae tuae.
HAB|3|12|In fremitu calcabis terram,in furore conteres gentes.
HAB|3|13|Egressus es in salutem populi tui,in salutem cum christo tuo.Percussisti caput de domo impii,denudasti fundamentum usque ad petram. - Selah.
HAB|3|14|Confodisti iaculis tuis caput bellatorum eius,venientium ut turbo ad dispergendum me;exsultatio eorum, sicut eius, qui devorat pauperem in abscondito.
HAB|3|15|Viam fecisti in mari equis tuis,in luto aquarum multarum.
HAB|3|16|Audivi, et conturbatus est venter meus,ad vocem contremuerunt labia mea. Ingreditur putredo in ossibus meis, et subter me vacillant gressus mei.Conquiescam in die tribulationis,ut ascendat super populum, qui invadit nos.
HAB|3|17|Ficus enim non florebit,et non erit fructus in vineis;mentietur opus olivae,et arva non afferent cibum;abscissum est de ovili pecus,et non est armentum in praesepibus.
HAB|3|18|Ego autem in Domino gaudeboet exsultabo in Deo salvatore meo.
HAB|3|19|Dominus Deus fortitudo meaet ponet pedes meos quasi cervorum et super excelsa mea deducet me.Magistro chori. Ad sonitum chordarum.
ZEPH|1|1|Verbum Domini, quod factum est ad Sophoniam filium Chusi filii Godoliae filii Amariae filii Ezechiae, in diebus Iosiae filii Amon regis Iudae.
ZEPH|1|2|" Auferens auferam omniaa facie terrae,dicit Dominus,
ZEPH|1|3|auferam hominem et pecus,auferam volatile caeliet pisces maris.Et ruinae impiorum erunt;et disperdam homines a facie terrae,dicit Dominus.
ZEPH|1|4|Et extendam manum meam super Iudamet super omnes habitantes Ierusalem;et disperdam de loco hoc reliquias Baalet nomina aedituorum cum sacerdotibus
ZEPH|1|5|et eos, qui adorant super tectamilitiam caeliet adorant et iurant in Dominoet iurant in Melchom,
ZEPH|1|6|et qui avertuntur de post tergum Domini,et qui non quaerunt Dominum nec investigant eum ".
ZEPH|1|7|Silete a facie Domini Dei,quia iuxta est dies Domini;quia praeparavit Dominus hostiam,sanctificavit vocatos suos.
ZEPH|1|8|" Et erit in die hostiae Domini:visitabo super principeset super filios regiset super omnes, qui induti suntveste peregrina;
ZEPH|1|9|et visitabo super omnem,qui arroganter ingreditur super limen in die illa,qui complent domum domini suiiniquitate et dolo.
ZEPH|1|10|Et erit in die illa,dicit Dominus,vox clamoris a porta Piscium,et ululatus ab urbe Nova,et contritio magna a collibus.
ZEPH|1|11|Ululate, habitatores Pilae,quia interiit omnis populus Chanaan,disperierunt omnes involuti argento.
ZEPH|1|12|Et erit in tempore illo:scrutabor Ierusalem in lucerniset visitabo super virosdefixos in faecibus suis,qui dicunt in cordibus suis:Non faciet bene Dominuset non faciet male".
ZEPH|1|13|Et erunt opes eorum in direptionem,et domus eorum in desertum;et aedificabunt domoset non habitabunt,et plantabunt vineaset non bibent vinum earum ".
ZEPH|1|14|Iuxta est dies Domini magnus,iuxta et velox nimis;vox diei Domini amara,tribulabitur ibi fortis.
ZEPH|1|15|Dies irae dies illa,dies tribulationis et angustiae,dies vastitatis et desolationis,dies tenebrarum et caliginis,dies nebulae et turbinis,
ZEPH|1|16|dies tubae et clangorissuper civitates munitaset super angulos excelsos.
ZEPH|1|17|Et tribulabo homines,et ambulabunt ut caeci,quia Domino peccaverunt;et effundetur sanguis eorum sicut humus,et viscera eorum sicut stercora.
ZEPH|1|18|Sed et argentum eorum et aurum eorumnon poterit liberare eosin die irae Domini;in igne zeli eiusdevorabitur omnis terra,quia consummationem cum festinatione facietcunctis habitantibus terram.
ZEPH|2|1|Convenite, congregamini,gens non amabilis,
ZEPH|2|2|priusquam dispergaminiquasi pulvis transeuntes,antequam veniat super vosira furoris Domini,antequam veniat super vosdies furoris Domini.
ZEPH|2|3|Quaerite Dominum,omnes mansueti terrae,qui iudicium eius estis operati;quaerite iustitiam, quaerite mansuetudinem,si quomodo abscondaminiin die furoris Domini.
ZEPH|2|4|Quia Gaza deserta erit,et Ascalon desolata,Azotum in meridie eicient,et Accaron eradicabitur.
ZEPH|2|5|Vae, qui habitatis funiculum maris, gens Cretensium!Verbum Domini super vos,Chanaan, terra Philisthinorum: Disperdam te,ita ut non sit inhabitator ".
ZEPH|2|6|Et erit funiculus marisrequies pastorum et caulae pecorum.
ZEPH|2|7|Et erit funiculus marisreliquiis domus Iudae:ibi pascentur,in domibus Ascalonis ad vesperam requiescent,quia visitabit eos Dominus Deus eorumet convertet sortem eorum.
ZEPH|2|8|" Audivi opprobrium Moabet blasphemias filiorum Ammon, qui exprobraverunt populo meoet magnificati sunt super terminos eorum.
ZEPH|2|9|Propterea vivo ego,dicit Dominus exercituum, Deus Israel,quia Moab ut Sodoma erit,et filii Ammon quasi Gomorra,possessio spinarum et acervi saliset desertum usque in aeternum;reliquiae populi mei diripient eos,et residui gentis meae possidebunt illos ".
ZEPH|2|10|Hoc eis eveniet pro superbia sua, quia blasphemaverunt et magnificati suntsuper populum Domini exercituum.
ZEPH|2|11|Horribilis Dominus super eos,quia attenuabit omnes deos terrae;et adorabunt eum, singuli de loco suo,omnes insulae gentium.
ZEPH|2|12|" Sed et vos, Aethiopes,interfecti gladio meo eritis ".
ZEPH|2|13|Et extendet manum suam super aquilonemet perdet Assyriam;et ponet Nineven in solitudinemet in aridam, quasi desertum.
ZEPH|2|14|Et accubabunt in medio eius greges,omne genus animalium.Et onocrotalus et ululain capitellis eius morabuntur;vox cantat in fenestra,corvus in limine,quoniam tabulatum cedrinum sublatum est.
ZEPH|2|15|Haec est civitas exsultans,habitans in confidentia,quae dicebat in corde suo: Ego sum, et extra me non est alia amplius! ".Quomodo facta est in desertum,cubile bestiae?Omnis, qui transit per eam,sibilabit et movebit manum suam.
ZEPH|3|1|Vae, provocatrix et inquinata,civitas violenta!
ZEPH|3|2|Non audivit vocem,non suscepit disciplinam;in Domino non est confisa,ad Deum suum non appropiavit.
ZEPH|3|3|Principes eius in medio eiusleones rugientes;iudices eius lupi deserti,ossa non relinquunt in mane.
ZEPH|3|4|Prophetae eius vaniloqui,viri fallaces;sacerdotes eius polluerunt sanctum, iniuste egerunt contra legem.
ZEPH|3|5|Dominus iustus in medio eiusnon faciet iniquitatem;mane, mane iudicium suum dabit, sicut lucem, quae non deficit;nescivit autem iniquus confusionem.
ZEPH|3|6|" Disperdidi gentes,dissipati sunt anguli earum;desertas feci vias eorum,dum non est qui transeat;desolatae sunt civitates eorum,non remanente viro nec ullo habitatore.
ZEPH|3|7|Dixi: Nunc timebis me,suscipies disciplinam!Et non evanescent ab oculis eius omnia, in quibus visitavi eam.Verumtamen acceleraverunt corrumpereomnes actiones suas.
ZEPH|3|8|Quapropter exspecta me,dicit Dominus,in die qua surgam ut testis;quia iudicium meum, ut congregem genteset colligam regna,ut effundam super eas indignationem meam,omnem iram furoris mei;in igne enim zeli meidevorabitur omnis terra.
ZEPH|3|9|Quia tunc reddam populislabium purum,ut invocent omnes in nomine Dominiet serviant ei umero uno.
ZEPH|3|10|Ultra flumina Aethiopiae,inde supplices mei,filii dispersorum meorumdeferent munus mihi.
ZEPH|3|11|In die illa non confunderissuper cunctis actionibus tuis,quibus praevaricata es in me;quia tunc auferam de medio tuimagniloquos superbos tuos,et non adicies exaltari ampliusin monte sancto meo.
ZEPH|3|12|Et derelinquam in medio tuipopulum pauperem et egenum ".Et sperabunt in nomine Dominireliquiae Israel.
ZEPH|3|13|Non facient iniquitatemnec loquentur mendacium;et non invenietur in ore eorumlingua dolosa,quoniam ipsi pascentur et accubabunt,et non erit qui exterreat.
ZEPH|3|14|Lauda, filia Sion;iubilate, Israel!Laetare et exsulta in omni corde,filia Ierusalem!
ZEPH|3|15|Abstulit Dominus iudicium tuum,avertit inimicos tuos;rex Israel, Dominus, in medio tui,non timebis malum ultra.
ZEPH|3|16|In die illa dicetur Ierusalem: Noli timere, Sion;ne dissolvantur manus tuae!
ZEPH|3|17|Dominus Deus tuus in medio tui,fortis ipse salvabit;gaudebit super te in laetitia,commotus in dilectione sua;exsultabit super te in laude
ZEPH|3|18|sicut in die conventus ". Auferam a te calamitatem,ut non ultra habeas super ea opprobrium.
ZEPH|3|19|Ecce ego interficiamomnes, qui afflixerunt tein tempore illo;et salvabo claudicantemet eam, quae eiecta fuerat, congregabo;et ponam eos in laudem et in nomen in omni terra confusionis eorum,
ZEPH|3|20|in tempore illo, quo adducam vos,et in tempore, quo congregabo vos. Dabo enim vos in nomen et in laudemomnibus populis terrae,cum convertero sortem vestramcoram oculis vestris ",dicit Dominus.
HAG|1|1|In anno secundo Darii regis, in mense sexto, in die prima men sis, factum est verbum Domini in manu Aggaei prophetae ad Zorobabel filium Salathiel ducem Iudae et ad Iesua filium Iosedec sacerdotem magnum dicens:
HAG|1|2|" Haec ait Dominus exercituum dicens: Populus iste dicit: "Nondum venit tempus domus Domini aedificandae" ".
HAG|1|3|Et factum est verbum Domini in manu Aggaei prophetae dicens:
HAG|1|4|" Numquid tempus vobis est, ut habitetis in domibus laqueatis, et domus ista deserta?
HAG|1|5|Et nunc haec dicit Dominus exercituum: Ponite corda vestra super vias vestras:
HAG|1|6|seminastis multum et intulistis parum, comedistis et non estis satiati, bibistis et non estis inebriati, operuistis vos et non estis calefacti, et, qui pro mercede operatus est, misit eam in sacculum pertusum.
HAG|1|7|Haec dicit Dominus exercituum: Ponite corda vestra super vias vestras.
HAG|1|8|Ascendite in montem, portate lignum et aedificate domum, et acceptabilis mihi erit et glorificabor, dicit Dominus.
HAG|1|9|Respexistis ad amplius, et ecce factum est minus; et intulistis in domum, et exsufflavi illud. Quam ob causam?, dicit Dominus exercituum. Quia domus mea deserta est, et vos festinatis unusquisque in domum suam.
HAG|1|10|Propter hoc super vos prohibiti sunt caeli, ne darent rorem, et terra prohibita est, ne daret fructum suum.
HAG|1|11|Et vocavi siccitatem super terram et super montes et super triticum et super vinum et super oleum et, quaecumque profert humus, et super homines et super iumenta et super omnem laborem manuum ".
HAG|1|12|Et audivit Zorobabel filius Salathiel et Iesua filius Iosedec sacerdos magnus et omnes reliquiae populi vocem Domini Dei sui et verba Aggaei prophetae, sicut misit eum Dominus Deus eorum ad ipsos; et timuit populus a facie Domini.
HAG|1|13|Et dixit Aggaeus nuntius Domini secundum mandatum Domini populo dicens: Ego vobiscum, dicit Dominus ".
HAG|1|14|Et suscitavit Dominus spiritum Zorobabel filii Salathiel ducis Iudae et spiritum Iesua filii Iosedec sacerdotis magni et spiritum reliquorum omnium de populo; et ingressi sunt et faciebant opus in domo Domini exercituum Dei sui.
HAG|1|15|In die vicesima et quarta mensis, in sexto mense, in anno secundo Darii regis.
HAG|2|1|In septimo mense, vicesima et prima mensis, factum est ver bum Domini in manu Aggaei prophetae dicens:
HAG|2|2|" Loquere ad Zorobabel filium Salathiel ducem Iudae et ad Iesua filium Iosedec sacerdotem magnum et ad reliquos populi dicens:
HAG|2|3|Quis in vobis est derelictus, qui vidit domum istam in gloria sua prima? Et quid vos videtis eam nunc? Numquid non ita est quasi non sit in oculis vestris?
HAG|2|4|Sed et nunc confortare, Zorobabel, dicit Dominus, et confortare, Iesua fili Iosedec sacerdos magne, et confortare, omnis popule terrae, dicit Dominus exercituum; et facite, quoniam ego vobiscum sum, dicit Dominus exercituum.
HAG|2|5|Verbum quod pepigi vobiscum, cum egrederemini de terra Aegypti, et spiritus meus stat in medio vestrum; nolite timere.
HAG|2|6|Quia haec dicit Dominus exercituum: Adhuc unum modicum est, et ego commovebo caelum et terram et mare et aridam.
HAG|2|7|Et movebo omnes gentes, et venient thesauri cunctarum gentium, et implebo domum istam gloria, dicit Dominus exercituum.
HAG|2|8|Meum est argentum et meum est aurum, dicit Dominus exercituum.
HAG|2|9|Maior erit gloria domus istius novissima plus quam prima, dicit Dominus exercituum; et in loco isto dabo pacem, dicit Dominus exercituum ".
HAG|2|10|In vicesima et quarta noni mensis, in anno secundo Darii, factum est verbum Domini ad Aggaeum prophetam dicens:
HAG|2|11|" Haec dicit Dominus exercituum: Interroga sacerdotes legem dicens:
HAG|2|12|Si tulerit homo carnem sanctificatam in ora vestimenti sui et tetigerit de summitate eius panem aut pulmentum aut vinum aut oleum aut omnem cibum, numquid sanctificabitur? ". Respondentes autem sacerdotes dixerunt: " Non.
HAG|2|13|Et dixit Aggaeus: " Si tetigerit pollutus cadavere omnia haec, numquid contaminabuntur? ". Et responderunt sacerdotes et dixerunt: " Contaminabuntur ".
HAG|2|14|Et respondit Aggaeus et dixit: " Sic populus iste et sic gens ista ante faciem meam, dicit Dominus, et sic omne opus manuum eorum et omnia, quae offerunt ibi, contaminata sunt.
HAG|2|15|Et nunc ponite corda vestra a die hac et supra: Antequam poneretur lapis super lapidem in templo Domini,
HAG|2|16|quid fuistis? Cum accederetis ad acervum viginti modiorum, erant decem; cum intraretis ad torcular, ut hauriretis quinquaginta lagenas, erant viginti.
HAG|2|17|Percussi vos ariditate et rubigine et grandine omnia opera manuum vestrarum, et non fuit in vobis qui reverteretur ad me, dicit Dominus.
HAG|2|18|Ponite corda vestra ex die ista et in futurum, a die vicesima et quarta noni mensis, a die, qua fundamenta iacta sunt templi Domini, ponite super cor vestrum.
HAG|2|19|Numquid adhuc semen in horreo est, et adhuc vinea et ficus et malogranatum et lignum olivae non portavit fructum? Ex die hac benedicam.
HAG|2|20|Et factum est verbum Domini secundo ad Aggaeum in vicesima et quarta mensis dicens:
HAG|2|21|" Loquere ad Zorobabel ducem Iudae dicens: Ego movebo caelum pariter et terram
HAG|2|22|et subvertam solium regnorum et conteram fortitudinem regnorum gentium et subvertam quadrigam et ascensores eius; et descendent equi et ascensores eorum, unusquisque percussus gladio fratris sui.
HAG|2|23|In die illo, dicit Dominus exercituum, assumam te, Zorobabel fili Salathiel, serve meus, dicit Dominus, et ponam te quasi signaculum, quia te elegi ", dicit Dominus exercituum.
ZECH|1|1|In mense octavo, in anno se cundo Darii, factum est verbum Domini ad Zachariam filium Barachiae filii Addo prophetam dicens:
ZECH|1|2|" Iratus est Dominus super patres vestros iracundia.
ZECH|1|3|Et dices ad eos: Haec dicit Dominus exercituum: Convertimini ad me, ait Dominus exercituum; et convertar ad vos, dicit Dominus exercituum.
ZECH|1|4|Ne sitis sicut patres vestri, ad quos clamabant prophetae priores dicentes: Haec dicit Dominus exercituum: Convertimini de viis vestris malis et de cogitationibus vestris malis; et non audierunt neque attenderunt ad me, dicit Dominus.
ZECH|1|5|Patres vestri ubi sunt? Et prophetae numquid in sempiternum vivent?
ZECH|1|6|Verumtamen verba mea et praecepta mea, quae mandavi servis meis prophetis, numquid non attigerunt patres vestros? Et conversi sunt et dixerunt: "Sicut cogitavit Dominus exercituum facere nobis, secundum vias nostras et secundum adinventiones nostras fecit nobis" ".
ZECH|1|7|In die vicesima et quarta undecimi mensis, qui est mensis Sabath, in anno secundo Darii, factum est verbum Domini ad Zachariam filium Barachiae filii Addo prophetam dicens:
ZECH|1|8|" Vidi per noctem, et ecce vir sedens super equum rufum et ipse stabat inter myrteta, quae erant in profundo; et post eum equi rufi, fulvi et albi.
ZECH|1|9|Et dixi: "Quid sunt isti, domine mi?". Et dixit ad me angelus, qui loquebatur in me: "Ego ostendam tibi quid sint isti".
ZECH|1|10|Et respondit vir, qui stabat inter myrteta, et dixit: "Isti sunt quos misit Dominus, ut perambularent terram".
ZECH|1|11|Et responderunt angelo Domini, qui stabat inter myrteta, et dixerunt: Perambulavimus terram, et ecce omnis terra habitatur et quiescit".
ZECH|1|12|Et respondit angelus Domini et dixit: "Domine exercituum, usquequo tu non misereberis Ierusalem et urbium Iudae, quibus iratus es? Iste septuagesimus annus est!".
ZECH|1|13|Et respondit Dominus angelo, qui loquebatur in me verba bona, verba consolatoria.
ZECH|1|14|Et dixit ad me angelus, qui loquebatur in me: "Clama dicens: Haec dixit Dominus exercituum: Zelatus sum Ierusalem et Sion zelo magno,
ZECH|1|15|sed ira magna ego irascor super gentes opulentas, quia ego iratus sum parum, ipsi vero adiuverunt in malum.
ZECH|1|16|Propterea haec dicit Dominus: Revertar ad Ierusalem in misericordiis. Domus mea aedificabitur in ea, ait Dominus exercituum, et perpendiculum extendetur super Ierusalem.
ZECH|1|17|Adhuc clama dicens: Haec dicit Dominus exercituum: Adhuc affluent civitates meae bonis, et consolabitur adhuc Dominus Sion et eliget adhuc Ierusalem".
ZECH|2|1|Et levavi oculos meos et vidi, et ecce quattuor cornua;
ZECH|2|2|et dixi ad angelum, qui loquebatur in me: "Quid sunt haec?". Et dixit ad me: "Haec sunt cornua, quae ventilaverunt Iudam et Israel et Ierusalem".
ZECH|2|3|Et ostendit mihi Dominus quattuor fabros;
ZECH|2|4|et dixi: "Quid isti veniunt facere?". Qui respondit dicens: "Haec sunt cornua, quae ventilaverunt Iudam per singulos viros, ut nemo eorum levaret caput suum; et venerunt isti deterrere ea, ut deiciant cornua gentium, quae levaverunt cornu super terram Iudae, ut dispergerent eam".
ZECH|2|5|Et levavi oculos meos et vidi; et ecce vir, et in manu eius funiculus mensorum.
ZECH|2|6|Et dixi: "Quo tu vadis?". Et dixit ad me: "Ut metiar Ierusalem et videam, quanta sit latitudo eius et quanta longitudo eius".
ZECH|2|7|Et ecce angelus, qui loquebatur in me, egrediebatur, et angelus alius egrediebatur in occursum eius;
ZECH|2|8|et dixit ad eum: "Curre, loquere ad puerum istum dicens: Absque muris habitabitur Ierusalem prae multitudine hominum et iumentorum in medio eius.
ZECH|2|9|Et ego ero ei, ait Dominus, murus ignis in circuitu et in gloria ero in medio eius.
ZECH|2|10|Heu, heu! Fugite de terra aquilonis, dicit Dominus, quoniam in quattuor ventos caeli dispersi vos, dicit Dominus.
ZECH|2|11|Heu, Sion, fuge, quae habitas apud filiam Babylonis!
ZECH|2|12|Quia haec dicit Dominus exercituum, cuius gloria misit me ad gentes, quae spoliaverunt vos: Qui tetigerit vos, tangit pupillam oculi mei.
ZECH|2|13|Quia ecce ego levo manum meam super eos, et erunt praeda servorum suorum; et cognoscetis quia Dominus exercituum misit me.
ZECH|2|14|Iubila et laetare, filia Sion,quia ecce ego venioet habitabo in medio tui,ait Dominus.
ZECH|2|15|Et applicabuntur gentes multaead Dominum in die illaet erunt ei in populum.Et habitabo in medio tui,et scies quia Dominus exercituummisit me ad te.
ZECH|2|16|Et possidebit Dominus Iudampartem suam super terram sanctamet eliget adhuc Ierusalem.
ZECH|2|17|Sileat omnis caro a facie Domini,quia consurrexit de habitaculo sancto suo".
ZECH|3|1|Et ostendit mihi Iesua sacer dotem magnum stantem coram angelo Domini; et Satan stabat a dextris eius, ut adversaretur ei.
ZECH|3|2|Et dixit angelus Domini ad Satan: "Increpet Dominus in te, Satan! Et increpet Dominus in te, qui elegit Ierusalem! Numquid non iste torris est erutus de igne?".
ZECH|3|3|Et Iesua erat indutus vestibus sordidis et stabat ante faciem angeli.
ZECH|3|4|Qui respondit et ait ad eos, qui stabant coram se, dicens: "Auferte vestimenta sordida ab eo". Et dixit ad eum: "Ecce, abstuli a te iniquitatem tuam; induam te mutatoriis".
ZECH|3|5|Et dixit: "Ponite cidarim mundam super caput eius". Et posuerunt cidarim mundam super caput eius et induerunt eum vestibus; et angelus Domini stabat.
ZECH|3|6|Et contestabatur angelus Domini Iesua dicens:
ZECH|3|7|"Haec dicit Dominus exercituum: Si in viis meis ambulaveris et ministerium meum custodieris, tu quoque iudicabis domum meam et custodies atria mea; et dabo tibi accessum inter eos, qui nunc hic assistunt.
ZECH|3|8|Audi, Iesua sacerdos magne, tu et amici tui, qui sedent coram te, quia viri portendentes sunt: Ecce enim ego adduco servum meum Germen.
ZECH|3|9|Quia ecce lapis, quem dedi coram Iesua: super lapidem unum septem oculi sunt; ecce ego caelabo sculpturam eius, ait Dominus exercituum, et auferam iniquitatem terrae illius in die una.
ZECH|3|10|In die illa, oraculum Domini exercituum, vocabit vir amicum suum subter vitem et subter ficum".
ZECH|4|1|Et reversus est angelus, qui loquebatur in me, et excitavit me quasi virum, qui excitatur de somno suo.
ZECH|4|2|Et dixit ad me: "Quid tu vides?". Et dixi: "Vidi: et ecce candelabrum aureum totum, et ampulla super caput ipsius, et septem lucernae eius super illud, et septena infusoria lucernis, quae erant super caput eius.
ZECH|4|3|Et duae olivae super illud, una a dextris ampullae et una a sinistris eius".
ZECH|4|4|Et respondi et aio ad angelum, qui loquebatur in me, dicens: "Quid sunt haec, domine mi?".
ZECH|4|5|Et respondit angelus, qui loquebatur in me, et dixit ad me: "Numquid nescis quid sunt haec?". Et dixi: "Non, domine mi".
ZECH|4|6|Et respondit et ait ad me dicens: "Hoc est verbum Domini ad Zorobabel dicens: Non in exercitu nec in robore sed in spiritu meo, dicit Dominus exercituum.
ZECH|4|7|Quis tu, mons magne, coram Zorobabel? Eris in planum. Et educet lapidem primarium inter clamores: Quam venustus!
ZECH|4|8|Et factum est verbum Domini ad me dicens:
ZECH|4|9|Manus Zorobabel fundaverunt domum istam et manus eius perficient eam, et scietis quia Dominus exercituum misit me ad vos.
ZECH|4|10|Quis enim despexit diem initiorum parvorum? Et laetabuntur et videbunt lapidem stanneum in manu Zorobabel. Septem illae oculi sunt Domini, qui discurrunt in universa terra".
ZECH|4|11|Et respondi et dixi ad eum: "Quid sunt duae olivae istae ad dexteram candelabri et ad sinistram eius?".
ZECH|4|12|Et respondi secundo et dixi ad eum: "Quid sunt duo rami olivarum, qui duabus fistulis aureis effundunt ex se aurum?".
ZECH|4|13|Et ait ad me dicens: "Numquid nescis quid sunt haec?". Et dixi: "Non, domine mi".
ZECH|4|14|Et dixit: "Isti sunt duo filii olei, qui assistunt Dominatori universae terrae".
ZECH|5|1|Et conversus sum et levavi ocu los meos et vidi: et ecce volu men volans.
ZECH|5|2|Et dixit ad me: "Quid tu vides?". Et dixi: "Ego video volumen volans; longitudo eius viginti cubitorum et latitudo eius decem cubitorum".
ZECH|5|3|Et dixit ad me: "Haec est maledictio, quae egreditur super faciem omnis terrae; quia omnis fur hinc iuxta illud expurgatur, et omnis periurus illinc iuxta illud expurgatur.
ZECH|5|4|Educo illud, dicit Dominus exercituum, et veniet ad domum furis et ad domum iurantis in nomine meo mendaciter; et commorabitur in medio domus eius, et consumet eam et ligna eius et lapides eius".
ZECH|5|5|Et egressus est angelus, qui loquebatur in me, et dixit ad me: "Leva, quaeso, oculos tuos et vide. Quid est hoc, quod egreditur?".
ZECH|5|6|Et dixi: "Quidnam est?". Et ait: "Haec est epha egrediens". Et dixit: Hoc est peccatum eorum in universa terra".
ZECH|5|7|Et ecce operculum plumbi elevatum est, et ecce mulier una sedens in medio ephae.
ZECH|5|8|Et dixit: "Haec est impietas". Et proiecit eam in epham et misit massam plumbeam in os eius.
ZECH|5|9|Et levavi oculos meos et vidi: et ecce duae mulieres egredientes, et ventus in alis earum, et habebant alas quasi alas milvi; et levaverunt epham inter terram et caelum.
ZECH|5|10|Et dixi ad angelum, qui loquebatur in me: "Quo istae deferunt epham?".
ZECH|5|11|Et dixit ad me: "Ut aedificetur ei domus in terra Sennaar; et, postquam constructa fuerit, ponetur ibi super basem suam".
ZECH|6|1|Et rursus levavi oculos meos et vidi: et ecce quattuor quadrigae egredientes de medio duorum montium; et montes, montes aerei.
ZECH|6|2|In quadriga prima equi rufi, et in quadriga secunda equi nigri,
ZECH|6|3|et in quadriga tertia equi albi, et in quadriga quarta equi varii.
ZECH|6|4|Et respondi et dixi ad angelum, qui loquebatur in me: "Quid sunt haec, domine mi?".
ZECH|6|5|Et respondit angelus et ait ad me: "Isti sunt quattuor venti caeli, qui egrediuntur, postquam steterunt coram Dominatore omnis terrae".
ZECH|6|6|In qua erant equi nigri, egrediebantur in terram aquilonis, et albi egressi sunt post eos, et varii egressi sunt ad terram austri.
ZECH|6|7|Et equi fortes exierunt et quaerebant ire et discurrere per terram. Et dixit: "Ite, perambulate terram". Et perambulaverunt terram.
ZECH|6|8|Et vocavit me et locutus est ad me dicens: "Ecce, qui egrediuntur in terram aquilonis requiescere fecerunt spiritum meum in terra aquilonis".
ZECH|6|9|Et factum est verbum Domini ad me dicens:
ZECH|6|10|"Sume ab his, qui de captivitate sunt, ab Holdai et a Thobia et ab Iedaia, et venies tu in die illa et intrabis domum Iosiae filii Sophoniae, qui venerunt de Babylone.
ZECH|6|11|Et sumes argentum et aurum et facies coronam et pones in capite Iesua filii Iosedec, sacerdotis magni,
ZECH|6|12|et loqueris ad eum dicens: Haec ait Dominus exercituum dicens: Ecce vir, Germen nomen eius; et in loco suo aliquid germinabit et aedificabit templum Domini.
ZECH|6|13|Et ipse exstruet templum Domini; et ipse portabit gloriam et sedebit et dominabitur super solio suo; et erit sacerdos ad dexteram eius, et consilium pacis erit inter illos duos.
ZECH|6|14|Et corona erit Helem et Thobiae et Iedaiae et Hen filio Sophoniae memoriale in templo Domini.
ZECH|6|15|Et qui procul sunt, venient et aedificabunt in templo Domini; et scietis quia Dominus exercituum misit me ad vos. Erit autem hoc, si oboedieritis voci Domini Dei vestri" ".
ZECH|7|1|Et factum est in anno quarto Darii regis, factum est verbum Domini ad Zachariam in quarta mensis noni, qui est Casleu.
ZECH|7|2|Et Bethel miserat Sarasar et Regemmelech et viros, qui erant cum eo, ad deprecandam faciem Domini,
ZECH|7|3|ut dicerent sacerdotibus domus Domini exercituum et prophetis loquentes: Numquid flendum est mihi in quinto mense vel ieiunandum, sicut iam feci multis annis? ".
ZECH|7|4|Et factum est verbum Domini exercituum ad me dicens:
ZECH|7|5|" Loquere ad omnem populum terrae et ad sacerdotes dicens: Cum ieiunaretis et plangeretis in quinto et septimo mense per hos septuaginta annos, numquid revera ieiunastis mihi?
ZECH|7|6|Et cum comedistis et bibistis, numquid non vobis comedistis et vobismetipsis bibistis?
ZECH|7|7|Numquid non sunt verba, quae locutus est Dominus in manu prophetarum priorum, cum adhuc Ierusalem habitaretur et esset opulenta, ipsa et urbes in circuitu eius, et Nageb habitaretur simul cum Sephela? ".
ZECH|7|8|Et factum est verbum Domini ad Zachariam dicens:
ZECH|7|9|" Haec ait Dominus exercituum dicens: Iudicium verum iudicate et misericordiam et miserationes facite unusquisque cum fratre suo;
ZECH|7|10|et viduam et pupillum et advenam et pauperem nolite calumniari, et malum unusquisque contra fratrem suum nolite cogitare in corde vestro.
ZECH|7|11|Et noluerunt attendere; et opposuerunt dorsum rebelle et aures suas aggravaverunt, ne audirent.
ZECH|7|12|Et cor suum posuerunt adamantem, ne audirent legem et verba, quae misit Dominus exercituum in spiritu suo per manum prophetarum priorum, et facta est indignatio magna a Domino exercituum.
ZECH|7|13|Et factum est, sicut cum clamaret, et ipsi non audierunt, sic clamabunt, et non exaudiam, dicit Dominus exercituum.
ZECH|7|14|Et disperdam eos per omnes gentes, quas nesciunt; et terra desolata est post eos, ita ut non esset transiens et revertens. Et posuerunt terram desiderabilem in desertum ".
ZECH|8|1|Et factum est verbum Domini exercituum dicens:
ZECH|8|2|" Haec dicit Dominus exercituum:Zelatus sum Sion zelo magnoet ardore magno zelatus sum eam.
ZECH|8|3|Haec dicit Dominus: Reversus sum ad Sion et habitabo in medio Ierusalem; et vocabitur Ierusalem civitas Veritatis, et mons Domini exercituum mons Sanctitatis.
ZECH|8|4|Haec dicit Dominus exercituum: Adhuc sedebunt senes et anus in plateis Ierusalem et unusquisque cum baculo suo in manu sua prae multitudine dierum;
ZECH|8|5|et plateae civitatis complebuntur pueris et puellis ludentibus in plateis eius.
ZECH|8|6|Haec dicit Dominus exercituum: Si videbitur difficile in oculis reliquiarum populi huius in diebus illis, numquid etiam in oculis meis difficile erit?, dicit Dominus exercituum.
ZECH|8|7|Haec dicit Dominus exercituum:Ecce ego salvabo populum meum de terra orientiset de terra occasus solis:
ZECH|8|8|et adducam eos,et habitabunt in medio Ierusalem;et erunt mihi in populum,et ego ero eis in Deumin veritate et iustitia.
ZECH|8|9|Haec dicit Dominus exercituum: Confortentur manus vestrae, qui auditis in his diebus sermones istos per os prophetarum in die, qua fundata est domus Domini exercituum, ut templum aedificaretur.
ZECH|8|10|Siquidem ante dies istosmerces hominis non erat,nec merces iumenti erat,neque introeunti neque exeuntierat pax prae tribulatione;et dimisi omnes homines,unumquemque contra proximum suum.
ZECH|8|11|Nunc autem non iuxta dies priores ego sumreliquiis populi huius,dicit Dominus exercituum;
ZECH|8|12|sed semen pacis erit:vinea dabit fructum suum,et terra dabit proventum suum,et possidere faciamreliquias populi huiusuniversa haec.
ZECH|8|13|Et erit: sicut eratis maledictio in gentibus, domus Iudae et domus Israel, sic salvabo vos, et eritis benedictio. Nolite timere; confortentur manus vestrae.
ZECH|8|14|Quia haec dicit Dominus exercituum: Sicut cogitavi, ut affligerem vos, cum ad iracundiam provocassent patres vestri me, dicit Dominus exercituum,
ZECH|8|15|et non sum misertus, sic conversus cogitavi in diebus istis, ut benefaciam Ierusalem et domui Iudae; nolite timere.
ZECH|8|16|Haec sunt ergo, quae facietis: Loquimini veritatem unusquisque cum proximo suo et iudicium pacis iudicate in portis vestris,
ZECH|8|17|et unusquisque malum contra amicum suum ne cogitetis in cordibus vestris et iuramentum mendax ne diligatis: omnia enim haec sunt quae odi, dicit Dominus.
ZECH|8|18|Et factum est verbum Domini exercituum ad me dicens:
ZECH|8|19|" Haec dicit Dominus exercituum: Ieiunium quarti et ieiunium quinti et ieiunium septimi et ieiunium decimi erit domui Iudae in gaudium et laetitiam et in sollemnitates praeclaras; veritatem tantum et pacem diligite.
ZECH|8|20|Haec dicit Dominus exercituum: Adhuc venient populi et habitatores civitatum magnarum,
ZECH|8|21|et ibunt habitatores unius ad alteram dicentes: "Eamus, ut deprecemur faciem Domini et quaeramus Dominum exercituum; vadam etiam ego".
ZECH|8|22|Et venient populi multi et gentes robustae ad quaerendum Dominum exercituum in Ierusalem et deprecandam faciem Domini.
ZECH|8|23|Haec dicit Dominus exercituum: In diebus illis apprehendent decem homines ex omnibus linguis gentium, apprehendent fimbriam viri Iudaei dicentes: "Ibimus vobiscum; audivimus enim quoniam Deus vobiscum est" ".
ZECH|9|1|Oraculum. Verbum Domini in terra Ha drachet Damasci requiei eius,quia Domini est oculus Aramsicut omnes tribus Israel.
ZECH|9|2|Emath quoque in terminis eiuset Tyrus et Sidon, quae sapiens est valde.
ZECH|9|3|Et aedificavit Tyrus munitionem suamet coacervavit argentum quasi pulveremet aurum ut lutum platearum.
ZECH|9|4|Ecce Dominus possidebit eamet percutiet in mari fortitudinem eius;et haec igni devorabitur.
ZECH|9|5|Videbit Ascalon et timebit,et Gaza dolore torquetur nimis,et Accaron, quoniam confusa est spes eius;et peribit rex de Gaza,et Ascalon non habitabitur.
ZECH|9|6|Et habitabit spurius in Azoto,et disperdam superbiam Philisthim.
ZECH|9|7|Et auferam sanguinem eius de ore eiuset abominationes eius de medio dentium eius,et relinquetur etiam ipse Deo nostro,et erit quasi dux in Iuda,et Accaron quasi Iebusaeus.
ZECH|9|8|Et circumdabo domum meam ut praesidiumcontra euntes et revertentes;et non transibit super eos ultra exactor,quia nunc vidi in oculis meis.
ZECH|9|9|Exsulta satis, filia Sion;iubila, filia Ierusalem.Ecce rex tuus venit tibiiustus et salvator ipse,pauper et sedens super asinumet super pullum filium asinae.
ZECH|9|10|Et disperdam currum ex Ephraimet equum de Ierusalem;et confringetur arcus belli,et loquetur pacem gentibus.Et imperium eius a mari usque ad mareet a flumine usque ad fines terrae.
ZECH|9|11|Tu quoque: in sanguine testamenti tuiextraho vinctos tuos de lacu,in quo non est aqua.
ZECH|9|12|Convertimini ad munitionem,vincti spei;hodie quoque annuntians:Duplicia reddam tibi.
ZECH|9|13|Nam extendi mihi Iudam quasi arcum,implevi Ephraim;et suscitabo filios tuos, Sion,super filios tuos, Graecia,et ponam te quasi gladium fortium.
ZECH|9|14|Et Dominus super eos videbitur,et exibit ut fulgur iaculum eius;et Dominus Deus in tuba canetet vadet in procellis austri.
ZECH|9|15|Dominus exercituum proteget eos;et devorabunt et conculcabunt lapides fundaeet bibent, agitabuntur quasi vinoet replebuntur ut phialae et quasi cornua altaris.
ZECH|9|16|Et salvabit eos Dominus Deus eorumin die illaut gregem populi sui,quia lapides coronaefulgebunt super terram eius.
ZECH|9|17|Quid enim bonum eius est,et quid pulchrum eius!Frumentum succrescere facit iuvenes,et mustum virgines.
ZECH|10|1|Petite a Domino pluviamin tempore pluviae serotinae.Dominus facit fulguraet pluviam imbris dabit eis,singulis herbam in agro.
ZECH|10|2|Quia theraphim loquuntur inania,et divini vident mendacium,et somnia loquuntur vana,vane consolantur;idcirco migrant quasi grex,affliguntur, quia non est eis pastor.
ZECH|10|3|Super pastores iratus est furor meus,et super hircos visitabo:certe visitat Dominus exercituumgregem suum, domum Iudae,et faciet eos quasi equum gloriae suaein bello.
ZECH|10|4|Ex ipso angulus,ex ipso paxillus,ex ipso arcus proelii,ex ipso egredietur omnis exactor simul.
ZECH|10|5|Et erunt quasi fortesconculcantes lutum viarum in proelioet bellabunt, quia Dominus cum eis; et confundentur ascensores equorum.
ZECH|10|6|Et confortabo domum Iudaeet domum Ioseph salvaboet reducam eos, quia miserebor eorum;et erunt, sicut non proiecissem eos:ego enim Dominus Deus eorum et exaudiam eos.
ZECH|10|7|Et erunt quasi fortes Ephraim,et laetabitur cor eorum quasi a vino,et filii eorum videbunt et laetabuntur,et exsultabit cor eorum in Domino.
ZECH|10|8|Sibilabo eis et congregabo illos,quia redemi eos,et multi erunt, sicut multi ante fuerant.
ZECH|10|9|Et seminabo eos in populis,et de longe recordabuntur mei;et alent filios suos et revertentur.
ZECH|10|10|Et reducam eos de terra Aegyptiet de Assyria congregabo eoset ad terram Galaad et Libani adducam eos,et non invenietur eis locus.
ZECH|10|11|Et transibunt per mare angustiae,et percutiet in mari fluctus,et exiccabuntur omnia profunda fluminis;et humiliabitur superbia Assyriae,et sceptrum Aegypti recedet.
ZECH|10|12|Confortabo eos in Domino,et in nomine eius ambulabunt ",dicit Dominus.
ZECH|11|1|Aperi, Libane, portas tuas,et comedat ignis cedros tuas.
ZECH|11|2|Ulula, abies, quia cecidit cedrus,quoniam magnifici vastati sunt;ululate, quercus Basan,quoniam corruit saltus impervius.
ZECH|11|3|Vox ululatus pastorum,quia vastata est magnificentia eorum;vox rugitus leonum,quoniam vastata est superbia Iordanis.
ZECH|11|4|Haec dicit Dominus Deus meus: " Pasce pecora occisionis.
ZECH|11|5|Quae, qui emunt, occidunt et non dolent; et, qui vendunt ea, dicunt: Benedictus Dominus! Dives factus sum". Et pastores eorum non miserentur eorum.
ZECH|11|6|Et ego non miserebor ultra super habitantes terram, dicit Dominus; ecce ego tradam homines, unumquemque in manu proximi sui et in manu regis sui; et concident terram, et non eruam de manu eorum ".
ZECH|11|7|Et ego pavi pecus occisionis pro mercatoribus gregis. Et assumpsi mihi duas virgas: unam vocavi Gratiam et alteram vocavi Funiculum; et pavi gregem.
ZECH|11|8|Et succidi tres pastores in mense uno, et taeduit eorum animam meam; siquidem et animam eorum taeduit mei.
ZECH|11|9|Et dixi: " Non pascam vos. Quae moritura est, moriatur; et, quae succidenda est, succidatur; et reliquae devorent unaquaeque carnem proximae suae ".
ZECH|11|10|Et tuli virgam meam, quae vocabatur Gratia, et abscidi eam, ut irritum facerem foedus meum, quod percussi cum omnibus populis.
ZECH|11|11|Et irritum factum est in die illa; et cognoverunt mercatores gregis, qui observabant me, quia verbum Domini est.
ZECH|11|12|Et dixi ad eos: " Si bonum est in oculis vestris, afferte mercedem meam et, si non, quiescite ". Et appenderunt mercedem meam triginta siclos argenteos.
ZECH|11|13|Et dixit Dominus ad me: " Proice illud in thesaurum, decorum pretium, quo appretiatus sum ab eis ".Et tuli triginta siclos argenteos et proieci illos in domum Domini in thesaurum.
ZECH|11|14|Et praecidi virgam meam secundam, quae appellabatur Funiculus, ut dissolverem germanitatem inter Iudam et Israel.
ZECH|11|15|Et dixit Dominus ad me: Adhuc sume tibi vasa pastoris stulti;
ZECH|11|16|quia ecce ego suscitabo pastorem in terra,qui perituram ovem non visitabit,dispersam non quaeretet contritam non sanabitet stantem non sustinebitet carnes pinguium comedetet ungulas earum confringet.
ZECH|11|17|Vae stulto meo pastoriderelinquenti gregem!Gladius super brachium eiuset super oculum dextrum eius;brachium eius ariditate siccetur,et oculus dexter eius tenebrescens obscuretur ".
ZECH|12|1|Oraculum. Verbum Domini super Israel et super Iudam. Oraculum Domini, qui extendit caelum et fundat terram et fingit spiritum hominis in eo:
ZECH|12|2|" Ecce ego pono Ierusalem pateram crapulae omnibus populis in circuitu. Hoc erit in obsidione contra Ierusalem.
ZECH|12|3|Et erit: in die illa ponam Ierusalem lapidem portandum cunctis populis; omnes portantes eam concisione lacerabuntur, et colligentur adversus eam omnes gentes terrae.
ZECH|12|4|In die illa, dicit Dominus, percutiam omnem equum in stuporem et ascensorem eius in amentiam; et super domum Iudae aperiam oculos meos et omnem equum populorum percutiam caecitate.
ZECH|12|5|Et dicent duces Iudae in corde suo: "Robur habitantium Ierusalem est in Domino exercituum, Deo eorum".
ZECH|12|6|In die illa ponam duces Iudae sicut ollam ignis super ligna et sicut facem ignis super fenum; et devorabunt ad dexteram et ad sinistram omnes populos in circuitu, et habitabitur Ierusalem rursus in loco suo.
ZECH|12|7|Et salvabit Dominus prius tabernacula Iudae, ut non elevetur gloria domus David et gloria habitantium Ierusalem contra Iudam.
ZECH|12|8|In die illa proteget Dominus habitatores Ierusalem; et erit, qui offenderit ex eis in die illa quasi David, et domus David quasi Deus, sicut angelus Domini in conspectu eorum.
ZECH|12|9|Et erit: in die illa quaeram conterere omnes gentes, quae veniunt contra Ierusalem,
ZECH|12|10|et effundam super domum David et super habitatores Ierusalem spiritum gratiae et precum; et aspicient ad me. Quem confixerunt, plangent quasi planctu super unigenitum et dolebunt super eum, ut doleri solet super primogenitum.
ZECH|12|11|In die illa magnus erit planctus in Ierusalem sicut planctus Adadremmon in campo Mageddo;
ZECH|12|12|et planget terra, singulae familiae seorsum:familia domus David seorsumet mulieres eorum seorsum;familia domus Nathan seorsumet mulieres eorum seorsum;
ZECH|12|13|familia domus Levi seorsumet mulieres eorum seorsum;familia Semei seorsumet mulieres eorum seorsum;
ZECH|12|14|omnes reliquae familiae, singulae familiae seorsumet mulieres eorum seorsum.
ZECH|13|1|In die illa erit fons patens domui David et habitantibus Ierusalem pro peccatis et immunditia.
ZECH|13|2|Et erit in die illa, dicit Dominus exercituum, disperdam nomina idolorum de terra, et non memorabuntur ultra; et pseudoprophetas et spiritum immundum auferam de terra.
ZECH|13|3|Et erit: cum prophetaverit quispiam ultra, dicent ei pater eius et mater eius, qui genuerunt eum: "Non vives, quia mendacium locutus es in nomine Domini"; et configent eum pater eius et mater eius, qui genuerunt eum, cum prophetaverit.
ZECH|13|4|Et erit: in die illa confundentur prophetae, unusquisque ex visione sua, cum prophetaverit; nec operientur pallio saccino, ut mentiantur,
ZECH|13|5|sed dicet: "Non sum propheta; homo operans terram ego sum, quoniam terra est possessio mea ab adulescentia mea".
ZECH|13|6|Et dicetur ei: "Quid sunt plagae istae in medio manuum tuarum?". Et dicet: "His plagatus sum in domo eorum, qui diligebant me".
ZECH|13|7|Framea, suscitare super pastorem meumet super virum cohaerentem mihi,dicit Dominus exercituum.Percute pastorem, et dispergentur oves,et convertam manum meam contra parvulos.
ZECH|13|8|Et erit in omni terra,dicit Dominus:partes duae in ea dispergentur et deficient,et tertia pars relinquetur in ea;
ZECH|13|9|et ducam tertiam partem per ignemet purgabo eos, sicut purgatur argentum,et probabo eos, sicut probatur aurum:ipse vocabit nomen meum,et ego exaudiam eum.Dicam: Populus meus est ille;et ipse dicet: "Dominus est Deus meus".
ZECH|14|1|Ecce venit dies Domino, et dividentur spolia tua in me dio tui,
ZECH|14|2|et congregabo omnes gentes ad Ierusalem in proelium, et capietur civitas, et vastabuntur domus, et mulieres violabuntur; et egredietur media pars civitatis in captivitatem, et reliquum populi non auferetur ex urbe.
ZECH|14|3|Et egredietur Dominus et proeliabitur contra gentes illas, sicut proeliatus est in die certaminis.
ZECH|14|4|Et stabunt pedes eius in die illa super montem Olivarum, qui est contra Ierusalem ad orientem; et scindetur mons Olivarum ex media parte sui ad orientem et ad occidentem, praerupto grandi valde, et separabitur medium montis ad aquilonem et medium eius ad meridiem.
ZECH|14|5|Et fugietis ad vallem montium eorum, quoniam vallis montium pertinget usque ad Iasol; et fugietis, sicut fugistis a facie terraemotus in diebus Oziae regis Iudae, et veniet Dominus Deus meus, omnesque sancti cum eo.
ZECH|14|6|Erit: in die illa non erit lux sed frigus et gelu;
ZECH|14|7|et erit dies una, quae nota est Domino, non dies neque nox; et in tempore vesperi erit lux.
ZECH|14|8|Et erit: in die illa exibunt aquae vivae de Ierusalem, medium earum ad mare orientale, et medium earum ad mare occidentale: in aestate et in hieme erunt.
ZECH|14|9|Et erit Dominus rex super omnem terram: in die illa erit Dominus unus, et erit nomen eius unum.
ZECH|14|10|Et revertetur omnis terra in desertum, a Gabaa usque ad Remmon ad austrum Ierusalem, quae exaltabitur et habitabitur in loco suo, a porta Beniamin usque ad locum portae Prioris, et usque ad portam Angulorum, et a turre Hananeel usque ad Torcularia regis.
ZECH|14|11|Et habitabunt in ea, et anathema non erit amplius; sed habitabitur Ierusalem secura.
ZECH|14|12|Et haec erit plaga, qua percutiet Dominus omnes gentes, quae pugnaverunt adversus Ierusalem: tabescet caro uniuscuiusque stantis super pedes suos, et oculi eius contabescent in foraminibus suis, et lingua eius contabescet in ore suo.
ZECH|14|13|In die illa erit tumultus Domini magnus in eis, et apprehendet vir manum proximi sui, et elevabitur manus eius super manum proximi sui.
ZECH|14|14|Sed et Iudas pugnabit in Ierusalem, et congregabuntur divitiae omnium gentium in circuitu, aurum et argentum et vestes multae nimis.
ZECH|14|15|Et sic erit ruina equi, muli, cameli et asini et omnium iumentorum, quae fuerint in castris illis, sicut ruina haec.
ZECH|14|16|Et omnes, qui reliqui fuerint de universis gentibus, quae venerunt contra Ierusalem, ascendent ab anno in annum, ut adorent Regem, Dominum exercituum, et celebrent festivitatem Tabernaculorum.
ZECH|14|17|Et erit: qui non ascenderit de familiis terrae ad Ierusalem, ut adoret Regem, Dominum exercituum, non erit super eos imber.
ZECH|14|18|Quod et si familia Aegypti non ascenderit et non venerit, super eos erit plaga, qua percutit Dominus gentes, quae non ascenderint ad celebrandam festivitatem Tabernaculorum.
ZECH|14|19|Haec erit poena Aegypti, et haec poena omnium gentium, quae non ascenderint ad celebrandam festivitatem Tabernaculorum.
ZECH|14|20|In die illa erit super tintinnabula equorum; "Sanctum Domino"; et erunt lebetes in domo Domini quasi phialae coram altari.
ZECH|14|21|Et erit omnis lebes in Ierusalem et in Iuda sanctificatus Domino exercituum; et venient omnes immolantes et sument ex eis et coquent in eis, et non erit mercator ultra in domo Domini exercituum in die illo ".
MAL|1|1|Oraculum. Verbum Domini ad Israel in manu Malachiae.
MAL|1|2|" Dilexi vos, dicit Dominus, et dixistis: "In quo dilexisti nos?". Nonne frater erat Esau Iacob?, dicit Dominus; et dilexi Iacob,
MAL|1|3|Esau autem odio habui et posui montes eius in solitudinem et hereditatem eius thoibus deserti.
MAL|1|4|Quod si dixerit Edom: "Destructi sumus, sed revertentes aedificabimus, quae destructa sunt", haec dicit Dominus exercituum: Isti aedificabunt, et ego destruam; et vocabuntur 'Termini impietatis' et 'Populus, cui iratus est Dominus usque in aeternum'.
MAL|1|5|Et oculi vestri videbunt, et vos dicetis: "Magnificatus est Dominus ultra terminos Israel".
MAL|1|6|Filius honorat patrem, et servus dominum suum. Si ergo pater ego sum, ubi est honor meus? Et si Dominus ego sum, ubi est timor meus?, dicit Dominus exercituum ad vos, o sacerdotes, qui despicitis nomen meum et dicitis: "In quo despeximus nomen tuum?".
MAL|1|7|Offertis super altare meum panem pollutum et dicitis: "In quo polluimus te?". In eo quod dicitis: "Mensa Domini contemptibilis est".
MAL|1|8|Si offeratis caecum ad immolandum, nonne malum est? Et si offeratis claudum et languidum, nonne malum est? Offer illud duci tuo, si placuerit ei, aut si susceperit faciem tuam!, dicit Dominus exercituum.
MAL|1|9|Sed nunc deprecamini vultum Dei, ut misereatur vestri! De manu enim vestra factum est hoc. Num suscipiet facies vestras?, dicit Dominus exercituum.
MAL|1|10|Quis est in vobis, qui claudat ostia, ne incendatis altare meum gratuito? Non est mihi voluntas in vobis, dicit Dominus exercituum; et munus non suscipiam de manu vestra.
MAL|1|11|Ab ortu enim solis usque ad occasum magnum est nomen meum in gentibus, et in omni loco sacrificatur et offertur nomini meo oblatio munda, quia magnum nomen meum in gentibus, dicit Dominus exercituum.
MAL|1|12|Vos autem polluistis illud in eo quod dicitis: "Mensa Domini contaminata est, et contemptibilis esca eius".
MAL|1|13|Et dicitis: "Quantus labor!", et despicitis illam, dicit Dominus exercituum. Et infertis de rapinis claudum et languidum et infertis sicut munus. Numquid suscipiam illud de manu vestra?, dicit Dominus.
MAL|1|14|Maledictus dolosus, qui habet in grege suo masculum et votum faciens immolat debile Domino. Quia Rex magnus ego, dicit Dominus exercituum, et nomen meum horribile in gentibus.
MAL|2|1|Et nunc ad vos mandatum hoc, o sacerdotes.
MAL|2|2|Si nolueritis audi re et si nolueritis ponere super cor, ut detis gloriam nomini meo, ait Dominus exercituum, mittam in vos maledictionem et maledicam benedictionibus vestris; et maledicam illis, quoniam non posuistis super cor.
MAL|2|3|Ecce ego abscindam vobis brachiumet dispergam stercus super vultum vestrum,stercus sollemnitatum vestrarum,et assumet vos secum;
MAL|2|4|et scietis quia misi ad vos mandatum istud,ut esset pactum meum cum Levi,dicit Dominus exercituum.
MAL|2|5|Pactum meum fuit cum eo vitae et pacis,et dedi haec ei simul cum timore, et timuit meet a facie nominis mei pavebat.
MAL|2|6|Lex veritatis fuit in ore eius,et iniquitas non est inventa in labiis eius;in pace et in aequitate ambulavit mecumet multos avertit ab iniquitate.
MAL|2|7|Labia enim sacerdotis custodiunt scientiam,et legem requirunt ex ore eius,quia angelus Domini exercituum est.
MAL|2|8|Vos autem recessistis de viaet scandalizastis plurimos in lege;irritum fecistis pactum Levi,dicit Dominus exercituum;
MAL|2|9|propter quod et ego dedi voscontemptibiles et humiles omnibus populis,sicut non servastis vias measet accepistis personam in lege.
MAL|2|10|Numquid non pater unus omnium nostrum? Numquid non Deus unus creavit nos? Quare ergo dolum facit unusquisque nostrum cum fratre suo, violans pactum patrum nostrorum?
MAL|2|11|Dolum fecit Iuda, et abominatio facta est in Israel et in Ierusalem, quia contaminavit Iuda sanctuarium Domini, quod diligit, et accepit uxorem filiam dei alieni.
MAL|2|12|Disperdet Dominus virum, qui fecerit hoc, filium et nepotem, de tabernaculis Iacob et de offerentibus munus Domino exercituum.
MAL|2|13|Et hoc rursum facitis: operitis lacrimis altare Domini, fletu et mugitu, ita ut non respiciam ultra ad sacrificium nec accipiam placabile quid de manu vestra;
MAL|2|14|et dicitis: "Quam ob causam?". Quia Dominus testificatus est inter te et uxorem adulescentiae tuae, cui tu factus es infidelis; et haec particeps tua et uxor foederis tui.
MAL|2|15|Nonne unitatem fecit carnis et spiritus? Et quid unitas quaerit nisi semen a Deo? Custodite ergo spiritum vestrum; et uxori adulescentiae tuae noli esse infidelis.
MAL|2|16|Si quis odio dimittit, dicit Dominus, Deus Israel, operit iniquitas vestimentum eius, dicit Dominus exercituum. Custodite spiritum vestrum et nolite esse infideles.
MAL|2|17|Laborare facitis Dominum in sermonibus vestris et dicitis: "In quo eum facimus laborare?". In eo quod dicitis: "Omnis, qui facit malum, bonus est in conspectu Domini, et tales ei placent" aut: "Ubi est Deus iudicii?".
MAL|3|1|Ecce ego mittam angelum meum, et praeparabit viam an te faciem meam; et statim veniet ad templum suum Dominator, quem vos quaeritis, et angelus testamenti, quem vos vultis. Ecce venit, dicit Dominus exercituum;
MAL|3|2|et quis poterit sustinere diem adventus eius, et quis stabit, cum apparebit? Ipse enim quasi ignis conflans et quasi herba fullonum;
MAL|3|3|et sedebit conflans et emundans argentum et purgabit filios Levi et colabit eos quasi aurum et quasi argentum, et erunt Domino offerentes sacrificia in iustitia.
MAL|3|4|Et placebit Domino sacrificium Iudae et Ierusalem sicut diebus pristinis et sicut annis antiquis.
MAL|3|5|Et accedam ad vos in iudicio; et ero testis velox maleficis et adulteris et periuris et, qui opprimunt mercennarios, viduas et pupillos et flectunt ius peregrinorum nec timuerunt me, dicit Dominus exercituum.
MAL|3|6|Ego enim Dominus et non mutatus sum;sed vos, filii lacob, nondum ad finem pervenistis.
MAL|3|7|A diebus enim patrum vestrorumrecessistis a praeceptis legitimis meis et non custodistis ea.Revertimini ad me,et revertar ad vos,dicit Dominus exercituum.Et dicitis: "In quo revertemur?".
MAL|3|8|Numquid homo potest defraudare Deum?Sed vos defraudatis me.Et dicitis: "In quo defraudavimus te?".In decimis et in primitiis.
MAL|3|9|Maledictione vos maledicti estis,quia me vos defraudatis, gens tota.
MAL|3|10|Inferte omnem decimam in horreum,et sit cibus in domo mea;et probate me super hoc,dicit Dominus exercituum:si non aperuero vobis cataractas caeliet effudero vobis benedictionem usque ad abundantiam
MAL|3|11|et increpabo pro vobis devorantem,et non corrumpet fructum terrae,nec erit sterilis vobis vinea in agro,dicit Dominus exercituum.
MAL|3|12|Et beatos vos dicent omnes gentes;eritis enim vos terra desiderabilis,dicit Dominus exercituum.
MAL|3|13|Invaluerunt super me verba vestra, dicit Dominus;
MAL|3|14|et dicitis: "Quid locuti sumus contra te?". Dicitis: "Vanum est servire Deo; et, quod emolumentum, quia custodivimus praecepta eius et quia ambulavimus tristes coram Domino exercituum?
MAL|3|15|Ergo nunc beatos dicimus arrogantes; siquidem aedificati sunt facientes impietatem et tentaverunt Deum et salvi facti sunt".
MAL|3|16|Tunc locuti sunt timentes Dominum, unusquisque cum proximo suo. Et attendit Dominus et audivit; et scriptus est liber memorabilium coram eo timentibus Dominum et cogitantibus nomen eius.
MAL|3|17|Erunt mihi, ait Dominus exercituum, in die, qua ego facio in peculium; et parcam eis, sicut parcit vir filio suo servienti sibi.
MAL|4|1|Rursum videbitis quid sit inter iustum et impium, inter servientem Deo et non servientem ei.
MAL|4|2|Ecce enim dies veniet succensa quasi caminus; et erunt omnes superbi et omnes facientes impietatem stipula; et inflammabit eos dies veniens, dicit Dominus exercituum, quae non derelinquet eis radicem et ramum.
MAL|4|3|Et orietur vobis timentibus nomen meum sol iustitiae et sanitas in pennis eius; et egrediemini et salietis sicut vituli saginati
MAL|4|4|et calcabitis impios, cum fuerint cinis sub planta pedum vestrorum in die, quam ego facio, dicit Dominus exercituum.
MAL|4|5|Mementote legis Moysi servi mei,cui mandaviin Horeb ad omnem Israelpraecepta et iudicia.
MAL|4|6|Ecce ego mittam vobisEliam prophetam,antequam veniat dies Dominimagnus et horribilis;
MAL|4|7|et convertet cor patrum ad filioset cor filiorum ad patres eorum,ne veniam et percutiamterram anathemate "
MATT|1|1|Liber generationis Iesu Christi filii David filii Abraham.
MATT|1|2|Abraham genuit Isaac, Isaac autem genuit Iacob, Iacob autem genuit Iudam et fratres eius,
MATT|1|3|Iudas autem genuit Phares et Zara de Thamar, Phares autem genuit Esrom, Esrom autem genuit Aram,
MATT|1|4|Aram autem genuit Aminadab, Aminadab autem genuit Naasson, Naasson autem genuit Salmon,
MATT|1|5|Salmon autem genuit Booz de Rahab, Booz autem genuit Obed ex Ruth, Obed autem genuit Iesse,
MATT|1|6|Iesse autem genuit David regem.David autem genuit Salomonem ex ea, quae fuit Uriae,
MATT|1|7|Salomon autem genuit Roboam, Roboam autem genuit Abiam, Abia autem genuit Asa,
MATT|1|8|Asa autem genuit Iosaphat, Iosaphat autem genuit Ioram, Ioram autem genuit Oziam,
MATT|1|9|Ozias autem genuit Ioatham, Ioatham autem genuit Achaz, Achaz autem genuit Ezechiam,
MATT|1|10|Ezechias autem genuit Manassen, Manasses autem genuit Amon, Amon autem genuit Iosiam,
MATT|1|11|Iosias autem genuit Iechoniam et fratres eius in transmigratione Babylonis.
MATT|1|12|Et post transmigrationem Babylonis Iechonias genuit Salathiel, Salathiel autem genuit Zorobabel,
MATT|1|13|Zorobabel autem genuit Abiud, Abiud autem genuit Eliachim, Eliachim autem genuit Azor,
MATT|1|14|Azor autem genuit Sadoc, Sadoc autem genuit Achim, Achim autem genuit Eliud,
MATT|1|15|Eliud autem genuit Eleazar, Eleazar autem genuit Matthan, Matthan autem genuit Iacob,
MATT|1|16|Iacob autem genuit Ioseph virum Mariae, de qua natus est Iesus, qui vocatur Christus.
MATT|1|17|Omnes ergo generationes ab Abraham usque ad David generationes quattuordecim; et a David usque ad transmigrationem Babylonis generationes quattuordecim; et a transmigratione Babylonis usque ad Christum generationes quattuordecim.
MATT|1|18|Iesu Christi autem generatio sic erat.Cum esset desponsata mater eius Maria Ioseph, antequam convenirent inventa est in utero habens de Spiritu Sancto.
MATT|1|19|Ioseph autem vir eius, cum esset iustus et nollet eam traducere, voluit occulte dimittere eam.
MATT|1|20|Haec autem eo cogitante, ecce angelus Domini in somnis apparuit ei dicens: " Ioseph fili David, noli timere accipere Mariam coniugem tuam. Quod enim in ea natum est, de Spiritu Sancto est;
MATT|1|21|pariet autem filium, et vocabis nomen eius Iesum: ipse enim salvum faciet populum suum a peccatis eorum ".
MATT|1|22|Hoc autem totum factum est, ut adimpleretur id, quod dictum est a Domino per prophetam dicentem:
MATT|1|23|" Ecce, virgo in utero habebit et pariet filium, et vocabunt nomen eius Emmanuel ", quod est interpretatum Nobiscum Deus.
MATT|1|24|Exsurgens autem Ioseph a somno fecit, sicut praecepit ei angelus Domini, et accepit coniugem suam;
MATT|1|25|et non cognoscebat eam, donec peperit filium, et vocavit nomen eius Iesum.
MATT|2|1|Cum autem natus esset Iesus in Bethlehem Iudaeae in diebus Herodis regis, ecce Magi ab oriente venerunt Hierosolymam
MATT|2|2|dicentes: " Ubi est, qui natus est, rex Iudaeorum? Vidimus enim stellam eius in oriente et venimus adorare eum ".
MATT|2|3|Audiens autem Herodes rex turbatus est et omnis Hierosolyma cum illo;
MATT|2|4|et congregans omnes principes sacerdotum et scribas populi, sciscitabatur ab eis ubi Christus nasceretur.
MATT|2|5|At illi dixerunt ei: " In Bethlehem Iudaeae. Sic enim scriptum est per prophetam:
MATT|2|6|"Et tu, Bethlehem terra Iudae,nequaquam minima es in principibus Iudae;ex te enim exiet dux,qui reget populum meum Israel" ".
MATT|2|7|Tunc Herodes, clam vocatis Magis, diligenter didicit ab eis tempus stellae, quae apparuit eis;
MATT|2|8|et mittens illos in Bethlehem dixit: " Ite et interrogate diligenter de puero; et cum inveneritis, renuntiate mihi, ut et ego veniens adorem eum.
MATT|2|9|Qui cum audissent regem, abierunt. Et ecce stella, quam viderant in oriente, antecedebat eos, usque dum veniens staret supra, ubi erat puer.
MATT|2|10|Videntes autem stellam gavisi sunt gaudio magno valde.
MATT|2|11|Et intrantes domum viderunt puerum cum Maria matre eius, et procidentes adoraverunt eum; et apertis thesauris suis, obtulerunt ei munera, aurum et tus et myrrham.
MATT|2|12|Et responso accepto in somnis, ne redirent ad Herodem, per aliam viam reversi sunt in regionem suam.
MATT|2|13|Qui cum recessissent, ecce angelus Domini apparet in somnis Ioseph dicens: " Surge et accipe puerum et matrem eius et fuge in Aegyptum et esto ibi, usque dum dicam tibi; futurum est enim ut Herodes quaerat puerum ad perdendum eum ".
MATT|2|14|Qui consurgens accepit puerum et matrem eius nocte et recessit in Aegyptum
MATT|2|15|et erat ibi usque ad obitum Herodis, ut adimpleretur, quod dictum est a Domino per prophetam dicentem: Ex Aegypto vocavi filium meum ".
MATT|2|16|Tunc Herodes videns quoniam illusus esset a Magis, iratus est valde et mittens occidit omnes pueros, qui erant in Bethlehem et in omnibus finibus eius, a bimatu et infra, secundum tempus, quod exquisierat a Magis.
MATT|2|17|Tunc adimpletum est, quod dictum est per Ieremiam prophetam dicentem:
MATT|2|18|" Vox in Rama audita est,ploratus et ululatus multus:Rachel plorans filios suos,et noluit consolari, quia non sunt ".
MATT|2|19|Defuncto autem Herode, ecce apparet angelus Domini in somnis Ioseph in Aegypto
MATT|2|20|dicens: " Surge et accipe puerum et matrem eius et vade in terram Israel; defuncti sunt enim, qui quaerebant animam pueri ".
MATT|2|21|Qui surgens accepit puerum et matrem eius et venit in terram Israel.
MATT|2|22|Audiens autem quia Archelaus regnaret in Iudaea pro Herode patre suo, timuit illuc ire; et admonitus in somnis, secessit in partes Galilaeae
MATT|2|23|et veniens habitavit in civitate, quae vocatur Nazareth, ut adimpleretur, quod dictum est per Prophetas: " Nazaraeus vocabitur ".
MATT|3|1|In diebus autem illis venit Ioannes Baptista praedicans in deserto Iudaeae
MATT|3|2|et dicens: " Paenitentiam agite; appropinquavit enim regnum caelorum ".
MATT|3|3|Hic est enim, qui dictus est per Isaiam prophetam dicentem: Vox clamantis in deserto:Parate viam Domini,rectas facite semitas eius!" ".
MATT|3|4|Ipse autem Ioannes habebat vestimentum de pilis cameli et zonam pelliceam circa lumbos suos; esca autem eius erat locustae et mel silvestre.
MATT|3|5|Tunc exibat ad eum Hierosolyma et omnis Iudaea et omnis regio circa Iordanem,
MATT|3|6|et baptizabantur in Iordane flumine ab eo, confitentes peccata sua.
MATT|3|7|Videns autem multos pharisaeorum et sadducaeorum venientes ad baptismum suum, dixit eis: " Progenies viperarum, quis demonstravit vobis fugere a futura ira?
MATT|3|8|Facite ergo fructum dignum paenitentiae
MATT|3|9|et ne velitis dicere intra vos: "Patrem habemus Abraham"; dico enim vobis quoniam potest Deus de lapidibus istis suscitare Abrahae filios.
MATT|3|10|Iam enim securis ad radicem arborum posita est; omnis ergo arbor, quae non facit fructum bonum, exciditur et in ignem mittitur.
MATT|3|11|Ego quidem vos baptizo in aqua in paenitentiam; qui autem post me venturus est, fortior me est, cuius non sum dignus calceamenta portare; ipse vos baptizabit in Spiritu Sancto et igni,
MATT|3|12|cuius ventilabrum in manu sua, et permundabit aream suam et congregabit triticum suum in horreum, paleas autem comburet igni inexstinguibili ".
MATT|3|13|Tunc venit Iesus a Galilaea in Iordanem ad Ioannem, ut baptizaretur ab eo.
MATT|3|14|Ioannes autem prohibebat eum dicens: " Ego a te debeo baptizari, et tu venis ad me? ".
MATT|3|15|Respondens autem Iesus dixit ei: " Sine modo, sic enim decet nos implere omnem iustitiam ". Tunc dimittit eum.
MATT|3|16|Baptizatus autem Iesus, confestim ascendit de aqua; et ecce aperti sunt ei caeli, et vidit Spiritum Dei descendentem sicut columbam et venientem super se.
MATT|3|17|Et ecce vox de caelis dicens: "Hic est Filius meus dilectus, in quomihi complacui ".
MATT|4|1|Tunc Iesus ductus est in de sertum a Spiritu, ut tentaretur a Diabolo.
MATT|4|2|Et cum ieiunasset quadraginta diebus et quadraginta noctibus, postea esuriit.
MATT|4|3|Et accedens tentator dixit ei: " Si Filius Dei es, dic, ut lapides isti panes fiant ".
MATT|4|4|Qui respondens dixit: Scriptum est:Non in pane solo vivet homo,sed in omni verbo, quod procedit de ore Dei" ".
MATT|4|5|Tunc assumit eum Diabolus in sanctam civitatem et statuit eum supra pinnaculum templi
MATT|4|6|et dicit ei: " Si Filius Dei es, mitte te deorsum. Scriptum est enim:Angelis suis mandabit de te,et in manibus tollent te,ne forte offendas ad lapidem pedem tuum" ".
MATT|4|7|Ait illi Iesus: " Rursum scriptum est: "Non tentabis Dominum Deum tuum".
MATT|4|8|Iterum assumit eum Diabolus in montem excelsum valde et ostendit ei omnia regna mundi et gloriam eorum
MATT|4|9|et dicit illi: " Haec tibi omnia dabo, si cadens adoraveris me".
MATT|4|10|Tunc dicit ei Iesus: Vade, Satanas! Scriptum est enim:Dominum Deum tuum adorabiset illi soli servies" ".
MATT|4|11|Tunc reliquit eum Diabolus, et ecce angeli accesserunt et ministrabant ei.
MATT|4|12|Cum autem audisset quod Ioannes traditus esset, secessit in Galilaeam.
MATT|4|13|Et relicta Nazareth, venit et habitavit in Capharnaum maritimam
MATT|4|14|in finibus Zabulon et Nephthali, ut impleretur, quod dictum est per Isaiam prophetam dicentem:
MATT|4|15|" Terra Zabulon et terra Nephthali,ad viam maris, trans Iordanem,Galilaea gentium;
MATT|4|16|populus, qui sedebat in tenebris,lucem vidit magnam,et sedentibus in regione et umbra mortislux orta est eis ".
MATT|4|17|Exinde coepit Iesus praedicare et dicere: " Paenitentiam agite; appropinquavit enim regnum caelorum ".
MATT|4|18|Ambulans autem iuxta mare Galilaeae, vidit duos fratres, Simonem, qui vocatur Petrus, et Andream fratrem eius, mittentes rete in mare; erant enim piscatores.
MATT|4|19|Et ait illis: " Venite post me, et faciam vos piscatores hominum ".
MATT|4|20|At illi continuo, relictis retibus, secuti sunt eum.
MATT|4|21|Et procedens inde vidit alios duos fratres, Iacobum Zebedaei et Ioannem fratrem eius, in navi cum Zebedaeo patre eorum reficientes retia sua; et vocavit eos.
MATT|4|22|Illi autem statim, relicta navi et patre suo, secuti sunt eum.
MATT|4|23|Et circumibat Iesus totam Galilaeam, docens in synagogis eorum et praedicans evangelium regni et sanans omnem languorem et omnem infirmitatem in populo.
MATT|4|24|Et abiit opinio eius in totam Syriam; et obtulerunt ei omnes male habentes, variis languoribus et tormentis comprehensos, et qui daemonia habebant, et lunaticos et paralyticos, et curavit eos.
MATT|4|25|Et secutae sunt eum turbae multae de Galilaea et Decapoli et Hierosolymis et Iudaea et de trans Iordanem.
MATT|5|1|Videns autem turbas, ascendit in montem; et cum sedisset, ac cesserunt ad eum discipuli eius;
MATT|5|2|et aperiens os suum docebat eos dicens:
MATT|5|3|" Beati pauperes spiritu, quoniam ipsorum est regnum caelorum.
MATT|5|4|Beati, qui lugent, quoniam ipsi consolabuntur.
MATT|5|5|Beati mites, quoniam ipsi possidebunt terram.
MATT|5|6|Beati, qui esuriunt et sitiunt iustitiam, quoniam ipsi saturabuntur.
MATT|5|7|Beati misericordes, quia ipsi misericordiam consequentur.
MATT|5|8|Beati mundo corde, quoniam ipsi Deum videbunt.
MATT|5|9|Beati pacifici, quoniam filii Dei vocabuntur.
MATT|5|10|Beati, qui persecutionem patiuntur propter iustitiam, quoniam ipsorum est regnum caelorum.
MATT|5|11|Beati estis cum maledixerint vobis et persecuti vos fuerint et dixerint omne malum adversum vos, mentientes, propter me.
MATT|5|12|Gaudete et exsultate, quoniam merces vestra copiosa est in caelis; sic enim persecuti sunt prophetas, qui fuerunt ante vos.
MATT|5|13|Vos estis sal terrae; quod si sal evanuerit, in quo salietur? Ad nihilum valet ultra, nisi ut mittatur foras et conculcetur ab hominibus.
MATT|5|14|Vos estis lux mundi. Non potest civitas abscondi supra montem posita;
MATT|5|15|neque accendunt lucernam et ponunt eam sub modio, sed super candelabrum, ut luceat omnibus, qui in domo sunt.
MATT|5|16|Sic luceat lux vestra coram hominibus, ut videant vestra bona opera et glorificent Patrem vestrum, qui in caelis est.
MATT|5|17|Nolite putare quoniam veni solvere Legem aut Prophetas; non veni solvere, sed adimplere.
MATT|5|18|Amen quippe dico vobis: Donec transeat caelum et terra, iota unum aut unus apex non praeteribit a Lege, donec omnia fiant.
MATT|5|19|Qui ergo solverit unum de mandatis istis minimis et docuerit sic homines, minimus vocabitur in regno caelorum; qui autem fecerit et docuerit, hic magnus vocabitur in regno caelorum.
MATT|5|20|Dico enim vobis: Nisi abundaverit iustitia vestra plus quam scribarum et pharisaeorum, non intrabitis in regnum caelorum.
MATT|5|21|Audistis quia dictum est antiquis: "Non occides; qui autem occiderit, reus erit iudicio".
MATT|5|22|Ego autem dico vobis: Omnis, qui irascitur fratri suo, reus erit iudicio; qui autem dixerit fratri suo: "Racha", reus erit concilio; qui autem dixerit: "Fatue", reus erit gehennae ignis.
MATT|5|23|Si ergo offeres munus tuum ad altare, et ibi recordatus fueris quia frater tuus habet aliquid adversum te,
MATT|5|24|relinque ibi munus tuum ante altare et vade, prius, reconciliare fratri tuo et tunc veniens offer munus tuum.
MATT|5|25|Esto consentiens adversario tuo cito, dum es in via cum eo, ne forte tradat te adversarius iudici, et iudex tradat te ministro, et in carcerem mittaris.
MATT|5|26|Amen dico tibi: Non exies inde, donec reddas novissimum quadrantem.
MATT|5|27|Audistis quia dictum est: "Non moechaberis".
MATT|5|28|Ego autem dico vobis: Omnis, qui viderit mulierem ad concupiscendum eam, iam moechatus est eam in corde suo.
MATT|5|29|Quod si oculus tuus dexter scandalizat te, erue eum et proice abs te; expedit enim tibi, ut pereat unum membrorum tuorum, quam totum corpus tuum mittatur in gehennam.
MATT|5|30|Et si dextera manus tua scandalizat te, abscide eam et proice abs te; expedit enim tibi, ut pereat unum membrorum tuorum, quam totum corpus tuum abeat in gehennam.
MATT|5|31|Dictum est autem: "Quicumque dimiserit uxorem suam, det illi libellum repudii".
MATT|5|32|Ego autem dico vobis: Omnis, qui dimiserit uxorem suam, excepta fornicationis causa, facit eam moechari; et, qui dimissam duxerit, adulterat.
MATT|5|33|Iterum audistis quia dictum est antiquis: "Non periurabis; reddes autem Domino iuramenta tua".
MATT|5|34|Ego autem dico vobis: Non iurare omnino, neque per caelum, quia thronus Dei est,
MATT|5|35|neque per terram, quia scabellum est pedum eius, neque per Hierosolymam, quia civitas est magni Regis;
MATT|5|36|neque per caput tuum iuraveris, quia non potes unum capillum album facere aut nigrum.
MATT|5|37|Sit autem sermo vester: "Est, est", "Non, non"; quod autem his abundantius est, a Malo est.
MATT|5|38|Audistis quia dictum est: "Oculum pro oculo et dentem pro dente".
MATT|5|39|Ego autem dico vobis: Non resistere malo; sed si quis te percusserit in dextera maxilla tua, praebe illi et alteram;
MATT|5|40|et ei, qui vult tecum iudicio contendere et tunicam tuam tollere, remitte ei et pallium;
MATT|5|41|et quicumque te angariaverit mille passus, vade cum illo duo.
MATT|5|42|Qui petit a te, da ei; et volenti mutuari a te, ne avertaris.
MATT|5|43|Audistis quia dictum est: "Diliges proximum tuum et odio habebis inimicum tuum".
MATT|5|44|Ego autem dico vobis: Diligite inimicos vestros et orate pro persequentibus vos,
MATT|5|45|ut sitis filii Patris vestri, qui in caelis est, quia solem suum oriri facit super malos et bonos et pluit super iustos et iniustos.
MATT|5|46|Si enim dilexeritis eos, qui vos diligunt, quam mercedem habetis? Nonne et publicani hoc faciunt?
MATT|5|47|Et si salutaveritis fratres vestros tantum, quid amplius facitis? Nonne et ethnici hoc faciunt?
MATT|5|48|Estote ergo vos perfecti, sicut Pater vester caelestis perfectus est.
MATT|6|1|Attendite, ne iustitiam vestram faciatis coram hominibus, ut vi deamini ab eis; alioquin mercedem non habetis apud Patrem vestrum, qui in caelis est.
MATT|6|2|Cum ergo facies eleemosynam, noli tuba canere ante te, sicut hypocritae faciunt in synagogis et in vicis, ut honorificentur ab hominibus. Amen dico vobis: Receperunt mercedem suam.
MATT|6|3|Te autem faciente eleemosynam, nesciat sinistra tua quid faciat dextera tua,
MATT|6|4|ut sit eleemosyna tua in abscondito, et Pater tuus, qui videt in abscondito, reddet tibi.
MATT|6|5|Et cum oratis, non eritis sicut hypocritae, qui amant in synagogis et in angulis platearum stantes orare, ut videantur ab hominibus. Amen dico vobis: Receperunt mercedem suam.
MATT|6|6|Tu autem cum orabis, intra in cubiculum tuum et, clauso ostio tuo, ora Patrem tuum, qui est in abscondito; et Pater tuus, qui videt in abscondito, reddet tibi.
MATT|6|7|Orantes autem nolite multum loqui sicut ethnici; putant enim quia in multiloquio suo exaudiantur.
MATT|6|8|Nolite ergo assimilari eis; scit enim Pater vester, quibus opus sit vobis, antequam petatis eum.
MATT|6|9|Sic ergo vos orabitis:Pater noster, qui es in caelis,sanctificetur nomen tuum,
MATT|6|10|adveniat regnum tuum,fiat voluntas tua,sicut in caelo, et in terra.
MATT|6|11|Panem nostrum supersubstantialem da nobis hodie;
MATT|6|12|et dimitte nobis debita nostra,sicut et nos dimittimus debitoribus nostris;
MATT|6|13|et ne inducas nos in tentationem,sed libera nos a Malo.
MATT|6|14|Si enim dimiseritis hominibus peccata eorum, dimittet et vobis Pater vester caelestis;
MATT|6|15|si autem non dimiseritis hominibus, nec Pater vester dimittet peccata vestra.
MATT|6|16|Cum autem ieiunatis, nolite fieri sicut hypocritae tristes; demoliuntur enim facies suas, ut pareant hominibus ieiunantes. Amen dico vobis: Receperunt mercedem suam.
MATT|6|17|Tu autem cum ieiunas, unge caput tuum et faciem tuam lava,
MATT|6|18|ne videaris hominibus ieiunans sed Patri tuo, qui est in abscondito; et Pater tuus, qui videt in abscondito, reddet tibi.
MATT|6|19|Nolite thesaurizare vobis thesauros in terra, ubi aerugo et tinea demolitur, et ubi fures effodiunt et furantur;
MATT|6|20|thesaurizate autem vobis thesauros in caelo, ubi neque aerugo neque tinea demolitur, et ubi fures non effodiunt nec furantur;
MATT|6|21|ubi enim est thesaurus tuus, ibi erit et cor tuum.
MATT|6|22|Lucerna corporis est oculus. Si ergo fuerit oculus tuus simplex, totum corpus tuum lucidum erit;
MATT|6|23|si autem oculus tuus nequam fuerit, totum corpus tuum tenebrosum erit. Si ergo lumen, quod in te est, tene brae sunt, tenebrae quantae erunt!
MATT|6|24|Nemo potest duobus dominis servire: aut enim unum odio habebit et alterum diliget, aut unum sustinebit et alterum contemnet; non potestis Deo servire et mammonae.
MATT|6|25|Ideo dico vobis: Ne solliciti sitis animae vestrae quid manducetis, neque corpori vestro quid induamini. Nonne anima plus est quam esca, et corpus quam vestimentum?
MATT|6|26|Respicite volatilia caeli, quoniam non serunt neque metunt neque congregant in horrea, et Pater vester caelestis pascit illa. Nonne vos magis pluris estis illis?
MATT|6|27|Quis autem vestrum cogitans potest adicere ad aetatem suam cubitum unum?
MATT|6|28|Et de vestimento quid solliciti estis? Considerate lilia agri quomodo crescunt: non laborant neque nent.
MATT|6|29|Dico autem vobis quoniam nec Salomon in omni gloria sua coopertus est sicut unum ex istis.
MATT|6|30|Si autem fenum agri, quod hodie est et cras in clibanum mittitur, Deus sic vestit, quanto magis vos, modicae fidei?
MATT|6|31|Nolite ergo solliciti esse dicentes: "Quid manducabimus?", aut: "Quid bibemus?", aut: "Quo operiemur?".
MATT|6|32|Haec enim omnia gentes inquirunt; scit enim Pater vester caelestis quia his omnibus indigetis.
MATT|6|33|Quaerite autem primum regnum Dei et iustitiam eius, et haec omnia adicientur vobis.
MATT|6|34|Nolite ergo esse solliciti in crastinum; crastinus enim dies sollicitus erit sibi ipse. Sufficit diei malitia sua.
MATT|7|1|Nolite iudicare, ut non iudice mini;
MATT|7|2|in quo enim iudicio iudi caveritis, iudicabimini, et in qua mensura mensi fueritis, metietur vobis.
MATT|7|3|Quid autem vides festucam in oculo fratris tui, et trabem in oculo tuo non vides?
MATT|7|4|Aut quomodo dices fratri tuo: "Sine, eiciam festucam de oculo tuo", et ecce trabes est in oculo tuo?
MATT|7|5|Hypocrita, eice primum trabem de oculo tuo, et tunc videbis eicere festucam de oculo fratris tui.
MATT|7|6|Nolite dare sanctum canibus neque mittatis margaritas vestras ante porcos, ne forte conculcent eas pedibus suis et conversi dirumpant vos.
MATT|7|7|Petite, et dabitur vobis; quaerite et invenietis; pulsate, et aperietur vobis.
MATT|7|8|Omnis enim qui petit, accipit; et, qui quaerit, invenit; et pulsanti aperietur.
MATT|7|9|Aut quis est ex vobis homo, quem si petierit filius suus panem, numquid lapidem porriget ei?
MATT|7|10|Aut si piscem petierit, numquid serpentem porriget ei?
MATT|7|11|Si ergo vos, cum sitis mali, nostis dona bona dare filiis vestris, quanto magis Pater vester, qui in caelis est, dabit bona petentibus se.
MATT|7|12|Omnia ergo, quaecumque vultis ut faciant vobis homines, ita et vos facite eis; haec est enim Lex et Prophetae.
MATT|7|13|Intrate per angustam portam, quia lata porta et spatiosa via, quae ducit ad perditionem, et multi sunt, qui intrant per eam;
MATT|7|14|quam angusta porta et arta via, quae ducit ad vitam, et pauci sunt, qui inveniunt eam!
MATT|7|15|Attendite a falsis prophetis, qui veniunt ad vos in vestimentis ovium, intrinsecus autem sunt lupi rapaces.
MATT|7|16|A fructibus eorum cognoscetis eos; numquid colligunt de spinis uvas aut de tribulis ficus?
MATT|7|17|Sic omnis arbor bona fructus bonos facit, mala autem arbor fructus malos facit;
MATT|7|18|non potest arbor bona fructus malos facere, neque arbor mala fructus bonos facere.
MATT|7|19|Omnis arbor, quae non facit fructum bonum, exciditur et in ignem mittitur.
MATT|7|20|Igitur ex fructibus eorum cognoscetis eos.
MATT|7|21|Non omnis, qui dicit mihi: "Domine, Domine", intrabit in regnum caelorum, sed qui facit voluntatem Patris mei, qui in caelis est.
MATT|7|22|Multi dicent mihi in illa die: "Domine, Domine, nonne in tuo nomine prophetavimus, et in tuo nomine daemonia eiecimus, et in tuo nomine virtutes multas fecimus?".
MATT|7|23|Et tunc confitebor illis: Numquam novi vos; discedite a me, qui operamini iniquitatem.
MATT|7|24|Omnis ergo, qui audit verba mea haec et facit ea, assimilabitur viro sapienti, qui aedificavit domum suam supra petram.
MATT|7|25|Et descendit pluvia, et venerunt flumina, et flaverunt venti et irruerunt in domum illam, et non cecidit; fundata enim erat supra petram.
MATT|7|26|Et omnis, qui audit verba mea haec et non facit ea, similis erit viro stulto, qui aedificavit domum suam supra arenam.
MATT|7|27|Et descendit pluvia, et venerunt flumina, et flaverunt venti et irruerunt in domum illam, et cecidit, et fuit ruina eius magna ".
MATT|7|28|Et factum est, cum consummasset Iesus verba haec, admirabantur turbae super doctrinam eius;
MATT|7|29|erat enim docens eos sicut potestatem habens, et non sicut scribae eorum.
MATT|8|1|Cum autem descendisset de monte, secutae sunt eum turbae multae.
MATT|8|2|Et ecce leprosus veniens adorabat eum dicens: " Domine, si vis, potes me mundare ".
MATT|8|3|Et extendens manum, tetigit eum dicens: " Volo, mundare! "; et confestim mundata est lepra eius.
MATT|8|4|Et ait illi Iesus: " Vide, nemini dixeris; sed vade, ostende te sacerdoti et offer munus, quod praecepit Moyses, in testimonium illis ".
MATT|8|5|Cum autem introisset Capharnaum, accessit ad eum centurio rogans eum
MATT|8|6|et dicens: " Domine, puer meus iacet in domo paralyticus et male torquetur ".
MATT|8|7|Et ait illi: " Ego veniam et curabo eum ".
MATT|8|8|Et respondens centurio ait: " Domine, non sum dignus, ut intres sub tectum meum, sed tantum dic verbo, et sanabitur puer meus.
MATT|8|9|Nam et ego homo sum sub potestate, habens sub me milites, et dico huic: Vade", et vadit; et alii: "Veni", et venit; et servo meo: "Fac hoc", et facit".
MATT|8|10|Audiens autem Iesus, miratus est et sequentibus se dixit: "Amen dico vobis: Apud nullum inveni tantam fidem in Israel!
MATT|8|11|Dico autem vobis quod multi ab oriente et occidente venient et recumbent cum Abraham et Isaac et Iacob in regno caelorum;
MATT|8|12|filii autem regni eicientur in tenebras exteriores: ibi erit fletus et stridor dentium ".
MATT|8|13|Et dixit Iesus centurioni: " Vade; sicut credidisti, fiat tibi ". Et sanatus est puer in hora illa.
MATT|8|14|Et cum venisset Iesus in domum Petri, vidit socrum eius iacentem et febricitantem;
MATT|8|15|et tetigit manum eius, et dimisit eam febris; et surrexit et ministrabat ei.
MATT|8|16|Vespere autem facto, obtulerunt ei multos daemonia habentes; et eiciebat spiritus verbo et omnes male habentes curavit,
MATT|8|17|ut adimpleretur, quod dictum est per Isaiam prophetam dicentem: Ipse infirmitates nostras accepitet aegrotationes portavit ".
MATT|8|18|Videns autem Iesus turbas multas circum se, iussit ire trans fretum.
MATT|8|19|Et accedens unus scriba ait illi: " Magister, sequar te, quocumque ieris ".
MATT|8|20|Et dicit ei Iesus: " Vulpes foveas habent, et volucres caeli tabernacula, Filius autem hominis non habet, ubi caput reclinet ".
MATT|8|21|Alius autem de discipulis eius ait illi: "Domine, permitte me primum ire et sepelire patrem meum ".
MATT|8|22|Iesus autem ait illi: " Sequere me et dimitte mortuos sepelire mortuos suos ".
MATT|8|23|Et ascendente eo in naviculam, secuti sunt eum discipuli eius.
MATT|8|24|Et ecce motus magnus factus est in mari, ita ut navicula operiretur fluctibus; ipse vero dormiebat.
MATT|8|25|Et accesserunt et suscitaverunt eum dicentes: " Domine, salva nos, perimus! ".
MATT|8|26|Et dicit eis: " Quid timidi estis, modicae fidei? ". Tunc surgens increpavit ventis et mari, et facta est tranquillitas magna.
MATT|8|27|Porro homines mirati sunt dicentes: " Qualis est hic, quia et venti et mare oboediunt ei? ".
MATT|8|28|Et cum venisset trans fretum in regionem Gadarenorum, occurrerunt ei duo habentes daemonia, de monumentis exeuntes, saevi nimis, ita ut nemo posset transire per viam illam.
MATT|8|29|Et ecce clamaverunt dicentes: " Quid nobis et tibi, Fili Dei? Venisti huc ante tempus torquere nos? ".
MATT|8|30|Erat autem longe ab illis grex porcorum multorum pascens.
MATT|8|31|Daemones autem rogabant eum dicentes: " Si eicis nos, mitte nos in gregem porcorum ".
MATT|8|32|Et ait illis: " Ite ". Et illi exeuntes abierunt in porcos; et ecce impetu abiit totus grex per praeceps in mare, et mortui sunt in aquis.
MATT|8|33|Pastores autem fugerunt et venientes in civitatem nuntiaverunt omnia et de his, qui daemonia habuerant.
MATT|8|34|Et ecce tota civitas exiit obviam Iesu, et viso eo rogabant, ut transiret a finibus eorum.
MATT|9|1|Et ascendens in naviculam transfretavit et venit in civita tem suam.
MATT|9|2|Et ecce offerebant ei paralyticum iacentem in lecto. Et videns Iesus fidem illorum, dixit paralytico: " Confide, fili; remittuntur peccata tua.
MATT|9|3|Et ecce quidam de scribis dixerunt intra se: " Hic blasphemat ".
MATT|9|4|Et cum vidisset Iesus cogitationes eorum, dixit: " Ut quid cogitatis mala in cordibus vestris?
MATT|9|5|Quid enim est facilius, dicere: "Dimittuntur peccata tua", aut dicere: Surge et ambula"?
MATT|9|6|Ut sciatis autem quoniam Filius hominis habet potestatem in terra dimittendi peccata - tunc ait paralytico -: Surge, tolle lectum tuum et vade in domum tuam ".
MATT|9|7|Et surrexit et abiit in domum suam.
MATT|9|8|Videntes autem turbae timuerunt et glorificaverunt Deum, qui dedit potestatem talem hominibus.
MATT|9|9|Et cum transiret inde Iesus, vidit hominem sedentem in teloneo, Matthaeum nomine, et ait illi: "Sequere me". Et surgens secutus est eum.
MATT|9|10|Et factum est, discumbente eo in domo, ecce multi publicani et peccatores venientes simul discumbebant cum Iesu et discipulis eius.
MATT|9|11|Et videntes pharisaei dicebant discipulis eius: " Quare cum publicanis et peccatoribus manducat magister vester? ".
MATT|9|12|At ille audiens ait: " Non est opus valentibus medico sed male habentibus.
MATT|9|13|Euntes autem discite quid est: "Misericordiam volo et non sacrificium". Non enim veni vocare iustos sed peccatores ".
MATT|9|14|Tunc accedunt ad eum discipuli Ioannis dicentes: " Quare nos et pharisaei ieiunamus frequenter, discipuli autem tui non ieiunant? ".
MATT|9|15|Et ait illis Iesus: " Numquid possunt convivae nuptiarum lugere, quamdiu cum illis est sponsus? Venient autem dies, cum auferetur ab eis sponsus, et tunc ieiunabunt.
MATT|9|16|Nemo autem immittit commissuram panni rudis in vestimentum vetus; tollit enim supplementum eius a vestimento, et peior scissura fit.
MATT|9|17|Neque mittunt vinum novum in utres veteres, alioquin rumpuntur utres, et vinum effunditur, et utres pereunt; sed vinum novum in utres novos mittunt, et ambo conservantur ".
MATT|9|18|Haec illo loquente ad eos, ecce princeps unus accessit et adorabat eum dicens: " Filia mea modo defuncta est; sed veni, impone manum tuam super eam, et vivet ".
MATT|9|19|Et surgens Iesus sequebatur eum et discipuli eius.
MATT|9|20|Et ecce mulier, quae sanguinis fluxum patiebatur duodecim annis, accessit retro et tetigit fimbriam vestimenti eius.
MATT|9|21|Dicebat enim intra se: " Si tetigero tantum vestimentum eius, salva ero.
MATT|9|22|At Iesus conversus et videns eam dixit: " Confide, filia; fides tua te salvam fecit ". Et salva facta est mulier ex illa hora.
MATT|9|23|Et cum venisset Iesus in domum principis et vidisset tibicines et turbam tumultuantem,
MATT|9|24|dicebat: " Recedite; non est enim mortua puella, sed dormit ". Et deridebant eum.
MATT|9|25|At cum eiecta esset turba, intravit et tenuit manum eius, et surrexit puella.
MATT|9|26|Et exiit fama haec in universam terram illam.
MATT|9|27|Et transeunte inde Iesu, secuti sunt eum duo caeci clamantes et dicentes: " Miserere nostri, fili David! ".
MATT|9|28|Cum autem venisset domum, accesserunt ad eum caeci, et dicit eis Iesus: Creditis quia possum hoc facere? ". Dicunt ei: "Utique, Domine".
MATT|9|29|Tunc tetigit oculos eorum dicens: "Secundum fidem vestram fiat vobis".
MATT|9|30|Et aperti sunt oculi illorum. Et comminatus est illis Iesus dicens: " Videte, ne quis sciat ".
MATT|9|31|Illi autem exeuntes diffamaverunt eum in universa terra illa.
MATT|9|32|Egressis autem illis, ecce obtulerunt ei hominem mutum, daemonium habentem.
MATT|9|33|Et eiecto daemone, locutus est mutus. Et miratae sunt turbae dicentes: Numquam apparuit sic in Israel! ".
MATT|9|34|Pharisaei autem dicebant: " In principe daemoniorum eicit daemones ".
MATT|9|35|Et circumibat Iesus civitates omnes et castella, docens in synagogis eorum et praedicans evangelium regni et curans omnem languorem et omnem infirmitatem.
MATT|9|36|Videns autem turbas, misertus est eis, quia erant vexati et iacentes sicut oves non habentes pastorem.
MATT|9|37|Tunc dicit discipulis suis: " Messis quidem multa, operarii autem pauci;
MATT|9|38|rogate ergo Dominum messis, ut mittat operarios in messem suam ".
MATT|10|1|Et convocatis Duodecim di scipulis suis, dedit illis pote statem spirituum immundorum, ut eicerent eos et curarent omnem languorem et omnem infirmitatem.
MATT|10|2|Duodecim autem apostolorum nomina sunt haec: primus Simon, qui dicitur Petrus, et Andreas frater eius, et Iacobus Zebedaei et Ioannes frater eius,
MATT|10|3|Philippus et Bartholomaeus, Thomas et Matthaeus publicanus, Iacobus Alphaei et Thaddaeus,
MATT|10|4|Simon Chananaeus et Iudas Iscariotes, qui et tradidit eum.
MATT|10|5|Hos Duodecim misit Iesus praecipiens eis et dicens: " In viam gentium ne abieritis et in civitates Samaritanorum ne intraveritis;
MATT|10|6|sed potius ite ad oves, quae perierunt domus Israel.
MATT|10|7|Euntes autem praedicate dicentes: "Appropinquavit regnum caelorum".
MATT|10|8|Infirmos curate, mortuos suscitate, leprosos mundate, daemones eicite; gratis accepistis, gratis date.
MATT|10|9|Nolite possidere aurum neque argentum neque pecuniam in zonis vestris,
MATT|10|10|non peram in via neque duas tunicas neque calceamenta neque virgam; dignus enim est operarius cibo suo.
MATT|10|11|In quamcumque civitatem aut castellum intraveritis, interrogate quis in ea dignus sit; et ibi manete donec exeatis.
MATT|10|12|Intrantes autem in domum, salutate eam;
MATT|10|13|et si quidem fuerit domus digna, veniat pax vestra super eam; si autem non fuerit digna, pax vestra ad vos revertatur.
MATT|10|14|Et quicumque non receperit vos neque audierit sermones vestros, exeuntes foras de domo vel de civitate illa, excutite pulverem de pedibus vestris.
MATT|10|15|Amen dico vobis: Tolerabilius erit terrae Sodomorum et Gomorraeorum in die iudicii quam illi civitati.
MATT|10|16|Ecce ego mitto vos sicut oves in medio luporum; estote ergo prudentes sicut serpentes et simplices sicut columbae.
MATT|10|17|Cavete autem ab hominibus; tradent enim vos in conciliis, et in synagogis suis flagellabunt vos;
MATT|10|18|et ad praesides et ad reges ducemini propter me in testimonium illis et gentibus.
MATT|10|19|Cum autem tradent vos, nolite cogitare quomodo aut quid loquamini; dabitur enim vobis in illa hora quid loquamini.
MATT|10|20|Non enim vos estis, qui loquimini, sed Spiritus Patris vestri, qui loquitur in vobis.
MATT|10|21|Tradet autem frater fratrem in mortem, et pater filium; et insurgent filii in parentes et morte eos afficient.
MATT|10|22|Et eritis odio omnibus propter nomen meum; qui autem perseveraverit in finem, hic salvus erit.
MATT|10|23|Cum autem persequentur vos in civitate ista, fugite in aliam; amen enim dico vobis: Non consummabitis civitates Israel, donec veniat Filius hominis.
MATT|10|24|Non est discipulus super magistrum nec servus super dominum suum.
MATT|10|25|Sufficit discipulo, ut sit sicut magister eius, et servus sicut dominus eius. Si patrem familias Beelzebul vocaverunt, quanto magis domesticos eius!
MATT|10|26|Ne ergo timueritis eos. Nihil enim est opertum, quod non revelabitur, et occultum, quod non scietur.
MATT|10|27|Quod dico vobis in tenebris, dicite in lumine; et, quod in aure auditis, praedicate super tecta.
MATT|10|28|Et nolite timere eos, qui occidunt corpus, animam autem non possunt occidere; sed potius eum timete, qui potest et animam et corpus perdere in gehenna.
MATT|10|29|Nonne duo passeres asse veneunt? Et unus ex illis non cadet super terram sine Patre vestro.
MATT|10|30|Vestri autem et capilli capitis omnes numerati sunt.
MATT|10|31|Nolite ergo timere; multis passeribus meliores estis vos.
MATT|10|32|Omnis ergo qui confitebitur me coram hominibus, confitebor et ego eum coram Patre meo, qui est in caelis;
MATT|10|33|qui autem negaverit me coram hominibus, negabo et ego eum coram Patre meo, qui est in caelis.
MATT|10|34|Nolite arbitrari quia venerim mittere pacem in terram; non veni pacem mittere sed gladium.
MATT|10|35|Veni enim separarehominem adversus patrem suumet filiam adversus matrem suamet nurum adversus socrum suam:
MATT|10|36|et inimici hominis domestici eius.
MATT|10|37|Qui amat patrem aut matrem plus quam me, non est me dignus; et, qui amat filium aut filiam super me, non est me dignus;
MATT|10|38|et, qui non accipit crucem suam et sequitur me, non est me dignus.
MATT|10|39|Qui invenerit animam suam, perdet illam; et, qui perdiderit animam suam propter me, inveniet eam.
MATT|10|40|Qui recipit vos, me recipit; et, qui me recipit, recipit eum, qui me misit.
MATT|10|41|Qui recipit prophetam in nomine prophetae, mercedem prophetae accipiet; et, qui recipit iustum in nomine iusti, mercedem iusti accipiet.
MATT|10|42|Et, quicumque potum dederit uni ex minimis istis calicem aquae frigidae tantum in nomine discipuli, amen dico vobis: Non perdet mercedem suam ".
MATT|11|1|Et factum est, cum consum masset Iesus praecipiens Duodecim discipulis suis, transiit inde, ut doceret et praedicaret in civitatibus eorum.
MATT|11|2|Ioannes autem, cum audisset in vinculis opera Christi, mittens per discipulos suos
MATT|11|3|ait illi: " Tu es qui venturus es, an alium exspectamus? ".
MATT|11|4|Et respondens Iesus ait illis: " Euntes renuntiate Ioanni, quae auditis et videtis:
MATT|11|5|caeci vident et claudi ambulant, leprosi mundantur et surdi audiunt et mortui resurgunt et pauperes evangelizantur;
MATT|11|6|et beatus est, qui non fuerit scandalizatus in me ".
MATT|11|7|Illis autem abeuntibus, coepit Iesus dicere ad turbas de Ioanne: " Quid existis in desertum videre? Arundinem vento agitatam?
MATT|11|8|Sed quid existis videre? Hominem mollibus vestitum? Ecce, qui mollibus vestiuntur, in domibus regum sunt.
MATT|11|9|Sed quid existis videre? Prophetam? Etiam, dico vobis, et plus quam prophetam.
MATT|11|10|Hic est, de quo scriptum est:Ecce ego mitto angelum meum ante faciem tuam,qui praeparabit viam tuam ante te".
MATT|11|11|Amen dico vobis: Non surrexit inter natos mulierum maior Ioanne Baptista; qui autem minor est in regno caelorum, maior est illo.
MATT|11|12|A diebus autem Ioannis Baptistae usque nunc regnum caelorum vim patitur, et violenti rapiunt illud.
MATT|11|13|Omnes enim Prophetae et Lex usque ad Ioannem prophetaverunt;
MATT|11|14|et si vultis recipere, ipse est Elias, qui venturus est.
MATT|11|15|Qui habet aures, audiat.
MATT|11|16|Cui autem similem aestimabo generationem istam? Similis est pueris sedentibus in foro, qui clamantes coaequalibus
MATT|11|17|dicunt:Cecinimus vobis, et non saltastis;lamentavimus, et non planxistis".
MATT|11|18|Venit enim Ioannes neque manducans neque bibens, et dicunt: "Daemonium habet!";
MATT|11|19|venit Filius hominis manducans et bibens, et dicunt: "Ecce homo vorax et potator vini, publicanorum amicus et peccatorum!". Et iustificata est sapientia ab operibus suis ".
MATT|11|20|Tunc coepit exprobrare civitatibus, in quibus factae sunt plurimae virtutes eius, quia non egissent paenitentiam:
MATT|11|21|" Vae tibi, Chorazin! Vae tibi, Bethsaida! Quia si in Tyro et Sidone factae essent virtutes, quae factae sunt in vobis, olim in cilicio et cinere paenitentiam egissent.
MATT|11|22|Verumtamen dico vobis: Tyro et Sidoni remissius erit in die iudicii quam vobis.
MATT|11|23|Et tu, Capharnaum, numquid usque in caelum exaltaberis? Usque in infernum descendes! Quia si in Sodomis factae fuissent virtutes, quae factae sunt in te, mansissent usque in hunc diem.
MATT|11|24|Verumtamen dico vobis: Terrae Sodomorum remissius erit in die iudicii quam tibi ".
MATT|11|25|In illo tempore respondens Iesus dixit: " Confiteor tibi, Pater, Domine caeli et terrae, quia abscondisti haec a sapientibus et prudentibus et revelasti ea parvulis.
MATT|11|26|Ita, Pater, quoniam sic fuit placitum ante te.
MATT|11|27|Omnia mihi tradita sunt a Patre meo; et nemo novit Filium nisi Pater, neque Patrem quis novit nisi Filius et cui voluerit Filius revelare.
MATT|11|28|Venite ad me, omnes, qui laboratis et onerati estis, et ego reficiam vos.
MATT|11|29|Tollite iugum meum super vos et discite a me, quia mitis sum et humilis corde, et invenietis requiem animabus vestris.
MATT|11|30|Iugum enim meum suave, et onus meum leve est ".
MATT|12|1|In illo tempore abiit Iesus sabbatis per sata; discipuli autem eius esurierunt et coeperunt vellere spicas et manducare.
MATT|12|2|Pharisaei autem videntes dixerunt ei: " Ecce discipuli tui faciunt, quod non licet facere sabbato ".
MATT|12|3|At ille dixit eis: " Non legistis quid fecerit David, quando esuriit, et qui cum eo erant?
MATT|12|4|Quomodo intravit in domum Dei et panes propositionis comedit, quod non licebat ei edere neque his, qui cum eo erant, nisi solis sacerdotibus?
MATT|12|5|Aut non legistis in Lege quia sabbatis sacerdotes in templo sabbatum violant et sine crimine sunt?
MATT|12|6|Dico autem vobis quia templo maior est hic.
MATT|12|7|Si autem sciretis quid est: "Misericordiam volo et non sacrificium", numquam condemnassetis innocentes.
MATT|12|8|Dominus est enim Filius hominis sabbati ".
MATT|12|9|Et cum inde transisset, venit in synagogam eorum;
MATT|12|10|et ecce homo manum habens aridam. Et interrogabant eum dicentes: " Licet sabbatis curare? ", ut accusarent eum.
MATT|12|11|Ipse autem dixit illis: " Quis erit ex vobis homo, qui habeat ovem unam et, si ceciderit haec sabbatis in foveam, nonne tenebit et levabit eam?
MATT|12|12|Quanto igitur melior est homo ove! Itaque licet sabbatis bene facere ".
MATT|12|13|Tunc ait homini: " Extende manum tuam ". Et extendit, et restituta est sana sicut altera.
MATT|12|14|Exeuntes autem pharisaei consilium faciebant adversus eum, quomodo eum perderent.
MATT|12|15|Iesus autem sciens secessit inde. Et secuti sunt eum multi, et curavit eos omnes
MATT|12|16|et comminatus est eis, ne manifestum eum facerent,
MATT|12|17|ut adimpleretur, quod dictum est per Isaiam prophetam dicentem:
MATT|12|18|" Ecce puer meus, quem elegi,dilectus meus, in quo bene placuit animae meae;ponam Spiritum meum super eum,et iudicium gentibus nuntiabit.
MATT|12|19|Non contendet neque clamabit,neque audiet aliquis in plateis vocem eius.
MATT|12|20|Arundinem quassatam non confringetet linum fumigans non exstinguet,donec eiciat ad victoriam iudicium;
MATT|12|21|et in nomine eius gentes sperabunt ".
MATT|12|22|Tunc oblatus est ei daemonium habens, caecus et mutus, et curavit eum, ita ut mutus loqueretur et videret.
MATT|12|23|Et stupebant omnes turbae et dicebant: " Numquid hic est filius David?.
MATT|12|24|Pharisaei autem audientes dixerunt: " Hic non eicit daemones nisi in Beelzebul, principe daemonum ".
MATT|12|25|Sciens autem cogitationes eorum dixit eis: " Omne regnum divisum contra se desolatur, et omnis civitas vel domus divisa contra se non stabit.
MATT|12|26|Et si Satanas Satanam eicit, adversus se divisus est; quomodo ergo stabit regnum eius?
MATT|12|27|Et si ego in Beelzebul eicio daemones, filii vestri in quo eiciunt? Ideo ipsi iudices erunt vestri.
MATT|12|28|Si autem in Spiritu Dei ego eicio daemones, igitur pervenit in vos regnum Dei.
MATT|12|29|Aut quomodo potest quisquam intrare in domum fortis et vasa eius diripere, nisi prius alligaverit fortem? Et tunc domum illius diripiet.
MATT|12|30|Qui non est mecum, contra me est; et, qui non congregat mecum, spargit.
MATT|12|31|Ideo dico vobis: Omne peccatum et blasphemia remittetur hominibus, Spiritus autem blasphemia non remittetur.
MATT|12|32|Et quicumque dixerit verbum contra Filium hominis, remittetur ei; qui autem dixerit contra Spiritum Sanctum, non remittetur ei neque in hoc saeculo neque in futuro.
MATT|12|33|Aut facite arborem bonam et fructum eius bonum, aut facite arborem malam et fructum eius malum: si quidem ex fructu arbor agnoscitur.
MATT|12|34|Progenies viperarum, quomodo potestis bona loqui, cum sitis mali? Ex abundantia enim cordis os loquitur.
MATT|12|35|Bonus homo de bono thesauro profert bona, et malus homo de malo thesauro profert mala.
MATT|12|36|Dico autem vobis: Omne verbum otiosum, quod locuti fuerint homines, reddent rationem de eo in die iudicii:
MATT|12|37|ex verbis enim tuis iustificaberis, et ex verbis tuis condemnaberis ".
MATT|12|38|Tunc responderunt ei quidam de scribis et pharisaeis dicentes: " Magister, volumus a te signum videre ".
MATT|12|39|Qui respondens ait illis: " Generatio mala et adultera signum requirit; et signum non dabitur ei, nisi signum Ionae prophetae.
MATT|12|40|Sicut enim fuit Ionas in ventre ceti tribus diebus et tribus noctibus, sic erit Filius hominis in corde terrae tribus diebus et tribus noctibus.
MATT|12|41|Viri Ninevitae surgent in iudicio cum generatione ista et condemnabunt eam, quia paenitentiam egerunt in praedicatione Ionae; et ecce plus quam Iona hic!
MATT|12|42|Regina austri surget in iudicio cum generatione ista et condemnabit eam, quia venit a finibus terrae audire sapientiam Salomonis; et ecce plus quam Salomon hic!
MATT|12|43|Cum autem immundus spiritus exierit ab homine, ambulat per loca arida quaerens requiem et non invenit.
MATT|12|44|Tunc dicit: "Revertar in domum meam unde exivi"; et veniens invenit vacantem, scopis mundatam et ornatam.
MATT|12|45|Tunc vadit et assumit secum septem alios spiritus nequiores se, et intrantes habitant ibi; et fiunt novissima hominis illius peiora prioribus. Sic erit et generationi huic pessimae ".
MATT|12|46|Adhuc eo loquente ad turbas, ecce mater et fratres eius stabant foris quaerentes loqui ei.
MATT|12|47|Dixit autem ei quidam: " Ecce mater tua et fratres tui foris stant quaerentes loqui tecum ".
MATT|12|48|At ille respondens dicenti sibi ait: " Quae est mater mea, et qui sunt fratres mei? ".
MATT|12|49|Et extendens manum suam in discipulos suos dixit: " Ecce mater mea et fratres mei.
MATT|12|50|Quicumque enim fecerit voluntatem Patris mei, qui in caelis est, ipse meus frater et soror et mater est ".
MATT|13|1|In illo die exiens Iesus de domo sedebat secus mare;
MATT|13|2|et congregatae sunt ad eum turbae multae, ita ut in naviculam ascendens sederet, et omnis turba stabat in litore.
MATT|13|3|Et locutus est eis multa in parabolis dicens: " Ecce exiit, qui seminat, seminare.
MATT|13|4|Et dum seminat, quaedam ceciderunt secus viam, et venerunt volucres et comederunt ea.
MATT|13|5|Alia autem ceciderunt in petrosa, ubi non habebant terram multam, et continuo exorta sunt, quia non habebant altitudinem terrae;
MATT|13|6|sole autem orto, aestuaverunt et, quia non habebant radicem, aruerunt.
MATT|13|7|Alia autem ceciderunt in spinas, et creverunt spinae et suffocaverunt ea.
MATT|13|8|Alia vero ceciderunt in terram bonam et dabant fructum: aliud centesimum, aliud sexagesimum, aliud tricesimum.
MATT|13|9|Qui habet aures, audiat ".
MATT|13|10|Et accedentes discipuli dixerunt ei: " Quare in parabolis loqueris eis?.
MATT|13|11|Qui respondens ait illis: " Quia vobis datum est nosse mysteria regni caelorum, illis autem non est datum.
MATT|13|12|Qui enim habet, dabitur ei, et abundabit; qui autem non habet, et quod habet, auferetur ab eo.
MATT|13|13|Ideo in parabolis loquor eis, quia videntes non vident et audientes non audiunt neque intellegunt;
MATT|13|14|et adimpletur eis prophetia Isaiae dicens:Auditu audietis et non intellegetiset videntes videbitis et non videbitis.
MATT|13|15|Incrassatum est enim cor populi huius,et auribus graviter audieruntet oculos suos clauserunt,ne quando oculis videantet auribus audiantet corde intellegant et convertantur,et sanem eos".
MATT|13|16|Vestri autem beati oculi, quia vident, et aures vestrae, quia audiunt.
MATT|13|17|Amen quippe dico vobis: Multi prophetae et iusti cupierunt videre, quae videtis, et non viderunt, et audire, quae auditis, et non audierunt!
MATT|13|18|Vos ergo audite parabolam seminantis.
MATT|13|19|Omnis, qui audit verbum regni et non intellegit, venit Malus et rapit, quod seminatum est in corde eius; hic est, qui secus viam seminatus est.
MATT|13|20|Qui autem supra petrosa seminatus est, hic est, qui verbum audit et continuo cum gaudio accipit illud,
MATT|13|21|non habet autem in se radicem, sed est temporalis; facta autem tribulatione vel persecutione propter verbum, continuo scandalizatur.
MATT|13|22|Qui autem est seminatus in spinis, hic est, qui verbum audit, et sollicitudo saeculi et fallacia divitiarum suffocat verbum, et sine fructu efficitur.
MATT|13|23|Qui vero in terra bona seminatus est, hic est, qui audit verbum et intellegit et fructum affert et facit aliud quidem centum, aliud autem sexaginta, porro aliud triginta ".
MATT|13|24|Aliam parabolam proposuit illis dicens: " Simile factum est regnum caelorum homini, qui seminavit bonum semen in agro suo.
MATT|13|25|Cum autem dormirent homines, venit inimicus eius et superseminavit zizania in medio tritici et abiit.
MATT|13|26|Cum autem crevisset herba et fructum fecisset, tunc apparuerunt et zizania.
MATT|13|27|Accedentes autem servi patris familias dixerunt ei: "Domine, nonne bonum semen seminasti in agro tuo? Unde ergo habet zizania?".
MATT|13|28|Et ait illis: "Inimicus homo hoc fecit". Servi autem dicunt ei: "Vis, imus et colligimus ea?".
MATT|13|29|Et ait: "Non; ne forte colligentes zizania eradicetis simul cum eis triticum,
MATT|13|30|sinite utraque crescere usque ad messem. Et in tempore messis dicam messoribus: Colligite primum zizania et alligate ea in fasciculos ad comburendum ea, triticum autem congregate in horreum meum" ".
MATT|13|31|Aliam parabolam proposuit eis dicens: " Simile est regnum caelorum grano sinapis, quod accipiens homo seminavit in agro suo.
MATT|13|32|Quod minimum quidem est omnibus seminibus; cum autem creverit, maius est holeribus et fit arbor, ita ut volucres caeli veniant et habitent in ramis eius ".
MATT|13|33|Aliam parabolam locutus est eis: " Simile est regnum caelorum fermento, quod acceptum mulier abscondit in farinae satis tribus, donec fermentatum est totum ".
MATT|13|34|Haec omnia locutus est Iesus in parabolis ad turbas; et sine parabola nihil loquebatur eis,
MATT|13|35|ut adimpleretur, quod dictum erat per prophetam dicentem: Aperiam in parabolis os meum,eructabo abscondita a constitutione mundi ".
MATT|13|36|Tunc, dimissis turbis, venit in domum, et accesserunt ad eum discipuli eius dicentes: " Dissere nobis parabolam zizaniorum agri ".
MATT|13|37|Qui respondens ait: " Qui seminat bonum semen, est Filius hominis;
MATT|13|38|ager autem est mundus; bonum vero semen, hi sunt filii regni; zizania autem filii sunt Mali;
MATT|13|39|inimicus autem, qui seminavit ea, est Diabolus; messis vero consummatio saeculi est; messores autem angeli sunt.
MATT|13|40|Sicut ergo colliguntur zizania et igni comburuntur, sic erit in consummatione saeculi:
MATT|13|41|mittet Filius hominis angelos suos, et colligent de regno eius omnia scandala et eos, qui faciunt iniquitatem,
MATT|13|42|et mittent eos in caminum ignis; ibi erit fletus et stridor dentium.
MATT|13|43|Tunc iusti fulgebunt sicut sol in regno Pa tris eorum. Qui habet aures, audiat.
MATT|13|44|Simile est regnum caelorum thesauro abscondito in agro; quem qui invenit homo abscondit et prae gaudio illius vadit et vendit universa, quae habet, et emit agrum illum.
MATT|13|45|Iterum simile est regnum caelorum homini negotiatori quaerenti bonas margaritas.
MATT|13|46|Inventa autem una pretiosa margarita, abiit et vendidit omnia, quae habuit, et emit eam.
MATT|13|47|Iterum simile est regnum caelorum sagenae missae in mare et ex omni genere congreganti;
MATT|13|48|quam, cum impleta esset, educentes secus litus et sedentes collegerunt bonos in vasa, malos autem foras miserunt.
MATT|13|49|Sic erit in consummatione saeculi: exibunt angeli et separabunt malos de medio iustorum
MATT|13|50|et mittent eos in caminum ignis; ibi erit fletus et stridor dentium.
MATT|13|51|Intellexistis haec omnia? ". Dicunt ei: " Etiam ".
MATT|13|52|Ait autem illis: " Ideo omnis scriba doctus in regno caelorum similis est homini patri familias, qui profert de thesauro suo nova et vetera ".
MATT|13|53|Et factum est, cum consummasset Iesus parabolas istas, transiit inde.
MATT|13|54|Et veniens in patriam suam, docebat eos in synagoga eorum, ita ut mirarentur et dicerent: " Unde huic sapientia haec et virtutes?
MATT|13|55|Nonne hic est fabri filius? Nonne mater eius dicitur Maria, et fratres eius Iacobus et Ioseph et Simon et Iudas?
MATT|13|56|Et sorores eius nonne omnes apud nos sunt? Unde ergo huic omnia ista?.
MATT|13|57|Et scandalizabantur in eo. Iesus autem dixit eis: " Non est propheta sine honore nisi in patria et in domo sua ".
MATT|13|58|Et non fecit ibi virtutes multas propter incredulitatem illorum.
MATT|14|1|In illo tempore audivit He rodes tetrarcha famam Iesu
MATT|14|2|et ait pueris suis: " Hic est Ioannes Baptista; ipse surrexit a mortuis, et ideo virtutes operantur in eo ".
MATT|14|3|Herodes enim tenuit Ioannem et alligavit eum et posuit in carcere propter Herodiadem uxorem Philippi fratris sui.
MATT|14|4|Dicebat enim illi Ioannes: " Non licet tibi habere eam ".
MATT|14|5|Et volens illum occidere, timuit populum, quia sicut prophetam eum habebant.
MATT|14|6|Die autem natalis Herodis saltavit filia Herodiadis in medio et placuit Herodi,
MATT|14|7|unde cum iuramento pollicitus est ei dare, quodcumque postulasset.
MATT|14|8|At illa, praemonita a matre sua: " Da mihi, inquit, hic in disco caput Ioannis Baptistae ".
MATT|14|9|Et contristatus rex propter iuramentum et eos, qui pariter recumbebant, iussit dari
MATT|14|10|misitque et decollavit Ioannem in carcere;
MATT|14|11|et allatum est caput eius in disco et datum est puellae, et tulit matri suae.
MATT|14|12|Et accedentes discipuli eius tulerunt corpus et sepelierunt illud et venientes nuntiaverunt Iesu.
MATT|14|13|Quod cum audisset Iesus, secessit inde in navicula in locum desertum seorsum; et cum audissent, turbae secutae sunt eum pedestres de civitatibus.
MATT|14|14|Et exiens vidit turbam multam et misertus est eorum et curavit languidos eorum.
MATT|14|15|Vespere autem facto, accesserunt ad eum discipuli dicentes: " Desertus est locus, et hora iam praeteriit; dimitte turbas, ut euntes in castella emant sibi escas ".
MATT|14|16|Iesus autem dixit eis: " Non habent necesse ire; date illis vos manducare ".
MATT|14|17|Illi autem dicunt ei: " Non habemus hic nisi quinque panes et duos pisces ".
MATT|14|18|Qui ait: " Afferte illos mihi huc ".
MATT|14|19|Et cum iussisset turbas discumbere supra fenum, acceptis quinque panibus et duobus piscibus, aspiciens in caelum benedixit et fregit et dedit discipulis panes, discipuli autem turbis.
MATT|14|20|Et manducaverunt omnes et saturati sunt; et tulerunt reliquias fragmentorum duodecim cophinos plenos.
MATT|14|21|Manducantium autem fuit numerus fere quinque milia virorum, exceptis mulieribus et parvulis.
MATT|14|22|Et statim iussit discipulos ascendere in naviculam et praecedere eum trans fretum, donec dimitteret turbas.
MATT|14|23|Et dimissis turbis, ascendit in montem solus orare. Vespere autem facto, solus erat ibi.
MATT|14|24|Navicula autem iam multis stadiis a terra distabat, fluctibus iactata; erat enim contrarius ventus.
MATT|14|25|Quarta autem vigilia noctis venit ad eos ambulans supra mare.
MATT|14|26|Discipuli autem, videntes eum supra mare ambulantem, turbati sunt dicentes: " Phantasma est ", et prae timore clamaverunt.
MATT|14|27|Statimque Iesus locutus est eis dicens: " Habete fiduciam, ego sum; nolite timere! ".
MATT|14|28|Respondens autem ei Petrus dixit: " Domine, si tu es, iube me venire ad te super aquas ".
MATT|14|29|At ipse ait: " Veni! ". Et descendens Petrus de navicula ambulavit super aquas et venit ad Iesum.
MATT|14|30|Videns vero ventum validum timuit et, cum coepisset mergi, clamavit dicens: " Domine, salvum me fac! ".
MATT|14|31|Continuo autem Iesus extendens manum apprehendit eum et ait illi: " Modicae fidei, quare dubitasti? ".
MATT|14|32|Et cum ascendissent in naviculam, cessavit ventus.
MATT|14|33|Qui autem in navicula erant, adoraverunt eum dicentes: " Vere Filius Dei es! ".
MATT|14|34|Et cum transfretassent, venerunt in terram Gennesaret.
MATT|14|35|Et cum cognovissent eum viri loci illius, miserunt in universam regionem illam et obtulerunt ei omnes male habentes,
MATT|14|36|et rogabant eum, ut vel fimbriam vestimenti eius tangerent; et, quicumque tetigerunt, salvi facti sunt.
MATT|15|1|Tunc accedunt ad Iesum ab Hierosolymis pharisaei et scribae dicentes:
MATT|15|2|" Quare discipuli tui transgrediuntur traditionem seniorum? Non enim lavant manus suas, cum panem manducant ".
MATT|15|3|Ipse autem respondens ait illis: " Quare et vos transgredimini mandatum Dei propter traditionem vestram?
MATT|15|4|Nam Deus dixit: "Honora patrem tuum et matrem" et: "Qui maledixerit patri vel matri, morte moriatur".
MATT|15|5|Vos autem dicitis: "Quicumque dixerit patri vel matri: Munus est, quodcumque ex me profuerit,
MATT|15|6|non honorificabit patrem suum"; et irritum fecistis verbum Dei propter traditionem vestram.
MATT|15|7|Hypocritae! Bene prophetavit de vobis Isaias dicens:
MATT|15|8|"Populus hic labiis me honorat,cor autem eorum longe est a me;
MATT|15|9|sine causa autem colunt medocentes doctrinas mandata homi num" ".
MATT|15|10|Et convocata ad se turba, dixit eis: " Audite et intellegite:
MATT|15|11|Non quod intrat in os, coinquinat hominem; sed quod procedit ex ore, hoc coinquinat hominem! ".
MATT|15|12|Tunc accedentes discipuli dicunt ei: " Scis quia pharisaei, audito verbo, scandalizati sunt? ".
MATT|15|13|At ille respondens ait: " Omnis plantatio, quam non plantavit Pater meus caelestis, eradicabitur.
MATT|15|14|Sinite illos: caeci sunt, duces caecorum. Caecus autem si caeco ducatum praestet, ambo in foveam cadent ".
MATT|15|15|Respondens autem Petrus dixit ei: " Edissere nobis parabolam istam ".
MATT|15|16|At ille dixit: " Adhuc et vos sine intellectu estis?
MATT|15|17|Non intellegitis quia omne quod in os intrat, in ventrem vadit et in secessum emittitur?
MATT|15|18|Quae autem procedunt de ore, de corde exeunt, et ea coinquinant hominem.
MATT|15|19|De corde enim exeunt cogitationes malae, homicidia, adulteria, fornicationes, furta, falsa testimonia, blasphemiae.
MATT|15|20|Haec sunt, quae coinquinant hominem; non lotis autem manibus manducare non coinquinat hominem ".
MATT|15|21|Et egressus inde Iesus, secessit in partes Tyri et Sidonis.
MATT|15|22|Et ecce mulier Chananaea a finibus illis egressa clamavit dicens: " Miserere mei, Domine, fili David! Filia mea male a daemonio vexatur ".
MATT|15|23|Qui non respondit ei verbum.Et accedentes discipuli eius rogabant eum dicentes: " Dimitte eam, quia clamat post nos ".
MATT|15|24|Ipse autem respondens ait: " Non sum missus nisi ad oves, quae perierunt domus Israel ".
MATT|15|25|At illa venit et adoravit eum dicens: " Domine, adiuva me! ".
MATT|15|26|Qui respondens ait: " Non est bonum sumere panem filiorum et mittere catellis ".
MATT|15|27|At illa dixit: " Etiam, Domine, nam et catelli edunt de micis, quae cadunt de mensa dominorum suorum ".
MATT|15|28|Tunc respondens Iesus ait illi: " O mulier, magna est fides tua! Fiat tibi, sicut vis ". Et sanata est filia illius ex illa hora.
MATT|15|29|Et cum transisset inde, Iesus venit secus mare Galilaeae et ascendens in montem sedebat ibi.
MATT|15|30|Et accesserunt ad eum turbae multae habentes secum claudos, caecos, debiles, mutos et alios multos et proiecerunt eos ad pedes eius, et curavit eos,
MATT|15|31|ita ut turba miraretur videntes mutos loquentes, debiles sanos et claudos ambulantes et caecos videntes. Et magnificabant Deum Israel.
MATT|15|32|Iesus autem convocatis discipulis suis dixit: " Misereor turbae, quia triduo iam perseverant mecum et non habent, quod manducent; et dimittere eos ieiunos nolo, ne forte deficiant in via ".
MATT|15|33|Et dicunt ei discipuli: " Unde nobis in deserto panes tantos, ut saturemus turbam tantam? ".
MATT|15|34|Et ait illis Iesus: " Quot panes habetis? ". At illi dixerunt: " Septem et paucos pisciculos ".
MATT|15|35|Et praecepit turbae, ut discumberet super terram;
MATT|15|36|et accipiens septem panes et pisces et gratias agens fregit et dedit discipulis, discipuli autem turbis.
MATT|15|37|Et comederunt omnes et saturati sunt; et, quod superfuit de fragmentis, tulerunt septem sportas plenas.
MATT|15|38|Erant autem, qui manducaverant, quattuor milia hominum extra mulieres et parvulos.
MATT|15|39|Et dimissis turbis, ascendit in naviculam et venit in fines Magadan.
MATT|16|1|Et accesserunt ad eum pharisaei et sadducaei tentantes et rogaverunt eum, ut signum de caelo ostenderet eis.
MATT|16|2|At ille respondens ait eis: " Facto vespere dicitis: "Serenum erit, rubicundum est enim caelum";
MATT|16|3|et mane: "Hodie tempestas, rutilat enim triste caelum". Faciem quidem caeli diiudicare nostis, signa autem temporum non potestis.
MATT|16|4|Generatio mala et adultera signum quaerit, et signum non dabitur ei, nisi signum Ionae ". Et, relictis illis, abiit.
MATT|16|5|Et cum venissent discipuli trans fretum, obliti sunt panes accipere.
MATT|16|6|Iesus autem dixit illis: " Intuemini et cavete a fermento pharisaeorum et sadducaeorum ".
MATT|16|7|At illi cogitabant inter se dicentes: " Panes non accepimus!".
MATT|16|8|Sciens autem Iesus dixit: " Quid cogitatis inter vos, modicae fidei, quia panes non habetis?
MATT|16|9|Nondum intellegitis neque recordamini quinque panum quinque milium hominum, et quot cophinos sumpsistis?
MATT|16|10|Neque septem panum quattuor milium hominum, et quot sportas sumpsistis?
MATT|16|11|Quomodo non intellegitis quia non de panibus dixi vobis? Sed cavete a fermento pharisaeorum et sadducaeorum ".
MATT|16|12|Tunc intellexerunt quia non dixerit cavendum a fermento panum sed a doctrina pharisaeorum et sadducaeorum.
MATT|16|13|Venit autem Iesus in partes Caesareae Philippi et interrogabat discipulos suos dicens: " Quem dicunt homines esse Filium hominis?".
MATT|16|14|At illi dixerunt: " Alii Ioannem Baptistam, alii autem Eliam, alii vero Ieremiam, aut unum ex prophetis ".
MATT|16|15|Dicit illis: " Vos autem quem me esse dicitis? ".
MATT|16|16|Respondens Simon Petrus dixit: " Tu es Christus, Filius Dei vivi ".
MATT|16|17|Respondens autem Iesus dixit ei: " Beatus es, Simon Bariona, quia caro et sanguis non revelavit tibi sed Pater meus, qui in caelis est.
MATT|16|18|Et ego dico tibi: Tu es Petrus, et super hanc petram aedificabo Ecclesiam meam; et portae inferi non praevalebunt adversum eam.
MATT|16|19|Tibi dabo claves regni caelorum; et quodcumque ligaveris super terram, erit ligatum in caelis, et quodcumque solveris super terram, erit solutum in caelis ".
MATT|16|20|Tunc praecepit discipulis, ut nemini dicerent quia ipse esset Christus.
MATT|16|21|Exinde coepit Iesus ostendere discipulis suis quia oporteret eum ire Hierosolymam et multa pati a senioribus et principibus sacerdotum et scribis et occidi et tertia die resurgere.
MATT|16|22|Et assumens eum Petrus coepit increpare illum dicens: " Absit a te, Domine; non erit tibi hoc ".
MATT|16|23|Qui conversus dixit Petro: " Vade post me, Satana! Scandalum es mihi, quia non sapis ea, quae Dei sunt, sed ea, quae hominum! ".
MATT|16|24|Tunc Iesus dixit discipulis suis: " Si quis vult post me venire, abneget semetipsum et tollat crucem suam et sequatur me.
MATT|16|25|Qui enim voluerit animam suam salvam facere, perdet eam; qui autem perdiderit animam suam propter me, inveniet eam.
MATT|16|26|Quid enim prodest homini, si mundum universum lucretur, animae vero suae detrimentum patiatur? Aut quam dabit homo commutationem pro anima sua?
MATT|16|27|Filius enim hominis venturus est in gloria Patris sui cum angelis suis, et tunc reddet unicuique secundum opus eius.
MATT|16|28|Amen dico vobis: Sunt quidam de hic stantibus, qui non gustabunt mortem, donec videant Filium hominis venientem in regno suo ".
MATT|17|1|Et post dies sex assumit Iesus Petrum et Iacobum et Ioan nem fratrem eius et ducit illos in montem excelsum seorsum.
MATT|17|2|Et transfiguratus est ante eos; et resplenduit facies eius sicut sol, vestimenta autem eius facta sunt alba sicut lux.
MATT|17|3|Et ecce apparuit illis Moyses et Elias cum eo loquentes.
MATT|17|4|Respondens autem Petrus dixit ad Iesum: " Domine, bonum est nos hic esse. Si vis, faciam hic tria tabernacula: tibi unum et Moysi unum et Eliae unum ".
MATT|17|5|Adhuc eo loquente, ecce nubes lucida obumbravit eos; et ecce vox de nube dicens: " Hic est Filius meus dilectus, in quo mihi bene complacui; ipsum audite ".
MATT|17|6|Et audientes discipuli ceciderunt in faciem suam et timuerunt valde.
MATT|17|7|Et accessit Iesus et tetigit eos dixitque eis: " Surgite et nolite timere ".
MATT|17|8|Levantes autem oculos suos, neminem viderunt nisi solum Iesum.
MATT|17|9|Et descendentibus illis de monte, praecepit eis Iesus dicens: " Nemini dixeritis visionem, donec Filius hominis a mortuis resurgat ".
MATT|17|10|Et interrogaverunt eum discipuli dicentes: " Quid ergo scribae dicunt quod Eliam oporteat primum venire? ".
MATT|17|11|At ille respondens ait: " Elias quidem venturus est et restituet omnia.
MATT|17|12|Dico autem vobis quia Elias iam venit, et non cognoverunt eum, sed fecerunt in eo, quaecumque voluerunt; sic et Filius hominis passurus est ab eis ".
MATT|17|13|Tunc intellexerunt discipuli quia de Ioanne Baptista dixisset eis.
MATT|17|14|Et cum venissent ad turbam, accessit ad eum homo genibus provolutus ante eum
MATT|17|15|et dicens: " Domine, miserere filii mei, quia lunaticus est et male patitur; nam saepe cadit in ignem et crebro in aquam.
MATT|17|16|Et obtuli eum discipulis tuis, et non potuerunt curare eum ".
MATT|17|17|Respondens autem Iesus ait: " O generatio incredula et perversa, quousque ero vobiscum? Usquequo patiar vos? Afferte huc illum ad me ".
MATT|17|18|Et increpavit eum Iesus, et exiit ab eo daemonium, et curatus est puer ex illa hora.
MATT|17|19|Tunc accesserunt discipuli ad Iesum secreto et dixerunt: " Quare nos non potuimus eicere illum? ".
MATT|17|20|Ille autem dicit illis: " Propter modicam fidem vestram. Amen quippe dico vobis: Si habueritis fidem sicutgranum sinapis, dicetis monti huic: "Transi hinc illuc!", et transibit, et nihil impossibile erit vobis ".
MATT|17|21|()
MATT|17|22|Conversantibus autem eis in Galilaea, dixit illis Iesus: " Filius hominis tradendus est in manus hominum,
MATT|17|23|et occident eum, et tertio die resurget ". Et contristati sunt vehementer.
MATT|17|24|Et cum venissent Capharnaum, accesserunt, qui didrachma accipiebant, ad Petrum et dixerunt: " Magister vester non solvit didrachma? ".
MATT|17|25|Ait: " Etiam". Et cum intrasset domum, praevenit eum Iesus dicens: " Quid tibi videtur, Simon? Reges terrae a quibus accipiunt tributum vel censum? A filiis suis an ab alienis? ".
MATT|17|26|Cum autem ille dixisset: " Ab alienis ", dixit illi Iesus: " Ergo liberi sunt filii.
MATT|17|27|Ut autem non scandalizemus eos, vade ad mare et mitte hamum; et eum piscem, qui primus ascenderit, tolle; et, aperto ore, eius invenies staterem. Illum sumens, da eis pro me et te ".
MATT|18|1|In illa hora accesserunt di scipuli ad Iesum dicentes: " Quis putas maior est in regno caelorum? ".
MATT|18|2|Et advocans parvulum, statuit eum in medio eorum
MATT|18|3|et dixit: " Amen dico vobis: Nisi conversi fueritis et efiiciamini sicut parvuli, non intrabitis in regnum caelorum.
MATT|18|4|Quicumque ergo humiliaverit se sicut parvulus iste, hic est maior in regno caelorum.
MATT|18|5|Et, qui susceperit unum parvulum talem in nomine meo, me suscipit.
MATT|18|6|Qui autem scandalizaverit unum de pusillis istis, qui in me credunt, expedit ei, ut suspendatur mola asinaria in collo eius et demergatur in profundum maris.
MATT|18|7|Vae mundo ab scandalis! Necesse est enim ut veniant scandala; verumtamen vae homini, per quem scandalum venit!
MATT|18|8|Si autem manus tua vel pes tuus scandalizat te, abscide eum et proice abs te: bonum tibi est ad vitam ingredi debilem vel claudum, quam duas manus vel duos pedes habentem mitti in ignem aeternum.
MATT|18|9|Et si oculus tuus scandalizat te, erue eum et proice abs te: bonum tibi est unoculum in vitam intrare, quam duos oculos habentem mitti in gehennam ignis.
MATT|18|10|Videte, ne contemnatis unum ex his pusillis; dico enim vobis quia angeli eorum in caelis sempervident faciem Patris mei, qui in caelis est.
MATT|18|11|()
MATT|18|12|Quid vobis videtur? Si fuerint alicui centum oves, et erraverit una ex eis, nonne relinquet nonaginta novem in montibus et vadit quaerere eam, quae erravit?
MATT|18|13|Et si contigerit ut inveniat eam, amen dico vobis quia gaudebit super eam magis quam super nonaginta novem, quae non erraverunt.
MATT|18|14|Sic non est voluntas ante Patrem vestrum, qui in caelis est, ut pereat unus de pusillis istis.
MATT|18|15|Si autem peccaverit in te frater tuus, vade, corripe eum inter te et ipsum solum. Si te audierit, lucratus es fratrem tuum;
MATT|18|16|si autem non audierit, adhibe tecum adhuc unum vel duos, ut in ore duorum testium vel trium stet omne verbum;
MATT|18|17|quod si noluerit audire eos, dic ecclesiae; si autem et ecclesiam noluerit audire, sit tibi sicut ethnicus et publicanus.
MATT|18|18|Amen dico vobis: Quaecumque alligaveritis super terram, erunt ligata in caelo; et, quaecumque solveritis super terram, erunt soluta in caelo.
MATT|18|19|Iterum dico vobis: Si duo ex vobis consenserint super terram de omni re, quamcumque petierint, fiet illis a Patre meo, qui in caelis est.
MATT|18|20|Ubi enim sunt duo vel tres congregati in nomine meo, ibi sum in medio eorum ".
MATT|18|21|Tunc accedens Petrus dixit ei: " Domine, quotiens peccabit in me frater meus, et dimittam ei? Usque septies? ".
MATT|18|22|Dicit illi Iesus: " Non dico tibi usque septies sed usque septuagies septies.
MATT|18|23|Ideo assimilatum est regnum caelorum homini regi, qui voluit rationem ponere cum servis suis.
MATT|18|24|Et cum coepisset rationem ponere, oblatus est ei unus, qui debebat decem milia talenta.
MATT|18|25|Cum autem non haberet, unde redderet, iussit eum dominus venumdari et uxorem et filios et omnia, quae habebat, et reddi.
MATT|18|26|Procidens igitur servus ille adorabat eum dicens: "Patientiam habe in me, et omnia reddam tibi".
MATT|18|27|Misertus autem dominus servi illius dimisit eum et debitum dimisit ei.
MATT|18|28|Egressus autem servus ille invenit unum de conservis suis, qui debebat ei centum denarios, et tenens suffocabat eum dicens: "Redde, quod debes!".
MATT|18|29|Procidens igitur conservus eius rogabat eum dicens: "Patientiam habe in me, et reddam tibi".
MATT|18|30|Ille autem noluit, sed abiit et misit eum in carcerem, donec redderet debitum.
MATT|18|31|Videntes autem conservi eius, quae fiebant, contristati sunt valde et venerunt et narraverunt domino suo omnia, quae facta erant.
MATT|18|32|Tunc vocavit illum dominus suus et ait illi: "Serve nequam, omne debitum illud dimisi tibi, quoniam rogasti me;
MATT|18|33|non oportuit et te misereri conservi tui, sicut et ego tui misertus sum?".
MATT|18|34|Et iratus dominus eius tradidit eum tortoribus, quoadusque redderet universum debitum.
MATT|18|35|Sic et Pater meus caelestis faciet vobis, si non remiseritis unusquisque fratri suo de cordibus vestris ".
MATT|19|1|Et factum est, cum consum masset Iesus sermones istos, migravit a Galilaea et venit in fines Iudaeae trans Iordanem.
MATT|19|2|Et secutae sunt eum turbae multae, et curavit eos ibi.
MATT|19|3|Et accesserunt ad eum pharisaei tentantes eum et dicentes: " Licet homini dimittere uxorem suam quacumque ex causa? ".
MATT|19|4|Qui respondens ait: " Non legistis quia, qui creavit ab initio, masculum et feminam fecit eos
MATT|19|5|et dixit: "Propter hoc dimittet homo patrem et matrem et adhaerebit uxori suae, et erunt duo in carne una?".
MATT|19|6|Itaque iam non sunt duo sed una caro. Quod ergo Deus coniunxit, homo non separet ".
MATT|19|7|Dicunt illi: " Quid ergo Moyses mandavit dari libellum repudii et dimittere? ".
MATT|19|8|Ait illis: " Moyses ad duritiam cordis vestri permisit vobis dimittere uxores vestras; ab initio autem non sic fuit.
MATT|19|9|Dico autem vobis quia quicumque dimiserit uxorem suam, nisi ob fornicationem, et aliam duxerit, moechatur ".
MATT|19|10|Dicunt ei discipuli eius: " Si ita est causa hominis cum uxore, non expedit nubere ".
MATT|19|11|Qui dixit eis: " Non omnes capiunt verbum istud, sed quibus datum est.
MATT|19|12|Sunt enim eunuchi, qui de matris utero sic nati sunt; et sunt eunuchi, qui facti sunt ab hominibus; et sunt eunuchi, qui seipsos castraverunt propter regnum caelorum. Qui potest capere, capiat ".
MATT|19|13|Tunc oblati sunt ei parvuli, ut manus eis imponeret et oraret; discipuli autem increpabant eis.
MATT|19|14|Iesus vero ait: " Sinite parvulos et nolite eos prohibere ad me venire; talium est enim regnum caelorum ".
MATT|19|15|Et cum imposuisset eis manus, abiit inde.
MATT|19|16|Et ecce unus accedens ait illi: " Magister, quid boni faciam, ut habeam vitam aeternam? ". Qui dixit ei:
MATT|19|17|" Quid me interrogas de bono? Unus est bonus. Si autem vis ad vitam ingredi, serva mandata ".
MATT|19|18|Dicit illi: " Quae? ". Iesus autem dixit: " Non homicidium facies, non adulterabis, non facies furtum, non falsum testimonium dices,
MATT|19|19|honora patrem et matrem et diliges proximum tuum sicut teipsum ".
MATT|19|20|Dicit illi adulescens: " Omnia haec custodivi. Quid adhuc mihi deest?.
MATT|19|21|Ait illi Iesus: " Si vis perfectus esse, vade, vende, quae habes, et da pauperibus, et habebis thesaurum in caelo; et veni, sequere me ".
MATT|19|22|Cum audisset autem adulescens verbum, abiit tristis; erat enim habens multas possessiones.
MATT|19|23|Iesus autem dixit discipulis suis: " Amen dico vobis: Dives difficile intrabit in regnum caelorum.
MATT|19|24|Et iterum dico vobis: Facilius est camelum per foramen acus transire, quam divitem intrare in regnum Dei ".
MATT|19|25|Auditis autem his, discipuli mirabantur valde dicentes: " Quis ergo poterit salvus esse? ".
MATT|19|26|Aspiciens autem Iesus dixit illis: " Apud homines hoc impossibile est, apud Deum autem omnia possibilia sunt ".
MATT|19|27|Tunc respondens Petrus dixit ei: " Ecce nos reliquimus omnia et secuti sumus te. Quid ergo erit nobis? ".
MATT|19|28|Iesus autem dixit illis: " Amen dico vobis quod vos, qui secuti estis me, in regeneratione, cum sederit Filius hominis in throno gloriae suae, sedebitis et vos super thronos duodecim, iudicantes duodecim tribus Israel.
MATT|19|29|Et omnis, qui reliquit domos vel fratres aut sorores aut patrem aut matrem aut filios aut agros propter nomen meum, centuplum accipiet et vitam aeternam possidebit.
MATT|19|30|Multi autem erunt primi novissimi, et novissimi primi.
MATT|20|1|Simile est enim regnum cae lorum homini patri familias, qui exiit primo mane conducere operarios in vineam suam;
MATT|20|2|conventione autem facta cum operariis ex denario diurno, misit eos in vineam suam.
MATT|20|3|Et egressus circa horam tertiam vidit alios stantes in foro otiosos
MATT|20|4|et illis dixit: "Ite et vos in vineam; et, quod iustum fuerit, dabo vobis".
MATT|20|5|Illi autem abierunt. Iterum autem exiit circa sextam et nonam horam et fecit similiter.
MATT|20|6|Circa undecimam vero exiit et invenit alios stantes et dicit illis: Quid hic statis tota die otiosi?".
MATT|20|7|Dicunt ei: "Quia nemo nos conduxit". Dicit illis: "Ite et vos in vineam".
MATT|20|8|Cum sero autem factum esset, dicit dominus vineae procuratori suo: " Voca operarios et redde illis mercedem incipiens a novissimis usque ad primos ".
MATT|20|9|Et cum venissent, qui circa undecimam horam venerant, acceperunt singuli denarium.
MATT|20|10|Venientes autem primi arbitrati sunt quod plus essent accepturi; acceperunt autem et ipsi singuli denarium.
MATT|20|11|Accipientes autem murmurabant adversus patrem familias
MATT|20|12|dicentes: "Hi novissimi una hora fecerunt, et pares illos nobis fecisti, qui portavimus pondus diei et aestum!".
MATT|20|13|At ille respondens uni eorum dixit: "Amice, non facio tibi iniuriam; nonne ex denario convenisti mecum?
MATT|20|14|Tolle, quod tuum est, et vade; volo autem et huic novissimo dare sicut et tibi.
MATT|20|15|Aut non licet mihi, quod volo, facere de meis? An oculus tuus nequam est, quia ego bonus sum?".
MATT|20|16|Sic erunt novissimi primi, et primi novissimi ".
MATT|20|17|Et ascendens Iesus Hierosolymam assumpsit Duodecim discipulos secreto et ait illis in via:
MATT|20|18|" Ecce ascendimus Hierosolymam, et Filius hominis tradetur principibus sacerdotum et scribis, et condemnabunt eum morte
MATT|20|19|et tradent eum gentibus ad illudendum et flagellandum et crucifigendum, et tertia die resurget ".
MATT|20|20|Tunc accessit ad eum mater filiorum Zebedaei cum filiis suis, adorans et petens aliquid ab eo.
MATT|20|21|Qui dixit ei: " Quid vis? ". Ait illi: " Dic ut sedeant hi duo filii mei unus ad dexteram tuam et unus ad sinistram in regno tuo ".
MATT|20|22|Respondens autem Iesus dixit: " Nescitis quid petatis. Potestis bibere calicem, quem ego bibiturus sum? ". Dicunt ei: " Possumus ".
MATT|20|23|Ait illis: " Calicem quidem meum bibetis, sedere autem ad dexteram meam et sinistram non est meum dare illud, sed quibus paratum est a Patre meo.
MATT|20|24|Et audientes decem indignati sunt de duobus fratribus.
MATT|20|25|Iesus autem vocavit eos ad se et ait: " Scitis quia principes gentium dominantur eorum et, qui magni sunt, potestatem exercent in eos.
MATT|20|26|Non ita erit inter vos, sed quicumque voluerit inter vos magnus fieri, erit vester minister;
MATT|20|27|et, quicumque voluerit inter vos primus esse, erit vester servus;
MATT|20|28|sicut Filius hominis non venit ministrari sed ministrare et dare animam suam redemptionem pro multis ".
MATT|20|29|Et egredientibus illis ab Iericho, secuta est eum turba multa.
MATT|20|30|Et ecce duo caeci sedentes secus viam audierunt quia Iesus transiret et clamaverunt dicentes: " Domine, miserere nostri, fili David! ".
MATT|20|31|Turba autem increpabat eos, ut tacerent; at illi magis clamabant dicentes: " Domine, miserere nostri, fili David! ".
MATT|20|32|Et stetit Iesus et vocavit eos et ait: " Quid vultis, ut faciam vobis?".
MATT|20|33|Dicunt illi: " Domine, ut aperiantur oculi nostri ".
MATT|20|34|Misertus autem Iesus, tetigit oculos eorum; et confestim viderunt et secuti sunt eum.
MATT|21|1|Et cum appropinquassent Hierosolymis et venissent Bethfage, ad montem Oliveti, tunc Iesus misit duos discipulos
MATT|21|2|dicens eis: " Ite in castellum, quod contra vos est, et statim invenietis asinam alligatam et pullum cum ea; solvite et adducite mihi.
MATT|21|3|Et si quis vobis aliquid dixerit, dicite: "Dominus eos necessarios habet", et confestim dimittet eos ".
MATT|21|4|Hoc autem factum est, ut impleretur, quod dictum est per prophetam dicentem:
MATT|21|5|" Dicite filiae Sion:Ecce Rex tuus venit tibi,mansuetus et sedens super asinamet super pullum filium subiugalis ".
MATT|21|6|Euntes autem discipuli fecerunt, sicut praecepit illis Iesus,
MATT|21|7|et adduxerunt asinam et pullum; et imposuerunt super eis vestimenta sua, et sedit super ea.
MATT|21|8|Plurima autem turba straverunt vestimenta sua in via; alii autem caedebant ramos de arboribus et sternebant in via.
MATT|21|9|Turbae autem, quae praecedebant eum et quae sequebantur, clamabant dicentes: " Hosanna filio David! Benedictus, qui venit in nomine Domini! Hosanna in altissimis! ".
MATT|21|10|Et cum intrasset Hierosolymam, commota est universa civitas dicens: " Quis est hic?".
MATT|21|11|Turbae autem dicebant: " Hic est Iesus propheta a Nazareth Galilaeae ".
MATT|21|12|Et intravit Iesus in templum et eiciebat omnes vendentes et ementes in templo, et mensas nummulariorum evertit et cathedras vendentium columbas,
MATT|21|13|et dicit eis: " Scriptum est: "Domus mea domus orationis vocabitur". Vos autem facitis eam speluncam latronum ".
MATT|21|14|Et accesserunt ad eum caeci et claudi in templo, et sanavit eos.
MATT|21|15|Videntes autem principes sacerdotum et scribae mirabilia, quae fecit, et pueros clamantes in templo et dicentes: " Hosanna filio David ", indignati sunt
MATT|21|16|et dixerunt ei: " Audis quid isti dicant? ". Iesus autem dicit eis: " Utique; numquam legistis: "Ex ore infantium et lactantium perfecisti laudem"? ".
MATT|21|17|Et relictis illis, abiit foras extra civitatem in Bethaniam ibique mansit.
MATT|21|18|Mane autem revertens in civitatem, esuriit.
MATT|21|19|Et videns fici arborem unam secus viam, venit ad eam; et nihil invenit in ea nisi folia tantum et ait illi: " Numquam ex te fructus nascatur in sempiternum ". Et arefacta est continuo ficulnea.
MATT|21|20|Et videntes discipuli mirati sunt dicentes: " Quomodo continuo aruit ficulnea? ".
MATT|21|21|Respondens autem Iesus ait eis: " Amen dico vobis: Si habueritis fidem et non haesitaveritis, non solum de ficulnea facietis, sed et si monti huic dixeritis: "Tolle et iacta te in mare", fiet.
MATT|21|22|Et omnia, quaecumque petieritis in oratione credentes, accipietis ".
MATT|21|23|Et cum venisset in templum, accesserunt ad eum docentem principes sacerdotum et seniores populi dicentes: " In qua potestate haec facis? Et quis tibi dedit hanc potestatem? ".
MATT|21|24|Respondens autem Iesus dixit illis: " Interrogabo vos et ego unum sermonem, quem si dixeritis mihi, et ego vobis dicam, in qua potestate haec facio:
MATT|21|25|Baptismum Ioannis unde erat? A caelo an ex hominibus? ". At illi cogitabant inter se dicentes: " Si dixerimus: "E caelo", dicet nobis: Quare ergo non credidistis illi?";
MATT|21|26|si autem dixerimus: "Ex hominibus", timemus turbam; omnes enim habent Ioannem sicut prophetam ".
MATT|21|27|Et respondentes Iesu dixerunt: " Nescimus ". Ait illis et ipse: " Nec ego dico vobis in qua potestate haec facio ".
MATT|21|28|" Quid autem vobis videtur? Homo quidam habebat duos filios. Et accedens ad primum dixit: "Fili, vade hodie, operare in vinea".
MATT|21|29|Ille autem respondens ait: "Nolo"; postea autem paenitentia motus abiit.
MATT|21|30|Accedens autem ad alterum dixit similiter. At ille respondens ait: "Eo, domine"; et non ivit.
MATT|21|31|Quis ex duobus fecit voluntatem patris? ". Dicunt: " Primus ". Dicit illis Iesus: " Amen dico vobis: Publicani et meretrices praecedunt vos in regnum Dei.
MATT|21|32|Venit enim ad vos Ioannes in via iustitiae, et non credidistis ei; publicani autem et meretrices crediderunt ei. Vos autem videntes nec paenitentiam habuistis postea, ut crederetis ei.
MATT|21|33|Aliam parabolam audite. Homo erat pater familias, qui plantavit vineam et saepem circumdedit ei et fodit in ea torcular et aedificavit turrim et locavit eam agricolis et peregre profectus est.
MATT|21|34|Cum autem tempus fructuum appropinquasset, misit servos suos ad agricolas, ut acciperent fructus eius.
MATT|21|35|Et agricolae, apprehensis servis eius, alium ceciderunt, alium occiderunt, alium vero lapidaverunt.
MATT|21|36|Iterum misit alios servos plures prioribus, et fecerunt illis similiter.
MATT|21|37|Novissime autem misit ad eos filium suum dicens: "Verebuntur filium meum".
MATT|21|38|Agricolae autem videntes filium dixerunt intra se: "Hic est heres. Venite, occidamus eum et habebimus hereditatem eius".
MATT|21|39|Et apprehensum eum eiecerunt extra vineam et occiderunt.
MATT|21|40|Cum ergo venerit dominus vineae, quid faciet agricolis illis? ".
MATT|21|41|Aiunt illi: " Malos male perdet et vineam locabit aliis agricolis, qui reddant ei fructum temporibus suis ".
MATT|21|42|Dicit illis Iesus: " Numquam legistis in Scripturis:Lapidem quem reprobaverunt aedificantes,hic factus est in caput anguli;a Domino factum est istudet est mirabile in oculis nostris"?
MATT|21|43|Ideo dico vobis quia auferetur a vobis regnum Dei et dabitur genti facienti fructus eius.
MATT|21|44|Et, qui ceciderit super lapidem istum confringetur; super quem vero ceciderit, conteret eum ".
MATT|21|45|Et cum audissent principes sacerdotum et pharisaei parabolas eius, cognoverunt quod de ipsis diceret;
MATT|21|46|et quaerentes eum tenere, timuerunt turbas, quoniam sicut prophetam eum habebant.
MATT|22|1|Et respondens Iesus dixit ite rum in parabolis eis dicens:
MATT|22|2|" Simile factum est regnum caelorum homini regi, qui fecit nuptias filio suo.
MATT|22|3|Et misit servos suos vocare invitatos ad nuptias, et nolebant venire.
MATT|22|4|Iterum misit alios servos dicens: "Dicite invitatis: Ecce prandium meum paravi, tauri mei et altilia occisa, et omnia parata; venite ad nuptias".
MATT|22|5|Illi autem neglexerunt et abierunt, alius in villam suam, alius vero ad negotiationem suam;
MATT|22|6|reliqui vero tenuerunt servos eius et contumelia affectos occiderunt.
MATT|22|7|Rex autem iratus est et, missis exercitibus suis, perdidit homicidas illos et civitatem illorum succendit.
MATT|22|8|Tunc ait servis suis: "Nuptiae quidem paratae sunt, sed qui invitati erant, non fuerunt digni;
MATT|22|9|ite ergo ad exitus viarum, et quoscumque inveneritis, vocate ad nuptias".
MATT|22|10|Et egressi servi illi in vias, congregaverunt omnes, quos invenerunt, malos et bonos; et impletae sunt nuptiae discumbentium.
MATT|22|11|Intravit autem rex, ut videret discumbentes, et vidit ibi hominem non vestitum veste nuptiali
MATT|22|12|et ait illi: "Amice, quomodo huc intrasti, non habens vestem nuptialem?". At ille obmutuit.
MATT|22|13|Tunc dixit rex ministris: "Ligate pedes eius et manus et mittite eum in tenebras exteriores: ibi erit fletus et stridor dentium".
MATT|22|14|Multi enim sunt vocati, pauci vero electi ".
MATT|22|15|Tunc abeuntes pharisaei consilium inierunt, ut caperent eum in sermone.
MATT|22|16|Et mittunt ei discipulos suos cum herodianis dicentes: " Magister, scimus quia verax es et viam Dei in veritate doces, et non est tibi cura de aliquo; non enim respicis personam hominum.
MATT|22|17|Dic ergo nobis quid tibi videatur: Licet censum dare Caesari an non? ".
MATT|22|18|Cognita autem Iesus nequitia eorum, ait: " Quid me tentatis, hypocritae?
MATT|22|19|Ostendite mihi nomisma census ". At illi obtulerunt ei denarium.
MATT|22|20|Et ait illis: " Cuius est imago haec et suprascriptio? ".
MATT|22|21|Dicunt ei: " Caesaris ". Tunc ait illis: " Reddite ergo, quae sunt Caesaris, Caesari et, quae sunt Dei, Deo ".
MATT|22|22|Et audientes mirati sunt et, relicto eo, abierunt.
MATT|22|23|In illo die accesserunt ad eum sadducaei, qui dicunt non esse resurrectionem, et interrogaverunt eum
MATT|22|24|dicentes: " Magister, Moyses dixit, si quis mortuus fuerit non habens filios, ut ducat frater eius uxorem illius et suscitet semen fratri suo.
MATT|22|25|Erant autem apud nos septem fratres: et primus, uxore ducta, defunctus est et non habens semen reliquit uxorem suam fratri suo;
MATT|22|26|similiter secundus et tertius usque ad septimum.
MATT|22|27|Novissime autem omnium mulier defuncta est.
MATT|22|28|In resurrectione ergo cuius erit de septem uxor? Omnes enim habuerunt eam ".
MATT|22|29|Respondens autem Iesus ait illis: " Erratis nescientes Scripturas neque virtutem Dei;
MATT|22|30|in resurrectione enim neque nubent neque nubentur, sed sunt sicut angeli in caelo.
MATT|22|31|De resurrectione autem mortuorum non legistis, quod dictum est vobis a Deo dicente:
MATT|22|32|"Ego sum Deus Abraham et Deus Isaac et Deus Iacob"? Non est Deus mortuorum sed viventium ".
MATT|22|33|Et audientes turbae mirabantur in doctrina eius.
MATT|22|34|Pharisaei autem audientes quod silentium imposuisset sadducaeis, convenerunt in unum.
MATT|22|35|Et interrogavit unus ex eis legis doctor tentans eum:
MATT|22|36|" Magister, quod est mandatum magnum in Lege? ".
MATT|22|37|Ait autem illi: " Diliges Dominum Deum tuum in toto corde tuo et in tota anima tua et in tota mente tua:
MATT|22|38|hoc est magnum et primum mandatum.
MATT|22|39|Secundum autem simile est huic: Diliges proximum tuum sicut teipsum.
MATT|22|40|In his duobus mandatis universa Lex pendet et Prophetae ".
MATT|22|41|Congregatis autem pharisaeis, interrogavit eos Iesus
MATT|22|42|dicens: " Quid vobis videtur de Christo? Cuius filius est? ". Dicunt ei: " David ".
MATT|22|43|Ait illis: " Quomodo ergo David in Spiritu vocat eum Dominum dicens:
MATT|22|44|"Dixit Dominus Domino meo: Sede a dextris meis,donec ponam inimicos tuos sub pedibus tuis"?
MATT|22|45|Si ergo David vocat eum Dominum, quomodo filius eius est? ".
MATT|22|46|Et nemo poterat respondere ei verbum, neque ausus fuit quisquam ex illa die eum amplius interrogare.
MATT|23|1|Tunc Iesus locutus est ad turbas et ad discipulos suos
MATT|23|2|dicens: " Super cathedram Moysis sederunt scribae et pharisaei.
MATT|23|3|Omnia ergo, quaecumque dixerint vobis, facite et servate; secundum opera vero eorum nolite facere: dicunt enim et non faciunt.
MATT|23|4|Alligant autem onera gravia et importabilia et imponunt in umeros hominum, ipsi autem digito suo nolunt ea movere.
MATT|23|5|Omnia vero opera sua faciunt, ut videantur ab hominibus: dilatant enim phylacteria sua et magnificant fimbrias,
MATT|23|6|amant autem primum recubitum in cenis et primas cathedras in synagogis
MATT|23|7|et salutationes in foro et vocari ab hominibus Rabbi.
MATT|23|8|Vos autem nolite vocari Rabbi; unus enim est Magister vester, omnes autem vos fratres estis.
MATT|23|9|Et Patrem nolite vocare vobis super terram, unus enim est Pater vester, caelestis.
MATT|23|10|Nec vocemini Magistri, quia Magister vester unus est, Christus.
MATT|23|11|Qui maior est vestrum, erit minister vester.
MATT|23|12|Qui autem se exaltaverit, humiliabitur; et, qui se humiliaverit, exaltabitur.
MATT|23|13|Vae autem vobis, scribae et pharisaei hypocritae, quia clauditis regnum caelorum ante homines! Vosenim non intratis nec introeuntes sinitis intrare.
MATT|23|14|()
MATT|23|15|Vae vobis, scribae et pharisaei hypocritae, quia circuitis mare et aridam, ut faciatis unum proselytum, et cum fuerit factus, facitis eum filium gehennae duplo quam vos!
MATT|23|16|Vae vobis, duces caeci, qui dicitis: "Quicumque iuraverit per templum, nihil est; quicumque autem iuraverit in auro templi, debet".
MATT|23|17|Stulti et caeci! Quid enim maius est: aurum an templum, quod sanctificat aurum?
MATT|23|18|Et: "Quicumque iuraverit in altari, nihil est; quicumque autem iuraverit in dono, quod est super illud, debet".
MATT|23|19|Caeci! Quid enim maius est: donum an altare, quod sanctificat donum?
MATT|23|20|Qui ergo iuraverit in altari, iurat in eo et in omnibus, quae super illud sunt;
MATT|23|21|et, qui iuraverit in templo, iurat in illo et in eo, qui inhabitat in ipso;
MATT|23|22|et, qui iuraverit in caelo, iurat in throno Dei et in eo, qui sedet super eum.
MATT|23|23|Vae vobis, scribae et pharisaei hypocritae, quia decimatis mentam et anethum et cyminum et reliquistis, quae graviora sunt legis: iudicium et misericordiam et fidem! Haec oportuit facere et illa non omittere.
MATT|23|24|Duces caeci, excolantes culicem, camelum autem glutientes.
MATT|23|25|Vae vobis, scribae et pharisaei hypocritae, quia mundatis, quod de foris est calicis et paropsidis, intus autem pleni sunt rapina et immunditia!
MATT|23|26|Pharisaee caece, munda prius, quod intus est calicis, ut fiat et id, quod de foris eius est, mundum.
MATT|23|27|Vae vobis, scribae et pharisaei hypocritae, quia similes estis sepulcris dealbatis, quae a foris quidem parent speciosa, intus vero plena sunt ossibus mortuorum et omni spurcitia!
MATT|23|28|Sic et vos a foris quidem paretis hominibus iusti, intus autem pleni estis hypocrisi et iniquitate.
MATT|23|29|Vae vobis, scribae et pharisaei hypocritae, qui aedificatis sepulcra prophetarum et ornatis monumenta iustorum
MATT|23|30|et dicitis: "Si fuissemus in diebus patrum nostrorum, non essemus socii eorum in sanguine prophetarum"!
MATT|23|31|Itaque testimonio estis vobismetipsis quia filii estis eorum, qui prophetas occiderunt.
MATT|23|32|Et vos implete mensuram patrum vestrorum.
MATT|23|33|Serpentes, genimina viperarum, quomodo fugietis a iudicio gehennae?
MATT|23|34|Ideo ecce ego mitto ad vos prophetas et sapientes et scribas; ex illis occidetis et crucifigetis et ex eis flagellabitis in synagogis vestris et persequemini de civitate in civitatem,
MATT|23|35|ut veniat super vos omnis sanguis iustus, qui effusus est super terram a sanguine Abel iusti usque ad sanguinem Zachariae filii Barachiae, quem occidistis inter templum et altare.
MATT|23|36|Amen dico vobis: Venient haec omnia super generationem istam.
MATT|23|37|Ierusalem, Ierusalem, quae occidis prophetas et lapidas eos, qui ad te missi sunt, quotiens volui congregare filios tuos, quemadmodum gallina congregat pullos suos sub alas, et noluistis!
MATT|23|38|Ecce relinquitur vobis domus vestra deserta!
MATT|23|39|Dico enim vobis: Non me videbitis amodo, donec dicatis: "Benedictus, qui venit in nomine Dominil" ".
MATT|24|1|Et egressus Iesus de templo ibat, et accesserunt discipuli eius, ut ostenderent ei aedificationes templi;
MATT|24|2|ipse autem respondens dixit eis: " Non videtis haec omnia? Amen dico vobis: Non relinquetur hic lapis super lapidem, qui non destruetur ".
MATT|24|3|Sedente autem eo super montem Oliveti, accesserunt ad eum discipuli secreto dicentes: " Dic nobis: Quando haec erunt, et quod signum adventus tui et consummationis saeculi? ".
MATT|24|4|Et respondens Iesus dixit eis: " Videte, ne quis vos seducat.
MATT|24|5|Multi enim venient in nomine meo dicentes: "Ego sum Christus", et multos seducent.
MATT|24|6|Audituri enim estis proelia et opiniones proeliorum. Videte, ne turbemini; oportet enim fieri, sed nondum est finis.
MATT|24|7|Consurget enim gens in gentem, et regnum in regnum, et erunt fames et terrae motus per loca;
MATT|24|8|haec autem omnia initia sunt dolorum.
MATT|24|9|Tunc tradent vos in tribulationem et occident vos, et eritis odio omnibus gentibus propter nomen meum.
MATT|24|10|Et tunc scandalizabuntur multi et invicem tradent et odio habebunt invicem;
MATT|24|11|et multi pseudoprophetae surgent et seducent multos.
MATT|24|12|Et, quoniam abundavit iniquitas, refrigescet caritas multorum;
MATT|24|13|qui autem permanserit usque in finem, hic salvus erit.
MATT|24|14|Et praedicabitur hoc evangelium regni in universo orbe in testimonium omnibus gentibus; et tunc veniet consummatio.
MATT|24|15|Cum ergo videritis abominationem desolationis, quae dicta est a Daniele propheta, stantem in loco sancto, qui legit, intellegat:
MATT|24|16|tunc qui in Iudaea sunt, fugiant ad montes;
MATT|24|17|qui in tecto, non descendat tollere aliquid de domo sua;
MATT|24|18|et, qui in agro, non revertatur tollere pallium suum.
MATT|24|19|Vae autem praegnantibus et nutrientibus in illis diebus!
MATT|24|20|Orate autem, ut non fiat fuga vestra hieme vel sabbato:
MATT|24|21|erit enim tunc tribulatio magna, qualis non fuit ab initio mundi usque modo neque fiet.
MATT|24|22|Et nisi breviati fuissent dies illi, non fieret salva omnis caro; sed propter electos breviabuntur dies illi.
MATT|24|23|Tunc si quis vobis dixerit: "Ecce hic Christus" aut: "Hic", nolite credere.
MATT|24|24|Surgent enim pseudochristi et pseudoprophetae et dabunt signa magna et prodigia, ita ut in errorem inducantur, si fieri potest, etiam electi.
MATT|24|25|Ecce praedixi vobis.
MATT|24|26|Si ergo dixerint vobis: "Ecce in deserto est", nolite exire; "Ecce in penetralibus", nolite credere;
MATT|24|27|sicut enim fulgur exit ab oriente et paret usque in occidentem, ita erit adventus Filii hominis.
MATT|24|28|Ubicumque fuerit corpus, illuc congregabuntur aquilae.
MATT|24|29|Statim autem post tribulationem dierum illorum, sol obscurabitur, et luna non dabit lumen suum, et stellae cadent de caelo, et virtutes caelorum commovebuntur.
MATT|24|30|Et tunc parebit signum Filii hominis in caelo, et tunc plangent omnes tribus terrae et videbunt Filium hominis venientem in nubibus caeli cum virtute et gloria multa;
MATT|24|31|et mittet angelos suos cum tuba magna, et congregabunt electos eius a quattuor ventis, a summis caelorum usque ad terminos eorum.
MATT|24|32|Ab arbore autem fici discite parabolam: cum iam ramus eius tener fuerit, et folia nata, scitis quia prope est aestas.
MATT|24|33|Ita et vos, cum videritis haec omnia, scitote quia prope est in ianuis.
MATT|24|34|Amen dico vobis: Non praeteribit haec generatio, donec omnia haec fiant.
MATT|24|35|Caelum et terra transibunt, verba vero mea non praeteribunt.
MATT|24|36|De die autem illa et hora nemo scit, neque angeli caelorum neque Filius, nisi Pater solus.
MATT|24|37|Sicut enim dies Noe, ita erit adventus Filii hominis.
MATT|24|38|Sicut enim erant in diebus ante diluvium comedentes et bibentes, nubentes et nuptum tradentes, usque ad eum diem, quo introivit in arcam Noe,
MATT|24|39|et non cognoverunt, donec venit diluvium et tulit omnes, ita erit et adventus Filii hominis.
MATT|24|40|Tunc duo erunt in agro: unus assumitur, et unus relinquitur;
MATT|24|41|duae molentes in mola: una assumitur, et una relinquitur.
MATT|24|42|Vigilate ergo, quia nescitis qua die Dominus vester venturus sit.
MATT|24|43|Illud autem scitote quoniam si sciret pater familias qua hora fur venturus esset, vigilaret utique et non sineret perfodi domum suam.
MATT|24|44|Ideo et vos estote parati, quia, qua nescitis hora, Filius hominis venturus est.
MATT|24|45|Quis putas est fidelis servus et prudens, quem constituit dominus supra familiam suam, ut det illis cibum in tempore?
MATT|24|46|Beatus ille servus, quem cum venerit dominus eius, invenerit sic facientem.
MATT|24|47|Amen dico vobis quoniam super omnia bona sua constituet eum.
MATT|24|48|Si autem dixerit malus servus ille in corde suo: "Moram facit dominus meus venire",
MATT|24|49|et coeperit percutere conservos suos, manducet autem et bibat cum ebriis,
MATT|24|50|veniet dominus servi illius in die, qua non sperat, et in hora, qua ignorat,
MATT|24|51|et dividet eum partemque eius ponet cum hypocritis; illic erit fletus et stridor dentium.
MATT|25|1|Tunc simile erit regnum cae lorum decem virginibus, quae accipientes lampades suas exierunt obviam sponso.
MATT|25|2|Quinque autem ex eis erant fatuae, et quinque prudentes.
MATT|25|3|Fatuae enim, acceptis lampadibus suis, non sumpserunt oleum secum;
MATT|25|4|prudentes vero acceperunt oleum in vasis cum lampadibus suis.
MATT|25|5|Moram autem faciente sponso, dormitaverunt omnes et dormierunt.
MATT|25|6|Media autem nocte clamor factus est: "Ecce sponsus! Exite obviam ei".
MATT|25|7|Tunc surrexerunt omnes virgines illae et ornaverunt lampades suas.
MATT|25|8|Fatuae autem sapientibus dixerunt: "Date nobis de oleo vestro, quia lampades nostrae exstinguuntur".
MATT|25|9|Responderunt prudentes dicentes: "Ne forte non sufficiat nobis et vobis, ite potius ad vendentes et emite vobis".
MATT|25|10|Dum autem irent emere, venit sponsus, et quae paratae erant, intraverunt cum eo ad nuptias; et clausa est ianua.
MATT|25|11|Novissime autem veniunt et reliquae virgines dicentes: "Domine, domine, aperi nobis".
MATT|25|12|At ille respondens ait: "Amen dico vobis: Nescio vos".
MATT|25|13|Vigilate itaque, quia nescitis diem neque horam.
MATT|25|14|Sicut enim homo peregre proficiscens vocavit servos suos et tradidit illis bona sua.
MATT|25|15|Et uni dedit quinque talenta, alii autem duo, alii vero unum, unicuique secundum propriam virtutem, et profectus est. Statim
MATT|25|16|abiit, qui quinque talenta acceperat, et operatus est in eis et lucratus est alia quinque;
MATT|25|17|similiter qui duo acceperat, lucratus est alia duo.
MATT|25|18|Qui autem unum acceperat, abiens fodit in terra et abscondit pecuniam domini sui.
MATT|25|19|Post multum vero temporis venit dominus servorum illorum et ponit rationem cum eis.
MATT|25|20|Et accedens, qui quinque talenta acceperat, obtulit alia quinque talenta dicens: "Domine, quinque talenta tradidisti mihi; ecce alia quinque superlucratus sum".
MATT|25|21|Ait illi dominus eius: "Euge, serve bone et fidelis. Super pauca fuisti fidelis; supra multa te constituam: intra in gaudium domini tui".
MATT|25|22|Accessit autem et qui duo talenta acceperat, et ait: "Domine, duo talenta tradidisti mihi; ecce alia duo lucratus sum".
MATT|25|23|Ait illi dominus eius: "Euge, serve bone et fidelis. Super pauca fuisti fidelis; supra multa te constituam: intra in gaudium domini tui".
MATT|25|24|Accedens autem et qui unum talentum acceperat, ait: "Domine, novi te quia homo durus es: metis, ubi non seminasti, et congregas, ubi non sparsisti;
MATT|25|25|et timens abii et abscondi talentum tuum in terra. Ecce habes, quod tuum est".
MATT|25|26|Respondens autem dominus eius dixit ei: "Serve male et piger! Sciebas quia meto, ubi non seminavi, et congrego, ubi non sparsi?
MATT|25|27|Oportuit ergo te mittere pecuniam meam nummulariis, et veniens ego recepissem, quod meum est cum usura.
MATT|25|28|Tollite itaque ab eo talentum et date ei, qui habet decem talenta:
MATT|25|29|omni enim habenti dabitur, et abundabit; ei autem, qui non habet, et quod habet, auferetur ab eo.
MATT|25|30|Et inutilem servum eicite in tenebras exteriores: illic erit fletus et stridor dentium".
MATT|25|31|Cum autem venerit Filius hominis in gloria sua, et omnes angeli cum eo, tunc sedebit super thronum gloriae suae.
MATT|25|32|Et congregabuntur ante eum omnes gentes; et separabit eos ab invicem, sicut pastor segregat oves ab haedis,
MATT|25|33|et statuet oves quidem a dextris suis, haedos autem a sinistris.
MATT|25|34|Tunc dicet Rex his, qui a dextris eius erunt: "Venite, benedicti Patris mei; possidete paratum vobis regnum a constitutione mundi.
MATT|25|35|Esurivi enim, et dedistis mihi manducare; sitivi, et dedistis mihi bibere; hospes eram, et collegistis me;
MATT|25|36|nudus, et operuistis me; infirmus, et visitastis me; in carcere eram, et venistis ad me".
MATT|25|37|Tunc respondebunt ei iusti dicentes: "Domine, quando te vidimus esurientem et pavimus, aut sitientem et dedimus tibi potum?
MATT|25|38|Quando autem te vidimus hospitem et collegimus, aut nudum et cooperuimus?
MATT|25|39|Quando autem te vidimus infirmum aut in carcere et venimus ad te?".
MATT|25|40|Et respondens Rex dicet illis: "Amen dico vobis: Quamdiu fecistis uni de his fratribus meis minimis, mihi fecistis".
MATT|25|41|Tunc dicet et his, qui a sinistris erunt: "Discedite a me, maledicti, in ignem aeternum, qui praeparatus est Diabolo et angelis eius.
MATT|25|42|Esurivi enim, et non dedistis mihi manducare; sitivi, et non dedistis mihi potum;
MATT|25|43|hospes eram, et non collegistis me; nudus, et non operuistis me; infirmus et in carcere, et non visitastis me".
MATT|25|44|Tunc respondebunt et ipsi dicentes: "Domine, quando te vidimus esurientem aut sitientem aut hospitem aut nudum aut infirmum vel in carcere et non ministravimus tibi?".
MATT|25|45|Tunc respondebit illis dicens: "Amen dico vobis: Quamdiu non fecistis uni de minimis his, nec mihi fecistis".
MATT|25|46|Et ibunt hi in supplicium aeternum, iusti autem in vitam aeternam ".
MATT|26|1|Et factum est, cum consum masset Iesus sermones hos omnes, dixit discipulis suis:
MATT|26|2|" Scitis quia post biduum Pascha fiet, et Filius hominis traditur, ut crucifigatur ".
MATT|26|3|Tunc congregati sunt principes sacerdotum et seniores populi in aulam principis sacerdotum, qui dicebatur Caiphas,
MATT|26|4|et consilium fecerunt, ut Iesum dolo tenerent et occiderent;
MATT|26|5|dicebant autem: " Non in die festo, ne tumultus fiat in populo ".
MATT|26|6|Cum autem esset Iesus in Bethania, in domo Simonis leprosi,
MATT|26|7|accessit ad eum mulier habens alabastrum unguenti pretiosi et effudit super caput ipsius recumbentis.
MATT|26|8|Videntes autem discipuli, indignati sunt dicentes: " Ut quid perditio haec?
MATT|26|9|Potuit enim istud venumdari multo et dari pauperibus ".
MATT|26|10|Sciens autem Iesus ait illis: " Quid molesti estis mulieri? Opus enim bonum operata est in me;
MATT|26|11|nam semper pauperes habetis vobiscum, me autem non semper habetis.
MATT|26|12|Mittens enim haec unguentum hoc supra corpus meum, ad sepeliendum me fecit.
MATT|26|13|Amen dico vobis: Ubicumque praedicatum fuerit hoc evangelium in toto mundo, dicetur et quod haec fecit in memoriam eius ".
MATT|26|14|Tunc abiit unus de Duodecim, qui dicebatur Iudas Iscariotes, ad principes sacerdotum
MATT|26|15|et ait: " Quid vultis mihi dare, et ego vobis eum tradam? ". At illi constituerunt ei triginta argenteos.
MATT|26|16|Et exinde quaerebat opportunitatem, ut eum traderet.
MATT|26|17|Prima autem Azymorum accesserunt discipuli ad Iesum dicentes: " Ubi vis paremus tibi comedere Pascha? ".
MATT|26|18|Ille autem dixit: " Ite in civitatem ad quendam et dicite ei: "Magister dicit: Tempus meum prope est; apud te facio Pascha cum discipulis meis" ".
MATT|26|19|Et fecerunt discipuli, sicut constituit illis Iesus, et paraverunt Pascha.
MATT|26|20|Vespere autem facto, discumbebat cum Duodecim.
MATT|26|21|Et edentibus illis, dixit: " Amen dico vobis: Unus vestrum me traditurus est ".
MATT|26|22|Et contristati valde, coeperunt singuli dicere ei: " Numquid ego sum, Domine? ".
MATT|26|23|At ipse respondens ait: " Qui intingit mecum manum in paropside, hic me tradet.
MATT|26|24|Filius quidem hominis vadit, sicut scriptum est de illo; vae autem homini illi, per quem Filius hominis traditur! Bonum erat ei, si natus non fuisset homo ille ".
MATT|26|25|Respondens autem Iudas, qui tradidit eum, dixit: " Numquid ego sum, Rabbi? ". Ait illi: " Tu dixisti ".
MATT|26|26|Cenantibus autem eis, accepit Iesus panem et benedixit ac fregit deditque discipulis et ait: " Accipite, comedite: hoc est corpus meum ".
MATT|26|27|Et accipiens calicem, gratias egit et dedit illis dicens: " Bibite ex hoc omnes:
MATT|26|28|hic est enim sanguis meus novi testamenti, qui pro multis effunditur in remissionem peccatorum.
MATT|26|29|Dico autem vobis: Non bibam amodo de hoc genimine vitis usque in diem illum, cum illud bibam vobiscum novum in regno Patris mei ".
MATT|26|30|Et hymno dicto, exierunt in montem Oliveti.
MATT|26|31|Tunc dicit illis Iesus: " Omnes vos scandalum patiemini in me in ista nocte. Scriptum est enim: "Percutiam pastorem, et dispergentur oves gregis".
MATT|26|32|Postquam autem resurrexero, praecedam vos in Galilaeam ".
MATT|26|33|Respondens autem Petrus ait illi: " Et si omnes scandalizati fuerint in te, ego numquam scandalizabor ".
MATT|26|34|Ait illi Iesus: " Amen dico tibi: In hac nocte, antequam gallus cantet, ter me negabis ".
MATT|26|35|Ait illi Petrus: " Etiam si oportuerit me mori tecum, non te negabo ". Similiter et omnes discipuli dixerunt.
MATT|26|36|Tunc venit Iesus cum illis in praedium, quod dicitur Gethsemani. Et dicit discipulis: " Sedete hic, donec vadam illuc et orem ".
MATT|26|37|Et assumpto Petro et duobus filiis Zebedaei, coepit contristari et maestus esse.
MATT|26|38|Tunc ait illis: " Tristis est anima mea usque ad mortem; sustinete hic et vigilate mecum ".
MATT|26|39|Et progressus pusillum, procidit in faciem suam orans et dicens: " Pater mi, si possibile est, transeat a me calix iste; verumtamen non sicut ego volo, sed sicut tu ".
MATT|26|40|Et venit ad discipulos et invenit eos dormientes; et dicit Petro: " Sic non potuistis una hora vigilare mecum?
MATT|26|41|Vigilate et orate, ut non intretis in tentationem; spiritus quidem promptus est, caro autem infirma ".
MATT|26|42|Iterum secundo abiit et oravit dicens: " Pater mi, si non potest hoc transire, nisi bibam illud, fiat voluntas tua ".
MATT|26|43|Et venit iterum et invenit eos dormientes: erant enim oculi eorum gravati.
MATT|26|44|Et relictis illis, iterum abiit et oravit tertio, eundem sermonem iterum dicens.
MATT|26|45|Tunc venit ad discipulos et dicit illis: " Dormite iam et requiescite; ecce appropinquavit hora, et Filius hominis traditur in manus peccatorum.
MATT|26|46|Surgite, eamus; ecce appropinquavit, qui me tradit ".
MATT|26|47|Et adhuc ipso loquente, ecce Iudas, unus de Duodecim, venit, et cum eo turba multa cum gladiis et fustibus, missi a principibus sacerdotum et senioribus populi.
MATT|26|48|Qui autem tradidit eum, dedit illis signum dicens: " Quemcumque osculatus fuero, ipse est; tenete eum! ".
MATT|26|49|Et confestim accedens ad Iesum dixit: " Ave, Rabbi! " et osculatus est eum.
MATT|26|50|Iesus autem dixit illi: " Amice, ad quod venisti! ". Tunc accesserunt et manus iniecerunt in Iesum et tenuerunt eum.
MATT|26|51|Et ecce unus ex his, qui erant cum Iesu, extendens manum exemit gladium suum et percutiens servum principis sacerdotum amputavit auriculam eius.
MATT|26|52|Tunc ait illi Iesus: " Converte gladium tuum in locum suum. Omnes enim, qui acceperint gladium, gladio peribunt.
MATT|26|53|An putas quia non possum rogare Patrem meum, et exhibebit mihi modo plus quam duodecim legiones angelorum?
MATT|26|54|Quomodo ergo implebuntur Scripturae quia sic oportet fieri? ".
MATT|26|55|In illa hora dixit Iesus turbis: " Tamquam ad latronem existis cum gladiis et fustibus comprehendere me? Cotidie sedebam docens in templo, et non me tenuistis ".
MATT|26|56|Hoc autem totum factum est, ut implerentur scripturae Prophetarum. Tunc discipuli omnes, relicto eo, fugerunt.
MATT|26|57|Illi autem tenentes Iesum duxerunt ad Caipham principem sacerdotum, ubi scribae et seniores convenerant.
MATT|26|58|Petrus autem sequebatur eum a longe usque in aulam principis sacerdotum; et ingressus intro sede bat cum ministris, ut videret finem.
MATT|26|59|Principes autem sacerdotum et omne concilium quaerebant falsum testimonium contra Iesum, ut eum morti traderent,
MATT|26|60|et non invenerunt, cum multi falsi testes accessissent. Novissime autem venientes duo
MATT|26|61|dixerunt: " Hic dixit: "Possum destruere templum Dei et post triduum aedificare illud" ".
MATT|26|62|Et surgens princeps sacerdotum ait illi: " Nihil respondes? Quid isti adversum te testificantur? ".
MATT|26|63|Iesus autem tacebat. Et princeps sacerdotum ait illi: " Adiuro te per Deum vivum, ut dicas nobis, si tu es Christus Filius Dei ".
MATT|26|64|Dicit illi Iesus: " Tu dixisti. Verumtamen dico vobis: Amodo videbitis Filium hominis sedentem a dextris Virtutis et venientem in nubibus caeli.
MATT|26|65|Tunc princeps sacerdotum scidit vestimenta sua dicens: " Blasphemavit! Quid adhuc egemus testibus? Ecce nunc audistis blasphemiam.
MATT|26|66|Quid vobis videtur? ". Illi autem respondentes dixerunt: " Reus est mortis! ".
MATT|26|67|Tunc exspuerunt in faciem eius et colaphis eum ceciderunt; alii autem palmas in faciem ei dederunt
MATT|26|68|dicentes: " Prophetiza nobis, Christe: Quis est, qui te percussit? ".
MATT|26|69|Petrus vero sedebat foris in atrio; et accessit ad eum una ancilla dicens: " Et tu cum Iesu Galilaeo eras! ".
MATT|26|70|At ille negavit coram omnibus dicens: " Nescio quid dicis! ".
MATT|26|71|Exeunte autem illo ad ianuam, vidit eum alia et ait his, qui erant ibi: Hic erat cum Iesu Nazareno! ".
MATT|26|72|Et iterum negavit cum iuramento: " Non novi hominem! ".
MATT|26|73|Post pusillum autem accesserunt, qui stabant, et dixerunt Petro: " Vere et tu ex illis es, nam et loquela tua manifestum te facit ".
MATT|26|74|Tunc coepit detestari et iurare: " Non novi hominem! ". Et continuo gallus cantavit;
MATT|26|75|et recordatus est Petrus verbi Iesu, quod dixerat: " Priusquam gallus cantet, ter me negabis ". Et egressus foras ploravit amare.
MATT|27|1|Mane autem facto, consi lium inierunt omnes princi pes sacerdotum et seniores populi adversus Iesum, ut eum morti traderent.
MATT|27|2|Et vinctum adduxerunt eum et tradiderunt Pilato praesidi.
MATT|27|3|Tunc videns Iudas, qui eum tradidit, quod damnatus esset, paenitentia ductus, rettulit triginta argenteos principibus sacerdotum et senioribus
MATT|27|4|dicens: " Peccavi tradens sanguinem innocentem ". At illi dixerunt: " Quid ad nos? Tu videris! ".
MATT|27|5|Et proiectis argenteis in templo, recessit et abiens laqueo se suspendit.
MATT|27|6|Principes autem sacerdotum, acceptis argenteis, dixerunt: " Non licet mittere eos in corbanam, quia pretium sanguinis est ".
MATT|27|7|Consilio autem inito, emerunt ex illis agrum Figuli in sepulturam peregrinorum.
MATT|27|8|Propter hoc vocatus est ager ille ager Sanguinis usque in hodiernum diem.
MATT|27|9|Tunc impletum est quod dictum est per Ieremiam prophetam di centem: " Et acceperunt triginta argenteos, pretium appretiati quem appretiaverunt a filiis Israel,
MATT|27|10|et dederunt eos in agrum Figuli, sicut constituit mihi Dominus ".
MATT|27|11|Iesus autem stetit ante praesidem; et interrogavit eum praeses dicens: Tu es Rex Iudaeorum? ". Dixit autem Iesus: " Tu dicis ".
MATT|27|12|Et cum accusaretur a principibus sacerdotum et senioribus, nihil respondit.
MATT|27|13|Tunc dicit illi Pilatus: " Non audis quanta adversum te dicant testimonia? ".
MATT|27|14|Et non respondit ei ad ullum verbum, ita ut miraretur praeses vehementer.
MATT|27|15|Per diem autem sollemnem consueverat praeses dimittere turbae unum vinctum, quem voluissent.
MATT|27|16|Habebant autem tunc vinctum insignem, qui dicebatur Barabbas.
MATT|27|17|Congregatis ergo illis dixit Pilatus: " Quem vultis dimittam vobis: Barabbam an Iesum, qui dicitur Christus? ".
MATT|27|18|Sciebat enim quod per invidiam tradidissent eum.
MATT|27|19|Sedente autem illo pro tribunali, misit ad illum uxor eius dicens: " Nihil tibi et iusto illi. Multa enim passa sum hodie per visum propter eum.
MATT|27|20|Principes autem sacerdotum et seniores persuaserunt turbis, ut peterent Barabbam, Iesum vero perderent.
MATT|27|21|Respondens autem praeses ait illis: " Quem vultis vobis de duobus dimittam? ". At illi dixerunt: " Barabbam! ".
MATT|27|22|Dicit illis Pilatus: " Quid igitur faciam de Iesu, qui dicitur Christus? ". Dicunt omnes: " Crucifigatur! ".
MATT|27|23|Ait autem: " Quid enim mali fecit? ". At illi magis clamabant dicentes: Crucifigatur! ".
MATT|27|24|Videns autem Pilatus quia nihil proficeret, sed magis tumultus fieret, accepta aqua, lavit manus coram turba dicens: " Innocens ego sum a sanguine hoc; vos videritis! ".
MATT|27|25|Et respondens universus populus dixit: " Sanguis eius super nos et super filios nostros ".
MATT|27|26|Tunc dimisit illis Barabbam; Iesum autem flagellatum tradidit, ut crucifigeretur.
MATT|27|27|Tunc milites praesidis suscipientes Iesum in praetorio congregaverunt ad eum universam cohortem.
MATT|27|28|Et exuentes eum, clamydem coccineam circumdederunt ei
MATT|27|29|et plectentes coronam de spinis posuerunt super caput eius et arundinem in dextera eius et, genu flexo ante eum, illudebant ei dicentes: " Ave, rex Iudaeorum! ".
MATT|27|30|Et exspuentes in eum acceperunt arundinem et percutiebant caput eius.
MATT|27|31|Et postquam illuserunt ei, exuerunt eum clamyde et induerunt eum vestimentis eius et duxerunt eum, ut crucifigerent.
MATT|27|32|Exeuntes autem invenerunt hominem Cyrenaeum nomine Simonem; hunc angariaverunt, ut tolleret crucem eius.
MATT|27|33|Et venerunt in locum, qui dicitur Golgotha, quod est Calvariae locus,
MATT|27|34|et dederunt ei vinum bibere cum felle mixtum; et cum gustasset, noluit bibere.
MATT|27|35|Postquam autem crucifixerunt eum, diviserunt vestimenta eius sortem mittentes
MATT|27|36|et sedentes servabant eum ibi.
MATT|27|37|Et imposuerunt super caput eius causam ipsius scriptam: " Hic est Iesus Rex Iudaeorum ".
MATT|27|38|Tunc crucifiguntur cum eo duo latrones: unus a dextris, et unus a sinistris.
MATT|27|39|Praetereuntes autem blasphemabant eum moventes capita sua
MATT|27|40|et dicentes: " Qui destruis templum et in triduo illud reaedificas, salva temetipsum; si Filius Dei es, descende de cruce! ".
MATT|27|41|Similiter et principes sacerdotum illudentes cum scribis et senioribus dicebant:
MATT|27|42|" Alios salvos fecit, seipsum non potest salvum facere. Rex Israel est; descendat nunc de cruce, et credemus in eum.
MATT|27|43|Confidit in Deo; liberet nunc, si vult eum. Dixit enim: "Dei Filius sum" ".
MATT|27|44|Idipsum autem et latrones, qui crucifixi erant cum eo, improperabant ei.
MATT|27|45|A sexta autem hora tenebrae factae sunt super universam terram usque ad horam nonam.
MATT|27|46|Et circa horam nonam clamavit Iesus voce magna dicens: " Eli, Eli, lema sabacthani? ", hoc est: " Deus meus, Deus meus, ut quid dereliquisti me?.
MATT|27|47|Quidam autem ex illic stantibus audientes dicebant: " Eliam vocat iste.
MATT|27|48|Et continuo currens unus ex eis acceptam spongiam implevit aceto et imposuit arundini et dabat ei bibere.
MATT|27|49|Ceteri vero dicebant: " Sine, videamus an veniat Elias liberans eum ".
MATT|27|50|Iesus autem iterum clamans voce magna emisit spiritum.
MATT|27|51|Et ecce velum templi scissum est a summo usque deorsum in duas partes, et terra mota est, et petrae scissae sunt;
MATT|27|52|et monumenta aperta sunt, et multa corpora sanctorum, qui dormierant, surrexerunt
MATT|27|53|et exeuntes de monumentis post resurrectionem eius venerunt in sanctam civitatem et apparuerunt multis.
MATT|27|54|Centurio autem et, qui cum eo erant custodientes Iesum, viso terrae motu et his, quae fiebant, timuerunt valde dicentes: " Vere Dei Filius erat iste! ".
MATT|27|55|Erant autem ibi mulieres multae a longe aspicientes, quae secutae erant Iesum a Galilaea ministrantes ei;
MATT|27|56|inter quas erat Maria Magdalene et Maria Iacobi et Ioseph mater et mater filiorum Zebedaei.
MATT|27|57|Cum sero autem factum esset, venit homo dives ab Arimathaea nomine Ioseph, qui et ipse discipulus erat Iesu.
MATT|27|58|Hic accessit ad Pilatum et petiit corpus Iesu. Tunc Pilatus iussit reddi.
MATT|27|59|Et accepto corpore, Ioseph involvit illud in sindone munda
MATT|27|60|et posuit illud in monumento suo novo, quod exciderat in petra, et advolvit saxum magnum ad ostium monumenti et abiit.
MATT|27|61|Erat autem ibi Maria Magdalene et altera Maria sedentes contra sepulcrum.
MATT|27|62|Altera autem die, quae est post Parascevem, convenerunt principes sacerdotum et pharisaei ad Pilatum
MATT|27|63|dicentes: " Domine, recordati sumus quia seductor ille dixit adhuc vivens: "Post tres dies resurgam".
MATT|27|64|Iube ergo custodiri sepulcrum usque in diem tertium, ne forte veniant discipuli eius et furentur eum et dicant plebi: "Surrexit a mortuis", et erit novissimus error peior priore ".
MATT|27|65|Ait illis Pilatus: " Habetis custodiam; ite, custodite, sicut scitis ".
MATT|27|66|Illi autem abeuntes munierunt sepulcrum, signantes lapidem, cum custodia.
MATT|28|1|Sero autem post sabbatum, cum illucesceret in primam sabbati, venit Maria Magdalene et altera Maria videre sepulcrum.
MATT|28|2|Et ecce terrae motus factus est magnus: angelus enim Domini descendit de caelo et accedens revolvit lapidem et sedebat super eum.
MATT|28|3|Erat autem aspectus eius sicut fulgur, et vestimentum eius candidum sicut nix.
MATT|28|4|Prae timore autem eius exterriti sunt custodes et facti sunt velut mortui.
MATT|28|5|Respondens autem angelus dixit mulieribus: " Nolite timere vos! Scio enim quod Iesum, qui crucifixus est, quaeritis.
MATT|28|6|Non est hic: surrexit enim, sicut dixit. Venite, videte locum, ubi positus erat.
MATT|28|7|Et cito euntes dicite discipulis eius: "Surrexit a mortuis et ecce praecedit vos in Galilaeam; ibi eum videbitis". Ecce dixi vobis ".
MATT|28|8|Et exeuntes cito de monumento cum timore et magno gaudio cucurrerunt nuntiare discipulis eius.
MATT|28|9|Et ecce Iesus occurrit illis dicens: " Avete ". Illae autem accesserunt et tenuerunt pedes eius et adoraverunt eum.
MATT|28|10|Tunc ait illis Iesus: " Nolite timere; ite, nuntiate fratribus meis, ut eant in Galilaeam et ibi me videbunt ".
MATT|28|11|Quae cum abiissent, ecce quidam de custodia venerunt in civitatem et nuntiaverunt principibus sacerdotum omnia, quae facta fuerant.
MATT|28|12|Et congregati cum senioribus, consilio accepto, pecuniam copiosam dederunt militibus
MATT|28|13|dicentes: " Dicite: "Discipuli eius nocte venerunt et furati sunt eum, nobis dormientibus".
MATT|28|14|Et si hoc auditum fuerit a praeside, nos suadebimus ei et securos vos faciemus ".
MATT|28|15|At illi, accepta pecunia, fecerunt, sicut erant docti. Et divulgatum est verbum istud apud Iudaeos usque in hodiernum diem.
MATT|28|16|Undecim autem discipuli abierunt in Galilaeam, in montem ubi constituerat illis Iesus,
MATT|28|17|et videntes eum adoraverunt; quidam autem dubitaverunt.
MATT|28|18|Et accedens Iesus locutus est eis dicens: " Data est mihi omnis potestas in caelo et in terra.
MATT|28|19|Euntes ergo docete omnes gentes, baptizantes eos in nomine Patris et Filii et Spiritus Sancti,
MATT|28|20|docentes eos servare omnia, quaecumque mandavi vobis. Et ecce ego vobiscum sum omnibus diebus usque ad consummationem saeculi ".
MARK|1|1|Initium evangelii Iesu Christi Filii Dei.
MARK|1|2|Sicut scriptum est in Isaia propheta: Ecce mitto angelum meum ante faciem tuam,qui praeparabit viam tuam;
MARK|1|3|vox clamantis in deserto:Parate viam Domini, rectas facite semitas eius" ",
MARK|1|4|fuit Ioannes Baptista in deserto praedicans baptismum paenitentiae in remissionem peccatorum.
MARK|1|5|Et egrediebatur ad illum omnis Iudaeae regio et Hierosolymitae universi et baptizabantur ab illo in Iordane flumine confitentes peccata sua.
MARK|1|6|Et erat Ioannes vestitus pilis cameli, et zona pellicea circa lumbos eius, et locustas et mel silvestre edebat.
MARK|1|7|Et praedicabat dicens: " Venit fortior me post me, cuius non sum dignus procumbens solvere corrigiam calceamentorum eius.
MARK|1|8|Ego baptizavi vos aqua; ille vero baptizabit vos in Spiritu Sancto ".
MARK|1|9|Et factum est in diebus illis, venit Iesus a Nazareth Galilaeae et baptizatus est in Iordane ab Ioanne.
MARK|1|10|Et statim ascendens de aqua vidit apertos caelos et Spiritum tamquam columbam descendentem in ipsum;
MARK|1|11|et vox facta est de caelis: " Tu es Filius meus dilectus; in te complacui ".
MARK|1|12|Et statim Spiritus expellit eum in desertum.
MARK|1|13|Et erat in deserto quadraginta diebus et tentabatur a Satana; eratque cum bestiis, et angeli ministrabant illi.
MARK|1|14|Postquam autem traditus est Ioannes, venit Iesus in Galilaeam praedicans evangelium Dei
MARK|1|15|et dicens: " Impletum est tempus, et appropinquavit regnum Dei; paenitemini et credite evangelio ".
MARK|1|16|Et praeteriens secus mare Galilaeae vidit Simonem et Andream fratrem Simonis mittentes in mare; erant enim piscatores.
MARK|1|17|Et dixit eis Iesus: " Venite post me, et faciam vos fieri piscatores hominum ".
MARK|1|18|Et protinus, relictis retibus, secuti sunt eum.
MARK|1|19|Et progressus pusillum vidit Iacobum Zebedaei et Ioannem fratrem eius, et ipsos in navi componentes retia,
MARK|1|20|et statim vocavit illos. Et, relicto patre suo Zebedaeo in navi cum mercennariis, abierunt post eum.
MARK|1|21|Et ingrediuntur Capharnaum. Et statim sabbatis ingressus synagogam docebat.
MARK|1|22|Et stupebant super doctrina eius: erat enim docens eos quasi potestatem habens et non sicut scribae.
MARK|1|23|Et statim erat in synagoga eorum homo in spiritu immundo; et exclamavit
MARK|1|24|dicens: " Quid nobis et tibi, Iesu Nazarene? Venisti perdere nos? Scio qui sis: Sanctus Dei ".
MARK|1|25|Et comminatus est ei Iesus dicens: " Obmutesce et exi de homine! ".
MARK|1|26|Et discerpens eum spiritus immundus et exclamans voce magna exivit ab eo.
MARK|1|27|Et mirati sunt omnes, ita ut conquirerent inter se dicentes: " Quidnam est hoc? Doctrina nova cum potestate; et spiritibus immundis imperat, et oboediunt ei ".
MARK|1|28|Et processit rumor eius statim ubique in omnem regionem Galilaeae.
MARK|1|29|Et protinus egredientes de synagoga venerunt in domum Simonis et Andreae cum Iacobo et Ioanne.
MARK|1|30|Socrus autem Simonis decumbebat febricitans; et statim dicunt ei de illa.
MARK|1|31|Et accedens elevavit eam apprehensa manu; et dimisit eam febris, et ministrabat eis.
MARK|1|32|Vespere autem facto, cum occidisset sol, afferebant ad eum omnes male habentes et daemonia habentes;
MARK|1|33|et erat omnis civitas congregata ad ianuam.
MARK|1|34|Et curavit multos, qui vexabantur variis languoribus, et daemonia multa eiecit et non sinebat loqui daemonia, quoniam sciebant eum.
MARK|1|35|Et diluculo valde mane surgens egressus est et abiit in desertum locum ibique orabat.
MARK|1|36|Et persecutus est eum Simon et qui cum illo erant;
MARK|1|37|et cum invenissent eum, dixerunt ei: " Omnes quaerunt te! ".
MARK|1|38|Et ait illis: " Eamus alibi in proximos vicos, ut et ibi praedicem: ad hoc enim veni ".
MARK|1|39|Et venit praedicans in synagogis eorum per omnem Galilaeam et daemonia eiciens.
MARK|1|40|Et venit ad eum leprosus deprecans eum et genu flectens et dicens ei: " Si vis, potes me mundare ".
MARK|1|41|Et misertus extendens manum suam tetigit eum et ait illi: " Volo, mundare! ";
MARK|1|42|et statim discessit ab eo lepra, et mundatus est.
MARK|1|43|Et infremuit in eum statimque eiecit illum
MARK|1|44|et dicit ei: "Vide, nemini quidquam dixeris; sed vade, ostende te sacerdoti et offer pro emundatione tua, quae praecepit Moyses, in testimonium illis ".
MARK|1|45|At ille egressus coepit praedicare multum et diffamare sermonem, ita ut iam non posset manifesto in civitatem introire, sed foris in desertis locis erat; et conveniebant ad eum undique.
MARK|2|1|Et iterum intravit Capharnaum post dies, et auditum est quod in domo esset.
MARK|2|2|Et convenerunt multi, ita ut non amplius caperentur neque ad ianuam, et loquebatur eis verbum.
MARK|2|3|Et veniunt ferentes ad eum paralyticum, qui a quattuor portabatur.
MARK|2|4|Et cum non possent offerre eum illi prae turba, nudaverunt tectum, ubi erat, et perfodientes summittunt grabatum, in quo paralyticus iacebat.
MARK|2|5|Cum vidisset autem Iesus fidem illorum, ait paralytico: " Fili, dimittuntur peccata tua ".
MARK|2|6|Erant autem illic quidam de scribis sedentes et cogitantes in cordibus suis:
MARK|2|7|" Quid hic sic loquitur? Blasphemat! Quis potest dimittere peccata nisi solus Deus? ".
MARK|2|8|Quo statim cognito Iesus spiritu suo quia sic cogitarent intra se, dicit illis: " Quid ista cogitatis in cordibus vestris?
MARK|2|9|Quid est facilius, dicere paralytico: "Dimittuntur peccata tua", an dicere: "Surge et tolle grabatum tuum et ambula"?
MARK|2|10|Ut autem sciatis quia potestatem habet Filius hominis interra dimittendi peccata - ait paralytico -:
MARK|2|11|Tibi dico: Surge, tolle grabatum tuum et vade in domum tuam ".
MARK|2|12|Et surrexit et protinus sublato grabato abiit coram omnibus, ita ut admirarentur omnes et glorificarent Deum dicentes: " Numquam sic vidimus!.
MARK|2|13|Et egressus est rursus ad mare; omnisque turba veniebat ad eum, et docebat eos.
MARK|2|14|Et cum praeteriret, vidit Levin Alphaei sedentem ad teloneum et ait illi: " Sequere me ". Et surgens secutus est eum.
MARK|2|15|Et factum est, cum accumberet in domo illius, et multi publicani et peccatores simul discumbebant cum Iesu et discipulis eius; erant enim multi et sequebantur eum.
MARK|2|16|Et scribae pharisaeorum, videntes quia manducaret cum peccatoribus et publicanis, dicebant discipulis eius: " Quare cum publicanis et peccatoribus manducat? ".
MARK|2|17|Et Iesus hoc audito ait illis: " Non necesse habent sani medicum, sed qui male habent; non veni vocare iustos sed peccatores ".
MARK|2|18|Et erant discipuli Ioannis et pharisaei ieiunantes. Et veniunt et dicunt illi: " Cur discipuli Ioannis et discipuli pharisaeorum ieiunant, tui autem discipuli non ieiunant? ".
MARK|2|19|Et ait illis Iesus: " Numquid possunt convivae nuptiarum, quamdiu sponsus cum illis est, ieiunare? Quanto tempore habent secum sponsum, non possunt ieiunare;
MARK|2|20|venient autem dies, cum auferetur ab eis sponsus, et tunc ieiunabunt in illa die.
MARK|2|21|Nemo assumentum panni rudis assuit vestimento veteri; alioquin supplementum aufert aliquid ab eo, novum a veteri, et peior scissura fit.
MARK|2|22|Et nemo mittit vinum novellum in utres veteres, alioquin dirumpet vinum utres et vinum perit et utres; sed vinum novum in utres novos ".
MARK|2|23|Et factum est, cum ipse sabbatis ambularet per sata, discipuli eius coeperunt praegredi vellentes spicas.
MARK|2|24|Pharisaei autem dicebant ei: " Ecce, quid faciunt sabbatis, quod non licet? ".
MARK|2|25|Et ait illis: " Numquam legistis quid fecerit David, quando necessitatem habuit et esuriit ipse et qui cum eo erant?
MARK|2|26|Quomodo introivit in domum Dei sub Abiathar principe sacerdotum et panes propositionis manducavit, quos non licet manducare nisi sacerdotibus, et dedit etiam eis, qui cum eo erant? ".
MARK|2|27|Et dicebat eis: " Sabbatum propter hominem factum est, et non homo propter sabbatum;
MARK|2|28|itaque dominus est Filius hominis etiam sabbati ".
MARK|3|1|Et introivit iterum in synago gam. Et erat ibi homo habens manum aridam;
MARK|3|2|et observabant eum, si sabbatis curaret illum, ut accusarent eum.
MARK|3|3|Et ait homini habenti manum aridam: " Surge in medium ".
MARK|3|4|Et dicit eis: " Licet sabbatis bene facere an male? Animam salvam facere an perdere? ". At illi tacebant.
MARK|3|5|Et circumspiciens eos cum ira, contristatus super caecitate cordis eorum, dicit homini: " Extende manum ". Et extendit, et restituta est manus eius.
MARK|3|6|Et exeuntes pharisaei statim cum herodianis consilium faciebant adversus eum quomodo eum perderent.
MARK|3|7|Et Iesus cum discipulis suis secessit ad mare. Et multa turba a Galilaea secuta est et a Iudaea
MARK|3|8|et ab Hierosolymis et ab Idumaea; et, qui trans Iordanem et circa Tyrum et Sidonem, multitudo magna, audientes, quae faciebat, venerunt ad eum.
MARK|3|9|Et dixit discipulis suis, ut navicula sibi praesto esset propter turbam, ne comprimerent eum.
MARK|3|10|Multos enim sanavit, ita ut irruerent in eum, ut illum tangerent, quotquot habebant plagas.
MARK|3|11|Et spiritus immundi, cum illum videbant, procidebant ei et clamabant dicentes: " Tu es Filius Dei! ".
MARK|3|12|Et vehementer comminabatur eis, ne manifestarent illum.
MARK|3|13|Et ascendit in montem et vocat ad se, quos voluit ipse, et venerunt ad eum.
MARK|3|14|Et fecit Duodecim, ut essent cum illo, et ut mitteret eos praedicare
MARK|3|15|habentes potestatem eiciendi daemonia:
MARK|3|16|et imposuit Simoni nomen Petrum;
MARK|3|17|et Iacobum Zebedaei et Ioannem fratrem Iacobi, et imposuit eis nomina Boanerges, quod est Filii tonitrui;
MARK|3|18|et Andream et Philippum et Bartholomaeum et Matthaeum et Thomam et Iacobum Alphaei et Thaddaeum et Simonem Chananaeum
MARK|3|19|et Iudam Iscarioth, qui et tradidit illum.
MARK|3|20|Et venit ad domum; et convenit iterum turba, ita ut non possent neque panem manducare.
MARK|3|21|Et cum audissent sui, exierunt tenere eum; dicebant enim: " In furorem versus est ".
MARK|3|22|Et scribae, qui ab Hierosolymis descenderant, dicebant: " Beelzebul habet " et: " In principe daemonum eicit daemonia ".
MARK|3|23|Et convocatis eis, in parabolis dicebat illis: " Quomodo potest Satanas Satanam eicere?
MARK|3|24|Et si regnum in se dividatur, non potest stare regnum illud;
MARK|3|25|et si domus in semetipsam dispertiatur, non poterit domus illa stare.
MARK|3|26|Et si Satanas consurrexit in semetipsum et dispertitus est, non potest stare, sed finem habet.
MARK|3|27|Nemo autem potest in domum fortis ingressus vasa eius diripere, nisi prius fortem alliget; et tunc domum eius diripiet.
MARK|3|28|Amen dico vobis: Omnia dimittentur filiis hominum peccata et blasphemiae, quibus blasphemaverint;
MARK|3|29|qui autem blasphemaverit in Spiritum Sanctum, non habet remissionem in aeternum, sed reus est aeterni delicti ".
MARK|3|30|Quoniam dicebant: " Spiritum immundum habet ".
MARK|3|31|Et venit mater eius et fratres eius, et foris stantes miserunt ad eum vocantes eum.
MARK|3|32|Et sedebat circa eum turba, et dicunt ei: " Ecce mater tua et fratres tui et sorores tuae foris quaerunt te ".
MARK|3|33|Et respondens eis ait: " Quae est mater mea et fratres mei? ".
MARK|3|34|Et circumspiciens eos, qui in circuitu eius sedebant, ait: " Ecce mater mea et fratres mei.
MARK|3|35|Qui enim fecerit voluntatem Dei, hic frater meus et soror mea et mater est ".
MARK|4|1|Et iterum coepit docere ad ma re. Et congregatur ad eum tur ba plurima, ita ut in navem ascendens sederet in mari, et omnis turba circa mare super terram erant.
MARK|4|2|Et docebat eos in parabolis multa et dicebat illis in doctrina sua:
MARK|4|3|" Audite. Ecce exiit seminans ad seminandum.
MARK|4|4|Et factum est, dum seminat, aliud cecidit circa viam, et venerunt volucres et comederunt illud.
MARK|4|5|Aliud cecidit super petrosa, ubi non habebat terram multam, et statim exortum est, quoniam non habebat altitudinem terrae;
MARK|4|6|et quando exortus est sol, exaestuavit et, eo quod non haberet radicem, exaruit.
MARK|4|7|Et aliud cecidit in spinas, et ascenderunt spinae et suffocaverunt illud, et fructum non dedit.
MARK|4|8|Et alia ceciderunt in terram bonam et dabant fructum: ascendebant et crescebant et afferebant unum triginta et unum sexaginta et unum centum ".
MARK|4|9|Et dicebat: " Qui habet aures audiendi, audiat ".
MARK|4|10|Et cum esset singularis, interrogaverunt eum hi, qui circa eum erant cum Duodecim, parabolas.
MARK|4|11|Et dicebat eis: " Vobis datum est mysterium regni Dei; illis autem, qui foris sunt, in parabolis omnia fiunt,
MARK|4|12|ut videntes videant et non videant,et audientes audiant et non intellegant,ne quando convertantur,et dimittatur eis ".
MARK|4|13|Et ait illis: " Nescitis parabolam hanc, et quomodo omnes parabolas cognoscetis?
MARK|4|14|Qui seminat, verbum seminat.
MARK|4|15|Hi autem sunt, qui circa viam, ubi seminatur verbum: et cum audierint, confestim venit Satanas et aufert verbum, quod seminatum est in eos.
MARK|4|16|Et hi sunt, qui super petrosa seminantur: qui cum audierint verbum, statim cum gaudio accipiunt illud
MARK|4|17|et non habent radicem in se, sed temporales sunt; deinde orta tribulatione vel persecutione propter verbum, confestim scandalizantur.
MARK|4|18|Et alii sunt, qui in spinis seminantur: hi sunt, qui verbum audierunt,
MARK|4|19|et aerumnae saeculi et deceptio divitiarum et circa reliqua concupiscentiae introeuntes suffocant verbum, et sine fructu efficitur.
MARK|4|20|Et hi sunt, qui super terram bonam seminati sunt: qui audiunt verbum et suscipiunt et fructificant unum triginta et unum sexaginta et unum centum.
MARK|4|21|Et dicebat illis: " Numquid venit lucerna, ut sub modio ponatur aut sub lecto? Nonne ut super candelabrum ponatur?
MARK|4|22|Non enim est aliquid absconditum, nisi ut manifestetur, nec factum est occultum, nisi ut in palam veniat.
MARK|4|23|Si quis habet aures audiendi, audiat ".
MARK|4|24|Et dicebat illis: " Videte quid audiatis. In qua mensura mensi fueritis, remetietur vobis et adicietur vobis.
MARK|4|25|Qui enim habet, dabitur illi; et, qui non habet, etiam quod habet, auferetur ab illo ".
MARK|4|26|Et dicebat: " Sic est regnum Dei, quemadmodum si homo iaciat sementem in terram
MARK|4|27|et dormiat et exsurgat nocte ac die, et semen germinet et increscat, dum nescit ille.
MARK|4|28|Ultro terra fructificat primum herbam, deinde spicam, deinde plenum frumentum in spica.
MARK|4|29|Et cum se produxerit fructus, statim mittit falcem, quoniam adest messis ".
MARK|4|30|Et dicebat: " Quomodo assimilabimus regnum Dei aut in qua parabola ponemus illud?
MARK|4|31|Sicut granum sinapis, quod cum seminatum fuerit in terra, minus est omnibus seminibus, quae sunt in terra;
MARK|4|32|et cum seminatum fuerit, ascendit et fit maius omnibus holeribus et facit ramos magnos, ita ut possint sub umbra eius aves caeli habitare ".
MARK|4|33|Et talibus multis parabolis loquebatur eis verbum, prout poterant audire;
MARK|4|34|sine parabola autem non loquebatur eis. Seorsum autem discipulis suis disserebat omnia.
MARK|4|35|Et ait illis illa die, cum sero esset factum: " Transeamus contra ".
MARK|4|36|Et dimittentes turbam, assumunt eum, ut erat in navi; et aliae naves erant cum illo.
MARK|4|37|Et exoritur procella magna venti, et fluctus se mittebant in navem, ita ut iam impleretur navis.
MARK|4|38|Et erat ipse in puppi supra cervical dormiens; et excitant eum et dicunt ei: " Magister, non ad te pertinet quia perimus? ".
MARK|4|39|Et exsurgens comminatus est vento et dixit mari: " Tace, obmutesce! ". Et cessavit ventus, et facta est tranquillitas magna.
MARK|4|40|Et ait illis: " Quid timidi estis? Necdum habetis fidem? ".
MARK|4|41|Et timuerunt magno timore et dicebant ad alterutrum: " Quis putas est iste, quia et ventus et mare oboediunt ei? ".
MARK|5|1|Et venerunt trans fretum maris in regionem Gerasenorum.
MARK|5|2|Et exeunte eo de navi, statim occurrit ei de monumentis homo in spiritu immundo,
MARK|5|3|qui domicilium habebat in monumentis; et neque catenis iam quisquam eum poterat ligare,
MARK|5|4|quoniam saepe compedibus et catenis vinctus dirupisset catenas et compedes comminuisset, et nemo poterat eum domare;
MARK|5|5|et semper nocte ac die in monumentis et in montibus erat clamans et concidens se lapidibus.
MARK|5|6|Et videns Iesum a longe cucurrit et adoravit eum
MARK|5|7|et clamans voce magna dicit: " Quid mihi et tibi, Iesu, fili Dei Altissimi? Adiuro te per Deum, ne me torqueas ".
MARK|5|8|Dicebat enim illi: " Exi, spiritus immunde, ab homine ".
MARK|5|9|Et interrogabat eum: " Quod tibi nomen est? ". Et dicit ei: " Legio nomen mihi est, quia multi sumus ".
MARK|5|10|Et deprecabatur eum multum, ne se expelleret extra regionem.
MARK|5|11|Erat autem ibi circa montem grex porcorum magnus pascens;
MARK|5|12|et deprecati sunt eum dicentes: " Mitte nos in porcos, ut in eos introeamus ".
MARK|5|13|Et concessit eis. Et exeuntes spiritus immundi introierunt in porcos. Et magno impetu grex ruit per praecipitium in mare, ad duo milia, et suffocabantur in mari.
MARK|5|14|Qui autem pascebant eos, fugerunt et nuntiaverunt in civitatem et in agros; et egressi sunt videre quid esset facti.
MARK|5|15|Et veniunt ad Iesum; et vident illum, qui a daemonio vexabatur, sedentem, vestitum et sanae mentis, eum qui legionem habuerat, et timuerunt.
MARK|5|16|Et qui viderant, narraverunt illis qualiter factum esset ei, qui daemonium habuerat, et de porcis.
MARK|5|17|Et rogare eum coeperunt, ut discederet a finibus eorum.
MARK|5|18|Cumque ascenderet navem, qui daemonio vexatus fuerat, deprecabatur eum, ut esset cum illo.
MARK|5|19|Et non admisit eum, sed ait illi: " Vade in domum tuam ad tuos et annuntia illis quanta tibi Dominus fecerit et misertus sit tui ".
MARK|5|20|Et abiit et coepit praedicare in Decapoli quanta sibi fecisset Iesus, et omnes mirabantur.
MARK|5|21|Et cum transcendisset Iesus in navi rursus trans fretum, convenit turba multa ad illum, et erat circa mare.
MARK|5|22|Et venit quidam de archisynagogis nomine Iairus et videns eum procidit ad pedes eius
MARK|5|23|et deprecatur eum multum dicens: " Filiola mea in extremis est; veni, impone manus super eam, ut salva sit et vivat ".
MARK|5|24|Et abiit cum illo. Et sequebatur eum turba multa et comprimebant illum.
MARK|5|25|Et mulier, quae erat in profluvio sanguinis annis duodecim
MARK|5|26|et fuerat multa perpessa a compluribus medicis et erogaverat omnia sua nec quidquam profecerat, sed magis deterius habebat,
MARK|5|27|cum audisset de Iesu, venit in turba retro et tetigit vestimentum eius;
MARK|5|28|dicebat enim: " Si vel vestimenta eius tetigero, salva ero ".
MARK|5|29|Et confestim siccatus est fons sanguinis eius, et sensit corpore quod sanata esset a plaga.
MARK|5|30|Et statim Iesus cognoscens in semetipso virtutem, quae exierat de eo, conversus ad turbam aiebat: " Quis tetigit vestimenta mea? ".
MARK|5|31|Et dicebant ei discipuli sui: " Vides turbam comprimentem te et dicis: Quis me tetigit?" ".
MARK|5|32|Et circumspiciebat videre eam, quae hoc fecerat.
MARK|5|33|Mulier autem timens et tremens, sciens quod factum esset in se, venit et procidit ante eum et dixit ei omnem veritatem.
MARK|5|34|Ille autem dixit ei: " Filia, fides tua te salvam fecit. Vade in pace et esto sana a plaga tua ".
MARK|5|35|Adhuc eo loquente, veniunt ab archisynagogo dicentes: " Filia tua mortua est; quid ultra vexas magistrum? ".
MARK|5|36|Iesus autem, verbo, quod dicebatur, audito, ait archisynagogo: " Noli timere; tantummodo crede! ".
MARK|5|37|Et non admisit quemquam sequi se nisi Petrum et Iacobum et Ioannem fratrem Iacobi.
MARK|5|38|Et veniunt ad domum archisynagogi; et videt tumultum et flentes et eiulantes multum,
MARK|5|39|et ingressus ait eis: " Quid turbamini et ploratis? Puella non est mortua, sed dormit ".
MARK|5|40|Et irridebant eum. Ipse vero, eiectis omnibus, assumit patrem puellae et matrem et, qui secum erant, et ingreditur, ubi erat puella;
MARK|5|41|et tenens manum puellae ait illi: " Talitha, qum! " - quod est interpretatum: " Puella, tibi dico: Surge! " -.
MARK|5|42|Et confestim surrexit puella et ambulabat; erat enim annorum duodecim. Et obstupuerunt continuo stupore magno.
MARK|5|43|Et praecepit illis vehementer, ut nemo id sciret, et dixit dari illi manducare.
MARK|6|1|Et egressus est inde et venit in patriam suam, et sequuntur il lum discipuli sui.
MARK|6|2|Et facto sabbato, coepit in synagoga docere; et multi audientes admirabantur dicentes: " Unde huic haec, et quae est sapientia, quae data est illi, et virtutes tales, quae per manus eius efficiuntur?
MARK|6|3|Nonne iste est faber, filius Mariae et frater Iacobi et Iosetis et Iudae et Simonis? Et nonne sorores eius hic nobiscum sunt? ". Et scandalizabantur in illo.
MARK|6|4|Et dicebat eis Iesus: " Non est propheta sine honore nisi in patria sua et in cognatione sua et in domo sua ".
MARK|6|5|Et non poterat ibi virtutem ullam facere, nisi paucos infirmos impositis manibus curavit;
MARK|6|6|et mirabatur propter incredulitatem eorum.Et circumibat castella in circuitu docens.
MARK|6|7|Et convocat Duodecim et coepit eos mittere binos et dabat illis potestatem in spiritus immundos;
MARK|6|8|et praecepit eis, ne quid tollerent in via nisi virgam tantum: non panem, non peram neque in zona aes,
MARK|6|9|sed ut calcearentur sandaliis et ne induerentur duabus tunicis.
MARK|6|10|Et dicebat eis: " Quocumque introieritis in domum, illic manete, donec exeatis inde.
MARK|6|11|Et quicumque locus non receperit vos nec audierint vos, exeuntes inde excutite pulverem de pedibus vestris in testimonium illis ".
MARK|6|12|Et exeuntes praedicaverunt, ut paenitentiam agerent;
MARK|6|13|et daemonia multa eiciebant et ungebant oleo multos aegrotos et sanabant.
MARK|6|14|Et audivit Herodes rex; manifestum enim factum est nomen eius. Et dicebant: " Ioannes Baptista resurrexit a mortuis, et propterea inoperantur virtutes in illo ".
MARK|6|15|Alii autem dicebant: " Elias est ". Alii vero dicebant: " Propheta est, quasi unus ex prophetis ".
MARK|6|16|Quo audito, Herodes aiebat: " Quem ego decollavi Ioannem, hic resurrexit! ".
MARK|6|17|Ipse enim Herodes misit ac tenuit Ioannem et vinxit eum in carcere propter Herodiadem uxorem Philippi fratris sui, quia duxerat eam.
MARK|6|18|Dicebat enim Ioannes Herodi: " Non licet tibi habere uxorem fratris tui.
MARK|6|19|Herodias autem insidiabatur illi et volebat occidere eum nec poterat:
MARK|6|20|Herodes enim metuebat Ioannem, sciens eum virum iustum et sanctum, et custodiebat eum, et, audito eo, multum haesitabat et libenter eum audiebat.
MARK|6|21|Et cum dies opportunus accidisset, quo Herodes natali suo cenam fecit principibus suis et tribunis et primis Galilaeae,
MARK|6|22|cumque introisset filia ipsius Herodiadis et saltasset, placuit Herodi simulque recumbentibus. Rex ait puellae: " Pete a me, quod vis, et dabo tibi ".
MARK|6|23|Et iuravit illi multum: " Quidquid petieris a me, dabo tibi, usque ad dimidium regni mei ".
MARK|6|24|Quae cum exisset, dixit matri suae: " Quid petam? ". At illa dixit: " Caput Ioannis Baptistae ".
MARK|6|25|Cumque introisset statim cum festinatione ad regem, petivit dicens: " Volo ut protinus des mihi in disco caput Ioannis Baptistae ".
MARK|6|26|Et contristatus rex, propter iusiurandum et propter recumbentes noluit eam decipere;
MARK|6|27|et statim misso spiculatore rex praecepit afferri caput eius. Et abiens decollavit eum in carcere
MARK|6|28|et attulit caput eius in disco; et dedit illud puellae, et puella dedit illud matri suae.
MARK|6|29|Quo audito, discipuli eius venerunt et tulerunt corpus eius et posuerunt illud in monumento.
MARK|6|30|Et convenientes apostoli ad Iesum renuntiaverunt illi omnia, quae egerant et docuerant.
MARK|6|31|Et ait illis: " Venite vos ipsi seorsum in desertum locum et requiescite pusillum ". Erant enim, qui veniebant et redibant, multi, et nec manducandi spatium habebant.
MARK|6|32|Et abierunt in navi in desertum locum seorsum.
MARK|6|33|Et viderunt eos abeuntes et cognoverunt multi; et pedestre de omnibus civitatibus concurrerunt illuc et praevenerunt eos.
MARK|6|34|Et exiens vidit multam turbam et misertus est super eos, quia erant sicut oves non habentes pastorem, et coepit docere illos multa.
MARK|6|35|Et cum iam hora multa facta esset, accesserunt discipuli eius dicentes: Desertus est locus hic, et hora iam est multa;
MARK|6|36|dimitte illos, ut euntes in villas et vicos in circuitu emant sibi, quod manducent ".
MARK|6|37|Respondens autem ait illis: " Date illis vos manducare ". Et dicunt ei: Euntes emamus denariis ducentis panes et dabimus eis manducare? ".
MARK|6|38|Et dicit eis: " Quot panes habetis? Ite, videte ". Et cum cognovissent, dicunt: " Quinque et duos pisces ".
MARK|6|39|Et praecepit illis, ut accumbere facerent omnes secundum contubernia super viride fenum.
MARK|6|40|Et discubuerunt secundum areas per centenos et per quinquagenos.
MARK|6|41|Et acceptis quinque panibus et duobus piscibus, intuens in caelum benedixit et fregit panes et dabat discipulis suis, ut ponerent ante eos; et duos pisces divisit omnibus.
MARK|6|42|Et manducaverunt omnes et saturati sunt;
MARK|6|43|et sustulerunt fragmenta duodecim cophinos plenos, et de piscibus.
MARK|6|44|Et erant, qui manducaverunt panes, quinque milia virorum.
MARK|6|45|Et statim coegit discipulos suos ascendere navem, ut praecederent trans fretum ad Bethsaidam, dum ipse dimitteret populum.
MARK|6|46|Et cum dimisisset eos, abiit in montem orare.
MARK|6|47|Et cum sero factum esset, erat navis in medio mari, et ipse solus in terra.
MARK|6|48|Et videns eos laborantes in remigando, erat enim ventus contrarius eis, circa quartam vigiliam noctis venit ad eos ambulans super mare et volebat praeterire eos.
MARK|6|49|At illi, ut viderunt eum ambulantem super mare, putaverunt phantasma esse et exclamaverunt;
MARK|6|50|omnes enim eum viderunt et conturbati sunt. Statim autem locutus est cum eis et dicit illis: " Confidite, ego sum; nolite timere! ".
MARK|6|51|Et ascendit ad illos in navem, et cessavit ventus. Et valde nimis intra se stupebant;
MARK|6|52|non enim intellexerant de panibus, sed erat cor illorum obcaecatum.
MARK|6|53|Et cum transfretassent in terram, pervenerunt Gennesaret et applicuerunt.
MARK|6|54|Cumque egressi essent de navi, continuo cognoverunt eum
MARK|6|55|et percurrentes universam regionem illam coeperunt in grabatis eos, qui se male habebant, circumferre, ubi audiebant eum esse.
MARK|6|56|Et quocumque introibat in vicos aut in civitates vel in villas, in plateis ponebant infirmos; et deprecabantur eum, ut vel fimbriam vestimenti eius tangerent; et, quotquot tangebant eum, salvi fiebant.
MARK|7|1|Et conveniunt ad eum pharisaei et quidam de scribis venientes ab Hierosolymis;
MARK|7|2|et cum vidissent quosdam ex discipulis eius communibus manibus, id est non lotis, manducare panes
MARK|7|3|- pharisaei enim et omnes Iudaei, nisi pugillo lavent manus, non manducant, tenentes traditionem seniorum;
MARK|7|4|et a foro nisi baptizentur, non comedunt; et alia multa sunt, quae acceperunt servanda: baptismata calicum et urceorum et aeramentorum et lectorum -
MARK|7|5|et interrogant eum pharisaei et scribae: " Quare discipuli tui non ambulant iuxta traditionem seniorum, sed communibus manibus manducant panem? ".
MARK|7|6|At ille dixit eis: " Bene prophetavit Isaias de vobis hypocritis, sicut scriptum est:Populus hic labiis me honorat,cor autem eorum longe est a me;
MARK|7|7|in vanum autem me coluntdocentes doctrinas praecepta hominum".
MARK|7|8|Relinquentes mandatum Dei tenetis traditionem hominum ".
MARK|7|9|Et dicebat illis: " Bene irritum facitis praeceptum Dei, ut traditionem vestram servetis.
MARK|7|10|Moyses enim dixit: "Honora patrem tuum et matrem tuam" et: "Qui maledixerit patri aut matri, morte moriatur";
MARK|7|11|vos autem dicitis: "Si dixerit homo patri aut matri: Corban, quod est donum, quodcumque ex me tibi profuerit",
MARK|7|12|ultra non permittitis ei facere quidquam patri aut matri
MARK|7|13|rescindentes verbum Dei per traditionem vestram, quam tradidistis; et similia huiusmodi multa facitis ".
MARK|7|14|Et advocata iterum turba, dicebat illis: " Audite me, omnes, et intellegite:
MARK|7|15|Nihil est extra hominem introiens in eum, quod possiteum coinquinare; sed quae de homine procedunt, illa sunt, quae coinquinant hominem! ".
MARK|7|16|()
MARK|7|17|Et cum introisset in domum a turba, interrogabant eum discipuli eius parabolam.
MARK|7|18|Et ait illis: " Sic et vos imprudentes estis? Non intellegitis quia omne extrinsecus introiens in hominem non potest eum coinquinare,
MARK|7|19|quia non introit in cor eius sed in ventrem et in secessum exit? ", purgans omnes escas.
MARK|7|20|Dicebat autem: " Quod de homine exit, illud coinquinat hominem;
MARK|7|21|ab intus enim de corde hominum cogitationes malae procedunt, fornicationes, furta, homicidia,
MARK|7|22|adulteria, avaritiae, nequitiae, dolus, impudicitia, oculus malus, blasphemia, superbia, stultitia:
MARK|7|23|omnia haec mala ab intus procedunt et coinquinant hominem ".
MARK|7|24|Inde autem surgens abiit in fines Tyri et Sidonis. Et ingressus domum neminem voluit scire et non potuit latere.
MARK|7|25|Sed statim ut audivit de eo mulier, cuius habebat filia spiritum immundum, veniens procidit ad pedes eius.
MARK|7|26|Erat autem mulier Graeca, Syrophoenissa genere. Et rogabat eum, ut daemonium eiceret de filia eius.
MARK|7|27|Et dicebat illi: " Sine prius saturari filios; non est enim bonum sumere panem filiorum et mittere catellis ".
MARK|7|28|At illa respondit et dicit ei: " Domine, etiam catelli sub mensa comedunt de micis puerorum ".
MARK|7|29|Et ait illi: " Propter hunc sermonem vade; exiit daemonium de filia tua.
MARK|7|30|Et cum abisset domum suam, invenit puellam iacentem supra lectum et daemonium exisse.
MARK|7|31|Et iterum exiens de finibus Tyri venit per Sidonem ad mare Galilaeae inter medios fines Decapoleos.
MARK|7|32|Et adducunt ei surdum et mutum et deprecantur eum, ut imponat illi manum.
MARK|7|33|Et apprehendens eum de turba seorsum misit digitos suos in auriculas eius et exspuens tetigit linguam eius
MARK|7|34|et suspiciens in caelum ingemuit et ait illi: " Effetha ", quod est: " Adaperire ".
MARK|7|35|Et statim apertae sunt aures eius, et solutum est vinculum linguae eius, et loquebatur recte.
MARK|7|36|Et praecepit illis, ne cui dicerent; quanto autem eis praecipiebat, tanto magis plus praedicabant.
MARK|7|37|Et eo amplius admirabantur dicentes: " Bene omnia fecit, et surdos facit audire et mutos loqui! ".
MARK|8|1|In illis diebus iterum cum turba multa esset nec haberent, quod manducarent, convocatis discipulis, ait illis:
MARK|8|2|" Misereor super turbam, quia iam triduo sustinent me nec habent, quod manducent;
MARK|8|3|et si dimisero eos ieiunos in domum suam, deficient in via; et quidam ex eis de longe venerunt ".
MARK|8|4|Et responderunt ei discipuli sui: " Unde istos poterit quis hic saturare panibus in solitudine? ".
MARK|8|5|Et interrogabat eos: " Quot panes habetis? ". Qui dixerunt: " Septem ".
MARK|8|6|Et praecipit turbae discumbere supra terram; et accipiens septem panes, gratias agens fregit et dabat discipulis suis, ut apponerent; et apposuerunt turbae.
MARK|8|7|Et habebant pisciculos paucos; et benedicens eos, iussit hos quoque apponi.
MARK|8|8|Et manducaverunt et saturati sunt; et sustulerunt, quod superaverat de fragmentis, septem sportas.
MARK|8|9|Erant autem quasi quattuor milia. Et dimisit eos.
MARK|8|10|Et statim ascendens navem cum discipulis suis venit in partes Dalmanutha.
MARK|8|11|Et exierunt pharisaei et coeperunt conquirere cum eo quaerentes ab illo signum de caelo, tentantes eum.
MARK|8|12|Et ingemiscens spiritu suo ait: " Quid generatio ista quaerit signum? Amen dico vobis: Non dabitur generationi isti signum ".
MARK|8|13|Et dimittens eos, iterum ascendens abiit trans fretum.
MARK|8|14|Et obliti sunt sumere panes et nisi unum panem non habebant secum in navi.
MARK|8|15|Et praecipiebat eis dicens: " Videte, cavete a fermento pharisaeorum et fermento Herodis! ".
MARK|8|16|Et disputabant ad invicem, quia panes non haberent.
MARK|8|17|Quo cognito, ait illis: " Quid disputatis, quia panes non habetis? Nondum cognoscitis nec intellegitis? Caecatum habetis cor vestrum?
MARK|8|18|Oculos habentes non videtis, et aures habentes non auditis? Nec recordamini,
MARK|8|19|quando quinque panes fregi in quinque milia, quot cophinos fragmentorum plenos sustulistis? ". Dicunt ei: " Duodecim ".
MARK|8|20|" Quando illos septem in quattuor milia, quot sportas plenas fragmentorum tulistis? ". Et dicunt ei: " Septem ".
MARK|8|21|Et dicebat eis: " Nondum intellegitis? ".
MARK|8|22|Et veniunt Bethsaida. Et adducunt ei caecum et rogant eum, ut illum tangat.
MARK|8|23|Et apprehendens manum caeci eduxit eum extra vicum; et exspuens in oculos eius, impositis manibus ei, interrogabat eum: " Vides aliquid? ".
MARK|8|24|Et aspiciens dicebat: " Video homines, quia velut arbores video ambulantes ".
MARK|8|25|Deinde iterum imposuit manus super oculos eius; et coepit videre et restitutus est et videbat clare omnia.
MARK|8|26|Et misit illum in domum suam dicens: " Nec in vicum introieris ".
MARK|8|27|Et egressus est Iesus et discipuli eius in castella Caesareae Philippi; et in via interrogabat discipulos suos dicens eis: " Quem me dicunt esse homines? ".
MARK|8|28|Qui responderunt illi dicentcs: " Ioannem Baptistam, alii Eliam, alii vero unum de prophetis ".
MARK|8|29|Et ipse interrogabat eos: " Vos vero quem me dicitis esse? ". Respondens Petrus ait ei: " Tu es Christus ".
MARK|8|30|Et comminatus est eis, ne cui dicerent de illo.
MARK|8|31|Et coepit docere illos: " Oportet Filium hominis multa pati et reprobari a senioribus et a summis sacerdotibus et scribis et occidi et post tres dies resurgere ";
MARK|8|32|et palam verbum loquebatur. Et apprehendens eum Petrus coepit increpare eum.
MARK|8|33|Qui conversus et videns discipulos suos comminatus est Petro et dicit: Vade retro me, Satana, quoniam non sapis, quae Dei sunt, sed quae sunt hominum ".
MARK|8|34|Et convocata turba cum discipulis suis, dixit eis: " Si quis vult post me sequi, deneget semetipsum et tollat crucem suam et sequatur me.
MARK|8|35|Qui enim voluerit animam suam salvam facere, perdet eam; qui autem perdiderit animam suam propter me et evangelium, salvam eam faciet.
MARK|8|36|Quid enim prodest homini, si lucretur mundum totum et detrimentum faciat animae suae?
MARK|8|37|Quid enim dabit homo commutationem pro anima sua?
MARK|8|38|Qui enim me confusus fuerit et mea verba in generatione ista adultera et peccatrice, et Filius hominis confundetur eum, cum venerit in gloria Patris sui cum angelis sanctis ".
MARK|9|1|Et dicebat illis: " Amen dico vobis: Sunt quidam de hic stan tibus, qui non gustabunt mortem, donec videant regnum Dei venisse in virtute ".
MARK|9|2|Et post dies sex assumit Iesus Petrum et Iacobum et Ioannem, et ducit illos in montem excelsum seorsum solos. Et transfiguratus est coram ipsis;
MARK|9|3|et vestimenta eius facta sunt splendentia, candida nimis, qualia fullo super terram non potest tam candida facere.
MARK|9|4|Et apparuit illis Elias cum Moyse, et erant loquentes cum Iesu.
MARK|9|5|Et respondens Petrus ait Iesu: " Rabbi, bonum est nos hic esse; et faciamus tria tabernacula: tibi unum et Moysi unum et Eliae unum ".
MARK|9|6|Non enim sciebat quid responderet; erant enim exterriti.
MARK|9|7|Et facta est nubes obumbrans eos, et venit vox de nube: " Hic est Filius meus dilectus; audite illum ".
MARK|9|8|Et statim circumspicientes neminem amplius viderunt nisi Iesum tantum secum.
MARK|9|9|Et descendentibus illis de monte, praecepit illis, ne cui, quae vidissent, narrarent, nisi cum Filius hominis a mortuis resurrexerit.
MARK|9|10|Et verbum continuerunt apud se, conquirentes quid esset illud: " a mortuis resurgere ".
MARK|9|11|Et interrogabant eum dicentes: " Quid ergo dicunt scribae quia Eliam oporteat venire primum? ".
MARK|9|12|Qui ait illis: " Elias veniens primo, restituit omnia; et quomodo scriptum est super Filio hominis, ut multa patiatur et contemnatur?
MARK|9|13|Sed dico vobis: Et Elias venit; et fecerunt illi, quaecumque volebant, sicut scriptum est de eo ".
MARK|9|14|Et venientes ad discipulos viderunt turbam magnam circa eos et scribas conquirentes cum illis.
MARK|9|15|Et confestim omnis populus videns eum stupefactus est, et accurrentes salutabant eum.
MARK|9|16|Et interrogavit eos: " Quid inter vos conquiritis? ".
MARK|9|17|Et respondit ei unus de turba: " Magister, attuli filium meum ad te habentem spiritum mutum;
MARK|9|18|et ubicumque eum apprehenderit, allidit eum, et spumat et stridet dentibus et arescit. Et dixi discipulis tuis, ut eicerent illum, et non potuerunt ".
MARK|9|19|Qui respondens eis dicit: " O generatio incredula, quamdiu apud vos ero? Quamdiu vos patiar? Afferte illum ad me ".
MARK|9|20|Et attulerunt illum ad eum. Et cum vidisset illum, spiritus statim conturbavit eum; et corruens in terram volutabatur spumans.
MARK|9|21|Et interrogavit patrem eius: " Quantum temporis est, ex quo hoc ei accidit? ". At ille ait: " Ab infantia;
MARK|9|22|et frequenter eum etiam in ignem et in aquas misit, ut eum perderet; sed si quid potes, adiuva nos, misertus nostri ".
MARK|9|23|Iesus autem ait illi: " "Si potes!". Omnia possibilia credenti ".
MARK|9|24|Et continuo exclamans pater pueri aiebat: " Credo; adiuva incredulitatem meam ".
MARK|9|25|Et cum videret Iesus concurrentem turbam, comminatus est spiritui immundo dicens illi: " Mute et surde spiritus, ego tibi praecipio: Exi ab eo et amplius ne introeas in eum ".
MARK|9|26|Et clamans et multum discerpens eum exiit; et factus est sicut mortuus, ita ut multi dicerent: " Mortuus est! ".
MARK|9|27|Iesus autem tenens manum eius elevavit illum, et surrexit.
MARK|9|28|Et cum introisset in domum, discipuli eius secreto interrogabant eum: " Quare nos non potuimus eicere eum? ".
MARK|9|29|Et dixit illis: " Hoc genus in nullo potest exire nisi in oratione ".
MARK|9|30|Et inde profecti peragrabant Galilaeam; nec volebat quemquam scire.
MARK|9|31|Docebat enim discipulos suos et dicebat illis: " Filius hominis traditur in manus hominum, et occident eum, et occisus post tres dies resurget ".
MARK|9|32|At illi ignorabant verbum et timebant eum interrogare.
MARK|9|33|Et venerunt Capharnaum. Qui cum domi esset, interrogabat eos: " Quid in via tractabatis? ".
MARK|9|34|At illi tacebant. Siquidem inter se in via disputaverant, quis esset maior.
MARK|9|35|Et residens vocavit Duodecim et ait illis: " Si quis vult primus esse, erit omnium novissimus et omnium minister ".
MARK|9|36|Et accipiens puerum, statuit eum in medio eorum; quem ut complexus esset, ait illis:
MARK|9|37|" Quisquis unum ex huiusmodi pueris receperit in nomine meo, me recipit; et, quicumque me susceperit, non me suscipit, sed eum qui me misit ".
MARK|9|38|Dixit illi Ioannes: " Magister, vidimus quendam in nomine tuo eicientem daemonia, et prohibebamus eum, quia non sequebatur nos ".
MARK|9|39|Iesus autem ait: " Nolite prohibere eum. Nemo est enim, qui faciat virtutem in nomine meo et possit cito male loqui de me;
MARK|9|40|qui enim non est adversum nos, pro nobis est.
MARK|9|41|Quisquis enim potum dederit vobis calicem aquae in nomine, quia Christi estis, amen dico vobis: Non perdet mercedem suam.
MARK|9|42|Et quisquis scandalizaverit unum ex his pusillis credentibus in me, bonum est ei magis, ut circumdetur mola asinaria collo eius, et in mare mittatur.
MARK|9|43|Et si scandalizaverit te manus tua, abscide illam: bonum est tibi debilem introire in vitam, quam duas manus habentem ire ingehennam, in ignem inexstinguibilem.
MARK|9|44|()
MARK|9|45|Et si pes tuus te scandalizat, amputa illum: bonum est tibi claudum introire in vitam,quam duos pedes habentem mitti in gehennam.
MARK|9|46|()
MARK|9|47|Et si oculus tuus scandalizat te, eice eum: bonum est tibi luscum introire in regnum Dei, quam duos oculos habentem mitti in gehennam,
MARK|9|48|ubi vermis eorum non moritur, et ignis non exstinguitur;
MARK|9|49|omnis enim igne salietur.
MARK|9|50|Bonum est sal; quod si sal insulsum fuerit, in quo illud condietis? Habete in vobis sal et pacem habete inter vos ".
MARK|10|1|Et inde exsurgens venit in fines Iudaeae ultra Iorda nem; et conveniunt iterum turbae ad eum, et, sicut consueverat, iterum docebat illos.
MARK|10|2|Et accedentes pharisaei interrogabant eum, si licet viro uxorem dimittere, tentantes eum.
MARK|10|3|At ille respondens dixit eis: " Quid vobis praecepit Moyses? ".
MARK|10|4|Qui dixerunt: " Moyses permisit libellum repudii scribere et dimittere.
MARK|10|5|Iesus autem ait eis: " Ad duritiam cordis vestri scripsit vobis praeceptum istud.
MARK|10|6|Ab initio autem creaturae masculum et feminam fecit eos.
MARK|10|7|Propter hoc relinquet homo patrem suum et matrem et adhaerebit ad uxorern suam,
MARK|10|8|et erunt duo in carne una; itaque iam non sunt duo sed una caro.
MARK|10|9|Quod ergo Deus coniunxit, homo non separet ".
MARK|10|10|Et domo iterum discipuli de hoc interrogabant eum.
MARK|10|11|Et dicit illis: " Quicumque dimiserit uxorem suam et aliam duxerit, adulterium committit in eam;
MARK|10|12|et si ipsa dimiserit virum suum et alii nupserit, moechatur ".
MARK|10|13|Et offerebant illi parvulos, ut tangeret illos; discipuli autem comminabantur eis.
MARK|10|14|At videns Iesus, indigne tulit et ait illis: " Sinite parvulos venire ad me. Ne prohibueritis eos; talium est enim regnum Dei.
MARK|10|15|Amen dico vobis: Quisquis non receperit regnum Dei velut parvulus, non intrabit in illud ".
MARK|10|16|Et complexans eos benedicebat imponens manus super illos.
MARK|10|17|Et cum egrederetur in viam, accurrens quidam et, genu flexo ante eum, rogabat eum: " Magister bone, quid faciam ut vitam aeternam percipiam? ".
MARK|10|18|Iesus autem dixit ei: " Quid me dicis bonum? Nemo bonus, nisi unus Deus.
MARK|10|19|Praecepta nosti: ne occidas, ne adulteres, ne fureris, ne falsum testimonium dixeris, ne fraudem feceris, honora patrem tuum et matrem ".
MARK|10|20|Ille autem dixit ei: " Magister, haec omnia conservavi a iuventute mea.
MARK|10|21|Iesus autem intuitus eum dilexit eum et dixit illi: " Unum tibi deest: vade, quaecumque habes, vende et da pauperibus et habebis thesaurum in caelo; et veni, sequere me ".
MARK|10|22|Qui contristatus in hoc verbo, abiit maerens: erat enim habens possessiones multas.
MARK|10|23|Et circumspiciens Iesus ait discipulis suis: " Quam difficile, qui pecunias habent, in regnum Dei introibunt ".
MARK|10|24|Discipuli autem obstupescebant in verbis eius. At Iesus rursus respondens ait illis: " Filii, quam diffficile est in regnum Dei introire.
MARK|10|25|Facilius est camelum per foramen acus transire quam divitem intrare in regnum Dei ".
MARK|10|26|Qui magis admirabantur dicentes ad semetipsos: " Et quis potest salvus fieri? ".
MARK|10|27|Intuens illos Iesus ait: " Apud homines impossibile est sed non apud Deum: omnia enim possibilia sunt apud Deum ".
MARK|10|28|Coepit Petrus ei dicere: " Ecce nos dimisimus omnia et secuti sumus te.
MARK|10|29|Ait Iesus: " Amen dico vobis: Nemo est, qui reliquerit domum aut fratres aut sorores aut matrem aut patrem aut filios aut agros propter me et propter evangelium,
MARK|10|30|qui non accipiat centies tantum nunc in tempore hoc, domos et fratres et sorores et matres et filios et agros cum persecutionibus, et in saeculo futuro vitam aeternam.
MARK|10|31|Multi autem erunt primi novissimi, et novissimi primi ".
MARK|10|32|Erant autem in via ascendentes in Hierosolymam, et praecedebat illos Iesus, et stupebant; illi autem sequentes timebant. Et assumens iterum Duodecim coepit illis dicere, quae essent ei eventura:
MARK|10|33|" Ecce ascendimus in Hierosolymam; et Filius hominis tradetur principibus sacerdotum et scribis, et damnabunt eum morte et tradent eum gentibus
MARK|10|34|et illudent ei et conspuent eum et flagellabunt eum et interficient eum, et post tres dies resurget ".
MARK|10|35|Et accedunt ad eum Iacobus et Ioannes filii Zebedaei dicentes ei: " Magister, volumus, ut quodcumque petierimus a te, facias nobis ".
MARK|10|36|At ille dixit eis: " Quid vultis, ut faciam vobis? ".
MARK|10|37|Illi autem dixerunt ei: " Da nobis, ut unus ad dexteram tuam et alius ad sinistram sedeamus in gloria tua ".
MARK|10|38|Iesus autem ait eis: " Nescitis quid petatis. Potestis bibere calicem, quem ego bibo, aut baptismum, quo ego baptizor, baptizari? ".
MARK|10|39|At illi dixerunt ei: " Possumus ". Iesus autem ait eis: " Calicem quidem, quem ego bibo, bibetis et baptismum, quo ego baptizor, baptizabimini;
MARK|10|40|sedere autem ad dexteram meam vel ad sinistram non est meum dare, sed quibus paratum est ".
MARK|10|41|Et audientes decem coeperunt indignari de Iacobo et Ioanne.
MARK|10|42|Et vocans eos Iesus ait illis: " Scitis quia hi, qui videntur principari gentibus, dominantur eis, et principes eorum potestatem habent ipsorum.
MARK|10|43|Non ita est autem in vobis, sed quicumque voluerit fieri maior inter vos, erit vester minister;
MARK|10|44|et, quicumque voluerit in vobis primus esse, erit omnium servus;
MARK|10|45|nam et Filius hominis non venit, ut ministraretur ei, sed ut ministraret et daret animam suam redemptionem pro multis ".
MARK|10|46|Et veniunt Ierichum. Et proficiscente eo de Iericho et discipulis eius et plurima multitudine, filius Timaei Bartimaeus caecus sedebat iuxta viam mendicans.
MARK|10|47|Qui cum audisset quia Iesus Nazarenus est, coepit clamare et dicere: " Fili David Iesu, miserere mei! ".
MARK|10|48|Et comminabantur ei multi, ut taceret; at ille multo magis clamabat: " Fili David, miserere mei! ".
MARK|10|49|Et stans Iesus dixit: " Vocate illum ". Et vocant caecum dicentes ei: " Animaequior esto. Surge, vocat te ".
MARK|10|50|Qui, proiecto vestimento suo, exsiliens venit ad Iesum.
MARK|10|51|Et respondens ei Iesus dixit: " Quid vis tibi faciam? ". Caecus autem dixit ei: " Rabboni, ut videam ".
MARK|10|52|Et Iesus ait illi: " Vade; fides tua te salvum fecit ". Et confestim vidit et sequebatur eum in via.
MARK|11|1|Et cum appropinquarent Hierosolymae, Bethphage et Bethaniae ad montem Olivarum, mittit duos ex discipulis suis
MARK|11|2|et ait illis: " Ite in castellum, quod est contra vos, et statim introeuntes illud invenietis pullum ligatum, super quem nemo adhuc hominum sedit; solvite illum et adducite.
MARK|11|3|Et si quis vobis dixerit: "Quid facitis hoc?", dicite: "Domino necessarius est, et continuo illum remittit iterum huc" ".
MARK|11|4|Et abeuntes invenerunt pullum ligatum ante ianuam foris in bivio et solvunt eum.
MARK|11|5|Et quidam de illic stantibus dicebant illis: " Quid facitis solventes pullum? ".
MARK|11|6|Qui dixerunt eis, sicut dixerat Iesus; et dimiserunt eis.
MARK|11|7|Et ducunt pullum ad Iesum et imponunt illi vestimenta sua; et sedit super eum.
MARK|11|8|Et multi vestimenta sua straverunt in via, alii autem frondes, quas exciderant in agris.
MARK|11|9|Et qui praeibant et qui sequebantur, clamabant: " Hosanna! Benedictus, qui venit in nomine Domini!
MARK|11|10|Benedictum, quod venit regnum patris nostri David! Hosanna in excelsis!.
MARK|11|11|Et introivit Hierosolymam in templum; et circumspectis omnibus, cum iam vespera esset hora, exivit in Bethaniam cum Duodecim.
MARK|11|12|Et altera die cum exirent a Bethania, esuriit.
MARK|11|13|Cumque vidisset a longe ficum habentem folia, venit si quid forte inveniret in ea; et cum venisset ad eam, nihil invenit praeter folia: non enim erat tempus ficorum.
MARK|11|14|Et respondens dixit ei: " Iam non amplius in aeternum quisquam fructum ex te manducet ". Et audiebant discipuli eius.
MARK|11|15|Et veniunt Hierosolymam. Et cum introisset in templum, coepit eicere vendentes et ementes in templo et mensas nummulariorum et cathedras vendentium columbas evertit;
MARK|11|16|et non sinebat, ut quisquam vas transferret per templum.
MARK|11|17|Et docebat dicens eis: " Non scriptum est: "Domus mea domus orationis vocabitur omnibus gentibus"? Vos autem fecistis eam speluncam latronum ".
MARK|11|18|Quo audito, principes sacerdotum et scribae quaerebant quomodo eum perderent; timebant enim eum, quoniam universa turba admirabatur super doctrina eius.
MARK|11|19|Et cum vespera facta esset, egrediebantur de civitate.
MARK|11|20|Et cum mane transirent, viderunt ficum aridam factam a radicibus.
MARK|11|21|Et recordatus Petrus dicit ei: " Rabbi, ecce ficus, cui maledixisti, aruit ".
MARK|11|22|Et respondens Iesus ait illis: " Habete fidem Dei!
MARK|11|23|Amen dico vobis: Quicumque dixerit huic monti: "Tollere et mittere in mare", et non haesitaverit in corde suo, sed crediderit quia, quod dixerit, fiat, fiet ei.
MARK|11|24|Propterea dico vobis: Omnia, quaecumque orantes petitis, credite quia iam accepistis, et erunt vobis.
MARK|11|25|Et cum statis in oratione, dimittite, si quid habetis adversus aliquem, ut etPater vester, qui in caelis est, dimittat vobis peccata vestra ".
MARK|11|26|()
MARK|11|27|Et veniunt rursus Hierosolymam. Et cum ambularet in templo, accedunt ad eum summi sacerdotes et scribae et seniores
MARK|11|28|et dicebant illi: " In qua potestate haec facis? Vel quis tibi dedit hanc potestatem, ut ista facias? ".
MARK|11|29|Iesus autem ait illis: " Interrogabo vos unum verbum, et respondete mihi; et dicam vobis, in qua potestate haec faciam:
MARK|11|30|Baptismum Ioannis de caelo erat an ex hominibus? Respondete mihi ".
MARK|11|31|At illi cogitabant secum dicentes: " Si dixerimus: "De caelo", dicet: Quare ergo non credidistis ei?";
MARK|11|32|si autem dixerimus: "Ex hominibus?" ". Timebant populum: omnes enim habebant Ioannem quia vere propheta esset.
MARK|11|33|Et respondentes dicunt Iesu: " Nescimus ". Et Iesus ait illis: " Neque ego dico vobis in qua potestate haec faciam ".
MARK|12|1|Et coepit illis in parabolis loqui: " Vineam pastinavit ho mo et circumdedit saepem et fodit lacum et aedificavit turrim et locavit eam agricolis et peregre profectus est.
MARK|12|2|Et misit ad agricolas in tempore servum, ut ab agricolis acciperet de fructu vineae;
MARK|12|3|qui apprehensum eum caeciderunt et dimiserunt vacuum.
MARK|12|4|Et iterum misit ad illos alium servum; et illum in capite vulneraverunt et contumeliis affecerunt.
MARK|12|5|Et alium misit, et illum occiderunt, et plures alios, quosdam caedentes, alios vero occidentes.
MARK|12|6|Adhuc unum habebat, filium dilectum. Misit illum ad eos novissimum dicens: "Reverebuntur filium meum".
MARK|12|7|Coloni autem illi dixerunt ad invicem: "Hic est heres. Venite, occidamus eum, et nostra erit hereditas".
MARK|12|8|Et apprehendentes eum occiderunt et eiecerunt extra vineam.
MARK|12|9|Quid ergo faciet dominus vineae? Veniet et perdet colonos et dabit vineam aliis.
MARK|12|10|Nec Scripturam hanc legistis: "Lapidem quem reprobaverunt aedificantes,hic factus est in caput anguli;
MARK|12|11|a Domino factum est istudet est mirabile in oculis nostris"? ".
MARK|12|12|Et quaerebant eum tenere et timuerunt turbam; cognoverunt enim quoniam ad eos parabolam hanc dixerit. Et relicto eo abierunt.
MARK|12|13|Et mittunt ad eum quosdam ex pharisaeis et herodianis, ut eum caperent in verbo.
MARK|12|14|Qui venientes dicunt ei: " Magister, scimus quia verax es et non curas quemquam; nec enim vides in faciem hominum, sed in veritate viam Dei doces. Licet dare tributum Caesari an non? Dabimus an non dabimus? ".
MARK|12|15|Qui sciens versutiam eorum ait illis: " Quid me tentatis? Afferte mihi denarium, ut videam ".
MARK|12|16|At illi attulerunt. Et ait illis: " Cuius est imago haec et inscriptio?. Illi autem dixerunt ei: " Caesaris ".
MARK|12|17|Iesus autem dixit illis: " Quae sunt Caesaris, reddite Caesari et, quae sunt Dei, Deo ". Et mirabantur super eo.
MARK|12|18|Et veniunt ad eum sadducaei, qui dicunt resurrectionem non esse, et interrogabant eum dicentes:
MARK|12|19|" Magister, Moyses nobis scripsit, ut si cuius frater mortuus fuerit et reliquerit uxorem et filium non reliquerit, accipiat frater eius uxorem et resuscitet semen fratri suo.
MARK|12|20|Septem fratres erant: et primus accepit uxorem et moriens non reliquit semen;
MARK|12|21|et secundus accepit eam et mortuus est, non relicto semine; et tertius similiter;
MARK|12|22|et septem non reliquerunt semen. Novissima omnium defuncta est et mulier.
MARK|12|23|In resurrectione, cum resurrexerint, cuius de his erit uxor? Septem enim habuerunt eam uxorem ".
MARK|12|24|Ait illis Iesus: " Non ideo erratis, quia non scitis Scripturas neque virtutem Dei?
MARK|12|25|Cum enim a mortuis resurrexerint, neque nubent neque nubentur, sed sunt sicut angeli in caelis.
MARK|12|26|De mortuis autem quod resurgant, non legistis in libro Moysis super rubum, quomodo dixerit illi Deus inquiens: "Ego sum Deus Abraham et Deus Isaac et Deus Iacob"?
MARK|12|27|Non est Deus mortuorum sed vivorum! Multum erratis ".
MARK|12|28|Et accessit unus de scribis, qui audierat illos conquirentes, videns quoniam bene illis responderit, interrogavit eum: " Quod est primum omnium mandatum? ".
MARK|12|29|Iesus respondit: " Primum est: "Audi, Israel: Dominus Deus noster Dominus unus est,
MARK|12|30|et diliges Dominum Deum tuum ex toto corde tuo et ex tota anima tua et ex tota mente tua et ex tota virtute tua".
MARK|12|31|Secundum est illud: "Diliges proximum tuum tamquam teipsum". Maius horum aliud mandatum non est ".
MARK|12|32|Et ait illi scriba: " Bene, Magister, in veritate dixisti: "Unus est, et non est alius praeter eum;
MARK|12|33|et diligere eum ex toto corde et ex toto intellectu et ex tota fortitudine" et: "Diligere proximum tamquam seipsum" maius est omnibus holocautomatibus et sacrificiis ".
MARK|12|34|Et Iesus videns quod sapienter respondisset, dixit illi: " Non es longe a regno Dei ". Et nemo iam audebat eum interrogare.
MARK|12|35|Et respondens Iesus dicebat docens in templo: " Quomodo dicunt scribae Christum filium esse David?
MARK|12|36|Ipse David dixit in Spiritu Sancto:Dixit Dominus Domino meo: Sede a dextris meis,donec ponam inimicos tuos sub pedibus tuis".
MARK|12|37|Ipse David dicit eum Dominum, et unde est filius eius? ". Et multa turba eum libenter audiebat.
MARK|12|38|Et dicebat in doctrina sua: " Cavete a scribis, qui volunt in stolis ambulare et salutari in foro
MARK|12|39|et in primis cathedris sedere in synagogis et primos discubitus in cenis;
MARK|12|40|qui devorant domos viduarum et ostentant prolixas orationes. Hi accipient amplius iudicium ".
MARK|12|41|Et sedens contra gazophylacium aspiciebat quomodo turba iactaret aes in gazophylacium; et multi divites iactabant multa.
MARK|12|42|Et cum venisset una vidua pauper, misit duo minuta, quod est quadrans.
MARK|12|43|Et convocans discipulos suos ait illis: " Amen dico vobis: Vidua haec pauper plus omnibus misit, qui miserunt in gazophylacium:
MARK|12|44|Omnes enim ex eo, quod abundabat illis, miserunt; haec vero de penuria sua omnia, quae habuit, misit, totum victum suum ".
MARK|13|1|Et cum egrederetur de tem plo, ait illi unus ex discipulis suis: " Magister, aspice quales lapides et quales structurae ".
MARK|13|2|Et Iesus ait illi: " Vides has magnas aedificationes? Hic non relinquetur lapis super lapidem, qui non destruatur ".
MARK|13|3|Et cum sederet in montem Olivarum contra templum, interrogabat eum separatim Petrus et Iacobus et Ioannes et Andreas:
MARK|13|4|" Dic nobis: Quando ista erunt, et quod signum erit, quando haec omnia incipient consummari? ".
MARK|13|5|Iesus autem coepit dicere illis: " Videte, ne quis vos seducat.
MARK|13|6|Multi venient in nomine meo dicentes: "Ego sum", et multos seducent.
MARK|13|7|Cum audieritis autem bella et opiniones bellorum, ne timueritis; oportet fieri sed nondum finis.
MARK|13|8|Exsurget enim gens super gentem, et regnum super regnum, erunt terrae motus per loca, erunt fames; initium dolorum haec.
MARK|13|9|Videte autem vosmetipsos. Tradent vos conciliis, et in synagogis vapulabitis et ante praesides et reges stabitis propter me in testimonium illis.
MARK|13|10|Et in omnes gentes primum oportet praedicari evangelium.
MARK|13|11|Et cum duxerint vos tradentes, nolite praecogitare quid loquamini, sed, quod datum vobis fuerit in illa hora, id loquimini: non enim estis vos loquentes sed Spiritus Sanctus.
MARK|13|12|Et tradet frater fratrem in mortem, et pater filium; et consurgent filii in parentes et morte afficient eos;
MARK|13|13|et eritis odio omnibus propter nomen meum. Qui autem sustinuerit in finem, hic salvus erit.
MARK|13|14|Cum autem videritis abominationem desolationis stantem, ubi non debet, qui legit, intellegat: tunc, qui in Iudaea sunt, fugiant in montes;
MARK|13|15|qui autem super tectum, ne descendat nec introeat, ut tollat quid de domo sua;
MARK|13|16|et, qui in agro erit, non revertatur retro tollere vestimentum suum.
MARK|13|17|Vae autem praegnantibus et nutrientibus in illis diebus!
MARK|13|18|Orate vero, ut hieme non fiat:
MARK|13|19|erunt enim dies illi tribulatio talis, qualis non fuit ab initio creaturae, quam condidit Deus, usque nunc, neque fiet.
MARK|13|20|Et nisi breviasset Dominus dies, non fuisset salva omnis caro. Sed propter electos, quos elegit, breviavit dies.
MARK|13|21|Et tunc, si quis vobis dixerit: "Ecce hic est Christus, ecce illic", ne credideritis.
MARK|13|22|Exsurgent enim pseudochristi et pseudoprophetae et dabunt signa et portenta ad seducendos, si potest fieri, electos.
MARK|13|23|Vos autem videte; praedixi vobis omnia.
MARK|13|24|Sed in illis diebus post tribulationem illam sol contenebrabitur, et luna non dabit splendorem suum,
MARK|13|25|et erunt stellae de caelo decidentes, et virtutes, quae sunt in caelis, movebuntur.
MARK|13|26|Et tunc videbunt Filium hominis venientem in nubibus cum virtute multa et gloria.
MARK|13|27|Et tunc mittet angelos et congregabit electos suos a quattuor ventis, a summo terrae usque ad summum caeli.
MARK|13|28|A ficu autem discite parabolam: cum iam ramus eius tener fuerit et germinaverit folia, cognoscitis quia in proximo sit aestas.
MARK|13|29|Sic et vos, cum videritis haec fieri, scitote quod in proximo sit in ostiis.
MARK|13|30|Amen dico vobis: Non transiet generatio haec, donec omnia ista fiant.
MARK|13|31|Caelum et terra transibunt, verba autem mea non transibunt.
MARK|13|32|De die autem illo vel hora nemo scit, neque angeli in caelo neque Filius, nisi Pater.
MARK|13|33|Videte, vigilate; nescitis enim, quando tempus sit.
MARK|13|34|Sicut homo, qui peregre profectus reliquit domum suam et dedit servis suis potestatem, unicuique opus suum, ianitori quoque praecepit, ut vigilaret.
MARK|13|35|Vigilate ergo; nescitis enim quando dominus domus veniat, sero an media nocte an galli cantu an mane;
MARK|13|36|ne, cum venerit repente, inveniat vos dormientes.
MARK|13|37|Quod autem vobis dico, omnibus dico: Vigilate! ".
MARK|14|1|Erat autem Pascha et Azy ma post biduum. Et quaerebant summi sacerdotes et scribae, quomodo eum dolo tenerent et occiderent;
MARK|14|2|dicebant enim: " Non in die festo, ne forte tumultus fieret populi ".
MARK|14|3|Et cum esset Bethaniae in domo Simonis leprosi et recumberet, venit mulier habens alabastrum unguenti nardi puri pretiosi; fracto alabastro, effudit super caput eius.
MARK|14|4|Erant autem quidam indigne ferentes intra semetipsos: " Ut quid perditio ista unguenti facta est?
MARK|14|5|Poterat enim unguentum istud veniri plus quam trecentis denariis et dari pauperibus ". Et fremebant in eam.
MARK|14|6|Iesus autem dixit: " Sinite eam; quid illi molesti estis? Bonum opus operata est in me.
MARK|14|7|Semper enim pauperes habetis vobiscum et, cum volueritis, potestis illis bene facere; me autem non semper habetis.
MARK|14|8|Quod habuit, operata est: praevenit ungere corpus meum in sepulturam.
MARK|14|9|Amen autem dico vobis: Ubicumque praedicatum fuerit evangelium in universum mundum, et, quod fecit haec, narrabitur in memoriam eius ".
MARK|14|10|Et Iudas Iscarioth, unus de Duodecim, abiit ad summos sacerdotes, ut proderet eum illis.
MARK|14|11|Qui audientes gavisi sunt et promiserunt ei pecuniam se daturos. Et quaerebat quomodo illum opportune traderet.
MARK|14|12|Et primo die Azymorum, quando Pascha immolabant, dicunt ei discipuli eius: " Quo vis eamus et paremus, ut manduces Pascha? ".
MARK|14|13|Et mittit duos ex discipulis suis et dicit eis: " Ite in civitatem, et occurret vobis homo lagoenam aquae baiulans; sequimini eum
MARK|14|14|et, quocumque introierit, dicite domino domus: "Magister dicit: Ubi est refectio mea, ubi Pascha cum discipulis meis manducem?".
MARK|14|15|Et ipse vobis demonstrabit cenaculum grande stratum paratum; et illic parate nobis ".
MARK|14|16|Et abierunt discipuli et venerunt in civitatem et invenerunt, sicut dixerat illis, et paraverunt Pascha.
MARK|14|17|Et vespere facto, venit cum Duodecim.
MARK|14|18|Et discumbentibus eis et manducantibus, ait Iesus: " Amen dico vobis: Unus ex vobis me tradet, qui manducat mecum ".
MARK|14|19|Coeperunt contristari et dicere ei singillatim: " Numquid ego? ".
MARK|14|20|Qui ait illis: " Unus ex Duodecim, qui intingit mecum in catino.
MARK|14|21|Nam Filius quidem hominis vadit, sicut scriptum est de eo. Vae autem homini illi, per quem Filius hominis traditur! Bonum est ei, si non esset natus homo ille ".
MARK|14|22|Et manducantibus illis, accepit panem et benedicens fregit et dedit eis et ait: " Sumite: hoc est corpus meum ".
MARK|14|23|Et accepto calice, gratias agens dedit eis; et biberunt ex illo omnes.
MARK|14|24|Et ait illis: " Hic est sanguis meus novi testamenti, qui pro multis effunditur.
MARK|14|25|Amen dico vobis: Iam non bibam de genimine vitis usque in diem illum, cum illud bibam novum in regno Dei ".
MARK|14|26|Et hymno dicto, exierunt in montem Olivarum.
MARK|14|27|Et ait eis Iesus: " Omnes scandalizabimini, quia scriptum est: Percutiam pastorem, et dispergentur oves".
MARK|14|28|Sed posteaquam resurrexero, praecedam vos in Galilaeam ".
MARK|14|29|Petrus autem ait ei: " Et si omnes scandalizati fuerint, sed non ego ".
MARK|14|30|Et ait illi Iesus: " Amen dico tibi: Tu hodie, in nocte hac, priusquam bis gallus vocem dederit, ter me es negaturus ".
MARK|14|31|At ille amplius loquebatur: " Et si oportuerit me commori tibi, non te negabo ". Similiter autem et omnes dicebant.
MARK|14|32|Et veniunt in praedium, cui nomen Gethsemani; et ait discipulis suis: " Sedete hic, donec orem ".
MARK|14|33|Et assumit Petrum et Iacobum et Ioannem secum et coepit pavere et taedere;
MARK|14|34|et ait illis: " Tristis est anima mea usque ad mortem; sustinete hic et vigilate ".
MARK|14|35|Et cum processisset paululum, procidebat super terram et orabat, ut, si fieri posset, transiret ab eo hora;
MARK|14|36|et dicebat: " Abba, Pater! Omnia tibi possibilia sunt. Transfer calicem hunc a me; sed non quod ego volo, sed quod tu ".
MARK|14|37|Et venit et invenit eos dormientes; et ait Petro: " Simon, dormis? Non potuisti una hora vigilare?
MARK|14|38|Vigilate et orate, ut non intretis in tentationem; spiritus quidem promptus, caro vero infirma ".
MARK|14|39|Et iterum abiens oravit, eundem sermonem dicens.
MARK|14|40|Et veniens denuo invenit eos dormientes; erant enim oculi illorum ingravati, et ignorabant quid responderent ei.
MARK|14|41|Et venit tertio et ait illis: " Dormite iam et requiescite? Sufficit, venit hora: ecce traditur Filius hominis in manus peccatorum.
MARK|14|42|Surgite, eamus; ecce, qui me tradit, prope est ".
MARK|14|43|Et confestim, adhuc eo loquente, venit Iudas unus ex Duodecim, et cum illo turba cum gladiis et lignis a summis sacerdotibus et scribis et senioribus.
MARK|14|44|Dederat autem traditor eius signum eis dicens: " Quemcumque osculatus fuero, ipse est; tenete eum et ducite caute ".
MARK|14|45|Et cum venisset, statim accedens ad eum ait: " Rabbi "; et osculatus est eum.
MARK|14|46|At illi manus iniecerunt in eum et tenuerunt eum.
MARK|14|47|Unus autem quidam de circumstantibus educens gladium percussit servum summi sacerdotis et amputavit illi auriculam.
MARK|14|48|Et respondens Iesus ait illis: " Tamquam ad latronem existis cum gladiis et lignis comprehendere me?
MARK|14|49|Cotidie eram apud vos in templo docens, et non me tenuistis; sed adimpleantur Scripturae ".
MARK|14|50|Et relinquentes eum omnes fugerunt.
MARK|14|51|Et adulescens quidam sequebatur eum amictus sindone super nudo, et tenent eum;
MARK|14|52|at ille, reiecta sindone, nudus profugit.
MARK|14|53|Et adduxerunt Iesum ad summum sacerdotem; et conveniunt omnes summi sacerdotes et seniores et scribae.
MARK|14|54|Et Petrus a longe secutus est eum usque intro in atrium summi sacerdotis et sedebat cum ministris et calefaciebat se ad ignem.
MARK|14|55|Summi vero sacerdotes et omne concilium quaerebant adversus Iesum testimonium, ut eum morte afficerent, nec inveniebant.
MARK|14|56|Multi enim testimonium falsum dicebant adversus eum, et convenientia testimonia non erant.
MARK|14|57|Et quidam surgentes falsum testimonium ferebant adversus eum dicentes:
MARK|14|58|" Nos audivimus eum dicentem: "Ego dissolvam templum hoc manu factum et intra triduum aliud non manu factum aedificabo" ".
MARK|14|59|Et ne ita quidem conveniens erat testimonium illorum.
MARK|14|60|Et exsurgens summus sacerdos in medium interrogavit Iesum dicens: " Non respondes quidquam ad ea, quae isti testantur adversum te? ".
MARK|14|61|Ille autem tacebat et nihil respondit. Rursum summus sacerdos interrogabat eum et dicit ei: " Tu es Christus filius Benedicti? ".
MARK|14|62|Iesus autem dixit: " Ego sum, et videbitis Filium hominis a dextris sedentem Virtutis et venientem cum nubibus caeli ".
MARK|14|63|Summus autem sacerdos scindens vestimenta sua ait: " Quid adhuc necessarii sunt nobis testes?
MARK|14|64|Audistis blasphemiam. Quid vobis videtur? ". Qui omnes condemnaverunt eum esse reum mortis.
MARK|14|65|Et coeperunt quidam conspuere eum et velare faciem eius et colaphis eum caedere et dicere ei: " Prophetiza "; et ministri alapis eum caedebant.
MARK|14|66|Et cum esset Petrus in atrio deorsum, venit una ex ancillis summi sacerdotis
MARK|14|67|et, cum vidisset Petrum calefacientem se, aspiciens illum ait: " Et tu cum hoc Nazareno, Iesu, eras! ".
MARK|14|68|At ille negavit dicens: " Neque scio neque novi quid tu dicas! ". Et exiit foras ante atrium, et gallus cantavit.
MARK|14|69|Et ancilla, cum vidisset illum, rursus coepit dicere circumstantibus: " Hic ex illis est! ".
MARK|14|70|At ille iterum negabat. Et post pusillum rursus, qui astabant, dicebant Petro: " Vere ex illis es, nam et Galilaeus es ".
MARK|14|71|Ille autem coepit anathematizare et iurare: " Nescio hominem istum, quem dicitis! ".
MARK|14|72|Et statim iterum gallus cantavit; et recordatus est Petrus verbi, sicut dixerat ei Iesus: " Priusquam gallus cantet bis, ter me negabis ". Et coepit flere.
MARK|15|1|Et confestim mane consilium facientes summi sacerdotes cum senioribus et scribis, id est universum concilium, vincientes Iesum duxerunt et tradiderunt Pilato.
MARK|15|2|Et interrogavit eum Pilatus: " Tu es rex Iudaeorum? ". At ille respondens ait illi: " Tu dicis ".
MARK|15|3|Et accusabant eum summi sacerdotes in multis.
MARK|15|4|Pilatus autem rursum interrogabat eum dicens: " Non respondes quidquam? Vide in quantis te accusant ".
MARK|15|5|Iesus autem amplius nihil respondit, ita ut miraretur Pilatus.
MARK|15|6|Per diem autem festum dimittere solebat illis unum ex vinctis, quem peterent.
MARK|15|7|Erat autem qui dicebatur Barabbas, vinctus cum seditiosis, qui in seditione fecerant homicidium.
MARK|15|8|Et cum ascendisset turba, coepit rogare, sicut faciebat illis.
MARK|15|9|Pilatus autem respondit eis et dixit: " Vultis dimittam vobis regem Iudaeorum? ".
MARK|15|10|Sciebat enim quod per invidiam tradidissent eum summi sacerdotes.
MARK|15|11|Pontifices autem concitaverunt turbam, ut magis Barabbam dimitteret eis.
MARK|15|12|Pilatus autem iterum respondens aiebat illis: " Quid ergo vultis faciam regi Iudaeorum? ".
MARK|15|13|At illi iterum clamaverunt: " Crucifige eum! ".
MARK|15|14|Pilatus vero dicebat eis: " Quid enim mali fecit? ". At illi magis clamaverunt: " Crucifige eum! ".
MARK|15|15|Pilatus autem, volens populo satisfacere, dimisit illis Barabbam et tradidit Iesum flagellis caesum, ut crucifigeretur.
MARK|15|16|Milites autem duxerunt eum intro in atrium, quod est praetorium, et convocant totam cohortem.
MARK|15|17|Et induunt eum purpuram et imponunt ei plectentes spineam coronam;
MARK|15|18|et coeperunt salutare eum: " Ave, rex Iudaeorum! ",
MARK|15|19|et percutiebant caput eius arundine et conspuebant eum et ponentes genua adorabant eum.
MARK|15|20|Et postquam illuserunt ei, exuerunt illum purpuram et induerunt eum vestimentis suis. Et educunt illum, ut crucifigerent eum.
MARK|15|21|Et angariant praetereuntem quempiam Simonem Cyrenaeum venientem de villa, patrem Alexandri et Rufi, ut tolleret crucem eius.
MARK|15|22|Et perducunt illum in Golgotha locum, quod est interpretatum Calvariae locus.
MARK|15|23|Et dabant ei myrrhatum vinum; ille autem non accepit.
MARK|15|24|Et crucifigunt eum et dividunt vestimenta eius, mittentes sortem super eis, quis quid tolleret.
MARK|15|25|Erat autem hora tertia, et crucifixerunt eum.
MARK|15|26|Et erat titulus causae eius inscriptus: " Rex Iudaeorum ".
MARK|15|27|Et cum eo crucifigunt duos latrones, unum a dextris et alium asinistris eius.
MARK|15|28|()
MARK|15|29|Et praetereuntes blasphemabant eum moventes capita sua et dicentes: " Vah, qui destruit templum et in tribus diebus aedificat;
MARK|15|30|salvum fac temetipsum descendens de cruce! ".
MARK|15|31|Similiter et summi sacerdotes ludentes ad alterutrum cum scribis dicebant: " Alios salvos fecit, seipsum non potest salvum facere.
MARK|15|32|Christus rex Israel descendat nunc de cruce, ut videamus et credamus ". Etiam qui cum eo crucifixi erant, conviciabantur ei.
MARK|15|33|Et, facta hora sexta, tenebrae factae sunt per totam terram usque in horam nonam.
MARK|15|34|Et hora nona exclamavit Iesus voce magna: " Heloi, Heloi, lema sabacthani? ", quod est interpretatum: " Deus meus, Deus meus, ut quid dereliquisti me? ".
MARK|15|35|Et quidam de circumstantibus audientes dicebant: " Ecce, Eliam vocat ".
MARK|15|36|Currens autem unus et implens spongiam aceto circumponensque calamo potum dabat ei dicens: " Sinite, videamus, si veniat Elias ad deponendum eum ".
MARK|15|37|Iesus autem, emissa voce magna, exspiravit.
MARK|15|38|Et velum templi scissum est in duo a sursum usque deorsum.
MARK|15|39|Videns autem centurio, qui ex adverso stabat, quia sic clamans exspirasset, ait: " Vere homo hic Filius Dei erat ".
MARK|15|40|Erant autem et mulieres de longe aspicientes, inter quas et Maria Magdalene et Maria Iacobi minoris et Iosetis mater et Salome,
MARK|15|41|quae, cum esset in Galilaea, sequebantur eum et ministrabant ei, et aliae multae, quae simul cum eo ascenderant Hierosolymam.
MARK|15|42|Et cum iam sero esset factum, quia erat Parasceve, quod est ante sabbatum,
MARK|15|43|venit Ioseph ab Arimathaea nobilis decurio, qui et ipse erat exspectans regnum Dei, et audacter introivit ad Pilatum et petiit corpus Iesu.
MARK|15|44|Pilatus autem miratus est si iam obisset, et, accersito centurione, interrogavit eum si iam mortuus esset,
MARK|15|45|et, cum cognovisset a centurione, donavit corpus Ioseph.
MARK|15|46|Is autem mercatus sindonem et deponens eum involvit sindone et posuit eum in monumento, quod erat excisum de petra, et advolvit lapidem ad ostium monumenti.
MARK|15|47|Maria autem Magdalene et Maria Iosetis aspiciebant, ubi positus esset.
MARK|16|1|Et cum transisset sabbatum, Maria Magdalene et Maria Iacobi et Salome emerunt aromata, ut venientes ungerent eum.
MARK|16|2|Et valde mane, prima sabbatorum, veniunt ad monumentum, orto iam sole.
MARK|16|3|Et dicebant ad invicem: " Quis revolvet nobis lapidem ab ostio monumenti? ".
MARK|16|4|Et respicientes vident revolutum lapidem; erat quippe magnus valde.
MARK|16|5|Et introeuntes in monumentum viderunt iuvenem sedentem in dextris, coopertum stola candida, et obstupuerunt.
MARK|16|6|Qui dicit illis: " Nolite expavescere! Iesum quaeritis Nazarenum crucifixum. Surrexit, non est hic; ecce locus, ubi posuerunt eum.
MARK|16|7|Sed ite, dicite discipulis eius et Petro: "Praecedit vos in Galilaeam. Ibi eum videbitis, sicut dixit vobis" ".
MARK|16|8|Et exeuntes fugerunt de monumento; invaserat enim eas tremor et pavor, et nemini quidquam dixerunt, timebant enim.
MARK|16|9|Surgens autem mane, prima sabbati, apparuit primo Mariae Magdalenae, de qua eiecerat septem daemonia.
MARK|16|10|Illa vadens nuntiavit his, qui cum eo fuerant, lugentibus et flentibus;
MARK|16|11|et illi audientes quia viveret et visus esset ab ea, non crediderunt.
MARK|16|12|Post haec autem duobus ex eis ambulantibus ostensus est in alia effigie euntibus in villam;
MARK|16|13|et illi euntes nuntiaverunt ceteris, nec illis crediderunt.
MARK|16|14|Novissime recumbentibus illis Undecim apparuit, et exprobravit incredulitatem illorum et duritiam cordis, quia his, qui viderant eum resuscitatum, non crediderant.
MARK|16|15|Et dixit eis: " Euntes in mundum universum praedicate evangelium omni creaturae.
MARK|16|16|Qui crediderit et baptizatus fuerit, salvus erit; qui vero non crediderit, condemnabitur.
MARK|16|17|Signa autem eos, qui crediderint, haec sequentur: in nomine meo daemonia eicient, linguis loquentur novis,
MARK|16|18|serpentes tollent, et, si mortiferum quid biberint, non eos nocebit, super aegrotos manus imponent, et bene habebunt ".
MARK|16|19|Et Dominus quidem Iesus, postquam locutus est eis, assumptus est in caelum et sedit a dextris Dei.
MARK|16|20|Illi autem profecti praedicaverunt ubique, Domino cooperante et sermonem confirmante, sequentibus signis.
LUKE|1|1|Quoniam quidem multi conati sunt ordinare narrationem, quae in nobis completae sunt, rerum,
LUKE|1|2|sicut tradiderunt nobis, qui ab initio ipsi viderunt et ministri fuerunt verbi,
LUKE|1|3|visum est et mihi, adsecuto a principio omnia, diligenter ex ordine tibi scribere, optime Theophile,
LUKE|1|4|ut cognoscas eorum verborum, de quibus eruditus es, firmitatem.
LUKE|1|5|Fuit in diebus Herodis regis Iudaeae sacerdos quidam nomine Zacharias de vice Abiae, et uxor illi de filiabus Aaron, et nomen eius Elisabeth.
LUKE|1|6|Erant autem iusti ambo ante Deum, incedentes in omnibus mandatis et iustificationibus Domini, irreprehensibiles.
LUKE|1|7|Et non erat illis filius, eo quod esset Elisabeth sterilis, et ambo processissent in diebus suis.
LUKE|1|8|Factum est autem, cum sacerdotio fungeretur in ordine vicis suae ante Deum,
LUKE|1|9|secundum consuetudinem sacerdotii sorte exiit, ut incensum poneret ingressus in templum Domini;
LUKE|1|10|et omnis multitudo erat populi orans foris hora incensi.
LUKE|1|11|Apparuit autem illi angelus Domini stans a dextris altaris incensi;
LUKE|1|12|et Zacharias turbatus est videns, et timor irruit super eum.
LUKE|1|13|Ait autem ad illum angelus: " Ne timeas, Zacharia, quoniam exaudita est deprecatio tua, et uxor tua Elisabeth pariet tibi filium, et vocabis nomen eius Ioannem.
LUKE|1|14|Et erit gaudium tibi et exsultatio, et multi in nativitate eius gaudebunt:
LUKE|1|15|erit enim magnus coram Domino et vinum et siceram non bibet et Spiritu Sancto replebitur adhuc ex utero matris suae
LUKE|1|16|et multos filiorum Israel convertet ad Dominum Deum ipsorum.
LUKE|1|17|Et ipse praecedet ante illum in spiritu et virtute Eliae, ut convertat corda patrum in filios et incredibiles ad prudentiam iustorum, parare Domino plebem perfectam ".
LUKE|1|18|Et dixit Zacharias ad angelum: " Unde hoc sciam? Ego enim sum senex, et uxor mea processit in diebus suis ".
LUKE|1|19|Et respondens angelus dixit ei: " Ego sum Gabriel, qui adsto ante Deum, et missus sum loqui ad te et haec tibi evangelizare.
LUKE|1|20|Et ecce: eris tacens et non poteris loqui usque in diem, quo haec fiant, pro eo quod non credidisti verbis meis, quae implebuntur in tempore suo ".
LUKE|1|21|Et erat plebs exspectans Zachariam, et mirabantur quod tardaret ipse in templo.
LUKE|1|22|Egressus autem non poterat loqui ad illos, et cognoverunt quod visionem vidisset in templo; et ipse erat innuens illis et permansit mutus.
LUKE|1|23|Et factum est, ut impleti sunt dies officii eius, abiit in domum suam.
LUKE|1|24|Post hos autem dies concepit Elisabeth uxor eius et occultabat se mensibus quinque dicens:
LUKE|1|25|" Sic mihi fecit Dominus in diebus, quibus respexit auferre opprobrium meum inter homines ".
LUKE|1|26|In mense autem sexto missus est angelus Gabriel a Deo in civitatem Galilaeae, cui nomen Nazareth,
LUKE|1|27|ad virginem desponsatam viro, cui nomen erat Ioseph de domo David, et nomen virginis Maria.
LUKE|1|28|Et ingressus ad eam dixit: " Ave, gratia plena, Dominus tecum ".
LUKE|1|29|Ipsa autem turbata est in sermone eius et cogitabat qualis esset ista salutatio.
LUKE|1|30|Et ait angelus ei: " Ne timeas, Maria; invenisti enim gratiam apud Deum.
LUKE|1|31|Et ecce concipies in utero et paries filium et vocabis nomen eius Iesum.
LUKE|1|32|Hic erit magnus et Filius Altissimi vocabitur, et dabit illi Dominus Deus sedem David patris eius,
LUKE|1|33|et regnabit super domum Iacob in aeternum, et regni eius non erit finis.
LUKE|1|34|Dixit autem Maria ad angelum: " Quomodo fiet istud, quoniam virum non cognosco? ".
LUKE|1|35|Et respondens angelus dixit ei: " Spiritus Sanctus superveniet in te, et virtus Altissimi obumbrabit tibi: ideoque et quod nascetur sanctum, vocabitur Filius Dei.
LUKE|1|36|Et ecce Elisabeth cognata tua et ipsa concepit filium in senecta sua, et hic mensis est sextus illi, quae vocatur sterilis,
LUKE|1|37|quia non erit impossibile apud Deum omne verbum ".
LUKE|1|38|Dixit autem Maria: " Ecce ancilla Domini; fiat mihi secundum verbum tuum ". Et discessit ab illa angelus.
LUKE|1|39|Exsurgens autem Maria in diebus illis abiit in montana cum festinatione in civitatem Iudae
LUKE|1|40|et intravit in domum Zachariae et salutavit Elisabeth.
LUKE|1|41|Et factum est, ut audivit salutationem Mariae Elisabeth, exsultavit infans in utero eius, et repleta est Spiritu Sancto Elisabeth
LUKE|1|42|et exclamavit voce magna et dixit: " Benedicta tu inter mulieres, et benedictus fructus ventris tui.
LUKE|1|43|Et unde hoc mihi, ut veniat mater Domini mei ad me?
LUKE|1|44|Ecce enim ut facta est vox salutationis tuae in auribus meis, exsultavit in gaudio infans in utero meo.
LUKE|1|45|Et beata, quae credidit, quoniam perficientur ea, quae dicta sunt ei a Domino ".
LUKE|1|46|Et ait Maria: Magnificat anima mea Dominum,
LUKE|1|47|et exsultavit spiritus meus in Deo salvatore meo,
LUKE|1|48|quia respexit humilitatem ancillae suae.Ecce enim ex hoc beatam me dicent omnes generationes,
LUKE|1|49|quia fecit mihi magna, qui potens est,et sanctum nomen eius,
LUKE|1|50|et misericordia eius in progenies et progeniestimentibus eum.
LUKE|1|51|Fecit potentiam in brachio suo,dispersit superbos mente cordis sui;
LUKE|1|52|deposuit potentes de sedeet exaltavit humiles;
LUKE|1|53|esurientes implevit boniset divites dimisit inanes.
LUKE|1|54|Suscepit Israel puerum suum,recordatus misericordiae,
LUKE|1|55|sicut locutus est ad patres nostros,Abraham et semini eius in saecula ".
LUKE|1|56|Mansit autem Maria cum illa quasi mensibus tribus et reversa est in domum suam.
LUKE|1|57|Elisabeth autem impletum est tempus pariendi, et peperit filium.
LUKE|1|58|Et audierunt vicini et cognati eius quia magnificavit Dominus misericordiam suam cum illa, et congratulabantur ei.
LUKE|1|59|Et factum est, in die octavo venerunt circumcidere puerum et vocabant eum nomine patris eius, Zachariam.
LUKE|1|60|Et respondens mater eius dixit: " Nequaquam, sed vocabitur Ioannes ".
LUKE|1|61|Et dixerunt ad illam: " Nemo est in cognatione tua, qui vocetur hoc nomine ".
LUKE|1|62|Innuebant autem patri eius quem vellet vocari eum.
LUKE|1|63|Et postulans pugillarem scripsit dicens: " Ioannes est nomen eius ". Et mirati sunt universi.
LUKE|1|64|Apertum est autem ilico os eius et lingua eius, et loquebatur benedicens Deum.
LUKE|1|65|Et factus est timor super omnes vicinos eorum, et super omnia montana Iudaeae divulgabantur omnia verba haec.
LUKE|1|66|Et posuerunt omnes, qui audierant, in corde suo dicentes: " Quid putas puer iste erit? ". Etenim manus Domini erat cum illo.
LUKE|1|67|Et Zacharias pater eius impletus est Spiritu Sancto et prophetavit dicens:
LUKE|1|68|" Benedictus Dominus, Deus Israel,quia visitavit et fecit redemptionem plebi suae
LUKE|1|69|et erexit cornu salutis nobisin domo David pueri sui,
LUKE|1|70|sicut locutus est per os sanctorum,qui a saeculo sunt, prophetarum eius,
LUKE|1|71|salutem ex inimicis nostriset de manu omnium, qui oderunt nos;
LUKE|1|72|ad faciendam misericordiam cum patribus nostriset memorari testamenti sui sancti,
LUKE|1|73|iusiurandum, quod iuravit ad Abraham patrem nostrum,daturum se nobis,
LUKE|1|74|ut sine timore, de manu inimicorum liberati,serviamus illi
LUKE|1|75|in sanctitate et iustitia coram ipsoomnibus diebus nostris.
LUKE|1|76|Et tu, puer, propheta Altissimi vocaberis:praeibis enim ante faciem Domini parare vias eius,
LUKE|1|77|ad dandam scientiam salutis plebi eiusin remissionem peccatorum eorum,
LUKE|1|78|per viscera misericordiae Dei nostri,in quibus visitabit nos oriens ex alto,
LUKE|1|79|illuminare his, qui in tenebris et in umbra mortis sedent,ad dirigendos pedes nostros in viam pacis ".
LUKE|1|80|Puer autem crescebat et confortabatur spiritu et erat in deserto usque in diem ostensionis suae ad Israel.
LUKE|2|1|Factum est autem, in diebus il lis exiit edictum a Caesare Au gusto, ut describeretur universus orbis.
LUKE|2|2|Haec descriptio prima facta est praeside Syriae Quirino.
LUKE|2|3|Et ibant omnes, ut profiterentur, singuli in suam civitatem.
LUKE|2|4|Ascendit autem et Ioseph a Galilaea de civitate Nazareth in Iudaeam in civitatem David, quae vocatur Bethlehem, eo quod esset de domo et familia David,
LUKE|2|5|ut profiteretur cum Maria desponsata sibi, uxore praegnante.
LUKE|2|6|Factum est autem, cum essent ibi, impleti sunt dies, ut pareret,
LUKE|2|7|et peperit filium suum primogenitum; et pannis eum involvit et reclinavit eum in praesepio, quia non erat eis locus in deversorio.
LUKE|2|8|Et pastores erant in regione eadem vigilantes et custodientes vigilias noctis supra gregem suum.
LUKE|2|9|Et angelus Domini stetit iuxta illos, et claritas Domini circumfulsit illos, et timuerunt timore magno.
LUKE|2|10|Et dixit illis angelus: " Nolite timere; ecce enim evangelizo vobis gaudium magnum, quod erit omni populo,
LUKE|2|11|quia natus est vobis hodie Salvator, qui est Christus Dominus, in civitate David.
LUKE|2|12|Et hoc vobis signum: invenietis infantem pannis involutum et positum in praesepio ".
LUKE|2|13|Et subito facta est cum angelo multitudo militiae caelestis laudantium Deum et dicentium:
LUKE|2|14|" Gloria in altissimis Deo,et super terram pax in hominibus bonae voluntatis ".
LUKE|2|15|Et factum est, ut discesserunt ab eis angeli in caelum, pastores loquebantur ad invicem: " Transeamus usque Bethlehem et videamus hoc verbum, quod factum est, quod Dominus ostendit nobis ".
LUKE|2|16|Et venerunt festinantes et invenerunt Mariam et Ioseph et infantem positum in praesepio.
LUKE|2|17|Videntes autem notum fecerunt verbum, quod dictum erat illis de puero hoc.
LUKE|2|18|Et omnes, qui audierunt, mirati sunt de his, quae dicta erant a pastoribus ad ipsos.
LUKE|2|19|Maria autem conservabat omnia verba haec conferens in corde suo.
LUKE|2|20|Et reversi sunt pastores glorificantes et laudantes Deum in omnibus, quae audierant et viderant, sicut dictum est ad illos.
LUKE|2|21|Et postquam consummati sunt dies octo, ut circumcideretur, vocatum est nomen eius Iesus, quod vocatum est ab angelo, priusquam in utero conciperetur.
LUKE|2|22|Et postquam impleti sunt dies purgationis eorum secundum legem Moysis, tulerunt illum in Hierosolymam, ut sisterent Domino,
LUKE|2|23|sicut scriptum est in lege Domini: " Omne masculinum adaperiens vulvam sanctum Domino vocabitur ",
LUKE|2|24|et ut darent hostiam secundum quod dictum est in lege Domini: par turturum aut duos pullos columbarum.
LUKE|2|25|Et ecce homo erat in Ierusalem, cui nomen Simeon, et homo iste iustus et timoratus, exspectans consolationem Israel, et Spiritus Sanctus erat super eum;
LUKE|2|26|et responsum acceperat ab Spiritu Sancto non visurum se mortem nisi prius videret Christum Domini.
LUKE|2|27|Et venit in Spiritu in templum. Et cum inducerent puerum Iesum parentes eius, ut facerent secundum consuetudinem legis pro eo,
LUKE|2|28|et ipse accepit eum in ulnas suas et benedixit Deum et dixit:
LUKE|2|29|" Nunc dimittis servum tuum, Domine,secundum verbum tuum in pace,
LUKE|2|30|quia viderunt oculi meisalutare tuum,
LUKE|2|31|quod parastiante faciem omnium populorum,
LUKE|2|32|lumen ad revelationem gentiumet gloriam plebis tuae Israel ".
LUKE|2|33|Et erat pater eius et mater mirantes super his, quae dicebantur de illo.
LUKE|2|34|Et benedixit illis Simeon et dixit ad Mariam matrem eius: " Ecce positus est hic in ruinam et resurrectionem multorum in Israel et in signum, cui contradicetur
LUKE|2|35|- et tuam ipsius animam pertransiet gladius - ut revelentur ex multis cordibus cogitationes ".
LUKE|2|36|Et erat Anna prophetissa, filia Phanuel, de tribu Aser. Haec processerat in diebus multis et vixerat cum viro annis septem a virginitate sua;
LUKE|2|37|et haec vidua usque ad annos octoginta quattuor, quae non discedebat de templo, ieiuniis et obsecrationibus serviens nocte ac die.
LUKE|2|38|Et haec ipsa hora superveniens confitebatur Deo et loquebatur de illo omnibus, qui exspectabant redemptionem Ierusalem.
LUKE|2|39|Et ut perfecerunt omnia secundum legem Domini, reversi sunt in Galilaeam in civitatem suam Nazareth.
LUKE|2|40|Puer autem crescebat et confortabatur plenus sapientia; et gratia Dei erat super illum.
LUKE|2|41|Et ibant parentes eius per omnes annos in Ierusalem in die festo Paschae.
LUKE|2|42|Et cum factus esset annorum duodecim, ascendentibus illis secundum consuetudinem diei festi,
LUKE|2|43|consummatisque diebus, cum redirent, remansit puer Iesus in Ierusalem, et non cognoverunt parentes eius.
LUKE|2|44|Existimantes autem illum esse in comitatu, venerunt iter diei et requirebant eum inter cognatos et notos;
LUKE|2|45|et non invenientes regressi sunt in Ierusalem requirentes eum.
LUKE|2|46|Et factum est, post triduum invenerunt illum in templo sedentem in medio doctorum, audientem illos et interrogantem eos;
LUKE|2|47|stupebant autem omnes, qui eum audiebant, super prudentia et responsis eius.
LUKE|2|48|Et videntes eum admirati sunt, et dixit Mater cius ad illum: " Fili, quid fecisti nobis sic? Ecce pater tuus et ego dolentes quaerebamus te ".
LUKE|2|49|Et ait ad illos: " Quid est quod me quaerebatis? Nesciebatis quia in his, quae Patris mei sunt, oportet me esse? ".
LUKE|2|50|Et ipsi non intellexerunt verbum, quod locutus est ad illos.
LUKE|2|51|Et descendit cum eis et venit Nazareth et erat subditus illis. Et mater eius conservabat omnia verba in corde suo.
LUKE|2|52|Et Iesus proficiebat sapientia et aetate et gratia apud Deum et homines.
LUKE|3|1|Anno autem quinto decimo im perii Tiberii Caesaris, procu rante Pontio Pilato Iudaeam, tetrarcha autem Galilaeae Herode, Philippo autem fratre eius tetrarcha Ituraeae et Trachonitidis regionis, et Lysania Abilinae tetrarcha,
LUKE|3|2|sub principe sacerdotum Anna et Caipha, factum est verbum Dei super Ioannem Zachariae filium in deserto.
LUKE|3|3|Et venit in omnem regionem circa Iordanem praedicans baptismum paenitentiae in remissionem peccatorum,
LUKE|3|4|sicut scriptum est in libro sermonum Isaiae prophetae: Vox clamantis in deserto:Parate viam Domini,rectas facite semitas eius.
LUKE|3|5|Omnis vallis implebitur,et omnis mons et collis humiliabitur;et erunt prava in directa,et aspera in vias planas:
LUKE|3|6|et videbit omnis caro salutare Dei" ".
LUKE|3|7|Dicebat ergo ad turbas, quae exibant, ut baptizarentur ab ipso: " Genimina viperarum, quis ostendit vobis fugere a ventura ira?
LUKE|3|8|Facite ergo fructus dignos paenitentiae et ne coeperitis dicere in vobis ipsis: "Patrem habemus Abraham"; dico enim vobis quia potest Deus de lapidibus istis suscitare Abrahae filios.
LUKE|3|9|Iam enim et securis ad radicem arborum posita est; omnis ergo arbor non faciens fructum bonum exciditur et in ignem mittitur ".
LUKE|3|10|Et interrogabant eum turbae dicentes: " Quid ergo faciemus? ".
LUKE|3|11|Respondens autem dicebat illis: " Qui habet duas tunicas, det non habenti; et, qui habet escas, similiter faciat ".
LUKE|3|12|Venerunt autem et publicani, ut baptizarentur, et dixerunt ad illum: " Magister, quid faciemus? ".
LUKE|3|13|At ille dixit ad eos: " Nihil amplius quam constitutum est vobis, faciatis ".
LUKE|3|14|Interrogabant autem eum et milites dicentes: " Quid faciemus et nos? ". Et ait illis: " Neminem concutiatis neque calumniam faciatis et contenti estote stipendiis vestris ".
LUKE|3|15|Existimante autem populo et cogitantibus omnibus in cordibus suis de Ioanne, ne forte ipse esset Christus,
LUKE|3|16|respondit Ioannes dicens omnibus: " Ego quidem aqua baptizo vos. Venit autem fortior me, cuius non sum dignus solvere corrigiam calceamentorum eius: ipse vos baptizabit in Spiritu Sancto et igni;
LUKE|3|17|cuius ventilabrum in manu eius ad purgandam aream suam et ad congregandum triticum in horreum suum, paleas autem comburet igni inexstinguibili ".
LUKE|3|18|Multa quidem et alia exhortans evangelizabat populum.
LUKE|3|19|Herodes autem tetrarcha, cum corriperetur ab illo de Herodiade uxore fratris sui et de omnibus malis, quae fecit Herodes,
LUKE|3|20|adiecit et hoc supra omnia et inclusit Ioannem in carcere.
LUKE|3|21|Factum est autem, cum baptizaretur omnis populus, et Iesu baptizato et orante, apertum est caelum,
LUKE|3|22|et descendit Spiritus Sanctus corporali specie sicut columba super ipsum; et vox de caelo facta est: " Tu es Filius meus dilectus; in te complacui mihi ".
LUKE|3|23|Et ipse Iesus erat incipiens quasi annorum triginta, ut putabatur, filius Ioseph, qui fuit Heli,
LUKE|3|24|qui fuit Matthat, qui fuit Levi, qui fuit Melchi, qui fuit Iannae, qui fuit Ioseph,
LUKE|3|25|qui fuit Matthathiae, qui fuit Amos, qui fuit Nahum, qui fuit Esli, qui fuit Naggae,
LUKE|3|26|qui fuit Maath, qui fuit Matthathiae, qui fuit Semei, qui fuit Iosech, qui fuit Ioda,
LUKE|3|27|qui fuit Ioanna, qui fuit Resa, qui fuit Zorobabel, qui fuit Salathiel, qui fuit Neri,
LUKE|3|28|qui fuit Melchi, qui fuit Addi, qui fuit Cosam, qui fuit Elmadam, qui fuit Her,
LUKE|3|29|qui fuit Iesu, qui fuit Eliezer, qui fuit Iorim, qui fuit Matthat, qui fuit Levi,
LUKE|3|30|qui fuit Simeon, qui fuit Iudae, qui fuit Ioseph, qui fuit Iona, qui fuit Eliachim,
LUKE|3|31|qui fuit Melea, qui fuit Menna, qui fuit Matthatha, qui fuit Nathan, qui fuit David,
LUKE|3|32|qui fuit Iesse, qui fuit Obed, qui fuit Booz, qui fuit Salmon, qui fuit Naasson,
LUKE|3|33|qui fuit Aminadab, qui fuit Admin, qui fuit Arni, qui fuit Esrom, qui fuit Phares, qui fuit Iudae,
LUKE|3|34|qui fuit Iacob, qui fuit Isaac, qui fuit Abrahae, qui fuit Thare, qui fuit Nachor,
LUKE|3|35|qui fuit Seruch, qui fuit Ragau, qui fuit Phaleg, qui fuit Heber, qui fuit Sala,
LUKE|3|36|qui fuit Cainan, qui fuit Arphaxad, qui fuit Sem, qui fuit Noe, qui fuit Lamech,
LUKE|3|37|qui fuit Mathusala, qui fuit Henoch, qui fuit Iared, qui fuit Malaleel, qui fuit Cainan,
LUKE|3|38|qui fuit Enos, qui fuit Seth, qui fuit Adam, qui fuit Dei.
LUKE|4|1|Iesus autem plenus Spiritu Sancto regressus est ab Iordane et agebatur in Spiritu in deserto
LUKE|4|2|diebus quadraginta et tentabatur a Diabolo. Et nihil manducavit in diebus illis et, consummatis illis, esuriit.
LUKE|4|3|Dixit autem illi Diabolus: " Si Filius Dei es, dic lapidi huic, ut panis fiat ".
LUKE|4|4|Et respondit ad illum Iesus: " Scriptum est: "Non in pane solo vivet homo" ".
LUKE|4|5|Et sustulit illum et ostendit illi omnia regna orbis terrae in momento temporis;
LUKE|4|6|et ait ei Diabolus: " Tibi dabo potestatem hanc universam et gloriam illorum, quia mihi tradita est, et, cui volo, do illam:
LUKE|4|7|tu ergo, si adoraveris coram me, erit tua omnis ".
LUKE|4|8|Et respondens Iesus dixit illi: " Scriptum est: "Dominum Deum tuum adorabis et illi soli servies" ".
LUKE|4|9|Duxit autem illum in Ierusalem et statuit eum supra pinnam templi et dixit illi: " Si Filius Dei es, mitte te hinc deorsum.
LUKE|4|10|Scriptum est enim:Angelis suis mandabit de te,ut conservent te"
LUKE|4|11|et: "In manibus tollent te,ne forte offendas ad lapidem pedem tuum" ".
LUKE|4|12|Et respondens Iesus ait illi: " Dictum est: "Non tentabis Dominum Deum tuum" ".
LUKE|4|13|Et consummata omni tentatione, Diabolus recessit ab illo usque ad tempus.
LUKE|4|14|Et regressus est Iesus in virtute Spiritus in Galilaeam. Et fama exiit per universam regionem de illo.
LUKE|4|15|Et ipse docebat in synagogis eorum et magnificabatur ab omnibus.
LUKE|4|16|Et venit Nazareth, ubi erat nutritus, et intravit secundum consuetudinem suam die sabbati in synagogam et surrexit legere.
LUKE|4|17|Et tradi tus est illi liber prophetae Isaiae; etut revolvit librum, invenit locum, ubi scriptum erat:
LUKE|4|18|" Spiritus Domini super me;propter quod unxit meevangelizare pauperibus,misit me praedicare captivis remissionemet caecis visum,dimittere confractos in remissione,
LUKE|4|19|praedicare annum Domini acceptum ".
LUKE|4|20|Et cum plicuisset librum, reddidit ministro et sedit; et omnium in synagoga oculi erant intendentes in eum.
LUKE|4|21|Coepit autem dicere ad illos: " Hodie impleta est haec Scriptura in auribus vestris ".
LUKE|4|22|Et omnes testimonium illi dabant et mirabantur in verbis gratiae, quae procedebant de ore ipsius, et dicebant: " Nonne hic filius est Ioseph? ".
LUKE|4|23|Et ait illis: " Utique dicetis mihi hanc similitudinem: "Medice, cura teipsum; quanta audivimus facta in Capharnaum, fac et hic in patria tua".
LUKE|4|24|Ait autem: " Amen dico vobis: Nemo propheta acceptus est in patria sua.
LUKE|4|25|In veritate autem dico vobis: Multae viduae erant in diebus Eliae in Israel, quando clausum est caelum annis tribus et mensibus sex, cum facta est fames magna in omni terra;
LUKE|4|26|et ad nullam illarum missus est Elias nisi in Sarepta Sidoniae ad mulierem viduam.
LUKE|4|27|Et multi leprosi erant in Israel sub Eliseo propheta; et nemo eorum mundatus est nisi Naaman Syrus ".
LUKE|4|28|Et repleti sunt omnes in synagoga ira haec audientes;
LUKE|4|29|et surrexerunt et eiecerunt illum extra civitatem et duxerunt illum usque ad supercilium montis, supra quem civitas illorum erat aedificata, ut praecipitarent eum.
LUKE|4|30|Ipse autem transiens per medium illorum ibat.
LUKE|4|31|Et descendit in Capharnaum civitatem Galilaeae. Et docebat illos sabbatis;
LUKE|4|32|et stupebant in doctrina eius, quia in potestate erat sermo ipsius.
LUKE|4|33|Et in synagoga erat homo habens spiritum daemonii immundi; et exclamavit voce magna:
LUKE|4|34|" Sine; quid nobis et tibi, Iesu Nazarene? Venisti perdere nos? Scio te qui sis: Sanctus Dei ".
LUKE|4|35|Et increpavit illi Iesus dicens: " Obmutesce et exi ab illo! ". Et cum proiecisset illum daemonium in medium, exiit ab illo nihilque illum nocuit.
LUKE|4|36|Et factus est pavor in omnibus; et colloquebantur ad invicem dicentes: Quod est hoc verbum, quia in potestate et virtute imperat immundis spiritibus, et exeunt? ".
LUKE|4|37|Et divulgabatur fama de illo in omnem locum regionis.
LUKE|4|38|Surgens autem de synagoga introivit in domum Simonis. Socrus autem Simonis tenebatur magna febri; et rogaverunt illum pro ea.
LUKE|4|39|Et stans super illam imperavit febri, et dimisit illam; et continuo surgens ministrabat illis.
LUKE|4|40|Cum sol autem occidisset, omnes, qui habebant infirmos variis languoribus, ducebant illos ad eum; at ille singulis manus imponens curabat eos.
LUKE|4|41|Exibant autem daemonia a multis clamantia et dicentia: " Tu es Filius Dei ". Et increpans non sinebat ea loqui, quia sciebant ipsum esse Christum.
LUKE|4|42|Facta autem die, egressus ibat in desertum locum; et turbae requirebant eum et venerunt usque ad ipsum et detinebant illum, ne discederet ab eis.
LUKE|4|43|Quibus ille ait: " Et aliis civitatibus oportet me evangelizare regnum Dei, quia ideo missus sum ".
LUKE|4|44|Et erat praedicans in synagogis Iudaeae.
LUKE|5|1|Factum est autem, cum turba urgeret illum et audiret verbum Dei, et ipse stabat secus stagnum Genesareth
LUKE|5|2|et vidit duas naves stantes secus stagnum; piscatores autem descenderant de illis et lavabant retia.
LUKE|5|3|Ascendens autem in unam navem, quae erat Simonis, rogavit eum a terra reducere pusillum; et sedens docebat de navicula turbas.
LUKE|5|4|Ut cessavit autem loqui, dixit ad Simonem: " Duc in altum et laxate retia vestra in capturam ".
LUKE|5|5|Et respondens Simon dixit: " Praeceptor, per totam noctem laborantes nihil cepimus; in verbo autem tuo laxabo retia ".
LUKE|5|6|Et cum hoc fecissent, concluserunt piscium multitudinem copiosam; rumpebantur autem retia eorum.
LUKE|5|7|Et annuerunt sociis, qui erant in alia navi, ut venirent et adiuvarent eos; et venerunt et impleverunt ambas naviculas, ita ut mergerentur.
LUKE|5|8|Quod cum videret Simon Petrus, procidit ad genua Iesu dicens: " Exi a me, quia homo peccator sum, Domine ".
LUKE|5|9|Stupor enim circumdederat eum et omnes, qui cum illo erant, in captura piscium, quos ceperant;
LUKE|5|10|similiter autem et Iacobum et Ioannem, filios Zebedaei, qui erant socii Simonis. Et ait ad Simonem Iesus: " Noli timere; ex hoc iam homines eris capiens ".
LUKE|5|11|Et subductis ad terram navibus, relictis omnibus, secuti sunt illum.
LUKE|5|12|Et factum est, cum esset in una civitatum, et ecce vir plenus lepra; et videns Iesum et procidens in faciem rogavit eum dicens: " Domine, si vis, potes me mundare ".
LUKE|5|13|Et extendens manum tetigit illum dicens: " Volo, mundare! "; et confestim lepra discessit ab illo.
LUKE|5|14|Et ipse praecepit illi, ut nemini diceret, sed: " Vade, ostende te sacerdoti et offer pro emundatione tua, sicut praecepit Moyses, in testimonium illis ".
LUKE|5|15|Perambulabat autem magis sermo de illo, et conveniebant turbae multae, ut audirent et curarentur ab infirmitatibus suis;
LUKE|5|16|ipse autem secedebat in desertis et orabat.
LUKE|5|17|Et factum est, in una dierum, et ipse erat docens, et erant pharisaei sedentes et legis doctores, qui venerant ex omni castello Galilaeae et Iudaeae et Ierusalem; et virtus Domini erat ei ad sanandum.
LUKE|5|18|Et ecce viri portantes in lecto hominem, qui erat paralyticus, et quaerebant eum inferre et ponere ante eum.
LUKE|5|19|Et non invenientes qua parte illum inferrent prae turba, ascenderunt supra tectum et per tegulas summiserunt illum cum lectulo in medium ante Iesum.
LUKE|5|20|Quorum fidem ut vidit, dixit: " Homo, remittuntur tibi peccata tua ".
LUKE|5|21|Et coeperunt cogitare scribae et pharisaei dicentes: " Quis est hic, qui loquitur blasphemias? Quis potest dimittere peccata nisi solus Deus?.
LUKE|5|22|Ut cognovit autem Iesus cogitationes eorum, respondens dixit ad illos: Quid cogitatis in cordibus vestris?
LUKE|5|23|Quid est facilius, dicere: "Dimittuntur tibi peccata tua", an dicere: Surge et ambula"?
LUKE|5|24|Ut autem sciatis quia Filius hominis potestatem habet in terra dimittere peccata - ait paralytico -: Tibi dico: Surge, tolle lectulum tuum et vade in domum tuam ".
LUKE|5|25|Et confestim surgens coram illis tulit, in quo iacebat, et abiit in domum suam magnificans Deum.
LUKE|5|26|Et stupor apprehendit omnes, et magnificabant Deum; et repleti sunt timore dicentes: " Vidimus mirabilia hodie ".
LUKE|5|27|Et post haec exiit et vidit publicanum nomine Levi sedentem ad teloneum et ait illi: " Sequere me ".
LUKE|5|28|Et relictis omnibus, surgens secutus est eum.
LUKE|5|29|Et fecit ei convivium magnum Levi in domo sua; et erat turba multa publicanorum et aliorum, qui cum illis erant discumbentes.
LUKE|5|30|Et murmurabant pharisaei et scribae eorum adversus discipulos eius dicentes: " Quare cum publicanis et peccatoribus manducatis et bibitis? ".
LUKE|5|31|Et respondens Iesus dixit ad illos: " Non egent, qui sani sunt, medico, sed qui male habent.
LUKE|5|32|Non veni vocare iustos sed peccatores in paenitentiam ".
LUKE|5|33|At illi dixerunt ad eum: " Discipuli Ioannis ieiunant frequenter et obsecrationes faciunt, similiter et pharisaeorum; tui autem edunt et bibunt ".
LUKE|5|34|Quibus Iesus ait: " Numquid potestis convivas nuptiarum, dum cum illis est sponsus, facere ieiunare?
LUKE|5|35|Venient autem dies; et cum ablatus fuerit ab illis sponsus, tunc ieiunabunt in illis diebus ".
LUKE|5|36|Dicebat autem et similitudinem ad illos: " Nemo abscindit commissuram a vestimento novo et immittit in vestimentum vetus; alioquin et novum rumpet, et veteri non conveniet commissura a novo.
LUKE|5|37|Et nemo mittit vinum novum in utres veteres; alioquin rumpet vinum novum utres et ipsum effundetur, et utres peribunt;
LUKE|5|38|sed vinum novum in utres novos mittendum est.
LUKE|5|39|Et nemo bibens vetus vult novum; dicit enim: "Vetus melius est!" ".
LUKE|6|1|Factum est autem in sabbato, cum transiret per sata, et velle bant discipuli eius spicas et manducabant confricantes manibus.
LUKE|6|2|Quidam autem pharisaeorum dixerunt: " Quid facitis, quod non licet in sabbatis? ".
LUKE|6|3|Et respondens Iesus ad eos dixit: " Nec hoc legistis, quod fecit David, cum esurisset ipse et qui cum eo erant?
LUKE|6|4|Quomodo intravit in domum Dei et panes propositionis sumpsit et manducavit et dedit his, qui cum ipso erant, quos non licet manducare nisi tantum sacerdotibus? ".
LUKE|6|5|Et dicebat illis: " Dominus est sabbati Filius hominis ".
LUKE|6|6|Factum est autem in alio sabbato, ut intraret in synagogam et doceret; et erat ibi homo, et manus eius dextra erat arida.
LUKE|6|7|Observabant autem illum scribae et pharisaei, si sabbato curaret, ut invenirent accusare illum.
LUKE|6|8|Ipse vero sciebat cogitationes eorum et ait homini, qui habebat manum aridam: " Surge et sta in medium ". Et surgens stetit.
LUKE|6|9|Ait autem ad illos Iesus: " Interrogo vos, si licet sabbato bene facere an male; animam salvam facere an perdere? ".
LUKE|6|10|Et circumspectis omnibus illis, dixit illi: " Extende manum tuam ". Et fecit; et restituta est manus eius.
LUKE|6|11|Ipsi autem repleti sunt insipientia et colloquebantur ad invicem quidnam facerent Iesu.
LUKE|6|12|Factum est autem in illis diebus, exiit in montem orare et erat pernoctans in oratione Dei.
LUKE|6|13|Et cum dies factus esset, vocavit discipulos suos et elegit Duodecim ex ipsis, quos et apostolos nominavit:
LUKE|6|14|Simonem, quem et cognominavit Petrum, et Andream fratrem eius et Iacobum et Ioannem et Philippum et Bartholomaeum
LUKE|6|15|et Matthaeum et Thomam et Iacobum Alphaei et Simonem, qui vocatur Zelotes,
LUKE|6|16|et Iudam Iacobi et Iudam Iscarioth, qui fuit proditor.
LUKE|6|17|Et descendens cum illis stetit in loco campestri, et turba multa discipulorum eius, et multitudo copiosa plebis ab omni Iudaea et Ierusalem et maritima Tyri et Sidonis,
LUKE|6|18|qui venerunt, ut audirent eum et sanarentur a languoribus suis; et, qui vexabantur a spiritibus immundis, curabantur.
LUKE|6|19|Et omnis turba quaerebant eum tangere, quia virtus de illo exibat et sanabat omnes.
LUKE|6|20|Et ipse, elevatis oculis suis in discipulos suos, dicebat: Beati pauperes, quia vestrum est regnum Dei.
LUKE|6|21|Beati, qui nunc esuritis, quia saturabimini.Beati, qui nunc fletis, quia ridebitis.
LUKE|6|22|Beati eritis, cum vos oderint homines et cum separaverint vos et exprobraverint et eiecerint nomen vestrum tamquam malum propter Filium hominis.
LUKE|6|23|Gaudete in illa die et exsultate, ecce enim merces vestra multa in caelo; secundum haec enim faciebant prophetis patres eorum.
LUKE|6|24|Verumtamen vae vobis divitibus, quia habetis consolationem vestram!
LUKE|6|25|Vae vobis, qui saturati estis nunc, quia esurietis!Vae vobis, qui ridetis nunc, quia lugebitis et flebitis!
LUKE|6|26|Vae, cum bene vobis dixerint omnes homines! Secundum haec enim faciebant pseudoprophetis patres eorum.
LUKE|6|27|Sed vobis dico, qui auditis: Diligite inimicos vestros, bene facite his, qui vos oderunt;
LUKE|6|28|benedicite male dicentibus vobis, orate pro calumniantibus vos.
LUKE|6|29|Ei, qui te percutit in maxillam, praebe et alteram; et ab eo, qui aufert tibi vestimentum, etiam tunicam noli prohibere.
LUKE|6|30|Omni petenti te tribue; et ab eo, qui aufert, quae tua sunt, ne repetas.
LUKE|6|31|Et prout vultis, ut faciant vobis homines, facite illis similiter.
LUKE|6|32|Et si diligitis eos, qui vos diligunt, quae vobis est gratia? Nam et peccatores diligentes se diligunt.
LUKE|6|33|Et si bene feceritis his, qui vobis bene faciunt, quae vobis est gratia? Si quidem et peccatores idem faciunt.
LUKE|6|34|Et si mutuum dederitis his, a quibus speratis recipere, quae vobis gratia est? Nam et peccatores peccatoribus fenerantur, ut recipiant aequalia.
LUKE|6|35|Verumtamen diligite inimicos vestros et bene facite et mutuum date nihil desperantes; et erit merces vestra multa, et eritis filii Altissimi, quia ipse benignus est super ingratos et malos.
LUKE|6|36|Estote misericordes, sicut et Pater vester misericors est.
LUKE|6|37|Et nolite iudicare et non iudicabimini; et nolite condemnare et non condemnabimini. Dimittite et dimittemini;
LUKE|6|38|date, et dabitur vobis: mensuram bonam, confertam, coagitatam, supereffluentem dabunt in sinum vestrum; eadem quippe mensura, qua mensi fueritis, remetietur vobis ".
LUKE|6|39|Dixit autem illis et similitudinem: " Numquid potest caecus caecum ducere? Nonne ambo in foveam cadent?
LUKE|6|40|Non est discipulus super magistrum; perfectus autem omnis erit sicut magister eius.
LUKE|6|41|Quid autem vides festucam in oculo fratris tui, trabem autem, quae in oculo tuo est, non consideras?
LUKE|6|42|Quomodo potes dicere fratri tuo: "Frater, sine eiciam festucam, quae est in oculo tuo", ipse in oculo tuo trabem non videns? Hypocrita, eice primum trabem de oculo tuo et tunc perspicies, ut educas festucam, quae est in oculo fratris tui.
LUKE|6|43|Non est enim arbor bona faciens fructum malum, neque iterum arbor mala faciens fructum bonum.
LUKE|6|44|Unaquaeque enim arbor de fructu suo cognoscitur; neque enim de spinis colligunt ficus, neque de rubo vindemiant uvam.
LUKE|6|45|Bonus homo de bono thesauro cordis profert bonum, et malus homo de malo profert malum: ex abundantia enim cordis os eius loquitur.
LUKE|6|46|Quid autem vocatis me: "Domine, Domine", et non facitis, quae dico?
LUKE|6|47|Omnis, qui venit ad me et audit sermones meos et facit eos, ostendam vobis cui similis sit:
LUKE|6|48|similis est homini aedificanti domum, qui fodit in altum et posuit fundamentum supra petram; inundatione autem facta, illisum est flumen domui illi et non potuit eam movere; bene enim aedificata erat.
LUKE|6|49|Qui autem audivit et non fecit, similis est homini aedificanti domum suam supra terram sine fundamento; in quam illisus est fluvius, et continuo cecidit, et facta est ruina domus illius magna ".
LUKE|7|1|Cum autem implesset omnia verba sua in aures plebis, intra vit Capharnaum.
LUKE|7|2|Centurionis autem cuiusdam servus male habens erat moriturus, qui illi erat pretiosus.
LUKE|7|3|Et cum audisset de Iesu, misit ad eum seniores Iudaeorum rogans eum, ut veniret et salvaret servum eius.
LUKE|7|4|At illi cum venissent ad Iesum, rogabant eum sollicite dicentes: " Dignus est, ut hoc illi praestes:
LUKE|7|5|diligit enim gentem nostram et synagogam ipse aedificavit nobis ".
LUKE|7|6|Iesus autem ibat cum illis. At cum iam non longe esset a domo, misit centurio amicos dicens ei: " Domine, noli vexari; non enim dignus sum, ut sub tectum meum intres,
LUKE|7|7|propter quod et meipsum non sum dignum arbitratus, ut venirem ad te; sed dic verbo, et sanetur puer meus.
LUKE|7|8|Nam et ego homo sum sub potestate constitutus, habens sub me milites, et dico huic: "Vade", et vadit; et alii: "Veni", et venit; et servo meo: "Fac hoc", et facit ".
LUKE|7|9|Quo audito, Iesus miratus est eum et conversus sequentibus se turbis dixit: " Dico vobis, nec in Israel tantam fidem inveni! ".
LUKE|7|10|Et reversi, qui missi fuerant, domum, invenerunt servum sanum.
LUKE|7|11|Et factum est, deinceps ivit in civitatem, quae vocatur Naim, et ibant cum illo discipuli eius et turba copiosa.
LUKE|7|12|Cum autem appropinquaret portae civitatis, et ecce defunctus efferebatur filius unicus matri suae; et haec vidua erat, et turba civitatis multa cum illa.
LUKE|7|13|Quam cum vidisset Dominus, misericordia motus super ea dixit illi: " Noli flere! ".
LUKE|7|14|Et accessit et tetigit loculum; hi autem, qui portabant, steterunt. Et ait: " Adulescens, tibi dico: Surge! ".
LUKE|7|15|Et resedit, qui erat mortuus, et coepit loqui; et dedit illum matri suae.
LUKE|7|16|Accepit autem omnes timor, et magnificabant Deum dicentes: " Propheta magnus surrexit in nobis " et: " Deus visitavit plebem suam ".
LUKE|7|17|Et exiit hic sermo in universam Iudaeam de eo et omnem circa regionem.
LUKE|7|18|Et nuntiaverunt Ioanni discipuli eius de omnibus his.
LUKE|7|19|Et convocavit duos de discipulis suis Ioannes et misit ad Dominum dicens: " Tu es qui venturus es, an alium exspectamus? ".
LUKE|7|20|Cum autem venissent ad eum viri, dixerunt: " Ioannes Baptista misit nos ad te dicens: "Tu es qui venturus es, an alium exspectamus?" ".
LUKE|7|21|In ipsa hora curavit multos a languoribus et plagis et spiritibus malis et caecis multis donavit visum.
LUKE|7|22|Et respondens dixit illis: " Euntes nuntiate Ioanni, quae vidistis et audistis: caeci vident, claudi ambulant, leprosi mundantur et surdi audiunt, mortui resurgunt, pauperes evangelizantur;
LUKE|7|23|et beatus est, quicumque non fuerit scandalizatus in me ".
LUKE|7|24|Et cum discessissent nuntii Ioannis, coepit dicere de Ioanne ad turbas: Quid existis in desertum videre? Arundinem vento moveri?
LUKE|7|25|Sed quid existis videre? Hominem mollibus vestimentis indutum? Ecce, qui in veste pretiosa sunt et deliciis, in domibus regum sunt.
LUKE|7|26|Sed quid existis videre? Prophetam? Utique, dico vobis, et plus quam prophetam.
LUKE|7|27|Hic est, de quo scriptum est:Ecce mitto angelum meum ante faciem tuam,qui praeparabit viam tuam ante te".
LUKE|7|28|Dico vobis: Maior inter natos mulierum Ioanne nemo est; qui autem minor est in regno Dei, maior est illo.
LUKE|7|29|Et omnis populus audiens et publicani iustificaverunt Deum, baptizati baptismo Ioannis;
LUKE|7|30|pharisaei autem et legis periti consilium Dei spreverunt in semetipsos, non baptizati ab eo.
LUKE|7|31|Cui ergo similes dicam homines generationis huius, et cui similes sunt?
LUKE|7|32|Similes sunt pueris sedentibus in foro et loquentibus ad invicem, quod dicit:Cantavimus vobis tibiis, et non saltastis;lamentavimus, et non plorastis!".
LUKE|7|33|Venit enim Ioannes Baptista neque manducans panem neque bibens vinum, et dicitis: "Daemonium habet!";
LUKE|7|34|venit Filius hominis manducans et bibens, et dicitis: "Ecce homo devorator et bibens vinum, amicus publicanorum et peccatorum!".
LUKE|7|35|Et iustificata est sapientia ab omnibus filiis suis ".
LUKE|7|36|Rogabat autem illum quidam de pharisaeis, ut manducaret cum illo; et ingressus domum pharisaei discubuit.
LUKE|7|37|Et ecce mulier, quae erat in civitate peccatrix, ut cognovit quod accubuit in domo pharisaei, attulit alabastrum unguenti;
LUKE|7|38|et stans retro secus pedes eius flens lacrimis coepit rigare pedes eius et capillis capitis sui tergebat, et osculabatur pedes eius et unguento ungebat.
LUKE|7|39|Videns autem pharisaeus, qui vocaverat eum, ait intra se dicens: " Hic si esset propheta, sciret utique quae et qualis mulier, quae tangit eum, quia peccatrix est ".
LUKE|7|40|Et respondens Iesus dixit ad illum: " Simon, habeo tibi aliquid dicere. At ille ait: " Magister, dic ".
LUKE|7|41|" Duo debitores erant cuidam feneratori: unus debebat denarios quingentos, alius quinquaginta.
LUKE|7|42|Non habentibus illis, unde redderent, donavit utrisque. Quis ergo eorum plus diliget eum? ".
LUKE|7|43|Respondens Simon dixit: " Aestimo quia is, cui plus donavit ". At ille dixit ei: " Recte iudicasti ".
LUKE|7|44|Et conversus ad mulierem, dixit Simoni: " Vides hanc mulierem? Intravi in domum tuam: aquam pedibus meis non dedisti; haec autem lacrimis rigavit pedes meos et capillis suis tersit.
LUKE|7|45|Osculum mihi non dedisti; haec autem, ex quo intravi, non cessavit osculari pedes meos.
LUKE|7|46|Oleo caput meum non unxisti; haec autem unguento unxit pedes meos.
LUKE|7|47|Propter quod dico tibi: Remissa sunt peccata eius multa, quoniam dilexit multum; cui autem minus dimittitur, minus diligit ".
LUKE|7|48|Dixit autem ad illam: " Remissa sunt peccata tua ".
LUKE|7|49|Et coeperunt, qui simul accumbebant, dicere intra se: " Quis est hic, qui etiam peccata dimittit?".
LUKE|7|50|Dixit autem ad mulierem: " Fides tua te salvam fecit; vade in pace! ".
LUKE|8|1|Et factum est deinceps, et ipse iter faciebat per civitatem et ca stellum praedicans et evangelizans regnum Dei; et Duodecim cum illo
LUKE|8|2|et mulieres aliquae, quae erant curatae ab spiritibus malignis et infirmitatibus: Maria, quae vocatur Magdalene, de qua daemonia septem exierant,
LUKE|8|3|et Ioanna uxor Chuza, procuratoris Herodis, et Susanna et aliae multae, quae ministrabant eis de facultatibus suis.
LUKE|8|4|Cum autem turba plurima conveniret, et de singulis civitatibus properarent ad eum, dixit per similitudinem:
LUKE|8|5|" Exiit, qui seminat, seminare semen suum. Et dum seminat ipse, aliud cecidit secus viam et conculcatum est, et volucres caeli comederunt illud.
LUKE|8|6|Et aliud cecidit super petram et natum aruit, quia non habebat umorem.
LUKE|8|7|Et aliud cecidit inter spinas, et simul exortae spinae suffocaverunt illud.
LUKE|8|8|Et aliud cecidit in terram bonam et ortum fecit fructum centuplum ". Haec dicens clamabat: " Qui habet aures audiendi, audiat ".
LUKE|8|9|Interrogabant autem eum discipuli eius, quae esset haec parabola.
LUKE|8|10|Quibus ipse dixit: " Vobis datum est nosse mysteria regni Dei, ceteris autem in parabolis, ut videntes non videant et audientes non intellegant.
LUKE|8|11|Est autem haec parabola: Semen est verbum Dei.
LUKE|8|12|Qui autem secus viam, sunt qui audiunt; deinde venit Diabolus et tollit verbum de corde eorum, ne credentes salvi fiant.
LUKE|8|13|Qui autem supra petram: qui cum audierint, cum gaudio suscipiunt verbum; et hi radices non habent, qui ad tempus credunt, et in tempore tentationis recedunt.
LUKE|8|14|Quod autem in spinis cecidit: hi sunt, qui audierunt et a sollicitudinibus et divitiis et voluptatibus vitae euntes suffocantur et non referunt fructum.
LUKE|8|15|Quod autem in bonam terram: hi sunt, qui in corde bono et optimo audientes verbum retinent et fructum afferunt in patientia.
LUKE|8|16|Nemo autem lucernam accendens operit eam vaso aut subtus lectum ponit, sed supra candelabrum ponit, ut intrantes videant lumen.
LUKE|8|17|Non enim est occultum, quod non manifestetur, nec absconditum, quod non cognoscatur et in palam veniat.
LUKE|8|18|Videte ergo quomodo audiatis: qui enim habet, dabitur illi; et, quicumque non habet, etiam quod putat se habere, auferetur ab illo ".
LUKE|8|19|Venerunt autem ad illum mater et fratres eius, et non poterant adire ad eum prae turba.
LUKE|8|20|Et nuntiatum est illi: " Mater tua et fratres tui stant foris volentes te videre ".
LUKE|8|21|Qui respondens dixit ad eos: " Mater mea et fratres mei hi sunt, qui verbum Dei audiunt et faciunt ".
LUKE|8|22|Factum est autem in una dierum, et ipse ascendit in navem et discipuli eius, et ait ad illos: " Transfretemus trans stagnum ". Et ascenderunt.
LUKE|8|23|Navigantibus autem illis, obdormivit. Et descendit procella venti in stagnum, et complebantur et periclitabantur.
LUKE|8|24|Accedentes autem suscitaverunt eum dicentes: " Praeceptor, praeceptor, perimus! ". At ille surgens increpavit ventum et tempestatem aquae, et cessaverunt, et facta est tranquillitas.
LUKE|8|25|Dixit autem illis: " Ubi est fides vestra? ". Qui timentes mirati sunt dicentes ad invicem: " Quis putas hic est, quia et ventis imperat et aquae, et oboediunt ei? ".
LUKE|8|26|Enavigaverunt autem ad regionem Gergesenorum, quae est contra Galilaeam.
LUKE|8|27|Et cum egressus esset ad terram, occurrit illi vir quidam de civitate, qui habebat daemonia et iam tempore multo vestimento non induebatur neque in domo manebat sed in monumentis.
LUKE|8|28|Is ut vidit Iesum, exclamans procidit ante illum et voce magna dixit: " Quid mihi et tibi est, Iesu, Fili Dei Altissimi? Obsecro te, ne me torqueas ".
LUKE|8|29|Praecipiebat enim spiritui immundo, ut exiret ab homine. Multis enim temporibus arripiebat illum, vinciebatur catenis et compedibus custoditus; et ruptis vinculis, agebatur a daemonio in deserta.
LUKE|8|30|Interrogavit autem illum Iesus dicens: " Quod tibi nomen est? ". At ille dixit: " Legio ", quia intraverunt daemonia multa in eum.
LUKE|8|31|Et rogabant eum, ne imperaret illis, ut in abyssum irent.
LUKE|8|32|Erat autem ibi grex porcorum multorum pascentium in monte; et rogaverunt eum, ut permitteret eis in illos ingredi. Et permisit illis.
LUKE|8|33|Exierunt ergo daemonia ab homine et intraverunt in porcos, et impetu abiit grex per praeceps in stagnum et suffocatus est.
LUKE|8|34|Quod ut viderunt factum, qui pascebant, fugerunt et nuntiaverunt in civitatem et in villas.
LUKE|8|35|Exierunt autem videre, quod factum est, et venerunt ad Iesum et invenerunt hominem sedentem, a quo daemonia exierant, vestitum ac sana mente ad pedes Iesu et timuerunt.
LUKE|8|36|Nuntiaverunt autem illis hi, qui viderant, quomodo sanus factus esset, qui a daemonio vexabatur.
LUKE|8|37|Et rogaverunt illum omnis multitudo regionis Gergesenorum, ut discederet ab ipsis, quia timore magno tenebantur. Ipse autem ascendens navem reversus est.
LUKE|8|38|Et rogabat illum vir, a quo daemonia exierant, ut cum eo esset. Dimisit autem eum dicens:
LUKE|8|39|" Redi domum tuam et narra quanta tibi fecit Deus ". Et abiit per universam civitatem praedicans quanta illi fecisset Iesus.
LUKE|8|40|Cum autem rediret Iesus, excepit illum turba; erant enim omnes exspectantes eum.
LUKE|8|41|Et ecce venit vir, cui nomen Iairus, et ipse princeps synagogae erat, et cecidit ad pedes Iesu rogans eum, ut intraret in domum eius,
LUKE|8|42|quia filia unica erat illi fere annorum duodecim, et haec moriebatur. Et dum iret, a turbis comprimebatur.
LUKE|8|43|Et mulier quaedam erat in fluxu sanguinis ab annis duodecim, quae in medicos erogaverat omnem substantiam suam nec ab ullo potuit curari;
LUKE|8|44|accessit retro et tetigit fimbriam vestimenti eius, et confestim stetit fluxus sanguinis eius.
LUKE|8|45|Et ait Iesus: " Quis est, qui me tetigit? ". Negantibus autem omnibus, dixit Petrus: " Praeceptor, turbae te comprimunt et affligunt ".
LUKE|8|46|At dixit Iesus: " Tetigit me aliquis; nam et ego novi virtutem de me exisse ".
LUKE|8|47|Videns autem mulier quia non latuit, tremens venit et procidit ante eum et ob quam causam tetigerit eum indicavit coram omni populo et quemadmodum confestim sanata sit.
LUKE|8|48|At ipse dixit illi: " Filia, fides tua te salvam fecit. Vade in pace ".
LUKE|8|49|Adhuc illo loquente, venit quidam e domo principis synagogae dicens: " Mortua est filia tua; noli amplius vexare magistrum ".
LUKE|8|50|Iesus autem, audito hoc verbo, respondit ei: " Noli timere; crede tantum, et salva erit ".
LUKE|8|51|Et cum venisset domum, non permisit intrare secum quemquam nisi Petrum et Ioannem et Iacobum et patrem puellae et matrem.
LUKE|8|52|Flebant autem omnes et plangebant illam. At ille dixit: " Nolite flere; non est enim mortua, sed dormit ".
LUKE|8|53|Et deridebant eum scientes quia mortua esset.
LUKE|8|54|Ipse autem tenens manum eius clamavit dicens: " Puella, surge! ".
LUKE|8|55|Et reversus est spiritus eius, et surrexit continuo; et iussit illi dari manducare.
LUKE|8|56|Et stupuerunt parentes eius, quibus praecepit, ne alicui dicerent, quod factum erat.
LUKE|9|1|Convocatis autem Duodecim, dedit illis virtutem et potesta tem super omnia daemonia, et ut languores curarent,
LUKE|9|2|et misit illos praedicare regnum Dei et sanare infirmos;
LUKE|9|3|et ait ad illos: " Nihil tuleritis in via, neque virgam neque peram neque panem neque pecuniam, neque duas tunicas habeatis.
LUKE|9|4|Et in quamcumque domum intraveritis, ibi manete et inde exite.
LUKE|9|5|Et quicumque non receperint vos, exeuntes de civitate illa pulverem pedum vestrorum excutite in testimonium supra illos ".
LUKE|9|6|Egressi autem circumibant per castella evangelizantes et curantes ubique.
LUKE|9|7|Audivit autem Herodes tetrarcha omnia, quae fiebant, et haesitabat, eo quod diceretur a quibusdam: " Ioannes surrexit a mortuis ";
LUKE|9|8|a quibusdam vero: " Elias apparuit "; ab aliis autem: " Propheta unus de antiquis surrexit ".
LUKE|9|9|Et ait Herodes: " Ioannem ego decollavi; quis autem est iste, de quo audio ego talia? ". Et quaerebat videre eum.
LUKE|9|10|Et reversi apostoli narraverunt illi, quaecumque fecerunt. Et assumptis illis, secessit seorsum ad civitatem, quae vocatur Bethsaida.
LUKE|9|11|Quod cum cognovissent turbae, secutae sunt illum. Et excepit illos et loquebatur illis de regno Dei et eos, qui cura indigebant, sanabat.
LUKE|9|12|Dies autem coeperat declinare; et accedentes Duodecim dixerunt illi: " Dimitte turbam, ut euntes in castella villasque, quae circa sunt, divertant et inveniant escas, quia hic in loco deserto sumus ".
LUKE|9|13|Ait autem ad illos: " Vos date illis manducare ". At illi dixerunt: " Non sunt nobis plus quam quinque panes et duo pisces, nisi forte nos eamus et emamus in omnem hanc turbam escas ".
LUKE|9|14|Erant enim fere viri quinque milia. Ait autem ad discipulos suos: " Facite illos discumbere per convivia ad quinquagenos ".
LUKE|9|15|Et ita fecerunt et discumbere fecerunt omnes.
LUKE|9|16|Acceptis autem quinque panibus et duobus piscibus, respexit in caelum et benedixit illis et fregit et dabat discipulis suis, ut ponerent ante turbam.
LUKE|9|17|Et manducaverunt et saturati sunt omnes; et sublatum est, quod superfuit illis, fragmentorum cophini duodecim.
LUKE|9|18|Et factum est, cum solus esset orans, erant cum illo discipuli, et interrogavit illos dicens: " Quem me dicunt esse turbae? ".
LUKE|9|19|At illi responderunt et dixerunt: " Ioannem Baptistam, alii autem Eliam, alii vero: Propheta unus de prioribus surrexit ".
LUKE|9|20|Dixit autem illis: " Vos autem quem me esse dicitis? ". Respondens Petrus dixit: " Christum Dei ".
LUKE|9|21|At ille increpans illos praecepit, ne cui dicerent hoc,
LUKE|9|22|dicens: " Oportet Filium hominis multa pati et reprobari a senioribus et principibus sacerdotum et scribis et occidi et tertia die resurgere ".
LUKE|9|23|Dicebat autem ad omnes: " Si quis vult post me venire, abneget semetipsum et tollat crucem suam cotidie et sequatur me.
LUKE|9|24|Qui enim voluerit animam suam salvam facere, perdet illam; qui autem perdiderit animam suam propter me, hic salvam faciet illam.
LUKE|9|25|Quid enim proficit homo, si lucretur universum mundum, se autem ipsum perdat vel detrimentum sui faciat?
LUKE|9|26|Nam qui me erubuerit et meos sermones, hunc Filius hominis erubescet, cum venerit in gloria sua et Patris et sanctorum angelorum.
LUKE|9|27|Dico autem vobis vere: Sunt aliqui hic stantes, qui non gustabunt mortem, donec videant regnum Dei ".
LUKE|9|28|Factum est autem post haec verba fere dies octo, et assumpsit Petrum et Ioannem et Iacobum et ascendit in montem, ut oraret.
LUKE|9|29|Et facta est, dum oraret, species vultus eius altera, et vestitus eius albus, refulgens.
LUKE|9|30|Et ecce duo viri loquebantur cum illo, et erant Moyses et Elias,
LUKE|9|31|qui visi in gloria dicebant exodum eius, quam completurus erat in Ierusalem.
LUKE|9|32|Petrus vero et qui cum illo gravati erant somno; et evigilantes viderunt gloriam eius et duos viros, qui stabant cum illo.
LUKE|9|33|Et factum est, cum discederent ab illo, ait Petrus ad Iesum: " Praeceptor, bonum est nos hic esse; et faciamus tria tabernacula: unum tibi et unum Moysi et unum Eliae ", nesciens quid diceret.
LUKE|9|34|Haec autem illo loquente, facta est nubes et obumbravit eos; et timuerunt intrantibus illis in nubem.
LUKE|9|35|Et vox facta est de nube dicens: " Hic est Filius meus electus; ipsum audite ".
LUKE|9|36|Et dum fieret vox, inventus est Iesus solus. Et ipsi tacuerunt et nemini dixerunt in illis diebus quidquam ex his, quae viderant.
LUKE|9|37|Factum est autem in sequenti die, descendentibus illis de monte, occurrit illi turba multa.
LUKE|9|38|Et ecce vir de turba exclamavit dicens: " Magister, obsecro te, respice in filium meum, quia unicus est mihi;
LUKE|9|39|et ecce spiritus apprehendit illum, et subito clamat, et dissipat eum cum spuma et vix discedit ab eo dilanians eum;
LUKE|9|40|et rogavi discipulos tuos, ut eicerent illum, et non potuerunt ".
LUKE|9|41|Respondens autem Iesus dixit: " O generatio infidelis et perversa, usquequo ero apud vos et patiar vos? Adduc huc filium tuum ".
LUKE|9|42|Et cum accederet, elisit illum daemonium et dissipavit. Et increpavit Iesus spiritum immundum et sanavit puerum et reddidit illum patri eius.
LUKE|9|43|Stupebant autem omnes in magnitudine Dei.Omnibusque mirantibus in omnibus, quae faciebat, dixit ad discipulos suos:
LUKE|9|44|" Ponite vos in auribus vestris sermones istos: Filius enim hominis futurum est ut tradatur in manus hominum ".
LUKE|9|45|At illi ignorabant verbum istud, et erat velatum ante eos, ut non sentirent illud, et time bant interrogare eum de hoc verbo.
LUKE|9|46|Intravit autem cogitatio in eos, quis eorum maior esset.
LUKE|9|47|At Iesus sciens cogitationem cordis illorum, apprehendens puerum statuit eum secus se
LUKE|9|48|et ait illis: " Quicumque susceperit puerum istum in nomine meo, me recipit; et, quicumque me receperit, recipit eum, qui me misit; nam qui minor est inter omnes vos, hic maior est ".
LUKE|9|49|Respondens autem Ioannes dixit: " Praeceptor, vidimus quendam in nomine tuo eicientem daemonia et prohibuimus eum, quia non sequitur nobiscum ".
LUKE|9|50|Et ait ad illum Iesus: " Nolite prohibere; qui enim non est adversus vos, pro vobis est ".
LUKE|9|51|Factum est autem, dum complerentur dies assumptionis eius, et ipse faciem suam firmavit, ut iret Ierusalem,
LUKE|9|52|et misit nuntios ante conspectum suum. Et euntes intraverunt in castellum Samaritanorum, ut pararent illi.
LUKE|9|53|Et non receperunt eum, quia facies eius erat euntis Ierusalem.
LUKE|9|54|Cum vidissent autem discipuli Iacobus et Ioannes, dixerunt: " Domine, vis dicamus, ut ignis descendat de caelo et consumat illos? ".
LUKE|9|55|Et conversus increpavit illos.
LUKE|9|56|Et ierunt in aliud castellum.
LUKE|9|57|Et euntibus illis in via, dixit quidam ad illum: " Sequar te, quocumque ieris ".
LUKE|9|58|Et ait illi Iesus: " Vulpes foveas habent, et volucres caeli nidos, Filius autem hominis non habet, ubi caput reclinet ".
LUKE|9|59|Ait autem ad alterum: " Sequere me ". Ille autem dixit: " Domine, permitte mihi primum ire et sepelire patrem meum ".
LUKE|9|60|Dixitque ei Iesus: " Sine, ut mortui sepeliant mortuos suos; tu autem vade, annuntia regnum Dei ".
LUKE|9|61|Et ait alter: " Sequar te, Domine, sed primum permitte mihi renuntiare his, qui domi sunt ".
LUKE|9|62|Ait ad illum Iesus: " Nemo mittens manum suam in aratrum et aspiciens retro, aptus est regno Dei ".
LUKE|10|1|Post haec autem designavit Dominus alios septuaginta duos et misit illos binos ante faciem suam in omnem civitatem et locum, quo erat ipse venturus.
LUKE|10|2|Et dicebat illis: " Messis quidem multa, operarii autem pauci; rogate ergo Dominum messis, ut mittat operarios in messem suam.
LUKE|10|3|Ite; ecce ego mitto vos sicut agnos inter lupos.
LUKE|10|4|Nolite portare sacculum neque peram neque calceamenta et neminem per viam salutaveritis.
LUKE|10|5|In quamcumque domum intraveritis, primum dicite: "Pax huic domui".
LUKE|10|6|Et si ibi fuerit filius pacis, requiescet super illam pax vestra; sin autem, ad vos revertetur.
LUKE|10|7|In eadem autem domo manete edentes et bibentes, quae apud illos sunt: dignus enim est operarius mercede sua. Nolite transire de domo in domum.
LUKE|10|8|Et in quamcumque civitatem intraveritis, et susceperint vos, manducate, quae apponuntur vobis,
LUKE|10|9|et curate infirmos, qui in illa sunt, et dicite illis: "Appropinquavit in vos regnum Dei".
LUKE|10|10|In quamcumque civitatem intraveritis, et non receperint vos, exeuntes in plateas eius dicite:
LUKE|10|11|"Etiam pulverem, qui adhaesit nobis ad pedes de civitate vestra, extergimus in vos; tamen hoc scitote, quia appropinquavit regnum Dei".
LUKE|10|12|Dico vobis quia Sodomis in die illa remissius erit quam illi civitati.
LUKE|10|13|Vae tibi, Chorazin! Vae tibi, Bethsaida! Quia si in Tyro et Sidone factae fuissent virtutes, quae in vobis factae sunt, olim in cilicio et cinere sedentes paeniterent.
LUKE|10|14|Verumtamen Tyro et Sidoni remissius erit in iudicio quam vobis.
LUKE|10|15|Et tu, Capharnaum, numquid usque in caelum exaltaberis? Usque ad infernum demergeris!
LUKE|10|16|Qui vos audit, me audit; et, qui vos spernit, me spernit; qui autem me spernit, spernit eum, qui me misit ".
LUKE|10|17|Reversi sunt autem septuaginta duo cum gaudio dicentes: " Domine, etiam daemonia subiciuntur nobis in nomine tuo! ".
LUKE|10|18|Et ait illis: " Videbam Satanam sicut fulgur de caelo cadentem.
LUKE|10|19|Ecce dedi vobis potestatem calcandi supra serpentes et scorpiones et supra omnem virtutem inimici; et nihil vobis nocebit.
LUKE|10|20|Verumtamen in hoc nolite gaudere, quia spiritus vobis subiciuntur; gaudete autem quod nomina vestra scripta sunt in caelis ".
LUKE|10|21|In ipsa hora exsultavit Spiritu Sancto et dixit: " Confiteor tibi, Pater, Domine caeli et terrae, quod abscondisti haec a sapientibus et prudentibus et revelasti ea parvulis; etiam, Pater, quia sic placuit ante te.
LUKE|10|22|Omnia mihi tradita sunt a Patre meo; et nemo scit qui sit Filius, nisi Pater, et qui sit Pater, nisi Filius et cui voluerit Filius revelare ".
LUKE|10|23|Et conversus ad discipulos seorsum dixit: " Beati oculi, qui vident, quae videtis.
LUKE|10|24|Dico enim vobis: Multi prophetae et reges voluerunt videre, quae vos videtis, et non viderunt, et audire, quae auditis, et non audierunt ".
LUKE|10|25|Et ecce quidam legis peritus surrexit tentans illum dicens: " Magister, quid faciendo vitam aeternam possidebo? ".
LUKE|10|26|At ille dixit ad eum: " In Lege quid scriptum est? Quomodo legis? ".
LUKE|10|27|Ille autem respondens dixit: " Diliges Dominum Deum tuum ex toto corde tuo et ex tota anima tua et ex omnibus viribus tuis et ex omni mente tua et proximum tuum sicut teipsum ".
LUKE|10|28|Dixitque illi: " Recte respondisti; hoc fac et vives ".
LUKE|10|29|Ille autem, volens iustificare seipsum, dixit ad Iesum: " Et quis est meus proximus? ".
LUKE|10|30|Suscipiens autem Iesus dixit: " Homo quidam descendebat ab Ierusalem in Iericho et incidit in latrones, qui etiam despoliaverunt eum et, plagis impositis, abierunt, semivivo relicto.
LUKE|10|31|Accidit autem, ut sacerdos quidam descenderet eadem via et, viso illo, praeterivit;
LUKE|10|32|similiter et Levita, cum esset secus locum et videret eum, pertransiit.
LUKE|10|33|Samaritanus autem quidam iter faciens, venit secus eum et videns eum misericordia motus est,
LUKE|10|34|et appropians alligavit vulnera eius infundens oleum et vinum; et imponens illum in iumentum suum duxit in stabulum et curam eius egit.
LUKE|10|35|Et altera die protulit duos denarios et dedit stabulario et ait: "Curam illius habe, et, quodcumque supererogaveris, ego, cum rediero, reddam tibi".
LUKE|10|36|Quis horum trium videtur tibi proximus fuisse illi, qui incidit in latrones? ".
LUKE|10|37|At ille dixit: " Qui fecit misericordiam in illum ". Et ait illi Iesus: Vade et tu fac similiter ".
LUKE|10|38|Cum autem irent, ipse intravit in quoddam castellum, et mulier quaedam Martha nomine excepit illum.
LUKE|10|39|Et huic erat soror nomine Maria, quae etiam sedens secus pedes Domini audiebat verbum illius.
LUKE|10|40|Martha autem satagebat circa frequens ministerium; quae stetit et ait: Domine, non est tibi curae quod soror mea reliquit me solam ministrare? Dic ergo illi, ut me adiuvet ".
LUKE|10|41|Et respondens dixit illi Dominus: " Martha, Martha, sollicita es et turbaris erga plurima,
LUKE|10|42|porro unum est necessarium; Maria enim optimam partem elegit, quae non auferetur ab ea ".
LUKE|11|1|Et factum est cum esset in loco quodam orans, ut cessa vit, dixit unus ex discipulis eius ad eum: " Domine, doce nos orare, sicut et Ioannes docuit discipulos suos ".
LUKE|11|2|Et ait illis: " Cum oratis, dicite:Pater, sanctificetur nomen tuum,adveniat regnum tuum;
LUKE|11|3|panem nostrum cotidianum da nobis cotidie,
LUKE|11|4|et dimitte nobis peccata nostra,si quidem et ipsi dimittimus omni debenti nobis,et ne nos inducas in tentationem ".
LUKE|11|5|Et ait ad illos: " Quis vestrum habebit amicum et ibit ad illum media nocte et dicet illi: "Amice, commoda mihi tres panes,
LUKE|11|6|quoniam amicus meus venit de via ad me, et non habeo, quod ponam ante illum";
LUKE|11|7|et ille de intus respondens dicat: "Noli mihi molestus esse; iam ostium clausum est, et pueri mei mecum sunt in cubili; non possum surgere et dare tibi".
LUKE|11|8|Dico vobis: Et si non dabit illi surgens, eo quod amicus eius sit, propter improbitatem tamen eius surget et dabit illi, quotquot habet necessarios.
LUKE|11|9|Et ego vobis dico: Petite, et dabitur vobis; quaerite, et invenietis; pulsate, et aperietur vobis.
LUKE|11|10|Omnis enim qui petit, accipit; et, qui quaerit, invenit; et pulsanti aperietur.
LUKE|11|11|Quem autem ex vobis patrem filius petierit piscem, numquid pro pisce serpentem dabit illi?
LUKE|11|12|Aut si petierit ovum, numquid porriget illi scorpionem?
LUKE|11|13|Si ergo vos, cum sitis mali, nostis dona bona dare filiis vestris, quanto magis Pater de caelo dabit Spiritum Sanctum petentibus se ".
LUKE|11|14|Et erat eiciens daemonium, et illud erat mutum; et factum est, cum daemonium exisset, locutus est mutus. Et admiratae sunt turbae;
LUKE|11|15|quidam autem ex eis dixerunt: " In Beelzebul principe daemoniorum eicit daemonia ".
LUKE|11|16|Et alii tentantes signum de caelo quaerebant ab eo.
LUKE|11|17|Ipse autem sciens cogitationes eorum dixit eis: " Omne regnum in seipsum divisum desolatur, et domus supra domum cadit.
LUKE|11|18|Si autem et Satanas in seipsum divisus est, quomodo stabit regnum ipsius? Quia dicitis in Beelzebul eicere me daemonia.
LUKE|11|19|Si autem ego in Beelzebul eicio daemonia, filii vestri in quo eiciunt? Ideo ipsi iudices vestri erunt.
LUKE|11|20|Porro si in digito Dei eicio daemonia, profecto pervenit in vos regnum Dei.
LUKE|11|21|Cum fortis armatus custodit atrium suum, in pace sunt ea, quae possidet;
LUKE|11|22|si autem fortior illo superveniens vicerit eum, universa arma eius auferet, in quibus confidebat, et spolia eius distribuet.
LUKE|11|23|Qui non est mecum, adversum me est; et, qui non colligit mecum, dispergit.
LUKE|11|24|Cum immundus spiritus exierit de homine, perambulat per loca inaquosa quaerens requiem; et non inveniens dicit: "Revertar in domum meam unde exivi".
LUKE|11|25|Et cum venerit, invenit scopis mundatam et exornatam.
LUKE|11|26|Et tunc vadit et assumit septem alios spiritus nequiores se, et ingressi habitant ibi; et sunt novissima hominis illius peiora prioribus.
LUKE|11|27|Factum est autem, cum haec diceret, extollens vocem quaedam mulier de turba dixit illi: " Beatus venter, qui te portavit, et ubera, quae suxisti! ".
LUKE|11|28|At ille dixit: " Quinimmo beati, qui audiunt verbum Dei et custodiunt!.
LUKE|11|29|Turbis autem concurrentibus, coepit dicere: " Generatio haec generatio nequam est; signum quaerit, et signum non dabitur illi, nisi signum Ionae.
LUKE|11|30|Nam sicut Ionas fuit signum Ninevitis, ita erit et Filius hominis generationi isti.
LUKE|11|31|Regina austri surget in iudicio cum viris generationis huius et condemnabit illos, quia venit a finibus terrae audire sapientiam Salomonis, et ecce plus Salomone hic.
LUKE|11|32|Viri Ninevitae surgent in iudicio cum generatione hac et condemnabunt illam, quia paenitentiam egerunt ad praedicationem Ionae, et ecce plus Iona hic.
LUKE|11|33|Nemo lucernam accendit et in abscondito ponit neque sub modio sed supra candelabrum, ut, qui ingrediuntur, lumen videant.
LUKE|11|34|Lucerna corporis est oculus tuus. Si oculus tuus fuerit simplex, totum corpus tuum lucidum erit; si autem nequam fuerit, etiam corpus tuum tenebrosum erit.
LUKE|11|35|Vide ergo, ne lumen, quod in te est, tenebrae sint.
LUKE|11|36|Si ergo corpus tuum totum lucidum fuerit non habens aliquam partem tenebrarum, erit lucidum totum, sicut quando lucerna in fulgore suo illuminat te ".
LUKE|11|37|Et cum loqueretur, rogavit illum quidam pharisaeus, ut pranderet apud se; et ingressus recubuit.
LUKE|11|38|Pharisaeus autem videns miratus est quod non baptizatus esset ante prandium.
LUKE|11|39|Et ait Dominus ad illum: " Nunc vos pharisaei, quod de foris est calicis et catini, mundatis; quod autem intus est vestrum, plenum est rapina et iniquitate.
LUKE|11|40|Stulti! Nonne, qui fecit, quod de foris est, etiam id, quod de intus est, fecit?
LUKE|11|41|Verumtamen, quae insunt, date eleemosynam; et ecce omnia munda sunt vobis.
LUKE|11|42|Sed vae vobis pharisaeis, quia decimatis mentam et rutam et omne holus et praeteritis iudicium et caritatem Dei! Haec autem oportuit facere et illa non omittere.
LUKE|11|43|Vae vobis pharisaeis, quia diligitis primam cathedram in synagogis et salutationes in foro!
LUKE|11|44|Vae vobis, quia estis ut monumenta, quae non parent, et homines ambulantes supra nesciunt! ".
LUKE|11|45|Respondens autem quidam ex legis peritis ait illi: " Magister, haec dicens etiam nobis contumeliam facis ".
LUKE|11|46|At ille ait: " Et vobis legis peritis: Vae, quia oneratis homines oneribus, quae portari non possunt, et ipsi uno digito vestro non tangitis sarcinas!
LUKE|11|47|Vae vobis, quia aedificatis monumenta prophetarum, patres autem vestri occiderunt illos!
LUKE|11|48|Profecto testificamini et consentitis operibus patrum vestrorum, quoniam ipsi quidem eos occiderunt, vos autem aedificatis.
LUKE|11|49|Propterea et sapientia Dei dixit: Mittam ad illos prophetas et apostolos, et ex illis occident et persequentur,
LUKE|11|50|ut requiratur sanguis omnium prophetarum, qui effusus est a constitutione mundi, a generatione ista,
LUKE|11|51|a sanguine Abel usque ad sanguinem Zachariae, qui periit inter altare et aedem. Ita dico vobis: Requiretur ab hac generatione.
LUKE|11|52|Vae vobis legis peritis, quia tulistis clavem scientiae! Ipsi non introistis et eos, qui introibant, prohibuistis ".
LUKE|11|53|Cum autem inde exisset, coeperunt scribae et pharisaei graviter insistere et eum allicere in sermone de multis
LUKE|11|54|insidiantes ei, ut caperent aliquid ex ore eius.
LUKE|12|1|Interea multis turbis cir cumstantibus, ita ut se invi cem conculcarent, coepit dicere ad discipulos suos primum: " Attendite a fermento pharisaeorum, quod est hypocrisis.
LUKE|12|2|Nihil autem opertum est, quod non reveletur, neque absconditum, quod non sciatur.
LUKE|12|3|Quoniam, quae in tenebris dixistis, in lumine audientur; et, quod in aurem locuti estis in cubiculis, praedicabitur in tectis.
LUKE|12|4|Dico autem vobis amicis meis: Ne terreamini ab his, qui occidunt corpus et post haec non habent amplius, quod faciant.
LUKE|12|5|Ostendam autem vobis quem timeatis: Timete eum, qui postquam occiderit, habet potestatem mittere in gehennam. Ita dico vobis: Hunc timete.
LUKE|12|6|Nonne quinque passeres veneunt dipundio? Et unus ex illis non est in oblivione coram Deo.
LUKE|12|7|Sed et capilli capitis vestri omnes numerati sunt. Nolite timere; multis passeribus pluris estis.
LUKE|12|8|Dico autem vobis: Omnis, quicumque confessus fuerit in me coram hominibus, et Filius hominis confitebitur in illo coram angelis Dei;
LUKE|12|9|qui autem negaverit me coram hominibus, denegabitur coram angelis Dei.
LUKE|12|10|Et omnis, qui dicet verbum in Filium hominis, remittetur illi; ei autem, qui in Spiritum Sanctum blasphemaverit, non remittetur.
LUKE|12|11|Cum autem inducent vos in synagogas et ad magistratus et potestates, nolite solliciti esse qualiter aut quid respondeatis aut quid dicatis:
LUKE|12|12|Spiritus enim Sanctus docebit vos in ipsa hora, quae oporteat dicere ".
LUKE|12|13|Ait autem quidam ei de turba: " Magister, dic fratri meo, ut dividat mecum hereditatem ".
LUKE|12|14|At ille dixit ei: " Homo, quis me constituit iudicem aut divisorem super vos? ".
LUKE|12|15|Dixitque ad illos: " Videte et cavete ab omni avaritia, quia si cui res abundant, vita eius non est ex his, quae possidet ".
LUKE|12|16|Dixit autem similitudinem ad illos dicens: " Hominis cuiusdam divitis uberes fructus ager attulit.
LUKE|12|17|Et cogitabat intra se dicens: "Quid faciam, quod non habeo, quo congregem fructus meos?".
LUKE|12|18|Et dixit: "Hoc faciam: destruam horrea mea et maiora aedificabo et illuc congregabo omne triticum et bona mea;
LUKE|12|19|et dicam animae meae: Anima, habes multa bona posita in annos plurimos; requiesce, comede, bibe, epulare".
LUKE|12|20|Dixit autem illi Deus: "Stulte! Hac nocte animam tuam repetunt a te; quae autem parasti, cuius erunt?".
LUKE|12|21|Sic est qui sibi thesaurizat et non fit in Deum dives ".
LUKE|12|22|Dixitque ad discipulos suos: " Ideo dico vobis: nolite solliciti esse animae quid manducetis, neque corpori quid vestiamini.
LUKE|12|23|Anima enim plus est quam esca, et corpus quam vestimentum.
LUKE|12|24|Considerate corvos, quia non seminant neque metunt, quibus non est cellarium neque horreum, et Deus pascit illos; quanto magis vos pluris estis volucribus.
LUKE|12|25|Quis autem vestrum cogitando potest adicere ad aetatem suam cubitum?
LUKE|12|26|Si ergo neque, quod minimum est, potestis, quid de ceteris solliciti estis?
LUKE|12|27|Considerate lilia quomodo crescunt: non laborant neque nent; dico autem vobis: Nec Salomon in omni gloria sua vestiebatur sicut unum ex istis.
LUKE|12|28|Si autem fenum, quod hodie in agro est et cras in clibanum mittitur, Deus sic vestit, quanto magis vos, pusillae fidei.
LUKE|12|29|Et vos nolite quaerere quid manducetis aut quid bibatis et nolite solliciti esse.
LUKE|12|30|Haec enim omnia gentes mundi quaerunt; Pater autem vester scit quoniam his indigetis.
LUKE|12|31|Verumtamen quaerite regnum eius; et haec adicientur vobis.
LUKE|12|32|Noli timere, pusillus grex, quia complacuit Patri vestro dare vobis regnum.
LUKE|12|33|Vendite, quae possidetis, et date eleemosynam. Facite vobis sacculos, qui non veterescunt, thesaurum non deficientem in caelis, quo fur non appropiat, neque tinea corrumpit;
LUKE|12|34|ubi enim thesaurus vester est, ibi et cor vestrum erit.
LUKE|12|35|Sint lumbi vestri praecincti et lucernae ardentes,
LUKE|12|36|et vos similes hominibus exspectantibus dominum suum, quando revertatur a nuptiis, ut, cum venerit et pulsaverit, confestim aperiant ei.
LUKE|12|37|Beati, servi illi, quos, cum venerit dominus, invenerit vigilantes. Amen dico vobis, quod praecinget se et faciet illos discumbere et transiens ministrabit illis.
LUKE|12|38|Et si venerit in secunda vigilia, et si in tertia vigilia venerit, et ita invenerit, beati sunt illi.
LUKE|12|39|Hoc autem scitote, quia, si sciret pater familias, qua hora fur veniret, non sineret perfodi domum suam.
LUKE|12|40|Et vos estote parati, quia, qua hora non putatis, Filius hominis venit.
LUKE|12|41|Ait autem Petrus: " Domine, ad nos dicis hanc parabolam an et ad omnes?.
LUKE|12|42|Et dixit Dominus: " Quis putas est fidelis dispensator et prudens, quem constituet dominus super familiam suam, ut det illis in tempore tritici mensuram?
LUKE|12|43|Beatus ille servus, quem, cum venerit dominus eius, invenerit ita facientem.
LUKE|12|44|Vere dico vobis: Supra omnia, quae possidet, constituet illum.
LUKE|12|45|Quod si dixerit servus ille in corde suo: "Moram facit dominus meus venire", et coeperit percutere pueros et ancillas et edere et bibere et inebriari,
LUKE|12|46|veniet dominus servi illius in die, qua non sperat, et hora, qua nescit, et dividet eum partemque eius cum infidelibus ponet.
LUKE|12|47|Ille autem servus, qui cognovit voluntatem domini sui et non praeparavit vel non fecit secundum voluntatem eius, vapulabit multis;
LUKE|12|48|qui autem non cognovit et fecit digna plagis, vapulabit paucis. Omni autem, cui multum datum est, multum quaeretur ab eo; et cui commendaverunt multum, plus petent ab eo.
LUKE|12|49|Ignem veni mittere in terram et quid volo? Si iam accensus esset!
LUKE|12|50|Baptisma autem habeo baptizari et quomodo coartor, usque dum perficiatur!
LUKE|12|51|Putatis quia pacem veni dare in terram? Non, dico vobis, sed separationem.
LUKE|12|52|Erunt enim ex hoc quinque in domo una divisi: tres in duo, et duo in tres;
LUKE|12|53|dividentur pater in filium et filius in patrem, mater in filiam et filia in matrem, socrus in nurum suam et nurus in socrum ".
LUKE|12|54|Dicebat autem et ad turbas: " Cum videritis nubem orientem ab occasu, statim dicitis: "Nimbus venit", et ita fit;
LUKE|12|55|et cum austrum flantem, dicitis: "Aestus erit", et fit.
LUKE|12|56|Hypocritae, faciem terrae et caeli nostis probare, hoc autem tempus quomodo nescitis probare?
LUKE|12|57|Quid autem et a vobis ipsis non iudicatis, quod iustum est?
LUKE|12|58|Cum autem vadis cum adversario tuo ad principem, in via da operam liberari ab illo, ne forte trahat te apud iudicem, et iudex tradat te exactori, et exactor mittat te in carcerem.
LUKE|12|59|Dico tibi: Non exies inde, donec etiam novissimum minutum reddas ".
LUKE|13|1|Aderant autem quidam ipso in tempore nuntiantes illi de Galilaeis, quorum sanguinem Pilatus miscuit cum sacrificiis eorum.
LUKE|13|2|Et respondens dixit illis: " Putatis quod hi Galilaei prae omnibus Galilaeis peccatores fuerunt, quia talia passi sunt?
LUKE|13|3|Non, dico vobis, sed, nisi paenitentiam egeritis, omnes similiter peribitis.
LUKE|13|4|Vel illi decem et octo, supra quos cecidit turris in Siloam et occidit eos, putatis quia et ipsi debitores fuerunt praeter omnes homines habitantes in Ierusalem?
LUKE|13|5|Non, dico vobis, sed, si non paenitentiam egeritis, omnes similiter peribitis ".
LUKE|13|6|Dicebat autem hanc similitudinem: " Arborem fici habebat quidam plantatam in vinea sua et venit quaerens fructum in illa et non invenit.
LUKE|13|7|Dixit autem ad cultorem vineae: "Ecce anni tres sunt, ex quo venio quaerens fructum in ficulnea hac et non invenio. Succide ergo illam. Ut quid etiam terram evacuat?".
LUKE|13|8|At ille respondens dicit illi: "Domine, dimitte illam et hoc anno, usque dum fodiam circa illam et mittam stercora,
LUKE|13|9|et si quidem fecerit fructum in futurum; sin autem succides eam" ".
LUKE|13|10|Erat autem docens in una synagogarum sabbatis.
LUKE|13|11|Et ecce mulier, quae habebat spiritum infirmitatis annis decem et octo et erat inclinata nec omnino poterat sursum respicere.
LUKE|13|12|Quam cum vidisset Iesus, vocavit et ait illi: " Mulier, dimissa es ab infirmitate tua ",
LUKE|13|13|et imposuit illi manus; et confestim erecta est et glorificabat Deum.
LUKE|13|14|Respondens autem archisynagogus, indignans quia sabbato curasset Iesus, dicebat turbae: " Sex dies sunt, in quibus oportet operari; in his ergo venite et curamini et non in die sabbati ".
LUKE|13|15|Respondit autem ad illum Dominus et dixit: " Hypocritae, unusquisque vestrum sabbato non solvit bovem suum aut asinum a praesepio et ducit adaquare?
LUKE|13|16|Hanc autem filiam Abrahae, quam alligavit Satanas ecce decem et octo annis, non oportuit solvi a vinculo isto die sabbati? ".
LUKE|13|17|Et cum haec diceret, erubescebant omnes adversarii eius, et omnis populus gaudebat in universis, quae gloriose fiebant ab eo.
LUKE|13|18|Dicebat ergo: " Cui simile est regnum Dei, et cui simile existimabo illud?
LUKE|13|19|Simile est grano sinapis, quod acceptum homo misit in hortum suum, et crevit et factum est in arborem, et volucres caeli requieverunt in ramis eius ".
LUKE|13|20|Et iterum dixit: " Cui simile aestimabo regnum Dei?
LUKE|13|21|Simile est fermento, quod acceptum mulier abscondit in farinae sata tria, donec fermentaretur totum ".
LUKE|13|22|Et ibat per civitates et castella docens et iter faciens in Hierosolymam.
LUKE|13|23|Ait autem illi quidam: " Domine, pauci sunt, qui salvantur? ". Ipse autem dixit ad illos:
LUKE|13|24|" Contendite intrare per angustam portam, quia multi, dico vobis, quaerent intrare et non poterunt.
LUKE|13|25|Cum autem surrexerit pater familias et clauserit ostium, et incipietis foris stare et pulsare ostium dicentes: "Domine, aperi nobis"; et respondens dicet vobis: "Nescio vos unde sitis".
LUKE|13|26|Tunc incipietis dicere: "Manducavimus coram te et bibimus, et in plateis nostris docuisti";
LUKE|13|27|et dicet loquens vobis: "Nescio vos unde sitis; discedite a me, omnes operarii iniquitatis".
LUKE|13|28|Ibi erit fletus et stridor dentium, cum videritis Abraham et Isaac et Iacob et omnes prophetas in regno Dei, vos autem expelli foras.
LUKE|13|29|Et venient ab oriente et occidente et aquilone et austro et accumbent in regno Dei.
LUKE|13|30|Et ecce sunt novissimi, qui erunt primi, et sunt primi, qui erunt novissimi ".
LUKE|13|31|In ipsa hora accesserunt quidam pharisaeorum dicentes illi: " Exi et vade hinc, quia Herodes vult te occidere ".
LUKE|13|32|Et ait illis: " Ite, dicite vulpi illi: "Ecce eicio daemonia et sanitates perficio hodie et cras et tertia consummor.
LUKE|13|33|Verumtamen oportet me hodie et cras et sequenti ambulare, quia non capit prophetam perire extra Ierusalem".
LUKE|13|34|Ierusalem, Ierusalem, quae occidis prophetas et lapidas eos, qui missi sunt ad te, quotiens volui congregare filios tuos, quemadmodum avis nidum suum sub pinnis, et noluistis.
LUKE|13|35|Ecce relinquitur vobis domus vestra. Dico autem vobis: Non videbitis me, donec veniat cum dicetis: "Benedictus, qui venit in nomine Domini" ".
LUKE|14|1|Et factum est, cum intraret in domum cuiusdam princi pis pharisaeorum sabbato manducare panem, et ipsi observabant eum.
LUKE|14|2|Et ecce homo quidam hydropicus erat ante illum.
LUKE|14|3|Et respondens Iesus dixit ad legis peritos et pharisaeos dicens: " Licet sabbato curare an non? ".
LUKE|14|4|At illi tacuerunt. Ipse vero apprehensum sanavit eum ac dimisit.
LUKE|14|5|Et ad illos dixit: " Cuius vestrum filius aut bos in puteum cadet, et non continuo extrahet illum die sabbati? ".
LUKE|14|6|Et non poterant ad haec respondere illi.
LUKE|14|7|Dicebat autem ad invitatos parabolam, intendens quomodo primos accubitus eligerent, dicens ad illos:
LUKE|14|8|" Cum invitatus fueris ab aliquo ad nuptias, non discumbas in primo loco, ne forte honoratior te sit invitatus ab eo,
LUKE|14|9|et veniens is qui te et illum vocavit, dicat tibi: "Da huic locum"; et tunc incipias cum rubore novissimum locum tenere.
LUKE|14|10|Sed cum vocatus fueris, vade, recumbe in novissimo loco, ut, cum venerit qui te invitavit, dicat tibi: "Amice, ascende superius"; tunc erit tibi gloria coram omnibus simul discumbentibus.
LUKE|14|11|Quia omnis, qui se exaltat, humiliabitur; et, qui se humiliat, exaltabitur ".
LUKE|14|12|Dicebat autem et ei, qui se invitaverat: " Cum facis prandium aut cenam, noli vocare amicos tuos neque fratres tuos neque cognatos neque vicinos divites, ne forte et ipsi te reinvitent, et fiat tibi retributio.
LUKE|14|13|Sed cum facis convivium, voca pauperes, debiles, claudos, caecos;
LUKE|14|14|et beatus eris, quia non habent retribuere tibi. Retribuetur enim tibi in resurrectione iustorum ".
LUKE|14|15|Haec cum audisset quidam de simul discumbentibus, dixit illi: " Beatus, qui manducabit panem in regno Dei ".
LUKE|14|16|At ipse dixit ei: " Homo quidam fecit cenam magnam et vocavit multos;
LUKE|14|17|et misit servum suum hora cenae dicere invitatis: "Venite, quia iam paratum est".
LUKE|14|18|Et coeperunt simul omnes excusare. Primus dixit ei: "Villam emi et necesse habeo exire et videre illam; rogo te, habe me excusatum".
LUKE|14|19|Et alter dixit: "Iuga boum emi quinque et eo probare illa; rogo te, habe me excusatum".
LUKE|14|20|Et alius dixit: "Uxorem duxi et ideo non possum venire".
LUKE|14|21|Et reversus servus nuntiavit haec domino suo. Tunc iratus pater familias dixit servo suo: "Exi cito in plateas et vicos civitatis et pauperes ac debiles et caecos et claudos introduc huc".
LUKE|14|22|Et ait servus: "Domine, factum est, ut imperasti, et adhuc locus est".
LUKE|14|23|Et ait dominus servo: "Exi in vias et saepes, et compelle intrare, ut impleatur domus mea.
LUKE|14|24|Dico autem vobis, quod nemo virorum illorum, qui vocati sunt, gustabit cenam meam" ".
LUKE|14|25|Ibant autem turbae multae cum eo; et conversus dixit ad illos:
LUKE|14|26|" Si quis venit ad me et non odit patrem suum et matrem et uxorem et filios et fratres et sorores, adhuc et animam suam, non potest esse meus discipulus.
LUKE|14|27|Et, qui non baiulat crucem suam et venit post me, non potest esse meus discipulus.
LUKE|14|28|Quis enim ex vobis volens turrem aedificare, non prius sedens computat sumptus, si habet ad perficiendum?
LUKE|14|29|Ne, posteaquam posuerit fundamentum et non potuerit perficere, omnes, qui vident, incipiant illudere ei
LUKE|14|30|dicentes: "Hic homo coepit aedificare et non potuit consummare".
LUKE|14|31|Aut quis rex, iturus committere bellum adversus alium regem, non sedens prius cogitat, si possit cum decem milibus occurrere ei, qui cum viginti milibus venit ad se?
LUKE|14|32|Alioquin, adhuc illo longe agente, legationem mittens rogat ea, quae pacis sunt.
LUKE|14|33|Sic ergo omnis ex vobis, qui non renuntiat omnibus, quae possidet, non potest meus esse discipulus.
LUKE|14|34|Bonum est sal; si autem sal quoque evanuerit, in quo condietur?
LUKE|14|35|Neque in terram neque in sterquilinium utile est, sed foras proiciunt illud. Qui habet aures audiendi, audiat ".
LUKE|15|1|Erant autem appropinquan tes ei omnes publicani et pec catores, ut audirent illum.
LUKE|15|2|Et murmurabant pharisaei et scribae dicentes: " Hic peccatores recipit et manducat cum illis ".
LUKE|15|3|Et ait ad illos parabolam istam dicens:
LUKE|15|4|" Quis ex vobis homo, qui habet centum oves et si perdiderit unam ex illis, nonne dimittit nonaginta novem in deserto et vadit ad illam, quae perierat, donec inveniat illam?
LUKE|15|5|Et cum invenerit eam, imponit in umeros suos gaudens
LUKE|15|6|et veniens domum convocat amicos et vicinos dicens illis: Congratulamini mihi, quia inveni ovem meam, quae perierat".
LUKE|15|7|Dico vobis: Ita gaudium erit in caelo super uno peccatore paenitentiam agente quam super nonaginta novem iustis, qui non indigent paenitentia.
LUKE|15|8|Aut quae mulier habens drachmas decem, si perdiderit drachmam unam, nonne accendit lucernam et everrit domum et quaerit diligenter, donec inveniat?
LUKE|15|9|Et cum invenerit, convocat amicas et vicinas dicens: "Congratulamini mihi, quia inveni drachmam, quam perdideram".
LUKE|15|10|Ita dico vobis: Gaudium fit coram angelis Dei super uno peccatore paenitentiam agente ".
LUKE|15|11|Ait autem: " Homo quidam habebat duos filios.
LUKE|15|12|Et dixit adulescentior ex illis patri: "Pater, da mihi portionem substantiae, quae me contingit". Et divisit illis substantiam.
LUKE|15|13|Et non post multos dies, congregatis omnibus, adulescentior filius peregre profectus est in regionem longinquam et ibi dissipavit substantiam suam vivendo luxuriose.
LUKE|15|14|Et postquam omnia consummasset, facta est fames valida in regione illa, et ipse coepit egere.
LUKE|15|15|Et abiit et adhaesit uni civium regionis illius, et misit illum in villam suam, ut pasceret porcos;
LUKE|15|16|et cupiebat saturari de siliquis, quas porci manducabant, et nemo illi dabat.
LUKE|15|17|In se autem reversus dixit: "Quanti mercennarii patris mei abundant panibus, ego autem hic fame pereo.
LUKE|15|18|Surgam et ibo ad patrem meum et dicam illi: Pater, peccavi in caelum et coram te
LUKE|15|19|et iam non sum dignus vocari filius tuus; fac me sicut unum de mercennariis tuis".
LUKE|15|20|Et surgens venit ad patrem suum.Cum autem adhuc longe esset, vidit illum pater ipsius et misericordia motus est et accurrens cecidit supra collum eius et osculatus est illum.
LUKE|15|21|Dixitque ei filius: "Pater, peccavi in caelum et coram te; iam non sum dignus vocari filius tuus".
LUKE|15|22|Dixit autem pater ad servos suos: "Cito proferte stolam primam et induite illum et date anulum in manum eius et calceamenta in pedes
LUKE|15|23|et adducite vitulum saginatum, occidite et manducemus et epulemur,
LUKE|15|24|quia hic filius meus mortuus erat et revixit, perierat et inventus est". Et coeperunt epulari.
LUKE|15|25|Erat autem filius eius senior in agro et, cum veniret et appropinquaret domui, audivit symphoniam et choros
LUKE|15|26|et vocavit unum de servis et interrogavit quae haec essent.
LUKE|15|27|Isque dixit illi: "Frater tuus venit, et occidit pater tuus vitulum saginatum, quia salvum illum recepit".
LUKE|15|28|Indignatus est autem et nolebat introire. Pater ergo illius egressus coepit rogare illum.
LUKE|15|29|At ille respondens dixit patri suo: "Ecce tot annis servio tibi et numquam mandatum tuum praeterii, et numquam dedisti mihi haedum, ut cum amicis meis epularer;
LUKE|15|30|sed postquam filius tuus hic, qui devoravit substantiam tuam cum meretricibus, venit, occidisti illi vitulum saginatum".
LUKE|15|31|At ipse dixit illi: "Fili, tu semper mecum es, et omnia mea tua sunt;
LUKE|15|32|epulari autem et gaudere oportebat, quia frater tuus hic mortuus erat et revixit, perierat et inventus est" ".
LUKE|16|1|Dicebat autem et ad disci pulos: " Homo quidam erat dives, qui habebat vilicum, et hic diffamatus est apud illum quasi dissipasset bona ipsius.
LUKE|16|2|Et vocavit illum et ait illi: "Quid hoc audio de te? Redde rationem vilicationis tuae; iam enim non poteris vilicare".
LUKE|16|3|Ait autem vilicus intra se: "Quid faciam, quia dominus meus aufert a me vilicationem? Fodere non valeo, mendicare erubesco.
LUKE|16|4|Scio quid faciam, ut, cum amotus fuero a vilicatione, recipiant me in domos suas".
LUKE|16|5|Convocatis itaque singulis debitoribus domini sui, dicebat primo: Quantum debes domino meo?".
LUKE|16|6|At ille dixit: "Centum cados olei". Dixitque illi: "Accipe cautionem tuam et sede cito, scribe quinquaginta".
LUKE|16|7|Deinde alii dixit: "Tu vero quantum debes?". Qui ait: "Centum coros tritici". Ait illi: "Accipe litteras tuas et scribe octoginta".
LUKE|16|8|Et laudavit dominus vilicum iniquitatis, quia prudenter fecisset, quia filii huius saeculi prudentiores filiis lucis in generatione sua sunt.
LUKE|16|9|Et ego vobis dico: Facite vobis amicos de mammona iniquitatis, ut, cum defecerit, recipiant vos in aeterna tabernacula.
LUKE|16|10|Qui fidelis est in minimo, et in maiori fidelis est; et, qui in modico iniquus est, et in maiori iniquus est.
LUKE|16|11|Si ergo in iniquo mammona fideles non fuistis, quod verum est, quis credet vobis?
LUKE|16|12|Et si in alieno fideles non fuistis, quod vestrum est, quis dabit vobis?
LUKE|16|13|Nemo servus potest duobus dominis servire: aut enim unum odiet et alterum diliget, aut uni adhaerebit et alterum contemnet. Non potestis Deo servire et mammonae ".
LUKE|16|14|Audiebant autem omnia haec pharisaei, qui erant avari, et deridebant illum.
LUKE|16|15|Et ait illis: " Vos estis, qui iustificatis vos coram hominibus; Deus autem novit corda vestra, quia, quod hominibus altum est, abominatio est ante Deum.
LUKE|16|16|Lex et Prophetae usque ad Ioannem; ex tunc regnum Dei evangelizatur, et omnis in illud vim facit.
LUKE|16|17|Facilius est autem caelum et terram praeterire, quam de Lege unum apicem cadere.
LUKE|16|18|Omnis, qui dimittit uxorem suam et ducit alteram, moechatur; et, qui dimissam a viro ducit, moechatur.
LUKE|16|19|Homo quidam erat dives et induebatur purpura et bysso et epulabatur cotidie splendide.
LUKE|16|20|Quidam autem pauper nomine Lazarus iacebat ad ianuam eius ulceribus plenus
LUKE|16|21|et cupiens saturari de his, quae cadebant de mensa divitis; sed et canes veniebant et lingebant ulcera eius.
LUKE|16|22|Factum est autem ut moreretur pauper et portaretur ab angelis in sinum Abrahae; mortuus est autem et dives et sepultus est.
LUKE|16|23|Et in inferno elevans oculos suos, cum esset in tormentis, videbat Abraham a longe et Lazarum in sinu eius.
LUKE|16|24|Et ipse clamans dixit: "Pater Abraham, miserere mei et mitte Lazarum, ut intingat extremum digiti sui in aquam, ut refrigeret linguam meam, quia crucior in hac flamma".
LUKE|16|25|At dixit Abraham: "Fili, recordare quia recepisti bona tua in vita tua, et Lazarus similiter mala; nunc autem hic consolatur, tu vero cruciaris.
LUKE|16|26|Et in his omnibus inter nos et vos chaos magnum firmatum est, ut hi, qui volunt hinc transire ad vos, non possint, neque inde ad nos transmeare".
LUKE|16|27|Et ait: "Rogo ergo te, Pater, ut mittas eum in domum patris mei
LUKE|16|28|- habeo enim quinque fratres - ut testetur illis, ne et ipsi veniant in locum hunc tormentorum".
LUKE|16|29|Ait autem Abraham: "Habent Moysen et Prophetas; audiant illos".
LUKE|16|30|At ille dixit: "Non, pater Abraham, sed si quis ex mortuis ierit ad eos, paenitentiam agent".
LUKE|16|31|Ait autem illi: "Si Moysen et Prophetas non audiunt, neque si quis ex mortuis resurrexerit, credent" ".
LUKE|17|1|Et ad discipulos suos ait: " Impossibile est ut non ve niant scandala; vae autem illi, per quem veniunt!
LUKE|17|2|Utilius est illi, si lapis molaris imponatur circa collum eius et proiciatur in mare, quam ut scandalizet unum de pusillis istis.
LUKE|17|3|Attendite vobis!Si peccaverit frater tuus, increpa illum et, si paenitentiam egerit, dimitte illi;
LUKE|17|4|et si septies in die peccaverit in te et septies conversus fuerit ad te dicens: "Paenitet me", dimittes illi ".
LUKE|17|5|Et dixerunt apostoli Domino: " Adauge nobis fidem! ".
LUKE|17|6|Dixit autem Dominus: " Si haberetis fidem sicut granum sinapis, diceretis huic arbori moro: "Eradicare et transplantare in mare", et oboediret vobis.
LUKE|17|7|Quis autem vestrum habens servum arantem aut pascentem, qui regresso de agro dicet illi: "Statim transi, recumbe",
LUKE|17|8|et non dicet ei: "Para, quod cenem, et praecinge te et ministra mihi, donec manducem et bibam, et post haec tu manducabis et bibes"?
LUKE|17|9|Numquid gratiam habet servo illi, quia fecit, quae praecepta sunt?
LUKE|17|10|Sic et vos, cum feceritis omnia, quae praecepta sunt vobis, dicite: Servi inutiles sumus; quod debuimus facere, fecimus" ".
LUKE|17|11|Et factum est, dum iret in Ierusalem, et ipse transibat per mediam Samariam et Galilaeam.
LUKE|17|12|Et cum ingrederetur quoddam castellum, occurrerunt ei decem viri leprosi, qui steterunt a longe
LUKE|17|13|et levaverunt vocem dicentes: " Iesu praeceptor, miserere nostri! ".
LUKE|17|14|Quos ut vidit, dixit: " Ite, ostendite vos sacerdotibus ". Et factum est, dum irent, mundati sunt.
LUKE|17|15|Unus autem ex illis, ut vidit quia sanatus est, regressus est cum magna voce magnificans Deum
LUKE|17|16|et cecidit in faciem ante pedes eius gratias agens ei; et hic erat Samaritanus.
LUKE|17|17|Respondens autem Iesus dixit: " Nonne decem mundati sunt? Et novem ubi sunt?
LUKE|17|18|Non sunt inventi qui redirent, ut darent gloriam Deo, nisi hic alienigena? ".
LUKE|17|19|Et ait illi: " Surge, vade; fides tua te salvum fecit ".
LUKE|17|20|Interrogatus autem a pharisaeis: " Quando venit regnum Dei? ", respondit eis et dixit: " Non venit regnum Dei cum observatione,
LUKE|17|21|neque dicent: "Ecce hic" aut: "Illic"; ecce enim regnum Dei intra vos est ".
LUKE|17|22|Et ait ad discipulos: " Venient dies, quando desideretis videre unum diem Filii hominis et non videbitis.
LUKE|17|23|Et dicent vobis: "Ecce hic", "Ecce illic"; nolite ire neque sectemini.
LUKE|17|24|Nam sicut fulgur coruscans de sub caelo in ea, quae sub caelo sunt, fulget, ita erit Filius hominis in die sua.
LUKE|17|25|Primum autem oportet illum multa pati et reprobari a generatione hac.
LUKE|17|26|Et sicut factum est in diebus Noe, ita erit et in diebus Filii hominis:
LUKE|17|27|edebant, bibebant, uxores ducebant, dabantur ad nuptias, usque in diem, qua intravit Noe in arcam, et venit diluvium et perdidit omnes.
LUKE|17|28|Similiter sicut factum est in diebus Lot: edebant, bibebant, emebant, vendebant, plantabant, aedificabant;
LUKE|17|29|qua die autem exiit Lot a Sodomis, pluit ignem et sulphur de caelo et omnes perdidit.
LUKE|17|30|Secundum haec erit, qua die Filius hominis revelabitur.
LUKE|17|31|In illa die, qui fuerit in tecto, et vasa eius in domo, ne descendat tollere illa; et, qui in agro, similiter non redeat retro.
LUKE|17|32|Memores estote uxoris Lot.
LUKE|17|33|Quicumque quaesierit animam suam salvam facere, perdet illam; et, quicumque perdiderit illam, vivificabit eam.
LUKE|17|34|Dico vobis: Illa nocte erunt duo in lecto uno:unus assumetur, et alter relinquetur;
LUKE|17|35|duae erunt molentes in unum: una assumetur, et altera relinquetur ". 36) 37 Respondentes dicunt illi: " Ubi, Domine? ". Qui dixit eis: " Ubicumque fuerit corpus, illuc congregabuntur et aquilae ".
LUKE|18|1|Dicebat autem parabolam ad illos, quoniam oportet semper orare et non deficere,
LUKE|18|2|dicens: " Iudex quidam erat in quadam civitate, qui Deum non timebat et hominem non reverebatur.
LUKE|18|3|Vidua autem erat in civitate illa et veniebat ad eum dicens: "Vindica me de adversario meo".
LUKE|18|4|Et nolebat per multum tempus; post haec autem dixit intra se: "Etsi Deum non timeo nec hominem revereor,
LUKE|18|5|tamen quia molesta est mihi haec vidua, vindicabo illam, ne in novissimo veniens suggillet me" ".
LUKE|18|6|Ait autem Dominus: " Audite quid iudex iniquitatis dicit;
LUKE|18|7|Deus autem non faciet vindictam electorum suorum clamantium ad se die ac nocte, et patientiam habebit in illis?
LUKE|18|8|Dico vobis: Cito faciet vindictam illorum. Verumtamen Filius hominis veniens, putas, inveniet fidem in terra? ".
LUKE|18|9|Dixit autem et ad quosdam, qui in se confidebant tamquam iusti et aspernabantur ceteros, parabolam istam:
LUKE|18|10|" Duo homines ascenderunt in templum, ut orarent: unus pharisaeus et alter publicanus.
LUKE|18|11|Pharisaeus stans haec apud se orabat: "Deus, gratias ago tibi, quia non sum sicut ceteri hominum, raptores, iniusti, adulteri, velut etiam hic publicanus;
LUKE|18|12|ieiuno bis in sabbato, decimas do omnium, quae possideo".
LUKE|18|13|Et publicanus a longe stans nolebat nec oculos ad caelum levare, sed percutiebat pectus suum dicens: "Deus, propitius esto mihi peccatori".
LUKE|18|14|Dico vobis: Descendit hic iustificatus in domum suam ab illo. Quia omnis, qui se exaltat, humiliabitur; et, qui se humiliat, exaltabitur ".
LUKE|18|15|Afferebant autem ad illum et infantes, ut eos tangeret; quod cum viderent, discipuli increpabant illos.
LUKE|18|16|Iesus autem convocans illos dixit: " Sinite pueros venire ad me et nolite eos vetare; talium est enim regnum Dei.
LUKE|18|17|Amen dico vobis: Quicumque non acceperit regnum Dei sicut puer, non intrabit in illud ".
LUKE|18|18|Et interrogavit eum quidam princeps dicens: " Magister bone, quid faciens vitam aeternam possidebo? ".
LUKE|18|19|Dixit autem ei Iesus: " Quid me dicis bonum? Nemo bonus nisi solus Deus.
LUKE|18|20|Mandata nosti: non moechaberis, non occides, non furtum facies, non falsum testimonium dices, honora patrem tuum et matrem ".
LUKE|18|21|Qui ait: " Haec omnia custodivi a iuventute ".
LUKE|18|22|Quo audito, Iesus ait ei: " Adhuc unum tibi deest: omnia, quaecumque habes, vende et da pauperibus et habebis thesaurum in caelo: et veni, sequere me ".
LUKE|18|23|His ille auditis, contristatus est, quia dives erat valde.
LUKE|18|24|Videns autem illum Iesus tristem factum dixit: " Quam difficile, qui pecunias habent, in regnum Dei intrant.
LUKE|18|25|Facilius est enim camelum per foramen acus transire, quam divitem intrare in regnum Dei ".
LUKE|18|26|Et dixerunt, qui audiebant: " Et quis potest salvus fieri? ".
LUKE|18|27|Ait autem illis: " Quae impossibilia sunt apud homi nes, possibilia sunt apud Deum ".
LUKE|18|28|Ait autem Petrus: " Ecce nos dimisimus nostra et secuti sumus te ".
LUKE|18|29|Qui dixit eis: " Amen dico vobis: Nemo est, qui reliquit domum aut uxorem aut fratres aut parentes aut filios propter regnum Dei,
LUKE|18|30|et non recipiat multo plura in hoc tempore et in saeculo venturo vitam aeternam ".
LUKE|18|31|Assumpsit autem Duodecim et ait illis: " Ecce ascendimus Ierusalem, et consummabuntur omnia, quae scripta sunt per Prophetas de Filio hominis:
LUKE|18|32|tradetur enim gentibus et illudetur et contumeliis afficietur et conspuetur;
LUKE|18|33|et, postquam flagellaverint, occident eum, et die tertia resurget ".
LUKE|18|34|Et ipsi nihil horum intellexerunt; et erat verbum istud absconditum ab eis, et non intellegebant, quae dicebantur.
LUKE|18|35|Factum est autem, cum appropinquaret Iericho, caecus quidam sedebat secus viam mendicans.
LUKE|18|36|Et cum audiret turbam praetereuntem, interrogabat quid hoc esset.
LUKE|18|37|Dixerunt autem ei: " Iesus Nazarenus transit ".
LUKE|18|38|Et clamavit dicens: " Iesu, fili David, miserere mei! ".
LUKE|18|39|Et qui praeibant, increpabant eum, ut taceret; ipse vero multo magis clamabat: " Fili David, miserere mei! ".
LUKE|18|40|Stans autem Iesus iussit illum adduci ad se. Et cum appropinquasset, interrogavit illum:
LUKE|18|41|" Quid tibi vis faciam? ". At ille dixit: " Domine, ut videam ".
LUKE|18|42|Et Iesus dixit illi: " Respice! Fides tua te salvum fecit ". 43 Et confestim vidit et sequebatur illum magnificans Deum. Et omnis plebs, ut vidit, dedit laudem Deo.
LUKE|19|1|Et ingressus perambulabat Iericho.
LUKE|19|2|Et ecce vir nomine Zacchaeus, et hic erat princeps publicanorum et ipse dives.
LUKE|19|3|Et quaerebat videre Iesum, quis esset, et non poterat prae turba, quia statura pusillus erat.
LUKE|19|4|Et praecurrens ascendit in arborem sycomorum, ut videret illum, quia inde erat transiturus.
LUKE|19|5|Et cum venisset ad locum, suspiciens Iesus dixit ad eum: " Zacchaee, festinans descende, nam hodie in domo tua oportet me manere ".
LUKE|19|6|Et festinans descendit et excepit illum gaudens.
LUKE|19|7|Et cum viderent, omnes murmurabant dicentes: " Ad hominem peccatorem divertit! ".
LUKE|19|8|Stans autem Zacchaeus dixit ad Dominum: " Ecce dimidium bonorum meorum, Domine, do pauperibus et, si quid aliquem defraudavi, reddo quadruplum ".
LUKE|19|9|Ait autem Iesus ad eum: " Hodie salus domui huic facta est, eo quod et ipse filius sit Abrahae;
LUKE|19|10|venit enim Filius hominis quaerere et salvum facere, quod perierat ".
LUKE|19|11|Haec autem illis audientibus, adiciens dixit parabolam, eo quod esset prope Ierusalem, et illi existimarent quod confestim regnum Dei manifestaretur.
LUKE|19|12|Dixit ergo: " Homo quidam nobilis abiit in regionem longinquam accipere sibi regnum et reverti.
LUKE|19|13|Vocatis autem decem servis suis, dedit illis decem minas et ait ad illos: "Negotiamini, dum venio".
LUKE|19|14|Cives autem eius oderant illum et miserunt legationem post illum dicentes: "Nolumus hunc regnare super nos!".
LUKE|19|15|Et factum est ut rediret, accepto regno, et iussit ad se vocari servos illos, quibus dedit pecuniam, ut sciret quantum negotiati essent.
LUKE|19|16|Venit autem primus dicens: "Domine, mina tua decem minas acquisivit".
LUKE|19|17|Et ait illi: "Euge, bone serve; quia in modico fidelis fuisti, esto potestatem habens supra decem civitates".
LUKE|19|18|Et alter venit dicens: "Mina tua, domine, fecit quinque minas".
LUKE|19|19|Et huic ait: "Et tu esto supra quinque civitates".
LUKE|19|20|Et alter venit dicens: "Domine, ecce mina tua, quam habui repositam in sudario;
LUKE|19|21|timui enim te, quia homo austerus es: tollis, quod non posuisti, et metis, quod non seminasti".
LUKE|19|22|Dicit ei: "De ore tuo te iudico, serve nequam! Sciebas quod ego austerus homo sum, tollens quod non posui et metens quod non seminavi?
LUKE|19|23|Et quare non dedisti pecuniam meam ad mensam? Et ego veniens cum usuris utique exegissem illud".
LUKE|19|24|Et adstantibus dixit: "Auferte ab illo minam et date illi, qui decem minas habet".
LUKE|19|25|Et dixerunt ei: "Domine, habet decem minas!".
LUKE|19|26|Dico vobis: "Omni habenti dabitur; ab eo autem, qui non habet, et, quod habet, auferetur.
LUKE|19|27|Verumtamen inimicos meos illos, qui noluerunt me regnare super se, adducite huc et interficite ante me! ".
LUKE|19|28|Et his dictis, praecedebat ascendens Hierosolymam.
LUKE|19|29|Et factum est, cum appropinquasset ad Bethfage et Bethaniam, ad montem, qui vocatur Oliveti, misit duos discipulos
LUKE|19|30|dicens: " Ite in castellum, quod contra est, in quod introeuntes invenietis pullum asinae alligatum, cui nemo umquam hominum sedit; solvite illum et adducite.
LUKE|19|31|Et si quis vos interrogaverit: "Quare solvitis?", sic dicetis: "Dominus eum necessarium habet" ".
LUKE|19|32|Abierunt autem, qui missi erant, et invenerunt, sicut dixit illis.
LUKE|19|33|Solventibus autem illis pullum, dixerunt domini eius ad illos: " Quid solvitis pullum? ".
LUKE|19|34|At illi dixerunt: " Dominus eum necessarium habet ".
LUKE|19|35|Et duxerunt illum ad Iesum; et iactantes vestimenta sua supra pullum, imposuerunt Iesum.
LUKE|19|36|Eunte autem illo, substernebant vestimenta sua in via.
LUKE|19|37|Et cum appropinquaret iam ad descensum montis Oliveti, coeperunt omnis multitudo discipulorum gaudentes laudare Deum voce magna super omnibus, quas viderant, virtutibus
LUKE|19|38|dicentes: Benedictus, qui venit rex in nomine Domini!Pax in caelo, et gloria in excelsis! ".
LUKE|19|39|Et quidam pharisaeorum de turbis dixerunt ad illum: " Magister, increpa discipulos tuos! ".
LUKE|19|40|Et respondens dixit: " Dico vobis: Si hi tacuerint, lapides clamabunt!.
LUKE|19|41|Et ut appropinquavit, videns civitatem flevit super illam
LUKE|19|42|dicens: " Si cognovisses et tu in hac die, quae ad pacem tibi! Nunc autem abscondita sunt ab oculis tuis.
LUKE|19|43|Quia venient dies in te, et circumdabunt te inimici tui vallo et obsidebunt te et coangustabunt te undique
LUKE|19|44|et ad terram prosternent te et filios tuos, qui in te sunt, et non relinquent in te lapidem super lapidem, eo quod non cognoveris tempus visitationis tuae ".
LUKE|19|45|Et ingressus in templum, coepit eicere vendentes
LUKE|19|46|dicens illis: " Scriptum est: "Et erit domus mea domus orationis". Vos autem fecistis illam speluncam latronum ".
LUKE|19|47|Et erat docens cotidie in templo. Principes autem sacerdotum et scribae et principes plebis quaerebant illum perdere
LUKE|19|48|et non inveniebant quid facerent; omnis enim populus suspensus erat audiens illum.
LUKE|20|1|Et factum est in una dierum, docente illo populum in tem plo et evangelizante, supervenerunt principes sacerdotum et scribae cum senioribus
LUKE|20|2|et aiunt dicentes ad illum: " Dic nobis: In qua potestate haec facis, aut quis est qui dedit tibi hanc potestatem? ".
LUKE|20|3|Respondens autem dixit ad illos: " Interrogabo vos et ego verbum; et dicite mihi:
LUKE|20|4|Baptismum Ioannis de caelo erat an ex hominibus? ".
LUKE|20|5|At illi cogitabant inter se dicentes: " Si dixerimus: "De caelo", dicet: Quare non credidistis illi?;
LUKE|20|6|si autem dixerimus: "Ex hominibus", plebs universa lapidabit nos; certi sunt enim Ioannem prophetam esse ".
LUKE|20|7|Et responderunt se nescire unde esset.
LUKE|20|8|Et Iesus ait illis: " Neque ego dico vobis in qua potestate haec facio.
LUKE|20|9|Coepit autem dicere ad plebem parabolam hanc: " Homo plantavit vineam et locavit eam colonis et ipse peregre fuit multis temporibus.
LUKE|20|10|Et in tempore misit ad cultores servum, ut de fructu vineae darent illi; cultores autem caesum dimiserunt eum inanem.
LUKE|20|11|Et addidit alterum servum mittere; illi autem hunc quoque caedentes et afficientes contumelia dimiserunt inanem.
LUKE|20|12|Et addidit tertium mittere; qui et illum vulnerantes eiecerunt.
LUKE|20|13|Dixit autem dominus vineae: "Quid faciam? Mittam filium meum dilectum; forsitan hunc verebuntur".
LUKE|20|14|Quem cum vidissent coloni, cogitaverunt inter se dicentes: "Hic est heres. Occidamus illum, ut nostra fiat hereditas".
LUKE|20|15|Et eiectum illum extra vineam occiderunt. Quid ergo faciet illis dominus vineae?
LUKE|20|16|Veniet et perdet colonos istos et dabit vineam aliis ".Quo audito, dixerunt: " Absit! ".
LUKE|20|17|Ille autem aspiciens eos ait: " Quid est ergo hoc, quod scriptum est:Lapidem quem reprobaverunt aedificantes,hic factus est in caput anguli"?
LUKE|20|18|Omnis, qui ceciderit supra illum lapidem, conquassabitur; supra quem autem ceciderit, comminuet illum ".
LUKE|20|19|Et quaerebant scribae et principes sacerdotum mittere in illum manus in illa hora et timuerunt populum; cognoverunt enim quod ad ipsos dixerit similitudinem istam.
LUKE|20|20|Et observantes miserunt insidiatores, qui se iustos simularent, ut caperent eum in sermone, et sic traderent illum principatui et potestati praesidis.
LUKE|20|21|Et interrogaverunt illum dicentes: " Magister, scimus quia recte dicis et doces et non accipis personam, sed in veritate viam Dei doces.
LUKE|20|22|Licet nobis dare tributum Caesari an non? ".
LUKE|20|23|Considerans autem dolum illorum dixit ad eos:
LUKE|20|24|" Ostendite mihi denarium. Cuius habet imaginem et inscriptionem? ".
LUKE|20|25|At illi dixerunt: " Caesaris ". Et ait illis: " Reddite ergo, quae Caesaris sunt, Caesari et, quae Dei sunt, Deo ".
LUKE|20|26|Et non potuerunt verbum eius reprehendere coram plebe et mirati in responso eius tacuerunt.
LUKE|20|27|Accesserunt autem quidam sadducaeorum, qui negant esse resurrectionem, et interrogaverunt eum
LUKE|20|28|dicentes: " Magister, Moyses scripsit nobis, si frater alicuius mortuus fuerit habens uxorem et hic sine filiis fuerit, ut accipiat eam frater eius uxorem et suscitet semen fratri suo.
LUKE|20|29|Septem ergo fratres erant: et primus accepit uxorem et mortuus est sine filiis;
LUKE|20|30|et sequens
LUKE|20|31|et tertius accepit illam, similiter autem et septem non reliquerunt filios et mortui sunt.
LUKE|20|32|Novissima mortua est et mulier.
LUKE|20|33|Mulier ergo in resurrectione cuius eorum erit uxor? Si quidem septem habuerunt eam uxorem ".
LUKE|20|34|Et ait illis Iesus: " Filii saeculi huius nubunt et traduntur ad nuptias;
LUKE|20|35|illi autem, qui digni habentur saeculo illo et resurrectione ex mortuis, neque nubunt neque ducunt uxores.
LUKE|20|36|Neque enim ultra mori possunt: aequales enim angelis sunt et filii sunt Dei, cum sint filii resurrectionis.
LUKE|20|37|Quia vero resurgant mortui, et Moyses ostendit secus rubum, sicut dicit: "Dominum Deum Abraham et Deum Isaac et Deum Iacob".
LUKE|20|38|Deus autem non est mortuorum sed vivorum: omnes enim vivunt ei ".
LUKE|20|39|Respondentes autem quidam scribarum dixerunt: " Magister, bene dixisti.
LUKE|20|40|Et amplius non audebant eum quidquam interrogare.
LUKE|20|41|Dixit autem ad illos: " Quomodo dicunt Christum filium David esse?
LUKE|20|42|Ipse enim David dicit in libro Psalmorum:Dixit Dominus Domino meo: Sede a dextris meis,
LUKE|20|43|donec ponam inimicos tuos scabellum pedum tuorum".
LUKE|20|44|David ergo Dominum illum vocat; et quomodo filius eius est? ".
LUKE|20|45|Audiente autem omni populo, dixit discipulis suis:
LUKE|20|46|" Attendite a scribis, qui volunt ambulare in stolis et amant salutationes in foro et primas cathedras in synagogis et primos discubitus in conviviis,
LUKE|20|47|qui devorant domos viduarum et simulant longam orationem. Hi accipient damnationem maiorem ".
LUKE|21|1|Respiciens autem vidit eos, qui mittebant munera sua in gazophylacium, divites.
LUKE|21|2|Vidit autem quandam viduam pauperculam mittentem illuc minuta duo
LUKE|21|3|et dixit: " Vere dico vobis: Vidua haec pauper plus quam omnes misit.
LUKE|21|4|Nam omnes hi ex abundantia sua miserunt in munera; haec autem ex inopia sua omnem victum suum, quem habebat, misit ".
LUKE|21|5|Et quibusdam dicentibus de templo, quod lapidibus bonis et donis ornatum, esset dixit:
LUKE|21|6|" Haec quae videtis, venient dies, in quibus non relinquetur lapis super lapidem, qui non destruatur ".
LUKE|21|7|Interrogaverunt autem illum dicentes: " Praeceptor, quando ergo haec erunt, et quod signum, cum fieri incipient? ".
LUKE|21|8|Qui dixit: " Videte, ne seducamini. Multi enim venient in nomine meo dicentes: "Ego sum" et: "Tempus appropinquavit". Nolite ergo ire post illos.
LUKE|21|9|Cum autem audieritis proelia et seditiones, nolite terreri; oportet enim primum haec fieri, sed non statim finis ".
LUKE|21|10|Tunc dicebat illis: " Surget gens contra gentem, et regnum adversus regnum;
LUKE|21|11|et terrae motus magni et per loca fames et pestilentiae erunt, terroresque et de caelo signa magna erunt.
LUKE|21|12|Sed ante haec omnia inicient vobis manus suas et persequentur tradentes in synagogas et custodias, et trahemini ad reges et praesides propter nomen meum;
LUKE|21|13|continget autem vobis in testimonium.
LUKE|21|14|Ponite ergo in cordibus vestris non praemeditari quemadmodum respondeatis;
LUKE|21|15|ego enim dabo vobis os et sapientiam, cui non poterunt resistere vel contradicere omnes adversarii vestri.
LUKE|21|16|Trademini autem et a parentibus et fratribus et cognatis et amicis, et morte afficient ex vobis,
LUKE|21|17|et eritis odio omnibus propter nomen meum.
LUKE|21|18|Et capillus de capite vestro non peribit.
LUKE|21|19|In patientia vestra possidebitis animas vestras.
LUKE|21|20|Cum autem videritis circumdari ab exercitu Ierusalem, tunc scitote quia appropinquavit desolatio eius.
LUKE|21|21|Tunc, qui in Iudaea sunt, fugiant in montes; et, qui in medio eius, discedant; et, qui in regionibus, non intrent in eam.
LUKE|21|22|Quia dies ultionis hi sunt, ut impleantur omnia, quae scripta sunt.
LUKE|21|23|Vae autem praegnantibus et nutrientibus in illis diebus! Erit enim pressura magna super terram et ira populo huic,
LUKE|21|24|et cadent in ore gladii et captivi ducentur in omnes gentes, et Ierusalem calcabitur a gentibus, donec impleantur tempora nationum.
LUKE|21|25|Et erunt signa in sole et luna et stellis, et super terram pressura gentium prae confusione sonitus maris et fluctuum,
LUKE|21|26|arescentibus hominibus prae timore et exspectatione eorum, quae supervenient orbi, nam virtutes caelorum movebuntur.
LUKE|21|27|Et tunc videbunt Filium hominis venientem in nube cum potestate et gloria magna.
LUKE|21|28|His autem fieri incipientibus, respicite et levate capita vestra, quoniam appropinquat redemptio vestra ".
LUKE|21|29|Et dixit illis similitudinem: " Videte ficulneam et omnes arbores:
LUKE|21|30|cum iam germinaverint, videntes vosmetipsi scitis quia iam prope est aestas.
LUKE|21|31|Ita et vos, cum videritis haec fieri, scitote quoniam prope est regnum Dei.
LUKE|21|32|Amen dico vobis: Non praeteribit generatio haec, donec omnia fiant.
LUKE|21|33|Caelum et terra transibunt, verba autem mea non transibunt.
LUKE|21|34|Attendite autem vobis, ne forte graventur corda vestra in crapula et ebrietate et curis huius vitae, et superveniat in vos repentina dies illa;
LUKE|21|35|tamquam laqueus enim superveniet in omnes, qui sedent super faciem omnis terrae.
LUKE|21|36|Vigilate itaque omni tempore orantes, ut possitis fugere ista omnia, quae futura sunt, et stare ante Filium hominis ".
LUKE|21|37|Erat autem diebus docens in templo, noctibus vero exiens morabatur in monte, qui vocatur Oliveti.
LUKE|21|38|Et omnis populus manicabat ad eum in templo audire eum.
LUKE|22|1|Appropinquabat autem dies festus Azymorum, qui dici tur Pascha.
LUKE|22|2|Et quaerebant principes sacerdotum et scribae quomodo eum interficerent; timebant vero plebem.
LUKE|22|3|Intravit autem Satanas in Iudam, qui cognominabatur Iscarioth, unum de Duodecim;
LUKE|22|4|et abiit et locutus est cum principibus sacerdotum et magistratibus, quemadmodum illum traderet eis.
LUKE|22|5|Et gavisi sunt et pacti sunt pecuniam illi dare.
LUKE|22|6|Et spopondit et quaerebat opportunitatem, ut eis traderet illum sine turba.
LUKE|22|7|Venit autem dies Azymorum, in qua necesse erat occidi Pascha.
LUKE|22|8|Et misit Petrum et Ioannem dicens: " Euntes parate nobis Pascha, ut manducemus ".
LUKE|22|9|At illi dixerunt ei: "Ubi vis paremus? ".
LUKE|22|10|Et dixit ad eos: " Ecce, introeuntibus vobis in civitatem, occurret vobis homo amphoram aquae portans; sequimini eum in domum, in quam intrat.
LUKE|22|11|Et dicetis patri familias domus: "Dicit tibi Magister: Ubi est deversorium, ubi Pascha cum discipulis meis manducem?".
LUKE|22|12|Ipse vobis ostendet cenaculum magnum stratum; ibi parate ".
LUKE|22|13|Euntes autem invenerunt, sicut dixit illis, et paraverunt Pascha.
LUKE|22|14|Et cum facta esset hora, discubuit, et apostoli cum eo.
LUKE|22|15|Et ait illis: " Desiderio desideravi hoc Pascha manducare vobiscum, antequam patiar.
LUKE|22|16|Dico enim vobis: Non manducabo illud, donec impleatur in regno Dei ".
LUKE|22|17|Et accepto calice, gratias egit et dixit: " Accipite hoc et dividite inter vos.
LUKE|22|18|Dico enim vobis: Non bibam amodo de generatione vitis, donec regnum Dei veniat ".
LUKE|22|19|Et accepto pane, gratias egit et fregit et dedit eis dicens: " Hoc est corpus meum, quod pro vobis datur. Hoc facite in meam commemorationem ".
LUKE|22|20|Similiter et calicem, postquam cenavit, dicens: " Hic calix novum testamentum est in sanguine meo, qui pro vobis funditur.
LUKE|22|21|Verumtamen ecce manus tradentis me mecum est in mensa;
LUKE|22|22|et quidem Filius hominis, secundum quod definitum est, vadit; verumtamen vae illi homini, per quem traditur! ".
LUKE|22|23|Et ipsi coeperunt quaerere inter se, quis esset ex eis, qui hoc facturus esset.
LUKE|22|24|Facta est autem et contentio inter eos, quis eorum videretur esse maior.
LUKE|22|25|Dixit autem eis: " Reges gentium dominantur eorum; et, qui potestatem habent super eos, benefici vocantur.
LUKE|22|26|Vos autem non sic, sed qui maior est in vobis, fiat sicut iunior; et, qui praecessor est, sicut ministrator.
LUKE|22|27|Nam quis maior est: qui recumbit, an qui ministrat? Nonne qui recumbit? Ego autem in medio vestrum sum, sicut qui ministrat.
LUKE|22|28|Vos autem estis, qui permansistis mecum in tentationibus meis;
LUKE|22|29|et ego dispono vobis, sicut disposuit mihi Pater meus regnum,
LUKE|22|30|ut edatis et bibatis super mensam meam in regno meo et sedeatis super thronos iudicantes duodecim tribus Israel.
LUKE|22|31|Simon, Simon, ecce Satanas expetivit vos, ut cribraret sicut triticum;
LUKE|22|32|ego autem rogavi pro te, ut non deficiat fides tua. Et tu, aliquando conversus, confirma fratres tuos ".
LUKE|22|33|Qui dixit ei: " Domine, tecum paratus sum et in carcerem et in mortem ire ".
LUKE|22|34|Et ille dixit: " Dico tibi, Petre, non cantabit hodie gallus, donec ter abneges nosse me ".
LUKE|22|35|Et dixit eis: " Quando misi vos sine sacculo et pera et calceamentis, numquid aliquid defuit vobis? ". At illi dixerunt: " Nihil ".
LUKE|22|36|Dixit ergo eis: " Sed nunc, qui habet sacculum, tollat, similiter et peram; et, qui non habet, vendat tunicam suam et emat gladium.
LUKE|22|37|Dico enim vobis: Hoc, quod scriptum est, oportet impleri in me, illud: Cum iniustis deputatus est". Etenim ea, quae sunt de me, adimpletionem habent ".
LUKE|22|38|At illi dixerunt: " Domine, ecce gladii duo hic ". At ille dixit eis: " Satis est ".
LUKE|22|39|Et egressus ibat secundum consuetudinem in montem Olivarum; secuti sunt autem illum et discipuli.
LUKE|22|40|Et cum pervenisset ad locum, dixit illis: " Orate, ne intretis in tentationem ".
LUKE|22|41|Et ipse avulsus est ab eis, quantum iactus est lapidis, et, positis genibus, orabat
LUKE|22|42|dicens: " Pater, si vis, transfer calicem istum a me; verumtamen non mea voluntas sed tua fiat ".
LUKE|22|43|Apparuit autem illi angelus de caelo confortans eum. Et factus in agonia prolixius orabat.
LUKE|22|44|Et factus est sudor eius sicut guttae sanguinis decurrentis in terram.
LUKE|22|45|Et cum surrexisset ab oratione et venisset ad discipulos, invenit eos dormientes prae tristitia
LUKE|22|46|et ait illis: " Quid dormitis? Surgite; orate, ne intretis in tentationem ".
LUKE|22|47|Adhuc eo loquente, ecce turba; et, qui vocabatur Iudas, unus de Duodecim, antecedebat eos et appropinquavit Iesu, ut oscularetur eum.
LUKE|22|48|Iesus autem dixit ei: " Iuda, osculo Filium hominis tradis? ".
LUKE|22|49|Videntes autem hi, qui circa ipsum erant, quod futurum erat, dixerunt: Domine, si percutimus in gladio? ".
LUKE|22|50|Et percussit unus ex illis servum principis sacerdotum et amputavit auriculam eius dextram.
LUKE|22|51|Respondens autem Iesus ait: " Sinite usque huc! ". Et cum tetigisset auriculam eius, sanavit eum.
LUKE|22|52|Dixit autem Iesus ad eos, qui venerant ad se principes sacerdotum et magistratus templi et seniores: " Quasi ad latronem existis cum gladiis et fustibus?
LUKE|22|53|Cum cotidie vobiscum fuerim in templo, non extendistis manus in me; sed haec est hora vestra et potestas tenebrarum ".
LUKE|22|54|Comprehendentes autem eum, duxerunt et introduxerunt in domum principis sacerdotum. Petrus vero sequebatur a longe.
LUKE|22|55|Accenso autem igni in medio atrio et circumsedentibus illis, sedebat Petrus in medio eorum.
LUKE|22|56|Quem cum vidisset ancilla quaedam sedentem ad lumen et eum fuisset intuita, dixit:
LUKE|22|57|" Et hic cum illo erat! ". At ille negavit eum dicens:
LUKE|22|58|" Mulier, non novi illum! ". Et post pusillum alius videns eum dixit: " Et tu de illis es! ". Petrus vero ait: " O homo, non sum! ".
LUKE|22|59|Et intervallo facto quasi horae unius, alius quidam affirmabat dicens: Vere et hic cum illo erat, nam et Galilaeus est! ".
LUKE|22|60|Et ait Petrus: " Homo, nescio quid dicis! ". Et continuo adhuc illo loquente cantavit gallus.
LUKE|22|61|Et conversus Dominus respexit Petrum; et recordatus est Petrus verbi Domini, sicut dixit ei: " Priusquam gallus cantet hodie, ter me negabis ".
LUKE|22|62|Et egressus foras flevit amare.
LUKE|22|63|Et viri, qui tenebant illum, illudebant ei caedentes;
LUKE|22|64|et velaverunt eum et interrogabant eum dicentes: " Prophetiza: Quis est, qui te percussit? ".
LUKE|22|65|Et alia multa blasphemantes dicebant in eum.
LUKE|22|66|Et ut factus est dies, convenerunt seniores plebis et principes sacerdotum et scribae et duxerunt illum in concilium suum
LUKE|22|67|dicentes: " Si tu es Christus, dic nobis ". Et ait illis: " Si vobis dixero, non credetis;
LUKE|22|68|si autem interrogavero, non respondebitis mihi.
LUKE|22|69|Ex hoc autem erit Filius hominis sedens a dextris virtutis Dei ".
LUKE|22|70|Dixerunt autem omnes: " Tu ergo es Filius Dei? ". Qui ait ad illos: " Vos dicitis quia ego sum ".
LUKE|22|71|At illi dixerunt: " Quid adhuc desideramus testimonium? Ipsi enim audivimus de ore eius! ".
LUKE|23|1|Et surgens omnis multitudo eorum duxerunt illum ad Pi latum.
LUKE|23|2|Coeperunt autem accusare illum dicentes: " Hunc invenimus subvertentem gentem nostram et prohibentem tributa dare Caesari et dicentem se Christum regem esse ".
LUKE|23|3|Pilatus autem interrogavit eum dicens: " Tu es rex Iudaeorum? ". At ille respondens ait: " Tu dicis ".
LUKE|23|4|Ait autem Pilatus ad principes sacerdotum et turbas: " Nihil invenio causae in hoc homine ".
LUKE|23|5|At illi invalescebant dicentes: " Commovet populum docens per universam Iudaeam et in cipiens a Galilaea usque huc! ".
LUKE|23|6|Pilatus autem audiens interrogavit si homo Galilaeus esset;
LUKE|23|7|et ut cognovit quod de Herodis potestate esset, remisit eum ad Herodem, qui et ipse Hierosolymis erat illis diebus.
LUKE|23|8|Herodes autem, viso Iesu, gavisus est valde; erat enim cupiens ex multo tempore videre eum, eo quod audiret de illo et sperabat signum aliquod videre ab eo fieri.
LUKE|23|9|Interrogabat autem illum multis sermonibus; at ipse nihil illi respondebat.
LUKE|23|10|Stabant etiam principes sacerdotum et scribae constanter accusantes eum.
LUKE|23|11|Sprevit autem illum Herodes cum exercitu suo et illusit indutum veste alba et remisit ad Pilatum.
LUKE|23|12|Facti sunt autem amici inter se Herodes et Pilatus in ipsa die; nam antea inimici erant ad invicem.
LUKE|23|13|Pilatus autem, convocatis principibus sacerdotum et magistratibus et plebe,
LUKE|23|14|dixit ad illos: " Obtulistis mihi hunc hominem quasi avertentem populum, et ecce ego coram vobis interrogans nullam causam inveni in homine isto ex his, in quibus eum accusatis,
LUKE|23|15|sedneque Herodes; remisit enim illum ad nos. Et ecce nihil dignum morte actum est ei.
LUKE|23|16|Emendatum ergo illum dimittam ".
LUKE|23|17|()
LUKE|23|18|Exclamavit autem universa turba dicens: " Tolle hunc et dimitte nobis Barabbam! ",
LUKE|23|19|qui erat propter seditionem quandam factam in civitate et homicidium missus in carcerem.
LUKE|23|20|Iterum autem Pilatus locutus est ad illos volens dimittere Iesum,
LUKE|23|21|at illi succlamabant dicentes: " Crucifige, crucifige illum! ".
LUKE|23|22|Ille autem tertio dixit ad illos: " Quid enim mali fecit iste? Nullam causam mortis invenio in eo; corripiam ergo illum et dimittam ".
LUKE|23|23|At illi instabant vocibus magnis postulantes, ut crucifigeretur, et invalescebant voces eorum.
LUKE|23|24|Et Pilatus adiudicavit fieri petitionem eorum:
LUKE|23|25|dimisit autem eum, qui propter seditionem et homicidium missus fuerat in carcerem, quem petebant; Iesum vero tradidit voluntati eorum.
LUKE|23|26|Et cum abducerent eum, apprehenderunt Simonem quendam Cyrenensem venientem de villa et imposuerunt illi crucem portare post Iesum.
LUKE|23|27|Sequebatur autem illum multa turba populi et mulierum, quae plangebant et lamentabant eum.
LUKE|23|28|Conversus autem ad illas Iesus dixit: " Filiae Ierusalem, nolite flere super me, sed super vos ipsas flete et super filios vestros,
LUKE|23|29|quoniam ecce venient dies, in quibus dicent: "Beatae steriles et ventres, qui non genuerunt, et ubera, quae non lactaverunt!".
LUKE|23|30|Tunc incipient dicere montibus: "Cadite super nos!", et collibus: Operite nos!",
LUKE|23|31|quia si in viridi ligno haec faciunt, in arido quid fiet? ".
LUKE|23|32|Ducebantur autem et alii duo nequam cum eo, ut interficerentur.
LUKE|23|33|Et postquam venerunt in locum, qui vocatur Calvariae, ibi crucifixerunt eum et latrones, unum a dextris et alterum a sinistris.
LUKE|23|34|Iesus autem dicebat: " Pater, dimitte illis, non enim sciunt quid faciunt ".Dividentes vero vestimenta eius miserunt sortes.
LUKE|23|35|Et stabat populus exspectans. Et deridebant illum et principes dicentes: " Alios salvos fecit; se salvum faciat, si hic est Christus Dei electus! ".
LUKE|23|36|Illudebant autem ei et milites accedentes, acetum offerentes illi
LUKE|23|37|et dicentes: " Si tu es rex Iudaeorum, salvum te fac! ".
LUKE|23|38|Erat autem et superscriptio super illum: " Hic est rex Iudaeorum ".
LUKE|23|39|Unus autem de his, qui pendebant, latronibus blasphemabat eum dicens: " Nonne tu es Christus? Salvum fac temetipsum et nos! ".
LUKE|23|40|Respondens autem alter increpabat illum dicens: " Neque tu times Deum, quod in eadem damnatione es?
LUKE|23|41|Et nos quidem iuste, nam digna factis recipimus! Hic vero nihil mali gessit ".
LUKE|23|42|Et dicebat: " Iesu, memento mei, cum veneris in regnum tuum ".
LUKE|23|43|Et dixit illi: " Amen dico tibi: Hodie mecum eris in paradiso ".
LUKE|23|44|Et erat iam fere hora sexta, et tenebrae factae sunt in universa terra usque in horam nonam,
LUKE|23|45|et obscuratus est sol, et velum templi scissum est medium.
LUKE|23|46|Et clamans voce magna Iesus ait: " Pater, in manus tuas commendo spiritum meum "; et haec dicens exspiravit.
LUKE|23|47|Videns autem centurio, quod factum fuerat, glorificavit Deum dicens: " Vere hic homo iustus erat! ".
LUKE|23|48|Et omnis turba eorum, qui simul aderant ad spectaculum istud et videbant, quae fiebant, percutientes pectora sua revertebantur.
LUKE|23|49|Stabant autem omnes noti eius a longe et mulieres, quae secutae erant eum a Galilaea, haec videntes.
LUKE|23|50|Et ecce vir nomine Ioseph, qui erat decurio, vir bonus et iustus
LUKE|23|51|Chic non consenserat consilio et actibus eorum - ab Arimathaea civitate Iudaeorum, qui exspectabat regnum Dei,
LUKE|23|52|hic accessit ad Pilatum et petiit corpus Iesu
LUKE|23|53|et depositum involvit sindone et posuit eum in monumento exciso, in quo nondum quisquam positus fuerat.
LUKE|23|54|Et dies erat Parasceves, et sabbatum illucescebat.
LUKE|23|55|Subsecutae autem mulieres, quae cum ipso venerant de Galilaea, viderunt monumentum et quemadmodum positum erat corpus eius;
LUKE|23|56|et revertentes paraverunt aromata et unguenta et sabbato quidem siluerunt secundum mandatum.
LUKE|24|1|Prima autem sabbatorum, valde diluculo venerunt ad monumentum portantes, quae paraverant, aromata.
LUKE|24|2|Et invenerunt lapidem revolutum a monumento;
LUKE|24|3|et ingressae non invenerunt corpus Domini Iesu.
LUKE|24|4|Et factum est, dum mente haesitarent de isto, ecce duo viri steterunt secus illas in veste fulgenti.
LUKE|24|5|Cum timerent autem et declinarent vultum in terram, dixerunt ad illas: " Quid quaeritis viventem cum mortuis?
LUKE|24|6|Non est hic, sed surrexit. Recordamini qualiter locutus est vobis, cum adhuc in Galilaea esset,
LUKE|24|7|dicens: "Oportet Filium hominis tradi in manus hominum peccatorum et crucifigi et die tertia resurgere" ".
LUKE|24|8|Et recordatae sunt verborum eius
LUKE|24|9|et regressae a monumento nuntiaverunt haec omnia illis Undecim et ceteris omnibus.
LUKE|24|10|Erat autem Maria Magdalene et Ioanna et Maria Iacobi; et ceterae cum eis dicebant ad apostolos haec.
LUKE|24|11|Et visa sunt ante illos sicut deliramentum verba ista, et non credebant illis.
LUKE|24|12|Petrus autem surgens cucurrit ad monumentum et procumbens videt linteamina sola; et rediit ad sua mirans, quod factum fuerat.
LUKE|24|13|Et ecce duo ex illis ibant ipsa die in castellum, quod erat in spatio stadiorum sexaginta ab Ierusalem nomine Emmaus;
LUKE|24|14|et ipsi loquebantur ad invicem de his omnibus, quae acciderant.
LUKE|24|15|Et factum est, dum fabularentur et secum quaererent, et ipse Iesus appropinquans ibat cum illis;
LUKE|24|16|oculi autem illorum tenebantur, ne eum agnoscerent.
LUKE|24|17|Et ait ad illos: " Qui sunt hi sermones, quos confertis ad invicem ambulantes? ". Et steterunt tristes.
LUKE|24|18|Et respondens unus, cui nomen Cleopas, dixit ei: " Tu solus peregrinus es in Ierusalem et non cognovisti, quae facta sunt in illa his diebus? ".
LUKE|24|19|Quibus ille dixit: " Quae? ". Et illi dixerunt ei: " De Iesu Nazareno, qui fuit vir propheta, potens in opere et sermone coram Deo et omni populo;
LUKE|24|20|et quomodo eum tradiderunt summi sacerdotes et principes nostri in damnationem mortis et crucifixerunt eum.
LUKE|24|21|Nos autem sperabamus, quia ipse esset redempturus Israel; at nunc super haec omnia tertia dies hodie quod haec facta sunt.
LUKE|24|22|Sed et mulieres quaedam ex nostris terruerunt nos, quae ante lucem fuerunt ad monumentum
LUKE|24|23|et, non invento corpore eius, venerunt dicentes se etiam visionem angelorum vidisse, qui dicunt eum vivere.
LUKE|24|24|Et abierunt quidam ex nostris ad monumentum et ita invenerunt, sicut mulieres dixerunt, ipsum vero non viderunt ".
LUKE|24|25|Et ipse dixit ad eos: " O stulti et tardi corde ad credendum in omnibus, quae locuti sunt Prophetae!
LUKE|24|26|Nonne haec oportuit pati Christum et intrare in gloriam suam? ".
LUKE|24|27|Et incipiens a Moyse et omnibus Prophetis interpretabatur illis in omnibus Scripturis, quae de ipso erant.
LUKE|24|28|Et appropinquaverunt castello, quo ibant, et ipse se finxit longius ire.
LUKE|24|29|Et coegerunt illum dicentes: " Mane nobiscum, quoniam advesperascit, et inclinata est iam dies ". Et intravit, ut maneret cum illis.
LUKE|24|30|Et factum est, dum recumberet cum illis, accepit panem et benedixit ac fregit et porrigebat illis.
LUKE|24|31|Et aperti sunt oculi eorum, et cognoverunt eum; et ipse evanuit ab eis.
LUKE|24|32|Et dixerunt ad invicem: " Nonne cor nostrum ardens erat in nobis, dum loqueretur nobis in via et aperiret nobis Scripturas? ".
LUKE|24|33|Et surgentes eadem hora regressi sunt in Ierusalem et invenerunt congregatos Undecim et eos, qui cum ipsis erant,
LUKE|24|34|dicentes: " Surrexit Dominus vere et apparuit Simoni ".
LUKE|24|35|Et ipsi narrabant, quae gesta erant in via, et quomodo cognoverunt eum in fractione panis.
LUKE|24|36|Dum haec autem loquuntur, ipse stetit in medio eorum et dicit eis: " Pax vobis! ".
LUKE|24|37|Conturbati vero et conterriti existimabant se spiritum videre.
LUKE|24|38|Et dixit eis: " Quid turbati estis, et quare cogitationes ascendunt in corda vestra?
LUKE|24|39|Videte manus meas et pedes meos, quia ipse ego sum! Palpate me et videte, quia spiritus carnem et ossa non habet, sicut me videtis habere ".
LUKE|24|40|Et cum hoc dixisset, ostendit eis manus et pedes.
LUKE|24|41|Adhuc autem illis non credentibus prae gaudio et mirantibus, dixit eis: Habetis hic aliquid, quod manducetur? ".
LUKE|24|42|At illi obtulerunt ei partem piscis assi.
LUKE|24|43|Et sumens, coram eis manducavit.
LUKE|24|44|Et dixit ad eos: " Haec sunt verba, quae locutus sum ad vos, cum adhuc essem vobiscum, quoniam necesse est impleri omnia, quae scripta sunt in Lege Moysis et Prophetis et Psalmis de me ".
LUKE|24|45|Tunc aperuit illis sensum, ut intellegerent Scripturas.
LUKE|24|46|Et dixit eis: " Sic scriptum est, Christum pati et resurgere a mortuis die tertia,
LUKE|24|47|et praedicari in nomine eius paenitentiam in remissionem peccatorum in omnes gentes, incipientibus ab Ierusalem.
LUKE|24|48|Vos estis testes horum.
LUKE|24|49|Et ecce ego mitto promissum Patris mei in vos; vos autem sedete in civitate, quoadusque induamini virtutem ex alto ".
LUKE|24|50|Eduxit autem eos foras usque in Bethaniam et, elevatis manibus suis, benedixit eis.
LUKE|24|51|Et factum est, dum benediceret illis, recessit ab eis et ferebatur in caelum.
LUKE|24|52|Et ipsi adoraverunt eum et regressi sunt in Ierusalem cum gaudio magno
LUKE|24|53|et erant semper in templo benedicentes Deum.
JOHN|1|1|In principio erat Verbum, et Verbum erat apud Deum, et Deus erat Verbum.
JOHN|1|2|Hoc erat in principio apud Deum.
JOHN|1|3|Omnia per ipsum facta sunt, et sine ipso factum est nihil, quod factum est;
JOHN|1|4|in ipso vita erat, et vita erat lux hominum,
JOHN|1|5|et lux in tenebris lucet, et tenebrae eam non comprehenderunt.
JOHN|1|6|Fuit homo missus a Deo, cui nomen erat Ioannes;
JOHN|1|7|hic venit in testimonium, ut testimonium perhiberet de lumine, ut omnes crederent per illum.
JOHN|1|8|Non erat ille lux, sed ut testimonium perhiberet de lumine.
JOHN|1|9|Erat lux vera, quae illuminat omnem hominem, veniens in mundum.
JOHN|1|10|In mundo erat, et mundus per ipsum factus est, et mundus eum non cognovit.
JOHN|1|11|In propria venit, et sui eum non receperunt.
JOHN|1|12|Quotquot autem acceperunt eum, dedit eis potestatem filios Dei fieri, his, qui credunt in nomine eius,
JOHN|1|13|qui non ex sanguinibus neque ex voluntate carnis neque ex voluntate viri, sed ex Deo nati sunt.
JOHN|1|14|Et Verbum caro factum est et habitavit in nobis; et vidimus gloriam eius, gloriam quasi Unigeniti a Patre, plenum gratiae et veritatis.
JOHN|1|15|Ioannes testimonium perhibet de ipso et clamat dicens: " Hic erat, quem dixi: Qui post me venturus est, ante me factus est, quia prior me erat ".
JOHN|1|16|Et de plenitudine eius nos omnes accepimus, et gratiam pro gratia;
JOHN|1|17|quia lex per Moysen data est, gratia et veritas per Iesum Christum facta est.
JOHN|1|18|Deum nemo vidit umquam; unigenitus Deus, qui est in sinum Patris, ipse enarravit.
JOHN|1|19|Et hoc est testimonium Ioannis, quando miserunt ad eum Iudaei ab Hierosolymis sacerdotes et Levitas, ut interrogarent eum: " Tu quis es? ".
JOHN|1|20|Et confessus est et non negavit; et confessus est: " Non sum ego Christus ".
JOHN|1|21|Et interrogaverunt eum: " Quid ergo? Elias es tu? ". Et dicit: " Non sum ". " Propheta es tu? ". Et respondit: " Non ".
JOHN|1|22|Dixerunt ergo ei: " Quis es? Ut responsum demus his, qui miserunt nos. Quid dicis de teipso? ".
JOHN|1|23|Ait: Ego vox clamantis in deserto:Dirigite viam Domini",sicut dixit Isaias propheta ".
JOHN|1|24|Et qui missi fuerant, erant ex pharisaeis;
JOHN|1|25|et interrogaverunt eum et dixerunt ei: " Quid ergo baptizas, si tu non es Christus neque Elias neque propheta? ".
JOHN|1|26|Respondit eis Ioannes dicens: " Ego baptizo in aqua; medius vestrum stat, quem vos non scitis,
JOHN|1|27|qui post me venturus est, cuius ego non sum dignus, ut solvam eius corrigiam calceamenti ".
JOHN|1|28|Haec in Bethania facta sunt trans Iordanem, ubi erat Ioannes baptizans.
JOHN|1|29|Altera die videt Iesum venientem ad se et ait: " Ecce agnus Dei, qui tollit peccatum mundi.
JOHN|1|30|Hic est, de quo dixi: Post me venit vir, qui ante me factus est, quia prior me erat.
JOHN|1|31|Et ego nesciebam eum, sed ut manifestetur Israel, propterea veni ego in aqua baptizans ".
JOHN|1|32|Et testimonium perhibuit Ioannes dicens: " Vidi Spiritum descendentem quasi columbam de caelo, et mansit super eum;
JOHN|1|33|et ego nesciebam eum, sed, qui misit me baptizare in aqua, ille mihi dixit: "Super quem videris Spiritum descendentem et manentem super eum, hic est qui baptizat in Spiritu Sancto".
JOHN|1|34|Et ego vidi et testimonium perhibui quia hic est Filius Dei ".
JOHN|1|35|Altera die iterum stabat Ioannes et ex discipulis eius duo,
JOHN|1|36|et respiciens Iesum ambulantem dicit: " Ecce agnus Dei ".
JOHN|1|37|Et audierunt eum duo discipuli loquentem et secuti sunt Iesum.
JOHN|1|38|Conversus autem Iesus et videns eos sequentes se dicit eis: " Quid quaeritis? ". Qui dixerunt ei: " Rabbi - quod dicitur interpretatum Magister - ubi manes? ".
JOHN|1|39|Dicit eis: " Venite et videbitis ". Venerunt ergo et viderunt, ubi maneret, et apud eum manserunt die illo; hora erat quasi decima.
JOHN|1|40|Erat Andreas, frater Simonis Petri, unus ex duobus, qui audierant ab Ioanne et secuti fuerant eum.
JOHN|1|41|Invenit hic primum fratrem suum Simonem et dicit ei: " Invenimus Messiam " - quod est interpretatum Christus C;
JOHN|1|42|adduxit eum ad Iesum. Intuitus eum Iesus dixit: " Tu es Simon filius Ioannis; tu vocaberis Cephas " - quod interpretatur Petrus C.
JOHN|1|43|In crastinum voluit exire in Galilaeam et invenit Philippum. Et dicit ei Iesus: " Sequere me ".
JOHN|1|44|Erat autem Philippus a Bethsaida, civitate Andreae et Petri.
JOHN|1|45|Invenit Philippus Nathanael et dicit ei: " Quem scripsit Moyses in Lege et Prophetae invenimus, Iesum filium Ioseph a Nazareth ".
JOHN|1|46|Et dixit ei Nathanael: " A Nazareth potest aliquid boni esse? ". Dicit ei Philippus: " Veni et vide ".
JOHN|1|47|Vidit Iesus Nathanael venientem ad se et dicit de eo: " Ecce vere Israelita, in quo dolus non est ".
JOHN|1|48|Dicit ei Nathanael: " Unde me nosti? ". Respondit Iesus et dixit ei: " Priusquam te Philippus vocaret, cum esses sub ficu, vidi te ".
JOHN|1|49|Respondit ei Nathanael: " Rabbi, tu es Filius Dei, tu rex es Israel! ".
JOHN|1|50|Respondit Iesus et dixit ei: " Quia dixi tibi: Vidi te sub ficu, credis? Maiora his videbis ".
JOHN|1|51|Et dicit ei: " Amen, amen dico vobis: Videbitis caelum apertum et angelos Dei ascendentes et descendentes supra Filium hominis ".
JOHN|2|1|Et die tertio nuptiae factae sunt in Cana Galilaeae, et erat mater Iesu ibi;
JOHN|2|2|vocatus est autem et Iesus et discipuli eius ad nuptias.
JOHN|2|3|Et deficiente vino, dicit mater Iesu ad eum: " Vinum non habent ".
JOHN|2|4|Et dicit ei Iesus: " Quid mihi et tibi, mulier? Nondum venit hora mea ".
JOHN|2|5|Dicit mater eius ministris: " Quodcumque dixerit vobis, facite ".
JOHN|2|6|Erant autem ibi lapideae hydriae sex positae secundum purificationem Iudaeorum, capientes singulae metretas binas vel ternas.
JOHN|2|7|Dicit eis Iesus: " Implete hydrias aqua ". Et impleverunt eas usque ad summum.
JOHN|2|8|Et dicit eis: " Haurite nunc et ferte architriclino ". Illi autem tulerunt.
JOHN|2|9|Ut autem gustavit architriclinus aquam vinum factam et non sciebat unde esset, ministri autem sciebant, qui haurierant aquam, vocat sponsum architriclinus
JOHN|2|10|et dicit ei: " Omnis homo primum bonum vinum ponit et, cum inebriati fuerint, id quod deterius est; tu servasti bonum vinum usque adhuc ".
JOHN|2|11|Hoc fecit initium signorum Iesus in Cana Galilaeae et manifestavit gloriam suam, et crediderunt in eum discipuli eius.
JOHN|2|12|Post hoc descendit Capharnaum ipse et mater eius et fratres eius et discipuli eius, et ibi manserunt non multis diebus.
JOHN|2|13|Et prope erat Pascha Iudaeorum, et ascendit Hierosolymam Iesus.
JOHN|2|14|Et invenit in templo vendentes boves et oves et columbas, et nummularios sedentes;
JOHN|2|15|et cum fecisset flagellum de funiculis, omnes eiecit de templo, oves quoque et boves, et nummulariorum effudit aes et mensas subvertit;
JOHN|2|16|et his, qui columbas vendebant, dixit: " Auferte ista hinc! Nolite facere domum Patris mei domum negotiationis ".
JOHN|2|17|Recordati sunt discipuli eius quia scriptum est: " Zelus domus tuae comedit me ".
JOHN|2|18|Responderunt ergo Iudaei et dixerunt ei: " Quod signum ostendis nobis, quia haec facis? ".
JOHN|2|19|Respondit Iesus et dixit eis: " Solvite templum hoc, et in tribus diebus excitabo illud ".
JOHN|2|20|Dixerunt ergo Iudaei: " Quadraginta et sex annis aedificatum est templum hoc, et tu tribus diebus excitabis illud? ".
JOHN|2|21|Ille autem dicebat de templo corporis sui.
JOHN|2|22|Cum ergo resurrexisset a mortuis, recordati sunt discipuli eius quia hoc dicebat, et crediderunt Scripturae et sermoni, quem dixit Iesus.
JOHN|2|23|Cum autem esset Hierosolymis in Pascha, in die festo, multi crediderunt in nomine eius, videntes signa eius, quae faciebat.
JOHN|2|24|Ipse autem Iesus non credebat semetipsum eis, eo quod ipse nosset omnes,
JOHN|2|25|et quia opus ei non erat, ut quis testimonium perhiberet de homine; ipse enim sciebat quid esset in homine.
JOHN|3|1|Erat autem homo ex pharisaeis, Nicodemus nomine, princeps Iudaeorum;
JOHN|3|2|hic venit ad eum nocte et dixit ei: " Rabbi, scimus quia a Deo venisti magister; nemo enim potest haec signa facere, quae tu facis, nisi fuerit Deus cum eo ".
JOHN|3|3|Respondit Iesus et dixit ei: " Amen, amen dico tibi: Nisi quis natus fuerit desuper, non potest videre regnum Dei ".
JOHN|3|4|Dicit ad eum Nicodemus: " Quomodo potest homo nasci, cum senex sit? Numquid potest in ventrem matris suae iterato introire et nasci? ".
JOHN|3|5|Respondit Iesus: " Amen, amen dico tibi: Nisi quis natus fuerit ex aqua et Spiritu, non potest introire in regnum Dei.
JOHN|3|6|Quod natum est ex carne, caro est; et, quod natum est ex Spiritu, spiritus est.
JOHN|3|7|Non mireris quia dixi tibi: Oportet vos nasci denuo.
JOHN|3|8|Spiritus, ubi vult, spirat, et vocem eius audis, sed non scis unde veniat et quo vadat; sic est omnis, qui natus est ex Spiritu ".
JOHN|3|9|Respondit Nicodemus et dixit ei: " Quomodo possunt haec fieri? ".
JOHN|3|10|Respondit Iesus et dixit ei: " Tu es magister Israel et haec ignoras?
JOHN|3|11|Amen, amen dico tibi: Quod scimus, loquimur et, quod vidimus, testamur; et testimonium nostrum non accipitis.
JOHN|3|12|Si terrena dixi vobis, et non creditis, quomodo, si dixero vobis caelestia, credetis?
JOHN|3|13|Et nemo ascendit in caelum, nisi qui descendit de caelo, Filius hominis.
JOHN|3|14|Et sicut Moyses exaltavit serpentem in deserto, ita exaltari oportet Filium hominis,
JOHN|3|15|ut omnis, qui credit, in ipso habeat vitam aeternam ".
JOHN|3|16|Sic enim dilexit Deus mundum, ut Filium suum unigenitum daret, ut omnis, qui credit in eum, non pereat, sed habeat vitam aeternam.
JOHN|3|17|Non enim misit Deus Filium in mundum, ut iudicet mundum, sed ut salvetur mundus per ipsum.
JOHN|3|18|Qui credit in eum, non iudicatur; qui autem non credit, iam iudicatus est, quia non credidit in nomen Unigeniti Filii Dei.
JOHN|3|19|Hoc est autem iudicium: Lux venit in mundum, et dilexerunt homines magis tenebras quam lucem; erant enim eorum mala opera.
JOHN|3|20|Omnis enim, qui mala agit, odit lucem et non venit ad lucem, ut non arguantur opera eius;
JOHN|3|21|qui autem facit veritatem, venit ad lucem, ut manifestentur eius opera, quia in Deo sunt facta.
JOHN|3|22|Post haec venit Iesus et discipuli eius in Iudaeam terram, et illic demorabatur cum eis et baptizabat.
JOHN|3|23|Erat autem et Ioannes baptizans in Enon iuxta Salim, quia aquae multae erant illic, et adveniebant et baptizabantur;
JOHN|3|24|nondum enim missus fuerat in carcerem Ioannes.
JOHN|3|25|Facta est ergo quaestio ex discipulis Ioannis cum Iudaeo de purificatione.
JOHN|3|26|Et venerunt ad Ioannem et dixerunt ei: " Rabbi, qui erat tecum trans Iordanem, cui tu testimonium perhibuisti, ecce hic baptizat, et omnes veniunt ad eum! ".
JOHN|3|27|Respondit Ioannes et dixit: " Non potest homo accipere quidquam, nisi fuerit ei datum de caelo.
JOHN|3|28|Ipsi vos mihi testimonium perhibetis, quod dixerim: Non sum ego Christus, sed: Missus sum ante illum.
JOHN|3|29|Qui habet sponsam, sponsus est; amicus autem sponsi, qui stat et audit eum, gaudio gaudet propter vocem sponsi. Hoc ergo gaudium meum impletum est.
JOHN|3|30|Illum oportet crescere, me autem minui ".
JOHN|3|31|Qui de sursum venit, supra omnes est; qui est de terra, de terra est et de terra loquitur. Qui de caelo venit, supra omnes est;
JOHN|3|32|et quod vidit et audivit, hoc testatur, et testimonium eius nemo accipit.
JOHN|3|33|Qui accipit eius testimonium, signavit quia Deus verax est.
JOHN|3|34|Quem enim misit Deus, verba Dei loquitur; non enim ad mensuram dat Spiritum.
JOHN|3|35|Pater diligit Filium et omnia dedit in manu eius.
JOHN|3|36|Qui credit in Filium, habet vitam aeternam; qui autem incredulus est Filio, non videbit vitam, sed ira Dei manet super eum.
JOHN|4|1|Ut ergo cognovit Iesus quia audierunt pharisaei quia Iesus plures discipulos facit et baptizat quam Ioannes
JOHN|4|2|- quamquam Iesus ipse non baptizaret sed discipuli eius -
JOHN|4|3|reliquit Iudaeam et abiit iterum in Galilaeam.
JOHN|4|4|Oportebat autem eum transire per Samariam.
JOHN|4|5|Venit ergo in civitatem Samariae, quae dicitur Sichar, iuxta praedium, quod dedit Iacob Ioseph filio suo;
JOHN|4|6|erat autem ibi fons Iacob. Iesus ergo fatigatus ex itinere sedebat sic super fontem; hora erat quasi sexta.
JOHN|4|7|Venit mulier de Samaria haurire aquam. Dicit ei Iesus: " Da mihi bibere;
JOHN|4|8|discipuli enim eius abierant in civitatem, ut cibos emerent.
JOHN|4|9|Dicit ergo ei mulier illa Samaritana: " Quomodo tu, Iudaeus cum sis, bibere a me poscis, quae sum mulier Samaritana? ". Non enim coutuntur Iudaei Samaritanis.
JOHN|4|10|Respondit Iesus et dixit ei: " Si scires donum Dei, et quis est, qui dicit tibi: "Da mihi bibere", tu forsitan petisses ab eo, et dedisset tibi aquam vivam ".
JOHN|4|11|Dicit ei mulier: " Domine, neque in quo haurias habes, et puteus altus est; unde ergo habes aquam vivam?
JOHN|4|12|Numquid tu maior es patre nostro Iacob, qui dedit nobis puteum, et ipse ex eo bibit et filii eius et pecora eius? ".
JOHN|4|13|Respondit Iesus et dixit ei: " Omnis, qui bibit ex aqua hac, sitiet iterum;
JOHN|4|14|qui autem biberit ex aqua, quam ego dabo ei, non sitiet in aeternum; sed aqua, quam dabo ei, fiet in eo fons aquae salientis in vitam aeternam.
JOHN|4|15|Dicit ad eum mulier: " Domine, da mihi hanc aquam, ut non sitiam neque veniam huc haurire ".
JOHN|4|16|Dicit ei: " Vade, voca virum tuum et veni huc ".
JOHN|4|17|Respondit mulier et dixit ei: " Non habeo virum ". Dicit ei Iesus: " Bene dixisti: "Non habeo virum";
JOHN|4|18|quinque enim viros habuisti, et nunc, quem habes, non est tuus vir. Hoc vere dixisti ".
JOHN|4|19|Dicit ei mulier: " Domine, video quia propheta es tu.
JOHN|4|20|Patres nostri in monte hoc adoraverunt, et vos dicitis quia in Hierosolymis est locus, ubi adorare oportet ".
JOHN|4|21|Dicit ei Iesus: " Crede mihi, mulier, quia venit hora, quando neque in monte hoc neque in Hierosolymis adorabitis Patrem.
JOHN|4|22|Vos adoratis, quod nescitis; nos adoramus, quod scimus, quia salus ex Iudaeis est.
JOHN|4|23|Sed venit hora, et nunc est, quando veri adoratores adorabunt Patrem in Spiritu et veritate; nam et Pater tales quaerit, qui adorent eum.
JOHN|4|24|Spiritus est Deus, et eos, qui adorant eum, in Spiritu et veritate oportet adorare ".
JOHN|4|25|Dicit ei mulier: " Scio quia Messias venit - qui dicitur Christus C; cum venerit ille, nobis annuntiabit omnia ".
JOHN|4|26|Dicit ei Iesus: " Ego sum, qui loquor tecum ".
JOHN|4|27|Et continuo venerunt discipuli eius et mirabantur quia cum muliere loquebatur; nemo tamen dixit: " Quid quaeris aut quid loqueris cum ea? ".
JOHN|4|28|Reliquit ergo hydriam suam mulier et abiit in civitatem et dicit illis hominibus:
JOHN|4|29|" Venite, videte hominem, qui dixit mihi omnia, quaecumque feci; numquid ipse est Christus? ".
JOHN|4|30|Exierunt de civitate et veniebant ad eum.
JOHN|4|31|Interea rogabant eum discipuli dicentes: " Rabbi, manduca ".
JOHN|4|32|Ille autem dixit eis: " Ego cibum habeo manducare, quem vos nescitis ".
JOHN|4|33|Dicebant ergo discipuli ad invicem: " Numquid aliquis attulit ei manducare? ".
JOHN|4|34|Dicit eis Iesus: " Meus cibus est, ut faciam voluntatem eius, qui misit me, et ut perficiam opus eius.
JOHN|4|35|Nonne vos dicitis: "Adhuc quattuor menses sunt, et messis venit"? Ecce dico vobis: Levate oculos vestros et videte regiones, quia albae sunt ad messem! Iam
JOHN|4|36|qui metit, mercedem accipit et congregat fructum in vitam aeternam, ut et qui seminat, simul gaudeat et qui metit.
JOHN|4|37|In hoc enim est verbum verum: Alius est qui seminat, et alius est qui metit.
JOHN|4|38|Ego misi vos metere, quod vos non laborastis; alii laboraverunt, et vos in laborem eorum introistis ".
JOHN|4|39|Ex civitate autem illa multi crediderunt in eum Samaritanorum propter verbum mulieris testimonium perhibentis: " Dixit mihi omnia, quaecumque feci! ".
JOHN|4|40|Cum venissent ergo ad illum Samaritani, rogaverunt eum, ut apud ipsos maneret; et mansit ibi duos dies.
JOHN|4|41|Et multo plures crediderunt propter sermonem eius;
JOHN|4|42|et mulieri dicebant: " Iam non propter tuam loquelam credimus; ipsi enim audivimus et scimus quia hic est vere Salvator mundi! ".
JOHN|4|43|Post duos autem dies exiit inde in Galilaeam;
JOHN|4|44|ipse enim Iesus testimonium perhibuit, quia propheta in sua patria honorem non habet.
JOHN|4|45|Cum ergo venisset in Galilaeam, exceperunt eum Galilaei, cum omnia vidissent, quae fecerat Hierosolymis in die festo; et ipsi enim venerant in diem festum.
JOHN|4|46|Venit ergo iterum in Cana Galilaeae, ubi fecit aquam vinum. Et erat quidam regius, cuius filius infirmabatur Capharnaum;
JOHN|4|47|hic, cum audisset quia Iesus advenerit a Iudaea in Galilaeam, abiit ad eum et rogabat, ut descenderet et sanaret filium eius; incipiebat enim mori.
JOHN|4|48|Dixit ergo Iesus ad eum: " Nisi signa et prodigia videritis, non credetis ".
JOHN|4|49|Dicit ad eum regius: " Domine, descende priusquam moriatur puer meus ".
JOHN|4|50|Dicit ei Iesus: " Vade. Filius tuus vivit ". Credidit homo sermoni, quem dixit ei Iesus, et ibat.
JOHN|4|51|Iam autem eo descendente, servi eius occurrerunt ei dicentes quia puer eius vivit.
JOHN|4|52|Interrogabat ergo horam ab eis, in qua melius habuerit. Dixerunt ergo ei: " Heri hora septima reliquit eum febris ".
JOHN|4|53|Cognovit ergo pater quia illa hora erat, in qua dixit ei Iesus: " Filius tuus vivit ", et credidit ipse et domus eius tota.
JOHN|4|54|Hoc iterum secundum signum fecit Iesus, cum venisset a Iudaea in Galilaeam.
JOHN|5|1|Post haec erat dies festus Iu daeorum, et ascendit Iesus Hie rosolymam.
JOHN|5|2|Est autem Hierosolymis, super Probatica, piscina, quae cognominatur HebraiceBethsatha, quinque porticus habens.
JOHN|5|3|In his iacebat multitudo languentium, caecorum, claudorum, aridorum.
JOHN|5|4|()
JOHN|5|5|Erat autem quidam homo ibi triginta et octo annos habens in infirmitate sua.
JOHN|5|6|Hunc cum vidisset Iesus iacentem, et cognovisset quia multum iam tempus habet, dicit ei: " Vis sanus fieri? ".
JOHN|5|7|Respondit ei languidus: " Domine, hominem non habeo, ut, cum turbata fuerit aqua, mittat me in piscinam; dum autem venio ego, alius ante me descendit ".
JOHN|5|8|Dicit ei Iesus: " Surge, tolle grabatum tuum et ambula ".
JOHN|5|9|Et statim sanus factus est homo et sustulit grabatum suum et ambulabat.Erat autem sabbatum in illo die.
JOHN|5|10|Dicebant ergo Iudaei illi, qui sanatus fuerat: " Sabbatum est, et non licet tibi tollere grabatum tuum ".
JOHN|5|11|Ille autem respondit eis: " Qui me fecit sanum, ille mihi dixit: "Tolle grabatum tuum et ambula" ".
JOHN|5|12|Interrogaverunt eum: " Quis est ille homo, qui dixit tibi: "Tolle et ambula"? ".
JOHN|5|13|Is autem, qui sanus fuerat effectus, nesciebat quis esset; Iesus enim declinavit a turba constituta in loco.
JOHN|5|14|Postea invenit eum Iesus in templo et dixit illi: " Ecce sanus factus es; iam noli peccare, ne deterius tibi aliquid contingat ".
JOHN|5|15|Abiit ille homo et nuntiavit Iudaeis quia Iesus esset, qui fecit eum sanum.
JOHN|5|16|Et propterea persequebantur Iudaei Iesum, quia haec faciebat in sabbato.
JOHN|5|17|Iesus autem respondit eis: " Pater meus usque modo operatur, et ego operor ".
JOHN|5|18|Propterea ergo magis quaerebant eum Iudaei interficere, quia non solum solvebat sabbatum, sed et Patrem suum dicebat Deum, aequalem se faciens Deo.
JOHN|5|19|Respondit itaque Iesus et dixit eis: " Amen, amen dico vobis: Non potest Filius a se facere quidquam, nisi quod viderit Patrem facientem; quaecumque enim ille faciat, haec et Filius similiter facit.
JOHN|5|20|Pater enim diligit Filium et omnia demonstrat ei, quae ipse facit, et maiora his demonstrabit ei opera, ut vos miremini.
JOHN|5|21|Sicut enim Pater suscitat mortuos et vivificat, sic et Filius, quos vult, vivificat.
JOHN|5|22|Neque enim Pater iudicat quemquam, sed iudicium omne dedit Filio,
JOHN|5|23|ut omnes honorificent Filium, sicut honorificant Patrem. Qui non honorificat Filium, non honorificat Patrem, qui misit illum.
JOHN|5|24|Amen, amen dico vobis: Qui verbum meum audit et credit ei, qui misit me, habet vitam aeternam et in iudicium non venit, sed transiit a morte in vitam.
JOHN|5|25|Amen, amen dico vobis: Venit hora, et nunc est, quando mortui audient vocem Filii Dei et, qui audierint, vivent.
JOHN|5|26|Sicut enim Pater habet vitam in semetipso, sic dedit et Filio vitam habere in semetipso;
JOHN|5|27|et potestatem dedit ei iudicium facere, quia Filius hominis est.
JOHN|5|28|Nolite mirari hoc, quia venit hora, in qua omnes, qui in monumentis sunt, audient vocem eius;
JOHN|5|29|et procedent, qui bona fecerunt, in resurrectionem vitae, qui vero mala egerunt, in resurrectionem iudicii.
JOHN|5|30|Non possum ego a meipso facere quidquam; sicut audio, iudico, et iudicium meum iustum est, quia non quaero voluntatem meam, sed voluntatem eius, qui misit me.
JOHN|5|31|Si ego testimonium perhibeo de meipso, testimonium meum non est verum;
JOHN|5|32|alius est, qui testimonium perhibet de me, et scio quia verum est testimonium, quod perhibet de me.
JOHN|5|33|Vos misistis ad Ioannem, et testimonium perhibuit veritati;
JOHN|5|34|ego autem non ab homine testimonium accipio, sed haec dico, ut vos salvi sitis.
JOHN|5|35|Ille erat lucerna ardens et lucens; vos autem voluistis exsultare ad horam in luce eius.
JOHN|5|36|Ego autem habeo testimonium maius Ioanne; opera enim, quae dedit mihi Pater, ut perficiam ea, ipsa opera, quae ego facio, testimonium perhibent de me, quia Pater me misit;
JOHN|5|37|et, qui misit me, Pater, ipse testimonium perhibuit de me. Neque vocem eius umquam audistis neque speciem eius vidistis;
JOHN|5|38|et verbum eius non habetis in vobis manens, quia, quem misit ille, huic vos non creditis.
JOHN|5|39|Scrutamini Scripturas, quia vos putatis in ipsis vitam aeternam habere; et illae sunt, quae testimonium perhibent de me.
JOHN|5|40|Et non vultis venire ad me, ut vitam habeatis.
JOHN|5|41|Gloriam ab hominibus non accipio,
JOHN|5|42|sed cognovi vos, quia dilectionem Dei non habetis in vobis.
JOHN|5|43|Ego veni in nomine Patris mei, et non accipitis me; si alius venerit in nomine suo, illum accipietis.
JOHN|5|44|Quomodo potestis vos credere, qui gloriam ab invicem accipitis, et gloriam, quae a solo est Deo, non quaeritis?
JOHN|5|45|Nolite putare quia ego accusaturus sim vos apud Patrem; est qui accuset vos: Moyses, in quo vos speratis.
JOHN|5|46|Si enim crederetis Moysi, crederetis forsitan et mihi; de me enim ille scripsit.
JOHN|5|47|Si autem illius litteris non creditis, quomodo meis verbis credetis? ".
JOHN|6|1|Post haec abiit Iesus trans mare Galilaeae, quod est Tiberiadis.
JOHN|6|2|Et sequebatur eum multitudo magna, quia videbant signa, quae faciebat super his, qui infirmabantur.
JOHN|6|3|Subiit autem in montem Iesus et ibi sedebat cum discipulis suis.
JOHN|6|4|Erat autem proximum Pascha, dies festus Iudaeorum.
JOHN|6|5|Cum sublevasset ergo oculos Iesus et vidisset quia multitudo magna venit ad eum, dicit ad Philippum: " Unde ememus panes, ut manducent hi? ".
JOHN|6|6|Hoc autem dicebat tentans eum; ipse enim sciebat quid esset facturus.
JOHN|6|7|Respondit ei Philippus: " Ducentorum denariorum panes non sufficiunt eis, ut unusquisque modicum quid accipiat! ".
JOHN|6|8|Dicit ei unus ex discipulis eius, Andreas frater Simonis Petri:
JOHN|6|9|" Est puer hic, qui habet quinque panes hordeaceos et duos pisces; sed haec quid sunt propter tantos? ".
JOHN|6|10|Dixit Iesus: " Facite homines discumbere ". Erat autem fenum multum in loco. Discubuerunt ergo viri numero quasi quinque milia.
JOHN|6|11|Accepit ergo panes Iesus et, cum gratias egisset, distribuit discumbentibus; similiter et ex piscibus, quantum volebant.
JOHN|6|12|Ut autem impleti sunt, dicit discipulis suis: " Colligite, quae superaverunt, fragmenta, ne quid pereat ".
JOHN|6|13|Collegerunt ergo et impleverunt duodecim cophinos fragmentorum ex quinque panibus hordeaceis, quae superfuerunt his, qui manducaverunt.
JOHN|6|14|Illi ergo homines, cum vidissent quod fecerat signum, dicebant: " Hic est vere propheta, qui venit in mundum! ".
JOHN|6|15|Iesus ergo, cum cognovisset quia venturi essent, ut raperent eum et facerent eum regem, secessit iterum in montem ipse solus.
JOHN|6|16|Ut autem sero factum est, descenderunt discipuli eius ad mare
JOHN|6|17|et, cum ascendissent navem, veniebant trans mare in Capharnaum. Et tenebrae iam factae erant, et nondum venerat ad eos Iesus.
JOHN|6|18|Mare autem, vento magno flante, exsurgebat.
JOHN|6|19|Cum remigassent ergo quasi stadia viginti quinque aut triginta, vident Iesum ambulantem super mare et proximum navi fieri, et timuerunt.
JOHN|6|20|Ille autem dicit eis: " Ego sum, nolite timere! ".
JOHN|6|21|Volebant ergo accipere eum in navem, et statim fuit navis ad terram, in quam ibant.
JOHN|6|22|Altera die turba, quae stabat trans mare, vidit quia navicula alia non erat ibi, nisi una, et quia non introisset cum discipulis suis Iesus in navem, sed soli discipuli eius abiissent;
JOHN|6|23|aliae supervenerunt naves a Tiberiade iuxta locum, ubi manducaverant panem, gratias agente Domino.
JOHN|6|24|Cum ergo vidisset turba quia Iesus non esset ibi neque discipuli eius, ascenderunt ipsi naviculas et venerunt Capharnaum quaerentes Iesum.
JOHN|6|25|Et cum invenissent eum trans mare, dixerunt ei: " Rabbi, quando huc venisti? ".
JOHN|6|26|Respondit eis Iesus et dixit: " Amen, amen dico vobis: Quaeritis me, non quia vidistis signa, sed quia manducastis ex panibus et saturati estis.
JOHN|6|27|Operamini non cibum, qui perit, sed cibum, qui permanet in vitam aeternam, quem Filius hominis vobis dabit; hunc enim Pater signavit Deus!.
JOHN|6|28|Dixerunt ergo ad eum: " Quid faciemus, ut operemur opera Dei? ".
JOHN|6|29|Respondit Iesus et dixit eis: " Hoc est opus Dei, ut credatis in eum, quem misit ille ".
JOHN|6|30|Dixerunt ergo ei: " Quod ergo tu facis signum, ut videamus et credamus tibi? Quid operaris?
JOHN|6|31|Patres nostri manna manducaverunt in deserto, sicut scriptum est: Panem de caelo dedit eis manducare" ".
JOHN|6|32|Dixit ergo eis Iesus: " Amen, amen dico vobis: Non Moyses dedit vobis panem de caelo, sed Pater meus dat vobis panem de caelo verum;
JOHN|6|33|panis enim Dei est, qui descendit de caelo et dat vitam mundo ".
JOHN|6|34|Dixerunt ergo ad eum: " Domine, semper da nobis panem hunc ".
JOHN|6|35|Dixit eis Iesus: " Ego sum panis vitae. Qui venit ad me, non esuriet; et, qui credit in me, non sitiet umquam.
JOHN|6|36|Sed dixi vobis, quia et vidistis me et non creditis.
JOHN|6|37|Omne, quod dat mihi Pater, ad me veniet; et eum, qui venit ad me, non eiciam foras,
JOHN|6|38|quia descendi de caelo, non ut faciam voluntatem meam sed voluntatem eius, qui misit me.
JOHN|6|39|Haec est autem voluntas eius, qui misit me, ut omne, quod dedit mihi, non perdam ex eo, sed resuscitem illud in novissimo die.
JOHN|6|40|Haec est enim voluntas Patris mei, ut omnis, qui videt Filium et credit in eum, habeat vitam aeternam; et resuscitabo ego eum in novissimo die ".
JOHN|6|41|Murmurabant ergo Iudaei de illo, quia dixisset: " Ego sum panis, qui de caelo descendi ",
JOHN|6|42|et dicebant: " Nonne hic est Iesus filius Ioseph, cuius nos novimus patrem et matrem? Quomodo dicit nunc: "De caelo descendi"? ".
JOHN|6|43|Respondit Iesus et dixit eis: " Nolite murmurare in invicem.
JOHN|6|44|Nemo potest venire ad me, nisi Pater, qui misit me, traxerit eum; et ego resuscitabo eum in novissimo die.
JOHN|6|45|Est scriptum in Prophetis: "Et erunt omnes docibiles Dei ". Omnis, qui audivit a Patre et didicit, venit ad me.
JOHN|6|46|Non quia Patrem vidit quisquam, nisi is qui est a Deo, hic vidit Patrem.
JOHN|6|47|Amen, amen dico vobis: Qui credit, habet vitam aeternam.
JOHN|6|48|Ego sum panis vitae.
JOHN|6|49|Patres vestri manducaverunt in deserto manna et mortui sunt.
JOHN|6|50|Hic est panis de caelo descendens, ut, si quis ex ipso manducaverit, non moriatur.
JOHN|6|51|Ego sum panis vivus, qui de caelo descendi. Si quis manducaverit ex hoc pane, vivet in aeternum; panis autem, quem ego dabo, caro mea est pro mundi vita ".
JOHN|6|52|Litigabant ergo Iudaei ad invicem dicentes: " Quomodo potest hic nobis carnem suam dare ad manducandum? ".
JOHN|6|53|Dixit ergo eis Iesus: " Amen, amen dico vobis: Nisi manducaveritis carnem Filii hominis et biberitis eius sanguinem, non habetis vitam in vobismetipsis.
JOHN|6|54|Qui manducat meam carnem et bibit meum sanguinem, habet vitam aeternam; et ego resuscitabo eum in novissimo die.
JOHN|6|55|Caro enim mea verus est cibus, et sanguis meus verus est potus.
JOHN|6|56|Qui manducat meam carnem et bibit meum sanguinem, in me manet, et ego in illo.
JOHN|6|57|Sicut misit me vivens Pater, et ego vivo propter Patrem; et, qui manducat me, et ipse vivet propter me.
JOHN|6|58|Hic est panis, qui de caelo descendit, non sicut manducaverunt patres et mortui sunt; qui manducat hunc panem, vivet in aeternum ".
JOHN|6|59|Haec dixit in synagoga docens in Capharnaum.
JOHN|6|60|Multi ergo audientes ex discipulis eius dixerunt: " Durus est hic sermo! Quis potest eum audire? ".
JOHN|6|61|Sciens autem Iesus apud semetipsum quia murmurarent de hoc discipuli eius, dixit eis: " Hoc vos scandalizat?
JOHN|6|62|Si ergo videritis Filium hominis ascendentem, ubi erat prius?
JOHN|6|63|Spiritus est, qui vivificat, caro non prodest quidquam; verba, quae ego locutus sum vobis, Spiritus sunt et vita sunt.
JOHN|6|64|Sed sunt quidam ex vobis, qui non credunt ". Sciebat enim ab initio Iesus, qui essent non credentes, et quis traditurus esset eum.
JOHN|6|65|Et dicebat: " Propterea dixi vobis: Nemo potest venire ad me, nisi fuerit ei datum a Patre ".
JOHN|6|66|Ex hoc multi discipulorum eius abierunt retro et iam non cum illo ambulabant.
JOHN|6|67|Dixit ergo Iesus ad Duodecim: " Numquid et vos vultis abire? ".
JOHN|6|68|Respondit ei Simon Petrus: " Domine, ad quem ibimus? Verba vitae aeternae habes;
JOHN|6|69|et nos credidimus et cognovimus quia tu es Sanctus Dei ".
JOHN|6|70|Respondit eis Iesus: " Nonne ego vos Duodecim elegi? Et ex vobis unus Diabolus est ".
JOHN|6|71|Dicebat autem Iudam Simonis Iscariotis; hic enim erat traditurus eum, cum esset unus ex Duodecim.
JOHN|7|1|Et post haec ambulabat Iesus in Galilaeam; non enim volebat in Iudaeam ambulare, quia quaerebant eum Iudaei interficere.
JOHN|7|2|Erat autem in proximo dies festus Iudaeorum, Scenopegia.
JOHN|7|3|Dixerunt ergo ad eum fratres eius: " Transi hinc et vade in Iudaeam, ut et discipuli tui videant opera tua, quae facis.
JOHN|7|4|Nemo quippe in occulto quid facit et quaerit ipse in palam esse. Si haec facis, manifesta teipsum mundo ".
JOHN|7|5|Neque enim fratres eius credebant in eum.
JOHN|7|6|Dicit ergo eis Iesus: " Tempus meum nondum adest, tempus autem vestrum semer est paratum.
JOHN|7|7|Non potest mundus odisse vos; me autem odit, quia ego testimonium perhibeo de illo, quia opera eius mala sunt.
JOHN|7|8|Vos ascendite ad diem festum; ego non ascendo ad diem festum istum, quia meum tempus nondum impletum est ".
JOHN|7|9|Haec autem cum dixisset, ipse mansit in Galilaea.
JOHN|7|10|Ut autem ascenderunt fratres eius ad diem festum, tunc et ipse ascendit, non manifeste sed quasi in occulto.
JOHN|7|11|Iudaei ergo quaerebant eum in die festo et dicebant: " Ubi est ille? ".
JOHN|7|12|Et murmur multus de eo erat in turba. Alii quidem dicebant: " Bonus est! "; alii autem dicebant: " Non, sed seducit turbam! ".
JOHN|7|13|Nemo tamen palam loquebatur de illo propter metum Iudaeorum.
JOHN|7|14|Iam autem die festo mediante, ascendit Iesus in templum et docebat.
JOHN|7|15|Mirabantur ergo Iudaei dicentes: " Quomodo hic litteras scit, cum non didicerit? ".
JOHN|7|16|Respondit ergo eis Iesus et dixit: " Mea doctrina non est mea sed eius, qui misit me.
JOHN|7|17|Si quis voluerit voluntatem eius facere, cognoscet de doctrina utrum ex Deo sit, an ego a meipso loquar.
JOHN|7|18|Qui a semetipso loquitur, gloriam propriam quaerit; qui autem quaerit gloriam eius, qui misit illum, hic verax est, et iniustitia in illo non est.
JOHN|7|19|Nonne Moyses dedit vobis legem? Et nemo ex vobis facit legem. Quid me quaeritis interficere? ".
JOHN|7|20|Respondit turba: " Daemonium habes! Quis te quaerit interficere? ".
JOHN|7|21|Respondit Iesus et dixit eis: " Unum opus feci, et omnes miramini.
JOHN|7|22|Propterea Moyses dedit vobis circumcisionem - non quia ex Moyse est sed ex patribus - et in sabbato circumciditis hominem.
JOHN|7|23|Si circumcisionem accipit homo in sabbato, ut non solvatur lex Moysis, mihi indignamini, quia totum hominem sanum feci in sabbato?
JOHN|7|24|Nolite iudicare secundum faciem, sed iustum iudicium iudicate ".
JOHN|7|25|Dicebant ergo quidam ex Hierosolymitis: " Nonne hic est, quem quaerunt interficere?
JOHN|7|26|Et ecce palam loquitur, et nihil ei dicunt. Numquid vere cognoverunt principes quia hic est Christus?
JOHN|7|27|Sed hunc scimus unde sit, Christus autem cum venerit, nemo scit unde sit ".
JOHN|7|28|Clamavit ergo docens in templo Iesus et dicens: " Et me scitis et unde sim scitis. Et a meipso non veni, sed est verus, qui misit me, quem vos non scitis.
JOHN|7|29|Ego scio eum, quia ab ipso sum, et ipse me misit ".
JOHN|7|30|Quaerebant ergo eum apprehendere, et nemo misit in illum manus, quia nondum venerat hora eius.
JOHN|7|31|De turba autem multi crediderunt in eum et dicebant: " Christus cum venerit, numquid plura signa faciet quam quae hic fecit? ".
JOHN|7|32|Audierunt pharisaei turbam murmurantem de illo haec et miserunt pontifices et pharisaei ministros, ut apprehenderent eum.
JOHN|7|33|Dixit ergo Iesus: " Adhuc modicum tempus vobiscum sum et vado ad eum, qui misit me.
JOHN|7|34|Quaeretis me et non invenietis; et ubi sum ego, vos non potestis venire.
JOHN|7|35|Dixerunt ergo Iudaei ad seipsos: " Quo hic iturus est, quia nos non inveniemus eum? Numquid in dispersionem Graecorum iturus est et docturus Graecos?
JOHN|7|36|Quis est hic sermo, quem dixit: "Quaeretis me et non invenietis" et: Ubi sum ego, vos non potestis venire"? ".
JOHN|7|37|In novissimo autem die magno festivitatis stabat Iesus et clamavit dicens: " Si quis sitit, veniat ad me et bibat,
JOHN|7|38|qui credit in me. Sicut dixit Scriptura, flumina de ventre eius fluent aquae vivae ".
JOHN|7|39|Hoc autem dixit de Spiritu, quem accepturi erant qui crediderant in eum. Nondum enim erat Spiritus, quia Iesus nondum fuerat glorificatus.
JOHN|7|40|Ex illa ergo turba, cum audissent hos sermones, dicebant: " Hic est vere propheta! ";
JOHN|7|41|alii dicebant: " Hic est Christus! "; quidam autem dicebant: " Numquid a Galilaea Christus venit?
JOHN|7|42|Nonne Scriptura dixit: "Ex semine David et de Bethlehem castello, ubi erat David, venit Christus"? ".
JOHN|7|43|Dissensio itaque facta est in turba propter eum.
JOHN|7|44|Quidam autem ex ipsis volebant apprehendere eum, sed nemo misit super illum manus.
JOHN|7|45|Venerunt ergo ministri ad pontifices et pharisaeos; et dixerunt eis illi: " Quare non adduxistis eum? ".
JOHN|7|46|Responderunt ministri: " Numquam sic locutus est homo ".
JOHN|7|47|Responderunt ergo eis pharisaei: " Numquid et vos seducti estis?
JOHN|7|48|Numquid aliquis ex principibus credidit in eum aut ex pharisaeis?
JOHN|7|49|Sed turba haec, quae non novit legem, maledicti sunt! ".
JOHN|7|50|Dicit Nicodemus ad eos, ille qui venit ad eum antea, qui unus erat ex ipsis:
JOHN|7|51|" Numquid lex nostra iudicat hominem, nisi audierit ab ipso prius et cognoverit quid faciat? ".
JOHN|7|52|Responderunt et dixerunt ei: " Numquid et tu ex Galilaea es? Scrutare et vide quia propheta a Galilaea non surgit! ".
JOHN|7|53|Et reversi sunt unusquisque in domum suam.
JOHN|8|1|Iesus autem perrexit in montem Oliveti.
JOHN|8|2|Diluculo autem iterum venit in templum, et omnis populus veniebat ad eum, et sedens docebat eos.
JOHN|8|3|Adducunt autem scribae et pharisaei mulierem in adulterio deprehensam et statuerunt eam in medio
JOHN|8|4|et dicunt ei: " Magister, haec mulier manifesto deprehensa est in adulterio.
JOHN|8|5|In lege autem Moyses mandavit nobis huiusmodi lapidare; tu ergo quid dicis? ".
JOHN|8|6|Hoc autem dicebant tentantes eum, ut possent accusare eum. Iesus autem inclinans se deorsum digito scribebat in terra.
JOHN|8|7|Cum autem perseverarent interrogantes eum, erexit se et dixit eis: " Qui sine peccato est vestrum, primus in illam lapidem mittat ";
JOHN|8|8|et iterum se inclinans scribebat in terra.
JOHN|8|9|Audientes autem unus post unum exibant, incipientes a senioribus, et remansit solus, et mulier in medio stans.
JOHN|8|10|Erigens autem se Iesus dixit ei: " Mulier, ubi sunt? Nemo te condemnavit? ".
JOHN|8|11|Quae dixit: " Nemo, Domine ". Dixit autem Iesus: " Nec ego te condemno; vade et amplius iam noli peccare ".
JOHN|8|12|Iterum ergo locutus est eis Iesus dicens: " Ego sum lux mundi; qui sequitur me, non ambulabit in tenebris, sed habebit lucem vitae ".
JOHN|8|13|Dixerunt ergo ei pharisaei: " Tu de teipso testimonium perhibes; testimonium tuum non est verum ".
JOHN|8|14|Respondit Iesus et dixit eis: " Et si ego testimonium perhibeo de meipso, verum est testimonium meum, quia scio unde veni et quo vado; vos autem nescitis unde venio aut quo vado.
JOHN|8|15|Vos secundum carnem iudicatis, ego non iudico quemquam.
JOHN|8|16|Et si iudico ego, iudicium meum verum est, quia solus non sum, sed ego et, qui me misit, Pater.
JOHN|8|17|Sed et in lege vestra scriptum est, quia duorum hominum testimonium verum est.
JOHN|8|18|Ego sum, qui testimonium perhibeo de meipso, et testimonium perhibet de me, qui misit me, Pater ".
JOHN|8|19|Dicebant ergo ei: " Ubi est Pater tuus? ". Respondit Iesus: " Neque me scitis neque Patrem meum; si me sciretis, forsitan et Patrem meum sciretis.
JOHN|8|20|Haec verba locutus est in gazophylacio docens in templo; et nemo apprehendit eum, quia necdum venerat hora eius.
JOHN|8|21|Dixit ergo iterum eis: " Ego vado, et quaeretis me et in peccato vestro moriemini! Quo ego vado, vos non potestis venire ".
JOHN|8|22|Dicebant ergo Iudaei: " Numquid interficiet semetipsum, quia dicit: Quo ego vado, vos non potestis venire"? ".
JOHN|8|23|Et dicebat eis: " Vos de deorsum estis, ego de supernis sum; vos de mundo hoc estis, ego non sum de hoc mundo.
JOHN|8|24|Dixi ergo vobis quia moriemini in peccatis vestris; si enim non credideritis quia ego sum, moriemini in peccatis vestris ".
JOHN|8|25|Dicebant ergo ei: " Tu quis es? ". Dixit eis Iesus: " In principio: id quod et loquor vobis!
JOHN|8|26|Multa habeo de vobis loqui et iudicare; sed, qui misit me, verax est, et ego, quae audivi ab eo, haec loquor ad mundum ".
JOHN|8|27|Non cognoverunt quia Patrem eis dicebat.
JOHN|8|28|Dixit ergo eis Iesus: " Cum exaltaveritis Filium hominis, tunc cognoscetis quia ego sum et a meipso facio nihil, sed, sicut docuit me Pater, haec loquor.
JOHN|8|29|Et qui me misit, mecum est; non reliquit me solum, quia ego, quae placita sunt ei, facio semper ".
JOHN|8|30|Haec illo loquente, multi crediderunt in eum.
JOHN|8|31|Dicebat ergo Iesus ad eos, qui crediderunt ei, Iudaeos: " Si vos manseritis in sermone meo, vere discipuli mei estis
JOHN|8|32|et cognoscetis veritatem, et veritas liberabit vos ".
JOHN|8|33|Responderunt ei: " Semen Abrahae sumus et nemini servivimus umquam! Quomodo tu dicis: "Liberi fietis"? ".
JOHN|8|34|Respondit eis Iesus: " Amen, amen dico vobis: Omnis, qui facit peccatum, servus est peccati.
JOHN|8|35|Servus autem non manet in domo in aeternum; filius manet in aeternum.
JOHN|8|36|Si ergo Filius vos liberaverit, vere liberi eritis.
JOHN|8|37|Scio quia semen Abrahae estis; sed quaeritis me interficere, quia sermo meus non capit in vobis.
JOHN|8|38|Ego, quae vidi apud Patrem, loquor; et vos ergo, quae audivistis a patre, facitis ".
JOHN|8|39|Responderunt et dixerunt ei: " Pater noster Abraham est ". Dicit eis Iesus: " Si filii Abrahae essetis, opera Abrahae faceretis.
JOHN|8|40|Nunc autem quaeritis me interficere, hominem, qui veritatem vobis locutus sum, quam audivi a Deo; hoc Abraham non fecit.
JOHN|8|41|Vos facitis opera patris vestri ". Dixerunt itaque ei: " Nos ex fornicatione non sumus nati; unum patrem habemus Deum! ".
JOHN|8|42|Dixit eis Iesus: " Si Deus pater vester esset, diligeretis me; ego enim ex Deo processi et veni; neque enim a meipso veni, sed ille me misit.
JOHN|8|43|Quare loquelam meam non cognoscitis? Quia non potestis audire sermonem meum.
JOHN|8|44|Vos ex patre Diabolo estis et desideria patris vestri vultis facere. Ille homicida erat ab initio et in veritate non stabat, quia non est veritas in eo. Cum loquitur mendacium, ex propriis loquitur, quia mendax est et pater eius.
JOHN|8|45|Ego autem quia veritatem dico, non creditis mihi.
JOHN|8|46|Quis ex vobis arguit me de peccato? Si veritatem dico, quare vos non creditis mihi?
JOHN|8|47|Qui est ex Deo, verba Dei audit; propterea vos non auditis, quia ex Deo non estis ".
JOHN|8|48|Responderunt Iudaei et dixerunt ei: " Nonne bene dicimus nos, quia Samaritanus es tu et daemonium habes? ".
JOHN|8|49|Respondit Iesus: " Ego daemonium non habeo, sed honorifico Patrem meum, et vos inhonoratis me.
JOHN|8|50|Ego autem non quaero gloriam meam; est qui quaerit et iudicat.
JOHN|8|51|Amen, amen dico vobis: Si quis sermonem meum servaverit, mortem non videbit in aeternum ".
JOHN|8|52|Dixerunt ergo ei Iudaei: " Nunc cognovimus quia daemonium habes. Abraham mortuus est et prophetae, et tu dicis: "Si quis sermonem meum servaverit, non gustabit mortem in aeternum".
JOHN|8|53|Numquid tu maior es patre nostro Abraham, qui mortuus est? Et prophetae mortui sunt! Quem teipsum facis? ".
JOHN|8|54|Respondit Iesus: " Si ego glorifico meipsum, gloria mea nihil est; est Pater meus, qui glorificat me, quem vos dicitis: "Deus noster est!",
JOHN|8|55|et non cognovistis eum. Ego autem novi eum. Et si dixero: Non scio eum, ero similis vobis, mendax; sed scio eum et sermonem eius servo.
JOHN|8|56|Abraham pater vester exsultavit, ut videret diem meum; et vidit et gavisus est ".
JOHN|8|57|Dixerunt ergo Iudaei ad eum: " Quinquaginta annos nondum habes et Abraham vidisti? ".
JOHN|8|58|Dixit eis Iesus: " Amen, amen dico vobis: Antequam Abraham fieret, ego sum ".
JOHN|8|59|Tulerunt ergo lapides, ut iacerent in eum; Iesus autem abscondit se et exivit de templo.
JOHN|9|1|Et praeteriens vidit hominem caecum a nativitate.
JOHN|9|2|Et interro gaverunt eum discipuli sui dicentes: " Rabbi, quis peccavit, hic aut parentes eius, ut caecus nasceretur? ".
JOHN|9|3|Respondit Iesus: " Neque hic peccavit neque parentes eius, sed ut manifestentur opera Dei in illo.
JOHN|9|4|Nos oportet operari opera eius, qui misit me, donec dies est; venit nox, quando nemo potest operari.
JOHN|9|5|Quamdiu in mundo sum, lux sum mundi ".
JOHN|9|6|Haec cum dixisset, exspuit in terram et fecit lutum ex sputo et linivit lutum super oculos eius
JOHN|9|7|et dixit ei: " Vade, lava in natatoria Siloae! " - quod interpretatur Missus C. Abiit ergo et lavit et venit videns.
JOHN|9|8|Itaque vicini et, qui videbant eum prius quia mendicus erat, dicebant: " Nonne hic est, qui sedebat et mendicabat? ";
JOHN|9|9|alii dicebant: " Hic est! "; alii dicebant: " Nequaquam, sed similis est eius! ". Ille dicebat: " Ego sum! ".
JOHN|9|10|Dicebant ergo ei: " Quomodo igitur aperti sunt oculi tibi? ".
JOHN|9|11|Respondit ille: " Homo, qui dicitur Iesus, lutum fecit et unxit oculos meos et dixit mihi: "Vade ad Siloam et lava! ". Abii ergo et lavi et vidi.
JOHN|9|12|Et dixerunt ei: " Ubi est ille? ". Ait: " Nescio ".
JOHN|9|13|Adducunt eum ad pharisaeos, qui caecus fuerat.
JOHN|9|14|Erat autem sabbatum, in qua die lutum fecit Iesus et aperuit oculos eius.
JOHN|9|15|Iterum ergo interrogabant et eum pharisaei quomodo vidisset. Ille autem dixit eis: " Lutum posuit super oculos meos, et lavi et video ".
JOHN|9|16|Dicebant ergo ex pharisaeis quidam: " Non est hic homo a Deo, quia sabbatum non custodit! "; alii autem dicebant: " Quomodo potest homo peccator haec signa facere? ". Et schisma erat in eis.
JOHN|9|17|Dicunt ergo caeco iterum: " Tu quid dicis de eo quia aperuit oculos tuos? ". Ille autem dixit: " Propheta est! ".
JOHN|9|18|Non crediderunt ergo Iudaei de illo quia caecus fuisset et vidisset, donec vocaverunt parentes eius, qui viderat.
JOHN|9|19|Et interrogaverunt eos dicentes: " Hic est filius vester, quem vos dicitis quia caecus natus est? Quomodo ergo nunc videt? ".
JOHN|9|20|Responderunt ergo parentes eius et dixerunt: " Scimus quia hic est filius noster et quia caecus natus est.
JOHN|9|21|Quomodo autem nunc videat nescimus, aut quis eius aperuit oculos nos nescimus; ipsum interrogate. Aetatem habet; ipse de se loquetur! ".
JOHN|9|22|Haec dixerunt parentes eius, quia timebant Iudaeos; iam enim conspiraverant Iudaei, ut, si quis eum confiteretur Christum, extra synagogam fieret.
JOHN|9|23|Propterea parentes eius dixerunt: " Aetatem habet; ipsum interrogate!.
JOHN|9|24|Vocaverunt ergo rursum hominem, qui fuerat caecus, et dixerunt ei: " Da gloriam Deo! Nos scimus quia hic homo peccator est ".
JOHN|9|25|Respondit ergo ille: " Si peccator est nescio; unum scio quia, caecus cum essem, modo video ".
JOHN|9|26|Dixerunt ergo illi: " Quid fecit tibi? Quomodo aperuit oculos tuos? ".
JOHN|9|27|Respondit eis: " Dixi vobis iam, et non audistis; quid iterum vultis audire? Numquid et vos vultis discipuli eius fieri? ".
JOHN|9|28|Et maledixerunt ei et dixerunt: " Tu discipulus illius es, nos autem Moysis discipuli sumus.
JOHN|9|29|Nos scimus quia Moysi locutus est Deus; hunc autem nescimus unde sit ".
JOHN|9|30|Respondit homo et dixit eis: " In hoc enim mirabile est, quia vos nescitis unde sit, et aperuit meos oculos!
JOHN|9|31|Scimus quia peccatores Deus non audit; sed, si quis Dei cultor est et voluntatem eius facit, hunc exaudit.
JOHN|9|32|A saeculo non est auditum quia aperuit quis oculos caeci nati;
JOHN|9|33|nisi esset hic a Deo, non poterat facere quidquam ".
JOHN|9|34|Responderunt et dixerunt ei: " In peccatis tu natus es totus et tu doces nos? ". Et eiecerunt eum foras.
JOHN|9|35|Audivit Iesus quia eiecerunt eum foras et, cum invenisset eum, dixit ei: " Tu credis in Filium hominis? ".
JOHN|9|36|Respondit ille et dixit: " Et quis est, Domine, ut credam in eum? ".
JOHN|9|37|Dixit ei Iesus: " Et vidisti eum; et, qui loquitur tecum, ipse est ".
JOHN|9|38|At ille ait: " Credo, Domine! "; et adoravit eum.
JOHN|9|39|Et dixit Iesus: " In iudicium ego in hunc mundum veni, ut, qui non vident, videant, et, qui vident, caeci fiant ".
JOHN|9|40|Audierunt haec ex pharisaeis, qui cum ipso erant, et dixerunt ei: " Numquid et nos caeci sumus? ".
JOHN|9|41|Dixit eis Iesus: " Si caeci essetis, non haberetis peccatum. Nunc vero dicitis: "Videmus!"; peccatum vestrum manet ".
JOHN|10|1|" Amen, amen dico vobis: Qui non intrat per ostium in ovile ovium, sed ascendit aliunde, ille fur est et latro;
JOHN|10|2|qui autem intrat per ostium, pastor est ovium.
JOHN|10|3|Huic ostiarius aperit, et oves vocem eius audiunt, et proprias oves vocat nominatim et educit eas.
JOHN|10|4|Cum proprias omnes emiserit, ante eas vadit, et oves illum sequuntur, quia sciunt vocem eius;
JOHN|10|5|alienum autem non sequentur, sed fugient ab eo, quia non noverunt vocem alienorum ".
JOHN|10|6|Hoc proverbium dixit eis Iesus; illi autem non cognoverunt quid esset, quod loquebatur eis.
JOHN|10|7|Dixit ergo iterum Iesus: " Amen, amen dico vobis: Ego sum ostium ovium.
JOHN|10|8|Omnes, quotquot venerunt ante me, fures sunt et latrones, sed non audierunt eos oves.
JOHN|10|9|Ego sum ostium; per me, si quis introierit, salvabitur et ingredietur et egredietur et pascua inveniet.
JOHN|10|10|Fur non venit, nisi ut furetur et mactet et perdat; ego veni, ut vitam habeant et abundantius habeant.
JOHN|10|11|Ego sum pastor bonus; bonus pastor animam suam ponit pro ovibus;
JOHN|10|12|mercennarius et, qui non est pastor, cuius non sunt oves propriae, videt lupum venientem et dimittit oves et fugit - et lupus rapit eas et dispergit -
JOHN|10|13|quia mercennarius est et non pertinet ad eum de ovibus.
JOHN|10|14|Ego sum pastor bonus et cognosco meas, et cognoscunt me meae,
JOHN|10|15|sicut cognoscit me Pater, et ego cognosco Patrem; et animam meam pono pro ovibus.
JOHN|10|16|Et alias oves habeo, quae non sunt ex hoc ovili, et illas oportet me adducere, et vocem meam audient et fient unus grex, unus pastor.
JOHN|10|17|Propterea me Pater diligit, quia ego pono animam meam, ut iterum sumam eam.
JOHN|10|18|Nemo tollit eam a me, sed ego pono eam a meipso. Potestatem habeo ponendi eam et potestatem habeo iterum sumendi eam. Hoc mandatum accepi a Patre meo ".
JOHN|10|19|Dissensio iterum facta est inter Iudaeos propter sermones hos.
JOHN|10|20|Dicebant autem multi ex ipsis: " Daemonium habet et insanit! Quid eum auditis? ".
JOHN|10|21|Alii dicebant: " Haec verba non sunt daemonium habentis! Numquid daemonium potest caecorum oculos aperire? ".
JOHN|10|22|Facta sunt tunc Encaenia in Hierosolymis. Hiems erat;
JOHN|10|23|et ambulabat Iesus in templo in porticu Salomonis.
JOHN|10|24|Circumdederunt ergo eum Iudaei et dicebant ei: " Quousque animam nostram tollis? Si tu es Christus, dic nobis palam! ".
JOHN|10|25|Respondit eis Iesus: " Dixi vobis, et non creditis; opera, quae ego facio in nomine Patris mei, haec testimonium perhibent de me.
JOHN|10|26|Sed vos non creditis, quia non estis ex ovibus meis.
JOHN|10|27|Oves meae vocem meam audiunt, et ego cognosco eas, et sequuntur me;
JOHN|10|28|et ego vitam aeternam do eis, et non peribunt in aeternum, et non rapiet eas quisquam de manu mea.
JOHN|10|29|Pater meus quod dedit mihi, maius omnibus est, et nemo potest rapere de manu Patris.
JOHN|10|30|Ego et Pater unum sumus ".
JOHN|10|31|Sustulerunt iterum lapides Iudaei, ut lapidarent eum.
JOHN|10|32|Respondit eis Iesus: " Multa opera bona ostendi vobis ex Patre; propter quod eorum opus me lapidatis? ".
JOHN|10|33|Responderunt ei Iudaei: " De bono opere non lapidamus te sed de blasphemia, et quia tu, homo cum sis, facis teipsum Deum ".
JOHN|10|34|Respondit eis Iesus: " Nonne scriptum est in lege vestra: "Ego dixi: Dii estis?".
JOHN|10|35|Si illos dixit deos, ad quos sermo Dei factus est, et non potest solvi Scriptura,
JOHN|10|36|quem Pater sanctificavit et misit in mundum, vos dicitis: Blasphemas!", quia dixi: Filius Dei sum?
JOHN|10|37|Si non facio opera Patris mei, nolite credere mihi;
JOHN|10|38|si autem facio, et si mihi non vultis credere, operibus credite, ut cognoscatis et sciatis quia in me est Pater, et ego in Patre ".
JOHN|10|39|Quaerebant ergo iterum eum prehendere; et exivit de manibus eorum.
JOHN|10|40|Et abiit iterum trans Iordanem in eum locum, ubi erat Ioannes baptizans primum, et mansit illic.
JOHN|10|41|Et multi venerunt ad eum et dicebant: " Ioannes quidem signum fecit nullum; omnia autem, quaecumque dixit Ioannes de hoc, vera erant ".
JOHN|10|42|Et multi crediderunt in eum illic.
JOHN|11|1|Erat autem quidam lan guens Lazarus a Bethania, de castello Mariae et Marthae sororis eius.
JOHN|11|2|Maria autem erat, quae unxit Dominum unguento et extersit pedes eius capillis suis, cuius frater Lazarus infirmabatur.
JOHN|11|3|Miserunt ergo sorores ad eum dicentes: " Domine, ecce, quem amas, infirmatur ".
JOHN|11|4|Audiens autem Iesus dixit: " Infirmitas haec non est ad mortem sed pro gloria Dei, ut glorificetur Filius Dei per eam ".
JOHN|11|5|Diligebat autem Iesus Martham et sororem eius et Lazarum.
JOHN|11|6|Ut ergo audivit quia infirmabatur, tunc quidem mansit in loco, in quo erat, duobus diebus;
JOHN|11|7|deinde post hoc dicit discipulis: " Eamus in Iudaeam iterum ".
JOHN|11|8|Dicunt ei discipuli: " Rabbi, nunc quaerebant te Iudaei lapidare, et iterum vadis illuc? ".
JOHN|11|9|Respondit Iesus: " Nonne duodecim horae sunt diei? Si quis ambulaverit in die, non offendit, quia lucem huius mundi videt;
JOHN|11|10|si quis autem ambulaverit in nocte, offendit, quia lux non est in eo ".
JOHN|11|11|Haec ait et post hoc dicit eis: " Lazarus amicus noster dormit, sed vado, ut a somno exsuscitem eum ".
JOHN|11|12|Dixerunt ergo ei discipuli: " Domine, si dormit, salvus erit ".
JOHN|11|13|Dixerat autem Iesus de morte eius, illi autem putaverunt quia de dormitione somni diceret.
JOHN|11|14|Tunc ergo dixit eis Iesus manifeste: " Lazarus mortuus est,
JOHN|11|15|et gaudeo propter vos, ut credatis, quoniam non eram ibi; sed eamus ad eum ".
JOHN|11|16|Dixit ergo Thomas, qui dicitur Didymus, ad condiscipulos: " Eamus et nos, ut moriamur cum eo! ".
JOHN|11|17|Venit itaque Iesus et invenit eum quattuor dies iam in monumento habentem.
JOHN|11|18|Erat autem Bethania iuxta Hierosolymam quasi stadiis quindecim.
JOHN|11|19|Multi autem ex Iudaeis venerant ad Martham et Mariam, ut consolarentur eas de fratre.
JOHN|11|20|Martha ergo ut audivit quia Iesus venit, occurrit illi; Maria autem domi sedebat.
JOHN|11|21|Dixit ergo Martha ad Iesum: " Domine, si fuisses hic, frater meus non esset mortuus!
JOHN|11|22|Sed et nunc scio quia, quaecumque poposceris a Deo, dabit tibi Deus ".
JOHN|11|23|Dicit illi Iesus: " Resurget frater tuus ".
JOHN|11|24|Dicit ei Martha: " Scio quia resurget in resurrectione in novissimo die.
JOHN|11|25|Dixit ei Iesus: " Ego sum resurrectio et vita. Qui credit in me, etsi mortuus fuerit, vivet;
JOHN|11|26|et omnis, qui vivit et credit in me, non morietur in aeternum. Credis hoc? ".
JOHN|11|27|Ait illi: " Utique, Domine; ego credidi quia tu es Christus Filius Dei, qui in mundum venisti ".
JOHN|11|28|Et cum haec dixisset, abiit et vocavit Mariam sororem suam silentio dicens: " Magister adest et vocat te ".
JOHN|11|29|Illa autem ut audivit, surrexit cito et venit ad eum;
JOHN|11|30|nondum enim venerat Iesus in castellum, sed erat adhuc in illo loco, ubi occurrerat ei Martha.
JOHN|11|31|Iudaei igitur, qui erant cum ea in domo et consolabantur eam, cum vidissent Mariam quia cito surrexit et exiit, secuti sunt eam putantes: " Vadit ad monumentum, ut ploret ibi ".
JOHN|11|32|Maria ergo, cum venisset ubi erat Iesus, videns eum cecidit ad pedes eius dicens ei: " Domine, si fuisses hic, non esset mortuus frater meus!.
JOHN|11|33|Iesus ergo, ut vidit eam plorantem et Iudaeos, qui venerant cum ea, plorantes, fremuit spiritu et turbavit seipsum
JOHN|11|34|et dixit: " Ubi posuistis eum? ". Dicunt ei: " Domine, veni et vide ".
JOHN|11|35|Lacrimatus est Iesus.
JOHN|11|36|Dicebant ergo Iudaei: " Ecce quomodo amabat eum! ".
JOHN|11|37|Quidam autem dixerunt ex ipsis: " Non poterat hic, qui aperuit oculos caeci, facere, ut et hic non moreretur? ".
JOHN|11|38|Iesus ergo rursum fremens in semetipso, venit ad monumentum; erat autem spelunca, et lapis superpositus erat ei.
JOHN|11|39|Ait Iesus: " Tollite lapidem! ". Dicit ei Martha, soror eius, qui mortuus fuerat: " Domine, iam foetet; quatriduanus enim est! ".
JOHN|11|40|Dicit ei Iesus: " Nonne dixi tibi quoniam, si credideris, videbis gloriam Dei? ".
JOHN|11|41|Tulerunt ergo lapidem. Iesus autem, elevatis sursum oculis, dixit: " Pater, gratias ago tibi quoniam audisti me.
JOHN|11|42|Ego autem sciebam quia semper me audis, sed propter populum, qui circumstat, dixi, ut credant quia tu me misisti ".
JOHN|11|43|Et haec cum dixisset, voce magna clamavit: " Lazare, veni foras! ".
JOHN|11|44|Prodiit, qui fuerat mortuus, ligatus pedes et manus institis; et facies illius sudario erat ligata. Dicit Iesus eis: " Solvite eum et sinite eum abire ".
JOHN|11|45|Multi ergo ex Iudaeis, qui venerant ad Mariam et viderant, quae fecit, crediderunt in eum;
JOHN|11|46|quidam autem ex ipsis abierunt ad pharisaeos et dixerunt eis, quae fecit Iesus.
JOHN|11|47|Collegerunt ergo pontifices et pharisaei concilium et dicebant: " Quid facimus, quia hic homo multa signa facit?
JOHN|11|48|Si dimittimus eum sic, omnes credent in eum, et venient Romani et tollent nostrum et locum et gentem! ".
JOHN|11|49|Unus autem ex ipsis, Caiphas, cum esset pontifex anni illius, dixit eis: " Vos nescitis quidquam
JOHN|11|50|nec cogitatis quia expedit vobis, ut unus moriatur homo pro populo, et non tota gens pereat! ".
JOHN|11|51|Hoc autem a semetipso non dixit; sed, cum esset pontifex anni illius, prophetavit quia Iesus moriturus erat pro gente
JOHN|11|52|et non tantum pro gente, sed et ut filios Dei, qui erant dispersi, congregaret in unum.
JOHN|11|53|Ab illo ergo die cogitaverunt, ut interficerent eum.
JOHN|11|54|Iesus ergo iam non in palam ambulabat apud Iudaeos, sed abiit inde in regionem iuxta desertum, in civitatem, quae dicitur Ephraim, et ibi morabatur cum discipulis.
JOHN|11|55|Proximum autem erat Pascha Iudaeorum, et ascenderunt multi Hierosolymam de regione ante Pascha, ut sanctificarent seipsos.
JOHN|11|56|Quaerebant ergo Iesum et colloquebantur ad invicem in templo stantes: " Quid videtur vobis? Numquid veniet ad diem festum? ".
JOHN|11|57|Dederant autem pontifices et pharisaei mandatum, ut, si quis cognoverit, ubi sit, indicet, ut apprehendant eum.
JOHN|12|1|Iesus ergo ante sex dies Paschae venit Bethaniam, ubi erat Lazarus, quem suscitavit a mortuis Iesus.
JOHN|12|2|Fecerunt ergo ei cenam ibi, et Martha ministrabat, Lazarus vero unus erat ex discumbentibus cum eo.
JOHN|12|3|Maria ergo accepit libram unguenti nardi puri, pretiosi, et unxit pedes Iesu et extersit capillis suis pedes eius; domus autem impleta est ex odore unguenti.
JOHN|12|4|Dicit autem Iudas Iscariotes, unus ex discipulis eius, qui erat eum traditurus:
JOHN|12|5|" Quare hoc unguentum non veniit trecentis denariis et datum est egenis?.
JOHN|12|6|Dixit autem hoc, non quia de egenis pertinebat ad eum, sed quia fur erat et, loculos habens, ea, quae mittebantur, portabat.
JOHN|12|7|Dixit ergo Iesus: " Sine illam, ut in diem sepulturae meae servet illud.
JOHN|12|8|Pauperes enim semper habetis vobiscum, me autem non semper habetis ".
JOHN|12|9|Cognovit ergo turba multa ex Iudaeis quia illic est, et venerunt non propter Iesum tantum, sed ut et Lazarum viderent, quem suscitavit a mortuis.
JOHN|12|10|Cogitaverunt autem principes sacerdotum, ut et Lazarum interficerent,
JOHN|12|11|quia multi propter illum abibant ex Iudaeis et credebant in Iesum.
JOHN|12|12|In crastinum turba multa, quae venerat ad diem festum, cum audissent quia venit Iesus Hierosolymam,
JOHN|12|13|acceperunt ramos palmarum et processerunt obviam ei et clamabant: Hosanna!Benedictus, qui venit in nomine Domini, et rex Israel! ".
JOHN|12|14|Invenit autem Iesus asellum et sedit super eum, sicut scriptum est:
JOHN|12|15|" Noli timere, filia Sion.Ecce rex tuus venitsedens super pullum asinae ".
JOHN|12|16|Haec non cognoverunt discipuli eius primum, sed quando glorificatus est Iesus, tunc recordati sunt quia haec erant scripta de eo, et haec fecerunt ei.
JOHN|12|17|Testimonium ergo perhibebat turba, quae erat cum eo, quando Lazarum vocavit de monumento et suscitavit eum a mortuis.
JOHN|12|18|Propterea et obviam venit ei turba, quia audierunt eum fecisse hoc signum.
JOHN|12|19|Pharisaei ergo dixerunt ad semetipsos: " Videtis quia nihil proficitis? Ecce mundus post eum abiit! ".
JOHN|12|20|Erant autem Graeci quidam ex his, qui ascenderant, ut adorarent in die festo;
JOHN|12|21|hi ergo accesserunt ad Philippum, qui erat a Bethsaida Galilaeae, et rogabant eum dicentes: " Domine, volumus Iesum videre ".
JOHN|12|22|Venit Philippus et dicit Andreae; venit Andreas et Philippus et dicunt Iesu.
JOHN|12|23|Iesus autem respondet eis dicens: " Venit hora, ut glorificetur Filius hominis.
JOHN|12|24|Amen, amen dico vobis: Nisi granum frumenti cadens in terram mortuum fuerit, ipsum solum manet; si autem mortuum fuerit, multum fructum affert.
JOHN|12|25|Qui amat animam suam, perdit eam; et, qui odit animam suam in hoc mundo, in vitam aeternam custodiet eam.
JOHN|12|26|Si quis mihi ministrat, me sequatur, et ubi sum ego, illic et minister meus erit; si quis mihi ministraverit, honorificabit eum Pater.
JOHN|12|27|Nunc anima mea turbata est. Et quid dicam? Pater, salvifica me ex hora hac? Sed propterea veni in horam hanc.
JOHN|12|28|Pater, glorifica tuum nomen! ". Venit ergo vox de caelo: " Et glorificavi et iterum glorificabo ".
JOHN|12|29|Turba ergo, quae stabat et audierat, dicebat tonitruum factum esse; alii dicebant: " Angelus ei locutus est ".
JOHN|12|30|Respondit Iesus et dixit: " Non propter me vox haec facta est sed propter vos.
JOHN|12|31|Nunc iudicium est huius mundi, nunc princeps huius mundi eicietur foras;
JOHN|12|32|et ego, si exaltatus fuero a terra, omnes traham ad meipsum ".
JOHN|12|33|Hoc autem dicebat significans, qua morte esset moriturus.
JOHN|12|34|Respondit ergo ei turba: " Nos audivimus ex Lege, quia Christus manet in aeternum; et quomodo tu dicis: "Oportet exaltari Filium hominis"? Quis est iste Filius hominis? ".
JOHN|12|35|Dixit ergo eis Iesus: " Adhuc modicum tempus lumen in vobis est. Ambulate, dum lucem habetis, ut non tenebrae vos comprehendant; et, qui ambulat in tenebris, nescit quo vadat.
JOHN|12|36|Dum lucem habetis, credite in lucem, ut filii lucis fiatis ". Haec locutus est Iesus et abiit et abscondit se ab eis.
JOHN|12|37|Cum autem tanta signa fecisset coram eis, non credebant in eum,
JOHN|12|38|ut sermo Isaiae prophetae impleretur, quem dixit: Domine, quis credidit auditui nostro,et brachium Domini cui revelatum est? ".
JOHN|12|39|Propterea non poterant credere, quia iterum dixit Isaias:
JOHN|12|40|" Excaecavit oculos eorumet induravit eorum cor,ut non videant oculiset intellegant corde et convertantur,et sanem eos ".
JOHN|12|41|Haec dixit Isaias, quia vidit gloriam eius et locutus est de eo.
JOHN|12|42|Verumtamen et ex principibus multi crediderunt in eum, sed propter pharisaeos non confitebantur, ut de synagoga non eicerentur;
JOHN|12|43|dilexerunt enim gloriam hominum magis quam gloriam Dei.
JOHN|12|44|Iesus autem clamavit et dixit: " Qui credit in me, non credit in me sed in eum, qui misit me;
JOHN|12|45|et, qui videt me, videt eum, qui misit me.
JOHN|12|46|Ego lux in mundum veni, ut omnis, qui credit in me, in tenebris non maneat.
JOHN|12|47|Et si quis audierit verba mea et non custodierit, ego non iudico eum; non enim veni, ut iudicem mundum, sed ut salvificem mundum.
JOHN|12|48|Qui spernit me et non accipit verba mea, habet, qui iudicet eum: sermo, quem locutus sum, ille iudicabit eum in novissimo die,
JOHN|12|49|quia ego ex meipso non sum locutus, sed, qui misit me, Pater, ipse mihi mandatum dedit quid dicam et quid loquar.
JOHN|12|50|Et scio quia mandatum eius vita aeterna est. Quae ergo ego loquor, sicut dixit mihi Pater, sic loquor ".
JOHN|13|1|Ante diem autem festum Pa schae, sciens Iesus quia venit eius hora, ut transeat ex hoc mundo ad Patrem, cum dilexisset suos, qui erant in mundo, in finem dilexit eos.
JOHN|13|2|Et in cena, cum Diabolus iam misisset in corde, ut traderet eum Iudas Simonis Iscariotis,
JOHN|13|3|sciens quia omnia dedit ei Pater in manus, et quia a Deo exivit et ad Deum vadit,
JOHN|13|4|surgit a cena et ponit vestimenta sua et, cum accepisset linteum, praecinxit se.
JOHN|13|5|Deinde mittit aquam in pelvem et coepit lavare pedes discipulorum et extergere linteo, quo erat praecinctus.
JOHN|13|6|Venit ergo ad Simonem Petrum. Dicit ei: " Domine, tu mihi lavas pedes?.
JOHN|13|7|Respondit Iesus et dixit ei: " Quod ego facio, tu nescis modo, scies autem postea ".
JOHN|13|8|Dicit ei Petrus: " Non lavabis mihi pedes in aeternum! ". Respondit Iesus ei: " Si non lavero te, non habes partem mecum ".
JOHN|13|9|Dicit ei Simon Petrus: " Domine, non tantum pedes meos sed et manus et caput! ".
JOHN|13|10|Dicit ei Iesus: " Qui lotus est, non indiget nisi ut pedes lavet, sed est mundus totus; et vos mundi estis sed non omnes ".
JOHN|13|11|Sciebat enim quisnam esset, qui traderet eum; propterea dixit: " Non estis mundi omnes ".
JOHN|13|12|Postquam ergo lavit pedes eorum et accepit vestimenta sua, cum recubuisset iterum, dixit eis: " Scitis quid fecerim vobis?
JOHN|13|13|Vos vocatis me: "Magister" et: "Domine", et bene dicitis; sum etenim.
JOHN|13|14|Si ergo ego lavi vestros pedes, Dominus et Magister, et vos debetis alter alterius lavare pedes.
JOHN|13|15|Exemplum enim dedi vobis, ut, quemadmodum ego feci vobis, et vos faciatis.
JOHN|13|16|Amen, amen dico vobis: Non est servus maior domino suo, neque apostolus maior eo, qui misit illum.
JOHN|13|17|Si haec scitis, beati estis, si facitis ea.
JOHN|13|18|Non de omnibus vobis dico, ego scio, quos elegerim, sed ut impleatur Scriptura: "Qui manducat meum panem, levavit contra me calcaneum suum".
JOHN|13|19|Amodo dico vobis priusquam fiat, ut credatis, cum factum fuerit, quia ego sum.
JOHN|13|20|Amen, amen dico vobis: Qui accipit, si quem misero, me accipit; qui autem me accipit, accipit eum, qui me misit ".
JOHN|13|21|Cum haec dixisset Iesus, turbatus est spiritu et protestatus est et dixit: " Amen, amen dico vobis: Unus ex vobis tradet me ".
JOHN|13|22|Aspiciebant ad invicem discipuli, haesitantes de quo diceret.
JOHN|13|23|Erat recumbens unus ex discipulis eius in sinu Iesu, quem diligebat Iesus.
JOHN|13|24|Innuit ergo huic Simon Petrus, ut interrogaret: " Quis est, de quo dicit? ".
JOHN|13|25|Cum ergo recumberet ille ita supra pectus Iesu, dicit ei: " Domine, quis est? ".
JOHN|13|26|Respondet Iesus: " Ille est, cui ego intinctam buccellam porrexero ". Cum ergo intinxisset buccellam, dat Iudae Simonis Iscariotis.
JOHN|13|27|Et post buccellam tunc introivit in illum Satanas. Dicit ergo ei Iesus: Quod facis, fac citius ".
JOHN|13|28|Hoc autem nemo scivit discumbentium ad quid dixerit ei;
JOHN|13|29|quidam enim putabant quia loculos habebat Iudas, quia dicit ei Iesus: " Eme ea, quae opus sunt nobis ad diem festum ", aut egenis ut aliquid daret.
JOHN|13|30|Cum ergo accepisset ille buccellam, exivit continuo; erat autem nox.
JOHN|13|31|Cum ergo exisset, dicit Iesus: " Nunc clarificatus est Filius hominis, et Deus clarificatus est in eo;
JOHN|13|32|si Deus clarificatus est in eo, et Deus clarificabit eum in semetipso et continuo clarificabit eum.
JOHN|13|33|Filioli, adhuc modicum vobiscum sum; quaeretis me, et sicut dixi Iudaeis: Quo ego vado, vos non potestis venire, et vobis dico modo.
JOHN|13|34|Mandatum novum do vobis, ut diligatis invicem; sicut dilexi vos, ut et vos diligatis invicem.
JOHN|13|35|In hoc cognoscent omnes quia mei discipuli estis: si dilectionem habueritis ad invicem ".
JOHN|13|36|Dicit ei Simon Petrus: " Domine, quo vadis? ". Respondit Iesus: " Quo vado, non potes me modo sequi, sequeris autem postea ".
JOHN|13|37|Dicit ei Petrus: " Domine, quare non possum te sequi modo? Animam meam pro te ponam ".
JOHN|13|38|Respondet Iesus: " Animam tuam pro me pones? Amen, amen dico tibi: Non cantabit gallus, donec me ter neges.
JOHN|14|1|Non turbetur cor vestrum. Creditis in Deum et in me credite.
JOHN|14|2|In domo Patris mei mansiones multae sunt; si quo minus, dixissem vobis, quia vado parare vobis locum?
JOHN|14|3|Et si abiero et praeparavero vobis locum, iterum venio et accipiam vos ad meipsum, ut, ubi sum ego, et vos sitis.
JOHN|14|4|Et quo ego vado, scitis viam ".
JOHN|14|5|Dicit ei Thomas: " Domine, nescimus quo vadis; quomodo possumus viam scire? ".
JOHN|14|6|Dicit ei Iesus: " Ego sum via et veritas et vita; nemo venit ad Patrem nisi per me.
JOHN|14|7|Si cognovistis me, et Patrem meum utique cognoscetis; et amodo cognoscitis eum et vidistis eum ".
JOHN|14|8|Dicit ei Philippus: " Domine, ostende nobis Patrem, et sufficit nobis ".
JOHN|14|9|Dicit ei Iesus: " Tanto tempore vobiscum sum, et non cognovisti me, Philippe? Qui vidit me, vidit Patrem. Quomodo tu dicis: "Ostende nobis Patrem"?
JOHN|14|10|Non credis quia ego in Patre, et Pater in me est? Verba, quae ego loquor vobis, a meipso non loquor; Pater autem in me manens facit opera sua.
JOHN|14|11|Credite mihi quia ego in Patre, et Pater in me est; alioquin propter opera ipsa credite.
JOHN|14|12|Amen, amen dico vobis: Qui credit in me, opera, quae ego facio, et ipse faciet et maiora horum faciet, quia ego ad Patrem vado.
JOHN|14|13|Et quodcumque petieritis in nomine meo, hoc faciam, ut glorificetur Pater in Filio;
JOHN|14|14|si quid petieritis me in nomine meo, ego faciam.
JOHN|14|15|Si diligitis me, mandata mea servabitis;
JOHN|14|16|et ego rogabo Patrem, et alium Paraclitum dabit vobis, ut maneat vobiscum in aeternum,
JOHN|14|17|Spiritum veritatis, quem mundus non potest accipere, quia non videt eum nec cognoscit. Vos cognoscitis eum, quia apud vos manet; et in vobis erit.
JOHN|14|18|Non relinquam vos orphanos; venio ad vos.
JOHN|14|19|Adhuc modicum, et mundus me iam non videt; vos autem videtis me, quia ego vivo et vos vivetis.
JOHN|14|20|In illo die vos cognoscetis quia ego sum in Patre meo, et vos in me, et ego in vobis.
JOHN|14|21|Qui habet mandata mea et servat ea, ille est, qui diligit me; qui autem diligit me, diligetur a Patre meo, et ego diligam eum et manifestabo ei meipsum ".
JOHN|14|22|Dicit ei Iudas, non ille Iscariotes: " Domine, et quid factum est, quia nobis manifestaturus es teipsum et non mundo? ".
JOHN|14|23|Respondit Iesus et dixit ei: " Si quis diligit me, sermonem meum servabit, et Pater meus diliget eum, et ad eum veniemus et mansionem apud eum faciemus;
JOHN|14|24|qui non diligit me, sermones meos non servat. Et sermo, quem auditis, non est meus, sed eius qui misit me, Patris.
JOHN|14|25|Haec locutus sum vobis apud vos manens.
JOHN|14|26|Paraclitus autem, Spiritus Sanctus, quem mittet Pater in nomine meo, ille vos docebit omnia et suggeret vobis omnia, quae dixi vobis.
JOHN|14|27|Pacem relinquo vobis, pacem meam do vobis; non quomodo mundus dat, ego do vobis. Non turbetur cor vestrum neque formidet.
JOHN|14|28|Audistis quia ego dixi vobis: Vado et venio ad vos. Si diligeretis me, gauderetis quia vado ad Patrem, quia Pater maior me est.
JOHN|14|29|Et nunc dixi vobis, priusquam fiat, ut, cum factum fuerit, credatis.
JOHN|14|30|Iam non multa loquar vobiscum, venit enim princeps mundi et in me non habet quidquam;
JOHN|14|31|sed, ut cognoscat mundus quia diligo Patrem, et sicut mandatum dedit mihi Pater, sic facio. Surgite, eamus hinc.
JOHN|15|1|Ego sum vitis vera, et Pater meus agricola est.
JOHN|15|2|Omnem palmitem in me non ferentem fructum tollit eum; et omnem, qui fert fructum, purgat eum, ut fructum plus afferat.
JOHN|15|3|Iam vos mundi estis propter sermonem, quem locutus sum vobis.
JOHN|15|4|Manete in me, et ego in vobis. Sicut palmes non potest ferre fructum a semetipso, nisi manserit in vite, sic nec vos, nisi in me manseritis.
JOHN|15|5|Ego sum vitis, vos palmites. Qui manet in me, et ego in eo, hic fert fructum multum, quia sine me nihil potestis facere.
JOHN|15|6|Si quis in me non manserit, missus est foras sicut palmes et aruit; et colligunt eos et in ignem mittunt, et ardent.
JOHN|15|7|Si manseritis in me, et verba mea in vobis manserint, quodcumque volueritis, petite, et fiet vobis.
JOHN|15|8|In hoc clarificatus est Pater meus, ut fructum multum afferatis et efficiamini mei discipuli.
JOHN|15|9|Sicut dilexit me Pater, et ego dilexi vos; manete in dilectione mea.
JOHN|15|10|Si praecepta mea servaveritis, manebitis in dilectione mea, sicut ego Patris mei praecepta servavi et maneo in eius dilectione.
JOHN|15|11|Haec locutus sum vobis, ut gaudium meum in vobis sit, et gaudium vestrum impleatur.
JOHN|15|12|Hoc est praeceptum meum, ut diligatis invicem, sicut dilexi vos;
JOHN|15|13|maiorem hac dilectionem nemo habet, ut animam suam quis ponat pro amicis suis.
JOHN|15|14|Vos amici mei estis, si feceritis, quae ego praecipio vobis.
JOHN|15|15|Iam non dico vos servos, quia servus nescit quid facit dominus eius; vos autem dixi amicos, quia omnia, quae audivi a Patre meo, nota feci vobis.
JOHN|15|16|Non vos me elegistis, sed ego elegi vos et posui vos, ut vos eatis et fructum afferatis, et fructus vester maneat, ut quodcumque petieritis Patrem in nomine meo, det vobis.
JOHN|15|17|Haec mando vobis, ut diligatis invicem.
JOHN|15|18|Si mundus vos odit, scitote quia me priorem vobis odio habuit.
JOHN|15|19|Si de mundo essetis, mundus, quod suum est, diligeret; quia vero de mundo non estis, sed ego elegi vos de mundo, propterea odit vos mundus.
JOHN|15|20|Mementote sermonis, quem ego dixi vobis: Non est servus maior domino suo. Si me persecuti sunt, et vos persequentur; si sermonem meum servaverunt, et vestrum servabunt.
JOHN|15|21|Sed haec omnia facient vobis propter nomen meum, quia nesciunt eum, qui misit me.
JOHN|15|22|Si non venissem et locutus fuissem eis, peccatum non haberent; nunc autem excusationem non habent de peccato suo.
JOHN|15|23|Qui me odit et Patrem meum odit.
JOHN|15|24|Si opera non fecissem in eis, quae nemo alius fecit, peccatum non haberent; nunc autem et viderunt et oderunt et me et Patrem meum.
JOHN|15|25|Sed ut impleatur sermo, qui in lege eorum scriptus est: "Odio me habuerunt gratis".
JOHN|15|26|Cum autem venerit Paraclitus, quem ego mittam vobis a Patre, Spiritum veritatis, qui a Patre procedit, ille testimonium perhibebit de me;
JOHN|15|27|sed et vos testimonium perhibetis, quia ab initio mecum estis.
JOHN|16|1|Haec locutus sum vobis, ut non scandalizemini.
JOHN|16|2|Absque synagogis facient vos; sed venit hora, ut omnis, qui interficit vos, arbitretur obsequium se praestare Deo.
JOHN|16|3|Et haec facient, quia non noverunt Patrem neque me.
JOHN|16|4|Sed haec locutus sum vobis, ut, cum venerit hora eorum, reminiscamini eorum, quia ego dixi vobis. Haec autem vobis ab initio non dixi, quia vobiscum eram.
JOHN|16|5|At nunc vado ad eum, qui me misit, et nemo ex vobis interrogat me: "Quo vadis?".
JOHN|16|6|Sed quia haec locutus sum vobis, tristitia implevit cor vestrum.
JOHN|16|7|Sed ego veritatem dico vobis: Expedit vobis, ut ego vadam. Si enim non abiero, Paraclitus non veniet ad vos; si autem abiero, mittam eum ad vos.
JOHN|16|8|Et cum venerit ille, arguet mundum de peccato et de iustitia et de iudicio:
JOHN|16|9|de peccato quidem, quia non credunt in me;
JOHN|16|10|de iustitia vero, quia ad Patrem vado, et iam non videtis me;
JOHN|16|11|de iudicio autem, quia princeps mundi huius iudicatus est.
JOHN|16|12|Adhuc multa habeo vobis dicere, sed non potestis portare modo.
JOHN|16|13|Cum autem venerit ille, Spiritus veritatis, deducet vos in omnem veritatem; non enim loquetur a semetipso, sed quaecumque audiet, loquetur et, quae ventura sunt, annuntiabit vobis.
JOHN|16|14|Ille me clarificabit, quia de meo accipiet et annuntiabit vobis.
JOHN|16|15|Omnia, quaecumque habet Pater, mea sunt; propterea dixi quia de meo accipit et annuntiabit vobis.
JOHN|16|16|Modicum, et iam non videtis me; et iterum modicum, et videbitis me ".
JOHN|16|17|Dixerunt ergo ex discipulis eius ad invicem: " Quid est hoc, quod dicit nobis: "Modicum, et non videtis me; et iterum modicum, et videbitis me" et: "Vado ad Patrem"? ".
JOHN|16|18|Dicebant ergo: " Quid est hoc, quod dicit: "Modicum"? Nescimus quid loquitur ".
JOHN|16|19|Cognovit Iesus quia volebant eum interrogare et dixit eis: " De hoc quaeritis inter vos, quia dixi: "Modicum, et non videtis me; et iterum modicum, et videbitis me"?
JOHN|16|20|Amen, amen dico vobis quia plorabitis et flebitis vos, mundus autem gaudebit; vos contristabimini, sed tristitia vestra vertetur in gaudium.
JOHN|16|21|Mulier, cum parit, tristitiam habet, quia venit hora eius; cum autem pepererit puerum, iam non meminit pressurae propter gaudium, quia natus est homo in mundum.
JOHN|16|22|Et vos igitur nunc quidem tristitiam habetis; iterum autem videbo vos, et gaudebit cor vestrum, et gaudium vestrum nemo tollit a vobis.
JOHN|16|23|Et in illo die me non rogabitis quidquam.Amen, amen dico vobis: Si quid petieritis Patrem in nomine meo, dabit vobis.
JOHN|16|24|Usque modo non petistis quidquam in nomine meo. Petite et accipietis, ut gaudium vestrum sit plenum.
JOHN|16|25|Haec in proverbiis locutus sum vobis; venit hora, cum iam non in proverbiis loquar vobis, sed palam de Patre annuntiabo vobis.
JOHN|16|26|Illo die in nomine meo petetis, et non dico vobis quia ego rogabo Patrem de vobis;
JOHN|16|27|ipse enim Pater amat vos, quia vos me amastis et credidistis quia ego a Deo exivi.
JOHN|16|28|Exivi a Patre et veni in mundum; iterum relinquo mundum et vado ad Patrem ".
JOHN|16|29|Dicunt discipuli eius: " Ecce nunc palam loqueris, et proverbium nullum dicis.
JOHN|16|30|Nunc scimus quia scis omnia, et non opus est tibi, ut quis te interroget; in hoc credimus quia a Deo existi ".
JOHN|16|31|Respondit eis Iesus: " Modo creditis?
JOHN|16|32|Ecce venit hora et iam venit, ut dispergamini unusquisque in propria et me solum relinquatis; et non sum solus, quia Pater mecum est.
JOHN|16|33|Haec locutus sum vobis, ut in me pacem habeatis; in mundo pressuram habetis, sed confidite, ego vici mundum ".
JOHN|17|1|Haec locutus est Iesus; et, sublevatis oculis suis in cae lum, dixit: " Pater, venit hora: clarifica Filium tuum, ut Filius clarificet te,
JOHN|17|2|sicut dedisti ei potestatem omnis carnis, ut omne, quod dedisti ei, det eis vitam aeternam.
JOHN|17|3|Haec est autem vita aeterna, ut cognoscant te solum verum Deum et, quem misisti, Iesum Christum.
JOHN|17|4|Ego te clarificavi super terram; opus consummavi, quod dedisti mihi, ut faciam;
JOHN|17|5|et nunc clarifica me tu, Pater, apud temetipsum claritate, quam habebam, priusquam mundus esset, apud te.
JOHN|17|6|Manifestavi nomen tuum hominibus, quos dedisti mihi de mundo. Tui erant, et mihi eos dedisti, et sermonem tuum servaverunt.
JOHN|17|7|Nunc cognoverunt quia omnia, quae dedisti mihi, abs te sunt,
JOHN|17|8|quia verba, quae dedisti mihi, dedi eis; et ipsi acceperunt et cognoverunt vere quia a te exivi et crediderunt quia tu me misisti.
JOHN|17|9|Ego pro eis rogo; non pro mundo rogo, sed pro his, quos dedisti mihi, quia tui sunt;
JOHN|17|10|et mea omnia tua sunt, et tua mea; et clarificatus sum in eis.
JOHN|17|11|Et iam non sum in mundo, et hi in mundo sunt, et ego ad te venio.Pater sancte, serva eos in nomine tuo, quod dedisti mihi, ut sint unum sicut nos.
JOHN|17|12|Cum essem cum eis, ego servabam eos in nomine tuo, quod dedisti mihi, et custodivi, et nemo ex his periit, nisi filius perditionis, ut Scriptura impleatur.
JOHN|17|13|Nunc autem ad te venio et haec loquor in mundo, ut habeant gaudium meum impletum in semetipsis.
JOHN|17|14|Ego dedi eis sermonem tuum, et mundus odio eos habuit, quia non sunt de mundo, sicut ego non sum de mundo.
JOHN|17|15|Non rogo, ut tollas eos de mundo, sed ut serves eos ex Malo.
JOHN|17|16|De mundo non sunt, sicut ego non sum de mundo.
JOHN|17|17|Sanctifica eos in veritate; sermo tuus veritas est.
JOHN|17|18|Sicut me misisti in mundum, et ego misi eos in mundum;
JOHN|17|19|et pro eis ego sanctifico meipsum, ut sint et ipsi sanctificati in veritate.
JOHN|17|20|Non pro his autem rogo tantum, sed et pro eis, qui credituri sunt per verbum eorum in me,
JOHN|17|21|ut omnes unum sint, sicut tu, Pater, in me et ego in te, ut et ipsi in nobis unum sint; ut mundus credat quia tu me misisti.
JOHN|17|22|Et ego claritatem, quam dedisti mihi, dedi illis, ut sint unum, sicut nos unum sumus;
JOHN|17|23|ego in eis, et tu in me, ut sint consummati in unum; ut cognoscat mundus, quia tu me misisti et dilexisti eos, sicut me dilexisti.
JOHN|17|24|Pater, quod dedisti mihi, volo, ut ubi ego sum, et illi sint mecum, ut videant claritatem meam, quam dedisti mihi, quia dilexisti me ante constitutionem mundi.
JOHN|17|25|Pater iuste, et mundus te non cognovit; ego autem te cognovi, et hi cognoverunt quia tu me misisti;
JOHN|17|26|et notum feci eis nomen tuum et notum faciam, ut dilectio, qua dilexisti me, in ipsis sit, et ego in ipsis ".
JOHN|18|1|Haec cum dixisset Iesus, egressus est cum discipulis suis trans torrentem Cedron, ubi erat hortus, in quem introivit ipse et discipuli eius.
JOHN|18|2|Sciebat autem et Iudas, qui tradebat eum, locum, quia frequenter Iesus convenerat illuc cum discipulis suis.
JOHN|18|3|Iudas ergo, cum accepisset cohortem et a pontificibus et pharisaeis ministros, venit illuc cum lanternis et facibus et armis.
JOHN|18|4|Iesus itaque sciens omnia, quae ventura erant super eum, processit et dicit eis: " Quem quaeritis? ".
JOHN|18|5|Responderunt ei: " Iesum Nazarenum ". Dicit eis: " Ego sum! ". Stabat autem et Iudas, qui tradebat eum, cum ipsis.
JOHN|18|6|Ut ergo dixit eis: " Ego sum! ", abierunt retrorsum et ceciderunt in terram.
JOHN|18|7|Iterum ergo eos interrogavit: " Quem quaeritis? ". Illi autem dixerunt: Iesum Nazarenum ".
JOHN|18|8|Respondit Iesus: " Dixi vobis: Ego sum! Si ergo me quaeritis, sinite hos abire ",
JOHN|18|9|ut impleretur sermo, quem dixit: " Quos dedisti mihi, non perdidi ex ipsis quemquam ".
JOHN|18|10|Simon ergo Petrus, habens gladium, eduxit eum et percussit pontificis servum et abscidit eius auriculam dextram. Erat autem nomen servo Malchus.
JOHN|18|11|Dixit ergo Iesus Petro: " Mitte gladium in vaginam; calicem, quem dedit mihi Pater, non bibam illum? ".
JOHN|18|12|Cohors ergo et tribunus et ministri Iudaeorum comprehenderunt Iesum et ligaverunt eum
JOHN|18|13|et adduxerunt ad Annam primum; erat enim socer Caiphae, qui erat pontifex anni illius.
JOHN|18|14|Erat autem Caiphas, qui consilium dederat Iudaeis: " Expedit unum hominem mori pro populo ".
JOHN|18|15|Sequebatur autem Iesum Simon Petrus et alius discipulus. Discipulus autem ille erat notus pontifici et introivit cum Iesu in atrium pontificis;
JOHN|18|16|Petrus autem stabat ad ostium foris. Exivit ergo discipulus alius, qui erat notus pontifici, et dixit ostiariae et introduxit Petrum.
JOHN|18|17|Dicit ergo Petro ancilla ostiaria: " Numquid et tu ex discipulis es hominis istius? ". Dicit ille: " Non sum! ".
JOHN|18|18|Stabant autem servi et ministri, qui prunas fecerant, quia frigus erat, et calefaciebant se; erat autem cum eis et Petrus stans et calefaciens se.
JOHN|18|19|Pontifex ergo interrogavit Iesum de discipulis suis et de doctrina eius.
JOHN|18|20|Respondit ei Iesus: " Ego palam locutus sum mundo; ego semper docui in synagoga et in templo, quo omnes Iudaei conveniunt, et in occulto locutus sum nihil.
JOHN|18|21|Quid me interrogas? Interroga eos, qui audierunt quid locutus sum ipsis; ecce hi sciunt, quae dixerim ego ".
JOHN|18|22|Haec autem cum dixisset, unus assistens ministrorum dedit alapam Iesu dicens: " Sic respondes pontifici? ".
JOHN|18|23|Respondit ei Iesus: " Si male locutus sum, testimonium perhibe de malo; si autem bene, quid me caedis? ".
JOHN|18|24|Misit ergo eum Annas ligatum ad Caipham pontificem.
JOHN|18|25|Erat autem Simon Petrus stans et calefaciens se. Dixerunt ergo ei: " Numquid et tu ex discipulis eius es? ". Negavit ille et dixit: " Non sum!.
JOHN|18|26|Dicit unus ex servis pontificis, cognatus eius, cuius abscidit Petrus auriculam: " Nonne ego te vidi in horto cum illo? ".
JOHN|18|27|Iterum ergo negavit Petrus; et statim gallus cantavit.
JOHN|18|28|Adducunt ergo Iesum a Caipha in praetorium. Erat autem mane. Et ipsi non introierunt in praetorium, ut non contaminarentur, sed manducarent Pascha.
JOHN|18|29|Exivit ergo Pilatus ad eos foras et dicit: " Quam accusationem affertis adversus hominem hunc? ".
JOHN|18|30|Responderunt et dixerunt ei: " Si non esset hic malefactor, non tibi tradidissemus eum ".
JOHN|18|31|Dixit ergo eis Pilatus: " Accipite eum vos et secundum legem vestram iudicate eum! ". Dixerunt ei Iudaei: " Nobis non licet interficere quemquam ",
JOHN|18|32|ut sermo Iesu impleretur, quem dixit, significans qua esset morte moriturus.
JOHN|18|33|Introivit ergo iterum in praetorium Pilatus et vocavit Iesum et dixit ei: " Tu es rex Iudaeorum? ".
JOHN|18|34|Respondit Iesus: " A temetipso tu hoc dicis, an alii tibi dixerunt de me? ".
JOHN|18|35|Respondit Pilatus: " Numquid ego Iudaeus sum? Gens tua et pontifices tradiderunt te mihi; quid fecisti? ".
JOHN|18|36|Respondit Iesus: " Regnum meum non est de mundo hoc; si ex hoc mundo esset regnum meum, ministri mei decertarent, ut non traderer Iudaeis; nunc autem meum regnum non est hinc ".
JOHN|18|37|Dixit itaque ei Pilatus: " Ergo rex es tu? ". Respondit Iesus: " Tu dicis quia rex sum. Ego in hoc natus sum et ad hoc veni in mundum, ut testimonium perhibeam veritati; omnis, qui est ex veritate, audit meam vocem ".
JOHN|18|38|Dicit ei Pilatus: " Quid est veritas? ". Et cum hoc dixisset, iterum exivit ad Iudaeos et dicit eis: " Ego nullam invenio in eo causam.
JOHN|18|39|Est autem consuetudo vobis, ut unum dimittam vobis in Pascha; vultis ergo dimittam vobis regem Iudaeorum? ".
JOHN|18|40|Clamaverunt ergo rursum dicentes: " Non hunc sed Barabbam! ". Erat autem Barabbas latro.
JOHN|19|1|Tunc ergo apprehendit Pi latus Iesum et flagellavit.
JOHN|19|2|Et milites, plectentes coronam de spinis, imposuerunt capiti eius et veste purpurea circumdederunt eum;
JOHN|19|3|et veniebant ad eum et dicebant: " Ave, rex Iudaeorum! ", et dabant ei alapas.
JOHN|19|4|Et exiit iterum Pilatus foras et dicit eis: " Ecce adduco vobis eum foras, ut cognoscatis quia in eo invenio causam nullam ".
JOHN|19|5|Exiit ergo Iesus foras, portans spineam coronam et purpureum vestimentum. Et dicit eis: " Ecce homo! ".
JOHN|19|6|Cum ergo vidissent eum pontifices et ministri, clamaverunt dicentes: " Crucifige, crucifige! ". Dicit eis Pilatus: " Accipite eum vos et crucifigite; ego enim non invenio in eo causam ".
JOHN|19|7|Responderunt ei Iudaei: " Nos legem habemus, et secundum legem debet mori, quia Filium Dei se fecit ".
JOHN|19|8|Cum ergo audisset Pilatus hunc sermonem, magis timuit
JOHN|19|9|et ingressus est praetorium iterum et dicit ad Iesum: " Unde es tu? ". Iesus autem responsum non dedit ei.
JOHN|19|10|Dicit ergo ei Pilatus: " Mihi non loqueris? Nescis quia potestatem habeo dimittere te et potestatem habeo crucifigere te? ".
JOHN|19|11|Respondit Iesus: " Non haberes potestatem adversum me ullam, nisi tibi esset datum desuper; propterea, qui tradidit me tibi, maius peccatum habet.
JOHN|19|12|Exinde quaerebat Pilatus dimittere eum; Iudaei autem clamabant dicentes: " Si hunc dimittis, non es amicus Caesaris! Omnis, qui se regem facit, contradicit Caesari ".
JOHN|19|13|Pilatus ergo, cum audisset hos sermones, adduxit foras Iesum et sedit pro tribunali in locum, qui dicitur Lithostrotos, Hebraice autem Gabbatha.
JOHN|19|14|Erat autem Parasceve Paschae, hora erat quasi sexta. Et dicit Iudaeis: Ecce rex vester! ".
JOHN|19|15|Clamaverunt ergo illi: " Tolle, tolle, crucifige eum! ". Dicit eis Pilatus: " Regem vestrum crucifigam? ". Responderunt pontifices: " Non habemus regem, nisi Caesarem ".
JOHN|19|16|Tunc ergo tradidit eis illum, ut crucifigeretur. Susceperunt ergo Iesum.
JOHN|19|17|Et baiulans sibi crucem exivit in eum, qui dicitur Calvariae locum, quod Hebraice dicitur Golgotha,
JOHN|19|18|ubi eum crucifixerunt et cum eo alios duos hinc et hinc, medium autem Iesum.
JOHN|19|19|Scripsit autem et titulum Pilatus et posuit super crucem; erat autem scriptum: " Iesus Nazarenus Rex Iudaeorum ".
JOHN|19|20|Hunc ergo titulum multi legerunt Iudaeorum, quia prope civitatem erat locus, ubi crucifixus est Iesus; et erat scriptum Hebraice, Latine, Graece.
JOHN|19|21|Dicebant ergo Pilato pontifices Iudaeorum: " Noli scribere: Rex Iudaeorum, sed: Ipse dixit: "Rex sum Iudaeorum" ".
JOHN|19|22|Respondit Pilatus: " Quod scripsi, scripsi! ".
JOHN|19|23|Milites ergo cum crucifixissent Iesum, acceperunt vestimenta eius et fecerunt quattuor partes, unicuique militi partem, et tunicam. Erat autem tunica inconsutilis, desuper contexta per totum.
JOHN|19|24|Dixerunt ergo ad invicem: " Non scindamus eam, sed sortiamur de illa,cuius sit ", ut Scriptura impleatur dicens: Partiti sunt vestimenta mea sibiet in vestem meam miserunt sortem ".Et milites quidem haec fecerunt.
JOHN|19|25|Stabant autem iuxta crucem Iesu mater eius et soror matris eius, Maria Cleopae, et Maria Magdalene.
JOHN|19|26|Cum vidisset ergo Iesus matrem et discipulum stantem, quem diligebat, dicit matri: " Mulier, ecce filius tuus ".
JOHN|19|27|Deinde dicit discipulo: " Ecce mater tua ". Et ex illa hora accepit eam discipulus in sua.
JOHN|19|28|Post hoc sciens Iesus quia iam omnia consummata sunt, ut consummaretur Scriptura, dicit: " Sitio ".
JOHN|19|29|Vas positum erat aceto plenum; spongiam ergo plenam aceto hyssopo circumponentes, obtulerunt ori eius.
JOHN|19|30|Cum ergo accepisset acetum, Iesus dixit: " Consummatum est! ". Et inclinato capite tradidit spiritum.
JOHN|19|31|Iudaei ergo, quoniam Parasceve erat, ut non remanerent in cruce corpora sabbato, erat enim magnus dies illius sabbati, rogaverunt Pilatum, ut frangerentur eorum crura, et tollerentur.
JOHN|19|32|Venerunt ergo milites et primi quidem fregerunt crura et alterius, qui crucifixus est cum eo;
JOHN|19|33|ad Iesum autem cum venissent, ut viderunt eum iam mortuum, non fregerunt eius crura,
JOHN|19|34|sed unus militum lancea latus eius aperuit, et continuo exivit sanguis et aqua.
JOHN|19|35|Et qui vidit, testimonium perhibuit, et verum est eius testimonium, et ille scit quia vera dicit, ut et vos credatis.
JOHN|19|36|Facta sunt enim haec, ut Scriptura impleatur: " Os non comminuetur eius,
JOHN|19|37|et iterum alia Scriptura dicit: " Videbunt in quem transfixerunt ".
JOHN|19|38|Post haec autem rogavit Pilatum Ioseph ab Arimathaea, qui erat discipulus Iesu, occultus autem propter metum Iudaeorum, ut tolleret corpus Iesu; et permisit Pilatus. Venit ergo et tulit corpus eius.
JOHN|19|39|Venit autem et Nicodemus, qui venerat ad eum nocte primum, ferens mixturam myrrhae et aloes quasi libras centum.
JOHN|19|40|Acceperunt ergo corpus Iesu et ligaverunt illud linteis cum aromatibus, sicut mos Iudaeis est sepelire.
JOHN|19|41|Erat autem in loco, ubi crucifixus est, hortus, et in horto monumentum novum, in quo nondum quisquam positus erat.
JOHN|19|42|Ibi ergo propter Parascevem Iudaeorum, quia iuxta erat monumentum, posuerunt Iesum.
JOHN|20|1|Prima autem sabbatorum Maria Magdalene venit ma ne, cum adhuc tenebrae essent, ad monumentum et videt lapidem sublatum a monumento.
JOHN|20|2|Currit ergo et venit ad Simonem Petrum et ad alium discipulum, quem amabat Iesus, et dicit eis: " Tulerunt Dominum de monumento, et nescimus, ubi posuerunt eum! ".
JOHN|20|3|Exiit ergo Petrus et ille alius discipulus, et veniebant ad monumentum.
JOHN|20|4|Currebant autem duo simul, et ille alius discipulus praecucurrit citius Petro et venit primus ad monumentum;
JOHN|20|5|et cum se inclinasset, videt posita linteamina, non tamen introivit.
JOHN|20|6|Venit ergo et Simon Petrus sequens eum et introivit in monumentum; et videt linteamina posita
JOHN|20|7|et sudarium, quod fuerat super caput eius, non cum linteaminibus positum, sed separatim involutum in unum locum.
JOHN|20|8|Tunc ergo introivit et alter discipulus, qui venerat primus ad monumentum, et vidit et credidit.
JOHN|20|9|Nondum enim sciebant Scripturam, quia oportet eum a mortuis resurgere.
JOHN|20|10|Abierunt ergo iterum ad semetipsos discipuli.
JOHN|20|11|Maria autem stabat ad monumentum foris plorans. Dum ergo fleret, inclinavit se in monumentum
JOHN|20|12|et videt duos angelos in albis sedentes, unum ad caput et unum ad pedes, ubi positum fuerat corpus Iesu.
JOHN|20|13|Et dicunt ei illi: " Mulier, quid ploras? ". Dicit eis: " Tulerunt Dominum meum, et nescio, ubi posuerunt eum ".
JOHN|20|14|Haec cum dixisset, conversa est retrorsum et videt Iesum stantem; et non sciebat quia Iesus est.
JOHN|20|15|Dicit ei Iesus: " Mulier, quid ploras? Quem quaeris? ". Illa, existimans quia hortulanus esset, dicit ei: " Domine, si tu sustulisti eum, dicito mihi, ubi posuisti eum, et ego eum tollam ".
JOHN|20|16|Dicit ei Iesus: " Maria! ". Conversa illa dicit ei Hebraice: " Rabbuni! - quod dicitur Magister C.
JOHN|20|17|Dicit ei Iesus: " Iam noli me tenere, nondum enim ascendi ad Patrem; vade autem ad fratres meos et dic eis: Ascendo ad Patrem meum et Patrem vestrum, et Deum meum et Deum vestrum ".
JOHN|20|18|Venit Maria Magdalene annuntians discipulis: " Vidi Dominum! ", et quia haec dixit ei.
JOHN|20|19|Cum esset ergo sero die illa prima sabbatorum, et fores essent clausae, ubi erant discipuli, propter metum Iudaeorum, venit Iesus et stetit in medio et dicit eis: " Pax vobis! ".
JOHN|20|20|Et hoc cum dixisset, ostendit eis manus et latus. Gavisi sunt ergo discipuli, viso Domino.
JOHN|20|21|Dixit ergo eis iterum: " Pax vobis! Sicut misit me Pater, et ego mitto vos ".
JOHN|20|22|Et cum hoc dixisset, insufflavit et dicit eis: " Accipite Spiritum Sanctum.
JOHN|20|23|Quorum remiseritis peccata, remissa sunt eis; quorum retinueritis, retenta sunt ".
JOHN|20|24|Thomas autem, unus ex Duodecim, qui dicitur Didymus, non erat cum eis, quando venit Iesus.
JOHN|20|25|Dicebant ergo ei alii discipuli: " Vidimus Dominum! ". Ille autem dixit eis: " Nisi videro in manibus eius signum clavorum et mittam digitum meum in signum clavorum et mittam manum meam in latus eius, non credam ".
JOHN|20|26|Et post dies octo iterum erant discipuli eius intus, et Thomas cum eis. Venit Iesus ianuis clausis et stetit in medio et dixit: " Pax vobis! ".
JOHN|20|27|Deinde dicit Thomae: " Infer digitum tuum huc et vide manus meas et affer manum tuam et mitte in latus meum; et noli fieri incredulus sed fidelis! ".
JOHN|20|28|Respondit Thomas et dixit ei: " Dominus meus et Deus meus! ".
JOHN|20|29|Dicit ei Iesus: " Quia vidisti me, credidisti. Beati, qui non viderunt et crediderunt! ".
JOHN|20|30|Multa quidem et alia signa fecit Iesus in conspectu discipulorum suorum, quae non sunt scripta in libro hoc;
JOHN|20|31|haec autem scripta sunt, ut credatis quia Iesus est Christus Filius Dei et ut credentes vitam habeatis in nomine eius.
JOHN|21|1|Postea manifestavit se ite rum Iesus discipulis ad mare Tiberiadis; manifestavit autem sic.
JOHN|21|2|Erant simul Simon Petrus et Thomas, qui dicitur Didymus, et Nathanael, qui erat a Cana Galilaeae, et filii Zebedaei et alii ex discipulis eius duo.
JOHN|21|3|Dicit eis Simon Petrus: " Vado piscari ". Dicunt ei: " Venimus et nos tecum ". Exierunt et ascenderunt in navem; et illa nocte nihil prendiderunt.
JOHN|21|4|Mane autem iam facto, stetit Iesus in litore; non tamen sciebant discipuli quia Iesus est.
JOHN|21|5|Dicit ergo eis Iesus: " Pueri, numquid pulmentarium habetis? ". Responderunt ei: " Non ".
JOHN|21|6|Ille autem dixit eis: " Mittite in dexteram navigii rete et invenietis. Miserunt ergo et iam non valebant illud trahere a multitudine piscium.
JOHN|21|7|Dicit ergo discipulus ille, quem diligebat Iesus, Petro: " Dominus est!. Simon ergo Petrus, cum audisset quia Dominus est, tunicam succinxit se, erat enim nudus, et misit se in mare;
JOHN|21|8|alii autem discipuli navigio venerunt, non enim longe erant a terra, sed quasi cubitis ducentis, trahentes rete piscium.
JOHN|21|9|Ut ergo descenderunt in terram, vident prunas positas et piscem superpositum et panem.
JOHN|21|10|Dicit eis Iesus: " Afferte de piscibus, quos prendidistis nunc ".
JOHN|21|11|Ascendit ergo Simon Petrus et traxit rete in terram, plenum magnis piscibus centum quinquaginta tribus; et cum tanti essent, non est scissum rete.
JOHN|21|12|Dicit eis Iesus: " Venite, prandete ". Nemo autem audebat discipulorum interrogare eum: " Tu quis es? ", scientes quia Dominus est.
JOHN|21|13|Venit Iesus et accipit panem et dat eis et piscem similiter.
JOHN|21|14|Hoc iam tertio manifestatus est Iesus discipulis, cum resurrexisset a mortuis.
JOHN|21|15|Cum ergo prandissent, dicit Simoni Petro Iesus: " Simon Ioannis, diligis me plus his? ". Dicit ei: " Etiam, Domine, tu scis quia amo te ". Dicit ei: " Pasce agnos meos ".
JOHN|21|16|Dicit ei iterum secundo: " Simon Ioannis, diligis me? ". Ait illi: " Etiam, Domine, tu scis quia amo te ". Dicit ei: " Pasce oves meas ".
JOHN|21|17|Dicit ei tertio: " Simon Ioannis, amas me? ". Contristatus est Petrus quia dixit ei tertio: " Amas me? ", et dicit ei: " Domine, tu omnia scis, tu cognoscis quia amo te ". Dicit ei: " Pasce oves meas.
JOHN|21|18|Amen, amen dico tibi: Cum esses iunior, cingebas teipsum et ambulabas, ubi volebas; cum autem senueris, extendes manus tuas, et alius te cinget et ducet, quo non vis ".
JOHN|21|19|Hoc autem dixit significans qua morte clarificaturus esset Deum. Et hoc cum dixisset, dicit ei: " Sequere me ".
JOHN|21|20|Conversus Petrus videt illum discipulum, quem diligebat Iesus, sequentem, qui et recubuit in cena super pectus eius et dixit: " Domine, quis est qui tradit te? ".
JOHN|21|21|Hunc ergo cum vidisset Petrus, dicit Iesu: " Domine, hic autem quid? ".
JOHN|21|22|Dicit ei Iesus: " Si eum volo manere donec veniam, quid ad te? Tu me sequere ".
JOHN|21|23|Exivit ergo sermo iste in fratres, quia discipulus ille non moritur. Non autem dixit ei Iesus: " Non moritur ", sed: " Si eum volo manere donec veniam, quid ad te? ".
JOHN|21|24|Hic est discipulus, qui testimonium perhibet de his et scripsit haec; et scimus quia verum est testimonium eius.
JOHN|21|25|Sunt autem et alia multa, quae fecit Iesus; quae, si scribantur per singula, nec ipsum arbitror mundum capere eos, qui scribendi sunt, libros.
ACTS|1|1|Primum quidem sermonem feci de omnibus, o Theophile, quae coepit Iesus facere et docere,
ACTS|1|2|usque in diem, qua, cum praecepisset apostolis per Spiritum Sanctum, quos elegit, assumptus est;
ACTS|1|3|quibus et praebuit seipsum vivum post passionem suam in multis argumentis, per dies quadraginta apparens eis et loquens ea, quae sunt de regno Dei.
ACTS|1|4|Et convescens praecepit eis ab Hierosolymis ne discederent, sed exspectarent promissionem Patris: " Quam audistis a me,
ACTS|1|5|quia Ioannes quidem baptizavit aqua, vos autem baptizabimini in Spiritu Sancto non post multos hos dies ".
ACTS|1|6|Igitur qui convenerant, interrogabant eum dicentes: " Domine, si in tempore hoc restitues regnum Israeli? ".
ACTS|1|7|Dixit autem eis: " Non est vestrum nosse tempora vel momenta, quae Pater posuit in sua potestate,
ACTS|1|8|sed accipietis virtutem, superveniente Sancto Spiritu in vos, et eritis mihi testes et in Ierusalem et in omni Iudaea et Samaria et usque ad ultimum terrae ".
ACTS|1|9|Et cum haec dixisset, videntibus illis, elevatus est, et nubes suscepit eum ab oculis eorum.
ACTS|1|10|Cumque intuerentur in caelum, eunte illo, ecce duo viri astiterunt iuxta illos in vestibus albis,
ACTS|1|11|qui et dixerunt: " Viri Galilaei, quid statis aspicientes in caelum? Hic Iesus, qui assumptus est a vobis in caelum, sic veniet quemadmodum vidistis eum euntem in caelum ".
ACTS|1|12|Tunc reversi sunt in Ierusalem a monte, qui vocatur Oliveti, qui est iuxta Ierusalem sabbati habens iter.
ACTS|1|13|Et cum introissent, in cenaculum ascenderunt, ubi manebant et Petrus et Ioannes et Iacobus et Andreas, Philippus et Thomas, Bartholomaeus et Matthaeus, Iacobus Alphaei et Simon Zelotes et Iudas Iacobi.
ACTS|1|14|Hi omnes erant perseverantes unanimiter in oratione cum mulieribus et Maria matre Iesu et fratribus eius.
ACTS|1|15|Et in diebus illis exsurgens Petrus in medio fratrum dixit - erat autem turba hominum simul fere centum viginti C:
ACTS|1|16|" Viri fratres, oportebat impleri Scripturam, quam praedixit Spiritus Sanctus per os David de Iuda, qui fuit dux eorum, qui comprehenderunt Iesum,
ACTS|1|17|quia connumeratus erat in nobis et sortitus est sortem ministerii huius.
ACTS|1|18|Hic quidem possedit agrum de mercede iniquitatis; et pronus factus crepuit medius, et diffusa sunt omnia viscera eius.
ACTS|1|19|Et notum factum est omnibus habitantibus Ierusalem, ita ut appellaretur ager ille lingua eorum Aceldamach, hoc est ager Sanguinis.
ACTS|1|20|Scriptum est enim in libro Psalmorum:Fiat commoratío eius deserta,et non sit qui inhabitet in ea"et: "Episcopatum eius accipiat alius".
ACTS|1|21|Oportet ergo ex his viris, qui nobiscum congregati erant in omni tempore, quo intravit et exivit inter nos Dominus Iesus,
ACTS|1|22|incipiens a baptismate Ioannis usque in diem, qua assumptus est a nobis, testem resurrectionis eius nobiscum fieri unum ex istis ".
ACTS|1|23|Et statuerunt duos, Ioseph, qui vocabatur Barsabbas, qui cognominatus est Iustus, et Matthiam.
ACTS|1|24|Et orantes dixerunt: " Tu, Domine, qui corda nosti omnium, ostende quem elegeris ex his duobus unum
ACTS|1|25|accipere locum ministerii huius et apostolatus, de quo praevaricatus est Iudas, ut abiret in locum suum ".
ACTS|1|26|Et dederunt sortes eis, et cecidit sors super Matthiam, et annumeratus est cum undecim apostolis.
ACTS|2|1|Et cum compleretur dies Pen tecostes, erant omnes pariter in eodem loco.
ACTS|2|2|Et factus est repente de caelo sonus tamquam advenientis spiritus vehementis et replevit totam domum, ubi erant sedentes.
ACTS|2|3|Et apparuerunt illis dispertitae linguae tamquam ignis, seditque supra singulos eorum;
ACTS|2|4|et repleti sunt omnes Spiritu Sancto et coeperunt loqui aliis linguis, prout Spiritus dabat eloqui illis.
ACTS|2|5|Erant autem in Ierusalem habitantes Iudaei, viri religiosi ex omni natione, quae sub caelo est;
ACTS|2|6|facta autem hac voce, convenit multitudo et confusa est, quoniam audiebat unusquisque lingua sua illos loquentes.
ACTS|2|7|Stupebant autem et mirabantur dicentes: " Nonne ecce omnes isti, qui loquuntur, Galilaei sunt?
ACTS|2|8|Et quomodo nos audimus unusquisque propria lingua nostra, in qua nati sumus?
ACTS|2|9|Parthi et Medi et Elamitae et qui habitant Mesopotamiam, Iudaeam quoque et Cappadociam, Pontum et Asiam,
ACTS|2|10|Phrygiam quoque et Pamphyliam, Aegyptum et partes Libyae, quae est circa Cyrenem, et advenae Romani,
ACTS|2|11|Iudaei quoque et proselyti, Cretes et Arabes, audimus loquentes eos nostris linguis magnalia Dei ".
ACTS|2|12|Stupebant autem omnes et haesitabant ad invicem dicentes: " Quidnam hoc vult esse? ";
ACTS|2|13|alii autem irridentes dicebant: " Musto pleni sunt isti ".
ACTS|2|14|Stans autem Petrus cum Undecim levavit vocem suam et locutus est eis: " Viri Iudaei et qui habitatis Ierusalem universi, hoc vobis notum sit, et auribus percipite verba mea.
ACTS|2|15|Non enim, sicut vos aestimatis, hi ebrii sunt, est enim hora diei tertia;
ACTS|2|16|sed hoc est, quod dictum est per prophetam Ioel:
ACTS|2|17|"Et erit: in novissimis diebus, dicit Deus,effundam de Spiritu meo super omnem carnem,et prophetabunt filii vestri et filiae vestrae,et iuvenes vestri visiones videbunt,et seniores vestri somnia somniabunt;
ACTS|2|18|et quidem super servos meos et super ancillas measin diebus illis effundam de Spiritu meo,et prophetabunt.
ACTS|2|19|Et dabo prodigia in caelo sursum et signa in terra deorsum,sanguinem et ignem et vaporem fumi;
ACTS|2|20|sol convertetur in tenebras,et luna in sanguinem,antequam veniat dies Dominimagnus et manifestus.
ACTS|2|21|Et erit:omnis quicumque invocaverit nomen Domini, salvus erit".
ACTS|2|22|Viri Israelitae, audite verba haec: Iesum Nazarenum, virum approbatum a Deo apud vos virtutibus et prodigiis et signis, quae fecit per illum Deus in medio vestri, sicut ipsi scitis,
ACTS|2|23|hunc definito consilio et praescientia Dei traditum per manum iniquorum affigentes interemistis,
ACTS|2|24|quem Deus suscitavit, solutis doloribus mortis, iuxta quod impossibile erat teneri illum ab ea.
ACTS|2|25|David enim dicit circa eum:Providebam Dominum coram me semper, quoniam a dextris meis est, ne commovear.
ACTS|2|26|Propter hoc laetatum est cor meum,et exsultavit lingua mea;insuper et caro mea requiescet in spe.
ACTS|2|27|Quoniam non derelinques animam meam in infernoneque dabis Sanctum tuum videre corruptionem.
ACTS|2|28|Notas fecisti mihi vias vitae,replebis me iucunditate cum facie tua".
ACTS|2|29|Viri fratres, liceat audenter dicere ad vos de patriarcha David, quoniam et defunctus est et sepultus est, et sepulcrum eius est apud nos usque in hodiernum diem;
ACTS|2|30|propheta igitur cum esset et sciret quia iure iurando iurasset illi Deus de fructu lumbi eius sedere super sedem eius,
ACTS|2|31|providens locutus est de resurrectione Christi, quia neque derelictus est in inferno, neque caro eius vidit corruptionem.
ACTS|2|32|Hunc Iesum resuscitavit Deus, cuius omnes nos testes sumus.
ACTS|2|33|Dextera igitur Dei exaltatus, et promissione Spiritus Sancti accepta a Patre, effudit hunc, quem vos videtis et auditis.
ACTS|2|34|Non enim David ascendit in caelos; dicit autem ipse:Dixit Dominus Domino meo: Sede a dextris meis,
ACTS|2|35|donec ponam inimicos tuos scabellum pedum tuorum".
ACTS|2|36|Certissime ergo sciat omnis domus Israel quia et Dominum eum et Christum Deus fecit, hunc Iesum, quem vos crucifixistis ".
ACTS|2|37|His auditis, compuncti sunt corde et dixerunt ad Petrum et reliquos apostolos: " Quid faciemus, viri fratres? ".
ACTS|2|38|Petrus vero ad illos: " Paenitentiam, inquit, agite, et baptizetur unusquisque vestrum in nomine Iesu Christi in remissionem peccatorum vestrorum, et accipietis donum Sancti Spiritus;
ACTS|2|39|vobis enim est repromissio et filiis vestris et omnibus, qui longe sunt, quoscumque advocaverit Dominus Deus noster ".
ACTS|2|40|Aliis etiam verbis pluribus testificatus est et exhortabatur eos dicens: " Salvamini a generatione ista prava ".
ACTS|2|41|Qui ergo, recepto sermone eius, baptizati sunt; et appositae sunt in il la die animae circiter tria milia.
ACTS|2|42|Erant autem perseverantes in doctrina apostolorum et communicatione, in fractione panis et orationibus.
ACTS|2|43|Fiebat autem omni animae timor; multa quoque prodigia et signa per apostolos fiebant.
ACTS|2|44|Omnes autem, qui crediderant, erant pariter et habebant omnia communia;
ACTS|2|45|et possessiones et substantias vendebant et dividebant illas omnibus, prout cuique opus erat;
ACTS|2|46|cotidie quoque perdurantes unanimiter in templo et frangentes circa domos panem, sumebant cibum cum exsultatione et simplicitate cordis,
ACTS|2|47|collaudantes Deum et habentes gratiam ad omnem plebem. Dominus autem augebat, qui salvi fierent cotidie in idipsum.
ACTS|3|1|Petrus autem et Ioannes ascen debant in templum ad horam orationis nonam.
ACTS|3|2|Et quidam vir, qui erat claudus ex utero matris suae, baiulabatur; quem ponebant cotidie ad portam templi, quae dicitur Speciosa, ut peteret eleemosynam ab introeuntibus in templum;
ACTS|3|3|is cum vidisset Petrum et Ioannem incipientes introire in templum, rogabat, ut eleemosynam acciperet.
ACTS|3|4|Intuens autem in eum Petrus cum Ioanne dixit: " Respice in nos ".
ACTS|3|5|At ille intendebat in eos, sperans se aliquid accepturum ab eis.
ACTS|3|6|Petrus autem dixit: " Argentum et aurum non est mihi; quod autem habeo, hoc tibi do: In nomine Iesu Christi Nazareni surge et ambula! ".
ACTS|3|7|Et apprehensa ei manu dextera, allevavit eum; et protinus consolidatae sunt bases eius et tali,
ACTS|3|8|et exsiliens stetit et ambulabat; et intravit cum illis in templum, ambulans et exsiliens et laudans Deum.
ACTS|3|9|Et vidit omnis populus eum ambulantem et laudantem Deum;
ACTS|3|10|cognoscebant autem illum quoniam ipse erat, qui ad eleemosynam sedebat ad Speciosam portam templi, et impleti sunt stupore et exstasi in eo, quod contigerat illi.
ACTS|3|11|Cum teneret autem Petrum et Ioannem, concurrit omnis populus ad eos ad porticum, qui appellatur Salomonis, stupentes.
ACTS|3|12|Videns autem Petrus respondit ad populum: " Viri Israelitae, quid miramini in hoc aut nos quid intuemini, quasi nostra virtute aut pietate fecerimus hunc ambulare?
ACTS|3|13|Deus Abraham et Deus Isaac et Deus Iacob, Deus patrum nostrorum, glorificavit puerum suum Iesum, quem vos quidem tradidistis et negastis ante faciem Pilati, iudicante illo dimitti;
ACTS|3|14|vos autem Sanctum et Iustum negastis et petistis virum homicidam donari vobis,
ACTS|3|15|ducem vero vitae interfecistis, quem Deus suscitavit a mortuis, cuius nos testes sumus.
ACTS|3|16|Et in fide nominis eius hunc, quem videtis et nostis, confirmavit nomen eius; et fides, quae per eum est, dedit huic integritatem istam in conspectu omnium vestrum.
ACTS|3|17|Et nunc, fratres, scio quia per ignorantiam fecistis, sicut et principes vestri;
ACTS|3|18|Deus autem, quae praenuntiavit per os omnium Prophetarum pati Christum suum, implevit sic.
ACTS|3|19|Paenitemini igitur et convertimini, ut deleantur vestra peccata,
ACTS|3|20|ut veniant tempora refrigerii a conspectu Domini, et mittat eum, qui praedestinatus est vobis Christus, Iesum,
ACTS|3|21|quem oportet caelum quidem suscipere usque in tempora restitutionis omnium, quae locutus est Deus per os sanctorum a saeculo suorum prophetarum.
ACTS|3|22|Moyses quidem dixit: "Prophetam vobis suscitabit Dominus Deus vester de fratribus vestris tamquam me; ipsum audietis iuxta omnia, quaecumque locutus fuerit vobis.
ACTS|3|23|Erit autem: omnis anima, quae non audierit prophetam illum, exterminabitur de plebe".
ACTS|3|24|Et omnes prophetae a Samuel et deinceps quotquot locuti sunt, etiam annuntiaverunt dies istos.
ACTS|3|25|Vos estis filii prophetarum et testamenti, quod disposuit Deus ad patres vestros dicens ad Abraham: "Et in semine tuo benedicentur omnes familiae terrae".
ACTS|3|26|Vobis primum Deus suscitans Puerum suum, misit eum benedicentem vobis in avertendo unumquemque a nequitiis vestris ".
ACTS|4|1|Loquentibus autem illis ad populum, supervenerunt eis sa cerdotes et magistratus templi et sadducaei,
ACTS|4|2|dolentes quod docerent populum et annuntiarent in Iesu resurrectionem ex mortuis;
ACTS|4|3|et iniecerunt in eos manus et posuerunt in custodiam in crastinum; erat enim iam vespera.
ACTS|4|4|Multi autem eorum, qui audierant verbum, crediderunt; et factus est numerus virorum quinque milia.
ACTS|4|5|Factum est autem in crastinum, ut congregarentur principes eorum et seniores et scribae in Ierusalem,
ACTS|4|6|et Annas princeps sacerdotum et Caiphas et Ioannes et Alexander et quotquot erant de genere sacerdotali,
ACTS|4|7|et statuentes eos in medio interrogabant: " In qua virtute aut in quo nomine fecistis hoc vos? ".
ACTS|4|8|Tunc Petrus repletus Spiritu Sancto dixit ad eos: " Principes populi et seniores,
ACTS|4|9|si nos hodie diiudicamur in benefacto hominis infirmi, in quo iste salvus factus est,
ACTS|4|10|notum sit omnibus vobis et omni plebi Israel quia in nomine Iesu Christi Nazareni, quem vos crucifixistis, quem Deus suscitavit a mortuis, in hoc iste astat coram vobis sanus.
ACTS|4|11|Hic estlapis, qui reprobatus est a vobis aedificatoribus,qui factus est in caput anguli.
ACTS|4|12|Et non est in alio aliquo salus, nec enim nomen aliud est sub caelo datum in hominibus, in quo oportet nos salvos fieri ".
ACTS|4|13|Videntes autem Petri fiduciam et Ioannis, et comperto quod homines essent sine litteris et idiotae, admirabantur et cognoscebant eos quoniam cum Iesu fuerant;
ACTS|4|14|hominem quoque videntes stantem cum eis, qui curatus fuerat, nihil poterant contradicere.
ACTS|4|15|Iubentes autem eos foras extra concilium secedere, conferebant ad invicem
ACTS|4|16|dicentes: " Quid faciemus hominibus istis? Quoniam quidem notum signum factum est per eos omnibus habitantibus in Ierusalem manifestum, et non possumus negare;
ACTS|4|17|sed ne amplius divulgetur in populum, comminemur eis, ne ultra loquantur in nomine hoc ulli hominum ".
ACTS|4|18|Et vocantes eos denuntiaverunt, ne omnino loquerentur neque docerent in nomine Iesu.
ACTS|4|19|Petrus vero et Ioannes respondentes dixerunt ad eos: " Si iustum est in conspectu Dei vos potius audire quam Deum, iudicate;
ACTS|4|20|non enim possumus nos, quae vidimus et audivimus, non loqui ".
ACTS|4|21|At illi ultra comminantes dimiserunt eos, nequaquam invenientes, quomodo punirent eos, propter populum, quia omnes glorificabant Deum in eo, quod acciderat;
ACTS|4|22|annorum enim erat amplius quadraginta homo, in quo factum erat signum istud sanitatis.
ACTS|4|23|Dimissi autem venerunt ad suos et annuntiaverunt quanta ad eos principes sacerdotum et seniores dixissent.
ACTS|4|24|Qui cum audissent, unanimiter levaverunt vocem ad Deum et dixerunt: " Domine, tu, qui fecisti caelum et terram et mare et omnia, quae in eis sunt,
ACTS|4|25|qui Spiritu Sancto per os patris nostri David pueri tui dixisti:Quare fremuerunt gentes,et populi meditati sunt inania?
ACTS|4|26|Astiterunt reges terrae,et principes convenerunt in unumadversus Dominum et adversus Christum eius".
ACTS|4|27|Convenerunt enim vere in civitate ista adversus sanctum puerum tuum Iesum, quem unxisti, Herodes et Pontius Pilatus cum gentibus et populis Israel
ACTS|4|28|facere, quaecumque manus tua et consilium praedestinavit fieri.
ACTS|4|29|Et nunc, Domine, respice in minas eorum et da servis tuis cum omni fiducia loqui verbum tuum,
ACTS|4|30|in eo quod manum tuam extendas ad sanitatem et signa et prodigia facienda per nomen sancti pueri tui Iesu ".
ACTS|4|31|Et cum orassent, motus est locus, in quo erant congregati, et repleti sunt omnes Sancto Spiritu et loquebantur verbum Dei cum fiducia.
ACTS|4|32|Multitudinis autem credentium erat cor et anima una, nec quisquam eorum, quae possidebant, aliquid suum esse dicebat, sed erant illis omnia communia.
ACTS|4|33|Et virtute magna reddebant apostoli testimonium resurrectionis Domini Iesu, et gratia magna erat super omnibus illis.
ACTS|4|34|Neque enim quisquam egens erat inter illos; quotquot enim possessores agrorum aut domorum erant, vendentes afferebant pretia eorum, quae vendebant,
ACTS|4|35|et ponebant ante pedes apostolorum; dividebatur autem singulis, prout cuique opus erat.
ACTS|4|36|Ioseph autem, qui cognominatus est Barnabas ab apostolis - quod est interpretatum filius Consolationis - Levites, Cyprius genere,
ACTS|4|37|cum haberet agrum, vendidit et attulit pecuniam et posuit ante pedes apostolorum.
ACTS|5|1|Vir autem quidam nomine Ananias cum Sapphira uxore sua vendidit agrum
ACTS|5|2|et subtraxit de pretio, conscia quoque uxore, et afferens partem quandam ad pedes apostolorum posuit.
ACTS|5|3|Dixit autem Petrus: " Anania, cur implevit Satanas cor tuum mentiri te Spiritui Sancto et subtrahere de pretio agri?
ACTS|5|4|Nonne manens tibi manebat et venumdatum in tua erat potestate? Quare posuisti in corde tuo hanc rem? Non es mentitus hominibus sed Deo! ".
ACTS|5|5|Audiens autem Ananias haec verba cecidit et exspiravit; et factus est timor magnus in omnes audientes.
ACTS|5|6|Surgentes autem iuvenes involverunt eum et efferentes sepelierunt.
ACTS|5|7|Factum est autem quasi horarum trium spatium, et uxor ipsius nesciens, quod factum fuerat, introivit.
ACTS|5|8|Respondit autem ei Petrus: " Dic mihi, si tanti agrum vendidistis? ". At illa dixit: " Etiam, tanti ".
ACTS|5|9|Petrus autem ad eam: " Quid est quod convenit vobis tentare Spiritum Domini? Ecce pedes eorum, qui sepelierunt virum tuum, ad ostium, et efferent te ".
ACTS|5|10|Confestim cecidit ante pedes eius et exspiravit; intrantes autem iuvenes invenerunt illam mortuam et efferentes sepelierunt ad virum suum.
ACTS|5|11|Et factus est timor magnus super universam ecclesiam et in omnes, qui audierunt haec.
ACTS|5|12|Per manus autem apostolorum fiebant signa et prodigia multa in plebe; et erant unanimiter omnes in porticu Salomonis.
ACTS|5|13|Ceterorum autem nemo audebat coniungere se illis, sed magnificabat eos populus;
ACTS|5|14|magis autem addebantur credentes Domino multitudines virorum ac mulierum,
ACTS|5|15|ita ut et in plateas efferrent infirmos et ponerent in lectulis et grabatis, ut, veniente Petro, saltem umbra illius obumbraret quemquam eorum.
ACTS|5|16|Concurrebat autem et multitudo vicinarum civitatum Ierusalem, afferentes aegros et vexatos ab spiritibus immundis, qui curabantur omnes.
ACTS|5|17|Exsurgens autem princeps sacerdotum et omnes, qui cum illo erant, quae est haeresis sadducaeorum, repleti sunt zelo
ACTS|5|18|et iniecerunt manus in apostolos et posuerunt illos in custodia publica.
ACTS|5|19|Angelus autem Domini per noctem aperuit ianuas carceris et educens eos dixit:
ACTS|5|20|" Ite et stantes loquimini in templo plebi omnia verba vitae huius ".
ACTS|5|21|Qui cum audissent, intraverunt diluculo in templum et docebant.Adveniens autem princeps sacerdotum et, qui cum eo erant, convocaverunt concilium et omnes seniores filiorum Israel et miserunt in carcerem, ut adducerentur illi.
ACTS|5|22|Cum venissent autem ministri, non invenerunt illos in carcere; reversi autem nuntiaverunt
ACTS|5|23|dicentes: " Carcerem invenimus clausum cum omni diligentia et custodes stantes ad ianuas; aperientes autem intus neminem invenimus! ".
ACTS|5|24|Ut audierunt autem hos sermones, magistratus templi et principes sacerdotum ambigebant de illis quidnam fieret illud.
ACTS|5|25|Adveniens autem quidam nuntiavit eis: " Ecce viri, quos posuistis in carcere, sunt in templo stantes et docentes populum ".
ACTS|5|26|Tunc abiens magistratus cum ministris adducebat illos, non per vim; timebant enim populum, ne lapidarentur.
ACTS|5|27|Et cum adduxissent illos, statuerunt in concilio. Et interrogavit eos princeps sacerdotum
ACTS|5|28|dicens: " Nonne praecipiendo praecepimus vobis, ne doceretis in nomine isto? Et ecce replevistis Ierusalem doctrina vestra et vultis inducere super nos sanguinem hominis istius ".
ACTS|5|29|Respondens autem Petrus et apostoli dixerunt: " Oboedire oportet Deo magis quam hominibus.
ACTS|5|30|Deus patrum nostrorum suscitavit Iesum, quem vos interemistis suspendentes in ligno;
ACTS|5|31|hunc Deus Ducem et Salvatorem exaltavit dextera sua ad dandam paenitentiam Israel et remissionem peccatorum.
ACTS|5|32|Et nos sumus testes horum verborum, et Spiritus Sanctus, quem dedit Deus oboedientibus sibi ".
ACTS|5|33|Haec cum audissent, dissecabantur et volebant interficere illos.
ACTS|5|34|Surgens autem quidam in concilio pharisaeus nomine Gamaliel, legis doctor honorabilis universae plebi, iussit foras ad breve homines fieri
ACTS|5|35|dixitque ad illos: " Viri Israelitae, attendite vobis super hominibus istis quid acturi sitis.
ACTS|5|36|Ante hos enim dies exstitit Theudas dicens esse se aliquem, cui consensit virorum numerus circiter quadringentorum; qui occisus est, et omnes, quicumque credebant ei, dissipati sunt et redacti sunt ad nihilum.
ACTS|5|37|Post hunc exstitit Iudas Galilaeus in diebus census et avertit populum post se; et ipse periit, et omnes, quotquot consentiebant ei, dispersi sunt.
ACTS|5|38|Et nunc dico vobis: Discedite ab hominibus istis et sinite illos. Quoniam si est ex hominibus consilium hoc aut opus hoc, dissolvetur;
ACTS|5|39|si vero ex Deo est, non poteritis dissolvere eos, ne forte et adversus Deum pugnantes inveniamini! ".Consenserunt autem illi
ACTS|5|40|et convocantes apostolos, caesis denuntiaverunt, ne loquerentur in nomine Iesu, et dimiserunt eos.
ACTS|5|41|Et illi quidem ibant gaudentes a conspectu concilii, quoniam digni habiti sunt pro nomine contumeliam pati;
ACTS|5|42|et omni die in templo et circa domos non cessabant docentes et evangelizantes Christum, Iesum.
ACTS|6|1|In diebus autem illis, crescente numero discipulorum, factus est murmur Graecorum adversus Hebraeos, eo quod neglegerentur in ministerio cotidiano viduae eorum.
ACTS|6|2|Convocantes autem Duodecim multitudinem discipulorum, dixerunt: " Non est aequum nos derelinquentes verbum Dei ministrare mensis;
ACTS|6|3|considerate vero, fratres, viros ex vobis boni testimonii septem plenos Spiritu et sapientia, quos constituemus super hoc opus;
ACTS|6|4|nos vero orationi et ministerio verbi instantes erimus ".
ACTS|6|5|Et placuit sermo coram omni multitudine; et elegerunt Stephanum, virum plenum fide et Spiritu Sancto, et Philippum et Prochorum et Nicanorem et Timonem et Parmenam et Nicolaum proselytum Antiochenum,
ACTS|6|6|quos statuerunt ante conspectum apostolorum, et orantes imposuerunt eis manus.
ACTS|6|7|Et verbum Dei crescebat, et multiplicabatur numerus discipulorum in Ierusalem valde; multa etiam turba sacerdotum oboediebat fidei.
ACTS|6|8|Stephanus autem plenus gratia et virtute faciebat prodigia et signa magna in populo.
ACTS|6|9|Surrexerunt autem quidam de synagoga, quae appellatur Libertinorum et Cyrenensium et Alexandrinorum et eorum, qui erant a Cilicia et Asia, disputantes cum Stephano;
ACTS|6|10|et non poterant resistere sapientiae et Spiritui, quo loquebatur.
ACTS|6|11|Tunc submiserunt viros, qui dicerent: " Audivimus eum dicentem verba blasphema in Moysen et Deum ";
ACTS|6|12|et commoverunt plebem et seniores et scribas, et concurrentes rapuerunt eum et adduxerunt in concilium
ACTS|6|13|et statuerunt testes falsos dicentes: " Homo iste non cessat loqui verba adversus locum sanctum et Legem;
ACTS|6|14|audivimus enim eum dicentem quoniam Iesus Nazarenus hic destruet locum istum et mutabit consuetudines, quas tradidit nobis Moyses ".
ACTS|6|15|Et intuentes eum omnes, qui sedebant in concilio, viderunt faciem eius tamquam faciem angeli.
ACTS|7|1|Dixit autem princeps sacerdo tum: " Si haec ita se habent? ".
ACTS|7|2|Qui ait: " Viri fratres et patres, audite. Deus gloriae apparuit patri nostro Abraham, cum esset in Mesopotamia, priusquam moraretur in Charran,
ACTS|7|3|et dixit ad illum: "Exi de terra tua et de cognatione tua et veni in terram, quam tibi monstravero".
ACTS|7|4|Tunc egressus de terra Chaldaeorum habitavit in Charran. Et inde, postquam mortuus est pater eius, transtulit illum in terram istam, in qua nunc vos habitatis;
ACTS|7|5|et non dedit illi hereditatem in ea nec passum pedis et repromisit dare illi eam in possessionem et semini eius post ipsum, cum non haberet filium.
ACTS|7|6|Locutus est autem sic Deus: "Erit semen eius accola in terra aliena, et servituti eos subicient et male tractabunt annis quadringentis;
ACTS|7|7|et gentem, cui servierint, iudicabo ego, dixit Deus; et post haec exibunt et deservient mihi in loco isto".
ACTS|7|8|Et dedit illi testamentum circumcisionis; et sic genuit Isaac et circumcidit eum die octava, et Isaac Iacob, et Iacob duodecim patriarchas.
ACTS|7|9|Et patriarchae aemulantes Ioseph vendiderunt in Aegyptum; et erat Deus cum eo
ACTS|7|10|et eripuit eum ex omnibus tribulationibus eius et dedit ei gratiam et sapientiam in conspectu pharaonis regis Aegypti; et constituit eum praepositum super Aegyptum et super omnem domum suam.
ACTS|7|11|Venit autem fames in universam Aegyptum et Chanaan et tribulatio magna, et non inveniebant cibos patres nostri.
ACTS|7|12|Cum audisset autem Iacob esse frumentum in Aegypto, misit patres nostros primum;
ACTS|7|13|et in secundo cognitus est Ioseph a fratribus suis, et manifestatum est pharaoni genus Ioseph.
ACTS|7|14|Mittens autem Ioseph accersivit Iacob patrem suum et omnem cognationem in animabus septuaginta quinque;
ACTS|7|15|et descendit Iacob in Aegyptum. Et defunctus est ipse et patres nostri;
ACTS|7|16|et translati sunt in Sichem et positi sunt in sepulcro, quod emit Abraham pretio argenti a filiis Hemmor in Sichem.
ACTS|7|17|Cum appropinquaret autem tempus repromissionis, quam confessus erat Deus Abrahae, crevit populus et multiplicatus est in Aegypto,
ACTS|7|18|quoadusque surrexit rex alius super Aegypto, qui non sciebat Ioseph.
ACTS|7|19|Hic circumveniens genus nostrum, afflixit patres, ut exponerent infantes suos, ne vivi servarentur.
ACTS|7|20|Eodem tempore natus est Moyses et erat formosus coram Deo; qui nutritus est tribus mensibus in domo patris.
ACTS|7|21|Exposito autem illo, sustulit eum filia pharaonis et enutrivit eum sibi in filium;
ACTS|7|22|et eruditus est Moyses in omni sapientia Aegyptiorum; et erat potens in verbis et in operibus suis.
ACTS|7|23|Cum autem impleretur ei quadraginta annorum tempus, ascendit in cor eius, ut visitaret fratres suos filios Israel.
ACTS|7|24|Et cum vidisset quendam iniuriam patientem, vindicavit et fecit ultionem ei, qui opprimebatur, percusso Aegyptio.
ACTS|7|25|Existimabat autem intellegere fratres, quoniam Deus per manum ipsius daret salutem illis; at illi non intellexerunt.
ACTS|7|26|Atque sequenti die apparuit illis litigantibus et reconciliabat eos in pacem dicens: "Viri, fratres estis; ut quid nocetis alterutrum?".
ACTS|7|27|Qui autem iniuriam faciebat proximo, reppulit eum dicens: "Quis te constituit principem et iudicem super nos?
ACTS|7|28|Numquid interficere me tu vis, quemadmodum interfecisti heri Aegyptium?".
ACTS|7|29|Fugit autem Moyses propter verbum istud; et factus est advena in terra Madian, ubi generavit filios duos.
ACTS|7|30|Et expletis annis quadraginta, apparuit illi in deserto montis Sinai angelus in ignis flamma rubi.
ACTS|7|31|Moyses autem videns admirabatur visum; accedente autem illo, ut consideraret, facta est vox Domini:
ACTS|7|32|"Ego Deus patrum tuorum, Deus Abraham et Isaac et Iacob". Tremefactus autem Moyses non audebat considerare.
ACTS|7|33|Dixit autem illi Dominus: "Solve calceamentum pedum tuorum; locus enim, in quo stas, terra sancta est.
ACTS|7|34|Videns vidi afflictionem populi mei, qui est in Aegypto, et gemitum eorum audivi et descendi liberare eos; et nunc veni, mittam te in Aegyptum".
ACTS|7|35|Hunc Moysen, quem negaverunt dicentes: "Quis te constituit principem et iudicem?", hunc Deus et principem et redemptorem misit cum manu angeli, qui apparuit illi in rubo.
ACTS|7|36|Hic eduxit illos faciens prodigia et signa in terra Aegypti et in Rubro mari et in deserto annis quadraginta.
ACTS|7|37|Hic est Moyses, qui dixit filiis Israel: "Prophetam vobis suscitabit Deus de fratribus vestris tamquam me".
ACTS|7|38|Hic est qui fuit in ecclesia in solitudine cum angelo, qui loquebatur ei in monte Sinai, et cum patribus nostris; qui accepit verba viva dare nobis;
ACTS|7|39|cui noluerunt oboedire patres nostri, sed reppulerunt et aversi sunt in cordibus suis in Aegyptum
ACTS|7|40|dicentes ad Aaron: "Fac nobis deos, qui praecedant nos; Moyses enim hic, qui eduxit nos de terra Aegypti, nescimus quid factum sit ei".
ACTS|7|41|Et vitulum fecerunt in illis diebus et obtulerunt hostiam simulacro et laetabantur in operibus manuum suarum.
ACTS|7|42|Convertit autem Deus et tradidit eos servire militiae caeli, sicut scriptum est in libro Prophetarum:Numquid victimas et hostias obtulistis mihiannis quadraginta in deserto, domus Israel?
ACTS|7|43|Et suscepistis tabernaculum Molochet sidus dei vestri Rhaephan,figuras, quas fecistis ad adorandum eas.Et transferam vos trans Babylonem".
ACTS|7|44|Tabernaculum testimonii erat patribus nostris in deserto, sicut disposuit, qui loquebatur ad Moysen, ut faceret illud secundum formam, quam viderat;
ACTS|7|45|quod et induxerunt suscipientes patres nostri cum Iesu in possessionem gentium, quas expulit Deus a facie patrum nostrorum, usque in diebus David,
ACTS|7|46|qui invenit gratiam ante Deum et petiit, ut inveniret tabernaculum domui Iacob.
ACTS|7|47|Salomon autem aedificavit illi domum.
ACTS|7|48|Sed non Altissimus in manufactis habitat, sicut propheta dicit:
ACTS|7|49|"Caelum mihi thronus est,terra autem scabellum pedum meorum.Quam domum aedificabitis mihi, dicit Dominus,aut quis locus requietionis meae?
ACTS|7|50|Nonne manus mea fecit haec omnia?".
ACTS|7|51|Duri cervice et incircumcisi cordibus et auribus, vos semper Spiritui Sancto resistitis; sicut patres vestri, et vos.
ACTS|7|52|Quem prophetarum non sunt persecuti patres vestri? Et occiderunt eos, qui praenuntiabant de adventu Iusti, cuius vos nunc proditores et homicidae fuistis,
ACTS|7|53|qui accepistis legem in dispositionibus angelorum et non custodistis ".
ACTS|7|54|Audientes autem haec, dissecabantur cordibus suis et stridebant dentibus in eum.
ACTS|7|55|Cum autem esset plenus Spiritu Sancto, intendens in caelum vidit gloriam Dei et Iesum stantem a dextris Dei
ACTS|7|56|et ait: " Ecce video caelos apertos et Filium hominis a dextris stantem Dei ".
ACTS|7|57|Exclamantes autem voce magna continuerunt aures suas et impetum fecerunt unanimiter in eum
ACTS|7|58|et eicientes extra civitatem lapidabant. Et testes deposuerunt vestimenta sua secus pedes adulescentis, qui vocabatur Saulus.
ACTS|7|59|Et lapidabant Stephanum invocantem et dicentem: " Domine Iesu, suscipe spiritum meum ".
ACTS|7|60|Positis autem genibus clamavit voce magna: " Domine, ne statuas illis hoc peccatum "; et cum hoc dixisset, obdormivit.
ACTS|8|1|Saulus autem erat consentiens neci eius. Facta est autem in illa die persecutio magna in ecclesiam, quae erat Hierosolymis; et omnes dispersi sunt per regiones Iudaeae et Samariae praeter apostolos.
ACTS|8|2|Sepelierunt autem Stephanum viri timorati et fecerunt planctum magnum super illum.
ACTS|8|3|Saulus vero devastabat ecclesiam, per domos intrans et trahens viros ac mulieres tradebat in custodiam.
ACTS|8|4|Igitur qui dispersi erant, pertransierunt evangelizantes verbum.
ACTS|8|5|Philippus autem descendens in civitatem Samariae praedicabat illis Christum.
ACTS|8|6|Intendebant autem turbae his, quae a Philippo dicebantur, unanimiter, audientes et videntes signa, quae faciebat:
ACTS|8|7|ex multis enim eorum, qui habebant spiritus immundos, clamantes voce magna exibant; multi autem paralytici et claudi curati sunt.
ACTS|8|8|Factum est autem magnum gaudium in illa civitate.
ACTS|8|9|Vir autem quidam nomine Simon iampridem erat in civitate magias faciens et dementans gentem Samariae, dicens esse se aliquem magnum;
ACTS|8|10|cui attendebant omnes a minimo usque ad maximum dicentes: " Hic est virtus Dei, quae vocatur Magna ".
ACTS|8|11|Attendebant autem eum, propter quod multo tempore magiis dementasset eos.
ACTS|8|12|Cum vero credidissent Philippo evangelizanti de regno Dei et nomine Iesu Christi, baptizabantur viri ac mulieres.
ACTS|8|13|Tunc Simon et ipse credidit et, cum baptizatus esset, adhaerebat Philippo; videns etiam signa et virtutes magnas fieri stupens admirabatur.
ACTS|8|14|Cum autem audissent apostoli, qui erant Hierosolymis, quia recepit Samaria verbum Dei, miserunt ad illos Petrum et Ioannem;
ACTS|8|15|qui cum descendissent, oraverunt pro ipsis, ut acciperent Spiritum Sanctum:
ACTS|8|16|nondum enim super quemquam illorum venerat, sed baptizati tantum erant in nomine Domini Iesu.
ACTS|8|17|Tunc imposuerunt manus super illos, et accipiebant Spiritum Sanctum.
ACTS|8|18|Cum vidisset autem Simon quia per impositionem manuum apostolorum daretur Spiritus, obtulit eis pecuniam
ACTS|8|19|dicens: " Date et mihi hanc potestatem, ut cuicumque imposuero manus, accipiat Spiritum Sanctum ".
ACTS|8|20|Petrus autem dixit ad eum: " Argentum tuum tecum sit in perditionem, quoniam donum Dei existimasti pecunia possideri!
ACTS|8|21|Non est tibi pars neque sors in verbo isto; cor enim tuum non est rectum coram Deo.
ACTS|8|22|Paenitentiam itaque age ab hac nequitia tua et roga Dominum, si forte remittatur tibi haec cogitatio cordis tui;
ACTS|8|23|in felle enim amaritudinis et obligatione iniquitatis video te esse ".
ACTS|8|24|Respondens autem Simon dixit: " Precamini vos pro me ad Dominum, ut nihil veniat super me horum, quae dixistis ".
ACTS|8|25|Et illi quidem testificati et locuti verbum Domini, redibant Hierosolymam et multis vicis Samaritanorum evangelizabant.
ACTS|8|26|Angelus autem Domini locutus est ad Philippum dicens: " Surge et vade contra meridianum ad viam, quae descendit ab Ierusalem in Gazam; haec est deserta ".
ACTS|8|27|Et surgens abiit; et ecce vir Aethiops eunuchus potens Candacis reginae Aethiopum, qui erat super omnem gazam eius, qui venerat adorare in Ierusalem
ACTS|8|28|et revertebatur sedens super currum suum et legebat prophetam Isaiam.
ACTS|8|29|Dixit autem Spiritus Philippo: " Accede et adiunge te ad currum istum.
ACTS|8|30|Accurrens autem Philippus audivit illum legentem Isaiam prophetam et dixit: " Putasne intellegis, quae legis? ".
ACTS|8|31|Qui ait: " Et quomodo possum, si non aliquis ostenderit mihi? ". Rogavitque Philippum, ut ascenderet et sederet secum.
ACTS|8|32|Locus autem Scripturae, quem legebat, erat hic: Tamquam ovis ad occisionem ductus estet sicut agnus coram tondente se sine voce,sic non aperit os suum.
ACTS|8|33|In humilitate eius iudicium eius sublatum est.Generationem illius quis enarrabit?Quoniam tollitur de terra vita eius ".
ACTS|8|34|Respondens autem eunuchus Philippo dixit: " Obsecro te, de quo propheta dicit hoc? De se an de alio aliquo? ".
ACTS|8|35|Aperiens autem Philippus os suum et incipiens a Scriptura ista, evangelizavit illi Iesum.
ACTS|8|36|Et dum irent per viam, venerunt ad quandam aquam; et ait eunuchus: " Ecce aqua; quid prohibet me baptizari? ".
ACTS|8|37|()
ACTS|8|38|Et iussit stare currum; et descenderunt uterque in aquam Philippus et eunuchus, et baptizavit eum.
ACTS|8|39|Cum autem ascendissent de aqua, Spiritus Domini rapuit Philippum, et amplius non vidit eum eunuchus; ibat autem per viam suam gaudens.
ACTS|8|40|Philippus autem inventus est in Azoto et pertransiens evangelizabat civitatibus cunctis, donec veniret Caesaream.
ACTS|9|1|Saulus autem, adhuc spirans minarum et caedis in discipulos Domini, accessit ad principem sacerdotum
ACTS|9|2|et petiit ab eo epistulas in Damascum ad synagogas, ut, si quos invenisset huius viae viros ac mulieres, vinctos perduceret in Ierusalem.
ACTS|9|3|Et cum iter faceret, contigit ut appropinquaret Damasco; et subito circumfulsit eum lux de caelo,
ACTS|9|4|et cadens in terram audivit vocem dicentem sibi: " Saul, Saul, quid me persequeris? ".
ACTS|9|5|Qui dixit: " Quis es, Domine? ". Et ille: " Ego sum Iesus, quem tu persequeris!
ACTS|9|6|Sed surge et ingredere civitatem, et dicetur tibi quid te oporteat facere ".
ACTS|9|7|Viri autem illi, qui comitabantur cum eo, stabant stupefacti, audientes quidem vocem, neminem autem videntes.
ACTS|9|8|Surrexit autem Saulus de terra; apertisque oculis, nihil videbat; ad manus autem illum trahentes introduxerunt Damascum.
ACTS|9|9|Et erat tribus diebus non videns et non manducavit neque bibit.
ACTS|9|10|Erat autem quidam discipulus Damasci nomine Ananias; et dixit ad illum in visu Dominus: " Anania ". At ille ait: " Ecce ego, Domine ".
ACTS|9|11|Et Dominus ad illum: " Surgens vade in vicum, qui vocatur Rectus, et quaere in domo Iudae Saulum nomine Tarsensem; ecce enim orat
ACTS|9|12|et vidit virum Ananiam nomine introeuntem et imponentem sibi manus, ut visum recipiat ".
ACTS|9|13|Respondit autem Ananias: " Domine, audivi a multis de viro hoc, quanta mala sanctis tuis fecerit in Ierusalem;
ACTS|9|14|et hic habet potestatem a principibus sacerdotum alligandi omnes, qui invocant nomen tuum ".
ACTS|9|15|Dixit autem ad eum Dominus: " Vade, quoniam vas electionis est mihi iste, ut portet nomen meum coram gentibus et regibus et filiis Israel;
ACTS|9|16|ego enim ostendam illi quanta oporteat eum pro nomine meo pati ".
ACTS|9|17|Et abiit Ananias; et introivit in domum et imponens ei manus dixit: " Saul frater, Dominus misit me, Iesus qui apparuit tibi in via, qua veniebas, ut videas et implearis Spiritu Sancto ".
ACTS|9|18|Et confestim ceciderunt ab oculis eius tamquam squamae, et visum recepit. Et surgens baptizatus est
ACTS|9|19|et, cum accepisset cibum, confortatus est.Fuit autem cum discipulis, qui erant Damasci, per dies aliquot;
ACTS|9|20|et continuo in synagogis praedicabat Iesum, quoniam hic est Filius Dei.
ACTS|9|21|Stupebant autem omnes, qui audiebant, et dicebant: " Nonne hic est, qui expugnabat in Ierusalem eos, qui invocabant nomen istud, et huc ad hoc venerat, ut vinctos illos duceret ad principes sacerdotum? ".
ACTS|9|22|Saulus autem magis convalescebat et confundebat Iudaeos, qui habitabant Damasci, affirmans quoniam hic est Christus.
ACTS|9|23|Cum implerentur autem dies multi, consilium fecerunt Iudaei, ut eum interficerent;
ACTS|9|24|notae autem factae sunt Saulo insidiae eorum. Custodiebant autem et portas die ac nocte, ut eum interficerent;
ACTS|9|25|accipientes autem discipuli eius nocte per murum dimiserunt eum submittentes in sporta.
ACTS|9|26|Cum autem venisset in Ierusalem, tentabat iungere se discipulis; et omnes timebant eum, non credentes quia esset discipulus.
ACTS|9|27|Barnabas autem apprehensum illum duxit ad apostolos et narravit illis quomodo in via vidisset Dominum, et quia locutus est ei, et quomodo in Damasco fiducialiter egerit in nomine Iesu.
ACTS|9|28|Et erat cum illis intrans et exiens in Ierusalem, fiducialiter agens in nomine Domini.
ACTS|9|29|Loquebatur quoque et disputabat cum Graecis; illi autem quaerebant occidere eum.
ACTS|9|30|Quod cum cognovissent, fratres deduxerunt eum Caesaream et dimiserunt Tarsum.
ACTS|9|31|Ecclesia quidem per totam Iudaeam et Galilaeam et Samariam habebat pacem; aedificabatur et ambulabat in timore Domini et consolatione Sancti Spiritus crescebat.
ACTS|9|32|Factum est autem Petrum, dum pertransiret universos, devenire et ad sanctos, qui habitabant Lyddae.
ACTS|9|33|Invenit autem ibi hominem quendam nomine Aeneam ab annis octo iacentem in grabato, qui erat paralyticus.
ACTS|9|34|Et ait illi Petrus: " Aenea, sanat te Iesus Christus; surge et sterne tibi ". Et continuo surrexit.
ACTS|9|35|Et viderunt illum omnes, qui inhabitabant Lyddam et Saron, qui conversi sunt ad Dominum.
ACTS|9|36|In Ioppe autem erat quaedam discipula nomine Tabitha, quae interpretata dicitur Dorcas; haec erat plena operibus bonis et eleemosynis, quas faciebat.
ACTS|9|37|Factum est autem in diebus illis ut infirmata moreretur; quam cum lavissent, posuerunt in cenaculo.
ACTS|9|38|Cum autem prope esset Lydda ab Ioppe, discipuli audientes quia Petrus esset in ea, miserunt duos viros ad eum rogantes: " Ne pigriteris venire usque ad nos! ".
ACTS|9|39|Exsurgens autem Petrus venit cum illis; et cum advenisset, duxerunt illum in cenaculum; et circumsteterunt illum omnes viduae flentes et ostendentes tunicas et vestes, quas faciebat Dorcas, cum esset cum illis.
ACTS|9|40|Eiectis autem omnibus foras Petrus, et ponens genua oravit et conversus ad corpus dixit: " Tabitha, surge! ". At illa aperuit oculos suos et, viso Petro, resedit.
ACTS|9|41|Dans autem illi manum erexit eam et, cum vocasset sanctos et viduas, exhibuit eam vivam.
ACTS|9|42|Notum autem factum est per universam Ioppen, et crediderunt multi in Domino.
ACTS|9|43|Factum est autem, ut dies multos moraretur in Ioppe apud quendam Simonem coriarium.
ACTS|10|1|Vir autem quidam in Cae sarea nomine Cornelius, cen turio cohortis, quae dicitur Italica,
ACTS|10|2|religiosus et timens Deum cum omni domo sua, faciens eleemosynas multas plebi et deprecans Deum semper,
ACTS|10|3|vidit in visu manifeste quasi hora nona diei angelum Dei introeuntem ad se et dicentem sibi: " Corneli ".
ACTS|10|4|At ille intuens eum et timore correptus dixit: " Quid est, domine? ". Dixit autem illi: " Orationes tuae et eleemosynae tuae ascenderunt in memoriam in conspectu Dei.
ACTS|10|5|Et nunc mitte viros in Ioppen et accersi Simonem quendam, qui cognominatur Petrus;
ACTS|10|6|hic hospitatur apud Simonem quendam coriarium, cui est domus iuxta mare.
ACTS|10|7|Ut autem discessit angelus, qui loquebatur illi, cum vocasset duos domesticos suos et militem religiosum ex his, qui illi parebant,
ACTS|10|8|et narrasset illis omnia, misit illos in Ioppen.
ACTS|10|9|Postera autem die, iter illis facientibus et appropinquantibus civitati, ascendit Petrus super tectum, ut oraret circa horam sextam.
ACTS|10|10|Et cum esuriret, voluit gustare; parantibus autem eis, cecidit super eum mentis excessus,
ACTS|10|11|et videt caelum apertum et descendens vas quoddam velut linteum magnum quattuor initiis submitti in terram,
ACTS|10|12|in quo erant omnia quadrupedia et serpentia terrae et volatilia caeli.
ACTS|10|13|Et facta est vox ad eum: " Surge, Petre, occide et manduca! ".
ACTS|10|14|Ait autem Petrus: " Nequaquam, Domine, quia numquam manducavi omne commune et immundum ".
ACTS|10|15|Et vox iterum secundo ad eum: " Quae Deus purificavit, ne tu commune dixeris ".
ACTS|10|16|Hoc autem factum est per ter, et statim receptum est vas in caelum.
ACTS|10|17|Et dum intra se haesitaret Petrus quidnam esset visio, quam vidisset, ecce viri, qui missi erant a Cornelio, inquirentes domum Simonis astiterunt ad ianuam
ACTS|10|18|et, cum vocassent, interrogabant si Simon, qui cognominatur Petrus, illic haberet hospitium.
ACTS|10|19|Petro autem cogitante de visione, dixit Spiritus ei: " Ecce viri tres quaerunt te;
ACTS|10|20|surge itaque et descende et vade cum eis nihil dubitans, quia ego misi illos ".
ACTS|10|21|Descendens autem Petrus ad viros dixit: " Ecce ego sum, quem quaeritis; quae causa est, propter quam venistis? ".
ACTS|10|22|Qui dixerunt: " Cornelius centurio, vir iustus et timens Deum et testimonium habens ab universa gente Iudaeorum, responsum accepit ab angelo sancto accersire te in domum suam et audire verba abs te ".
ACTS|10|23|Invitans igitur eos recepit hospitio.Sequenti autem die, surgens profectus est cum eis, et quidam ex fratribus ab Ioppe comitati sunt eum.
ACTS|10|24|Altera autem die introivit Caesaream; Cornelius vero exspectabat illos, convocatis cognatis suis et necessariis amicis.
ACTS|10|25|Et factum est, cum introisset Petrus, obvius ei Cornelius procidens ad pedes adoravit.
ACTS|10|26|Petrus vero levavit eum dicens: " Surge, et ego ipse homo sum ".
ACTS|10|27|Et loquens cum illo intravit et invenit multos, qui convenerant;
ACTS|10|28|dixitque ad illos: " Vos scitis quomodo illicitum sit viro Iudaeo coniungi aut accedere ad alienigenam. Et mihi ostendit Deus neminem communem aut immundum dicere hominem;
ACTS|10|29|propter quod sine dubitatione veni accersitus. Interrogo ergo quam ob causam accersistis me ".
ACTS|10|30|Et Cornelius ait: " A nudius quarta die usque in hanc horam orans eram hora nona in domo mea, et ecce vir stetit ante me in veste candida
ACTS|10|31|et ait: "Corneli, exaudita est oratio tua, et eleemosynae tuae commemoratae sunt in conspectu Dei.
ACTS|10|32|Mitte ergo in Ioppen et accersi Simonem, qui cognominatur Petrus; hic hospitatur in domo Simonis coriarii iuxta mare".
ACTS|10|33|Confestim igitur misi ad te, et tu bene fecisti veniendo. Nunc ergo omnes nos in conspectu Dei adsumus audire omnia, quaecumque tibi praecepta sunt a Domino ".
ACTS|10|34|Aperiens autem Petrus os dixit: " In veritate comperio quoniam non est personarum acceptor Deus,
ACTS|10|35|sed in omni gente, qui timet eum et operatur iustitiam, acceptus est illi.
ACTS|10|36|Verbum misit filiis Israel evangelizans pacem per Iesum Christum; hic est omnium Dominus.
ACTS|10|37|Vos scitis quod factum est verbum per universam Iudaeam incipiens a Galilaea post baptismum, quod praedicavit Ioannes:
ACTS|10|38|Iesum a Nazareth, quomodo unxit eum Deus Spiritu Sancto et virtute, qui pertransivit benefaciendo et sanando omnes oppressos a Diabolo, quoniam Deus erat cum illo.
ACTS|10|39|Et nos testes sumus omnium, quae fecit in regione Iudaeorum et Ierusalem; quem et occiderunt suspendentes in ligno.
ACTS|10|40|Hunc Deus suscitavit tertia die et dedit eum manifestum fieri
ACTS|10|41|non omni populo, sed testibus praeordinatis a Deo, nobis, qui manducavimus et bibimus cum illo postquam resurrexit a mortuis;
ACTS|10|42|et praecepit nobis praedicare populo et testificari quia ipse est, qui constitutus est a Deo iudex vivorum et mortuorum.
ACTS|10|43|Huic omnes Prophetae testimonium perhibent remissionem peccatorum accipere per nomen eius omnes, qui credunt in eum ".
ACTS|10|44|Adhuc loquente Petro verba haec, cecidit Spiritus Sanctus super omnes, qui audiebant verbum.
ACTS|10|45|Et obstupuerunt, qui ex circumcisione fideles, qui venerant cum Petro, quia et in nationes gratia Spiritus Sancti effusa est;
ACTS|10|46|audiebant enim illos loquentes linguis et magnificantes Deum. Tunc respondit Petrus:
ACTS|10|47|" Numquid aquam quis prohibere potest, ut non baptizentur hi, qui Spiritum Sanctum acceperunt sicut et nos? ".
ACTS|10|48|Et iussit eos in nomine Iesu Christi baptizari. Tunc rogaverunt eum, ut maneret aliquot diebus.
ACTS|11|1|Audierunt autem apostoli et fratres, qui erant in Iudaea, quoniam et gentes receperunt verbum Dei.
ACTS|11|2|Cum ascendisset autem Petrus in Ierusalem, disceptabant adversus illum, qui erant ex circumcisione,
ACTS|11|3|dicentes: " Introisti ad viros praeputium habentes et manducasti cum illis! ".
ACTS|11|4|Incipiens autem Petrus exponebat illis ex ordine dicens:
ACTS|11|5|" Ego eram in civitate Ioppe orans et vidi in excessu mentis visionem, descendens vas quoddam velut linteum magnum quattuor initiis submitti de caelo et venit usque ad me;
ACTS|11|6|in quod intuens considerabam et vidi quadrupedia terrae et bestias et reptilia et volatilia caeli.
ACTS|11|7|Audivi autem et vocem dicentem mihi: "Surgens, Petre, occide et manduca!".
ACTS|11|8|Dixi autem: Nequaquam, Domine, quia commune aut immundum numquam introivit in os meum.
ACTS|11|9|Respondit autem vox secundo de caelo: "Quae Deus mundavit, tu ne commune dixeris".
ACTS|11|10|Hoc autem factum est per ter, et retracta sunt rursum omnia in caelum.
ACTS|11|11|Et ecce confestim tres viri astiterunt in domo, in qua eramus, missi a Caesarea ad me.
ACTS|11|12|Dixit autem Spiritus mihi, ut irem cum illis nihil haesitans. Venerunt autem mecum et sex fratres isti, et ingressi sumus in domum viri.
ACTS|11|13|Narravit autem nobis quomodo vidisset angelum ad domum suam stantem et dicentem: "Mitte in Ioppen et accersi Simonem, qui cognominatur Petrus,
ACTS|11|14|qui loquetur tibi verba, in quibus salvus eris tu et universa domus tua".
ACTS|11|15|Cum autem coepissem loqui, decidit Spiritus Sanctus super eos, sicut et super nos in initio.
ACTS|11|16|Recordatus sum autem verbi Domini, sicut dicebat: "Ioannes quidem baptizavit aqua, vos autem baptizabimini in Spiritu Sancto".
ACTS|11|17|Si ergo aequale donum dedit illis Deus sicut et nobis, qui credidimus in Dominum Iesum Christum, ego quis eram qui possem prohibere Deum? ".
ACTS|11|18|His autem auditis, acquieverunt et glorificaverunt Deum dicentes: " Ergo et gentibus Deus paenitentiam ad vitam dedit ".
ACTS|11|19|Et illi quidem, qui dispersi fuerant a tribulatione, quae facta fuerat sub Stephano, perambulaverunt usque Phoenicen et Cyprum et Antiochiam, nemini loquentes verbum; nisi solis Iudaeis.
ACTS|11|20|Erant autem quidam ex eis viri Cyprii et Cyrenaei, qui, cum introissent Antiochiam, loquebantur et ad Graecos evangelizantes Dominum Iesum.
ACTS|11|21|Et erat manus Domini cum eis; multusque numerus credentium conversus est ad Dominum.
ACTS|11|22|Auditus est autem sermo in auribus ecclesiae, quae erat in Ierusalem, super istis, et miserunt Barnabam usque Antiochiam;
ACTS|11|23|qui cum pervenisset et vidisset gratiam Dei, gavisus est et hortabatur omnes proposito cordis permanere in Domino,
ACTS|11|24|quia erat vir bonus et plenus Spiritu Sancto et fide. Et apposita est turba multa Domino.
ACTS|11|25|Profectus est autem Tarsum, ut quaereret Saulum;
ACTS|11|26|quem cum invenisset, perduxit Antiochiam. Factum est autem eis, ut annum totum conversarentur in ecclesia et docerent turbam multam, et cognominarentur primum Antiochiae discipuli Christiani.
ACTS|11|27|In his autem diebus supervenerunt ab Hierosolymis prophetae Antiochiam;
ACTS|11|28|et surgens unus ex eis nomine Agabus significavit per Spiritum famem magnam futuram in universo orbe terrarum; quae facta est sub Claudio.
ACTS|11|29|Discipuli autem, prout quis habebat, proposuerunt singuli eorum in ministerium mittere habitantibus in Iudaea fratribus;
ACTS|11|30|quod et fecerunt, mittentes ad presbyteros per manum Barnabae et Sauli.
ACTS|12|1|Illo autem tempore, misit Herodes rex manus, ut affli geret quosdam de ecclesia.
ACTS|12|2|Occidit autem Iacobum fratrem Ioannis gladio.
ACTS|12|3|Videns autem quia placeret Iudaeis, apposuit apprehendere et Petrum - erant autem dies Azymorum -
ACTS|12|4|quem cum apprehendisset, misit in carcerem tradens quattuor quaternionibus militum custodire eum, volens post Pascha producere eum populo.
ACTS|12|5|Et Petrus quidem servabatur in carcere; oratio autem fiebat sine intermissione ab ecclesia ad Deum pro eo.
ACTS|12|6|Cum autem producturus eum esset Herodes, in ipsa nocte erat Petrus dormiens inter duos milites vinctus catenis duabus, et custodes ante ostium custodiebant carcerem.
ACTS|12|7|Et ecce angelus Domini astitit, et lumen refulsit in habitaculo; percusso autem latere Petri, suscitavit eum dicens: " Surge velociter! ". Et ceciderunt catenae de manibus eius.
ACTS|12|8|Dixit autem angelus ad eum: " Praecingere et calcea te sandalia tua! ". Et fecit sic. Et dicit illi: " Circumda tibi vestimentum tuum et sequere me! ".
ACTS|12|9|Et exiens sequebatur et nesciebat quia verum est, quod fiebat per angelum; aestimabat autem se visum videre.
ACTS|12|10|Transeuntes autem primam custodiam et secundam venerunt ad portam ferream, quae ducit ad civitatem, quae ultro aperta est eis, et exeuntes processerunt vicum unum, et continuo discessit angelus ab eo.
ACTS|12|11|Et Petrus ad se reversus dixit: " Nunc scio vere quia misit Dominus angelum suum et eripuit me de manu Herodis et de omni exspectatione plebis Iudaeorum ".
ACTS|12|12|Consideransque venit ad domum Mariae matris Ioannis, qui cognominatur Marcus, ubi erant multi congregati et orantes.
ACTS|12|13|Pulsante autem eo ostium ianuae, processit puella ad audiendum, nomine Rhode;
ACTS|12|14|et ut cognovit vocem Petri, prae gaudio non aperuit ianuam, sed intro currens nuntiavit stare Petrum ante ianuam.
ACTS|12|15|At illi dixerunt ad eam: " Insanis! ". Illa autem affirmabat sic se habere. Illi autem dicebant: " Angelus eius est ".
ACTS|12|16|Petrus autem perseverabat pulsans; cum autem aperuissent, viderunt eum et obstupuerunt.
ACTS|12|17|Annuens autem eis manu, ut tacerent, enarravit quomodo Dominus eduxisset eum de carcere dixitque: " Nuntiate Iacobo ct fratribus haec ". Et egressus abiit in alium locum.
ACTS|12|18|Facta autem die, erat non parva turbatio inter milites, quidnam de Petro factum esset.
ACTS|12|19|Herodes autem, cum requisisset eum et non invenisset, interrogatis custodibus, iussit eos abduci; descendensque a Iudaea in Caesaream ibi commorabatur.
ACTS|12|20|Erat autem iratus Tyriis et Sidoniis; at illi unanimes venerunt ad eum et, persuaso Blasto, qui erat super cubiculum regis, postulabant pacem, eo quod aleretur regio eorum ab annona regis.
ACTS|12|21|Statuto autem die, Herodes, vestitus veste regia, sedens pro tribunalicontionabatur ad eos;
ACTS|12|22|populus autem acclamabat: " Dei vox et non hominis! ".
ACTS|12|23|Confestim autem percussit eum angelus Domini, eo quod non dedisset gloriam Deo; et consumptus a vermibus exspiravit.
ACTS|12|24|Verbum autem Dei crescebat et multiplicabatur.
ACTS|12|25|Barnabas autem et Saulus reversi sunt in Ierusalem expleto ministerio, assumpto Ioanne, qui cognominatus est Marcus.
ACTS|13|1|Erant autem in ecclesia, quae erat Antiochiae, pro phetae et doctores: Barnabas et Simeon, qui vocabatur Niger, et Lucius Cyrenensis et Manaen, qui erat Herodis tetrarchae collactaneus, et Saulus.
ACTS|13|2|Ministrantibus autem illis Domino et ieiunantibus, dixit Spiritus Sanctus: " Separate mihi Barnabam et Saulum in opus, ad quod vocavi eos ".
ACTS|13|3|Tunc ieiunantes et orantes imponentesque eis manus dimiserunt illos.
ACTS|13|4|Et ipsi quidem missi ab Spiritu Sancto devenerunt Seleuciam et inde navigaverunt Cyprum
ACTS|13|5|et, cum venissent Salamina, praedicabant verbum Dei in synagogis Iudaeorum; habebant autem et Ioannem ministrum.
ACTS|13|6|Et cum perambulassent universam insulam usque Paphum, invenerunt quendam virum magum pseudoprophetam Iudaeum, cui nomen Bariesu,
ACTS|13|7|qui erat cum proconsule Sergio Paulo, viro prudente. Hic, accitis Barnaba et Saulo, quaesivit audire verbum Dei;
ACTS|13|8|resistebat autem illis Elymas, magus, sic enim interpretatur nomen eius, quaerens avertere proconsulem a fide.
ACTS|13|9|Saulus autem, qui et Paulus, repletus Spiritu Sancto, intuens in eum
ACTS|13|10|dixit: " O plene omni dolo et omni fallacia, fili Diaboli, inimice omnis iustitiae, non desines subvertere vias Domini rectas?
ACTS|13|11|Et nunc, ecce manus Domini super te; et eris caecus, non videns solem usque ad tempus ". Et confestim cecidit in eum caligo et tenebrae, et circumiens quaerebat, qui eum manum darent.
ACTS|13|12|Tunc proconsul, cum vidisset factum, credidit admirans super doctrinam Domini.
ACTS|13|13|Et cum a Papho navigassent, qui erant cum Paulo, venerunt Pergen Pamphyliae; Ioannes autem discedens ab eis reversus est Hierosolymam.
ACTS|13|14|Illi vero pertranseuntes, a Perge venerunt Antiochiam Pisidiae, et ingressi synagogam die sabbatorum sederunt.
ACTS|13|15|Post lectionem autem Legis et Prophetarum, miserunt principes synagogae ad eos dicentes: " Viri fratres, si quis est in vobis sermo exhortationis ad plebem, dicite! ".
ACTS|13|16|Surgens autem Paulus et manu silentium indicens ait: " Viri Israelitae et qui timetis Deum, audite.
ACTS|13|17|Deus plebis huius Israel elegit patres nostros et plebem exaltavit, cum essent incolae in terra Aegypti, et in brachio excelso eduxit eos ex ea;
ACTS|13|18|et per quadraginta fere annorum tempus mores eorum sustinuit in deserto;
ACTS|13|19|et destruens gentes septem in terra Chanaan sorte distribuit terram eorum,
ACTS|13|20|quasi quadringentos et quinquaginta annos. Et post haec dedit iudices usque ad Samuel prophetam.
ACTS|13|21|Et exinde postulaverunt regem, et dedit illis Deus Saul filium Cis, virum de tribu Beniamin, annis quadraginta.
ACTS|13|22|Et amoto illo, suscitavit illis David in regem, cui et testimonium perhibens dixit: "Inveni David filium Iesse, virum secundum cor meum, qui faciet omnes voluntates meas".
ACTS|13|23|Huius Deus ex semine secundum promissionem eduxit Israel salvatorem Iesum,
ACTS|13|24|praedicante Ioanne ante adventum eius baptismum paenitentiae omni populo Israel.
ACTS|13|25|Cum impleret autem Ioannes cursum suum, dicebat: "Quid me arbitramini esse? Non sum ego; sed ecce venit post me, cuius non sum dignus calceamenta pedum solvere".
ACTS|13|26|Viri fratres, filii generis Abraham et qui in vobis timent Deum, nobis verbum salutis huius missum est.
ACTS|13|27|Qui enim habitabant Ierusalem et principes eorum, hunc ignorantes et voces Prophetarum, quae per omne sabbatum leguntur, iudicantes impleverunt;
ACTS|13|28|et nullam causam mortis invenientes petierunt a Pilato, ut interficeretur;
ACTS|13|29|cumque consummassent omnia, quae de eo scripta erant, deponentes eum de ligno posuerunt in monumento.
ACTS|13|30|Deus vero suscitavit eum a mortuis;
ACTS|13|31|qui visus est per dies multos his, qui simul ascenderant cum eo de Galilaea in Ierusalem, qui nunc sunt testes eius ad plebem.
ACTS|13|32|Et nos vobis evangelizamus eam, quae ad patres promissio facta est,
ACTS|13|33|quoniam hanc Deus adimplevit filiis eorum, nobis resuscitans Iesum, sicut et in Psalmo secundo scriptum est:Filius meus es tu; ego hodie genui te".
ACTS|13|34|Quod autem suscitaverit eum a mortuis, amplius iam non reversurum in corruptionem, ita dixit: "Dabo vobis sancta David fidelia".
ACTS|13|35|Ideoque et in alio dicit:Non dabis Sanctum tuum videre corruptionem".
ACTS|13|36|David enim sua generatione cum administrasset voluntati Dei, dormivit et appositus est ad patres suos et vidit corruptionem;
ACTS|13|37|quem vero Deus suscitavit, non vidit corruptionem.
ACTS|13|38|Notum igitur sit vobis, viri fratres, quia per hunc vobis remissio peccatorum annuntiatur; ab omnibus, quibus non potuistis in lege Moysi iustificari,
ACTS|13|39|in hoc omnis, qui credit, iustificatur.
ACTS|13|40|Videte ergo, ne superveniat, quod dictum est in Prophetis:
ACTS|13|41|"Videte, contemptores,et admiramini et disperdimini,quia opus operor ego in diebus vestris,opus, quod non credetis, si quis enarraverit vobis!" ".
ACTS|13|42|Exeuntibus autem illis, rogabant, ut sequenti sabbato loquerentur sibi verba haec.
ACTS|13|43|Cumque dimissa esset synagoga, secuti sunt multi Iudaeorum et colentium proselytorum Paulum et Barnabam, qui loquentes suadebant eis, ut permanerent in gratia Dei.
ACTS|13|44|Sequenti vero sabbato paene universa civitas convenit audire verbum Domini.
ACTS|13|45|Videntes autem turbas Iudaei, repleti sunt zelo; et contradicebant his, quae a Paulo dicebantur, blasphemantes.
ACTS|13|46|Tunc audenter Paulus et Barnabas dixerunt: " Vobis oportebat primum loqui verbum Dei; sed quoniam repellitis illud et indignos vos iudicatis aeternae vitae, ecce convertimur ad gentes.
ACTS|13|47|Sic enim praecepit nobis Dominus:Posui te in lumen gentium,ut sis in salutem usque ad extremum terrae" ".
ACTS|13|48|Audientes autem gentes gaudebant et glorificabant verbum Domini, et crediderunt, quotquot erant praeordinati ad vitam aeternam;
ACTS|13|49|ferebatur autem verbum Domini per universam regionem.
ACTS|13|50|Iudaei autem concitaverunt honestas inter colentes mulieres et primos civitatis et excitaverunt persecutionem in Paulum et Barnabam et eiecerunt eos de finibus suis.
ACTS|13|51|At illi, excusso pulvere pedum in eos, venerunt Iconium;
ACTS|13|52|discipuli quoque replebantur gaudio et Spiritu Sancto.
ACTS|14|1|Factum est autem Iconii, ut eodem modo introirent syna gogam Iudaeorum et ita loquerentur, ut crederet Iudaeorum et Graecorum copiosa multitudo.
ACTS|14|2|Qui vero increduli fuerunt Iudaei, suscitaverunt et exacerbaverunt animas gentium adversus fratres.
ACTS|14|3|Multo igitur tempore demorati sunt, fiducialiter agentes in Domino, testimonium perhibente verbo gratiae suae, dante signa et prodigia fieri per manus eorum.
ACTS|14|4|Divisa est autem multitudo civitatis: et quidam quidem erant cum Iudaeis, quidam vero cum apostolis.
ACTS|14|5|Cum autem factus esset impetus gentilium et Iudaeorum cum principibus suis, ut contumeliis afficerent et lapidarent eos,
ACTS|14|6|intellegentes confugerunt ad civitates Lycaoniae, Lystram et Derben et ad regionem in circuitu
ACTS|14|7|et ibi evangelizantes erant.
ACTS|14|8|Et quidam vir in Lystris infirmus pedibus sedebat, claudus ex utero matris suae, qui numquam ambulaverat.
ACTS|14|9|Hic audivit Paulum loquentem; qui intuitus eum et videns quia haberet fidem, ut salvus fieret,
ACTS|14|10|dixit magna voce: " Surge super pedes tuos rectus! ". Et exsilivit et ambulabat.
ACTS|14|11|Turbae autem cum vidissent, quod fecerat Paulus, levaverunt vocem suam Lycaonice dicentes: " Dii similes facti hominibus descenderunt ad nos! ";
ACTS|14|12|et vocabant Barnabam Iovem, Paulum vero Mercurium, quoniam ipse erat dux verbi.
ACTS|14|13|Sacerdos quoque templi Iovis, quod erat ante civitatem, tauros et coronas ad ianuas afferens cum populis, volebat sacrificare.
ACTS|14|14|Quod ubi audierunt apostoli Barnabas et Paulus, conscissis tunicis suis, exsilierunt in turbam clamantes
ACTS|14|15|et dicentes: " Viri, quid haec facitis? Et nos mortales sumus similes vobis homines, evangelizantes vobis ab his vanis converti ad Deum vivum, qui fecit caelum et terram et mare et omnia, quae in eis sunt.
ACTS|14|16|Qui in praeteritis generationibus permisit omnes gentes ambulare in viis suis;
ACTS|14|17|et quidem non sine testimonio semetipsum reliquit benefaciens, de caelo dans vobis pluvias et tempora fructifera, implens cibo et laetitia corda vestra ".
ACTS|14|18|Et haec dicentes vix sedaverunt turbas, ne sibi immolarent.
ACTS|14|19|Supervenerunt autem ab Antiochia et Iconio Iudaei et persuasis turbis lapidantesque Paulum trahebant extra civitatem aestimantes eum mortuum esse.
ACTS|14|20|Circumdantibus autem eum discipulis, surgens intravit civitatem. Et postera die profectus est cum Barnaba in Derben.
ACTS|14|21|Cumque evangelizassent civitati illi et docuissent multos, reversi sunt Lystram et Iconium et Antiochiam
ACTS|14|22|confirmantes animas discipulorum, exhortantes, ut permanerent in fide, et quoniam per multas tribulationes oportet nos intrare in regnum Dei.
ACTS|14|23|Et cum ordinassent illis per singulas ecclesias presbyteros et orassent cum ieiunationibus, commendaverunt eos Domino, in quem crediderant.
ACTS|14|24|Transeuntesque Pisidiam venerunt Pamphyliam;
ACTS|14|25|et loquentes in Perge verbum descenderunt in Attaliam.
ACTS|14|26|Et inde navigaverunt Antiochiam, unde erant traditi gratiae Dei in opus, quod compleverunt.
ACTS|14|27|Cum autem venissent et congregassent ecclesiam, rettulerunt quanta fecisset Deus cum illis et quia aperuisset gentibus ostium fidei.
ACTS|14|28|Morati sunt autem tempus non modicum cum discipulis.
ACTS|15|1|Et quidam descendentes de Iudaea docebant fratres: " Nisi circumcidamini secundum morem Moysis, non potestis salvi fieri ".
ACTS|15|2|Facta autem seditione et conquisitione non minima Paulo et Barnabae adversum illos, statuerunt, ut ascenderent Paulus et Barnabas et quidam alii ex illis ad apostolos et presbyteros in Ierusalem super hac quaestione.
ACTS|15|3|Illi igitur deducti ab ecclesia pertransiebant Phoenicen et Samariam narrantes conversionem gentium et faciebant gaudium magnum omnibus fratribus.
ACTS|15|4|Cum autem venissent Hierosolymam, suscepti sunt ab ecclesia et apostolis et presbyteris et annuntiaverunt quanta Deus fecisset cum illis.
ACTS|15|5|Surrexerunt autem quidam de haeresi pharisaeorum, qui crediderant, dicentes: " Oportet circumcidere eos, praecipere quoque servare legem Moysis! ".
ACTS|15|6|Conveneruntque apostoli et presbyteri videre de verbo hoc.
ACTS|15|7|Cum autem magna conquisitio fieret, surgens Petrus dixit ad eos: " Viri fratres, vos scitis quoniam ab antiquis diebus in vobis elegit Deus per os meum audire gentes verbum evangelii et credere;
ACTS|15|8|et qui novit corda, Deus, testimonium perhibuit illis dans Spiritum Sanctum sicut et nobis;
ACTS|15|9|et nihil discrevit inter nos et illos fide purificans corda eorum.
ACTS|15|10|Nunc ergo quid tentatis Deum imponere iugum super cervicem discipulorum, quod neque patres nostri neque nos portare potuimus?
ACTS|15|11|Sed per gratiam Domini Iesu credimus salvari quemadmodum et illi ".
ACTS|15|12|Tacuit autem omnis multitudo, et audiebant Barnabam et Paulum narrantes quanta fecisset Deus signa et prodigia in gentibus per eos.
ACTS|15|13|Et postquam tacuerunt, respondit Iacobus dicens: " Viri fratres, audite me.
ACTS|15|14|Simeon narravit quemadmodum primum Deus visitavit sumere ex gentibus populum nomini suo;
ACTS|15|15|et huic concordant verba Prophetarum, sicut scriptum est:
ACTS|15|16|"Post haec revertaret reaedificabo tabernaculum David, quod decidit,et diruta eius reaedificabo et erigam illud.
ACTS|15|17|ut requirant reliqui hominum Dominumet omnes gentes, super quas invocatum est nomen meum,dicit Dominus faciens haec
ACTS|15|18|nota a saeculo".
ACTS|15|19|Propter quod ego iudico non inquietari eos, qui ex gentibus convertuntur ad Deum,
ACTS|15|20|sed scribere ad eos, ut abstineant se a contaminationibus simulacrorum et fornicatione et suffocato et sanguine.
ACTS|15|21|Moyses enim a generationibus antiquis habet in singulis civitatibus, qui eum praedicent in synagogis, ubi per omne sabbatum legitur ".
ACTS|15|22|Tunc placuit apostolis et presbyteris cum omni ecclesia electos viros ex eis mittere Antiochiam cum Paulo et Barnaba: Iudam, qui cognominatur Barsabbas, et Silam, viros primos in fratribus,
ACTS|15|23|scribentes per manum eorum: " Apostoli et presbyteri fratres his, qui sunt Antiochiae et Syriae et Ciliciae, fratribus ex gentibus, salutem!
ACTS|15|24|Quoniam audivimus quia quidam ex nobis, quibus non mandavimus, exeuntes turbaverunt vos verbis evertentes animas vestras,
ACTS|15|25|placuit nobis collectis in unum eligere viros et mittere ad vos cum carissimis nobis Barnaba et Paulo,
ACTS|15|26|hominibus, qui tradiderunt animas suas pro nomine Domini nostri Iesu Christi.
ACTS|15|27|Misimus ergo Iudam et Silam, qui et ipsi verbis referent eadem.
ACTS|15|28|Visum est enim Spiritui Sancto et nobis nihil ultra imponere vobis oneris quam haec necessario:
ACTS|15|29|abstinere ab idolothytis et sanguine et suffocatis et fornicatione; a quibus custodientes vos bene agetis. Valete ".
ACTS|15|30|Illi igitur dimissi descenderunt Antiochiam et, congregata multitudine, tradiderunt epistulam;
ACTS|15|31|quam cum legissent, gavisi sunt super consolatione.
ACTS|15|32|Iudas quoque et Silas, cum et ipsi essent prophetae, verbo plurimo consolati sunt fratres et confirmaverunt.
ACTS|15|33|Facto autem tempore, dimissi sunt cum pace a fratribus ad eos, qui miserant illos.
ACTS|15|34|()
ACTS|15|35|Paulus autem et Barnabas demorabantur Antiochiae docentes et evangelizantes cum aliis pluribus verbum Domini.
ACTS|15|36|Post aliquot autem dies dixit ad Barnabam Paulus: " Revertentes visitemus fratres per universas civitates, in quibus praedicavimus verbum Domini, quomodo se habeant ".
ACTS|15|37|Barnabas autem volebat secum assumere et Ioannem, qui cognominatur Marcus;
ACTS|15|38|Paulus autem iudicabat eum, qui discessisset ab eis a Pamphylia et non isset cum eis in opus, non debere recipi eum.
ACTS|15|39|Facta est autem exacerbatio, ita ut discederent ab invicem, et Barnabas, assumpto Marco, navigaret Cyprum.
ACTS|15|40|Paulus vero, electo Sila, profectus est, traditus gratiae Domini a fratribus;
ACTS|15|41|perambulabat autem Syriam et Ciliciam confirmans ecclesias.
ACTS|16|1|Pervenit autem in Derben et Lystram. Et ecce discipulus quidam erat ibi nomine Timotheus, filius mulieris Iudaeae fidelis, patre autem Graeco;
ACTS|16|2|huic testimonium reddebant, qui in Lystris erant et Iconii fratres.
ACTS|16|3|Hunc voluit Paulus secum proficisci et assumens circumcidit eum propter Iudaeos, qui erant in illis locis; sciebant enim omnes quod pater eius Graecus esset.
ACTS|16|4|Cum autem pertransirent civitates, tradebant eis custodire dogmata, quae erant decreta ab apostolis et presbyteris, qui essent Hierosolymis.
ACTS|16|5|Ecclesiae quidem confirmabantur fide et abundabant numero cotidie.
ACTS|16|6|Transierunt autem Phrygiam et Galatiae regionem, vetati a Sancto Spiritu loqui verbum in Asia;
ACTS|16|7|cum venissent autem circa Mysiam, tentabant ire Bithyniam, et non permisit eos Spiritus Iesu;
ACTS|16|8|cum autem praeterissent Mysiam, descenderunt Troadem.
ACTS|16|9|Et visio per noctem Paulo ostensa est: vir Macedo quidam erat stans et deprecans eum et dicens: " Transiens in Macedoniam, adiuva nos! ".
ACTS|16|10|Ut autem visum vidit, statim quaesivimus proficisci in Macedoniam, certi facti quia vocasset nos Deus evangelizare eis.
ACTS|16|11|Navigantes autem a Troade recto cursu venimus Samothraciam et sequenti die Neapolim
ACTS|16|12|et inde Philippos, quae est prima partis Macedoniae civitas, colonia. Eramus autem in hac urbe diebus aliquot commorantes.
ACTS|16|13|Die autem sabbatorum egressi sumus foras portam iuxta flumen, ubi putabamus orationem esse, et sedentes loquebamur mulieribus, quae convenerant.
ACTS|16|14|Et quaedam mulier nomine Lydia, purpuraria civitatis Thyatirenorum colens Deum, audiebat, cuius Dominus aperuit cor intendere his, quae dicebantur a Paulo.
ACTS|16|15|Cum autem baptizata esset et domus eius, deprecata est dicens: " Si iudicastis me fidelem Domino esse, introite in domum meam et manete "; et coegit nos.
ACTS|16|16|Factum est autem, euntibus nobis ad orationem, puellam quandam habentem spiritum pythonem obviare nobis, quae quaestum magnum praestabat dominis suis divinando.
ACTS|16|17|Haec subsecuta Paulum et nos clamabat dicens: " Isti homines servi Dei Altissimi sunt, qui annuntiant vobis viam salutis ".
ACTS|16|18|Hoc autem faciebat multis diebus. Dolens autem Paulus et conversus spiritui dixit: " Praecipio tibi in nomine Iesu Christi exire ab ea "; et exiit eadem hora.
ACTS|16|19|Videntes autem domini eius quia exivit spes quaestus eorum, apprehendentes Paulum et Silam traxerunt in forum ad principes;
ACTS|16|20|et producentes eos magistratibus dixerunt: " Hi homines conturbant civitatem nostram, cum sint Iudaei,
ACTS|16|21|et annuntiant mores, quos non licet nobis suscipere neque facere, cum simus Romani ".
ACTS|16|22|Et concurrit plebs adversus eos; et magistratus, scissis tunicis eorum, iusserunt virgis caedi
ACTS|16|23|et, cum multas plagas eis imposuissent, miserunt eos in carcerem, praecipientes custodi, ut caute custodiret eos;
ACTS|16|24|qui cum tale praeceptum accepisset, misit eos in interiorem carcerem et pedes eorum strinxit in ligno.
ACTS|16|25|Media autem nocte, Paulus et Silas orantes laudabant Deum, et audiebant eos, qui in custodia erant;
ACTS|16|26|subito vero terraemotus factus est magnus, ita ut moverentur fundamenta carceris, et aperta sunt statim ostia omnia, et universorum vincula soluta sunt.
ACTS|16|27|Expergefactus autem custos carceris et videns apertas ianuas carceris, evaginato gladio volebat se interficere, aestimans fugisse vinctos.
ACTS|16|28|Clamavit autem Paulus magna voce dicens: " Nihil feceris tibi mali; universi enim hic sumus ".
ACTS|16|29|Petitoque lumine, intro cucurrit et tremefactus procidit Paulo et Silae;
ACTS|16|30|et producens eos foras ait: " Domini, quid me oportet facere, ut salvus fiam? ".
ACTS|16|31|At illi dixerunt: " Crede in Domino Iesu et salvus eris tu et domus tua.
ACTS|16|32|Et locuti sunt ei verbum Domini cum omnibus, qui erant in domo eius.
ACTS|16|33|Et tollens eos in illa hora noctis lavit eos a plagis, et baptizatus est ipse et omnes eius continuo;
ACTS|16|34|cumque perduxisset eos in domum, apposuit mensam et laetatus est cum omni domo sua credens Deo.
ACTS|16|35|Et cum dies factus esset, miserunt magistratus lictores dicentes: " Dimitte homines illos! ".
ACTS|16|36|Nuntiavit autem custos carceris verba haec Paulo: " Miserunt magistratus, ut dimittamini; nunc igitur exeuntes ite in pace ".
ACTS|16|37|Paulus autem dixit eis: " Caesos nos publice, indemnatos, cum homines Romani essemus, miserunt in carcerem; et nunc occulte nos eiciunt? Non ita, sed veniant et ipsi nos educant ".
ACTS|16|38|Nuntiaverunt autem magistratibus lictores verba haec. Timueruntque audito quod Romani essent;
ACTS|16|39|et venientes deprecati sunt eos et educentes rogabant, ut egrederentur urbem.
ACTS|16|40|Exeuntes autem de carcere introierunt ad Lydiam et, visis fratribus, consolati sunt eos et profecti sunt.
ACTS|17|1|Cum autem perambulassent Amphipolim et Apolloniam, venerunt Thessalonicam, ubi erat synagoga Iudaeorum.
ACTS|17|2|Secundum consuetudinem autem suam Paulus introivit ad eos et per sabbata tria disserebat eis de Scripturis
ACTS|17|3|adaperiens et comprobans quia Christum oportebat pati et resurgere a mortuis, et: " Hic est Christus, Iesus, quem ego annuntio vobis ".
ACTS|17|4|Et quidam ex eis crediderunt et adiuncti sunt Paulo et Silae et de colentibus Graecis multitudo magna et mulieres nobiles non paucae.
ACTS|17|5|Zelantes autem Iudaei assumentesque de foro viros quosdam malos et turba facta concitaverunt civitatem; et assistentes domui Iasonis quaerebant eos producere in populum.
ACTS|17|6|Et cum non invenissent eos, trahebant Iasonem et quosdam fratres ad politarchas clamantes: " Qui orbem concitaverunt, isti et huc venerunt,
ACTS|17|7|quos suscepit Iason; et hi omnes contra decreta Caesaris faciunt, regem alium dicentes esse, Iesum ".
ACTS|17|8|Concitaverunt autem plebem et politarchas audientes haec;
ACTS|17|9|et accepto satis ab Iasone et a ceteris, dimiserunt eos.
ACTS|17|10|Fratres vero confestim per noctem dimiserunt Paulum et Silam in Beroeam; qui cum advenissent, in synagogam Iudaeorum introierunt.
ACTS|17|11|Hi autem erant nobiliores eorum, qui sunt Thessalonicae, qui susceperunt verbum cum omni aviditate, cotidie scrutantes Scripturas, si haec ita se haberent.
ACTS|17|12|Et multi quidem crediderunt ex eis et Graecarum mulierum honestarum et virorum non pauci.
ACTS|17|13|Cum autem cognovissent in Thessalonica Iudaei quia et Beroeae annuntiatum est a Paulo verbum Dei, venerunt et illuc commoventes et turbantes multitudinem.
ACTS|17|14|Statimque tunc Paulum dimiserunt fratres, ut iret usque ad mare; Silas autem et Timotheus remanserunt ibi.
ACTS|17|15|Qui autem deducebant Paulum, perduxerunt usque Athenas; et accepto mandato ad Silam et Timotheum, ut quam celerrime venirent ad illum, profecti sunt.
ACTS|17|16|Paulus autem cum Athenis eos exspectaret, irritabatur spiritus eius in ipso videns idololatriae deditam civitatem.
ACTS|17|17|Disputabat igitur in synagoga cum Iudaeis et colentibus et in foro per omnes dies ad eos, qui aderant.
ACTS|17|18|Quidam autem ex Epicureis et Stoicis philosophi disserebant cum eo. Et quidam dicebant: " Quid vult seminiverbius hic dicere? "; alii vero: " Novorum daemoniorum videtur annuntiator esse ", quia Iesum et resurrectionem evangelizabat.
ACTS|17|19|Et apprehensum eum ad Areopagum duxerunt dicentes: " Possumus scire quae est haec nova, quae a te dicitur, doctrina?
ACTS|17|20|Mira enim quaedam infers auribus nostris; volumus ergo scire quidnam velint haec esse ".
ACTS|17|21|Athenienses autem omnes et advenae hospites ad nihil aliud vacabant nisi aut dicere aut audire aliquid novi.
ACTS|17|22|Stans autem Paulus in medio Areopagi ait: " Viri Athenienses, per omnia quasi superstitiosiores vos video;
ACTS|17|23|praeteriens enim et videns simulacra vestra inveni et aram, in qua scriptum erat: "Ignoto deo". Quod ergo ignorantes colitis, hoc ego annuntio vobis.
ACTS|17|24|Deus, qui fecit mundum et omnia, quae in eo sunt, hic, caeli et terrae cum sit Dominus, non in manufactis templis inhabitat
ACTS|17|25|nec manibus humanis colitur indigens aliquo, cum ipse det omnibus vitam et inspirationem et omnia;
ACTS|17|26|fecitque ex uno omne genus hominum inhabitare super universam faciem terrae, definiens statuta tempora et terminos habitationis eorum,
ACTS|17|27|quaerere Deum, si forte attrectent eum et inveniant, quamvis non longe sit ab unoquoque nostrum.
ACTS|17|28|In ipso enim vivimus et movemur et sumus, sicut et quidam vestrum poetarum dixerunt:Ipsius enim et genus sumus".
ACTS|17|29|Genus ergo cum simus Dei, non debemus aestimare auro aut argento aut lapidi, sculpturae artis et cogitationis hominis, divinum esse simile.
ACTS|17|30|Et tempora quidem ignorantiae despiciens Deus, nunc annuntiat hominibus, ut omnes ubique paenitentiam agant,
ACTS|17|31|eo quod statuit diem, in qua iudicaturus est orbem in iustitia in viro, quem constituit, fidem praebens omnibus suscitans eum a mortuis ".
ACTS|17|32|Cum audissent autem resurrectionem mortuorum, quidam quidem irridebant, quidam vero dixerunt: " Audiemus te de hoc iterum ".
ACTS|17|33|Sic Paulus exivit de medio eorum.
ACTS|17|34|Quidam vero viri adhaerentes ei crediderunt; in quibus et Dionysius Areopagita et mulier nomine Damaris et alii cum eis.
ACTS|18|1|Post haec discedens ab Athe nis venit Corinthum.
ACTS|18|2|Et in veniens quendam Iudaeum nomine Aquilam, Ponticum genere, qui nuper venerat ab Italia, et Priscillam uxorem eius, eo quod praecepisset Claudius discedere omnes Iudaeos a Roma, accessit ad eos
ACTS|18|3|et, quia eiusdem erat artis, manebat apud eos et operabatur; erant autem scenofactoriae artis.
ACTS|18|4|Disputabat autem in synagoga per omne sabbatum suadebatque Iudaeis et Graecis.
ACTS|18|5|Cum venissent autem de Macedonia Silas et Timotheus, instabat verbo Paulus testificans Iudaeis esse Christum Iesum.
ACTS|18|6|Contradicentibus autem eis et blasphemantibus, excutiens vestimenta dixit ad eos: " Sanguis vester super caput vestrum! Mundus ego. Ex hoc nunc ad gentes vadam ".
ACTS|18|7|Et migrans inde intravit in domum cuiusdam nomine Titi Iusti, colentis Deum, cuius domus erat coniuncta synagogae.
ACTS|18|8|Crispus autem archisynagogus credidit Domino cum omni domo sua, et multi Corinthiorum audientes credebant et baptizabantur.
ACTS|18|9|Dixit autem Dominus nocte per visionem Paulo: " Noli timere, sed loquere et ne taceas,
ACTS|18|10|quia ego sum tecum, et nemo apponetur tibi, ut noceat te, quoniam populus est mihi multus in hac civitate ".
ACTS|18|11|Sedit autem annum et sex menses docens apud eos verbum Dei.
ACTS|18|12|Gallione autem proconsule Achaiae, insurrexerunt uno animo Iudaei in Paulum et adduxerunt eum ad tribunal
ACTS|18|13|dicentes: " Contra legem hic persuadet hominibus colere Deum ".
ACTS|18|14|Incipiente autem Paulo aperire os, dixit Gallio ad Iudaeos: " Si quidem esset iniquum aliquid aut facinus pessimum, o Iudaei, merito vos sustinerem;
ACTS|18|15|si vero quaestiones sunt de verbo et nominibus et lege vestra, vos ipsi videritis; iudex ego horum nolo esse ".
ACTS|18|16|Et minavit eos a tribunali.
ACTS|18|17|Apprehendentes autem omnes Sosthenen, principem synagogae, percutiebant ante tribunal; et nihil horum Gallioni curae erat.
ACTS|18|18|Paulus vero, cum adhuc sustinuisset dies multos, fratribus valefaciens navigabat Syriam, et cum eo Priscilla et Aquila, qui sibi totonderat in Cenchreis caput; habebat enim votum.
ACTS|18|19|Deveneruntque Ephesum, et illos ibi reliquit; ipse vero ingressus synagogam disputabat cum Iudaeis.
ACTS|18|20|Rogantibus autem eis, ut ampliore tempore maneret, non consensit,
ACTS|18|21|sed valefaciens et dicens: " Iterum revertar ad vos Deo volente ", navigavit ab Epheso;
ACTS|18|22|et descendens Caesaream ascendit et salutavit ecclesiam et descendit Antiochiam.
ACTS|18|23|Et facto ibi aliquanto tempore, profectus est perambulans ex ordine Galaticam regionem et Phrygiam, confirmans omnes discipulos.
ACTS|18|24|Iudaeus autem quidam Apollo nomine, Alexandrinus natione, vir eloquens, devenit Ephesum, potens in Scripturis.
ACTS|18|25|Hic erat catechizatus viam Domini; et fervens spiritu loquebatur et docebat diligenter ea, quae sunt de Iesu, sciens tantum baptisma Ioannis.
ACTS|18|26|Hic ergo coepit fiducialiter agere in synagoga; quem cum audissent Priscilla et Aquila, assumpserunt eum et diligentius exposuerunt ei viam Dei.
ACTS|18|27|Cum autem vellet transire in Achaiam, exhortati fratres scripserunt discipulis, ut susciperent eum; qui cum venisset, contulit multum his, qui crediderant per gratiam;
ACTS|18|28|vehementer enim Iudaeos revincebat publice, ostendens per Scripturas esse Christum Iesum.
ACTS|19|1|Factum est autem, cum Apollo esset Corinthi, ut Paulus, peragratis superioribus partibus, veniret Ephesum et inveniret quosdam discipulos;
ACTS|19|2|dixitque ad eos: " Si Spiritum Sanctum accepistis credentes? ". At illi ad eum: " Sed neque, si Spiritus Sanctus est, audivimus ".
ACTS|19|3|Ille vero ait: " In quo ergo baptizati estis? ". Qui dixerunt: " In Ioannis baptismate ".
ACTS|19|4|Dixit autem Paulus: " Ioannes baptizavit baptisma paenitentiae, populo dicens in eum, qui venturus esset post ipsum ut crederent, hoc est in Iesum ".
ACTS|19|5|His auditis, baptizati sunt in nomine Domini Iesu;
ACTS|19|6|et cum imposuisset illis manus Paulus, venit Spiritus Sanctus super eos, et loquebantur linguis et prophetabant.
ACTS|19|7|Erant autem omnes viri fere duodecim.
ACTS|19|8|Introgressus autem synagogam cum fiducia loquebatur per tres menses disputans et suadens de regno Dei.
ACTS|19|9|Cum autem quidam indurarentur et non crederent maledicentes viam coram multitudine, discedens ab eis segregavit discipulos, cotidie disputans in schola Tyranni.
ACTS|19|10|Hoc autem factum est per biennium, ita ut omnes, qui habitabant in Asia, audirent verbum Domini, Iudaei atque Graeci.
ACTS|19|11|Virtutesque non quaslibet Deus faciebat per manus Pauli,
ACTS|19|12|ita ut etiam super languidos deferrentur a corpore eius sudaria vel semicinctia, et recederent ab eis languores, et spiritus nequam egrederentur.
ACTS|19|13|Tentaverunt autem quidam et de circumeuntibus Iudaeis exorcistis invocare super eos, qui habebant spiritus malos, nomen Domini Iesu dicentes: " Adiuro vos per Iesum, quem Paulus praedicat ".
ACTS|19|14|Erant autem cuiusdam Scevae Iudaei principis sacerdotum septem filii, qui hoc faciebant.
ACTS|19|15|Respondens autem spiritus nequam dixit eis: " Iesum novi et Paulum scio; vos autem qui estis? ".
ACTS|19|16|Et insiliens homo in eos, in quo erat spiritus malus, dominatus amborum invaluit contra eos, ita ut nudi et vulnerati effugerent de domo illa.
ACTS|19|17|Hoc autem notum factum est omnibus Iudaeis atque Graecis, qui habitabant Ephesi, et cecidit timor super omnes illos, et magnificabatur nomen Domini Iesu.
ACTS|19|18|Multique credentium veniebant confitentes et annuntiantes actus suos.
ACTS|19|19|Multi autem ex his, qui fuerant curiosa sectati, conferentes libros combusserunt coram omnibus; et computaverunt pretia illorum et invenerunt argenti quinquaginta milia.
ACTS|19|20|Ita fortiter verbum Domini crescebat et convalescebat.
ACTS|19|21|His autem expletis, proposuit Paulus in Spiritu, transita Macedonia et Achaia, ire Hierosolymam, dicens: " Postquam fuero ibi, oportet me et Romam videre ".
ACTS|19|22|Mittens autem in Macedoniam duos ex ministrantibus sibi, Timotheum et Erastum, ipse remansit ad tempus in Asia.
ACTS|19|23|Facta est autem in illo tempore turbatio non minima de via.
ACTS|19|24|Demetrius enim quidam nomine, argentarius, faciens aedes argenteas Dianae praestabat artificibus non modicum quaestum;
ACTS|19|25|quos congregans et eos, qui eiusmodi erant opifices, dixit: " Viri, scitis quia de hoc artificio acquisitio est nobis;
ACTS|19|26|et videtis et auditis quia non solum Ephesi, sed paene totius Asiae Paulus hic suadens avertit multam turbam dicens quoniam non sunt dii, qui manibus fiunt.
ACTS|19|27|Non solum autem haec periclitatur nobis pars in redargutionem venire, sed et magnae deae Dianae templum in nihilum reputari, et destrui incipiet maiestas eius, quam tota Asia et orbis colit ".
ACTS|19|28|His auditis, repleti sunt ira et clamabant dicentes: " Magna Diana Ephesiorum! ";
ACTS|19|29|et impleta est civitas confusione, et impetum fecerunt uno animo in theatrum, rapto Gaio et Aristarcho Macedonibus, comitibus Pauli.
ACTS|19|30|Paulo autem volente intrare in populum, non permiserunt discipuli;
ACTS|19|31|quidam autem de Asiarchis, qui erant amici eius, miserunt ad eum rogantes, ne se daret in theatrum.
ACTS|19|32|Alii autem aliud clamabant; erat enim ecclesia confusa, et plures nesciebant qua ex causa convenissent.
ACTS|19|33|De turba autem instruxerunt Alexandrum, propellentibus eum Iudaeis; Alexander ergo, manu silentio postulato, volebat rationem reddere populo.
ACTS|19|34|Quem ut cognoverunt Iudaeum esse, vox facta est una omnium quasi per horas duas clamantium: " Magna Diana Ephesiorum ".
ACTS|19|35|Et cum sedasset scriba turbam, dixit: " Viri Ephesii, quis enim est hominum, qui nesciat Ephesiorum civitatem cultricem esse magnae Dianae et simulacri a Iove delapsi?
ACTS|19|36|Cum ergo his contradici non possit, oportet vos sedatos esse et nihil temere agere.
ACTS|19|37|Adduxistis enim homines istos neque sacrilegos neque blasphemantes deam nostram.
ACTS|19|38|Quod si Demetrius et, qui cum eo sunt, artifices habent adversus aliquem causam, conventus forenses aguntur, et proconsules sunt: accusent invicem.
ACTS|19|39|Si quid autem ulterius quaeritis, in legitima ecclesia poterit absolvi.
ACTS|19|40|Nam et periclitamur argui seditionis hodiernae, cum nullus obnoxius sit, de quo non possimus reddere rationem concursus istius ". Et cum haec dixisset, dimisit ecclesiam.
ACTS|20|1|Postquam autem cessavit tumultus, accersitis Paulus discipulis et exhortatus eos, valedixit et profectus est, ut iret in Macedoniam.
ACTS|20|2|Cum autem perambulasset partes illas et exhortatus eos fuisset multo sermone, venit ad Graeciam;
ACTS|20|3|cumque fecisset menses tres, factae sunt illi insidiae a Iudaeis navigaturo in Syriam, habuitque consilium, ut reverteretur per Macedoniam.
ACTS|20|4|Comitabatur autem eum Sopater Pyrrhi Beroeensis, Thessalonicensium vero Aristarchus et Secundus et Gaius Derbeus et Timotheus, Asiani vero Tychicus et Trophimus.
ACTS|20|5|Hi cum praecessissent, sustinebant nos Troade;
ACTS|20|6|nos vero navigavimus post dies Azymorum a Philippis et venimus ad eos Troadem in diebus quinque, ubi demorati sumus diebus septem.
ACTS|20|7|In una autem sabbatorum, cum convenissemus ad frangendum panem, Paulus disputabat eis, profecturus in crastinum, protraxitque sermonem usque in mediam noctem.
ACTS|20|8|Erant autem lampades copiosae in cenaculo, ubi eramus congregati;
ACTS|20|9|sedens autem quidam adulescens nomine Eutychus super fenestram, cum mergeretur somno gravi, disputante diutius Paulo, eductus somno cecidit de tertio cenaculo deorsum et sublatus est mortuus.
ACTS|20|10|Cum descendisset autem Paulus, incubuit super eum et complexus dixit: " Nolite turbari, anima enim ipsius in eo est! ".
ACTS|20|11|Ascendens autem frangensque panem et gustans satisque allocutus usque in lucem, sic profectus est.
ACTS|20|12|Adduxerunt autem puerum viventem et consolati sunt non minime.
ACTS|20|13|Nos autem praecedentes navi enavigavimus in Asson, inde suscepturi Paulum; sic enim disposuerat volens ipse per terram iter facere.
ACTS|20|14|Cum autem convenisset nos in Asson, assumpto eo, venimus Mitylenen
ACTS|20|15|et inde navigantes sequenti die pervenimus contra Chium et alia applicuimus Samum et sequenti venimus Miletum.
ACTS|20|16|Proposuerat enim Paulus transnavigare Ephesum, ne qua mora illi fieret in Asia; festinabat enim, si possibile sibi esset, ut diem Pentecosten faceret Hierosolymis.
ACTS|20|17|A Mileto autem mittens Ephesum convocavit presbyteros ecclesiae.
ACTS|20|18|Qui cum venissent ad eum, dixit eis: " Vos scitis a prima die, qua ingressus sum in Asiam, qualiter vobiscum per omne tempus fuerim,
ACTS|20|19|serviens Domino cum omni humilitate et lacrimis et tentationibus, quae mihi acciderunt in insidiis Iudaeorum;
ACTS|20|20|quomodo nihil subtraxerim utilium, quominus annuntiarem vobis et docerem vos publice et per domos,
ACTS|20|21|testificans Iudaeis atque Graecis in Deum paenitentiam et fidem in Dominum nostrum Iesum.
ACTS|20|22|Et nunc ecce alligatus ego Spiritu vado in Ierusalem, quae in ea eventura sint mihi ignorans,
ACTS|20|23|nisi quod Spiritus Sanctus per omnes civitates protestatur mihi dicens quoniam vincula et tribulationes me manent.
ACTS|20|24|Sed nihili facio animam meam pretiosam mihi, dummodo consummem cursum meum et ministerium, quod accepi a Domino Iesu, testificari evangelium gratiae Dei.
ACTS|20|25|Et nunc ecce ego scio quia amplius non videbitis faciem meam vos omnes, per quos transivi praedicans regnum;
ACTS|20|26|quapropter contestor vos hodierna die, quia mundus sum a sanguine omnium;
ACTS|20|27|non enim subterfugi, quominus annuntiarem omne consilium Dei vobis.
ACTS|20|28|Attendite vobis et universo gregi, in quo vos Spiritus Sanctus posuit episcopos, pascere ecclesiam Dei, quam acquisivit sanguine suo.
ACTS|20|29|Ego scio quoniam intrabunt post discessionem meam lupi graves in vos non parcentes gregi;
ACTS|20|30|et ex vobis ipsis exsurgent viri loquentes perversa, ut abstrahant discipulos post se.
ACTS|20|31|Propter quod vigilate, memoria retinentes quoniam per triennium nocte et die non cessavi cum lacrimis monens unumquemque vestrum.
ACTS|20|32|Et nunc commendo vos Deo et verbo gratiae ipsius, qui potens est aedificare et dare hereditatem in sanctificatis omnibus.
ACTS|20|33|Argentum aut aurum aut vestem nullius concupivi;
ACTS|20|34|ipsi scitis quoniam ad ea, quae mihi opus erant et his, qui mecum sunt, ministraverunt manus istae.
ACTS|20|35|Omnia ostendi vobis quoniam sic laborantes oportet suscipere infirmos, ac meminisse verborum Domini Iesu, quoniam ipse dixit: "Beatius est magis dare quam accipere!" ".
ACTS|20|36|Et cum haec dixisset, positis genibus suis, cum omnibus illis oravit.
ACTS|20|37|Magnus autem fletus factus est omnium; et procumbentes super collum Pauli osculabantur eum
ACTS|20|38|dolentes maxime in verbo, quod dixerat, quoniam amplius faciem eius non essent visuri. Et deducebant eum ad navem.
ACTS|21|1|Cum autem factum esset, ut navigaremus abstracti ab eis, recto cursu venimus Cho et sequenti die Rhodum et inde Patara;
ACTS|21|2|et cum invenissemus navem transfretantem in Phoenicen, ascendentes navigavimus.
ACTS|21|3|Cum paruissemus autem Cypro, et relinquentes eam ad sinistram navigabamus in Syriam et venimus Tyrum, ibi enim navis erat expositura onus.
ACTS|21|4|Inventis autem discipulis, mansimus ibi diebus septem; qui Paulo dicebant per Spiritum, ne iret Hierosolymam.
ACTS|21|5|Et explicitis diebus, profecti ibamus, deducentibus nos omnibus cum uxoribus et filiis usque foras civitatem; et positis genibus in litore orantes,
ACTS|21|6|valefecimus invicem et ascendimus in navem; illi autem redierunt in sua.
ACTS|21|7|Nos vero, navigatione explicita, a Tyro devenimus Ptolemaida et, salutatis fratribus, mansimus die una apud illos.
ACTS|21|8|Alia autem die profecti venimus Caesaream et intrantes in domum Philippi evangelistae, qui erat de septem, mansimus apud eum.
ACTS|21|9|Huic autem erant filiae quattuor virgines prophetantes.
ACTS|21|10|Et cum moraremur plures dies, supervenit quidam a Iudaea propheta nomine Agabus;
ACTS|21|11|is cum venisset ad nos et tulisset zonam Pauli, alligans sibi pedes et manus dixit: " Haec dicit Spiritus Sanctus: Virum, cuius est zona haec, sic alligabunt in Ierusalem Iudaei et tradent in manus gentium ".
ACTS|21|12|Quod cum audissemus, rogabamus nos et, qui loci illius erant, ne ipse ascenderet Ierusalem.
ACTS|21|13|Tunc respondit Paulus: " Quid facitis flentes et affligentes cor meum? Ego enim non solum alligari sed et mori in Ierusalem paratus sum propter nomen Domini Iesu ".
ACTS|21|14|Et cum ei suadere non possemus, quievimus dicentes: " Domini voluntas fiat! ".
ACTS|21|15|Post dies autem istos praeparati ascendebamus Hierosolymam;
ACTS|21|16|venerunt autem et ex discipulis a Caesarea nobiscum adducentes apud quem hospitaremur, Mnasonem quendam Cyprium, antiquum discipulum.
ACTS|21|17|Et cum venissemus Hierosolymam, libenter exceperunt nos fratres.
ACTS|21|18|Sequenti autem die introibat Paulus nobiscum ad Iacobum, omnesque collecti sunt presbyteri.
ACTS|21|19|Quos cum salutasset, narrabat per singula, quae fecisset Deus in gentibus per ministerium ipsius.
ACTS|21|20|At illi cum audissent, glorificabant Deum dixeruntque ei: " Vides, frater, quot milia sint in Iudaeis, qui crediderunt, et omnes aemulatores sunt legis;
ACTS|21|21|audierunt autem de te quia discessionem doceas a Moyse omnes, qui per gentes sunt, Iudaeos, dicens non debere circumcidere eos filios suos neque secundum consuetudines ambulare.
ACTS|21|22|Quid ergo est? Utique audient te supervenisse.
ACTS|21|23|Hoc ergo fac, quod tibi dicimus. Sunt nobis viri quattuor votum habentes super se;
ACTS|21|24|his assumptis, sanctifica te cum illis et impende pro illis, ut radant capita, et scient omnes quia, quae de te audierunt, nihil sunt, sed ambulas et ipse custodiens legem.
ACTS|21|25|De his autem, qui crediderunt, gentibus nos scripsimus iudicantes, ut abstineant ab idolothyto et sanguine et suffocato et fornicatione ".
ACTS|21|26|Tunc Paulus, assumptis viris, postera die purificatus cum illis intravit in templum annuntians expletionem dierum purificationis, donec offerretur pro unoquoque eorum oblatio.
ACTS|21|27|Dum autem septem dies consummarentur, hi, qui de Asia erant, Iudaei cum vidissent eum in templo, concitaverunt omnem turbam et iniecerunt ei manus
ACTS|21|28|clamantes: " Viri Israelitae, adiuvate! Hic est homo, qui adversus populum et legem et locum hunc omnes ubique docens, insuper et Graecos induxit in templum et polluit sanctum locum istum ".
ACTS|21|29|Viderant enim Trophimum Ephesium in civitate cum ipso, quem aestimabant quoniam in templum induxisset Paulus.
ACTS|21|30|Commotaque est civitas tota, et facta est concursio populi, et apprehendentes Paulum trahebant eum extra templum, et statim clausae sunt ianuae.
ACTS|21|31|Quaerentibus autem eum occidere, nuntiatum est tribuno cohortis quia tota confunditur Ierusalem,
ACTS|21|32|qui statim, assumptis militibus et centurionibus, decucurrit ad illos; qui cum vidissent tribunum et milites, cessaverunt percutere Paulum.
ACTS|21|33|Tunc accedens tribunus apprehendit eum et iussit alligari catenis duabus et interrogabat quis esset et quid fecisset.
ACTS|21|34|Alii autem aliud clamabant in turba; et cum non posset certum cognoscere prae tumultu, iussit duci eum in castra.
ACTS|21|35|Et cum venisset ad gradus, contigit ut portaretur a militibus propter vim turbae;
ACTS|21|36|sequebatur enim multitudo populi clamantes: " Tolle eum! ".
ACTS|21|37|Et cum coepisset induci in castra, Paulus dicit tribuno: " Si licet mihi loqui aliquid ad te? ". Qui dixit: " Graece nosti?
ACTS|21|38|Nonne tu es Aegyptius, qui ante hos dies tumultum concitasti et eduxisti in desertum quattuor milia virorum sicariorum? ".
ACTS|21|39|Et dixit Paulus: " Ego homo sum quidem Iudaeus a Tarso Ciliciae, non ignotae civitatis municeps; rogo autem te, permitte mihi loqui ad populum.
ACTS|21|40|Et cum ille permisisset, Paulus stans in gradibus annuit manu ad plebem et, magno silentio facto, allocutus est Hebraea lingua dicens:
ACTS|22|1|" Viri fratres et patres, audi te a me, quam ad vos nunc reddo, rationem.
ACTS|22|2|Cum audissent autem quia Hebraea lingua loquebatur ad illos, magis praestiterunt silentium. Et dixit:
ACTS|22|3|" Ego sum vir Iudaeus, natus Tarso Ciliciae, enutritus autem in ista civitate, secus pedes Gamaliel eruditus iuxta veritatem paternae legis, aemulator Dei, sicut et vos omnes estis hodie.
ACTS|22|4|Qui hanc viam persecutus sum usque ad mortem, alligans et tradens in custodias viros ac mulieres,
ACTS|22|5|sicut et princeps sacerdotum testimonium mihi reddit et omne concilium; a quibus et epistulas accipiens ad fratres, Damascum pergebam, ut adducerem et eos, qui ibi essent, vinctos in Ierusalem, uti punirentur.
ACTS|22|6|Factum est autem, eunte me et appropinquante Damasco, circa mediam diem subito de caelo circumfulsit me lux copiosa;
ACTS|22|7|et decidi in terram et audivi vocem dicentem mihi: "Saul, Saul, quid me persequeris?".
ACTS|22|8|Ego autem respondi: "Quis es, Domine?". Dixitque ad me: "Ego sum Iesus Nazarenus, quem tu persequeris".
ACTS|22|9|Et, qui mecum erant, lumen quidem viderunt, vocem autem non audierunt eius, qui loquebatur mecum.
ACTS|22|10|Et dixi: "Quid faciam, Domine?". Dominus autem dixit ad me: "Surgens vade Damascum, et ibi tibi dicetur de omnibus, quae statutum est tibi, ut faceres".
ACTS|22|11|Et cum non viderem prae claritate luminis illius, ad manum deductus a comitibus veni Damascum.
ACTS|22|12|Ananias autem quidam vir religiosus secundum legem, testimonium habens ab omnibus habitantibus Iudaeis,
ACTS|22|13|veniens ad me et astans dixit mihi: "Saul frater, respice!". Et ego eadem hora respexi in eum.
ACTS|22|14|At ille dixit: "Deus patrum nostrorum praeordinavit te, ut cognosceres voluntatem eius et videres Iustum et audires vocem ex ore eius,
ACTS|22|15|quia eris testis illi ad omnes homines eorum, quae vidisti et audisti.
ACTS|22|16|Et nunc quid moraris? Exsurgens baptizare et ablue peccata tua, invocato nomine ipsius".
ACTS|22|17|Factum est autem, revertenti mihi in Ierusalem et oranti in templo fieri me in stupore mentis
ACTS|22|18|et videre illum dicentem mihi: "Festina et exi velociter ex Ierusalem, quoniam non recipient testimonium tuum de me".
ACTS|22|19|Et ego dixi: "Domine, ipsi sciunt quia ego eram concludens in carcerem et caedens per synagogas eos, qui credebant in te;
ACTS|22|20|et cum funderetur sanguis Stephani testis tui, et ipse astabam et consentiebam et custodiebam vestimenta interficientium illum".
ACTS|22|21|Et dixit ad me: "Vade, quoniam ego in nationes longe mittam te" ".
ACTS|22|22|Audiebant autem eum usque ad hoc verbum et levaverunt vocem suam dicentes: " Tolle de terra eiusmodi, non enim fas est eum vivere! ".
ACTS|22|23|Vociferantibus autem eis et proicientibus vestimenta sua et pulverem iactantibus in aerem,
ACTS|22|24|iussit tribunus induci eum in castra dicens flagellis eum interrogari, ut sciret propter quam causam sic acclamarent ei.
ACTS|22|25|Et cum astrinxissent eum loris, dixit astanti centurioni Paulus: " Si hominem Romanum et indemnatum licet vobis flagellare? ".
ACTS|22|26|Quo audito, centurio accedens ad tribunum nuntiavit dicens: " Quid acturus es? Hic enim homo Romanus est ".
ACTS|22|27|Accedens autem tribunus dixit illi: " Dic mihi, tu Romanus es? ". At ille dixit: " Etiam ".
ACTS|22|28|Et respondit tribunus: " Ego multa summa civitatem hanc consecutus sum. Et Paulus ait: " Ego autem et natus sum ".
ACTS|22|29|Protinus ergo discesserunt ab illo, qui eum interrogaturi erant; tribunus quoque timuit, postquam rescivit quia Romanus esset, et quia alligasset eum.
ACTS|22|30|Postera autem die, volens scire diligenter qua ex causa accusaretur a Iudaeis, solvit eum et iussit principes sacerdotum convenire et omne concilium et producens Paulum statuit coram illis.
ACTS|23|1|Intendens autem concilium Paulus ait: " Viri fratres, ego omni conscientia bona conversatus sum ante Deum usque in hodiernum diem ".
ACTS|23|2|Princeps autem sacerdotum Ananias praecepit astantibus sibi percutere os eius.
ACTS|23|3|Tunc Paulus ad eum dixit: " Percutiet te Deus, paries dealbate! Et tu sedes iudicans me secundum legem et contra legem iubes me percuti? ".
ACTS|23|4|Et, qui astabant, dixerunt: " Summum sacerdotem Dei maledicis?".
ACTS|23|5|Dixit autem Paulus: " Nesciebam, fratres, quia princeps est sacerdotum; scriptum est enim: "Principem populi tui non maledices" ".
ACTS|23|6|Sciens autem Paulus quia una pars esset sadducaeorum, et altera pharisaeorum, exclamabat in concilio: " Viri fratres, ego pharisaeus sum, filius pharisaeorum; de spe et resurrectione mortuorum ego iudicor ".
ACTS|23|7|Et cum haec diceret, facta est dissensio inter pharisaeos et sadducaeos; et divisa est multitudo.
ACTS|23|8|Sadducaei enim dicunt non esse resurrectionem neque angelum neque spiritum; pharisaei autem utrumque confitentur.
ACTS|23|9|Factus est autem clamor magnus; et surgentes scribae quidam partis pharisaeorum pugnabant dicentes: " Nihil mali invenimus in homine isto: quod si spiritus locutus est ei aut angelus ";
ACTS|23|10|et cum magna dissensio facta esset, timens tribunus ne discerperetur Paulus ab ipsis, iussit milites descendere, ut raperent eum de medio eorum ac deducerent in castra.
ACTS|23|11|Sequenti autem nocte, assistens ei Dominus ait: " Constans esto! Sicut enim testificatus es, quae sunt de me, in Ierusalem, sic te oportet et Romae testificari ".
ACTS|23|12|Facta autem die, faciebant concursum Iudaei et devoverunt se dicentes neque manducaturos neque bibituros, donec occiderent Paulum.
ACTS|23|13|Erant autem plus quam quadraginta, qui hanc coniurationem fecerant;
ACTS|23|14|qui accedentes ad principes sacerdotum et seniores dixerunt: " Devotione devovimus nos nihil gustaturos, donec occidamus Paulum.
ACTS|23|15|Nunc ergo vos notum facite tribuno cum concilio, ut producat illum ad vos, tamquam aliquid certius cognituri de eo; nos vero, priusquam appropiet, parati sumus interficere illum ".
ACTS|23|16|Quod cum audisset filius sororis Pauli insidias, venit et intravit in castra nuntiavitque Paulo.
ACTS|23|17|Vocans autem Paulus ad se unum ex centurionibus ait: " Adulescentem hunc perduc ad tribunum, habet enim aliquid indicare illi ".
ACTS|23|18|Et ille quidem assumens eum duxit ad tribunum et ait: " Vinctus Paulus vocans rogavit me hunc adulescentem perducere ad te, habentem aliquid loqui tibi ".
ACTS|23|19|Apprehendens autem tribunus manum illius, secessit cum eo seorsum et interrogabat: " Quid est, quod habes indicare mihi? ".
ACTS|23|20|Ille autem dixit: " Iudaei constituerunt rogare te, ut crastina die Paulum producas in concilium, quasi aliquid certius inquisiturum sit de illo.
ACTS|23|21|Tu ergo ne credideris illis; insidiantur enim ei ex eis viri amplius quadraginta, qui se devoverunt non manducare neque bibere, donec interficiant eum; et nunc parati sunt exspectantes promissum tuum ".
ACTS|23|22|Tribunus igitur dimisit adulescentem praecipiens, ne cui eloqueretur quoniam " haec nota mihi fecisti ".
ACTS|23|23|Et vocatis duobus centurionibus, dixit: " Parate milites ducentos, ut eant usque Caesaream, et equites septuaginta et lancearios ducentos, a tertia hora noctis,
ACTS|23|24|et iumenta praeparate ", ut imponentes Paulum salvum perducerent ad Felicem praesidem,
ACTS|23|25|scribens epistulam habentem formam hanc:
ACTS|23|26|" Claudius Lysias optimo praesidi Felici salutem.
ACTS|23|27|Virum hunc comprehensum a Iudaeis et incipientem interfici ab eis, superveniens cum exercitu eripui, cognito quia Romanus est.
ACTS|23|28|Volensque scire causam, propter quam accusabant illum, deduxi in concilium eorum;
ACTS|23|29|quem inveni accusari de quaestionibus legis ipsorum, nihil vero dignum morte aut vinculis habentem crimen.
ACTS|23|30|Et cum mihi perlatum esset de insidiis, quae in virum pararentur, confestim misi ad te denuntians et accusatoribus, ut dicant adversum eum apud te ".
ACTS|23|31|Milites ergo, secundum praeceptum sibi assumentes Paulum, duxerunt per noctem in Antipatridem;
ACTS|23|32|et postera die, dimissis equitibus, ut abirent cum eo, reversi sunt ad castra.
ACTS|23|33|Qui cum venissent Caesaream et tradidissent epistulam praesidi, statuerunt ante illum et Paulum.
ACTS|23|34|Cum legisset autem et interrogasset de qua provincia esset, et cognoscens quia de Cilicia:
ACTS|23|35|" Audiam te, inquit, cum et accusatores tui venerint "; iussitque in praetorio Herodis custodiri eum.
ACTS|24|1|Post quinque autem dies, descendit princeps sacerdo tum Ananias cum senioribus quibusdam et Tertullo quodam oratore, qui adierunt praesidem adversus Paulum.
ACTS|24|2|Et citato eo, coepit accusare Tertullus dicens: " Cum in multa pace agamus per te, et multa corrigantur genti huic per tuam providentiam,
ACTS|24|3|semper et ubique suscipimus, optime Felix, cum omni gratiarum actione.
ACTS|24|4|Ne diutius autem te protraham, oro, breviter audias nos pro tua clementia.
ACTS|24|5|Invenimus enim hunc hominem pestiferum et concitantem seditiones omnibus Iudaeis, qui sunt in universo orbe, et auctorem seditionis sectae Nazarenorum,
ACTS|24|6|qui etiam templum violare conatus est, quem et apprehendimus,
ACTS|24|7|()
ACTS|24|8|a quo poteris ipse diiudicans de omnibus istis cognoscere, de quibus nos accusamus eum ".
ACTS|24|9|Adiecerunt autem et Iudaei dicentes haec ita se habere.
ACTS|24|10|Respondit autem Paulus, annuente sibi praeside dicere: " Ex multis annis esse te iudicem genti huic sciens bono animo de causa mea rationem reddam,
ACTS|24|11|cum possis cognoscere quia non plus sunt dies mihi quam duodecim, ex quo ascendi adorare in Ierusalem,
ACTS|24|12|et neque in templo invenerunt me cum aliquo disputantem aut concursum facientem turbae neque in synagogis neque in civitate,
ACTS|24|13|neque probare possunt tibi, de quibus nunc accusant me.
ACTS|24|14|Confiteor autem hoc tibi, quod secundum viam, quam dicunt haeresim, sic deservio patrio Deo credens omnibus, quae secundum Legem sunt et in Prophetis scripta,
ACTS|24|15|spem habens in Deum, quam et hi ipsi exspectant, resurrectionem futuram iustorum et iniquorum.
ACTS|24|16|In hoc et ipse studeo sine offendiculo conscientiam habere ad Deum et ad homines semper.
ACTS|24|17|Post annos autem plures, eleemosynas facturus in gentem meam veni et oblationes;
ACTS|24|18|in quibus invenerunt me purificatum in templo, non cum turba neque cum tumultu;
ACTS|24|19|quidam autem ex Asia Iudaei, quos oportebat apud te praesto esse et accusare, si quid haberent adversum me;
ACTS|24|20|aut hi ipsi dicant quid invenerint iniquitatis, cum starem in concilio,
ACTS|24|21|nisi de una hac voce, qua clamavi inter eos stans: De resurrectione mortuorum ego iudicor hodie apud vos! ".
ACTS|24|22|Distulit autem illos Felix certissime sciens ea, quae de hac via sunt, dicens: " Cum tribunus Lysias descenderit, cognoscam causam vestram ",
ACTS|24|23|iubens centurioni custodiri eum et habere mitigationem, nec quemquam prohibere de suis ministrare ei.
ACTS|24|24|Post aliquot autem dies, adveniens Felix cum Drusilla uxore sua, quae erat Iudaea, vocavit Paulum et audivit ab eo de fide, quae est in Christum Iesum.
ACTS|24|25|Disputante autem illo de iustitia et continentia et de iudicio futuro, timefactus Felix respondit: " Quod nunc attinet, vade; tempore autem opportuno accersiam te ",
ACTS|24|26|simul et sperans quia pecunia daretur sibi a Paulo; propter quod et frequenter accersiens eum loquebatur cum eo.
ACTS|24|27|Biennio autem expleto, accepit successorem Felix Porcium Festum; volensque gratiam praestare Iudaeis, Felix reliquit Paulum vinctum.
ACTS|25|1|Festus ergo cum venisset in provinciam, post triduum ascendit Hierosolymam a Caesarea;
ACTS|25|2|adieruntque eum principes sacerdotum et primi Iudaeorum adversus Paulum, et rogabant eum
ACTS|25|3|postulantes gratiam adversum eum, ut iuberet perduci eum in Ierusalem, insidias tendentes, ut eum interficerent in via.
ACTS|25|4|Festus igitur respondit servari Paulum in Caesarea, se autem maturius profecturum:
ACTS|25|5|" Qui ergo in vobis, ait, potentes sunt, descendentes simul, si quod est in viro crimen, accusent eum ".
ACTS|25|6|Demoratus autem inter eos dies non amplius quam octo aut decem, descendit Caesaream; et altera die sedit pro tribunali et iussit Paulum adduci.
ACTS|25|7|Qui cum perductus esset, circumsteterunt eum, qui ab Hierosolyma descenderant, Iudaei, multas et graves causas obicientes, quas non poterant probare,
ACTS|25|8|Paulo rationem reddente: " Neque in legem Iudaeorum neque in templum neque in Caesarem quidquam peccavi ".
ACTS|25|9|Festus autem volens Iudaeis gratiam praestare, respondens Paulo dixit: " Vis Hierosolymam ascendere et ibi de his iudicari apud me? ".
ACTS|25|10|Dixit autem Paulus: " Ad tribunal Caesaris sto, ubi me oportet iudicari. Iudaeis nihil nocui, sicut et tu melius nosti.
ACTS|25|11|Si ergo iniuste egi et dignum morte aliquid feci, non recuso mori; si vero nihil est eorum, quae hi accusant me, nemo potest me illis donare. Caesarem appello! ".
ACTS|25|12|Tunc Festus cum consilio locutus respondit: " Caesarem appellasti; ad Caesarem ibis ".
ACTS|25|13|Et cum dies aliquot transacti essent, Agrippa rex et Berenice descenderunt Caesaream et salutaverunt Festum.
ACTS|25|14|Et cum dies plures ibi demorarentur, Festus regi indicavit de Paulo dicens: " Vir quidam est derelictus a Felice vinctus,
ACTS|25|15|de quo, cum essem Hierosolymis, adierunt me principes sacerdotum et seniores Iudaeorum postulantes adversus illum damnationem;
ACTS|25|16|ad quos respondi, quia non est consuetudo Romanis donare aliquem hominem, priusquam is, qui accusatur, praesentes habeat accusatores locumque defendendi se ab accusatione accipiat.
ACTS|25|17|Cum ergo huc convenissent, sine ulla dilatione sequenti die sedens pro tribunali iussi adduci virum;
ACTS|25|18|de quo, cum stetissent accusatores, nullam causam deferebant, de quibus ego suspicabar malis;
ACTS|25|19|quaestiones vero quasdam de sua superstitione habebant adversus eum et de quodam Iesu defuncto, quem affirmabat Paulus vivere.
ACTS|25|20|Haesitans autem ego de huiusmodi quaestione, dicebam si vellet ire Hierosolymam et ibi iudicari de istis.
ACTS|25|21|Paulo autem appellante, ut servaretur ad Augusti cognitionem, iussi servari eum, donec mittam eum ad Caesarem ".
ACTS|25|22|Agrippa autem ad Festum: " Volebam et ipse hominem audire! ". " Cras, inquit, audies eum ".
ACTS|25|23|Altera autem die, cum venisset Agrippa et Berenice cum multa ambitione, et introissent in auditorium cum tribunis et viris principalibus civitatis, et iubente Festo, adductus est Paulus.
ACTS|25|24|Et dicit Festus: " Agrippa rex et omnes, qui simul adestis nobiscum viri, videtis hunc, de quo omnis multitudo Iudaeorum interpellavit me Hierosolymis et hic, clamantes non oportere eum vivere amplius.
ACTS|25|25|Ego vero comperi nihil dignum eum morte fecisse, ipso autem hoc appellante Augustum, iudicavi mittere.
ACTS|25|26|De quo quid certum scribam domino, non habeo; propter quod produxi eum ad vos et maxime ad te, rex Agrippa, ut, interrogatione facta, habeam quid scribam;
ACTS|25|27|sine ratione enim mihi videtur mittere vinctum et causas eius non significare ".
ACTS|26|1|Agrippa vero ad Paulum ait: " Permittitur tibi loqui pro temetipso ". Tunc Paulus, extenta manu, coepit rationem reddere:
ACTS|26|2|" De omnibus, quibus accusor a Iudaeis, rex Agrippa, aestimo me beatum, apud te cum sim defensurus me hodie,
ACTS|26|3|maxime te sciente omnia, quae apud Iudaeos sunt consuetudines et quaestiones; propter quod, obsecro, patienter me audias.
ACTS|26|4|Et quidem vitam meam a iuventute, quae ab initio fuit in gente mea et in Hierosolymis, noverunt omnes Iudaei;
ACTS|26|5|praescientes me ab initio, si velint testimonium perhibere, quoniam secundum diligentissimam sectam nostrae religionis vixi pharisaeus.
ACTS|26|6|Et nunc propter spem eius, quae ad patres nostros repromissionis facta est a Deo, sto iudicio subiectus,
ACTS|26|7|in quam duodecim tribus nostrae cum perseverantia nocte ac die deservientes sperant devenire; de qua spe accusor a Iudaeis, rex!
ACTS|26|8|Quid incredibile iudicatur apud vos, si Deus mortuos suscitat?
ACTS|26|9|Et ego quidem existimaveram me adversus nomen Iesu Nazareni debere multa contraria agere;
ACTS|26|10|quod et feci Hierosolymis, et multos sanctorum ego in carceribus inclusi, a principibus sacerdotum potestate accepta, et cum occiderentur, detuli sententiam;
ACTS|26|11|et per omnes synagogas frequenter puniens eos compellebam blasphemare, et abundantius insaniens in eos persequebar usque in exteras civitates.
ACTS|26|12|In quibus, dum irem Damascum cum potestate et permissu principum sacerdotum,
ACTS|26|13|die media in via vidi, rex, de caelo supra splendorem solis circumfulgens me lumen et eos, qui mecum simul ibant;
ACTS|26|14|omnesque nos cum decidissemus in terram, audivi vocem loquentem mihi Hebraica lingua: "Saul, Saul, quid me persequeris? Durum est tibi contra stimulum calcitrare".
ACTS|26|15|Ego autem dixi: "Quis es, Domine?". Dominus autem dixit: "Ego sum Iesus, quem tu persequeris.
ACTS|26|16|Sed exsurge et sta super pedes tuos; ad hoc enim apparui tibi, ut constituam te ministrum et testem eorum, quae vidisti, et eorum, quibus apparebo tibi,
ACTS|26|17|eripiens te de populo et de gentibus, in quas ego mitto te
ACTS|26|18|aperire oculos eorum, ut convertantur a tenebris ad lucem et de potestate Satanae ad Deum, ut accipiant remissionem peccatorum et sortem inter sanctificatos per fidem, quae est in me".
ACTS|26|19|Unde, rex Agrippa, non fui incredulus caelestis visionis,
ACTS|26|20|sed his, qui sunt Damasci primum et Hierosolymis, et in omnem regionem Iudaeae et gentibus annuntiabam, ut paenitentiam agerent et converterentur ad Deum digna paenitentiae opera facientes.
ACTS|26|21|Hac ex causa me Iudaei, cum essem in templo comprehensum, tentabant interficere.
ACTS|26|22|Auxilium igitur assecutus a Deo usque in hodiernum diem sto testificans minori atque maiori, nihil extra dicens quam ea, quae Prophetae sunt locuti futura esse et Moyses:
ACTS|26|23|si passibilis Christus, si primus ex resurrectione mortuorum lumen annuntiaturus est populo et gentibus ".
ACTS|26|24|Sic autem eo rationem reddente, Festus magna voce dixit: " Insanis, Paule; multae te litterae ad insaniam convertunt! ".
ACTS|26|25|At Paulus: " Non insanio, inquit, optime Feste, sed veritatis et sobrietatis verba eloquor.
ACTS|26|26|Scit enim de his rex, ad quem et audenter loquor; latere enim eum nihil horum arbitror, neque enim in angulo hoc gestum est.
ACTS|26|27|Credis, rex Agrippa, Prophetis? Scio quia credis ".
ACTS|26|28|Agrippa autem ad Paulum: " In modico suades me Christianum fieri! ".
ACTS|26|29|Et Paulus: " Optarem apud Deum et in modico et in magno non tantum te sed et omnes hos, qui audiunt me hodie, fieri tales, qualis et ego sum, exceptis vinculis his! ".
ACTS|26|30|Et exsurrexit rex et praeses et Berenice et qui assidebant eis;
ACTS|26|31|et cum secessissent, loquebantur ad invicem dicentes: " Nihil morte aut vinculis dignum quid facit homo iste ".
ACTS|26|32|Agrippa autem Festo dixit: " Dimitti poterat homo hic, si non appellasset Caesarem ".
ACTS|27|1|Ut autem iudicatum est na vigare nos in Italiam, tradiderunt et Paulum et quosdam alios vinctos centurioni nomine Iulio, cohortis Augustae.
ACTS|27|2|Ascendentes autem navem Hadramyttenam, incipientem navigare circa Asiae loca, sustulimus, perseverante nobiscum Aristarcho Macedone Thessalonicensi;
ACTS|27|3|sequenti autem die, devenimus Sidonem, et humane tractans Iulius Paulum permisit ad amicos ire et curam sui agere.
ACTS|27|4|Et inde cum sustulissemus, subnavigavimus Cypro, propterea quod essent venti contrarii;
ACTS|27|5|et pelagus Ciliciae et Pamphyliae navigantes venimus Myram, quae est Lyciae.
ACTS|27|6|Et ibi inveniens centurio navem Alexandrinam navigantem in Italiam transposuit nos in eam.
ACTS|27|7|Et cum multis diebus tarde navigaremus et vix devenissemus contra Cnidum, prohibente nos vento, subnavigavimus Cretae secundum Salmonem;
ACTS|27|8|et vix iuxta eam navigantes venimus in locum quendam, qui vocatur Boni Portus, cui iuxta erat civitas Lasaea.
ACTS|27|9|Multo autem tempore peracto, et cum iam non esset tuta navigatio, eo quod et ieiunium iam praeterisset, monebat Paulus
ACTS|27|10|dicens eis: " Viri, video quoniam cum iniuria et multo damno non solum oneris et navis sed etiam animarum nostrarum incipit esse navigatio ".
ACTS|27|11|Centurio autem gubernatori et nauclero magis credebat quam his, quae a Paulo dicebantur.
ACTS|27|12|Et cum aptus portus non esset ad hiemandum, plurimi statuerunt consilium enavigare inde, si quo modo possent devenientes Phoenicen hiemare, portum Cretae respicientem ad africum et ad caurum.
ACTS|27|13|Aspirante autem austro, aestimantes propositum se tenere, cum sustulissent, propius legebant Cretam.
ACTS|27|14|Non post multum autem misit se contra ipsam ventus typhonicus, qui vocatur euroaquilo;
ACTS|27|15|cumque arrepta esset navis et non posset conari in ventum, data nave flatibus, ferebamur.
ACTS|27|16|Insulam autem quandam decurrentes, quae vocatur Cauda, potuimus vix obtinere scapham,
ACTS|27|17|qua sublata, adiutoriis utebantur accingentes navem; et timentes, ne in Syrtim inciderent, submisso vase, sic ferebantur.
ACTS|27|18|Valide autem nobis tempestate iactatis, sequenti die iactum fecerunt
ACTS|27|19|et tertia die suis manibus armamenta navis proiecerunt.
ACTS|27|20|Neque sole autem neque sideribus apparentibus per plures dies, et tempestate non exigua imminente, iam auferebatur spes omnis salutis nostrae.
ACTS|27|21|Et cum multa ieiunatio fuisset, tunc stans Paulus in medio eorum dixit: Oportebat quidem, o viri, audito me, non tollere a Creta lucrique facere iniuriam hanc et iacturam.
ACTS|27|22|Et nunc suadeo vobis bono animo esse, nulla enim amissio animae erit ex vobis praeterquam navis;
ACTS|27|23|astitit enim mihi hac nocte angelus Dei, cuius sum ego, cui et deservio,
ACTS|27|24|dicens: "Ne timeas, Paule; Caesari te oportet assistere, et ecce donavit tibi Deus omnes, qui navigant tecum".
ACTS|27|25|Propter quod bono animo estote, viri; credo enim Deo, quia sic erit, quemadmodum dictum est mihi.
ACTS|27|26|In insulam autem quandam oportet nos incidere ".
ACTS|27|27|Sed posteaquam quarta decima nox supervenit, cum ferremur in Hadria, circa mediam noctem suspicabantur nautae apparere sibi aliquam regionem.
ACTS|27|28|Qui submittentes bolidem invenerunt passus viginti; et pusillum inde separati et rursum submittentes invenerunt passus quindecim;
ACTS|27|29|timentes autem, ne in aspera loca incideremus, de puppi mittentes ancoras quattuor optabant diem fieri.
ACTS|27|30|Nautis vero quaerentibus fugere de navi, cum demisissent scapham in mare sub obtentu, quasi a prora inciperent ancoras extendere,
ACTS|27|31|dixit Paulus centurioni et militibus: " Nisi hi in navi manserint, vos salvi fieri non potestis ".
ACTS|27|32|Tunc absciderunt milites funes scaphae et passi sunt eam excidere.
ACTS|27|33|Donec autem lux inciperet fieri, rogabat Paulus omnes sumere cibum dicens: " Quarta decima hodie die exspectantes ieiuni permanetis nihil accipientes;
ACTS|27|34|propter quod rogo vos accipere cibum, hoc enim pro salute vestra est, quia nullius vestrum capillus de capite peribit ".
ACTS|27|35|Et cum haec dixisset et sumpsisset panem, gratias egit Deo in conspectu omnium et, cum fregisset, coepit manducare.
ACTS|27|36|Animaequiores autem facti omnes et ipsi assumpserunt cibum.
ACTS|27|37|Eramus vero universae animae in navi ducentae septuaginta sex.
ACTS|27|38|Et satiati cibo alleviabant navem iactantes triticum in mare.
ACTS|27|39|Cum autem dies factus esset, terram non agnoscebant; sinum vero quendam considerabant habentem litus, in quem cogitabant, si possent, eicere navem.
ACTS|27|40|Et cum ancoras abstulissent, committebant mari simul laxantes iuncturas gubernaculorum et, levato artemone, secundum flatum aurae tendebant ad litus.
ACTS|27|41|Et cum incidissent in locum dithalassum, impegerunt navem; et prora quidem fixa manebat immobilis, puppis vero solvebatur a vi fluctuum.
ACTS|27|42|Militum autem consilium fuit, ut custodias occiderent, ne quis, cum enatasset, effugeret;
ACTS|27|43|centurio autem volens servare Paulum prohibuit eos a consilio iussitque eos, qui possent natare, mittere se primos et ad terram exire
ACTS|27|44|et ceteros, quosdam in tabulis, quosdam vero super ea, quae de navi essent; et sic factum est ut omnes evaderent ad terram.
ACTS|28|1|Et cum evasissemus, tunc cognovimus quia Melita in sula vocatur.
ACTS|28|2|Barbari vero praestabant non modicam humanitatem nobis; accensa enim pyra, suscipiebant nos omnes propter imbrem, qui imminebat, et frigus.
ACTS|28|3|Cum congregasset autem Paulus sarmentorum aliquantam multitudinem et imposuisset super ignem, vipera, a calore cum processisset, invasit manum eius.
ACTS|28|4|Ut vero viderunt barbari pendentem bestiam de manu eius, ad invicem dicebant: " Utique homicida est homo hic, qui cum evaserit de mari, Ultio non permisit vivere ".
ACTS|28|5|Et ille quidem excutiens bestiam in ignem, nihil mali passus est;
ACTS|28|6|at illi exspectabant eum in tumorem convertendum aut subito casurum et mori. Diu autem illis exspectantibus et videntibus nihil mali in eo fieri, convertentes se dicebant eum esse deum.
ACTS|28|7|In locis autem illis erant praedia principis insulae nomine Publii, qui nos suscipiens triduo benigne hospitio recepit.
ACTS|28|8|Contigit autem patrem Publii febribus et dysenteria vexatum iacere, ad quem Paulus intravit et, cum orasset et imposuisset ei manus, sanavit eum.
ACTS|28|9|Quo facto, et ceteri, qui in insula habebant infirmitates, accedebant et curabantur;
ACTS|28|10|qui etiam multis honoribus nos honoraverunt et navigantibus imposuerunt, quae necessaria erant.
ACTS|28|11|Post menses autem tres, navigavimus in navi Alexandrina, quae in insula hiemaverat, cui erat insigne Castorum.
ACTS|28|12|Et cum venissemus Syracusam, mansimus ibi triduo;
ACTS|28|13|inde solventes devenimus Rhegium. Et post unum diem, superveniente austro, secunda die venimus Puteolos,
ACTS|28|14|ubi, inventis fratribus, rogati sumus manere apud eos dies septem; et sic venimus Romam.
ACTS|28|15|Et inde cum audissent de nobis fratres, occurrerunt nobis usque ad Appii Forum et Tres Tabernas; quos cum vidisset Paulus, gratias agens Deo, accepit fiduciam.
ACTS|28|16|Cum introissemus autem Romam, permissum est Paulo manere sibimet cum custodiente se milite.
ACTS|28|17|Factum est autem, ut post tertium diem convocaret primos Iudaeorum; cumque convenissent dicebat eis: " Ego, viri fratres, nihil adversus plebem faciens aut mores paternos, vinctus ab Hierosolymis traditus sum in manus Romanorum,
ACTS|28|18|qui cum interrogationem de me habuissent, volebant dimittere, eo quod nulla causa esset mortis in me;
ACTS|28|19|contradicentibus autem Iudaeis, coactus sum appellare Caesarem, non quasi gentem meam habens aliquid accusare.
ACTS|28|20|Propter hanc igitur causam rogavi vos videre et alloqui; propter spem enim Israel catena hac circumdatus sum ".
ACTS|28|21|At illi dixerunt ad eum: " Nos neque litteras accepimus de te a Iudaea, neque adveniens aliquis fratrum nuntiavit aut locutus est quid de te malum.
ACTS|28|22|Rogamus autem a te audire quae sentis; nam de secta hac notum est nobis quia ubique ei contradicitur ".
ACTS|28|23|Cum constituissent autem illi diem, venerunt ad eum in hospitium plures, quibus exponebat testificans regnum Dei suadensque eos de Iesu ex Lege Moysis et Prophetis a mane usque ad vesperam.
ACTS|28|24|Et quidam credebant his, quae dicebantur, quidam vero non credebant;
ACTS|28|25|cumque invicem non essent consentientes, discedebant, dicente Paulo unum verbum: " Bene Spiritus Sanctus locutus est per Isaiam prophetam ad patres vestros
ACTS|28|26|dicens:Vade ad populum istum et dic:Auditu audietis et non intellegetis,et videntes videbitis et non perspicietis.
ACTS|28|27|Incrassatum est enim cor populi huius,et auribus graviter audieruntet oculos suos compresserunt,ne forte videant oculiset auribus audiantet corde intellegant et convertantur,et sanabo illos".
ACTS|28|28|Notum ergo sit vobis quoniam gentibus missum est hoc salutare Dei; ipsi et audient! ".
ACTS|28|29|()
ACTS|28|30|Mansit autem biennio toto in suo conducto; et suscipiebat omnes, qui ingrediebantur ad eum,
ACTS|28|31|praedicans regnum Dei et docens quae sunt de Domino Iesu Christo cum omni fiducia sine prohibitione.
ROM|1|1|Paulus servus Christi Iesu, vo catus apostolus, segregatus in evangelium Dei,
ROM|1|2|quod ante promiserat per prophetas suos in Scripturis sanctis
ROM|1|3|de Filio suo, qui factus est ex semine David secundum carnem,
ROM|1|4|qui constitutus est Filius Dei in virtute secundum Spiritum sanctificationis ex resurrectione mortuorum, Iesu Christo Domino nostro,
ROM|1|5|per quem accepimus gratiam et apostolatum ad oboeditionem fidei in omnibus gentibus pro nomine eius,
ROM|1|6|in quibus estis et vos vocati Iesu Christi,
ROM|1|7|omnibus, qui sunt Romae dilectis Dei, vocatis sanctis: gratia vobis et pax a Deo Patre nostro et Domino Iesu Christo.
ROM|1|8|Primum quidem gratias ago Deo meo per Iesum Christum pro omnibus vobis, quia fides vestra annuntiatur in universo mundo;
ROM|1|9|testis enim mihi est Deus, cui servio in spiritu meo in evangelio Filii eius, quomodo sine intermissione memoriam vestri faciam
ROM|1|10|semper in orationibus meis obsecrans, si quo modo tandem aliquando prosperum iter habeam in voluntate Dei veniendi ad vos.
ROM|1|11|Desidero enim videre vos, ut aliquid impertiar gratiae vobis spiritalis ad confirmandos vos,
ROM|1|12|id est una vobiscum consolari per eam, quae invicem est, fidem vestram atque meam.
ROM|1|13|Nolo autem vos ignorare, fratres, quia saepe proposui venire ad vos et prohibitus sum usque adhuc, ut aliquem fructum habeam et in vobis, sicut et in ceteris gentibus.
ROM|1|14|Graecis ac barbaris, sapientibus et insipientibus debitor sum.
ROM|1|15|Itaque, quod in me est, promptus sum et vobis, qui Romae estis, evangelizare.
ROM|1|16|Non enim erubesco evangelium: virtus enim Dei est in salutem omni credenti, Iudaeo primum et Graeco.
ROM|1|17|Iustitia enim Dei in eo revelatur ex fide in fidem, sicut scriptum est: Iustus autem ex fide vivet ".
ROM|1|18|Revelatur enim ira Dei de caelo super omnem impietatem et iniustitiam hominum, qui veritatem in iniustitia detinent,
ROM|1|19|quia, quod noscibile est Dei, manifestum est in illis; Deus enim illis manifestavit.
ROM|1|20|Invisibilia enim ipsius a creatura mundi per ea, quae facta sunt, intellecta conspiciuntur, sempiterna eius et virtus et divinitas, ut sint inexcusabiles;
ROM|1|21|quia, cum cognovissent Deum, non sicut Deum glorificaverunt aut gratias egerunt, sed evanuerunt in cogitationibus suis, et obscuratum est insipiens cor eorum.
ROM|1|22|Dicentes se esse sapientes, stulti facti sunt,
ROM|1|23|et mutaverunt gloriam incorruptibilis Dei in similitudinem imaginis corruptibilis hominis et volucrum et quadrupedum et serpentium.
ROM|1|24|Propter quod tradidit illos Deus in concupiscentiis cordis eorum in immunditiam, ut ignominia afficiant corpora sua in semetipsis,
ROM|1|25|qui commutaverunt veritatem Dei in mendacio et coluerunt et servierunt creaturae potius quam Creatori, qui est benedictus in saecula. Amen.
ROM|1|26|Propterea tradidit illos Deus in passiones ignominiae. Nam et feminae eorum immutaverunt naturalem usum in eum, qui est contra naturam;
ROM|1|27|similiter et masculi, relicto naturali usu feminae, exarserunt in desideriis suis in invicem, masculi in masculos turpitudinem operantes et mercedem, quam oportuit, erroris sui in semetipsis recipientes.
ROM|1|28|Et sicut non probaverunt Deum habere in notitia, tradidit eos Deus in reprobum sensum, ut faciant, quae non conveniunt,
ROM|1|29|repletos omni iniquitate, malitia, avaritia, nequitia, plenos invidia, homicidio, contentione, dolo, malignitate, susurrones,
ROM|1|30|detractores, Deo odibiles, contumeliosos, superbos, elatos, inventores malorum, parentibus non oboedientes,
ROM|1|31|insipientes, incompositos, sine affectione, sine misericordia.
ROM|1|32|Qui cum iudicium Dei cognovissent, quoniam qui talia agunt, digni sunt morte, non solum ea faciunt, sed et consentiunt facientibus.
ROM|2|1|Propter quod inexcusabilis es, o homo omnis, qui iudicas. In quo enim iudicas alterum, teipsum condemnas; eadem enim agis, qui iudicas.
ROM|2|2|Scimus enim quoniam iudicium Dei est secundum veritatem in eos, qui talia agunt.
ROM|2|3|Existimas autem hoc, o homo, qui iudicas eos, qui talia agunt, et facis ea, quia tu effugies iudicium Dei?
ROM|2|4|An divitias benignitatis eius et patientiae et longanimitatis contemnis, ignorans quoniam benignitas Dei ad paenitentiam te adducit?
ROM|2|5|Secundum duritiam autem tuam et impaenitens cor thesaurizas tibi iram in die irae et revelationis iusti iudicii Dei,
ROM|2|6|qui reddet unicuique secundum opera eius:
ROM|2|7|his quidem, qui secundum patientiam boni operis gloriam et honorem et incorruptionem quaerunt, vitam aeternam;
ROM|2|8|his autem, qui ex contentione et non oboediunt veritati, oboediunt autem iniquitati, ira et indignatio.
ROM|2|9|Tribulatio et angustia in omnem animam hominis operantis malum, Iudaei primum et Graeci;
ROM|2|10|gloria autem et honor et pax omni operanti bonum, Iudaeo primum et Graeco.
ROM|2|11|Non est enim personarum acceptio apud Deum!
ROM|2|12|Quicumque enim sine lege peccaverunt, sine lege et peribunt; et, quicumque in lege peccaverunt, per legem iudicabuntur.
ROM|2|13|Non enim auditores legis iusti sunt apud Deum, sed factores legis iustificabuntur.
ROM|2|14|Cum enim gentes, quae legem non habent, naturaliter, quae legis sunt, faciunt, eiusmodi legem non habentes ipsi sibi sunt lex;
ROM|2|15|qui ostendunt opus legis scriptum in cordibus suis, testimonium simul reddente illis conscientia ipsorum, et inter se invicem cogitationibus accusantibus aut etiam defendentibus,
ROM|2|16|in die, cum iudicabit Deus occulta hominum secundum evangelium meum per Christum Iesum.
ROM|2|17|Si autem tu Iudaeus cognominaris et requiescis in lege et gloriaris in Deo,
ROM|2|18|et nosti Voluntatem et discernis potiora instructus per legem,
ROM|2|19|et confidis teipsum ducem esse caecorum, lumen eorum, qui in tenebris sunt,
ROM|2|20|eruditorem insipientium, magistrum infantium, habentem formam scientiae et veritatis in lege.
ROM|2|21|Qui ergo alium doces, teipsum non doces? Qui praedicas non furandum, furaris?
ROM|2|22|Qui dicis non moechandum, moecharis? Qui abominaris idola, templa spolias?
ROM|2|23|Qui in lege gloriaris, per praevaricationem legis Deum inhonoras?
ROM|2|24|" Nomen enim Dei propter vos blasphematur inter gentes ", sicut scriptum est.
ROM|2|25|Circumcisio quidem prodest, si legem observes; si autem praevaricator legis sis, circumcisio tua praeputium facta est.
ROM|2|26|Si igitur praeputium iustitias legis custodiat, nonne praeputium illius in circumcisionem reputabitur?
ROM|2|27|Et iudicabit, quod ex natura est praeputium legem consummans, te, qui per litteram et circumcisionem praevaricator legis es.
ROM|2|28|Non enim qui manifesto Iudaeus est, neque quae manifesto in carne circumcisio,
ROM|2|29|sed qui in abscondito Iudaeus est, et circumcisio cordis in spiritu non littera, cuius laus non ex hominibus sed ex Deo est.
ROM|3|1|Quid ergo amplius est Iudaeo, aut quae utilitas circumcisionis?
ROM|3|2|Multum per omnem modum. Primum quidem, quia credita sunt illis eloquia Dei.
ROM|3|3|Quid enim, si quidam non crediderunt? Numquid incredulitas illorum fidem Dei evacuabit?
ROM|3|4|Absit! Exstet autem Deus verax, omnis autem homo mendax, sicut scriptum est: " Ut iustificeris in sermonibus tuis et vincas cum iudicaris ".
ROM|3|5|Si autem iniustitia nostra iustitiam Dei commendat, quid dicemus? Numquid iniustus Deus, qui infert iram? Secundum hominem dico.
ROM|3|6|Absit! Alioquin quomodo iudicabit Deus mundum?
ROM|3|7|Si enim veritas Dei in meo mendacio abundavit in gloriam ipsius, quid adhuc et ego tamquam peccator iudicor?
ROM|3|8|Et non, sicut blasphemamur, et sicut aiunt quidam nos dicere: " Faciamus mala, ut veniant bona "? Quorum damnatio iusta est.
ROM|3|9|Quid igitur? Praecellimus eos? Nequaquam! Antea enim causati sumus Iudaeos et Graecos omnes sub peccato esse,
ROM|3|10|sicut scriptum est: Non est iustus quisquam,
ROM|3|11|non est intellegens, non est requirens Deum.
ROM|3|12|Omnes declinaverunt, simul inutiles facti sunt;non est qui faciat bonum, non est usque ad unum.
ROM|3|13|Sepulcrum patens est guttur eorum,linguis suis dolose agebant,venenum aspidum sub labiis eorum,
ROM|3|14|quorum os maledictione et amaritudine plenum est;
ROM|3|15|veloces pedes eorum ad effundendum sanguinem,
ROM|3|16|contritio et infelicitas in viis eorum,
ROM|3|17|et viam pacis non cognoverunt.
ROM|3|18|Non est timor Dei ante oculos eorum ".
ROM|3|19|Scimus autem quoniam, quaecumque lex loquitur, his, qui in lege sunt, loquitur, ut omne os obstruatur, et obnoxius fiat omnis mundus Deo;
ROM|3|20|quia ex operibus legis non iustificabitur omnis caro coram illo, per legem enim cognitio peccati.
ROM|3|21|Nunc autem sine lege iustitia Dei manifestata est, testificata a Lege et Prophetis,
ROM|3|22|iustitia autem Dei per fidem Iesu Christi, in omnes, qui credunt. Non enim est distinctio:
ROM|3|23|omnes enim peccaverunt et egent gloria Dei,
ROM|3|24|iustificati gratis per gratiam ipsius per redemptionem, quae est in Christo Iesu;
ROM|3|25|quem proposuit Deus propitiatorium per fidem in sanguine ipsius ad ostensionem iustitiae suae, cum praetermisisset praecedentia delicta
ROM|3|26|in sustentatione Dei, ad ostensionem iustitiae eius in hoc tempore, ut sit ipse iustus et iustificans eum, qui ex fide est Iesu.
ROM|3|27|Ubi est ergo gloriatio? Exclusa est. Per quam legem? Operum? Non, sed per legem fidei.
ROM|3|28|Arbitramur enim iustificari hominem per fidem sine operibus legis.
ROM|3|29|An Iudaeorum Deus tantum? Nonne et gentium? Immo et gentium,
ROM|3|30|quoniam quidem unus Deus, qui iustificabit circumcisionem ex fide et praeputium per fidem.
ROM|3|31|Legem ergo destruimus per fidem? Absit, sed legem statuimus.
ROM|4|1|Quid ergo dicemus invenisse Abraham progenitorem no strum secundum carnem?
ROM|4|2|Si enim Abraham ex operibus iustificatus est, habet gloriam sed non apud Deum.
ROM|4|3|Quid enim Scriptura dicit? " Credidit autem Abraham Deo, et reputatum est illi ad iustitiam ".
ROM|4|4|Ei autem, qui operatur, merces non reputatur secundum gratiam sed secundum debitum;
ROM|4|5|ei vero, qui non operatur, sed credit in eum, qui iustificat impium, reputatur fides eius ad iustitiam,
ROM|4|6|sicut et David dicit beatitudinem hominis, cui Deus reputat iustitiam sine operibus:
ROM|4|7|" Beati, quorum remissae sunt iniquitates,et quorum tecta sunt peccata.
ROM|4|8|Beatus vir, cui non imputabit Dominus peccatum ".
ROM|4|9|Beatitudo ergo haec in circumcisione an etiam in praeputio? Dicimus enim: " Reputata est Abrahae fides ad iustitiam ".
ROM|4|10|Quomodo ergo reputata est? In circumcisione an in praeputio? Non in circumcisione sed in praeputio:
ROM|4|11|et signum accepit circumcisionis, signaculum iustitiae fidei, quae fuit in praeputio, ut esset pater omnium credentium per praeputium, ut reputetur illis iustitia,
ROM|4|12|et pater circumcisionis his non tantum, qui ex circumcisione sunt, sed et qui sectantur vestigia eius, quae fuit in praeputio, fidei patris nostri Abrahae.
ROM|4|13|Non enim per legem promissio Abrahae aut semini eius, ut heres esset mundi, sed per iustitiam fidei;
ROM|4|14|si enim qui ex lege heredes sunt, exinanita est fides, et abolita est promissio.
ROM|4|15|Lex enim iram operatur; ubi autem non est lex, nec praevaricatio.
ROM|4|16|Ideo ex fide, ut secundum gratiam, ut firma sit promissio omni semini, non ei, qui ex lege est solum, sed et ei, qui ex fide est Abrahae - qui est pater omnium nostrum,
ROM|4|17|sicut scriptum est: " Patrem multarum gentium posui te " C, ante Deum, cui credidit, qui vivificat mortuos et vocat ea, quae non sunt, quasi sint;
ROM|4|18|qui contra spem in spe credidit, ut fieret pater multarum gentium, secundum quod dictum est: " Sic erit semen tuum ".
ROM|4|19|Et non infirmatus fide consideravit corpus suum iam emortuum, cum fere centum annorum esset, et emortuam vulvam Sarae;
ROM|4|20|in repromissione autem Dei non haesitavit diffidentia, sed confortatus est fide, dans gloriam Deo,
ROM|4|21|et plenissime sciens quia, quod promisit, potens est et facere.
ROM|4|22|Ideo et reputatum est illi ad iustitiam.
ROM|4|23|Non est autem scriptum tantum propter ipsum: reputatum est illi,
ROM|4|24|sed et propter nos, quibus reputabitur, credentibus in eum, qui suscitavit Iesum Dominum nostrum a mortuis,
ROM|4|25|qui traditus est propter delicta nostra et suscitatus est propter iustificationem nostram.
ROM|5|1|Iustificati igitur ex fide, pacem habemus ad Deum per Domi num nostrum Iesum Christum,
ROM|5|2|per quem et accessum habemus fide in gratiam istam, in qua stamus et gloriamur in spe gloriae Dei.
ROM|5|3|Non solum autem, sed et gloriamur in tribulationibus, scientes quod tribulatio patientiam operatur,
ROM|5|4|patientia autem probationem, probatio vero spem;
ROM|5|5|spes autem non confundit, quia caritas Dei diffusa est in cordibus nostris per Spiritum Sanctum, qui datus est nobis.
ROM|5|6|Adhuc enim Christus, cum adhuc infirmi essemus, secundum tempus pro impiis mortuus est.
ROM|5|7|Vix enim pro iusto quis moritur; nam pro bono forsitan quis et audeat mori.
ROM|5|8|Commendat autem suam caritatem Deus in nos, quoniam, cum adhuc peccatores essemus, Christus pro nobis mortuus est.
ROM|5|9|Multo igitur magis iustificati nunc in sanguine ipsius, salvi erimus ab ira per ipsum!
ROM|5|10|Si enim, cum inimici essemus, reconciliati sumus Deo per mortem Filii eius, multo magis reconciliati salvi erimus in vita ipsius;
ROM|5|11|non solum autem, sed et gloriamur in Deo per Dominum nostrum Iesum Christum, per quem nunc reconciliationem accepimus.
ROM|5|12|Propterea, sicut per unum hominem peccatum in hunc mundum intravit, et per peccatum mors, et ita in omnes homines mors pertransiit, eo quod omnes peccaverunt.
ROM|5|13|Usque ad legem enim peccatum erat in mundo; peccatum autem non imputatur, cum lex non est,
ROM|5|14|sed regnavit mors ab Adam usque ad Moysen etiam in eos, qui non peccaverunt in similitudine praevaricationis Adae, qui est figura futuri.
ROM|5|15|Sed non sicut delictum, ita et donum; si enim unius delicto multi mortui sunt, multo magis gratia Dei et donum in gratia unius hominis Iesu Christi in multos abundavit.
ROM|5|16|Et non sicut per unum, qui peccavit, ita et donum; nam iudicium ex uno in condemnationem, gratia autem ex multis delictis in iustificationem.
ROM|5|17|Si enim unius delicto mors regnavit per unum, multo magis, qui abundantiam gratiae et donationis iustitiae accipiunt, in vita regnabunt per unum Iesum Christum.
ROM|5|18|Igitur sicut per unius delictum in omnes homines in condemnationem, sic et per unius iustitiam in omnes homines in iustificationem vitae;
ROM|5|19|sicut enim per inoboedientiam unius hominis peccatores constituti sunt multi, ita et per unius oboeditionem iusti constituentur multi.
ROM|5|20|Lex autem subintravit, ut abundaret delictum; ubi autem abundavit peccatum, superabundavit gratia,
ROM|5|21|ut sicut regnavit peccatum in morte, ita et gratia regnet per iustitiam in vitam aeternam per Iesum Christum Dominum nostrum.
ROM|6|1|Quid ergo dicemus? Perma nebimus in peccato, ut gratia abundet?
ROM|6|2|Absit! Qui enim mortui sumus peccato, quomodo adhuc vivemus in illo?
ROM|6|3|An ignoratis quia, quicumque baptizati sumus in Christum Iesum, in mortem ipsius baptizati sumus?
ROM|6|4|Consepulti ergo sumus cum illo per baptismum in mortem, ut quemadmodum suscitatus est Christus a mortuis per gloriam Patris, ita et nos in novitate vitae ambulemus.
ROM|6|5|Si enim complantati facti sumus similitudini mortis eius, sed et resurrectionis erimus;
ROM|6|6|hoc scientes quia vetus homo noster simul crucifixus est, ut destruatur corpus peccati, ut ultra non serviamus peccato.
ROM|6|7|Qui enim mortuus est, iustificatus est a peccato.
ROM|6|8|Si autem mortui sumus cum Christo, credimus quia simul etiam vivemus cum eo;
ROM|6|9|scientes quod Christus suscitatus ex mortuis iam non moritur, mors illi ultra non dominatur.
ROM|6|10|Quod enim mortuus est, peccato mortuus est semel; quod autem vivit, vivit Deo.
ROM|6|11|Ita et vos existimate vos mortuos quidem esse peccato, viventes autem Deo in Christo Iesu.
ROM|6|12|Non ergo regnet peccatum in vestro mortali corpore, ut oboediatis concupiscentiis eius,
ROM|6|13|neque exhibeatis membra vestra arma iniustitiae peccato, sed exhibete vos Deo tamquam ex mortuis viventes et membra vestra arma iustitiae Deo.
ROM|6|14|Peccatum enim vobis non dominabitur; non enim sub lege estis sed sub gratia.
ROM|6|15|Quid ergo? Peccabimus, quoniam non sumus sub lege sed sub gratia? Absit!
ROM|6|16|Nescitis quoniam, cui exhibetis vos servos ad oboedientiam, servi estis eius, cui oboeditis, sive peccati ad mortem, sive oboeditionis ad iustitiam?
ROM|6|17|Gratias autem Deo quod fuistis servi peccati, oboedistis autem ex corde in eam formam doctrinae, in quam traditi estis,
ROM|6|18|liberati autem a peccato servi facti estis iustitiae.
ROM|6|19|Humanum dico propter infirmitatem carnis vestrae. Sicut enim exhibuistis membra vestra servientia immunditiae et iniquitati ad iniquitatem, ita nunc exhibete membra vestra servientia iustitiae ad sanctificationem.
ROM|6|20|Cum enim servi essetis peccati, liberi eratis iustitiae.
ROM|6|21|Quem ergo fructum habebatis tunc, in quibus nunc erubescitis? Nam finis illorum mors!
ROM|6|22|Nunc vero liberati a peccato, servi autem facti Deo, habetis fructum vestrum in sanctificationem, finem vero vitam aeternam!
ROM|6|23|Stipendia enim peccati mors, donum autem Dei vita aeterna in Christo Iesu Domino nostro.
ROM|7|1|An ignoratis, fratres - scienti bus enim legem loquor - quia lex in homine dominatur, quanto tempore vivit?
ROM|7|2|Nam quae sub viro est mulier, viventi viro alligata est lege; si autem mortuus fuerit vir, soluta est a lege viri.
ROM|7|3|Igitur, vivente viro, vocabitur adultera, si fuerit alterius viri; si autem mortuus fuerit vir, libera est a lege, ut non sit adultera, si fuerit alterius viri.
ROM|7|4|Itaque, fratres mei, et vos mortificati estis legi per corpus Christi, ut sitis alterius, eius qui ex mortuis suscitatus est, ut fructificaremus Deo.
ROM|7|5|Cum enim essemus in carne, passiones peccatorum, quae per legem sunt, operabantur in membris nostris, ut fructificarent morti;
ROM|7|6|nunc autem soluti sumus a lege, mortui ei, in qua detinebamur, ita ut serviamus in novitate Spiritus et non in vetustate litterae.
ROM|7|7|Quid ergo dicemus? Lex peccatum est? Absit! Sed peccatum non cognovi, nisi per legem; nam concupiscentiam nescirem, nisi lex diceret: " Non concupisces ".
ROM|7|8|Occasione autem accepta, peccatum per mandatum operatum est in me omnem concupiscentiam; sine lege enim peccatum mortuum erat.
ROM|7|9|Ego autem vivebam sine lege aliquando; sed, cum venisset mandatum, peccatum revixit,
ROM|7|10|ego autem mortuus sum; et inventum est mihi mandatum, quod erat ad vitam, hoc esse ad mortem;
ROM|7|11|nam peccatum, occasione accepta, per mandatum seduxit me et per illud occidit.
ROM|7|12|Itaque lex quidem sancta, et mandatum sanctum et iustum et bonum.
ROM|7|13|Quod ergo bonum est, mihi factum est mors? Absit! Sed peccatum, ut appareat peccatum, per bonum mihi operatum est mortem; ut fiat supra modum peccans peccatum per mandatum.
ROM|7|14|Scimus enim quod lex spiritalis est; ego autem carnalis sum, venumdatus sub peccato.
ROM|7|15|Quod enim operor, non intellego; non enim, quod volo, hoc ago, sed quod odi, illud facio.
ROM|7|16|Si autem, quod nolo, illud facio, consentio legi quoniam bona.
ROM|7|17|Nunc autem iam non ego operor illud, sed, quod habitat in me, peccatum.
ROM|7|18|Scio enim quia non habitat in me, hoc est in carne mea, bonum; nam velle adiacet mihi, operari autem bonum, non!
ROM|7|19|Non enim, quod volo bonum, facio, sed, quod nolo malum, hoc ago.
ROM|7|20|Si autem, quod nolo, illud facio, iam non ego operor illud, sed, quod habitat in me, peccatum.
ROM|7|21|Invenio igitur hanc legem volenti mihi facere bonum, quoniam mihi malum adiacet.
ROM|7|22|Condelector enim legi Dei secundum interiorem hominem;
ROM|7|23|video autem aliam legem in membris meis repugnantem legi mentis meae et captivantem me in lege peccati, quae est in membris meis.
ROM|7|24|Infelix ego homo! Quis me liberabit de corpore mortis huius?
ROM|7|25|Gratias autem Deo per Iesum Christum Dominum nostrum! Igitur ego ipse mente servio legi Dei, carne autem legi peccati.
ROM|8|1|Nihil ergo nunc damnationis est his, qui sunt in Christo Iesu;
ROM|8|2|lex enim Spiritus vitae in Christo Iesu liberavit te a lege peccati et mortis.
ROM|8|3|Nam, quod impossibile erat legi, in quo infirmabatur per carnem, Deus Filium suum mittens in similitudine carnis peccati et pro peccato, damnavit peccatum in carne,
ROM|8|4|ut iustitia legis impleretur in nobis, qui non secundum carnem ambulamus sed secundum Spiritum.
ROM|8|5|Qui enim secundum carnem sunt, quae carnis sunt, sapiunt; qui vero secundum Spiritum, quae sunt Spiritus.
ROM|8|6|Nam sapientia carnis mors, sapientia autem Spiritus vita et pax;
ROM|8|7|quoniam sapientia carnis inimicitia est in Deum, legi enim Dei non subicitur nec enim potest.
ROM|8|8|Qui autem in carne sunt, Deo placere non possunt.
ROM|8|9|Vos autem in carne non estis sed in Spiritu, si tamen Spiritus Dei habitat in vobis. Si quis autem Spiritum Christi non habet, hic non est eius.
ROM|8|10|Si autem Christus in vobis est, corpus quidem mortuum est propter peccatum, Spiritus vero vita propter iustitiam.
ROM|8|11|Quod si Spiritus eius, qui suscitavit Iesum a mortuis, habitat in vobis, qui suscitavit Christum a mortuis vivificabit et mortalia corpora vestra per inhabitantem Spiritum suum in vobis.
ROM|8|12|Ergo, fratres, debitores sumus non carni, ut secundum carnem vivamus.
ROM|8|13|Si enim secundum carnem vixeritis, moriemini; si autem Spiritu opera corporis mortificatis, vivetis.
ROM|8|14|Quicumque enim Spiritu Dei aguntur, hi filii Dei sunt.
ROM|8|15|Non enim accepistis spiritum servitutis iterum in timorem, sed accepistis Spiritum adoptionis filiorum, in quo clamamus: " Abba, Pater!.
ROM|8|16|Ipse Spiritus testimonium reddit una cum spiritu nostro, quod sumus filii Dei.
ROM|8|17|Si autem filii, et heredes: heredes quidem Dei, coheredes autem Christi, si tamen compatimur, ut et conglorificemur.
ROM|8|18|Existimo enim quod non sunt condignae passiones huius temporis ad futuram gloriam, quae revelanda est in nobis.
ROM|8|19|Nam exspectatio creaturae revelationem filiorum Dei exspectat;
ROM|8|20|vanitati enim creatura subiecta est, non volens sed propter eum, qui subiecit, in spem,
ROM|8|21|quia et ipsa creatura liberabitur a servitute corruptionis in libertatem gloriae filiorum Dei.
ROM|8|22|Scimus enim quod omnis creatura congemiscit et comparturit usque adhuc;
ROM|8|23|non solum autem, sed et nos ipsi primitias Spiritus habentes, et ipsi intra nos gemimus adoptionem filiorum exspectantes, redemptionem corporis nostri.
ROM|8|24|Spe enim salvi facti sumus; spes autem, quae videtur, non est spes; nam, quod videt, quis sperat?
ROM|8|25|Si autem, quod non videmus, speramus, per patientiam exspectamus.
ROM|8|26|Similiter autem et Spiritus adiuvat infirmitatem nostram; nam quid oremus, sicut oportet, nescimus, sed ipse Spiritus interpellat gemitibus inenarrabilibus;
ROM|8|27|qui autem scrutatur corda, scit quid desideret Spiritus, quia secundum Deum postulat pro sanctis.
ROM|8|28|Scimus autem quoniam diligentibus Deum omnia cooperantur in bonum, his, qui secundum propositum vocati sunt.
ROM|8|29|Nam, quos praescivit, et praedestinavit conformes fieri imaginis Filii eius, ut sit ipse primogenitus in multis fratribus;
ROM|8|30|quos autem praedestinavit, hos et vocavit; et quos vocavit, hos et iustificavit; quos autem iustificavit, illos et glorificavit.
ROM|8|31|Quid ergo dicemus ad haec? Si Deus pro nobis, quis contra nos?
ROM|8|32|Qui Filio suo non pepercit, sed pro nobis omnibus tradidit illum, quomodo non etiam cum illo omnia nobis donabit?
ROM|8|33|Quis accusabit adversus electos Dei? Deus, qui iustificat?
ROM|8|34|Quis est qui condemnet? Christus Iesus, qui mortuus est, immo qui suscitatus est, qui et est ad dexteram Dei, qui etiam interpellat pro nobis?
ROM|8|35|Quis nos separabit a caritate Christi? Tribulatio an angustia an persecutio an fames an nuditas an periculum an gladius?
ROM|8|36|Sicut scriptum est: Propter te mortificamur tota die,aestimati sumus ut oves occisionis ".
ROM|8|37|Sed in his omnibus supervincimus per eum, qui dilexit nos.
ROM|8|38|Certus sum enim quia neque mors neque vita neque angeli neque principatus neque instantia neque futura neque virtutes
ROM|8|39|neque altitudo neque profundum neque alia quaelibet creatura poterit nos separare a caritate Dei, quae est in Christo Iesu Domino nostro.
ROM|9|1|Veritatem dico in Christo, non mentior, testimonium mihi per hibente conscientia mea in Spiritu Sancto,
ROM|9|2|quoniam tristitia est mihi magna, et continuus dolor cordi meo.
ROM|9|3|Optarem enim ipse ego anathema esse a Christo pro fratribus meis, cognatis meis secundum carnem,
ROM|9|4|qui sunt Israelitae, quorum adoptio est filiorum et gloria et testamenta et legislatio et cultus et promissiones,
ROM|9|5|quorum sunt patres, et ex quibus Christus secundum carnem: qui est super omnia Deus benedictus in saecula. Amen.
ROM|9|6|Non autem quod exciderit verbum Dei. Non enim omnes, qui ex Israel, hi sunt Israel;
ROM|9|7|neque quia semen sunt Abrahae, omnes filii, sed: " In Isaac vocabitur tibi semen ".
ROM|9|8|Id est, non qui filii carnis, hi filii Dei, sed qui filii sunt promissionis, aestimantur semen;
ROM|9|9|promissionis enim verbum hoc est: " Secundum hoc tempus veniam, et erit Sarae filius ".
ROM|9|10|Non solum autem, sed et Rebecca ex uno concubitum habens, Isaac patre nostro;
ROM|9|11|cum enim nondum nati fuissent aut aliquid egissent bonum aut malum, ut secundum electionem propositum Dei maneret,
ROM|9|12|non ex operibus sed ex vocante dictum est ei: " Maior serviet minori ";
ROM|9|13|sicut scriptum est: " Iacob dilexi, Esau autem odio habui ".
ROM|9|14|Quid ergo dicemus? Numquid iniustitia apud Deum? Absit!
ROM|9|15|Moysi enim dicit: " Miserebor, cuius misereor, et misericordiam praestabo, cui misericordiam praesto ".
ROM|9|16|Igitur non volentis neque currentis sed miserentis Dei.
ROM|9|17|Dicit enim Scriptura pharaoni: " In hoc ipsum excitavi te, ut ostendam in te virtutem meam, et ut annuntietur nomen meum in universa terra ".
ROM|9|18|Ergo, cuius vult, miseretur et, quem vult, indurat.
ROM|9|19|Dices itaque mihi: " Quid ergo adhuc queritur? Voluntati enim eius quis restitit? ".
ROM|9|20|O homo, sed tu quis es, qui respondeas Deo? Numquid dicet figmentum ei, qui se finxit: " Quid me fecisti sic? ".
ROM|9|21|An non habet potestatem figulus luti ex eadem massa facere aliud quidem vas in honorem, aliud vero in ignominiam?
ROM|9|22|Quod si volens Deus ostendere iram et notam facere potentiam suam, sustinuit in multa patientia vasa irae aptata in interitum;
ROM|9|23|et ut ostenderet divitias gloriae suae in vasa misericordiae, quae praeparavit in gloriam,
ROM|9|24|quos et vocavit nos non solum ex Iudaeis sed etiam ex gentibus?
ROM|9|25|Sicut et in Osee dicit: Vocabo Non plebem meam Plebem meamet Non dilectam Dilectam.
ROM|9|26|Et erit: in loco, ubi dictum est eis:Non plebs mea vos",ibi vocabuntur Filii Dei vivi ".
ROM|9|27|Isaias autem clamat pro Israel: " Si fuerit numerus filiorum Israel tamquam arena maris, reliquiae salvae fient.
ROM|9|28|Verbum enim consummans et brevians faciet Dominus super terram ".
ROM|9|29|Et sicut praedixit Isaias: Nisi Dominus Sabaoth reliquisset nobis semen,sicut Sodoma facti essemuset sicut Gomorra similes fuissemus ".
ROM|9|30|Quid ergo dicemus? Quod gentes, quae non sectabantur iustitiam, apprehenderunt iustitiam, iustitiam autem, quae ex fide est;
ROM|9|31|Israel vero sectans legem iustitiae in legem non pervenit.
ROM|9|32|Quare? Quia non ex fide sed quasi ex operibus; offenderunt in lapidem offensionis,
ROM|9|33|sicut scriptum est: Ecce pono in Sion lapidem offensionis et petram scandali;et, qui credit in eo, non confundetur ".
ROM|10|1|Fratres, voluntas quidem cordis mei et obsecratio ad Deum pro illis in salutem.
ROM|10|2|Testimonium enim perhibeo illis quod aemulationem Dei habent sed non secundum scientiam;
ROM|10|3|ignorantes enim Dei iustitiam et suam iustitiam quaerentes statuere, iustitiae Dei non sunt subiecti;
ROM|10|4|finis enim legis Christus ad iustitiam omni credenti.
ROM|10|5|Moyses enim scribit de iustitia, quae ex lege est: " Qui fecerit homo, vivet in eis ".
ROM|10|6|Quae autem ex fide est iustitia, sic dicit: " Ne dixeris in corde tuo: Quis ascendet in caelum?", id est Christum deducere;
ROM|10|7|aut: " Quis descendet in abyssum? ", hoc est Christum ex mortuis revocare.
ROM|10|8|Sed quid dicit? " Prope te est verbum, in ore tuo et in corde tuo "; hoc est verbum fidei, quod praedicamus.
ROM|10|9|Quia si confitearis in ore tuo: " Dominum Iesum! ", et in corde tuo credideris quod Deus illum excitavit ex mortuis, salvus eris.
ROM|10|10|Corde enim creditur ad iustitiam, ore autem confessio fit in salutem.
ROM|10|11|Dicit enim Scriptura: Omnis, qui credit in illo, non confundetur ".
ROM|10|12|Non enim est distinctio Iudaei et Graeci, nam idem Dominus omnium, dives in omnes, qui invocant illum:
ROM|10|13|Omnis enim, quicumque invocaverit nomen Domini, salvus erit.
ROM|10|14|Quomodo ergo invocabunt, in quem non crediderunt? Aut quomodo credent ei, quem non audierunt? Quomodo autem audient sine praedicante?
ROM|10|15|Quomodo vero praedicabunt nisi mittantur? Sicut scriptum est: Quam speciosi pedes evangelizantium bona ".
ROM|10|16|Sed non omnes oboedierunt evangelio; Isaias enim dicit: Domine, quis credidit auditui nostro? ".
ROM|10|17|Ergo fides ex auditu, auditus autem per verbum Christi.
ROM|10|18|Sed dico: Numquid non audierunt? Quin immo,in omnem terram exiit sonus eorum,et in fines orbis terrae verba eorum.
ROM|10|19|Sed dico: Numquid Israel non cognovit? Primus Moyses dicit: Ego ad aemulationem vos adducam per Non gentem:per gentem insipientem ad iram vos provocabo ".
ROM|10|20|Isaias autem audet et dicit: " Inventus sum in non quaerentibus me; palam apparui his, qui me non interrogabant ".
ROM|10|21|Ad Israel autem dicit: " Tota die expandi manus meas ad populum non credentem et contradicentem ".
ROM|11|1|Dico ergo: Numquid repulit Deus populum suum? Absit! Nam et ego Israelita sum, ex semine Abraham, tribu Beniamin.
ROM|11|2|Non reppulit Deus plebem suam, quam praescivit. An nescitis in Elia quid dicit Scriptura? Quemadmodum interpellat Deum adversus Israel:
ROM|11|3|" Domine, prophetas tuos occiderunt, altaria tua suffoderunt, et ego relictus sum solus, et quaerunt animam meam ".
ROM|11|4|Sed quid dicit illi responsum divinum? Reliqui mihi septem milia virorum, qui non curvaverunt genu Baal ".
ROM|11|5|Sic ergo et in hoc tempore reliquiae secundum electionem gratiae factae sunt.
ROM|11|6|Si autem gratia, iam non ex operibus, alioquin gratia iam non est gratia.
ROM|11|7|Quid ergo? Quod quaerit Israel, hoc non est consecutus, electio autem consecuta est; ceteri vero excaecati sunt,
ROM|11|8|sicut scriptum est: Dedit illis Deus spiritum soporis,oculos, ut non videant,et aures, ut non audiant,usque in hodiernum diem ".
ROM|11|9|Et David dicit: Fiat mensa eorum in laqueum et in captionemet in scandalum et in retributionem illis.
ROM|11|10|Obscurentur oculi eorum, ne videant,et dorsum illorum semper incurva! ".
ROM|11|11|Dico ergo: Numquid sic offenderunt, ut caderent? Absit! Sed illorum casu salus gentibus, ut illi ad aemulationem adducantur.
ROM|11|12|Quod si casus illorum divitiae sunt mundi, et deminutio eorum divitiae gentium, quanto magis plenitudo eorum!
ROM|11|13|Vobis autem dico gentibus: Quantum quidem ego sum gentium apostolus, ministerium meum honorifico,
ROM|11|14|si quo modo ad aemulandum provocem carnem meam et salvos faciam aliquos ex illis.
ROM|11|15|Si enim amissio eorum reconciliatio est mundi, quae assumptio, nisi vita ex mortuis?
ROM|11|16|Quod si primitiae sanctae sunt, et massa; et si radix sancta, et rami.
ROM|11|17|Quod si aliqui ex ramis fracti sunt, tu autem, cum oleaster esses, insertus es in illis et consocius radicis pinguedinis olivae factus es,
ROM|11|18|noli gloriari adversus ramos; quod si gloriaris, non tu radicem portas, sed radix te.
ROM|11|19|Dices ergo: " Fracti sunt rami, ut ego inserar ".
ROM|11|20|Bene; incredulitate fracti sunt, tu autem fide stas. Noli altum sapere, sed time:
ROM|11|21|si enim Deus naturalibus ramis non pepercit, ne forte nec tibi parcat.
ROM|11|22|Vide ergo bonitatem et severitatem Dei: in eos quidem, qui ceciderunt, severitatem; in te autem bonitatem Dei, si permanseris in bonitate, alioquin et tu excideris.
ROM|11|23|Sed et illi, si non permanserint in incredulitate, inserentur; potens est enim Deus iterum inserere illos!
ROM|11|24|Nam si tu ex naturali excisus es oleastro et contra naturam insertus es in bonam olivam, quanto magis hi, qui secundum naturam sunt, inserentur suae olivae.
ROM|11|25|Nolo enim vos ignorare, fratres, mysterium hoc, ut non sitis vobis ipsis sapientes, quia caecitas ex parte contigit in Israel, donec plenitudo gentium intraret,
ROM|11|26|et sic omnis Israel salvus fiet, sicut scriptum est: Veniet ex Sion, qui eripiat,avertet impietates ab Iacob;
ROM|11|27|et hoc illis a me testamentum,cum abstulero peccata eorum ".
ROM|11|28|Secundum evangelium quidem inimici propter vos, secundum electionem autem carissimi propter patres;
ROM|11|29|sine paenitentia enim sunt dona et vocatio Dei!
ROM|11|30|Sicut enim aliquando vos non credidistis Deo, nunc autem misericordiam consecuti estis propter illorum incredulitatem,
ROM|11|31|ita et isti nunc non crediderunt propter vestram misericordiam, ut et ipsi nunc misericordiam consequantur.
ROM|11|32|Conclusit enim Deus omnes in incredulitatem, ut omnium misereatur!
ROM|11|33|O altitudo divitiarum et sapientiae et scientiae Dei! Quam incomprehensibilia sunt iudicia eius, et investigabiles viae eius!
ROM|11|34|Quis enim cognovit sensum Domini?Aut quis consiliarius eius fuit?
ROM|11|35|Aut quis prior dedit illi,et retribuetur ei?
ROM|11|36|Quoniam ex ipso et per ipsum et in ipsum omnia. Ipsi gloria in saecula. Amen.
ROM|12|1|Obsecro itaque vos, fratres, per misericordiam Dei, ut exhibeatis corpora vestra hostiam viventem, sanctam, Deo placentem, rationabile obsequium vestrum;
ROM|12|2|et nolite conformari huic saeculo, sed transformamini renovatione mentis, ut probetis quid sit voluntas Dei, quid bonum et bene placens et perfectum.
ROM|12|3|Dico enim per gratiam, quae data est mihi, omnibus, qui sunt inter vos, non altius sapere quam oportet sapere, sed sapere ad sobrietatem, unicuique sicut Deus divisit mensuram fidei.
ROM|12|4|Sicut enim in uno corpore multa membra habemus, omnia autem membra non eundem actum habent,
ROM|12|5|ita multi unum corpus sumus in Christo, singuli autem alter alterius membra.
ROM|12|6|Habentes autem donationes secundum gratiam, quae data est nobis, differentes: sive prophetiam, secundum rationem fidei;
ROM|12|7|sive ministerium, in ministrando; sive qui docet, in doctrina;
ROM|12|8|sive qui exhortatur, in exhortando; qui tribuit, in simplicitate; qui praeest, in sollicitudine; qui miseretur, in hilaritate.
ROM|12|9|Dilectio sine simulatione. Odientes malum, adhaerentes bono;
ROM|12|10|caritate fraternitatis invicem diligentes, honore invicem praevenientes,
ROM|12|11|sollicitudine non pigri, spiritu ferventes, Domino servientes,
ROM|12|12|spe gaudentes, in tribulatione patientes, orationi instantes,
ROM|12|13|necessitatibus sanctorum communicantes, hospitalitatem sectantes.
ROM|12|14|Benedicite persequentibus; benedicite et nolite maledicere!
ROM|12|15|Gaudere cum gaudentibus, flere cum flentibus.
ROM|12|16|Idipsum invicem sentientes, non alta sapientes, sed humilibus consentientes. Nolite esse prudentes apud vosmetipsos.
ROM|12|17|Nulli malum pro malo reddentes; providentes bona coram omnibus hominibus;
ROM|12|18|si fieri potest, quod ex vobis est, cum omnibus hominibus pacem habentes;
ROM|12|19|non vosmetipsos vindicantes, carissimi, sed date locum irae, scriptum est enim: " Mihi vindicta, ego retribuam ", dicit Dominus.
ROM|12|20|Sed si esurierit inimicus tuus, ciba illum; si sitit, potum da illi. Hoc enim faciens, carbones ignis congeres super caput eius.
ROM|12|21|Noli vinci a malo, sed vince in bono malum.
ROM|13|1|Omnis anima potestatibus sublimioribus subdita sit. Non est enim potestas nisi a Deo; quae autem sunt, a Deo ordinatae sunt.
ROM|13|2|Itaque, qui resistit potestati, Dei ordinationi resistit; qui autem resistunt ipsi, sibi damnationem acquirent.
ROM|13|3|Nam principes non sunt timori bono operi sed malo. Vis autem non timere potestatem? Bonum fac, et habebis laudem ex illa;
ROM|13|4|Dei enim ministra est tibi in bonum. Si autem malum feceris, time; non enim sine causa gladium portat; Dei enim ministra est, vindex in iram ei, qui malum agit.
ROM|13|5|Ideo necesse est subditos esse, non solum propter iram sed et propter conscientiam.
ROM|13|6|Ideo enim et tributa praestatis; ministri enim Dei sunt in hoc ipsum instantes.
ROM|13|7|Reddite omnibus debita: cui tributum tributum, cui vectigal vectigal, cui timorem timorem, cui honorem honorem.
ROM|13|8|Nemini quidquam debeatis, nisi ut invicem diligatis: qui enim diligit proximum, legem implevit.
ROM|13|9|Nam: Non adulterabis, Non occides, Non furaberis, Non concupisces, et si quod est aliud mandatum, in hoc verbo recapitulatur: Diliges proximum tuum tamquam teipsum.
ROM|13|10|Dilectio proximo malum non operatur; plenitudo ergo legis est dilectio.
ROM|13|11|Et hoc scientes tempus, quia hora est iam vos de somno surgere; nunc enim propior est nobis salus quam cum credidimus.
ROM|13|12|Nox processit, dies autem appropiavit. Abiciamus ergo opera tenebrarum et induamur arma lucis.
ROM|13|13|Sicut in die honeste ambulemus: non in comissationibus et ebrietatibus, non in cubilibus et impudicitiis, non in contentione et aemulatione;
ROM|13|14|sed induite Dominum Iesum Christum et carnis curam ne feceritis in concupiscentiis.
ROM|14|1|Infirmum autem in fide assumite, non in disceptatio nibus cogitationum.
ROM|14|2|Alius enim credit manducare omnia; qui autem infirmus est, holus manducat.
ROM|14|3|Is qui manducat, non manducantem non spernat; et, qui non manducat, manducantem non iudicet, Deus enim illum assumpsit.
ROM|14|4|Tu quis es, qui iudices alienum servum? Suo domino stat aut cadit; stabit autem, potens est enim Dominus statuere illum.
ROM|14|5|Nam alius iudicat inter diem et diem, alius iudicat omnem diem; unusquisque in suo sensu abundet.
ROM|14|6|Qui sapit diem, Domino sapit; et, qui manducat, Domino manducat, gratias enim agit Deo; et, qui non manducat, Domino non manducat et gratias agit Deo.
ROM|14|7|Nemo enim nostrum sibi vivit, et nemo sibi moritur;
ROM|14|8|sive enim vivimus, Domino vivimus, sive morimur, Domino morimur. Sive ergo vivimus, sive morimur, Domini sumus.
ROM|14|9|In hoc enim Christus et mortuus est et vixit, ut et mortuorum et vivorum dominetur.
ROM|14|10|Tu autem, quid iudicas fratrem tuum? Aut tu, quare spernis fratrem tuum? Omnes enim stabimus ante tribunal Dei;
ROM|14|11|scriptum est enim: Vivo ego, dicit Dominus,mihi flectetur omne genu,et omnis lingua confitebitur Deo ".
ROM|14|12|Itaque unusquisque nostrum pro se rationem reddet Deo.
ROM|14|13|Non ergo amplius invicem iudicemus, sed hoc iudicate magis, ne ponatis offendiculum fratri vel scandalum.
ROM|14|14|Scio et certus sum in Domino Iesu, quia nihil commune per seipsum, nisi ei, qui existimat quid commune esse, illi commune est.
ROM|14|15|Si enim propter cibum frater tuus contristatur, iam non secundum caritatem ambulas. Noli cibo tuo illum perdere, pro quo Christus mortuus est!
ROM|14|16|Non ergo blasphemetur bonum vestrum!
ROM|14|17|Non est enim regnum Dei esca et potus, sed iustitia et pax et gaudium in Spiritu Sancto;
ROM|14|18|qui enim in hoc servit Christo, placet Deo et probatus est hominibus.
ROM|14|19|Itaque, quae pacis sunt, sectemur et quae aedificationis sunt in invicem.
ROM|14|20|Noli propter escam destruere opus Dei! Omnia quidem munda sunt, sed malum est homini, qui per offendiculum manducat.
ROM|14|21|Bonum est non manducare carnem et non bibere vinum neque id, in quo frater tuus offendit.
ROM|14|22|Tu, quam fidem habes, penes temetipsum habe coram Deo. Beatus, qui non iudicat semetipsum in eo quod probat.
ROM|14|23|Qui autem discernit si manducaverit, damnatus est, quia non ex fide; omne autem, quod non ex fide, peccatum est.
ROM|15|1|Debemus autem nos fir miores imbecillitates infir morum sustinere et non nobis placere.
ROM|15|2|Unusquisque nostrum proximo placeat in bonum ad aedificationem;
ROM|15|3|etenim Christus non sibi placuit, sed sicut scriptum est: " Improperia improperantium tibi ceciderunt super me ".
ROM|15|4|Quaecumque enim antea scripta sunt, ad nostram doctrinam scripta sunt, ut per patientiam et consolationem Scripturarum spem habeamus.
ROM|15|5|Deus autem patientiae et solacii det vobis idipsum sapere in alterutrum secundum Christum Iesum,
ROM|15|6|ut unanimes uno ore glorificetis Deum et Patrem Domini nostri Iesu Christi.
ROM|15|7|Propter quod suscipite invicem, sicut et Christus suscepit vos, in gloriam Dei.
ROM|15|8|Dico enim Christum ministrum fuisse circumcisionis propter veritatem Dei ad confirmandas promissiones patrum;
ROM|15|9|gentes autem propter misericordiam glorificare Deum, sicut scriptum est: Propter hoc confitebor tibi in gentibus et nomini tuo cantabo ".
ROM|15|10|Et iterum dicit: " Laetamini, gentes, cum plebe eius ".
ROM|15|11|Et iterum: Laudate, omnes gentes, Dominum,et magnificent eum omnes populi ".
ROM|15|12|Et rursus Isaias ait: Erit radix Iesse,et qui exsurget regere gentes:in eo gentes sperabunt ".
ROM|15|13|Deus autem spei repleat vos omni gaudio et pace in credendo, ut abundetis in spe in virtute Spiritus Sancti.
ROM|15|14|Certus sum autem, fratres mei, et ego ipse de vobis, quoniam et ipsi pleni estis bonitate, repleti omni scientia, ita ut possitis et alterutrum monere.
ROM|15|15|Audacius autem scripsi vobis ex parte, tamquam in memoriam vos reducens propter gratiam, quae data est mihi a Deo,
ROM|15|16|ut sim minister Christi Iesu ad gentes, consecrans evangelium Dei, ut fiat oblatio gentium accepta, sanctificata in Spiritu Sancto.
ROM|15|17|Habeo igitur gloriationem in Christo Iesu ad Deum;
ROM|15|18|non enim audebo aliquid loqui eorum, quae per me non effecit Christus in oboedientiam gentium, verbo et factis,
ROM|15|19|in virtute signorum et prodigiorum, in virtute Spiritus, ita ut ab Ierusalem et per circuitum usque in Illyricum repleverim evangelium Christi,
ROM|15|20|sic autem contendens praedicare evangelium, non ubi nominatus est Christus, ne super alienum fundamentum aedificarem,
ROM|15|21|sed sicut scriptum est: Quibus non est annuntiatum de eo, videbunt;et, qui non audierunt, intellegent ".
ROM|15|22|Propter quod et impediebar plurimum venire ad vos;
ROM|15|23|nunc vero ulterius locum non habens in his regionibus, cupiditatem autem habens veniendi ad vos ex multis iam annis,
ROM|15|24|cum in Hispaniam proficisci coepero, spero enim quod praeteriens videam vos et a vobis deducar illuc, si vobis primum ex parte fruitus fuero.
ROM|15|25|Nunc autem proficiscor in Ierusalem ministrare sanctis;
ROM|15|26|probaverunt enim Macedonia et Achaia communicationem aliquam facere in pauperes sanctorum, qui sunt in Ierusalem.
ROM|15|27|Placuit enim eis, et debitores sunt eorum; nam si spiritalibus eorum communicaverunt gentes, debent et in carnalibus ministrare eis.
ROM|15|28|Hoc igitur cum consummavero et assignavero eis fructum hunc, proficiscar per vos in Hispaniam;
ROM|15|29|scio autem quoniam veniens ad vos, in abundantia benedictionis Christi veniam.
ROM|15|30|Obsecro autem vos, fratres, per Dominum nostrum Iesum Christum et per caritatem Spiritus, ut concertemini mecum in orationibus pro me ad Deum,
ROM|15|31|ut liberer ab infidelibus, qui sunt in Iudaea, et ministerium meum pro Ierusalem acceptum sit sanctis,
ROM|15|32|ut veniens ad vos in gaudio per voluntatem Dei refrigerer vobiscum.
ROM|15|33|Deus autem pacis sit cum omnibus vobis. Amen.
ROM|16|1|Commendo autem vobis Phoebem sororem nostram, quae est ministra ecclesiae, quae est Cenchreis,
ROM|16|2|ut eam suscipiatis in Domino digne sanctis et assistatis ei in quocumque negotio vestri indiguerit; etenim ipsa astitit multis et mihi ipsi.
ROM|16|3|Salutate Priscam et Aquilam adiutores meos in Christo Iesu,
ROM|16|4|qui pro anima mea suas cervices supposuerunt, quibus non solus ego gratias ago sed et cunctae ecclesiae gentium;
ROM|16|5|et domesticam eorum ecclesiam.Salutate Epaenetum dilectum mihi, primitias Asiae in Christo.
ROM|16|6|Salutate Mariam, quae multum laboravit in vobis.
ROM|16|7|Salutate Andronicum et Iuniam cognatos meos et concaptivos meos, qui sunt nobiles in apostolis, qui et ante me fuerunt in Christo.
ROM|16|8|Salutate Ampliatum dilectissimum mihi in Domino.
ROM|16|9|Salutate Urbanum adiutorem nostrum in Christo et Stachyn dilectum meum.
ROM|16|10|Salutate Apellem probatum in Christo. Salutate eos, qui sunt ex Aristobuli.
ROM|16|11|Salutate Herodionem cognatum meum. Salutate eos, qui sunt ex Narcissi, qui sunt in Domino.
ROM|16|12|Salutate Tryphaenam et Tryphosam, quae laborant in Domino. Salutate Persidam carissimam, quae multum laboravit in Domino.
ROM|16|13|Salutate Rufum electum in Domino et matrem eius et meam.
ROM|16|14|Salutate Asyncritum, Phlegonta, Hermen, Patrobam, Hermam et, qui cum eis sunt, fratres.
ROM|16|15|Salutate Philologum et Iuliam, Nereum et sororem eius et Olympam et omnes, qui cum eis sunt, sanctos.
ROM|16|16|Salutate invicem in osculo sancto. Salutant vos omnes ecclesiae Christi.
ROM|16|17|Rogo autem vos, fratres, ut observetis eos, qui dissensiones et offendicula praeter doctrinam, quam vos didicistis, faciunt, et declinate ab illis;
ROM|16|18|huiusmodi enim Domino nostro Christo non serviunt sed suo ventri, et per dulces sermones et benedictiones seducunt corda innocentium.
ROM|16|19|Vestra enim oboedientia ad omnes pervenit; gaudeo igitur in vobis, sed volo vos sapientes esse in bono et simplices in malo.
ROM|16|20|Deus autem pacis conteret Satanam sub pedibus vestris velociter.Gratia Domini nostri Iesu vobiscum.
ROM|16|21|Salutat vos Timotheus adiutor meus et Lucius et Iason et Sosipater cognati mei.
ROM|16|22|Saluto vos ego Tertius, qui scripsi epistulam in Domino.
ROM|16|23|Salutat vos Gaius hospes meus et universae ecclesiae. Salutat vos Erastus arcarius civitatis et Quartus frater.
ROM|16|24|()
ROM|16|25|Ei autem, qui potens est vos confirmare iuxta evangelium meum et praedicationem Iesu Christi secundum revelationem mysterii temporibus aeternis taciti,
ROM|16|26|manifestati autem nunc, et per scripturas Prophetarum secundum praeceptum aeterni Dei ad oboeditionem fidei in cunctis gentibus patefacti,
ROM|16|27|soli sapienti Deo per Iesum Christum, cui gloria in saecula. Amen.
1COR|1|1|Paulus, vocatus apostolus Christi Iesu per voluntatem Dei, et Sosthenes frater
1COR|1|2|ecclesiae Dei, quae est Corinthi, sanctificatis in Christo Iesu, vocatis sanctis cum omnibus, qui invocant nomen Domini nostri Iesu Christi in omni loco ipsorum et nostro:
1COR|1|3|gratia vobis et pax a Deo Patre nostro et Domino Iesu Christo.
1COR|1|4|Gratias ago Deo meo semper pro vobis in gratia Dei, quae data est vobis in Christo Iesu,
1COR|1|5|quia in omnibus divites facti estis in illo, in omni verbo et in omni scientia,
1COR|1|6|sicut testimonium Christi confirmatum est in vobis,
1COR|1|7|ita ut nihil vobis desit in ulla donatione, exspectantibus revelationem Domini nostri Iesu Christi;
1COR|1|8|qui et confirmabit vos usque ad finem sine crimine in die Domini nostri Iesu Christi.
1COR|1|9|Fidelis Deus, per quem vocati estis in communionem Filii eius Iesu Christi Domini nostri.
1COR|1|10|Obsecro autem vos, fratres, per nomen Domini nostri Iesu Christi, ut idipsum dicatis omnes, et non sint in vobis schismata, sitis autem perfecti in eodem sensu et in eadem sententia.
1COR|1|11|Significatum est enim mihi de vobis, fratres mei, ab his, qui sunt Chloes, quia contentiones inter vos sunt.
1COR|1|12|Hoc autem dico, quod unusquisque vestrum dicit: " Ego quidem sum Pauli, " Ego autem Apollo ", " Ego vero Cephae ", " Ego autem Christi ".
1COR|1|13|Divisus est Christus? Numquid Paulus crucifixus est pro vobis, aut in nomine Pauli baptizati estis?
1COR|1|14|Gratias ago Deo quod neminem vestrum baptizavi, nisi Crispum et Gaium,
1COR|1|15|ne quis dicat quod in nomine meo baptizati sitis.
1COR|1|16|Baptizavi autem et Stephanae domum; ceterum nescio si quem alium baptizaverim.
1COR|1|17|Non enim misit me Christus baptizare, sed evangelizare; non in sapientia verbi, ut non evacuetur crux Christi.
1COR|1|18|Verbum enim crucis pereuntibus quidem stultitia est; his autem, qui salvi fiunt, id est nobis, virtus Dei est.
1COR|1|19|Scriptum est enim: Perdam sapientiam sapientiumet prudentiam prudentium reprobabo ".
1COR|1|20|Ubi sapiens? Ubi scriba? Ubi conquisitor huius saeculi? Nonne stultam fecit Deus sapientiam huius mundi?
1COR|1|21|Nam quia in Dei sapientia non cognovit mundus per sapientiam Deum, placuit Deo per stultitiam praedicationis salvos facere credentes.
1COR|1|22|Quoniam et Iudaei signa petunt, et Graeci sapientiam quaerunt,
1COR|1|23|nos autem praedicamus Christum crucifixum, Iudaeis quidem scandalum, gentibus autem stultitiam;
1COR|1|24|ipsis autem vocatis, Iudaeis atque Graecis, Christum Dei virtutem et Dei sapientiam;
1COR|1|25|quia quod stultum est Dei, sapientius est hominibus, et, quod infirmum est Dei, fortius est hominibus.
1COR|1|26|Videte enim vocationem vestram, fratres; quia non multi sapientes secundum carnem, non multi potentes, non multi nobiles;
1COR|1|27|sed, quae stulta sunt mundi, elegit Deus, ut confundat sapientes, et infirma mundi elegit Deus, ut confundat fortia,
1COR|1|28|et ignobilia mundi et contemptibilia elegit Deus, quae non sunt, ut ea, quae sunt, destrueret,
1COR|1|29|ut non glorietur omnis caro in conspectu Dei.
1COR|1|30|Ex ipso autem vos estis in Christo Iesu, qui factus est sapientia nobis a Deo et iustitia et sanctificatio et redemptio,
1COR|1|31|ut quemadmodum scriptum est: Qui gloriatur, in Domino glorietur ".
1COR|2|1|Et ego, cum venissem ad vos, fratres, veni non per sublimita tem sermonis aut sapientiae annuntians vobis mysterium Dei.
1COR|2|2|Non enim iudicavi scire me aliquid inter vos nisi Iesum Christum et hunc crucifixum.
1COR|2|3|Et ego in infirmitate et timore et tremore multo fui apud vos,
1COR|2|4|et sermo meus et praedicatio mea non in persuasibilibus sapientiae verbis sed in ostensione Spiritus et virtutis,
1COR|2|5|ut fides vestra non sit in sapientia hominum sed in virtute Dei.
1COR|2|6|Sapientiam autem loquimur inter perfectos, sapientiam vero non huius saeculi neque principum huius saeculi, qui destruuntur,
1COR|2|7|sed loquimur Dei sapientiam in mysterio, quae abscondita est, quam praedestinavit Deus ante saecula in gloriam nostram,
1COR|2|8|quam nemo principum huius saeculi cognovit; si enim cognovissent, numquam Dominum gloriae crucifixissent.
1COR|2|9|Sed sicut scriptum est: " Quod oculus non vidit, nec auris audivit, nec in cor hominis ascendit, quae praeparavit Deus his, qui diligunt illum ".
1COR|2|10|Nobis autem revelavit Deus per Spiritum; Spiritus enim omnia scrutatur, etiam profunda Dei.
1COR|2|11|Quis enim scit hominum, quae sint hominis, nisi spiritus hominis, qui in ipso est? Ita et, quae Dei sunt, nemo cognovit nisi Spiritus Dei.
1COR|2|12|Nos autem non spiritum mundi accepimus, sed Spiritum, qui ex Deo est, ut sciamus, quae a Deo donata sunt nobis;
1COR|2|13|quae et loquimur non in doctis humanae sapientiae sed in doctis Spiritus verbis, spiritalibus spiritalia comparantes.
1COR|2|14|Animalis autem homo non percipit, quae sunt Spiritus Dei, stultitia enim sunt illi, et non potest intellegere, quia spiritaliter examinantur;
1COR|2|15|spiritalis autem iudicat omnia, et ipse a nemine iudicatur.
1COR|2|16|Quis enim cognovit sensum Domini,qui instruat eum?Nos autem sensum Christi habemus.
1COR|3|1|Et ego, fratres, non potui vobis loqui quasi spiritalibus sed qua si carnalibus, tamquam parvulis in Christo.
1COR|3|2|Lac vobis potum dedi, non escam, nondum enim poteratis. Sed ne nunc quidem potestis,
1COR|3|3|adhuc enim estis carnales. Cum enim sit inter vos zelus et contentio, nonne carnales estis et secundum hominem ambulatis?
1COR|3|4|Cum enim quis dicit: " Ego quidem sum Pauli ", alius autem: " Ego Apollo, nonne homines estis?
1COR|3|5|Quid igitur est Apollo? Quid vero Paulus? Ministri, per quos credidistis, et unicuique sicut Dominus dedit.
1COR|3|6|Ego plantavi, Apollo rigavit, sed Deus incrementum dedit;
1COR|3|7|itaque neque qui plantat, est aliquid, neque qui rigat, sed qui incrementum dat, Deus.
1COR|3|8|Qui plantat autem et qui rigat unum sunt; unusquisque autem propriam mercedem accipiet secundum suum laborem.
1COR|3|9|Dei enim sumus adiutores: Dei agri cultura estis, Dei aedificatio estis.
1COR|3|10|Secundum gratiam Dei, quae data est mihi, ut sapiens architectus fundamentum posui; alius autem superaedificat. Unusquisque autem videat quomodo superaedificet;
1COR|3|11|fundamentum enim aliud nemo potest ponere praeter id, quod positum est, qui est Iesus Christus.
1COR|3|12|Si quis autem superaedificat supra fundamentum aurum, argentum, lapides pretiosos, ligna, fenum, stipulam,
1COR|3|13|uniuscuiusque opus manifestum erit; dies enim declarabit: quia in igne revelatur, et uniuscuiusque opus quale sit ignis probabit.
1COR|3|14|Si cuius opus manserit, quod superaedificavit, mercedem accipiet;
1COR|3|15|si cuius opus arserit, detrimentum patietur, ipse autem salvus erit, sic tamen quasi per ignem.
1COR|3|16|Nescitis quia templum Dei estis, et Spiritus Dei habitat in vobis?
1COR|3|17|Si quis autem templum Dei everterit, evertet illum Deus; templum enim Dei sanctum est, quod estis vos.
1COR|3|18|Nemo se seducat; si quis videtur sapiens esse inter vos in hoc saeculo, stultus fiat, ut sit sapiens.
1COR|3|19|Sapientia enim huius mundi stultitia est apud Deum. Scriptum est enim: Qui apprehendit sapientes in astutia eorum ";
1COR|3|20|et iterum: Dominus novit cogitationes sapientium,quoniam vanae sunt ".
1COR|3|21|Itaque nemo glorietur in hominibus. Omnia enim vestra sunt,
1COR|3|22|sive Paulus sive Apollo sive Cephas sive mundus sive vita sive mors sive praesentia sive futura, omnia enim vestra sunt,
1COR|3|23|vos autem Christi, Christus autem Dei.
1COR|4|1|Sic nos existimet homo ut mi nistros Christi et dispensatores mysteriorum Dei.
1COR|4|2|Hic iam quaeritur inter dispensatores, ut fidelis quis inveniatur.
1COR|4|3|Mihi autem pro minimo est, ut a vobis iudicer aut ab humano die. Sed neque meipsum iudico;
1COR|4|4|nihil enim mihi conscius sum, sed non in hoc iustificatus sum. Qui autem iudicat me, Dominus est!
1COR|4|5|Itaque nolite ante tempus quidquam iudicare, quoadusque veniat Dominus, qui et illuminabit abscondita tenebrarum et manifestabit consilia cordium; et tunc laus erit unicuique a Deo.
1COR|4|6|Haec autem, fratres, transfiguravi in me et Apollo propter vos, ut in nobis discatis illud: " Ne supra quae scripta sunt ", ne unus pro alio inflemini adversus alterum.
1COR|4|7|Quis enim te discernit? Quid autem habes, quod non accepisti? Si autem accepisti, quid gloriaris, quasi non acceperis?
1COR|4|8|Iam saturati estis, iam divites facti estis. Sine nobis regnastis; et utinam regnaretis, ut et nos vobiscum regnaremus.
1COR|4|9|Puto enim, Deus nos apostolos novissimos ostendit tamquam morti destinatos, quia spectaculum facti sumus mundo et angelis et hominibus.
1COR|4|10|Nos stulti propter Christum, vos autem prudentes in Christo; nos infirmi, vos autem fortes; vos gloriosi, nos autem ignobiles.
1COR|4|11|Usque in hanc horam et esurimus et sitimus et nudi sumus et colaphis caedimur et instabiles sumus
1COR|4|12|et laboramus operantes manibus nostris; maledicti benedicimus, persecutionem passi sustinemus,
1COR|4|13|blasphemati obsecramus; tamquam purgamenta mundi facti sumus, omnium peripsema, usque adhuc.
1COR|4|14|Non ut confundam vos, haec scribo, sed ut quasi filios meos carissimos moneam;
1COR|4|15|nam si decem milia paedagogorum habeatis in Christo, sed non multos patres, nam in Christo Iesu per evangelium ego vos genui.
1COR|4|16|Rogo ergo vos: imitatorcs mei estote!
1COR|4|17|Ideo misi ad vos Timotheum, qui est filius meus carissimus et fidelis in Domino, qui vos commonefaciat vias meas, quae sunt in Christo, sicut ubique in omni ecclesia doceo.
1COR|4|18|Tamquam non venturus sim ad vos, sic inflati sunt quidam;
1COR|4|19|veniam autem cito ad vos, si Dominus voluerit, et cognoscam non sermonem eorum, qui inflati sunt, sed virtutem;
1COR|4|20|non enim in sermone est regnum Dei sed in virtute.
1COR|4|21|Quid vultis? In virga veniam ad vos an in caritate et spiritu mansuetudinis?
1COR|5|1|Omnino auditur inter vos for nicatio, et talis fornicatio qualis nec inter gentes, ita ut uxorem patris aliquis habeat.
1COR|5|2|Et vos inflati estis et non magis luctum habuistis, ut tollatur de medio vestrum, qui hoc opus fecit?
1COR|5|3|Ego quidem absens corpore, praesens autem spiritu, iam iudicavi ut praesens eum, qui sic operatus est,
1COR|5|4|in nomine Domini nostri Iesu, congregatis vobis et meo spiritu cum virtute Domini nostri Iesu,
1COR|5|5|tradere huiusmodi Satanae in interitum carnis, ut spiritus salvus sit in die Domini.
1COR|5|6|Non bona gloriatio vestra. Nescitis quia modicum fermentum totam massam corrumpit?
1COR|5|7|Expurgate vetus fermentum, ut sitis nova consparsio, sicut estis azymi. Etenim Pascha nostrum immolatus est Christus!
1COR|5|8|Itaque festa celebremus, non in fermento veteri neque in fermento malitiae et nequitiae, sed in azymis sinceritatis et veritatis.
1COR|5|9|Scripsi vobis in epistula: Ne commisceamini fornicariis.
1COR|5|10|Non utique fornicariis huius mundi aut avaris aut rapacibus aut idolis servientibus, alioquin debueratis de hoc mundo exisse!
1COR|5|11|Nunc autem scripsi vobis non commisceri, si is, qui frater nominatur, est fornicator aut avarus aut idolis serviens aut maledicus aut ebriosus aut rapax; cum eiusmodi nec cibum sumere.
1COR|5|12|Quid enim mihi de his, qui foris sunt, iudicare? Nonne de his, qui intus sunt, vos iudicatis?
1COR|5|13|Nam eos, qui foris sunt, Deus iudicabit. Auferte malum ex vobis ipsis!
1COR|6|1|Audet aliquis vestrum habens negotium adversus alterum iu dicari apud iniquos et non apud sanctos?
1COR|6|2|An nescitis quoniam sancti de mundo iudicabunt? Et si in vobis iudicabitur mundus, indigni estis minimis iudiciis?
1COR|6|3|Nescitis quoniam angelos iudicabimus, quanto magis saecularia?
1COR|6|4|Saecularia igitur iudicia si habueritis, contemptibiles, qui sunt in ecclesia, illos constituite ad iudicandum?
1COR|6|5|Ad verecundiam vestram dico! Sic non est inter vos sapiens quisquam, qui possit iudicare inter fratrem suum?
1COR|6|6|Sed frater cum fratre iudicio contendit, et hoc apud infideles?
1COR|6|7|Iam quidem omnino defectio est vobis, quod iudicia habetis inter vosmetipsos! Quare non magis iniuriam accipitis, quare non magis fraudem patimini?
1COR|6|8|Sed vos iniuriam facitis et fraudatis, et hoc fratribus!
1COR|6|9|An nescitis quia iniqui regnum Dei non possidebunt? Nolite errare: neque fornicarii neque idolis servientes neque adulteri neque molles neque masculorum concubitores
1COR|6|10|neque fures neque avari, non ebriosi, non maledici, non rapaces regnum Dei possidebunt.
1COR|6|11|Et haec quidam fuistis. Sed abluti estis, sed sanctificati estis, sed iustificati estis in nomine Domini Iesu Christi et in Spiritu Dei nostri!
1COR|6|12|" Omnia mihi licent! ". Sed non omnia expediunt. " Omnia mihi licent!. Sed ego sub nullius redigar potestate.
1COR|6|13|" Esca ventri, et venter escis! ". Deus autem et hunc et has destruet. Corpus autem non fornicationi sed Domino, et Dominus corpori;
1COR|6|14|Deus vero et Dominum suscitavit et nos suscitabit per virtutem suam.
1COR|6|15|Nescitis quoniam corpora vestra membra Christi sunt? Tollens ergo membra Christi faciam membra meretricis? Absit!
1COR|6|16|An nescitis quoniam, qui adhaeret meretrici, unum corpus est? " Erunt enim, inquit, duo in carne una ".
1COR|6|17|Qui autem adhaeret Domino, unus Spiritus est.
1COR|6|18|Fugite fornicationem! Omne peccatum, quodcumque fecerit homo, extra corpus est; qui autem fornicatur, in corpus suum peccat.
1COR|6|19|An nescitis quoniam corpus vestrum templum est Spiritus Sancti, qui in vobis est, quem habetis a Deo, et non estis vestri?
1COR|6|20|Empti enim estis pretio! Glorificate ergo Deum in corpore vestro.
1COR|7|1|De quibus autem scripsistis, bo num est homini mulierem non non tangere;
1COR|7|2|propter fornicationes autem unusquisque suam uxorem habeat, et unaquaeque suum virum habeat.
1COR|7|3|Uxori vir debitum reddat; similiter autem et uxor viro.
1COR|7|4|Mulier sui corporis potestatem non habet sed vir; similiter autem et vir sui corporis potestatem non habet sed mulier.
1COR|7|5|Nolite fraudare invicem, nisi forte ex consensu ad tempus, ut vacetis orationi et iterum sitis in idipsum, ne tentet vos Satanas propter incontinentiam vestram.
1COR|7|6|Hoc autem dico secundum indulgentiam, non secundum imperium.
1COR|7|7|Volo autem omnes homines esse sicut meipsum; sed unusquisque proprium habet donum ex Deo: alius quidem sic, alius vero sic.
1COR|7|8|Dico autem innuptis et viduis: Bonum est illis si sic maneant, sicut et ego;
1COR|7|9|quod si non se continent, nubant. Melius est enim nubere quam uri.
1COR|7|10|His autem, qui matrimonio iuncti sunt, praecipio, non ego sed Dominus, uxorem a viro non discedere
1COR|7|11|- quod si discesserit, maneat innupta aut viro suo reconcilietur - et virum uxorem non dimittere.
1COR|7|12|Ceteris autem ego dico, non Dominus: Si quis frater uxorem habet infidelem, et haec consentit habitare cum illo, non dimittat illam;
1COR|7|13|et si qua mulier habet virum infidelem, et hic consentit habitare cum illa, non dimittat virum.
1COR|7|14|Sanctificatus est enim vir infidelis in muliere, et sanctificata est mulier infidelis in fratre. Alioquin filii vestri immundi essent; nunc autem sancti sunt.
1COR|7|15|Quod si infidelis discedit, discedat. Non est enim servituti subiectus frater aut soror in eiusmodi; in pace autem vocavit nos Deus.
1COR|7|16|Quid enim scis, mulier, si virum salvum facies? Aut quid scis, vir, si mulierem salvam facies?
1COR|7|17|Nisi unicuique, sicut divisit Dominus, unumquemque, sicut vocavit Deus, ita ambulet; et sic in omnibus ecclesiis doceo.
1COR|7|18|Circumcisus aliquis vocatus est? Non adducat praeputium! In praeputio aliquis vocatus est? Non circumcidatur!
1COR|7|19|Circumcisio nihil est, et praeputium nihil est, sed observatio mandatorum Dei.
1COR|7|20|Unusquisque, in qua vocatione vocatus est, in ea permaneat.
1COR|7|21|Servus vocatus es? Non sit tibi curae; sed et si potes liber fieri, magis utere!
1COR|7|22|Qui enim in Domino vocatus est servus, libertus est Domini; similiter, qui liber vocatus est, servus est Christi!
1COR|7|23|Pretio empti estis! Nolite fieri servi hominum.
1COR|7|24|Unusquisque, in quo vocatus est, fratres, in hoc maneat apud Deum.
1COR|7|25|De virginibus autem praeceptum Domini non habeo; consilium autem do, tamquam misericordiam consecutus a Domino, ut sim fidelis.
1COR|7|26|Existimo ergo hoc bonum esse propter instantem necessitatem, quoniam bonum est homini sic esse.
1COR|7|27|Alligatus es uxori? Noli quaerere solutionem. Solutus es ab uxore? Noli quaerere uxorem.
1COR|7|28|Si autem acceperis uxorem, non peccasti; et si nupserit virgo, non peccavit. Tribulationem tamen carnis habebunt huiusmodi, ego autem vobis parco.
1COR|7|29|Hoc itaque dico, fratres, tempus breviatum est; reliquum est, ut et qui habent uxores, tamquam non habentes sint,
1COR|7|30|et qui flent, tamquam non flentes, et qui gaudent, tamquam non gaudentes, et qui emunt, tamquam non possidentes,
1COR|7|31|et qui utuntur hoc mundo, tamquam non abutentes; praeterit enim figura huius mundi.
1COR|7|32|Volo autem vos sine sollicitudine esse. Qui sine uxore est, sollicitus est, quae Domini sunt, quomodo placeat Domino;
1COR|7|33|qui autem cum uxore est, sollicitus est, quae sunt mundi, quomodo placeat uxori,
1COR|7|34|et divisus est. Et mulier innupta et virgo cogitat, quae Domini sunt, ut sit sancta et corpore et spiritu; quae autem nupta est, cogitat, quae sunt mundi, quomodo placeat viro.
1COR|7|35|Porro hoc ad utilitatem vestram dico, non ut laqueum vobis iniciam, sed ad id quod honestum est, et ut assidue cum Domino sitis sine distractione.
1COR|7|36|Si quis autem turpem se videri existimat super virgine sua, quod sit superadulta, et ita oportet fieri, quod vult, faciat; non peccat: nubant.
1COR|7|37|Qui autem statuit in corde suo firmus, non habens necessitatem, potestatem autem habet suae voluntatis, et hoc iudicavit in corde suo servare virginem suam, bene faciet;
1COR|7|38|igitur et, qui matrimonio iungit virginem suam, bene facit; et, qui non iungit, melius faciet.
1COR|7|39|Mulier alligata est, quanto tempore vir eius vivit; quod si dormierit vir eius, libera est, cui vult nubere, tantum in Domino.
1COR|7|40|Beatior autem erit, si sic permanserit secundum meum consilium; puto autem quod et ego Spiritum Dei habeo.
1COR|8|1|De idolothytis autem, scimus quia omnes scientiam habemus. Scientia inflat, caritas vero aedificat.
1COR|8|2|Si quis se existimat scire aliquid, nondum cognovit, quemadmodum oporteat eum scire;
1COR|8|3|si quis autem diligit Deum, hic cognitus est ab eo.
1COR|8|4|De esu igitur idolothytorum, scimus quia nullum idolum est in mundo, et quod nullus deus nisi Unus.
1COR|8|5|Nam et si sunt, qui dicantur dii sive in caelo sive in terra, si quidem sunt dii multi et domini multi,
1COR|8|6|nobis tamen unus Deus Pater, ex quo omnia et nos in illum, et unus Dominus Iesus Christus, per quem omnia et nos per ipsum.
1COR|8|7|Sed non in omnibus est scientia; quidam autem consuetudine usque nunc idoli quasi idolothytum manducant, et conscientia ipsorum, cum sit infirma, polluitur.
1COR|8|8|Esca autem nos non commendat Deo; neque si non manducaverimus, deficiemus, neque si manducaverimus, abundabimus.
1COR|8|9|Videte autem, ne forte haec licentia vestra offendiculum fiat infirmis.
1COR|8|10|Si enim quis viderit eum, qui habet scientiam, in idolio recumbentem, nonne conscientia eius, cum sit infirma, aedificabitur ad manducandum idolothyta?
1COR|8|11|Peribit enim infirmus in tua scientia, frater, propter quem Christus mortuus est!
1COR|8|12|Sic autem peccantes in fratres et percutientes conscientiam eorum infirmam, in Christum peccatis.
1COR|8|13|Quapropter si esca scandalizat fratrem meum, non manducabo carnem in aeternum, ne fratrem meum scandalizem.
1COR|9|1|Non sum liber? Non sum apo stolus? Nonne Iesum Dominum nostrum vidi? Non opus meum vos estis in Domino?
1COR|9|2|Si aliis non sum apostolus, sed tamen vobis sum; nam signaculum apostolatus mei vos estis in Domino.
1COR|9|3|Mea defensio apud eos, qui me interrogant, haec est.
1COR|9|4|Numquid non habemus potestatem manducandi et bibendi?
1COR|9|5|Numquid non habemus potestatem sororem mulierem circumducendi, sicut et ceteri apostoli et fratres Domini et Cephas?
1COR|9|6|Aut solus ego et Barnabas non habemus potestatem non operandi?
1COR|9|7|Quis militat suis stipendiis umquam? Quis plantat vineam et fructum eius non edit? Aut quis pascit gregem et de lacte gregis non manducat?
1COR|9|8|Numquid secundum hominem haec dico? An et lex haec non dicit?
1COR|9|9|Scriptum est enim in Lege Moysis: " Non alligabis os bovi trituranti ". Numquid de bobus cura est Deo?
1COR|9|10|An propter nos utique dicit? Nam propter nos scripta sunt, quoniam debet in spe, qui arat, arare; et, qui triturat, in spe fructus percipiendi.
1COR|9|11|Si nos vobis spiritalia seminavimus, magnum est, si nos carnalia vestra metamus?
1COR|9|12|Si alii potestatis vestrae participes sunt, non potius nos? Sed non usi sumus hac potestate, sed omnia sustinemus, ne quod offendiculum demus evangelio Christi.
1COR|9|13|Nescitis quoniam, qui sacra operantur, quae de sacrario sunt, edunt; qui altari deserviunt, cum altari participantur?
1COR|9|14|Ita et Dominus ordinavit his, qui evangelium annuntiant, de evangelio vivere.
1COR|9|15|Ego autem nullo horum usus sum. Non scripsi autem haec, ut ita fiant in me; bonum est enim mihi magis mori quam ut gloriam meam quis evacuet.
1COR|9|16|Nam si evangelizavero, non est mihi gloria; necessitas enim mihi incumbit. Vae enim mihi est, si non evangelizavero!
1COR|9|17|Si enim volens hoc ago, mercedem habeo; si autem invitus, dispensatio mihi credita est.
1COR|9|18|Quae est ergo merces mea? Ut evangelium praedicans sine sumptu ponam evangelium, ut non abutar potestate mea in evangelio.
1COR|9|19|Nam cum liber essem ex omnibus, omnium me servum feci, ut plures lucri facerem.
1COR|9|20|Et factus sum Iudaeis tamquam Iudaeus, ut Iudaeos lucrarer; his, qui sub lege sunt, quasi sub lege essem, cum ipse non essem sub lege, ut eos, qui sub lege erant, lucri facerem;
1COR|9|21|his, qui sine lege erant, tamquam sine lege essem, cum sine lege Dei non essem, sed in lege essem Christi, ut lucri facerem eos, qui sine lege erant;
1COR|9|22|factus sum infirmis infirmus, ut infirmos lucri facerem; omnibus omnia factus sum, ut aliquos utique facerem salvos.
1COR|9|23|Omnia autem facio propter evangelium, ut comparticeps eius efficiar.
1COR|9|24|Nescitis quod hi, qui in stadio currunt, omnes quidem currunt, sed unus accipit bravium? Sic currite, ut comprehendatis.
1COR|9|25|Omnis autem, qui in agone contendit, ab omnibus se abstinet; et illi quidem, ut corruptibilem coronam accipiant, nos autem incorruptam.
1COR|9|26|Ego igitur sic curro non quasi in incertum, sic pugno non quasi aerem verberans;
1COR|9|27|sed castigo corpus meum et in servitutem redigo, ne forte, cum aliis praedicaverim, ipse reprobus efficiar.
1COR|10|1|Nolo enim vos ignorare, fra tres, quoniam patres nostri omnes sub nube fuerunt et omnes mare transierunt
1COR|10|2|et omnes in Moyse baptizati sunt in nube et in mari
1COR|10|3|et omnes eandem escam spiritalem manducaverunt
1COR|10|4|et omnes eundem potum spiritalem biberunt; bibebant autem de spiritali, consequente eos, petra; petra autem erat Christus.
1COR|10|5|Sed non in pluribus eorum complacuit sibi Deus, nam prostrati sunt in deserto.
1COR|10|6|Haec autem figurae fuerunt nostrae, ut non simus concupiscentes malorum, sicut et illi concupierunt.
1COR|10|7|Neque idolorum cultores efficiamini, sicut quidam ex ipsis; quemadmodum scriptum est: " Sedit populus manducare et bibere, et surrexerunt ludere.
1COR|10|8|Neque fornicemur, sicut quidam ex ipsis fornicati sunt, et ceciderunt una die viginti tria milia.
1COR|10|9|Neque tentemus Christum, sicut quidam eorum tentaverunt et a serpentibus perierunt.
1COR|10|10|Neque murmuraveritis, sicut quidam eorum murmuraverunt et perierunt ab exterminatore.
1COR|10|11|Haec autem in figura contingebant illis; scripta sunt autem ad correptionem nostram, in quos fines saeculorum devenerunt.
1COR|10|12|Itaque, qui se existimat stare, videat, ne cadat.
1COR|10|13|Tentatio vos non apprehendit nisi humana; fidelis autem Deus, qui non patietur vos tentari super id quod potestis, sed faciet cum tentatione etiam proventum, ut possitis sustinere.
1COR|10|14|Propter quod, carissimi mihi, fugite ab idolorum cultura.
1COR|10|15|Ut prudentibus loquor; vos iudicate, quod dico:
1COR|10|16|Calix benedictionis, cui benedicimus, nonne communicatio sanguinis Christi est? Et panis, quem frangimus, nonne communicatio corporis Christi est?
1COR|10|17|Quoniam unus panis, unum corpus multi sumus, omnes enim de uno pane participamur.
1COR|10|18|Videte Israel secundum carnem: nonne, qui edunt hostias, communicantes sunt altari?
1COR|10|19|Quid ergo dico? Quod idolothytum sit aliquid? Aut quod idolum sit aliquid?
1COR|10|20|Sed, quae immolant, daemoniis immolant et non Deo; nolo autem vos communicantes fieri daemoniis.
1COR|10|21|Non potestis calicem Domini bibere et calicem daemoniorum; non potestis mensae Domini participes esse et mensae daemoniorum.
1COR|10|22|An aemulamur Dominum? Numquid fortiores illo sumus?
1COR|10|23|" Omnia licent! ". Sed non omnia expediunt. " Omnia licent! ". Sed non omnia aedificant.
1COR|10|24|Nemo, quod suum est, quaerat, sed quod alterius.
1COR|10|25|Omne, quod in macello venit, manducate, nihil interrogantes propter conscientiam;
1COR|10|26|Domini enim est terra, et plenitudo eius.
1COR|10|27|Si quis vocat vos infidelium, et vultis ire, omne, quod vobis apponitur, manducate, nihil interrogantes propter conscientiam.
1COR|10|28|Si quis autem vobis dixerit: " Hoc immolaticium est idolis ", nolite manducare, propter illum, qui indicavit, et propter conscientiam;
1COR|10|29|conscientiam autem dico non tuam ipsius sed alterius. Ut quid enim libertas mea iudicatur ab alia conscientia?
1COR|10|30|Si ego cum gratia participo, quid blasphemor pro eo, quod gratias ago?
1COR|10|31|Sive ergo manducatis sive bibitis sive aliud quid facitis, omnia in gloriam Dei facite.
1COR|10|32|Sine offensione estote Iudaeis et Graecis et ecclesiae Dei,
1COR|10|33|sicut et ego per omnia omnibus placeo, non quaerens, quod mihi utile est, sed quod multis, ut salvi fiant.
1COR|11|1|Imitatores mei estote, sicut et ego Christi.
1COR|11|2|Laudo autem vos quod omnia mei memores estis et, sicut tradidi vobis, traditiones meas tenetis.
1COR|11|3|Volo autem vos scire quod omnis viri caput Christus est, caput autem mulieris vir, caput vero Christi Deus.
1COR|11|4|Omnis vir orans aut prophetans velato capite deturpat caput suum;
1COR|11|5|omnis autem mulier orans aut prophetans non velato capite deturpat caput suum; unum est enim atque si decalvetur.
1COR|11|6|Nam si non velatur mulier, et tondeatur! Si vero turpe est mulieri tonderi aut decalvari, veletur.
1COR|11|7|Vir quidem non debet velare caput, quoniam imago et gloria est Dei; mulier autem gloria viri est.
1COR|11|8|Non enim vir ex muliere est, sed mulier ex viro;
1COR|11|9|etenim non est creatus vir propter mulierem, sed mulier propter virum.
1COR|11|10|Ideo debet mulier potestatem habere supra caput propter angelos.
1COR|11|11|Verumtamen neque mulier sine viro, neque vir sine muliere in Domino;
1COR|11|12|nam sicut mulier de viro, ita et vir per mulierem, omnia autem ex Deo.
1COR|11|13|In vobis ipsi iudicate: Decet mulierem non velatam orare Deum?
1COR|11|14|Nec ipsa natura docet vos quod vir quidem, si comam nutriat, ignominia est illi;
1COR|11|15|mulier vero, si comam nutriat, gloria est illi? Quoniam coma pro velamine ei data est.
1COR|11|16|Si quis autem videtur contentiosus esse, nos talem consuetudinem non habemus, neque ecclesiae Dei.
1COR|11|17|Hoc autem praecipio, non laudans quod non in melius sed in deterius convenitis.
1COR|11|18|Primum quidem convenientibus vobis in ecclesia, audio scissuras inter vos esse et ex parte credo.
1COR|11|19|Nam oportet et haereses inter vos esse, ut et, qui probati sunt, manifesti fiant in vobis.
1COR|11|20|Convenientibus ergo vobis in unum, non est dominicam cenam manducare;
1COR|11|21|unusquisque enim suam cenam praesumit in manducando, et alius quidem esurit, alius autem ebrius est.
1COR|11|22|Numquid domos non habetis ad manducandum et bibendum? Aut ecclesiam Dei contemnitis et confunditis eos, qui non habent? Quid dicam vobis? Laudabo vos? In hoc non laudo!
1COR|11|23|Ego enim accepi a Domino, quod et tradidi vobis, quoniam Dominus Iesus, in qua nocte tradebatur, accepit panem
1COR|11|24|et gratias agens fregit et dixit: " Hoc est corpus meum, quod pro vobis est; hoc facite in meam commemorationem ";
1COR|11|25|similiter et calicem, postquam cenatum est, dicens: " Hic calix novum testamentum est in meo sanguine; hoc facite, quotiescumque bibetis, in meam commemorationem ".
1COR|11|26|Quotiescumque enim manducabitis panem hunc et calicem bibetis, mortem Domini annuntiatis, donec veniat.
1COR|11|27|Itaque, quicumque manducaverit panem vel biberit calicem Domini indigne, reus erit corporis et sanguinis Domini.
1COR|11|28|Probet autem seipsum homo, et sic de pane illo edat et de calice bibat;
1COR|11|29|qui enim manducat et bibit, iudicium sibi manducat et bibit non diiudicans corpus.
1COR|11|30|Ideo inter vos multi infirmi et imbecilles et dormiunt multi.
1COR|11|31|Quod si nosmetipsos diiudicaremus, non utique iudicaremur;
1COR|11|32|dum iudicamur autem, a Domino corripimur, ut non cum hoc mundo damnemur
1COR|11|33|Itaque, fratres mei, cum convenitis ad manducandum, invicem exspectate.
1COR|11|34|Si quis esurit, domi manducet, ut non in iudicium conveniatis. Cetera autem, cum venero, disponam.
1COR|12|1|De spiritalibus autem, fra tres, nolo vos ignorare.
1COR|12|2|Scitis quoniam, cum gentes essetis, ad simulacra muta, prout ducebamini, euntes.
1COR|12|3|Ideo notum vobis facio quod nemo in Spiritu Dei loquens dicit: " Anathema Iesus! "; et nemo potest dicere: " Dominus Iesus ", nisi in Spiritu Sancto.
1COR|12|4|Divisiones vero gratiarum sunt, idem autem Spiritus;
1COR|12|5|et divisiones ministrationum sunt, idem autem Dominus;
1COR|12|6|et divisiones operationum sunt, idem vero Deus, qui operatur omnia in omnibus.
1COR|12|7|Unicuique autem datur manifestatio Spiritus ad utilitatem.
1COR|12|8|Alii quidem per Spiritum datur sermo sapientiae, alii autem sermo scientiae secundum eundem Spiritum,
1COR|12|9|alteri fides in eodem Spiritu, alii donationes sanitatum in uno Spiritu,
1COR|12|10|alii operationes virtutum, alii prophetatio, alii discretio spirituum, alii genera linguarum, alii interpretatio linguarum;
1COR|12|11|haec autem omnia operatur unus et idem Spiritus, dividens singulis prout vult.
1COR|12|12|Sicut enim corpus unum est et membra habet multa, omnia autem membra corporis, cum sint multa, unum corpus sunt, ita et Christus;
1COR|12|13|etenim in uno Spiritu omnes nos in unum corpus baptizati sumus, sive Iudaei sive Graeci sive servi sive liberi, et omnes unum Spiritum potati sumus.
1COR|12|14|Nam et corpus non est unum membrum sed multa.
1COR|12|15|Si dixerit pes: "Non sum manus, non sum de corpore ", non ideo non est de corpore;
1COR|12|16|et si dixerit auris: " Non sum oculus, non sum de corpore ", non ideo non est de corpore.
1COR|12|17|Si totum corpus oculus est, ubi auditus? Si totum auditus, ubi odoratus?
1COR|12|18|Nunc autem posuit Deus membra, unumquodque eorum in corpore, sicut voluit.
1COR|12|19|Quod si essent omnia unum membrum, ubi corpus?
1COR|12|20|Nunc autem multa quidem membra, unum autem corpus.
1COR|12|21|Non potest dicere oculus manui: " Non es mihi necessaria! "; aut iterum caput pedibus: " Non estis mihi necessarii! ".
1COR|12|22|Sed multo magis, quae videntur membra corporis infirmiora esse, necessaria sunt;
1COR|12|23|et, quae putamus ignobiliora membra esse corporis, his honorem abundantiorem circumdamus; et, quae inhonesta sunt nostra, abundantiorem honestatem habent,
1COR|12|24|honesta autem nostra nullius egent. Sed Deus temperavit corpus, ei, cui deerat, abundantiorem tribuendo honorem,
1COR|12|25|ut non sit schisma in corpore, sed idipsum pro invicem sollicita sint membra.
1COR|12|26|Et sive patitur unum membrum, compatiuntur omnia membra; sive glorificatur unum membrum, congaudent omnia membra.
1COR|12|27|Vos autem estis corpus Christi et membra ex parte.
1COR|12|28|Et quosdam quidem posuit Deus in ecclesia primum apostolos, secundo prophetas, tertio doctores, deinde virtutes, exinde donationes curationum, opitulationes, gubernationes, genera linguarum.
1COR|12|29|Numquid omnes apostoli? Numquid omnes prophetae? Numquid omnes doctores? Numquid omnes virtutes?
1COR|12|30|Numquid omnes donationes habent curationum? Numquid omnes linguis loquuntur? Numquid omnes interpretantur?
1COR|12|31|Aemulamini autem charismata maiora. Et adhuc excellentiorem viam vobis demonstro.
1COR|13|1|Si linguis hominum loquar et angelorum, caritatem au tem non habeam, factus sum velut aes sonans aut cymbalum tinniens.
1COR|13|2|Et si habuero prophetiam et noverim mysteria omnia et omnem scientiam, et si habuero omnem fidem, ita ut montes transferam, caritatem autem non habuero, nihil sum.
1COR|13|3|Et si distribuero in cibos omnes facultates meas et si tradidero corpus meum, ut glorier, caritatem autem non habuero, nihil mihi prodest.
1COR|13|4|Caritas patiens est, benigna est caritas, non aemulatur, non agit superbe, non inflatur,
1COR|13|5|non est ambitiosa, non quaerit, quae sua sunt, non irritatur, non cogitat malum,
1COR|13|6|non gaudet super iniquitatem, congaudet autem veritati;
1COR|13|7|omnia suffert, omnia credit, omnia sperat, omnia sustinet.
1COR|13|8|Caritas numquam excidit. Sive prophetiae, evacuabuntur; sive linguae, cessabunt; sive scientia, destruetur.
1COR|13|9|Ex parte enim cognoscimus et ex parte prophetamus;
1COR|13|10|cum autem venerit, quod perfectum est, evacuabitur, quod ex parte est.
1COR|13|11|Cum essem parvulus, loquebar ut parvulus, sapiebam ut parvulus, cogitabam ut parvulus; quando factus sum vir, evacuavi, quae erant parvuli.
1COR|13|12|Videmus enim nunc per speculum in aenigmate, tunc autem facie ad faciem; nunc cognosco ex parte, tunc autem cognoscam, sicut et cognitus sum.
1COR|13|13|Nunc autem manet fides, spes, caritas, tria haec; maior autem ex his est caritas.
1COR|14|1|Sectamini caritatem, aemu lamini spiritalia, magis au tem, ut prophetetis.
1COR|14|2|Qui enim loquitur lingua, non hominibus loquitur sed Deo; nemo enim audit, spiritu autem loquitur mysteria.
1COR|14|3|Qui autem prophetat, hominibus loquitur aedificationem et exhortationem et consolationes.
1COR|14|4|Qui loquitur lingua, semetipsum aedificat; qui autem prophetat, ecclesiam aedificat.
1COR|14|5|Volo autem omnes vos loqui linguis, magis autem prophetare; maior autem est qui prophetat, quam qui loquitur linguis, nisi forte interpretetur, ut ecclesia aedificationem accipiat.
1COR|14|6|Nunc autem, fratres, si venero ad vos linguis loquens, quid vobis prodero, nisi vobis loquar aut in revelatione aut in scientia aut in prophetia aut in doctrina?
1COR|14|7|Tamen, quae sine anima sunt vocem dantia, sive tibia sive cithara, nisi distinctionem sonituum dederint, quomodo scietur quod tibia canitur, aut quod citharizatur?
1COR|14|8|Etenim si incertam vocem det tuba, quis parabit se ad bellum?
1COR|14|9|Ita et vos per linguam nisi manifestum sermonem dederitis, quomodo scietur id, quod dicitur? Eritis enim in aera loquentes.
1COR|14|10|Tam multa, ut puta, genera linguarum sunt in mundo, et nihil sine voce est.
1COR|14|11|Si ergo nesciero virtutem vocis, ero ei, qui loquitur, barbarus; et, qui loquitur, mihi barbarus.
1COR|14|12|Sic et vos, quoniam aemulatores estis spirituum, ad aedificationem ecclesiae quaerite, ut abundetis.
1COR|14|13|Et ideo, qui loquitur lingua, oret, ut interpretetur.
1COR|14|14|Nam si orem lingua, spiritus meus orat, mens autem mea sine fructu est.
1COR|14|15|Quid ergo est? Orabo spiritu, orabo et mente; psallam spiritu, psallam et mente.
1COR|14|16|Ceterum si benedixeris in spiritu, qui supplet locum idiotae, quomodo dicet " Amen! " super tuam benedictionem, quoniam quid dicas nescit?
1COR|14|17|Nam tu quidem bene gratias agis, sed alter non aedificatur.
1COR|14|18|Gratias ago Deo, quod omnium vestrum magis linguis loquor;
1COR|14|19|sed in ecclesia volo quinque verba sensu meo loqui, ut et alios instruam, quam decem milia verborum in lingua.
1COR|14|20|Fratres, nolite pueri effici sensibus, sed malitia parvuli estote; sensibus autem perfecti estote.
1COR|14|21|In lege scriptum est: In aliis linguis et in labiis aliorumloquar populo huic,et nec sic exaudient me ",dicit Dominus.
1COR|14|22|Itaque linguae in signum sunt non fidelibus sed infidelibus, prophetia autem non infidelibus sed fidelibus.
1COR|14|23|Si ergo conveniat universa ecclesia in unum, et omnes linguis loquantur, intrent autem idiotae aut infideles, nonne dicent quod insanitis?
1COR|14|24|Si autem omnes prophetent, intret autem quis infidelis vel idiota, convincitur ab omnibus, diiudicatur ab omnibus,
1COR|14|25|occulta cordis eius manifesta fiunt; et ita cadens in faciem adorabit Deum pronuntians: " Vere Deus in vobis est! ".
1COR|14|26|Quid ergo est, fratres? Cum convenitis, unusquisque psalmum habet, doctrinam habet, apocalypsim habet, linguam habet, interpretationem habet: omnia ad aedificationem fiant.
1COR|14|27|Sive lingua quis loquitur, secundum duos aut ut multum tres, et per partes, et unus interpretetur;
1COR|14|28|si autem non fuerit interpres, taceat in ecclesia, sibi autem loquatur et Deo.
1COR|14|29|Prophetae duo aut tres dicant, et ceteri diiudicent;
1COR|14|30|quod si alii revelatum fuerit sedenti, prior taceat.
1COR|14|31|Potestis enim omnes per singulos prophetare, ut omnes discant, et omnes exhortentur;
1COR|14|32|et spiritus prophetarum prophetis subiecti sunt;
1COR|14|33|non enim est dissensionis Deus sed pacis.Sicut in omnibus ecclesiis sanctorum,
1COR|14|34|mulieres in ecclesiis taceant, non enim permittitur eis loqui; sed subditae sint, sicut et Lex dicit.
1COR|14|35|Si quid autem volunt discere, domi viros suos interrogent; turpe est enim mulieri loqui in ecclesia.
1COR|14|36|An a vobis verbum Dei processit aut in vos solos pervenit?
1COR|14|37|Si quis videtur propheta esse aut spiritalis, cognoscat, quae scribo vobis, quia Domini est mandatum.
1COR|14|38|Si quis autem ignorat, ignorabitur.
1COR|14|39|Itaque, fratres mei, aemulamini prophetare et loqui linguis nolite prohibere;
1COR|14|40|omnia autem honeste et secundum ordinem fiant.
1COR|15|1|Notum autem vobis facio, fratres, evangelium, quod evangelizavi vobis, quod et accepistis, in quo et statis,
1COR|15|2|per quod et salvamini, qua ratione evangelizaverim vobis, si tenetis, nisi si frustra credidistis!
1COR|15|3|Tradidi enim vobis in primis, quod et accepi, quoniam Christus mortuus est pro peccatis nostris secundum Scripturas
1COR|15|4|et quia sepultus est et quia suscitatus est tertia die secundum Scripturas
1COR|15|5|et quia visus est Cephae et post haec Duodecim;
1COR|15|6|deinde visus est plus quam quingentis fratribus simul, ex quibus plures manent usque adhuc, quidam autem dormierunt;
1COR|15|7|deinde visus est Iacobo, deinde apostolis omnibus;
1COR|15|8|novissime autem omnium, tamquam abortivo, visus est et mihi.
1COR|15|9|Ego enim sum minimus apostolorum, qui non sum dignus vocari apostolus, quoniam persecutus sum ecclesiam Dei;
1COR|15|10|gratia autem Dei sum id, quod sum, et gratia eius in me vacua non fuit, sed abundantius illis omnibus laboravi; non ego autem, sed gratia Dei mecum.
1COR|15|11|Igitur sive ego sive illi, sic praedicamus, et sic credidistis.
1COR|15|12|Si autem Christus praedicatur quod suscitatus est a mortuis, quomodo quidam dicunt in vobis quoniam resurrectio mortuorum non est?
1COR|15|13|Si autem resurrectio mortuorum non est, neque Christus suscitatus est!
1COR|15|14|Si autem Christus non suscitatus est, inanis est ergo praedicatio nostra, inanis est et fides vestra;
1COR|15|15|invenimur autem et falsi testes Dei, quoniam testimonium diximus adversus Deum quod suscitaverit Christum, quem non suscitavit, si revera mortui non resurgunt.
1COR|15|16|Nam si mortui non resurgunt, neque Christus resurrexit;
1COR|15|17|quod si Christus non resurrexit, stulta est fides vestra; adhuc estis in peccatis vestris.
1COR|15|18|Ergo et, qui dormierunt in Christo, perierunt.
1COR|15|19|Si in hac vita tantum in Christo sperantes sumus, miserabiliores sumus omnibus hominibus.
1COR|15|20|Nunc autem Christus resurrexit a mortuis, primitiae dormientium.
1COR|15|21|Quoniam enim per hominem mors, et per hominem resurrectio mortuorum:
1COR|15|22|sicut enim in Adam omnes moriuntur, ita et in Christo omnes vivificabuntur.
1COR|15|23|Unusquisque autem in suo ordine: primitiae Christus; deinde hi, qui sunt Christi, in adventu eius;
1COR|15|24|deinde finis, cum tradiderit regnum Deo et Patri, cum evacuaverit omnem principatum et omnem potestatem et virtutem.
1COR|15|25|Oportet autem illum regnare, donec ponat omnes inimicos sub pedibus eius.
1COR|15|26|Novissima autem inimica destruetur mors;
1COR|15|27|omnia enim subiecit sub pedibus eius. Cum autem dicat: "Omnia subiecta sunt", sine dubio praeter eum, qui subiecit ei omnia.
1COR|15|28|Cum autem subiecta fuerint illi omnia, tunc ipse Filius subiectus erit illi, qui sibi subiecit omnia, ut sit Deus omnia in omnibus.
1COR|15|29|Alioquin quid facient, qui baptizantur pro mortuis? Si omnino mortui non resurgunt, ut quid et baptizantur pro illis?
1COR|15|30|Ut quid et nos periclitamur omni hora?
1COR|15|31|Cotidie morior, utique per vestram gloriationem, fratres, quam habeo in Christo Iesu Domino nostro!
1COR|15|32|Si secundum hominem ad bestias pugnavi Ephesi, quid mihi prodest? Si mortui non resurgunt, manducemus et bibamus, cras enim moriemur.
1COR|15|33|Noli te seduci: " Corrumpunt mores bonos colloquia mala ".
1COR|15|34|Evigilate iuste et nolite peccare! Ignorantiam enim Dei quidam ha bent; ad reverentiam vobis loquor.
1COR|15|35|Sed dicet aliquis: " Quomodo resurgunt mortui? Quali autem corpore veniunt? ".
1COR|15|36|Insipiens! Tu, quod seminas, non vivificatur, nisi prius moriatur;
1COR|15|37|et, quod seminas, non corpus, quod futurum est, seminas sed nudum granum, ut puta tritici aut alicuius ceterorum.
1COR|15|38|Deus autem dat illi corpus sicut voluit, et unicuique seminum proprium corpus.
1COR|15|39|Non omnis caro eadem caro, sed alia hominum, alia caro pecorum, alia caro volucrum, alia autem piscium.
1COR|15|40|Et corpora caelestia et corpora terrestria, sed alia quidem caelestium gloria, alia autem terrestrium.
1COR|15|41|Alia claritas solis, alia claritas lunae et alia claritas stellarum; stella enim a stella differt in claritate.
1COR|15|42|Sic et resurrectio mortuorum: seminatur in corruptione, resurgit in incorruptione;
1COR|15|43|seminatur in ignobilitate, resurgit in gloria; seminatur in infirmitate, resurgit in virtute;
1COR|15|44|seminatur corpus animale, resurgit corpus spiritale.Si est corpus animale, est et spiritale.
1COR|15|45|Sic et scriptum est: " Factus est primus homo Adam in animam viventem; novissimus Adam in Spiritum vivificantem.
1COR|15|46|Sed non prius, quod spiritale est, sed quod animale est; deinde quod spiritale.
1COR|15|47|Primus homo de terra terrenus, secundus homo de caelo.
1COR|15|48|Qualis terrenus, tales et terreni, et qualis caelestis, tales et caelestes;
1COR|15|49|et sicut portavimus imaginem terreni, portabimus et imaginem caelestis.
1COR|15|50|Hoc autem dico, fratres, quoniam caro et sanguis regnum Dei possidere non possunt, neque corruptio incorruptelam possidebit.
1COR|15|51|Ecce mysterium vobis dico: Non omnes quidem dormiemus, sed omnes immutabimur,
1COR|15|52|in momento, in ictu oculi, in novissima tuba; canet enim, et mortui suscitabuntur incorrupti, et nos immutabimur.
1COR|15|53|Oportet enim corruptibile hoc induere incorruptelam, et mortale induere immortalitatem.
1COR|15|54|Cum autem corruptibile hoc induerit incorruptelam, et mortale hoc induerit immortalitatem, tunc fiet sermo, qui scriptus est: " Absorpta est mors in victoria.
1COR|15|55|Ubi est, mors, victoria tua?Ubi est, mors, stimulus tuus? ".
1COR|15|56|Stimulus autem mortis peccatum est, virtus vero peccati lex.
1COR|15|57|Deo autem gratias, qui dedit nobis victoriam per Dominum nostrum Iesum Christum.
1COR|15|58|Itaque, fratres mei dilecti, stabiles estote, immobiles, abundantes in opere Domini semper, scientes quod labor vester non est inanis in Domino.
1COR|16|1|De collectis autem, quae fiunt in sanctos, sicut ordina vi ecclesiis Galatiae, ita et vos facite.
1COR|16|2|Per primam sabbati unusquisque vestrum apud se ponat recondens, quod ei beneplacuerit, ut non, cum venero, tunc collectae fiant.
1COR|16|3|Cum autem praesens fuero, quos probaveritis, per epistulas hos mittam perferre gratiam vestram in Ierusalem;
1COR|16|4|quod si dignum fuerit, ut et ego eam, mecum ibunt.
1COR|16|5|Veniam autem ad vos, cum Macedoniam pertransiero, nam Macedoniam pertransibo;
1COR|16|6|apud vos autem forsitan manebo vel etiam hiemabo, ut vos me deducatis, quocumque iero.
1COR|16|7|Nolo enim vos modo in transitu videre; spero enim me aliquantum temporis manere apud vos, si Dominus permiserit.
1COR|16|8|Permanebo autem Ephesi usque ad Pentecosten;
1COR|16|9|ostium enim mihi apertum est magnum et efficax, et adversarii multi.
1COR|16|10|Si autem venerit Timotheus, videte, ut sine timore sit apud vos, opus enim Domini operatur, sicut et ego;
1COR|16|11|ne quis ergo illum spernat. Deducite autem illum in pace, ut veniat ad me; exspecto enim illum cum fratribus.
1COR|16|12|De Apollo autem fratre, multum rogavi eum, ut veniret ad vos cum fratribus, et utique non fuit voluntas, ut nunc veniret; veniet autem, cum ei opportunum fuerit.
1COR|16|13|Vigilate, state in fide, viriliter agite, confortamini;
1COR|16|14|omnia vestra in caritate fiant.
1COR|16|15|Obsecro autem vos, fratres: nostis domum Stephanae, quoniam sunt primitiae Achaiae et in ministerium sanctorum ordinaverunt seipsos;
1COR|16|16|ut et vos subditi sitis eiusmodi et omni cooperanti et laboranti.
1COR|16|17|Gaudeo autem in praesentia Stephanae et Fortunati et Achaici, quoniam id quod vobis deerat, ipsi suppleverunt;
1COR|16|18|refecerunt enim et meum spiritum et vestrum. Cognoscite ergo, qui eiusmodi sunt.
1COR|16|19|Salutant vos ecclesiae Asiae. Salutant vos in Domino multum Aquila et Prisca cum domestica sua ecclesia.
1COR|16|20|Salutant vos fratres omnes. Salutate invicem in osculo sancto.
1COR|16|21|Salutatio mea manu Pauli.
1COR|16|22|Si quis non amat Dominum, sit anathema. Marana tha!
1COR|16|23|Gratia Domini Iesu vobiscum.
1COR|16|24|Caritas mea cum omnibus vobis in Christo Iesu.
2COR|1|1|Paulus, apostolus Christi Iesu per voluntatem Dei, et Timo theus frater ecclesiae Dei, quae est Corinthi, cum sanctis omnibus, qui sunt in universa Achaia:
2COR|1|2|gratia vobis et pax a Deo Patre nostro et Domino Iesu Christo.
2COR|1|3|Benedictus Deus et Pater Domini nostri Iesu Christi, Pater misericordiarum et Deus totius consolationis,
2COR|1|4|qui consolatur nos in omni tribulatione nostra, ut possimus et ipsi consolari eos, qui in omni pressura sunt, per exhortationem, qua exhortamur et ipsi a Deo;
2COR|1|5|quoniam, sicut abundant passiones Christi in nobis, ita per Christum abundat et consolatio nostra.
2COR|1|6|Sive autem tribulamur, pro vestra exhortatione et salute; sive exhortamur, pro vestra exhortatione, quae operatur in tolerantia earundem passionum, quas et nos patimur.
2COR|1|7|Et spes nostra firma pro vobis, scientes quoniam, sicut socii passionum estis, sic eritis et consolationis.
2COR|1|8|Non enim volumus ignorare vos, fratres, de tribulatione nostra, quae facta est in Asia, quoniam supra modum gravati sumus supra virtutem, ita ut taederet nos etiam vivere;
2COR|1|9|sed ipsi in nobis ipsis responsum mortis habuimus, ut non simus fidentes in nobis sed in Deo, qui suscitat mortuos:
2COR|1|10|qui de tanta morte eripuit nos et eruet, in quem speramus, et adhuc eripiet;
2COR|1|11|adiuvantibus et vobis in oratione pro nobis, ut propter eam, quae ex multis personis in nos est, donationem, per multos gratiae agantur pro nobis.
2COR|1|12|Nam gloria nostra haec est, testimonium conscientiae nostrae, quod in simplicitate et sinceritate Dei et non in sapientia carnali, sed in gratia Dei conversati sumus in mundo, abundantius autem ad vos.
2COR|1|13|Non enim alia scribimus vobis quam quae legitis aut etiam cognoscitis; spero autem quod usque in finem cognoscetis,
2COR|1|14|sicut et cognovistis nos ex parte, quia gloria vestra sumus, sicut et vos nostra in die Domini nostri Iesu.
2COR|1|15|Et hac confidentia volui prius venire ad vos, ut secundam gratiam haberetis,
2COR|1|16|et per vos transire in Macedoniam et iterum a Macedonia venire ad vos et a vobis deduci in Iudaeam.
2COR|1|17|Cum hoc ergo voluissem, numquid levitate usus sum? Aut, quae cogito, secundum carnem cogito, ut sit apud me " Est, est " et " Non, non "?
2COR|1|18|Fidelis autem Deus, quia sermo noster, qui fit apud vos, non est " Est et " Non "!
2COR|1|19|Dei enim Filius Iesus Christus, qui in vobis per nos praedicatus est, per me et Silvanum et Timotheum, non fuit " Est " et " Non ", sed " Est " in illo fuit.
2COR|1|20|Quotquot enim promissiones Dei sunt, in illo " Est "; ideo et per ipsum Amen " Deo ad gloriam per nos.
2COR|1|21|Qui autem confirmat nos vobiscum in Christum et qui unxit nos, Deus,
2COR|1|22|et qui signavit nos et dedit arrabonem Spiritus in cordibus nostris.
2COR|1|23|Ego autem testem Deum invoco in animam meam, quod parcens vobis non veni ultra Corinthum.
2COR|1|24|Non quia dominamur fidei vestrae, sed adiutores sumus gaudii vestri, nam fide stetistis.
2COR|2|1|Statui autem hoc ipse apud me, ne iterum in tristitia venirem ad vos;
2COR|2|2|si enim ego contristo vos, et quis est qui me laetificet, nisi qui contristatur ex me?
2COR|2|3|Et hoc ipsum scripsi, ut non, cum venero, tristitiam habeam de quibus oportebat me gaudere, confidens in omnibus vobis, quia meum gaudium omnium vestrum est.
2COR|2|4|Nam ex multa tribulatione et angustia cordis scripsi vobis per multas lacrimas, non ut contristemini, sed ut sciatis quam carita tem habeo abundantius in vos.
2COR|2|5|Si quis autem contristavit, non me contristavit, sed ex parte, ut non onerem, omnes vos.
2COR|2|6|Sufficit illi, qui eiusmodi est, obiurgatio haec, quae fit a pluribus,
2COR|2|7|ita ut e contra magis donetis et consolemini, ne forte abundantiore tristitia absorbeatur, qui eiusmodi est.
2COR|2|8|Propter quod obsecro vos, ut confirmetis in illum caritatem;
2COR|2|9|ideo enim et scripsi, ut cognoscam probationem vestram, an in omnibus oboedientes sitis.
2COR|2|10|Cui autem aliquid donatis, et ego; nam et ego, quod donavi, si quid donavi, propter vos in persona Christi,
2COR|2|11|ut non circumveniamur a Satana; non enim ignoramus cogitationes eius.
2COR|2|12|Cum venissem autem Troadem ob evangelium Christi, et ostium mihi apertum esset in Domino,
2COR|2|13|non habui requiem spiritui meo, eo quod non invenerim Titum fratrem meum, sed valefaciens eis profectus sum in Macedoniam.
2COR|2|14|Deo autem gratias, qui semper triumphat nos in Christo et odorem notitiae suae manifestat per nos in omni loco.
2COR|2|15|Quia Christi bonus odor sumus Deo in his, qui salvi fiunt, et in his, qui pereunt:
2COR|2|16|aliis quidem odor ex morte in mortem, aliis autem odor ex vita in vitam. Et ad haec quis idoneus?
2COR|2|17|Non enim sumus sicut plurimi adulterantes verbum Dei, sed sicut ex sinceritate, sed sicut ex Deo coram Deo in Christo loquimur.
2COR|3|1|Incipimus iterum nosmetipsos commendare? Aut numquid egemus, sicut quidam, commendaticiis epistulis ad vos aut ex vobis?
2COR|3|2|Epistula nostra vos estis, scripta in cordibus nostris, quae scitur et legitur ab omnibus hominibus;
2COR|3|3|manifestati quoniam epistula estis Christi ministrata a nobis, scripta non atramento sed Spiritu Dei vivi, non in tabulis lapideis sed in tabulis cordis carnalibus.
2COR|3|4|Fiduciam autem talem habemus per Christum ad Deum.
2COR|3|5|Non quod sufficientes simus cogitare aliquid a nobis quasi ex nobis, sed sufficientia nostra ex Deo est,
2COR|3|6|qui et idoneos nos fecit ministros Novi Testamenti, non litterae sed Spiritus: littera enim occidit, Spiritus autem vivificat.
2COR|3|7|Quod si ministratio mortis, litteris deformata in lapidibus, fuit in gloria, ita ut non possent intendere filii Israel in faciem Moysis propter gloriam vultus eius, quae evacuatur,
2COR|3|8|quomodo non magis ministratio Spiritus erit in gloria?
2COR|3|9|Nam si ministerium damnationis gloria est, multo magis abundat ministerium iustitiae in gloria.
2COR|3|10|Nam nec glorificatum est, quod claruit in hac parte, propter excellentem gloriam;
2COR|3|11|si enim, quod evacuatur, per gloriam est, multo magis, quod manet, in gloria est.
2COR|3|12|Habentes igitur talem spem multa fiducia utimur,
2COR|3|13|et non sicut Moyses: ponebat velamen super faciem suam, ut non intenderent filii Israel in finem illius quod evacuatur.
2COR|3|14|Sed obtusi sunt sensus eorum. Usque in hodiernum enim diem idipsum velamen in lectione Veteris Testamenti manet non revelatum, quoniam in Christo evacuatur;
2COR|3|15|sed usque in hodiernum diem, cum legitur Moyses, velamen est positum super cor eorum.
2COR|3|16|Quando autem conversus fuerit ad Dominum, aufertur velamen.
2COR|3|17|Dominus autem Spiritus est; ubi autem Spiritus Domini, ibi libertas.
2COR|3|18|Nos vero omnes revelata facie gloriam Domini speculantes, in eandem imaginem transformamur a claritate in clarita tem tamquam a Domini Spiritu.
2COR|4|1|Ideo habentes hanc ministra tionem, iuxta quod misericor diam consecuti sumus, non deficimus,
2COR|4|2|sed abdicavimus occulta dedecoris non ambulantes in astutia neque adulterantes verbum Dei, sed in manifestatione veritatis commendantes nosmetipsos ad omnem conscientiam hominum coram Deo.
2COR|4|3|Quod si etiam velatum est evangelium nostrum, in his, qui pereunt, est velatum;
2COR|4|4|in quibus deus huius saeculi excaecavit mentes infidelium, ut non fulgeat illuminatio evangelii gloriae Christi, qui est imago Dei.
2COR|4|5|Non enim nosmetipsos praedicamus sed Iesum Christum Dominum; nos autem servos vestros per Iesum.
2COR|4|6|Quoniam Deus, qui dixit: " De tenebris lux splendescat ", ipse illuxit in cordibus nostris ad illuminationem scientiae claritatis Dei in facie Iesu Christi.
2COR|4|7|Habemus autem thesaurum istum in vasis fictilibus, ut sublimitas sit virtutis Dei et non ex nobis.
2COR|4|8|In omnibus tribulationem patimur, sed non angustiamur; aporiamur, sed non destituimur;
2COR|4|9|persecutionem patimur, sed non derelinquimur; deicimur, sed non perimus;
2COR|4|10|semper mortificationem Iesu in corpore circumferentes, ut et vita Iesu in corpore nostro manifestetur.
2COR|4|11|Semper enim nos, qui vivimus, in mortem tradimur propter Iesum, ut et vita Iesu manifestetur in carne nostra mortali.
2COR|4|12|Ergo mors in nobis operatur, vita autem in vobis.
2COR|4|13|Habentes autem eundem spiritum fidei, sicut scriptum est: " Credidi, propter quod locutus sum ", et nos credimus, propter quod et loquimur,
2COR|4|14|scientes quoniam, qui suscitavit Dominum Iesum, et nos cum Iesu suscitabit et constituet vobiscum.
2COR|4|15|Omnia enim propter vos, ut gratia abundans per multos gratiarum actionem abundare faciat in gloriam Dei.
2COR|4|16|Propter quod non deficimus, sed licet is, qui foris est, noster homo corrumpitur, tamen is, qui intus est, noster renovatur de die in diem.
2COR|4|17|Id enim, quod in praesenti est, leve tribulationis nostrae supra modum in sublimitatem aeternum gloriae pondus operatur nobis,
2COR|4|18|non contemplantibus nobis, quae videntur, sed quae non videntur; quae enim videntur, temporalia sunt, quae autem non videntur, aeterna sunt.
2COR|5|1|Scimus enim quoniam, si terre stris domus nostra huius taber naculi dissolvatur, aedificationem ex Deo habemus domum non manufactam, aeternam in caelis.
2COR|5|2|Nam et in hoc ingemiscimus, habitationem nostram, quae de caelo est, superindui cupientes,
2COR|5|3|si tamen et exspoliati, non nudi inveniamur.
2COR|5|4|Nam et, qui sumus in tabernaculo, ingemiscimus gravati, eo quod nolumus exspoliari, sed supervestiri, ut absorbeatur, quod mortale est, a vita.
2COR|5|5|Qui autem effecit nos in hoc ipsum, Deus, qui dedit nobis arrabonem Spiritus.
2COR|5|6|Audentes igitur semper et scientes quoniam, dum praesentes sumus in corpore, peregrinamur a Domino;
2COR|5|7|per fidem enim ambulamus et non per speciem.
2COR|5|8|Audemus autem et bonam voluntatem habemus magis peregrinari a corpore et praesentes esse ad Dominum.
2COR|5|9|Et ideo contendimus sive praesentes sive absentes placere illi.
2COR|5|10|Omnes enim nos manifestari oportet ante tribunal Christi, ut referat unusquisque pro eis, quae per corpus gessit, sive bonum sive malum.
2COR|5|11|Scientes ergo timorem Domini hominibus suademus, Deo autem manifesti sumus; spero autem et in conscientiis vestris manifestos nos esse.
2COR|5|12|Non iterum nos commendamus vobis, sed occasionem damus vobis gloriandi pro nobis, ut habeatis ad eos, qui in facie gloriantur et non in corde.
2COR|5|13|Sive enim mente excedimus, Deo; sive sobrii sumus, vobis.
2COR|5|14|Caritas enim Christi urget nos, aestimantes, hoc, quoniam, si unus pro omnibus mortuus est, ergo omnes mortui sunt;
2COR|5|15|et pro omnibus mortuus est, ut et, qui vivunt, iam non sibi vivant, sed ei, qui pro ipsis mortuus est et resurrexit.
2COR|5|16|Itaque nos ex hoc neminem novimus secundum carnem; et si cognovimus secundum carnem Christum, sed nunc iam non novimus.
2COR|5|17|Si quis ergo in Christo, nova creatura; vetera transierunt, ecce, facta sunt nova.
2COR|5|18|Omnia autem ex Deo, qui reconciliavit nos sibi per Christum et dedit nobis ministerium reconciliationis,
2COR|5|19|quoniam quidem Deus erat in Christo mundum reconcilians sibi, non reputans illis delicta ipsorum; et posuit in nobis verbum reconciliationis.
2COR|5|20|Pro Christo ergo legatione fungimur, tamquam Deo exhortante per nos. Obsecramus pro Christo, reconciliamini Deo.
2COR|5|21|Eum, qui non noverat peccatum, pro nobis peccatum fecit, ut nos efficeremur iustitia Dei in ipso.
2COR|6|1|Adiuvantes autem et exhor tamur, ne in vacuum gratiam Dei recipiatis
2COR|6|2|- ait enim: Tempore accepto exaudivi teet in die salutis adiuvi te ";ecce nunc tempus acceptabile, ecce nunc dies salutis -
2COR|6|3|nemini dantes ullam offensionem, ut non vituperetur ministerium,
2COR|6|4|sed in omnibus exhibentes nosmetipsos sicut Dei ministros in multa patientia, in tribulationibus, in necessitatibus, in angustiis,
2COR|6|5|in plagis, in carceribus, in seditionibus, in laboribus, in vigiliis, in ieiuniis,
2COR|6|6|in castitate, in scientia, in longanimitate, in suavitate, in Spiritu Sancto, in caritate non ficta,
2COR|6|7|in verbo veritatis, in virtute Dei; per arma iustitiae a dextris et sinistris,
2COR|6|8|per gloriam et ignobilitatem, per infamiam et bonam famam; ut seductores, et veraces;
2COR|6|9|sicut qui ignoti, et cogniti; quasi morientes, et ecce vivimus; ut castigati, et non mortificati;
2COR|6|10|quasi tristes, semper autem gaudentes; sicut egentes, multos autem locupletantes; tamquam nihil habentes, et omnia possidentes.
2COR|6|11|Os nostrum patet ad vos, o Corinthii, cor nostrum dilatatum est.
2COR|6|12|Non angustiamini in nobis, sed angustiamini in visceribus vestris;
2COR|6|13|eandem autem habentes remunerationem, tamquam filiis dico, dilatamini et vos.
2COR|6|14|Nolite iugum ducere cum infidelibus! Quae enim participatio iustitiae cum iniquitate? Aut quae societas luci ad tenebras?
2COR|6|15|Quae autem conventio Christi cum Beliar, aut quae pars fideli cum infideli?
2COR|6|16|Qui autem consensus templo Dei cum idolis? Vos enim estis templum Dei vivi; sicut dicit Deus: Inhabitabo in illis et inambulaboet ero illorum Deus, et ipsi erunt mihi populus.
2COR|6|17|Propter quod exite de medio eorumet separamini, dicit Dominus,et immundum ne tetigeritis;et ego recipiam vos
2COR|6|18|et ero vobis in Patrem,et vos eritis mihi in filios et filias,dicit Dominus omnipotens ".
2COR|7|1|Has igitur habentes promissio nes, carissimi, mundemus nos ab omni inquinamento carnis et spiritus, perficientes sanctificationem in timore Dei.
2COR|7|2|Capite nos! Neminem laesimus, neminem corrupimus, neminem circumvenimus.
2COR|7|3|Non ad condemnationem dico; praedixi enim quod in cordibus nostris estis ad commoriendum et ad convivendum.
2COR|7|4|Multa mihi fiducia est apud vos, multa mihi gloriatio pro vobis; repletus sum consolatione, superabundo gaudio in omni tribulatione nostra.
2COR|7|5|Nam et cum venissemus Macedoniam, nullam requiem habuit caro nostra, sed omnem tribulationem passi: foris pugnae, intus timores.
2COR|7|6|Sed qui consolatur humiles, consolatus est nos Deus in adventu Titi;
2COR|7|7|non solum autem in adventu eius sed etiam in solacio, quo consolatus est in vobis, referens nobis vestrum desiderium, vestrum fletum, vestram aemulationem pro me, ita ut magis gauderem.
2COR|7|8|Quoniam etsi contristavi vos in epistula, non me paenitet; etsi paeniteret - video quod epistula illa, etsi ad horam, vos contristavit -
2COR|7|9|nunc gaudeo, non quia contristati estis, sed quia contristati estis ad paenitentiam; contristati enim estis secundum Deum, ut in nullo detrimentum patiamini ex nobis.
2COR|7|10|Quae enim secundum Deum tristitia, paenitentiam in salutem stabilem operatur; saeculi autem tristitia mortem operatur.
2COR|7|11|Ecce enim hoc ipsum secundum Deum contristari: quantam in vobis operatum est sollicitudinem, sed defensionem, sed indignationem, sed timorem, sed desiderium, sed aemulationem, sed vindictam! In omnibus exhibuistis vos incontaminatos esse negotio.
2COR|7|12|Igitur etsi scripsi vobis, non propter eum, qui fecit iniuriam, nec propter eum, qui passus est, sed ad manifestandam sollicitudinem vestram, quam pro nobis habetis, ad vos coram Deo.
2COR|7|13|Ideo consolati sumus.In consolatione autem nostra abundantius magis gavisi sumus super gaudium Titi, quia refectus est spiritus eius ab omnibus vobis;
2COR|7|14|et si quid apud illum de vobis gloriatus sum, non sum confusus, sed sicut omnia vobis in veritate locuti sumus, ita et gloriatio nostra, quae fuit ad Titum, veritas facta est.
2COR|7|15|Et viscera eius abundantius in vos sunt, reminiscentis omnium vestrum oboedientiam, quomodo cum timore et tremore excepistis eum.
2COR|7|16|Gaudeo quod in omnibus confido in vobis.
2COR|8|1|Notam autem facimus vobis, fratres, gratiam Dei, quae data est in ecclesiis Macedoniae,
2COR|8|2|quod in multo experimento tribulationis abundantia gaudii ipsorum et altissima paupertas eorum abundavit in divitias simplicitatis eorum;
2COR|8|3|quia secundum virtutem, testimonium reddo, et supra virtutem voluntarii fuerunt
2COR|8|4|cum multa exhortatione obsecrantes nos gratiam et communicationem ministerii, quod fit in sanctos.
2COR|8|5|Et non sicut speravimus, sed semetipsos dederunt primum Domino, deinde nobis per voluntatem Dei,
2COR|8|6|ita ut rogaremus Titum, ut, quemadmodum coepit, ita et perficiat in vos etiam gratiam istam.
2COR|8|7|Sed sicut in omnibus abundatis, fide et sermone et scientia et omni sollicitudine et caritate ex nobis in vobis, ut et in hac gratia abundetis.
2COR|8|8|Non quasi imperans dico, sed per aliorum sollicitudinem etiam vestrae caritatis ingenitum bonum comprobans;
2COR|8|9|scitis enim gratiam Domini nostri Iesu Christi, quoniam propter vos egenus factus est, cum esset dives, ut illius inopia vos divites essetis.
2COR|8|10|Et consilium in hoc do. Hoc enim vobis utile est, qui non solum facere, sed et velle coepistis ab anno priore;
2COR|8|11|nunc vero et facto perficite, ut, quemadmodum promptus est animus velle, ita sit et perficere ex eo, quod habetis.
2COR|8|12|Si enim voluntas prompta est, secundum id quod habet, accepta est, non secundum quod non habet.
2COR|8|13|Non enim, ut aliis sit remissio, vobis autem tribulatio; sed ex aequalitate
2COR|8|14|in praesenti tempore vestra abundantia illorum inopiam suppleat, ut et illorum abundantia vestram inopiam suppleat, ut fiat aequalitas, sicut scriptum est:
2COR|8|15|" Qui multum, non abundavit; et, qui modicum, non minoravit ".
2COR|8|16|Gratias autem Deo, qui dedit eandem sollicitudinem pro vobis in corde Titi,
2COR|8|17|quoniam exhortationem quidem suscepit, sed, cum sollicitior esset, sua voluntate profectus est ad vos.
2COR|8|18|Misimus etiam cum illo fratrem, cuius laus est in evangelio per omnes ecclesias
2COR|8|19|- non solum autem, sed et ordinatus ab ecclesiis comes noster cum hac gratia, quae ministratur a nobis ad Domini gloriam et destinatam voluntatem nostram -
2COR|8|20|devitantes hoc, ne quis nos vituperet in hac plenitudine, quae ministratur a nobis;
2COR|8|21|providemus enim bona non solum coram Domino sed etiam coram hominibus.
2COR|8|22|Misimus autem cum illis et fratrem nostrum, quem probavimus in multis saepe sollicitum esse, nunc autem multo sollicitiorem, confidentia multa in vos.
2COR|8|23|Sive pro Tito, est socius meus et in vos adiutor; sive fratres nostri, apostoli ecclesiarum, gloria Christi.
2COR|8|24|Ostensionem ergo, quae est caritatis vestrae et nostrae gloriationis pro vobis, in illos ostendite in faciem ecclesiarum.
2COR|9|1|Nam de ministerio, quod fit in sanctos, superfluum est mihi scribere vobis;
2COR|9|2|scio enim promptum animum vestrum, pro quo de vobis glorior apud Macedonas, quoniam Achaia parata est ab anno praeterito, et vestra aemulatio provocavit plurimos.
2COR|9|3|Misi autem fratres, ut ne, quod gloriamur de vobis, evacuetur in hac parte, ut, quemadmodum dixi, parati sitis,
2COR|9|4|ne, cum venerint mecum Macedones et invenerint vos imparatos, erubescamus nos, ut non dicam vos, in hac substantia.
2COR|9|5|Necessarium ergo existimavi rogare fratres, ut praeveniant ad vos et praeparent repromissam benedictionem vestram, ut haec sit parata sic quasi benedictio, non quasi avaritia.
2COR|9|6|Hoc autem: qui parce seminat, parce et metet; et, qui seminat in benedictionibus, in benedictionibus et metet.
2COR|9|7|Unusquisque prout destinavit corde suo, non ex tristitia aut ex necessitate; hilarem enim datorem diligit Deus.
2COR|9|8|Potens est autem Deus omnem gratiam abundare facere in vobis, ut, in omnibus semper omnem sufficientiam habentes, abundetis in omne opus bonum,
2COR|9|9|sicut scriptum est: Dispersit, dedit pauperibus;iustitia eius manet in aeternum ".
2COR|9|10|Qui autem administrat semen seminanti, et panem ad manducandum praestabit et multiplicabit semen vestrum et augebit incrementa frugum iustitiae vestrae.
2COR|9|11|In omnibus locupletati in omnem simplicitatem, quae operatur per nos gratiarum actionem Deo
2COR|9|12|- quoniam ministerium huius officii non solum supplet ea, quae desunt sanctis, sed etiam abundat per multas gratiarum actiones Deo -
2COR|9|13|per probationem ministerii huius glorificantes Deum in oboedientia confessionis vestrae in evangelium Christi et simplicitate communionis in illos et in omnes,
2COR|9|14|et ipsorum obsecratione pro vobis, desiderantium vos propter eminentem gratiam Dei in vobis.
2COR|9|15|Gratias Deo super inenarrabili dono eius.
2COR|10|1|Ipse autem ego Paulus obse cro vos per mansuetudinem et modestiam Christi, qui in facie quidem humilis inter vos, absens autem confido in vobis;
2COR|10|2|rogo autem, ne praesens audeam per eam confidentiam, quae existimo audere in quosdam, qui arbitrantur nos tamquam secundum carnem ambulemus.
2COR|10|3|In carne enim ambulantes, non secundum carnem militamus
2COR|10|4|- nam arma militiae nostrae non carnalia sed potentia Deo ad destructionem munitionum - consilia destruentes
2COR|10|5|et omnem altitudinem extollentem se adversus scientiam Dei, et in captivitatem redigentes omnem intellectum in obsequium Christi,
2COR|10|6|et in promptu habentes ulcisci omnem inoboedientiam, cum impleta fuerit vestra oboedientia.
2COR|10|7|Quae secundum faciem sunt, videte. Si quis confidit sibi Christi se esse, hoc cogitet iterum apud se, quia sicut ipse Christi est, ita et nos.
2COR|10|8|Nam et si amplius aliquid gloriatus fuero de potestate nostra, quam dedit Dominus in aedificationem et non in destructionem vestram, non erubescam,
2COR|10|9|ut non existimer tamquam terrere vos per epistulas;
2COR|10|10|quoniam quidem " Epistulae - inquiunt - graves sunt et fortes, praesentia autem corporis infirma, et sermo contemptibilis ".
2COR|10|11|Hoc cogitet, qui eiusmodi est, quia quales sumus verbo per epistulas absentes, tales et praesentes in facto.
2COR|10|12|Non enim audemus inserere aut comparare nos quibusdam, qui seipsos commendant; sed ipsi se in semetipsis metientes et comparantes semetipsos sibi, non intellegunt.
2COR|10|13|Nos autem non ultra mensuram gloriabimur sed secundum mensuram regulae, quam impertitus est nobis Deus, mensuram pertingendi usque ad vos.
2COR|10|14|Non enim quasi non pertingentes ad vos superextendimus nosmetipsos, usque ad vos enim pervenimus in evangelio Christi;
2COR|10|15|non ultra mensuram gloriantes in alienis laboribus, spem autem habentes, crescente fide vestra, in vobis magnificari secundum regulam nostram in abundantiam,
2COR|10|16|ad evangelizandum in iis, quae ultra vos sunt, et non in aliena regula gloriari in his, quae praeparata sunt.
2COR|10|17|Qui autem gloriatur, in Domino glorietur;
2COR|10|18|non enim qui seipsum commendat, ille probatus est, sed quem Dominus commendat.
2COR|11|1|Utinam sustineretis modi cum quid insipientiae meae; sed et supportate me!
2COR|11|2|Aemulor enim vos Dei aemulatione; despondi enim vos uni viro virginem castam exhibere Christo.
2COR|11|3|Timeo autem, ne, sicut serpens Evam seduxit astutia sua, ita corrumpantur sensus vestri a simplicitate et castitate, quae est in Christum.
2COR|11|4|Nam si is qui venit, alium Christum praedicat, quem non praedicavimus, aut alium Spiritum accipitis, quem non accepistis, aut aliud evangelium, quod non recepistis, recte pateremini.
2COR|11|5|Existimo enim nihil me minus fecisse magnis apostolis;
2COR|11|6|nam etsi imperitus sermone, sed non scientia, in omni autem manifestantes in omnibus ad vos.
2COR|11|7|Aut numquid peccatum feci meipsum humilians, ut vos exaltemini, quoniam gratis evangelium Dei evangelizavi vobis?
2COR|11|8|Alias ecclesias exspoliavi accipiens stipendium ad ministerium vestrum
2COR|11|9|et, cum essem apud vos et egerem, nulli onerosus fui; nam, quod mihi deerat, suppleverunt fratres, qui venerunt a Macedonia; et in omnibus sine onere me vobis servavi et servabo.
2COR|11|10|Est veritas Christi in me, quoniam haec gloria non infringetur in me in regionibus Achaiae.
2COR|11|11|Quare? Quia non diligo vos? Deus scit!
2COR|11|12|Quod autem facio et faciam, ut amputem occasionem eorum, qui volunt occasionem, ut in quo gloriantur, inveniantur sicut et nos.
2COR|11|13|Nam eiusmodi pseudoapostoli, operarii subdoli, transfigurantes se in apostolos Christi.
2COR|11|14|Et non mirum, ipse enim Satanas transfigurat se in angelum lucis;
2COR|11|15|non est ergo magnum, si et ministri eius transfigurentur velut ministri iustitiae, quorum finis erit secundum opera ipsorum.
2COR|11|16|Iterum dico, ne quis me putet insipientem esse; alioquin velut insipientem accipite me, ut et ego modicum quid glorier.
2COR|11|17|Quod loquor, non loquor secundum Dominum, sed quasi in insipientia, in hac substantia gloriationis.
2COR|11|18|Quoniam multi gloriantur secundum carnem, et ego gloriabor.
2COR|11|19|Libenter enim suffertis insipientes, cum sitis ipsi sapientes;
2COR|11|20|sustinetis enim, si quis vos in servitutem redigit, si quis devorat, si quis accipit, si quis extollitur, si quis in faciem vos caedit.
2COR|11|21|Secundum ignobilitatem dico, quasi nos infirmi fuerimus; in quo quis audet, in insipientia dico, audeo et ego.
2COR|11|22|Hebraei sunt? Et ego. Israelitae sunt? Et ego. Semen Abrahae sunt? Et ego.
2COR|11|23|Ministri Christi sunt? Minus sapiens dico, plus ego: in laboribus plurimis, in carceribus abundantius, in plagis supra modum, in mortibus frequenter;
2COR|11|24|a Iudaeis quinquies quadragenas una minus accepi,
2COR|11|25|ter virgis caesus sum, semel lapidatus sum, ter naufragium feci, nocte et die in profundo maris fui;
2COR|11|26|in itineribus saepe, periculis fluminum, periculis latronum, periculis ex genere, periculis ex gentibus, periculis in civitate, periculis in solitudine, periculis in mari, periculis in falsis fratribus;
2COR|11|27|in labore et aerumna, in vigiliis saepe, in fame et siti, in ieiuniis frequenter, in frigore et nuditate;
2COR|11|28|praeter illa, quae extrinsecus sunt, instantia mea cotidiana, sollicitudo omnium ecclesiarum.
2COR|11|29|Quis infirmatur, et non infirmor? Quis scandalizatur, et ego non uror?
2COR|11|30|Si gloriari oportet, quae infirmitatis meae sunt, gloriabor.
2COR|11|31|Deus et Pater Domini Iesu scit, qui est benedictus in saecula, quod non mentior.
2COR|11|32|Damasci praepositus gentis Aretae regis custodiebat civitatem Damascenorum, ut me comprehenderet;
2COR|11|33|et per fenestram in sporta dimissus sum per murum et effugi manus eius.
2COR|12|1|Gloriari oportet; non expedit quidem, veniam autem ad visiones et revelationes Domini.
2COR|12|2|Scio hominem in Christo ante annos quattuordecim - sive in corpore nescio, sive extra corpus nescio, Deus scit - raptum eiusmodi usque ad tertium caelum.
2COR|12|3|Et scio huiusmodi hominem - sive in corpore sive extra corpus nescio, Deus scit -
2COR|12|4|quoniam raptus est in paradisum et audivit arcana verba, quae non licet homini loqui.
2COR|12|5|Pro eiusmodi gloriabor; pro me autem nihil gloriabor nisi in infirmitatibus meis.
2COR|12|6|Nam, et si voluero gloriari, non ero insipiens, veritatem enim dicam; parco autem, ne quis in me existimet supra id, quod videt me aut audit ex me,
2COR|12|7|et ex magnitudine revelationum. Propter quod, ne extollar, datus est mihi stimulus carni, angelus Satanae, ut me colaphizet, ne extollar.
2COR|12|8|Propter quod ter Dominum rogavi, ut discederet a me;
2COR|12|9|et dixit mihi: " Sufficit tibi gratia mea, nam virtus in infirmitate perficitur ". Libentissime igitur potius gloriabor in infirmitatibus meis, ut inhabitet in me virtus Christi.
2COR|12|10|Propter quod placeo mihi in infirmitatibus, in contumeliis, in necessitatibus, in persecutionibus et in angustiis, pro Christo; cum enim infirmor, tunc potens sum.
2COR|12|11|Factus sum insipiens. Vos me coegistis; ego enim debui a vobis commendari. Nihil enim minus fui ab his, qui sunt supra modum apostoli, tametsi nihil sum;
2COR|12|12|signa tamen apostoli facta sunt super vos in omni patientia, signis quoque et prodigiis et virtutibus.
2COR|12|13|Quid est enim quod minus habuistis prae ceteris ecclesiis, nisi quod ego ipse non gravavi vos? Donate mihi hanc iniuriam.
2COR|12|14|Ecce tertio hoc paratus sum venire ad vos et non ero gravis vobis; non enim quaero, quae vestra sunt, sed vos; nec enim debent filii parentibus thesaurizare, sed parentes filiis.
2COR|12|15|Ego autem libentissime impendam et superimpendar ipse pro animabus vestris. Si plus vos diligo, minus diligar?
2COR|12|16|Esto quidem, ego vos non gravavi; sed cum essem astutus, dolo vos cepi.
2COR|12|17|Numquid per aliquem eorum, quos misi ad vos, circumveni vos?
2COR|12|18|Rogavi Titum et misi cum illo fratrem; numquid Titus vos circumvenit? Nonne eodem spiritu ambulavimus? Nonne iisdem vestigiis?
2COR|12|19|Olim putatis quod excusemus nos apud vos? Coram Deo in Christo loquimur; omnia autem, carissimi, propter vestram aedificationem.
2COR|12|20|Timeo enim, ne forte, cum venero, non quales volo, inveniam vos, et ego inveniar a vobis, qualem non vultis; ne forte contentiones, aemulationes, animositates, dissensiones, detractiones, susurrationes, inflationes, seditiones sint;
2COR|12|21|ne iterum, cum venero, humiliet me Deus meus apud vos, et lugeam multos ex his, qui ante peccaverunt et non egerunt paenitentiam super immunditia et fornicatione et impudicitia, quam gesserunt.
2COR|13|1|Ecce tertio hoc venio ad vos; in ore duorum vel trium testium stabit omne verbum.
2COR|13|2|Praedixi et praedico, ut praesens bis et nunc absens his, qui ante peccaverunt, et ceteris omnibus, quoniam, si venero iterum, non parcam,
2COR|13|3|quoniam experimentum quaeritis eius, qui in me loquitur, Christi, qui in vos non infirmatur, sed potens est in vobis.
2COR|13|4|Nam etsi crucifixus est ex infirmitate, sed vivit ex virtute Dei. Nam et nos infirmi sumus in illo, sed vivemus cum eo ex virtute Dei in vos.
2COR|13|5|Vosmetipsos tentate, si estis in fide; ipsi vos probate. An non cognoscitis vos ipsos, quia Iesus Christus in vobis est? Nisi forte reprobi estis.
2COR|13|6|Spero autem quod cognoscetis quia nos non sumus reprobi.
2COR|13|7|Oramus autem Deum, ut nihil mali faciatis, non ut nos probati pareamus, sed ut vos, quod bonum est, faciatis, nos autem ut reprobi simus.
2COR|13|8|Non enim possumus aliquid adversus veritatem, sed pro veritate.
2COR|13|9|Gaudemus enim, quando nos infirmi sumus, vos autem potentes estis; hoc et oramus, vestram consummationem.
2COR|13|10|Ideo haec absens scribo, ut non praesens durius agam secundum potestatem, quam Dominus dedit mihi in aedificationem et non in destructionem.
2COR|13|11|De cetero, fratres, gaudete, perfecti estote, exhortamini invicem, idem sapite, pacem habete, et Deus dilectionis et pacis erit vobiscum.
2COR|13|12|Salutate invicem in osculo sancto. Salutant vos sancti omnes.
2COR|13|13|Gratia Domini Iesu Christi et caritas Dei et communicatio Sancti Spiritus cum omnibus vobis.
GAL|1|1|Paulus apostolus, non ab ho minibus neque per hominem, sed per Iesum Christum et Deum Patrem, qui suscitavit eum a mortuis,
GAL|1|2|et, qui mecum sunt, omnes fratres ecclesiis Galatiae:
GAL|1|3|gratia vobis et pax a Deo Patre nostro et Domino Iesu Christo,
GAL|1|4|qui dedit semetipsum pro peccatis nostris, ut eriperet nos de praesenti saeculo nequam secundum voluntatem Dei et Patris nostri,
GAL|1|5|cui gloria in saecula saeculorum. Amen.
GAL|1|6|Miror quod tam cito transferimini ab eo, qui vos vocavit in gratia Christi, in aliud evangelium;
GAL|1|7|quod non est aliud, nisi sunt aliqui, qui vos conturbant et volunt convertere evangelium Christi.
GAL|1|8|Sed licet nos aut angelus de caelo evangelizet vobis praeterquam quod evangelizavimus vobis, anathema sit!
GAL|1|9|Sicut praediximus, et nunc iterum dico: Si quis vobis evangelizaverit praeter id, quod accepistis, anathema sit!
GAL|1|10|Modo enim hominibus suadeo aut Deo? Aut quaero hominibus placere? Si adhuc hominibus placerem, Christi servus non essem!
GAL|1|11|Notum enim vobis facio, fratres, evangelium, quod evangelizatum est a me, quia non est secundum hominem;
GAL|1|12|neque enim ego ab homine accepi illud neque didici sed per revelationem Iesu Christi.
GAL|1|13|Audistis enim conversationem meam aliquando in Iudaismo, quoniam supra modum persequebar ecclesiam Dei et expugnabam illam;
GAL|1|14|et proficiebam in Iudaismo supra multos coaetaneos in genere meo, abundantius aemulator exsistens paternarum mearum traditionum.
GAL|1|15|Cum autem placuit Deo, qui me segregavit de utero matris meae et vocavit per gratiam suam,
GAL|1|16|ut revelaret Filium suum in me, ut evangelizarem illum in gentibus, continuo non contuli cum carne et sanguine
GAL|1|17|neque ascendi Hierosolymam ad antecessores meos apostolos; sed abii in Arabiam et iterum reversus sum Damascum.
GAL|1|18|Deinde post annos tres, ascendi Hierosolymam videre Cepham et mansi apud eum diebus quindecim;
GAL|1|19|alium autem apostolorum non vidi, nisi Iacobum fratrem Domini.
GAL|1|20|Quae autem scribo vobis, ecce coram Deo quia non mentior.
GAL|1|21|Deinde veni in partes Syriae et Ciliciae.
GAL|1|22|Eram autem ignotus facie ecclesiis Iudaeae, quae sunt in Christo;
GAL|1|23|tantum autem auditum habebant: " Qui persequebatur nos aliquando, nunc evangelizat fidem, quam aliquando expugnabat ",
GAL|1|24|et in me glorificabant Deum.
GAL|2|1|Deinde post annos quattuor decim, iterum ascendi Hieroso lymam cum Barnaba, assumpto et Tito;
GAL|2|2|ascendi autem secundum revelationem; et contuli cum illis evangelium, quod praedico in gentibus, seorsum autem his, qui observabantur, ne forte in vacuum currerem aut cucurrissem.
GAL|2|3|Sed neque Titus, qui mecum erat, cum esset Graecus, compulsus est circumcidi.
GAL|2|4|Sed propter subintroductos falsos fratres, qui subintroierunt explorare libertatem nostram, quam habemus in Christo Iesu, ut nos in servitutem redigerent;
GAL|2|5|quibus neque ad horam cessimus subicientes nos, ut veritas evangelii permaneat apud vos.
GAL|2|6|Ab his autem, qui videbantur esse aliquid - quales aliquando fuerint, nihil mea interest; Deus personam hominis non accipit - mihi enim, qui observabantur, nihil contulerunt,
GAL|2|7|sed e contra, cum vidissent quod creditum est mihi evangelium praeputii, sicut Petro circumcisionis
GAL|2|8|- qui enim operatus est Petro in apostolatum circumcisionis, operatus est et mihi inter gentes -
GAL|2|9|et cum cognovissent gratiam, quae data est mihi, Iacobus et Cephas et Ioannes, qui videbantur columnae esse, dexteras dederunt mihi et Barnabae communionis, ut nos in gentes, ipsi autem in circumcisionem;
GAL|2|10|tantum ut pauperum memores essemus, quod etiam sollicitus fui hoc ipsum facere.
GAL|2|11|Cum autem venisset Cephas Antiochiam, in faciem ei restiti, quia reprehensibilis erat.
GAL|2|12|Prius enim quam venirent quidam ab Iacobo, cum gentibus comedebat; cum autem venissent, subtrahebat et segregabat se, timens eos, qui ex circumcisione erant.
GAL|2|13|Et simulationi eius consenserunt ceteri Iudaei, ita ut et Barnabas simul abduceretur illorum simulatione.
GAL|2|14|Sed cum vidissem quod non recte ambularent ad veritatem evangelii, dixi Cephae coram omnibus: " Si tu, cum Iudaeus sis, gentiliter et non Iudaice vivis, quomodo gentes cogis iudaizare? ".
GAL|2|15|Nos natura Iudaei et non ex gentibus peccatores,
GAL|2|16|scientes autem quod non iustificatur homo ex operibus legis, nisi per fidem Iesu Christi, et nos in Christum Iesum credidimus, ut iustificemur ex fide Christi et non ex operibus legis, quoniam ex operibus legis non iustificabitur omnis caro.
GAL|2|17|Quodsi quaerentes iustificari in Christo, inventi sumus et ipsi peccatores, numquid Christus peccati minister est? Absit!
GAL|2|18|Si enim, quae destruxi, haec iterum aedifico, praevaricatorem me constituo.
GAL|2|19|Ego enim per legem legi mortuus sum, ut Deo vivam. Christo confixus sum cruci;
GAL|2|20|vivo autem iam non ego, vivit vero in me Christus; quod autem nunc vivo in carne, in fide vivo Filii Dei, qui dilexit me et tradidit seipsum pro me.
GAL|2|21|Non irritam facio gratiam Dei; si enim per legem iustitia, ergo Christus gratis mortuus est.
GAL|3|1|O insensati Galatae, quis vos fascinavit, ante quorum oculos Iesus Christus descriptus est crucifixus?
GAL|3|2|Hoc solum volo a vobis discere: Ex operibus legis Spiritum accepistis an ex auditu fidei?
GAL|3|3|Sic stulti estis? Cum Spiritu coeperitis, nunc carne consummamini?
GAL|3|4|Tanta passi estis sine causa? Si tamen et sine causa!
GAL|3|5|Qui ergo tribuit vobis Spiritum et operatur virtutes in vobis, ex operibus legis an ex auditu fidei?
GAL|3|6|Sicut Abraham credidit Deo, et reputatum est ei ad iustitiam.
GAL|3|7|Cognoscitis ergo quia qui ex fide sunt, hi sunt filii Abrahae.
GAL|3|8|Providens autem Scriptura, quia ex fide iustificat gentes Deus, praenuntiavit Abrahae: "Benedicentur in te omnes gentes".
GAL|3|9|Igitur, qui ex fide sunt, benedi cuntur cum fideli Abraham.
GAL|3|10|Quicumque enim ex operibus legis sunt, sub maledicto sunt; scriptum est enim: " Maledictus omnis, qui non permanserit in omnibus, quae scripta sunt in libro legis, ut faciat ea ".
GAL|3|11|Quoniam autem in lege nemo iustificatur apud Deum manifestum est, quia iustus ex fide vivet;
GAL|3|12|lex autem non est ex fide; sed, qui fecerit ea, vivet in illis.
GAL|3|13|Christus nos redemit de maledicto legis factus pro nobis maledictum, quia scriptum est: " Maledictus omnis, qui pendet in ligno ",
GAL|3|14|ut in gentes benedictio Abrahae fieret in Christo Iesu, ut promissionem Spiritus accipiamus per fidem.
GAL|3|15|Fratres, secundum hominem dico, tamen hominis confirmatum testamentum nemo irritum facit aut superordinat.
GAL|3|16|Abrahae autem dictae sunt promissiones et semini eius. Non dicit: " Et seminibus ", quasi in multis, sed quasi in uno: "Et semini tuo", qui est Christus.
GAL|3|17|Hoc autem dico: Testamentum confirmatum a Deo, quae post quadringentos et triginta annos facta est lex, non irritum facit ad evacuandam promissionem.
GAL|3|18|Nam si ex lege hereditas, iam non ex promissione; Abrahae autem per promissionem donavit Deus.
GAL|3|19|Quid igitur lex? Propter transgressiones apposita est, donec veniret semen, cui promissum est, ordinata per angelos in manu mediatoris.
GAL|3|20|Mediator autem unius non est, Deus autem unus est.
GAL|3|21|Lex ergo adversus promissa Dei? Absit. Si enim data esset lex, quae posset vivificare, vere ex lege esset iustitia.
GAL|3|22|Sed conclusit Scriptura omnia sub peccato, ut promissio ex fide Iesu Christi daretur credentibus.
GAL|3|23|Prius autem quam veniret fides, sub lege custodiebamur conclusi in eam fidem, quae revelanda erat.
GAL|3|24|Itaque lex paedagogus noster fuit in Christum, ut ex fide iustificemur;
GAL|3|25|at ubi venit fides, iam non sumus sub paedagogo.
GAL|3|26|Omnes enim filii Dei estis per fidem in Christo Iesu.
GAL|3|27|Quicumque enim in Christum baptizati estis, Christum induistis:
GAL|3|28|non est Iudaeus neque Graecus, non est servus neque liber, non est masculus et femina; omnes enim vos unus estis in Christo Iesu.
GAL|3|29|Si autem vos Christi, ergo Abrahae semen estis, secundum promissionem heredes.
GAL|4|1|Dico autem: Quanto tempore heres parvulus est, nihil differt a servo, cum sit dominus omnium,
GAL|4|2|sed sub tutoribus est et actoribus usque ad praefinitum tempus a patre.
GAL|4|3|Ita et nos, cum essemus parvuli, sub elementis mundi eramus servientes;
GAL|4|4|at ubi venit plenitudo temporis, misit Deus Filium suum, factum ex muliere, factum sub lege,
GAL|4|5|ut eos, qui sub lege erant, redimeret, ut adoptionem filiorum reciperemus.
GAL|4|6|Quoniam autem estis filii, misit Deus Spiritum Filii sui in corda nostra clamantem: " Abba, Pater! ".
GAL|4|7|Itaque iam non es servus sed filius; quod si filius, et heres per Deum.
GAL|4|8|Sed tunc quidem ignorantes Deum, his, qui natura non sunt dii, servistis;
GAL|4|9|nunc autem, cum cognoveritis Deum, immo cogniti sitis a Deo, quomodo convertimini iterum ad infirma et egena elementa, quibus rursus ut antea servire vultis?
GAL|4|10|Dies observatis et menses et tempora et annos!
GAL|4|11|Timeo vos, ne forte sine causa laboraverim in vobis.
GAL|4|12|Estote sicut ego, quia et ego sicut vos; fratres, obsecro vos. Nihil me laesistis;
GAL|4|13|scitis autem quia per infirmitatem carnis pridem vobis evangelizavi,
GAL|4|14|et tentationem vestram in carne mea non sprevistis neque respuistis, sed sicut angelum Dei excepistis me, sicut Christum Iesum.
GAL|4|15|Ubi est ergo beatitudo vestra? Testimonium enim perhibeo vobis, quia, si fieri posset, oculos vestros eruissetis et dedissetis mihi.
GAL|4|16|Ergo inimicus vobis factus sum, verum dicens vobis?
GAL|4|17|Aemulantur vos non bene, sed excludere vos volunt, ut illos aemulemini.
GAL|4|18|Bonum est autem aemulari in bono semper, et non tantum cum praesens sum apud vos,
GAL|4|19|filioli mei, quos iterum parturio, donec formetur Christus in vobis!
GAL|4|20|Vellem autem esse apud vos modo et mutare vocem meam, quoniam incertus sum in vobis.
GAL|4|21|Dicite mihi, qui sub lege vultis esse: Legem non auditis?
GAL|4|22|Scriptum est enim quoniam Abraham duos filios habuit, unum de ancilla et unum de libera.
GAL|4|23|Sed qui de ancilla, secundum carnem natus est; qui autem de libera, per promissionem.
GAL|4|24|Quae sunt per allegoriam dicta; ipsae enim sunt duo Testamenta, unum quidem a monte Sinai, in servitutem generans, quod est Agar.
GAL|4|25|Illud vero Agar mons est Sinai in Arabia, respondet autem Ierusalem, quae nunc est; servit enim cum filiis suis.
GAL|4|26|Illa autem, quae sursum est Ierusalem, libera est, quae est mater nostra;
GAL|4|27|scriptum est enim: Laetare, sterilis, quae non paris,erumpe et exclama, quae non parturis,quia multi filii desertaemagis quam eius, quae habet virum ".
GAL|4|28|Vos autem, fratres, secundum Isaac promissionis filii estis.
GAL|4|29|Sed quomodo tunc, qui secundum carnem natus fuerat, persequebatur eum, qui secundum spiritum, ita et nunc.
GAL|4|30|Sed quid dicit Scriptura? " Eice ancillam et filium eius; non enim heres erit filius ancillae cum filio liberae ".
GAL|4|31|Itaque, fratres, non sumus ancillae filii sed liberae.
GAL|5|1|Hac libertate nos Christus liberavit; state igitur et nolite iterum iugo servitutis detineri.
GAL|5|2|Ecce ego Paulus dico vobis quoniam, si circumcidamini, Christus vobis nihil proderit.
GAL|5|3|Testificor autem rursum omni homini circumcidenti se quoniam debitor est universae legis faciendae.
GAL|5|4|Evacuati estis a Christo, qui in lege iustificamini, a gratia excidistis.
GAL|5|5|Nos enim Spiritu ex fide spem iustitiae exspectamus.
GAL|5|6|Nam in Christo Iesu neque circumcisio aliquid valet neque praeputium, sed fides, quae per caritatem operatur.
GAL|5|7|Currebatis bene; quis vos impedivit veritati non oboedire?
GAL|5|8|Haec persuasio non est ex eo, qui vocat vos.
GAL|5|9|Modicum fermentum totam massam corrumpit.
GAL|5|10|Ego confido in vobis in Domino, quod nihil aliud sapietis; qui autem conturbat vos, portabit iudicium, quicumque est ille.
GAL|5|11|Ego autem, fratres, si circumcisionem adhuc praedico, quid adhuc persecutionem patior? Ergo evacuatum est scandalum crucis.
GAL|5|12|Utinam et abscidantur, qui vos conturbant!
GAL|5|13|Vos enim in libertatem vocati estis, fratres; tantum ne libertatem in occasionem detis carni, sed per caritatem servite invicem.
GAL|5|14|Omnis enim lex in uno sermone impletur, in hoc: Diliges proximum tuum sicut teipsum.
GAL|5|15|Quod si invicem mordetis et devoratis, videte, ne ab invicem consumamini!
GAL|5|16|Dico autem: Spiritu ambulate et concupiscentiam carnis ne perfeceritis.
GAL|5|17|Caro enim concupiscit adversus Spiritum, Spiritus autem adversus carnem; haec enim invicem adversantur, ut non, quaecumque vultis, illa faciatis.
GAL|5|18|Quod si Spiritu ducimini, non estis sub lege.
GAL|5|19|Manifesta autem sunt opera carnis, quae sunt fornicatio, immunditia, luxuria,
GAL|5|20|idolorum servitus, veneficia, inimicitiae, contentiones, aemulationes, irae, rixae, dissensiones, sectae,
GAL|5|21|invidiae, ebrietates, comissationes et his similia; quae praedico vobis, sicut praedixi, quoniam, qui talia agunt, regnum Dei non consequentur.
GAL|5|22|Fructus autem Spiritus est caritas, gaudium, pax, longanimitas, benignitas, bonitas, fides,
GAL|5|23|mansuetudo, continentia; adversus huiusmodi non est lex.
GAL|5|24|Qui autem sunt Christi Iesu, carnem crucifixerunt cum vitiis et concupiscentiis.
GAL|5|25|Si vivimus Spiritu, Spiritu et ambulemus.
GAL|5|26|Non efficiamur inanis gloriae cupidi, invicem provocantes, invicem invidentes.
GAL|6|1|Fratres, et si praeoccupatus fuerit homo in aliquo delicto, vos, qui spiritales estis, huiusmodi instruite in spiritu lenitatis, considerans teipsum, ne et tu tenteris.
GAL|6|2|Alter alterius onera portate et sic adimplebitis legem Christi.
GAL|6|3|Nam si quis existimat se aliquid esse, cum sit nihil, ipse se seducit;
GAL|6|4|opus autem suum probet unusquisque et sic in semetipso tantum gloriationem habebit et non in altero.
GAL|6|5|Unusquisque enim onus suum portabit.
GAL|6|6|Communicet autem is, qui catechizatur verbum, ei qui se catechizat, in omnibus bonis.
GAL|6|7|Nolite errare: Deus non irridetur. Quae enim seminaverit homo, haec et metet;
GAL|6|8|quoniam, qui seminat in carne sua, de carne metet corruptionem; qui autem seminat in Spiritu, de Spiritu metet vitam aeternam.
GAL|6|9|Bonum autem facientes infatigabiles, tempore enim suo metemus non deficientes.
GAL|6|10|Ergo dum tempus habemus, operemur bonum ad omnes, maxime autem ad domesticos fidei.
GAL|6|11|Videte qualibus litteris scripsi vobis mea manu.
GAL|6|12|Quicumque volunt placere in carne, hi cogunt vos circumcidi, tantum ut crucis Christi persecutionem non patiantur;
GAL|6|13|neque enim, qui circumciduntur, legem custodiunt, sed volunt vos circumcidi, ut in carne vestra glorientur.
GAL|6|14|Mihi autem absit gloriari, nisi in cruce Domini nostri Iesu Christi, per quem mihi mundus crucifixus est, et ego mundo.
GAL|6|15|Neque enim circumcisio aliquid est neque praeputium sed nova creatura.
GAL|6|16|Et quicumque hanc regulam secuti fuerint, pax super illos et misericordia et super Israel Dei.
GAL|6|17|De cetero nemo mihi molestus sit; ego enim stigmata Iesu in super corpore meo porto.
GAL|6|18|Gratia Domini nostri Iesu Christi cum spiritu vestro, fratres. Amen.
EPH|1|1|Paulus, apostolus Christi Iesu per voluntatem Dei, sanctis, qui sunt Ephesi, et fidelibus in Christo Iesu:
EPH|1|2|gratia vobis et pax a Deo Patre nostro et Domino Iesu Christo.
EPH|1|3|Benedictus Deus et Pater Domini nostri Iesu Christi,qui benedixit nos in omni benedictione spiritali in caelestibus in Christo,
EPH|1|4|sicut elegit nos in ipso ante mundi constitutionem,ut essemus sancti et immaculati in conspectu eius in caritate;
EPH|1|5|qui praedestinavit nos in adoptionem filiorumper Iesum Christum in ipsum,secundum beneplacitum voluntatis suae,
EPH|1|6|in laudem gloriae gratiae suae,in qua gratificavit nos in Dilecto,
EPH|1|7|in quo habemus redemptionem per sanguinem eius,remissionem peccatorum,secundum divitias gratiae eius,
EPH|1|8|quam superabundare fecit in nobisin omni sapientia et prudentia,
EPH|1|9|notum faciens nobis mysterium voluntatis suae,secundum beneplacitum eius, quod proposuit in eo,
EPH|1|10|in dispensationem plenitudinis temporum:recapitulare omnia in Christo,quae in caelis et quae in terra, in ipso;
EPH|1|11|in quo etiam sorte vocati sumus, praedestinati secundum propositum eius, qui omnia operatur secundum consilium voluntatis suae,
EPH|1|12|ut simus in laudem gloriae eius, qui ante speravimus in Christo;
EPH|1|13|in quo et vos cum audissetis verbum veritatis, evangelium salutis vestrae, in quo et credentes signati estis Spiritu promissionis Sancto,
EPH|1|14|qui est arrabo hereditatis nostrae in redemptionem acquisitionis, in laudem gloriae ipsius.
EPH|1|15|Propterea et ego audiens fidem vestram, quae est in Domino Iesu, et dilectionem in omnes sanctos,
EPH|1|16|non cesso gratias agens pro vobis memoriam faciens in orationibus meis,
EPH|1|17|ut Deus Domini nostri Iesu Christi, Pater gloriae, det vobis Spiritum sapientiae et revelationis in agnitione eius,
EPH|1|18|illuminatos oculos cordis vestri, ut sciatis quae sit spes vocationis eius, quae divitiae gloriae hereditatis eius in sanctis,
EPH|1|19|et quae sit supereminens magnitudo virtutis eius in nos, qui credimus, secundum operationem potentiae virtutis eius,
EPH|1|20|quam operatus est in Christo, suscitans illum a mortuis et constituens ad dexteram suam in caelestibus
EPH|1|21|supra omnem principatum et potestatem et virtutem et dominationem et omne nomen, quod nominatur non solum in hoc saeculo sed et in futuro;
EPH|1|22|et omnia subiecit sub pedibus eius et ipsum dedit caput supra omnia ecclesiae,
EPH|1|23|quae est corpus ipsius, plenitudo eius, qui omnia in omnibus adimpletur.
EPH|2|1|Et vos, cum essetis mortui de lictis et peccatis vestris,
EPH|2|2|in qui bus aliquando ambulastis secundum saeculum mundi huius, secundum principem potestatis aeris, spiritus, qui nunc operatur in filios diffidentiae;
EPH|2|3|in quibus et nos omnes aliquando conversati sumus in concupiscentiis carnis nostrae, facientes voluntates carnis et cogitationum, et eramus natura filii irae, sicut et ceteri.
EPH|2|4|Deus autem, qui dives est in misericordia, propter nimiam caritatem suam, qua dilexit nos,
EPH|2|5|et cum essemus mortui peccatis, convivificavit nos Christo - gratia estis salvati -
EPH|2|6|et conresuscitavit et consedere fecit in caelestibus in Christo Iesu,
EPH|2|7|ut ostenderet in saeculis supervenientibus abundantes divitias gratiae suae in bonitate super nos in Christo Iesu.
EPH|2|8|Gratia enim estis salvati per fidem; et hoc non ex vobis, Dei donum est:
EPH|2|9|non ex operibus, ut ne quis glorietur.
EPH|2|10|Ipsius enim sumus factura, creati in Christo Iesu in opera bona, quae praeparavit Deus, ut in illis ambulemus.
EPH|2|11|Propter quod memores estote, quod aliquando vos gentes in carne, qui dicimini praeputium ab ea, quae dicitur circumcisio in carne manufacta,
EPH|2|12|quia eratis illo in tempore sine Christo, alienati a conversatione Israel et extranei testamentorum promissionis, spem non habentes et sine Deo in mundo.
EPH|2|13|Nunc autem in Christo Iesu vos, qui aliquando eratis longe, facti estis prope in sanguine Christi.
EPH|2|14|Ipse est enim pax nostra, qui fecit utraque unum et medium parietem maceriae solvit, inimicitiam, in carne sua,
EPH|2|15|legem mandatorum in decretis evacuans, ut duos condat in semetipso in unum novum hominem, faciens pacem,
EPH|2|16|et reconciliet ambos in uno corpore Deo per crucem, interficiens inimicitiam in semetipso.
EPH|2|17|Et veniens evangelizavit pacem vobis, qui longe fuistis, et pacem his, qui prope;
EPH|2|18|quoniam per ipsum habemus accessum ambo in uno Spiritu ad Patrem.
EPH|2|19|Ergo iam non estis extranei et advenae, sed estis concives sanctorum et domestici Dei,
EPH|2|20|superaedificati super fundamentum apostolorum et prophetarum, ipso summo angulari lapide Christo Iesu,
EPH|2|21|in quo omnis aedificatio compacta crescit in templum sanctum in Domino,
EPH|2|22|in quo et vos coaedificamini in habitaculum Dei in Spiritu.
EPH|3|1|Huius rei gratia, ego Paulus, vinctus Christi Iesu pro vobis gentibus -
EPH|3|2|si tamen audistis dispensationem gratiae Dei, quae data est mihi pro vobis,
EPH|3|3|quoniam secundum revelationem notum mihi factum est mysterium, sicut supra scripsi in brevi,
EPH|3|4|prout potestis legentes intellegere prudentiam meam in mysterio Christi,
EPH|3|5|quod aliis generationibus non innotuit filiis hominum, sicuti nunc revelatum est sanctis apostolis eius et prophetis in Spiritu,
EPH|3|6|esse gentes coheredes et concorporales et comparticipes promissionis in Christo Iesu per evangelium,
EPH|3|7|cuius factus sum minister secundum donum gratiae Dei, quae data est mihi secundum operationem virtutis eius.
EPH|3|8|Mihi omnium sanctorum minimo data est gratia haec: gentibus evangelizare investigabiles divitias Christi
EPH|3|9|et illuminare omnes, quae sit dispensatio mysterii absconditi a saeculis in Deo, qui omnia creavit,
EPH|3|10|ut innotescat nunc principatibus et potestatibus in caelestibus per ecclesiam multiformis sapientia Dei,
EPH|3|11|secundum propositum saeculorum, quod fecit in Christo Iesu Domino nostro,
EPH|3|12|in quo habemus fiduciam et accessum in confidentia per fidem eius.
EPH|3|13|Propter quod peto, ne deficiatis in tribulationibus meis pro vobis, quae est gloria vestra.
EPH|3|14|Huius rei gratia flecto genua mea ad Patrem,
EPH|3|15|ex quo omnis paternitas in caelis et in terra nominatur,
EPH|3|16|ut det vobis secundum divitias gloriae suae virtute corroborari per Spiritum eius in interiorem hominem,
EPH|3|17|habitare Christum per fidem in cordibus vestris, in caritate radicati et fundati,
EPH|3|18|ut valeatis comprehendere cum omnibus sanctis quae sit latitudo et longitudo et sublimitas et profundum,
EPH|3|19|scire etiam supereminentem scientiae caritatem Christi, ut impleamini in omnem plenitudinem Dei.
EPH|3|20|Ei autem, qui potens est supra omnia facere superabundanter quam petimus aut intellegimus, secundum virtutem, quae operatur in nobis,
EPH|3|21|ipsi gloria in ecclesia et in Christo Iesu in omnes generationes saeculi saeculorum. Amen.
EPH|4|1|Obsecro itaque vos ego, vinctus in Domino, ut digne ambuletis vocatione, qua vocati estis,
EPH|4|2|cum omni humilitate et mansuetudine, cum longanimitate, supportantes invicem in caritate,
EPH|4|3|solliciti servare unitatem spiritus in vinculo pacis;
EPH|4|4|unum corpus et unus Spiritus, sicut et vocati estis in una spe vocationis vestrae;
EPH|4|5|unus Dominus, una fides, unum baptisma;
EPH|4|6|unus Deus et Pater omnium, qui super omnes et per omnia et in omnibus.
EPH|4|7|Unicuique autem nostrum data est gratia secundum mensuram donationis Christi.
EPH|4|8|Propter quod dicit: Ascendens in altum captivam duxit captivitatem,dedit dona hominibus ".
EPH|4|9|Illud autem " ascendit " quid est, nisi quia et descendit in inferiores partes terrae?
EPH|4|10|Qui descendit, ipse est et qui ascendit super omnes caelos, ut impleret omnia.
EPH|4|11|Et ipse dedit quosdam quidem apostolos, quosdam autem prophetas, alios vero evangelistas, alios autem pastores et doctores
EPH|4|12|ad instructionem sanctorum in opus ministerii, in aedificationem corporis Christi,
EPH|4|13|donec occurramus omnes in unitatem fidei et agnitionis Filii Dei, in virum perfectum, in mensuram aetatis plenitudinis Christi,
EPH|4|14|ut iam non simus parvuli fluctuantes et circumacti omni vento doctrinae in fallacia hominum, in astutia ad circumventionem erroris;
EPH|4|15|veritatem autem facientes in caritate crescamus in illum per omnia, qui est caput Christus,
EPH|4|16|ex quo totum corpus compactum et conexum per omnem iuncturam subministrationis secundum operationem in mensura uniuscuiusque partis augmentum corporis facit in aedificationem sui in caritate.
EPH|4|17|Hoc igitur dico et testificor in Domino, ut iam non ambuletis, sicut et gentes ambulant in vanitate sensus sui
EPH|4|18|tenebris obscuratum habentes intellectum, alienati a vita Dei propter ignorantiam, quae est in illis propter caecitatem cordis ipsorum;
EPH|4|19|qui indolentes semetipsos tradiderunt impudicitiae in operationem immunditiae omnis in avaritia.
EPH|4|20|Vos autem non ita didicistis Christum,
EPH|4|21|si tamen illum audistis et in ipso edocti estis, sicut est veritas in Iesu:
EPH|4|22|deponere vos secundum pristinam conversationem veterem hominem, qui corrumpitur secundum desideria erroris,
EPH|4|23|renovari autem spiritu mentis vestrae
EPH|4|24|et induere novum hominem, qui secundum Deum creatus est in iustitia et sanctitate veritatis.
EPH|4|25|Propter quod deponentes mendacium loquimini veritatem unusquisque cum proximo suo, quoniam sumus invicem membra.
EPH|4|26|Irascimini et nolite peccare; sol non occidat super iracundiam vestram,
EPH|4|27|et nolite locum dare Diabolo.
EPH|4|28|Qui furabatur, iam non furetur, magis autem laboret operando manibus bonum, ut habeat unde tribuat necessitatem patienti.
EPH|4|29|Omnis sermo malus ex ore vestro non procedat, sed si quis bonus ad aedificationem opportunitatis, ut det gratiam audientibus.
EPH|4|30|Et nolite contristare Spiritum Sanctum Dei, in quo signati estis in diem redemptionis.
EPH|4|31|Omnis amaritudo et ira et indignatio et clamor et blasphemia tollatur a vobis cum omni malitia.
EPH|4|32|Estote autem invicem benigni, misericordes, donantes invicem, sicut et Deus in Christo donavit vobis.
EPH|5|1|Estote ergo imitatores Dei, sicut filii carissimi,
EPH|5|2|et ambulate in dilectione, sicut et Christus dilexit nos et tradidit seipsum pro nobis oblationem et hostiam Deo in odorem suavitatis.
EPH|5|3|Fornicatio autem et omnis immunditia aut avaritia nec nominetur in vobis, sicut decet sanctos,
EPH|5|4|et turpitudo et stultiloquium aut scurrilitas, quae non decent, sed magis gratiarum actio.
EPH|5|5|Hoc enim scitote intellegentes quod omnis fornicator aut immundus aut avarus, id est idolorum cultor, non habet hereditatem in regno Christi et Dei.
EPH|5|6|Nemo vos decipiat inanibus verbis; propter haec enim venit ira Dei in filios diffidentiae.
EPH|5|7|Nolite ergo effici comparticipes eorum;
EPH|5|8|eratis enim aliquando tenebrae, nunc autem lux in Domino. Ut filii lucis ambulate
EPH|5|9|- fructus enim lucis est in omni bonitate et iustitia et veritate -
EPH|5|10|probantes quid sit beneplacitum Domino;
EPH|5|11|et nolite communicare operibus infructuosis tenebrarum, magis autem et redarguite;
EPH|5|12|quae enim in occulto fiunt ab ipsis, turpe est et dicere;
EPH|5|13|omnia autem, quae arguuntur, a lumine manifestantur,
EPH|5|14|omne enim, quod manifestatur, lumen est. Propter quod dicit: " Surge, qui dormis, et exsurge a mortuis, et illuminabit te Christus ".
EPH|5|15|Videte itaque caute quomodo ambuletis, non quasi insipientes sed ut sapientes,
EPH|5|16|redimentes tempus, quoniam dies mali sunt.
EPH|5|17|Propterea nolite fieri imprudentes, sed intellegite, quae sit voluntas Domini.
EPH|5|18|Et nolite inebriari vino, in quo est luxuria, sed implemini Spiritu
EPH|5|19|loquentes vobismetipsis in psalmis et hymnis et canticis spiritalibus, cantantes et psallentes in cordibus vestris Domino.
EPH|5|20|Gratias agentes semper pro omnibus in nomine Domini nostri Iesu Christi Deo et Patri,
EPH|5|21|subiecti invicem in timore Christi.
EPH|5|22|Mulieres viris suis sicut Domino,
EPH|5|23|quoniam vir caput est mulieris, sicut et Christus caput est ecclesiae, ipse salvator corporis.
EPH|5|24|Sed ut ecclesia subiecta est Christo, ita et mulieres viris in omnibus.
EPH|5|25|Viri, diligite uxores, sicut et Christus dilexit ecclesiam et seipsum tradidit pro ea,
EPH|5|26|ut illam sanctificaret mundans lavacro aquae in verbo,
EPH|5|27|ut exhiberet ipse sibi gloriosam ecclesiam non habentem maculam aut rugam aut aliquid eiusmodi, sed ut sit sancta et immaculata.
EPH|5|28|Ita et viri debent diligere uxores suas ut corpora sua. Qui suam uxorem diligit, seipsum diligit;
EPH|5|29|nemo enim umquam carnem suam odio habuit, sed nutrit et fovet eam sicut et Christus ecclesiam,
EPH|5|30|quia membra sumus corporis eius.
EPH|5|31|Propter hoc relinquet homo patrem et matrem et adhaerebit uxori suae, et erunt duo in carne una.
EPH|5|32|Mysterium hoc magnum est; ego autem dico de Christo et ecclesia!
EPH|5|33|Verumtamen et vos singuli unusquisque suam uxorem sicut seipsum diligat; uxor autem timeat virum.
EPH|6|1|Filii, oboedite parentibus vestris in Domino; hoc enim est iu stum.
EPH|6|2|Honora patrem tuum et matrem, quod est mandatum primum cum promissione,
EPH|6|3|ut bene sit tibi, et sis longaevus super terram.
EPH|6|4|Et, patres, nolite ad iracundiam provocare filios vestros, sed educate illos in disciplina et correptione Domini.
EPH|6|5|Servi, oboedite dominis carnalibus cum timore et tremore, in simplicitate cordis vestri, sicut Christo;
EPH|6|6|non ad oculum servientes, quasi hominibus placentes, sed ut servi Christi facientes voluntatem Dei ex animo;
EPH|6|7|cum bona voluntate servientes, sicut Domino et non hominibus,
EPH|6|8|scientes quoniam unusquisque, si quid fecerit bonum, hoc percipiet a Domino, sive servus sive liber.
EPH|6|9|Et, domini, eadem facite illis, remittentes minas, scientes quia et illorum et vester Dominus est in caelis, et personarum acceptio non est apud eum.
EPH|6|10|De cetero confortamini in Domino et in potentia virtutis eius.
EPH|6|11|Induite armaturam Dei, ut possitis stare adversus insidias Diaboli.
EPH|6|12|Quia non est nobis colluctatio adversus sanguinem et carnem sed adversus principatus, adversus potestates, adversus mundi rectores tenebrarum harum, adversus spiritalia nequitiae in caelestibus.
EPH|6|13|Propterea accipite armaturam Dei, ut possitis resistere in die malo et, omnibus perfectis, stare.
EPH|6|14|State ergo succincti lumbos vestros in veritate et induti loricam iustitiae
EPH|6|15|et calceati pedes in praeparatione evangelii pacis,
EPH|6|16|inomnibus sumentes scutum fidei, in quo possitis omnia tela Maligni ignea exstinguere;
EPH|6|17|et galeam salutis assumite et gladium Spiritus, quod est verbum Dei;
EPH|6|18|per omnem orationem et obsecrationem orantes omni tempore in Spiritu, et in ipso vigilantes in omni instantia et obsecratione pro omnibus sanctis
EPH|6|19|et pro me, ut detur mihi sermo in aperitione oris mei cum fiducia notum facere mysterium evangelii,
EPH|6|20|pro quo legatione fungor in catena, ut in ipso audeam, prout oportet me, loqui.
EPH|6|21|Ut autem et vos sciatis, quae circa me sunt, quid agam, omnia nota vobis faciet Tychicus, carissimus frater et fidelis minister in Domino,
EPH|6|22|quem misi ad vos in hoc ipsum, ut cognoscatis, quae circa nos sunt, et consoletur corda vestra.
EPH|6|23|Pax fratribus et caritas cum fide a Deo Patre et Domino Iesu Christo.
EPH|6|24|Gratia cum omnibus, qui diligunt Dominum nostrum Iesum Christum in incorruptione.
PHIL|1|1|Paulus et Timotheus servi Christi Iesu omnibus sanctis in Christo Iesu, qui sunt Philippis, cum episcopis et diaconis:
PHIL|1|2|gratia vobis et pax a Deo Patre nostro et Domino Iesu Christo.
PHIL|1|3|Gratias ago Deo meo in omni memoria vestri,
PHIL|1|4|semper in omni oratione mea pro omnibus vobis cum gaudio deprecationem faciens
PHIL|1|5|super communione vestra in evangelio a prima die usque nunc;
PHIL|1|6|confidens hoc ipsum, quia, qui coepit in vobis opus bonum, perficiet usque in diem Christi Iesu;
PHIL|1|7|sicut est mihi iustum hoc sentire pro omnibus vobis, eo quod habeam in corde vos et in vinculis meis et in defensione et confirmatione evangelii socios gratiae meae omnes vos esse.
PHIL|1|8|Testis enim mihi Deus, quomodo cupiam omnes vos in visceribus Christi Iesu.
PHIL|1|9|Et hoc oro, ut caritas vestra magis ac magis abundet in scientia et omni sensu,
PHIL|1|10|ut probetis potiora, ut sitis sinceri et sine offensa in diem Christi,
PHIL|1|11|repleti fructu iustitiae, qui est per Iesum Christum, in gloriam et laudem Dei.
PHIL|1|12|Scire autem vos volo, fratres, quia, quae circa me sunt, magis ad profectum venerunt evangelii,
PHIL|1|13|ita ut vincula mea manifesta fierent in Christo in omni praetorio et in ceteris omnibus;
PHIL|1|14|et plures e fratribus in Domino confidentes vinculis meis, abundantius audere sine timore verbum loqui.
PHIL|1|15|Quidam quidem et propter invidiam et contentionem, quidam autem et propter bonam voluntatem Christum praedicant;
PHIL|1|16|hi quidem ex caritate scientes quoniam in defensionem evangelii positus sum,
PHIL|1|17|illi autem ex contentione Christum annuntiant, non sincere, existimantes pressuram se suscitare vinculis meis.
PHIL|1|18|Quid enim? Dum omni modo, sive sub obtentu sive in veritate, Christus annuntietur, et in hoc gaudeo; sed et gaudebo,
PHIL|1|19|scio enim quia hoc mihi proveniet in salutem per vestram orationem et subministrationem Spiritus Iesu Christi,
PHIL|1|20|secundum exspectationem et spem meam quia in nullo confundar, sed in omni fiducia, sicut semper et nunc, magnificabitur Christus in corpore meo, sive per vitam sive per mortem.
PHIL|1|21|Mihi enim vivere Christus est et mori lucrum.
PHIL|1|22|Quod si vivere in carne, hic mihi fructus operis est, et quid eligam ignoro.
PHIL|1|23|Coartor autem ex his duobus: desiderium habens dissolvi et cum Christo esse, multo magis melius;
PHIL|1|24|permanere autem in carne, magis necessarium est propter vos.
PHIL|1|25|Et hoc confidens, scio quia manebo et permanebo omnibus vobis ad profectum vestrum et gaudium fidei,
PHIL|1|26|ut gloriatio vestra abundet in Christo Iesu in me, per meum adventum iterum ad vos.
PHIL|1|27|Tantum digne evangelio Christi conversamini, ut sive cum venero et videro vos, sive absens audiam de vobis quia statis in uno Spiritu unanimes, concertantes fide evangelii;
PHIL|1|28|et in nullo perterriti ab adversariis, quod est illis indicium perditionis, vobis autem salutis, et hoc a Deo;
PHIL|1|29|quia vobis hoc donatum est pro Christo, non solum ut in eum credatis, sed ut etiam pro illo patiamini
PHIL|1|30|idem certamen habentes, quale vidistis in me et nunc auditis in me.
PHIL|2|1|Si qua ergo consolatio in Christo, si quod solacium cari tatis, si qua communio spiritus, si quae viscera et miserationes,
PHIL|2|2|implete gaudium meum, ut idem sapiatis, eandem caritatem habentes, unanimes, id ipsum sapientes;
PHIL|2|3|nihil per contentionem neque per inanem gloriam, sed in humilitate superiores sibi invicem arbitrantes;
PHIL|2|4|non, quae sua sunt, singuli considerantes, sed et ea, quae aliorum.
PHIL|2|5|Hoc sentite in vobis, quod et in Christo Iesu:
PHIL|2|6|qui cum in forma Dei esset,non rapinam arbitratus est esse se aequalem Deo,
PHIL|2|7|sed semetipsum exinanivit formam servi accipiens,in similitudinem hominum factus;et habitu inventus ut homo,
PHIL|2|8|humiliavit semetipsum factus oboediens usque ad mortem,mortem autem crucis.
PHIL|2|9|Propter quod et Deus illum exaltavitet donavit illi nomen,quod est super omne nomen,
PHIL|2|10|ut in nomine Iesu omne genu flectaturcaelestium et terrestrium et infernorum,
PHIL|2|11|et omnis lingua confiteatur Dominus Iesus Christus! ",in gloriam Dei Patris.
PHIL|2|12|Itaque, carissimi mei, sicut semper oboedistis, non ut in praesentia mei tantum sed multo magis nunc in absentia mea, cum metu et tremore vestram salutem operamini;
PHIL|2|13|Deus est enim, qui operatur in vobis et velle et perficere pro suo beneplacito.
PHIL|2|14|Omnia facite sine murmurationibus et haesitationibus,
PHIL|2|15|ut efficiamini sine querela et simplices, filii Dei sine reprehensione in medio generationis pravae et perversae, inter quos lucetis sicut luminaria in mundo,
PHIL|2|16|verbum vitae firmiter tenentes ad gloriam meam in die Christi, quia non in vacuum cucurri neque in vacuum laboravi.
PHIL|2|17|Sed et si delibor supra sacrificium et obsequium fidei vestrae, gaudeo et congaudeo omnibus vobis;
PHIL|2|18|idipsum autem et vos gaudete et congaudete mihi.
PHIL|2|19|Spero autem in Domino Iesu Timotheum cito me mittere ad vos, ut et ego bono animo sim, cognitis, quae circa vos sunt.
PHIL|2|20|Neminem enim habeo tam unanimem, qui sincere pro vobis sollicitus sit;
PHIL|2|21|omnes enim sua quaerunt, non quae sunt Iesu Christi.
PHIL|2|22|Probationem autem eius cognoscitis, quoniam sicut patri filius mecum servivit in evangelium.
PHIL|2|23|Hunc igitur spero me mittere, mox ut videro, quae circa me sunt;
PHIL|2|24|confido autem in Domino, quoniam et ipse cito veniam.
PHIL|2|25|Necessarium autem existimavi Epaphroditum fratrem et cooperatorem et commilitonem meum, vestrum autem apostolum et ministrum necessitatis meae, mittere ad vos,
PHIL|2|26|quoniam omnes vos desiderabat et maestus erat, propterea quod audieratis illum infirmatum.
PHIL|2|27|Nam et infirmatus est usque ad mortem, sed Deus misertus est eius; non solum autem eius, verum et mei, ne tristitiam super tristitiam haberem.
PHIL|2|28|Festinantius ergo misi illum, ut, viso eo, iterum gaudeatis, et ego sine tristitia sim.
PHIL|2|29|Excipite itaque illum in Domino cum omni gaudio et eiusmodi cum honore habetote,
PHIL|2|30|quoniam propter opus Christi usque ad mortem accessit in interitum tradens animam suam, ut suppleret id, quod vobis deerat ministerii erga me.
PHIL|3|1|De cetero, fratres mei, gaudete in Domino. Eadem vobis scribe re mihi quidem non pigrum, vobis autem securum.
PHIL|3|2|Videte canes, videte malos operarios, videte concisionem!
PHIL|3|3|Nos enim sumus circumcisio, qui Spiritu Dei servimus et gloriamur in Christo Iesu et non in carne fiduciam habentes,
PHIL|3|4|quamquam ego habeam confidentiam et in carne. Si quis alius videtur confidere in carne, ego magis:
PHIL|3|5|circumcisus octava die, ex genere Israel, de tribu Beniamin, Hebraeus ex Hebraeis, secundum legem pharisaeus,
PHIL|3|6|secundum aemulationem persequens ecclesiam, secundum iustitiam, quae in lege est, conversatus sine querela.
PHIL|3|7|Sed, quae mihi erant lucra, haec arbitratus sum propter Christum detrimentum.
PHIL|3|8|Verumtamen existimo omnia detrimentum esse propter eminentiam scientiae Christi Iesu Domini mei, propter quem omnia detrimentum feci et arbitror ut stercora, ut Christum lucrifaciam
PHIL|3|9|et inveniar in illo non habens meam iustitiam, quae ex lege est, sed illam, quae per fidem est Christi, quae ex Deo est iustitia in fide;
PHIL|3|10|ad cognoscendum illum et virtutem resurrectionis eius et communionem passionum illius, conformans me morti eius,
PHIL|3|11|si quo modo occurram ad resurrectionem, quae est ex mortuis.
PHIL|3|12|Non quod iam acceperim aut iam perfectus sim; persequor autem si umquam comprehendam, sicut et comprehensus sum a Christo Iesu.
PHIL|3|13|Fratres, ego me non arbitror comprehendisse; unum autem: quae quidem retro sunt, obliviscens, ad ea vero, quae ante sunt, extendens me
PHIL|3|14|ad destinatum persequor, ad bravium supernae vocationis Dei in Christo Iesu.
PHIL|3|15|Quicumque ergo perfecti, hoc sentiamus; et si quid aliter sapitis, et hoc vobis Deus revelabit;
PHIL|3|16|verumtamen, ad quod pervenimus, in eodem ambulemus.
PHIL|3|17|Coimitatores mei estote, fratres, et observate eos, qui ita ambulant, sicut habetis formam nos.
PHIL|3|18|Multi enim ambulant, quos saepe dicebam vobis, nunc autem et flens dico, inimicos crucis Christi,
PHIL|3|19|quorum finis interitus, quorum deus venter et gloria in confusione ipsorum, qui terrena sapiunt.
PHIL|3|20|Noster enim municipatus in caelis est, unde etiam salvatorem exspectamus Dominum Iesum Christum,
PHIL|3|21|qui transfigurabit corpus humilitatis nostrae, ut illud conforme faciat corpori gloriae suae secundum operationem, qua possit etiam subicere sibi omnia.
PHIL|4|1|Itaque, fratres mei carissimi et desideratissimi, gaudium et co rona mea, sic state in Domino, carissimi!
PHIL|4|2|Evodiam rogo et Syntychen deprecor idipsum sapere in Domino.
PHIL|4|3|Etiam rogo et te, germane compar, adiuva illas, quae mecum concertaverunt in evangelio cum Clemente et ceteris adiutoribus meis, quorum nomina sunt in libro vitae.
PHIL|4|4|Gaudete in Domino semper. Iterum dico: Gaudete!
PHIL|4|5|Modestia vestra nota sit omnibus hominibus. Dominus prope.
PHIL|4|6|Nihil solliciti sitis, sed in omnibus oratione et obsecratione cum gratiarum actione petitiones vestrae innotescant apud Deum.
PHIL|4|7|Et pax Dei, quae exsuperat omnem sensum, custodiet corda vestra et intellegentias vestras in Christo Iesu.
PHIL|4|8|De cetero, fratres, quaecumque sunt vera, quaecumque pudica, quaecumque iusta, quaecumque casta, quaecumque amabilia, quaecumque bonae famae, si qua virtus et si qua laus, haec cogitate;
PHIL|4|9|quae et didicistis et accepistis et audistis et vidistis in me, haec agite; et Deus pacis erit vobiscum.
PHIL|4|10|Gavisus sum autem in Domino vehementer, quoniam tandem aliquando refloruistis pro me sentire, sicut et sentiebatis, opportunitate autem carebatis.
PHIL|4|11|Non quasi propter penuriam dico, ego enim didici, in quibus sum, sufficiens esse.
PHIL|4|12|Scio et humiliari, scio et abundare; ubique et in omnibus institutus sum et satiari et esurire et abundare et penuriam pati.
PHIL|4|13|Omnia possum in eo, qui me confortat.
PHIL|4|14|Verumtamen bene fecistis communicantes tribulationi meae.
PHIL|4|15|Scitis autem et vos, Philippenses, quod in principio evangelii, quando profectus sum a Macedonia, nulla mihi ecclesia communicavit in ratione dati et accepti, nisi vos soli;
PHIL|4|16|quia et Thessalonicam et semel et bis in usum mihi misistis.
PHIL|4|17|Non quia quaero datum, sed requiro fructum, qui abundet in rationem vestram.
PHIL|4|18|Accepi autem omnia et abundo; repletus sum acceptis ab Epaphrodito, quae misistis odorem suavitatis, hostiam acceptam, placentem Deo.
PHIL|4|19|Deus autem meus implebit omne desiderium vestrum secundum divitias suas in gloria in Christo Iesu.
PHIL|4|20|Deo autem et Patri nostro gloria in saecula saeculorum. Amen.
PHIL|4|21|Salutate omnem sanctum in Christo Iesu. Salutant vos, qui mecum sunt, fratres.
PHIL|4|22|Salutant vos omnes sancti, maxime autem, qui de Caesaris domo sunt.
PHIL|4|23|Gratia Domini Iesu Christi cum spiritu vestro. Amen.
COL|1|1|Paulus, apostolus Christi Iesu per voluntatem Dei, et Timo theus frater
COL|1|2|his, qui sunt Colossis, sanctis et fidelibus fratribus in Christo: gratia vobis et pax a Deo Patre nostro.
COL|1|3|Gratias agimus Deo Patri Domini nostri Iesu Christi semper pro vobis orantes,
COL|1|4|audientes fidem vestram in Christo Iesu et dilectionem, quam habetis in sanctos omnes,
COL|1|5|propter spem, quae reposita est vobis in caelis, quam ante audistis in verbo veritatis evangelii,
COL|1|6|quod pervenit ad vos, sicut et in universo mundo est fructificans et crescens, sicut et in vobis, ex ea die, qua audistis et cognovistis gratiam Dei in veritate;
COL|1|7|sicut didicistis ab Epaphra carissimo conservo nostro, qui est fidelis pro nobis minister Christi,
COL|1|8|qui etiam manifestavit nobis dilectionem vestram in Spiritu.
COL|1|9|Ideo et nos, ex qua die audivimus, non cessamus pro vobis orantes et postulantes, ut impleamini agnitione voluntatis eius in omni sapientia et intellectu spiritali,
COL|1|10|ut ambuletis digne Domino per omnia placentes, in omni opere bono fructificantes et crescentes in scientia Dei,
COL|1|11|in omni virtute confortati secundum potentiam claritatis eius in omnem patientiam et longanimitatem, cum gaudio
COL|1|12|gratias agentes Patri,qui idoneos vos fecit in partem sortis sanctorum in lumine;
COL|1|13|qui eripuit nos de potestate tenebrarumet transtulit in regnum Filii dilectionis suae,
COL|1|14|in quo habemus redemptionem,remissionem peccatorum;
COL|1|15|qui est imago Dei invisibilis,primogenitus omnis creaturae,
COL|1|16|quia in ipso condita sunt universa in caelis et in terra,visibilia et invisibilia,sive throni sive dominationessive principatus sive potestates.Omnia per ipsum et in ipsum creata sunt,
COL|1|17|et ipse est ante omnia,et omnia in ipso constant.
COL|1|18|Et ipse est caput corporis ecclesiae;qui est principium, primogenitus ex mortuis,ut sit in omnibus ipse primatum tenens,
COL|1|19|quia in ipso complacuit omnem plenitudinem habitare
COL|1|20|et per eum reconciliare omnia in ipsum,pacificans per sanguinem crucis eius,sive quae in terris sive quae in caelis sunt.
COL|1|21|Et vos, cum essetis aliquando alienati et inimici sensu in operibus malis,
COL|1|22|nunc autem reconciliavit in corpore carnis eius per mortem exhibere vos sanctos et immaculatos et irreprehensibiles coram ipso;
COL|1|23|si tamen permanetis in fide fundati et stabiles et immobiles a spe evangelii, quod audistis, quod praedicatum est in universa creatura, quae sub caelo est, cuius factus sum ego Paulus minister.
COL|1|24|Nunc gaudeo in passionibus pro vobis et adimpleo, ea quae desunt passionum Christi in carne mea pro corpore eius, quod est ecclesia,
COL|1|25|cuius factus sum ego minister secundum dispensationem Dei, quae data est mihi in vos, ut impleam verbum Dei;
COL|1|26|mysterium, quod absconditum fuit a saeculis et generationibus, nunc autem manifestatum est sanctis eius,
COL|1|27|quibus voluit Deus notas facere divitias gloriae mysterii huius in gentibus, quod est Christus in vobis, spes gloriae;
COL|1|28|quem nos annuntiamus, commonentes omnem hominem et docentes omnem hominem in omni sapientia, ut exhibeamus omnem hominem perfectum in Christo;
COL|1|29|ad quod et laboro certando secundum operationem eius, quae operatur in me in virtute.
COL|2|1|Volo enim vos scire qualem sollicitudinem habeam pro vo bis et pro his, qui sunt Laodiciae, et quicumque non viderunt faciem meam in carne,
COL|2|2|ut consolentur corda ipsorum instructi in caritate et in omnes divitias plenitudinis intellectus, in agnitionem mysterii Dei, Christi,
COL|2|3|in quo sunt omnes thesauri sapientiae et scientiae absconditi.
COL|2|4|Hoc dico, ut nemo vos decipiat in subtilitate sermonum.
COL|2|5|Nam etsi corpore absens sum, sed spiritu vobiscum sum, gaudens et videns ordinem vestrum et firmamentum eius, quae in Christum est, fidei vestrae.
COL|2|6|Sicut ergo accepistis Christum Iesum Dominum, in ipso ambulate,
COL|2|7|radicati et superaedificati in ipso et confirmati fide, sicut didicistis, abundantes in gratiarum actione.
COL|2|8|Videte, ne quis vos depraedetur per philosophiam et inanem fallaciam secundum traditionem hominum, secundum elementa mundi et non secundum Christum;
COL|2|9|quia in ipso inhabitat omnis plenitudo divinitatis corporaliter,
COL|2|10|et estis in illo repleti, qui est caput omnis principatus et potestatis;
COL|2|11|in quo et circumcisi estis circumcisione non manufacta in exspoliatione corporis carnis, in circumcisione Christi;
COL|2|12|consepulti ei in baptismo, in quo et conresuscitati estis per fidem operationis Dei, qui suscitavit illum a mortuis;
COL|2|13|et vos, cum mortui essetis in delictis et praeputio carnis vestrae, convivificavit cum illo, donans nobis omnia delicta,
COL|2|14|delens, quod adversum nos erat, chirographum decretis, quod erat contrarium nobis, et ipsum tulit de medio affigens illud cruci;
COL|2|15|exspolians principatus et potestates traduxit confidenter, triumphans illos in semetipso.
COL|2|16|Nemo ergo vos iudicet in cibo aut in potu aut ex parte diei festi aut neomeniae aut sabbatorum,
COL|2|17|quae sunt umbra futurorum, corpus autem Christi.
COL|2|18|Nemo vos bravio defraudet complacens sibi in humilitate et religione angelorum propter ea, quae vidit, ingrediens, frustra inflatus sensu carnis suae
COL|2|19|et non tenens caput, ex quo totum corpus per nexus et coniunctiones subministratum et compaginatum crescit in augmentum Dei.
COL|2|20|Si mortui estis cum Christo ab elementis mundi, quid tamquam viventes in mundo decretis subicimini:
COL|2|21|" Ne tetigeris neque gustaveris neque contrectaveris ",
COL|2|22|quae sunt omnia in corruptionem ipso usu secundum praecepta et doctrinas hominum?
COL|2|23|Quae sunt rationem quidem habentia sapientiae in superstitione et humilitate, et non parcendo corpori, non in honore aliquo ad saturitatem carnis.
COL|3|1|Igitur, si conresurrexistis Chri sto, quae sursum sunt quaerite, ubi Christus est in dextera Dei sedens;
COL|3|2|quae sursum sunt sapite, non quae supra terram.
COL|3|3|Mortui enim estis, et vita vestra abscondita est cum Christo in Deo!
COL|3|4|Cum Christus apparuerit, vita vestra, tunc et vos apparebitis cum ipso in gloria.
COL|3|5|Mortificate ergo membra, quae sunt super terram: fornicationem, immunditiam, libidinem, concupiscentiam malam et avaritiam, quae est simulacrorum servitus,
COL|3|6|propter quae venit ira Dei super filios incredulitatis;
COL|3|7|in quibus et vos ambulastis aliquando, cum viveretis in illis.
COL|3|8|Nunc autem deponite et vos omnia: iram, indignationem, malitiam, blasphemiam, turpem sermonem de ore vestro;
COL|3|9|nolite mentiri invicem, qui exuistis vos veterem hominem cum actibus eius
COL|3|10|et induistis novum, eum, qui renovatur in agnitionem secundum imaginem eius, qui creavit eum,
COL|3|11|ubi non est Graecus et Iudaeus, circumcisio et praeputium, barbarus, Scytha, servus, liber, sed omnia et in omnibus Christus.
COL|3|12|Induite vos ergo, sicut electi Dei, sancti et dilecti, viscera misericordiae, benignitatem, humilitatem, mansuetudinem, longanimitatem,
COL|3|13|supportantes invicem et donantes vobis ipsis, si quis adversus aliquem habet querelam; sicut et Dominus donavit vobis, ita et vos;
COL|3|14|super omnia autem haec: caritatem, quod est vinculum perfectionis.
COL|3|15|Et pax Christi dominetur in cordibus vestris, ad quam et vocati estis in uno corpore. Et grati estote.
COL|3|16|Verbum Christi habitet in vobis abundanter, in omni sapientia docentes et commonentes vosmetipsos psalmis, hymnis, canticis spiritalibus, in gratia cantantes in cordibus vestris Deo;
COL|3|17|et omne, quodcumque facitis in verbo aut in opere, omnia in nomine Domini Iesu gratias agentes Deo Patri per ipsum.
COL|3|18|Mulieres, subditae estote viris, sicut oportet in Domino.
COL|3|19|Viri, diligite uxores et nolite amari esse ad illas.
COL|3|20|Filii, oboedite parentibus per omnia; hoc enim placitum est in Domino.
COL|3|21|Patres, nolite ad indignationem provocare filios vestros, ut non pusillo animo fiant.
COL|3|22|Servi, oboedite per omnia dominis carnalibus, non ad oculum servientes, quasi hominibus placentes, sed in simplicitate cordis, timentes Dominum.
COL|3|23|Quodcumque facitis, ex animo operamini sicut Domino et non hominibus,
COL|3|24|scientes quod a Domino accipietis retributionem hereditatis. Domino Christo servite;
COL|3|25|qui enim iniuriam facit, recipiet id quod inique gessit, et non est personarum acceptio.
COL|4|1|Domini, quod iustum est et aequum, servis praestate, scien tes quoniam et vos Dominum habetis in caelo.
COL|4|2|Orationi instate, vigilantes in ea in gratiarum actione,
COL|4|3|orantes simul et pro nobis, ut Deus aperiat nobis ostium sermonis ad loquendum mysterium Christi, propter quod etiam vinctus sum,
COL|4|4|ut manifestem illud, ita ut oportet me loqui.
COL|4|5|In sapientia ambulate ad eos, qui foris sunt, tempus redimentes.
COL|4|6|Sermo vester semper sit in gratia, sale conditus, ut sciatis quomodo oporteat vos unicuique respondere.
COL|4|7|Quae circa me sunt, omnia vobis nota faciet Tychicus, carissimus frater et fidelis minister et conservus in Domino,
COL|4|8|quem misi ad vos ad hoc ipsum, ut cognoscatis, quae circa nos sunt, et consoletur corda vestra,
COL|4|9|cum Onesimo fideli et carissimo fratre, qui est ex vobis; omnia, quae hic aguntur, nota facient vobis.
COL|4|10|Salutat vos Aristarchus concaptivus meus et Marcus consobrinus Barnabae, de quo accepistis mandata - si venerit ad vos, excipite illum -
COL|4|11|et Iesus, qui dicitur Iustus, qui sunt ex circumcisione; hi soli adiutores in regno Dei, qui mihi fuerunt solacio.
COL|4|12|Salutat vos Epaphras, qui ex vobis est, servus Christi Iesu, semper certans pro vobis in orationibus, ut stetis perfecti et impleti in omni voluntate Dei.
COL|4|13|Testimonium enim illi perhibeo, quod habet multum laborem pro vobis et pro his, qui sunt Laodiciae et qui Hierapoli.
COL|4|14|Salutat vos Lucas, medicus carissimus, et Demas.
COL|4|15|Salutate fratres, qui sunt Laodiciae, et Nympham et, quae in domo eius est, ecclesiam.
COL|4|16|Et cum lecta fuerit apud vos epistula, facite ut et in Laodicensium ecclesia legatur, et eam, quae ex Laodicia est, vos quoque legatis.
COL|4|17|Et dicite Archippo: " Vide ministerium, quod accepisti in Domino, ut illud impleas ".
COL|4|18|Salutatio mea manu Pauli. Memores estote vinculorum meorum.Gratia vobiscum.
1THESS|1|1|Paulus et Silvanus et Timo theus ecclesiae Thessalonicen sium in Deo Patre et Domino Iesu Christo: gratia vobis et pax.
1THESS|1|2|Gratias agimus Deo semper pro omnibus vobis, memoriam facientes in orationibus nostris, sine intermissione;
1THESS|1|3|memores operis fidei vestrae et laboris caritatis et sustinentiae spei Domini nostri Iesu Christi ante Deum et Patrem nostrum;
1THESS|1|4|scientes, fratres, dilecti a Deo, electionem vestram,
1THESS|1|5|quia evangelium nostrum non fuit ad vos in sermone tantum sed et in virtute et in Spiritu Sancto et in plenitudine multa, sicut scitis quales fuerimus vobis propter vos.
1THESS|1|6|Et vos imitatores nostri facti estis et Domini, excipientes verbum in tribulatione multa cum gaudio Spiritus Sancti,
1THESS|1|7|ita ut facti sitis forma omnibus credentibus in Macedonia et in Achaia.
1THESS|1|8|A vobis enim diffamatus est sermo Domini non solum in Macedonia et in Achaia, sed in omni loco fides vestra, quae est ad Deum, profecta est, ita ut non sit nobis necesse quidquam loqui;
1THESS|1|9|ipsi enim de nobis annuntiant qualem introitum habuerimus ad vos, et quomodo conversi estis ad Deum a simulacris, servire Deo vivo et vero
1THESS|1|10|et exspectare Filium eius de caelis, quem suscitavit ex mortuis, Iesum, qui eripit nos ab ira ventura.
1THESS|2|1|Nam ipsi scitis, fratres, introi tum nostrum ad vos, quia non inanis fuit;
1THESS|2|2|sed ante passi et contumeliis affecti, sicut scitis, in Philippis, fiduciam habuimus in Deo nostro loqui ad vos evangelium Dei in multa sollicitudine.
1THESS|2|3|Exhortatio enim nostra non ex errore neque ex immunditia neque in dolo,
1THESS|2|4|sed sicut probati sumus a Deo, ut crederetur nobis evangelium, ita loquimur non quasi hominibus placentes, sed Deo, qui probat corda nostra.
1THESS|2|5|Neque enim aliquando fuimus in sermone adulationis, sicut scitis, neque sub praetextu avaritiae, Deus testis,
1THESS|2|6|nec quaerentes ab hominibus gloriam, neque a vobis neque ab aliis;
1THESS|2|7|cum possemus oneri esse ut Christi apostoli, sed facti sumus parvuli in medio vestrum, tamquam si nutrix foveat filios suos;
1THESS|2|8|ita desiderantes vos, cupide volebamus tradere vobis non solum evangelium Dei sed etiam animas nostras, quoniam carissimi nobis facti estis.
1THESS|2|9|Memores enim estis, fratres, laboris nostri et fatigationis; nocte et die operantes, ne quem vestrum gravaremus, praedicavimus in vobis evangelium Dei.
1THESS|2|10|Vos testes estis et Deus, quam sancte et iuste et sine querela vobis, qui credidistis, fuimus;
1THESS|2|11|sicut scitis qualiter unumquemque vestrum, tamquam pater filios suos,
1THESS|2|12|deprecantes vos et consolantes testificati sumus, ut ambularetis digne Deo, qui vocat vos in suum regnum et gloriam.
1THESS|2|13|Ideo et nos gratias agimus Deo sine intermissione, quoniam cum accepissetis a nobis verbum auditus Dei, accepistis non ut verbum hominum sed, sicut est vere, verbum Dei, quod et operatur in vobis, qui creditis.
1THESS|2|14|Vos enim imitatores facti estis, fratres, ecclesiarum Dei, quae sunt in Iudaea in Christo Iesu; quia eadem passi estis et vos a contribulibus vestris, sicut et ipsi a Iudaeis,
1THESS|2|15|qui et Dominum occiderunt Iesum et prophetas et nos persecuti sunt et Deo non placent et omnibus hominibus adversantur,
1THESS|2|16|prohibentes nos gentibus loqui, ut salvae fiant, ut impleant peccata sua semper. Pervenit autem ira Dei super illos usque in finem.
1THESS|2|17|Nos autem, fratres, desolati a vobis ad tempus horae, facie non corde, abundantius festinavimus faciem vestram videre cum multo desiderio.
1THESS|2|18|Propter quod voluimus venire ad vos, ego quidem Paulus et semel et iterum; et impedivit nos Satanas.
1THESS|2|19|Quae est enim nostra spes aut gaudium aut corona gloriae - nonne et vos ante Dominum nostrum Iesum in adventu eius?
1THESS|2|20|Vos enim estis gloria nostra et gaudium.
1THESS|3|1|Propter quod non sustinentes amplius, placuit nobis, ut relin queremur Athenis soli,
1THESS|3|2|et misimus Timotheum, fratrem nostrum et cooperatorem Dei in evangelio Christi, ad confirmandos vos et exhortandos pro fide vestra,
1THESS|3|3|ut nemo turbetur in tribulationibus istis. Ipsi enim scitis quod in hoc positi sumus;
1THESS|3|4|nam et cum apud vos essemus, praedicebamus vobis passuros nos tribulationes, sicut et factum est et scitis.
1THESS|3|5|Propterea et ego amplius non sustinens, misi ad cognoscendam fidem vestram, ne forte tentaverit vos is qui tentat, et inanis fiat labor noster.
1THESS|3|6|Nunc autem, veniente Timotheo ad nos a vobis et annuntiante nobis fidem et caritatem vestram, et quia memoriam nostri habetis bonam semper, desiderantes nos videre, sicut nos quoque vos;
1THESS|3|7|ideo consolati sumus, fratres, propter vos in omni necessitate et tribulatione nostra per vestram fidem;
1THESS|3|8|quoniam nunc vivimus, si vos statis in Domino.
1THESS|3|9|Quam enim gratiarum actionem possumus Deo retribuere pro vobis in omni gaudio, quo gaudemus propter vos ante Deum nostrum,
1THESS|3|10|nocte et die abundantius orantes, ut videamus faciem vestram et compleamus ea, quae desunt fidei vestrae?
1THESS|3|11|Ipse autem Deus et Pater noster et Dominus noster Iesus dirigat viam nostram ad vos;
1THESS|3|12|vos autem Dominus abundare et superabundare faciat caritate in invicem et in omnes, quemadmodum et nos in vos;
1THESS|3|13|ad confirmanda corda vestra sine querela in sanctitate ante Deum et Patrem nostrum, in adventu Domini nostri Iesu cum omnibus sanctis eius. Amen.
1THESS|4|1|De cetero ergo, fratres, rogamus vos et obsecramus in Domino Iesu, ut - quemadmodum accepistis a nobis quomodo vos oporteat ambulare et placere Deo, sicut et ambulatis - ut abundetis magis.
1THESS|4|2|Scitis enim, quae praecepta dederimus vobis per Dominum Iesum.
1THESS|4|3|Haec est enim voluntas Dei, sanctificatio vestra,
1THESS|4|4|ut abstineatis a fornicatione; ut sciat unusquisque vestrum suum vas possidere in sanctificatione et honore,
1THESS|4|5|non in passione desiderii, sicut et gentes, quae ignorant Deum;
1THESS|4|6|ut ne quis supergrediatur neque circumveniat in negotio fratrem suum, quoniam vindex est Dominus de his omnibus, sicut et praediximus vobis et testificati sumus.
1THESS|4|7|Non enim vocavit nos Deus in immunditiam sed in sanctificationem.
1THESS|4|8|Itaque, qui spernit, non hominem spernit sed Deum, qui etiam dat Spiritum suum Sanctum in vos.
1THESS|4|9|De caritate autem fraternitatis non necesse habetis, ut vobis scribam; ipsi enim vos a Deo edocti estis, ut diligatis invicem;
1THESS|4|10|etenim facitis illud in omnes fratres in universa Macedonia. Rogamus autem vos, fratres, ut abundetis magis;
1THESS|4|11|et operam detis, ut quieti sitis et ut vestrum negotium agatis et operemini manibus vestris, sicut praecipimus vobis;
1THESS|4|12|ut honeste ambuletis ad eos, qui foris sunt, et nullius aliquid desideretis.
1THESS|4|13|Nolumus autem vos ignorare, fratres, de dormientibus, ut non contristemini sicut et ceteri, qui spem non habent.
1THESS|4|14|Si enim credimus quod Iesus mortuus est et resurrexit, ita et Deus eos, qui dormierunt, per Iesum adducet cum eo.
1THESS|4|15|Hoc enim vobis dicimus in verbo Domini, quia nos, qui vivimus, qui relinquimur in adventum Domini, non praeveniemus eos, qui dormierunt;
1THESS|4|16|quoniam ipse Dominus in iussu, in voce archangeli et in tuba Dei descendet de caelo, et mortui, qui in Christo sunt, resurgent primi;
1THESS|4|17|deinde nos, qui vivimus, qui relinquimur, simul rapiemur cum illis in nubibus obviam Domino in aera, et sic semper cum Domino erimus.
1THESS|4|18|Itaque consolamini invicem in verbis istis.
1THESS|5|1|De temporibus autem et mo mentis, fratres, non indigetis, ut scribatur vobis;
1THESS|5|2|ipsi enim diligenter scitis quia dies Domini, sicut fur in nocte, ita veniet.
1THESS|5|3|Cum enim dixerint: " Pax et securitas ", tunc repentinus eis superveniet interitus, sicut dolor in utero habenti, et non effugient.
1THESS|5|4|Vos autem, fratres, non estis in tenebris, ut vos dies ille tamquam fur comprehendat;
1THESS|5|5|omnes enim vos filii lucis estis et filii diei. Non sumus noctis neque tenebrarum;
1THESS|5|6|igitur non dormiamus sicut ceteri, sed vigilemus et sobrii simus.
1THESS|5|7|Qui enim dormiunt, nocte dormiunt; et, qui ebrii sunt, nocte inebriantur.
1THESS|5|8|Nos autem, qui diei sumus, sobrii simus, induti loricam fidei et caritatis et galeam spem salutis;
1THESS|5|9|quoniam non posuit nos Deus in iram sed in acquisitionem salutis per Dominum nostrum Iesum Christum,
1THESS|5|10|qui mortuus est pro nobis, ut sive vigilemus sive dormiamus, simul cum illo vivamus.
1THESS|5|11|Propter quod consolamini invicem et aedificate alterutrum, sicut et facitis.
1THESS|5|12|Rogamus autem vos, fratres, ut noveritis eos, qui laborant inter vos et praesunt vobis in Domino et monent vos,
1THESS|5|13|ut habeatis illos superabundanter in caritate propter opus illorum. Pacem habete inter vos.
1THESS|5|14|Hortamur autem vos, fratres: corripite inquietos, consolamini pusillanimes, suscipite infirmos, longanimes estote ad omnes.
1THESS|5|15|Videte, ne quis malum pro malo alicui reddat, sed semper, quod bonum est, sectamini et in invicem et in omnes.
1THESS|5|16|Semper gaudete,
1THESS|5|17|sine intermissione orate,
1THESS|5|18|in omnibus gratias agite; haec enim voluntas Dei est in Christo Iesu erga vos.
1THESS|5|19|Spiritum nolite exstinguere,
1THESS|5|20|prophetias nolite spernere;
1THESS|5|21|omnia autem probate, quod bonum est tenete,
1THESS|5|22|ab omni specie mala abstinete vos.
1THESS|5|23|Ipse autem Deus pacis sanctificet vos per omnia, et integer spiritus vester et anima et corpus sine querela in adventu Domini nostri Iesu Christi servetur.
1THESS|5|24|Fidelis est, qui vocat vos, qui etiam faciet.
1THESS|5|25|Fratres, orate etiam pro nobis.
1THESS|5|26|Salutate fratres omnes in osculo sancto.
1THESS|5|27|Adiuro vos per Dominum, ut legatur epistula omnibus fratribus.
1THESS|5|28|Gratia Domini nostri Iesu Christi vobiscum.
2THESS|1|1|Paulus et Silvanus et Timo theus ecclesiae Thessalonicen sium in Deo Patre nostro et Domino Iesu Christo:
2THESS|1|2|gratia vobis et pax a Deo Patre nostro et Domino Iesu Christo.
2THESS|1|3|Gratias agere debemus Deo semper pro vobis, fratres, sicut dignum est, quoniam supercrescit fides vestra, et abundat caritas uniuscuiusque omnium vestrum in invicem,
2THESS|1|4|ita ut et nos ipsi in vobis gloriemur in ecclesiis Dei pro patientia vestra et fide in omnibus persecutionibus vestris et tribulationibus, quas sustinetis,
2THESS|1|5|indicium iusti iudicii Dei, ut digni habeamini regno Dei, pro quo et patimini;
2THESS|1|6|si quidem iustum est apud Deum retribuere tribulationem his, qui vos tribulant,
2THESS|1|7|et vobis, qui tribulamini, requiem nobiscum in revelatione Domini Iesu de caelo cum angelis virtutis eius,
2THESS|1|8|in igne flammae, dantis vindictam his, qui non noverunt Deum et qui non oboediunt evangelio Domini nostri Iesu;
2THESS|1|9|qui poenas dabunt interitu aeterno a facie Domini et a gloria virtutis eius,
2THESS|1|10|cum venerit glorificari in sanctis suis et admirabilis fieri in omnibus, qui crediderunt; quia creditum est testimonium nostrum super vos in die illo.
2THESS|1|11|Ad quod etiam oramus semper pro vobis, ut dignetur vos vocatione sua Deus noster et impleat omnem voluntatem bonitatis et opus fidei in virtute;
2THESS|1|12|ut glorificetur nomen Domini nostri Iesu Christi in vobis, et vos in illo, secundum gratiam Dei nostri et Domini Iesu Christi.
2THESS|2|1|Rogamus autem vos, fratres, circa adventum Domini nostri Iesu Christi et nostram congregationem in ipsum,
2THESS|2|2|ut non cito moveamini a sensu neque terreamini, neque per spiritum neque per verbum neque per epistulam tamquam per nos, quasi instet dies Domini.
2THESS|2|3|Ne quis vos seducat ullo modo; quoniam, nisi venerit discessio primum, et revelatus fuerit homo iniquitatis, filius perditionis,
2THESS|2|4|qui adversatur et extollitur supra omne, quod dicitur Deus aut quod colitur, ita ut in templo Dei sedeat, ostendens se quia sit Deus.
2THESS|2|5|Non retinetis quod, cum adhuc essem apud vos, haec dicebam vobis?
2THESS|2|6|Et nunc quid detineat scitis, ut ipse reveletur in suo tempore.
2THESS|2|7|Nam mysterium iam operatur iniquitatis; tantum qui tenet nunc, donec de medio fiat.
2THESS|2|8|Et tunc revelabitur ille iniquus, quem Dominus Iesus interficiet spiritu oris sui et destruet illustratione adventus sui,
2THESS|2|9|eum, cuius est adventus secundum operationem Satanae in omni virtute et signis et prodigiis mendacibus
2THESS|2|10|et in omni seductione iniquitatis his, qui pereunt, eo quod caritatem veritatis non receperunt, ut salvi fierent.
2THESS|2|11|Et ideo mittit illis Deus operationem erroris, ut credant mendacio,
2THESS|2|12|ut iudicentur omnes, qui non crediderunt veritati, sed consenserunt iniquitati.
2THESS|2|13|Nos autem debemus gratias agere Deo semper pro vobis, fratres, dilecti a Domino, quod elegerit vos Deus primitias in salutem, in sanctificatione Spiritus et fide veritatis;
2THESS|2|14|ad quod et vocavit vos per evangelium nostrum in acquisitionem gloriae Domini nostri Iesu Christi.
2THESS|2|15|Itaque, fratres, state et tenete traditiones, quas didicistis sive per sermonem sive per epistulam nostram.
2THESS|2|16|Ipse autem Dominus noster Iesus Christus et Deus Pater noster, qui dilexit nos et dedit consolationem aeternam et spem bonam in gratia,
2THESS|2|17|consoletur corda vestra et confirmet in omni opere et sermone bono.
2THESS|3|1|De cetero, fratres, orate pro nobis, ut sermo Domini currat et glorificetur sicut et apud vos,
2THESS|3|2|et ut liberemur ab importunis et malis hominibus; non enim omnium est fides.
2THESS|3|3|Fidelis autem Dominus est, qui confirmabit vos et custodiet a Malo.
2THESS|3|4|Confidimus autem de vobis in Domino, quoniam, quae praecipimus, et facitis et facietis.
2THESS|3|5|Dominus autem dirigat corda vestra in caritatem Dei et patientiam Christi.
2THESS|3|6|Praecipimus autem vobis, fratres, in nomine Domini nostri Iesu Christi, ut subtrahatis vos ab omni fratre ambulante inordinate et non secundum traditionem, quam acceperunt a nobis.
2THESS|3|7|Ipsi enim scitis quemadmodum oporteat imitari nos, quoniam non inordinati fuimus inter vos
2THESS|3|8|neque gratìs panem manducavimus ab aliquo sed in labore et fatigatione, nocte et die operantes, ne quem vestrum gravaremus;
2THESS|3|9|non quasi non habuerimus potestatem, sed ut nosmetipsos formam daremus vobis ad imitandum nos.
2THESS|3|10|Nam et cum essemus apud vos, hoc praecipiebamus vobis: Si quis non vult operari, nec manducet.
2THESS|3|11|Audimus enim inter vos quosdam ambulare inordinate, nihil operantes sed curiose agentes;
2THESS|3|12|his autem, qui eiusmodi sunt, praecipimus et obsecramus in Domino Iesu Christo, ut cum quiete operantes suum panem manducent.
2THESS|3|13|Vos autem, fratres, nolite deficere benefacientes.
2THESS|3|14|Quod si quis non oboedit verbo nostro per epistulam, hunc notate, non commisceamini cum illo, ut confundatur;
2THESS|3|15|et nolite quasi inimicum existimare, sed corripite ut fratrem.
2THESS|3|16|Ipse autem Dominus pacis det vobis pacem sempiternam in omni modo. Dominus cum omnibus vobis.
2THESS|3|17|Salutatio mea manu Pauli, quod est signum in omni epistula; ita scribo.
2THESS|3|18|Gratia Domini nostri Iesu Christi cum omnibus vobis.
1TIM|1|1|Paulus, apostolus Christi Iesu secundum praeceptum Dei sal vatoris nostri et Christi Iesu spei nostrae,
1TIM|1|2|Timotheo germano filio in fide: gratia, misericordia, pax a Deo Patre et Christo Iesu Domino nostro.
1TIM|1|3|Sicut rogavi te, ut remaneres Ephesi, cum irem in Macedoniam, ut praeciperes quibusdam, ne aliter docerent
1TIM|1|4|neque intenderent fabulis et genealogiis interminatis, quae quaestiones praestant magis quam dispensationem Dei, quae est in fide;
1TIM|1|5|finis autem praecepti est caritas de corde puro et conscientia bona et fide non ficta,
1TIM|1|6|a quibus quidam aberrantes conversi sunt in vaniloquium,
1TIM|1|7|volentes esse legis doctores, non intellegentes neque quae loquuntur neque de quibus affirmant.
1TIM|1|8|Scimus autem quia bona est lex, si quis ea legitime utatur,
1TIM|1|9|sciens hoc quia iusto lex non est posita sed iniustis et non subiectis, impiis et peccatoribus, sceleratis et contaminatis, patricidis et matricidis, homicidis,
1TIM|1|10|fornicariis, masculorum concubitoribus, plagiariis, mendacibus, periuris et si quid aliud sanae doctrinae adversatur,
1TIM|1|11|secundum evangelium gloriae beati Dei, quod creditum est mihi.
1TIM|1|12|Gratiam habeo ei, qui me confortavit, Christo Iesu Domino nostro, quia fidelem me existimavit ponens in ministerio,
1TIM|1|13|qui prius fui blasphemus et persecutor et contumeliosus; sed misericordiam consecutus sum, quia ignorans feci in incredulitate;
1TIM|1|14|superabundavit autem gratia Domini nostri cum fide et dilectione, quae sunt in Christo Iesu.
1TIM|1|15|Fidelis sermo et omni acceptione dignus: Christus Iesus venit in mundum peccatores salvos facere; quorum primus ego sum,
1TIM|1|16|sed ideo misericordiam consecutus sum, ut in me primo ostenderet Christus Iesus omnem longanimitatem, ad informationem eorum, qui credituri sunt illi in vitam aeternam.
1TIM|1|17|Regi autem saeculorum, incorruptibili, invisibili, soli Deo honor et gloria in saecula saeculorum. Amen.
1TIM|1|18|Hoc praeceptum commendo tibi, fili Timothee, secundum praecedentes super te prophetias, ut milites in illis bonam militiam
1TIM|1|19|habens fidem et bonam conscientiam, quam quidam repellentes circa fidem naufragaverunt;
1TIM|1|20|ex quibus est Hymenaeus et Alexander, quos tradidi Satanae, ut discant non blasphemare.
1TIM|2|1|Obsecro igitur primo omnium fieri obsecrationes, orationes, postulationes, gratiarum actiones pro omnibus hominibus,
1TIM|2|2|pro regibus et omnibus, qui in sublimitate sunt, ut quietam et tranquillam vitam agamus in omni pietate et castitate.
1TIM|2|3|Hoc bonum est et acceptum coram salvatore nostro Deo,
1TIM|2|4|qui omnes homines vult salvos fieri et ad agnitionem veritatis venire.
1TIM|2|5|Unus enim Deus, unus et mediator Dei et hominum, homo Christus Iesus,
1TIM|2|6|qui dedit redemptionem semetipsum pro omnibus, testimonium temporibus suis;
1TIM|2|7|in quod positus sum ego praedicator et apostolus - veritatem dico, non mentior - doctor gentium in fide et veritate.
1TIM|2|8|Volo ergo viros orare in omni loco levantes puras manus sine ira et disceptatione;
1TIM|2|9|similiter et mulieres in habitu ornato cum verecundia et sobrietate ornantes se, non in tortis crinibus et auro aut margaritis vel veste pretiosa,
1TIM|2|10|sed, quod decet mulieres, profitentes pietatem per opera bona.
1TIM|2|11|Mulier in tranquillitate discat cum omni subiectione;
1TIM|2|12|docere autem mulieri non permitto neque dominari in virum, sed esse in tranquillitate.
1TIM|2|13|Adam enim primus formatus est, deinde Eva;
1TIM|2|14|et Adam non est seductus, mulier autem seducta in praevaricatione fuit.
1TIM|2|15|Salvabitur autem per filiorum generationem, si permanserint in fide et dilectione et sanctificatione cum sobrietate.
1TIM|3|1|Fidelis sermo: si quis episco patum appetit, bonum opus de siderat.
1TIM|3|2|Oportet ergo episcopum irreprehensibilem esse, unius uxoris virum, sobrium, prudentem, ornatum, hospitalem, doctorem,
1TIM|3|3|non vinolentum, non percussorem sed modestum, non litigiosum, non cupidum,
1TIM|3|4|suae domui bene praepositum, filios habentem in subiectione cum omni castitate
1TIM|3|5|- si quis autem domui suae praeesse nescit, quomodo ecclesiae Dei curam habebit? C,
1TIM|3|6|non neophytum, ne in superbia elatus in iudicium incidat Diaboli.
1TIM|3|7|Oportet autem illum et testimonium habere bonum ab his, qui foris sunt, ut non in opprobrium incidat et laqueum Diaboli.
1TIM|3|8|Diaconos similiter pudicos, non bilingues, non multo vino deditos, non turpe lucrum sectantes,
1TIM|3|9|habentes mysterium fidei in conscientia pura.
1TIM|3|10|Et hi autem probentur primum, deinde ministrent nullum crimen habentes.
1TIM|3|11|Mulieres similiter pudicas, non detrahentes, sobrias, fideles in omnibus.
1TIM|3|12|Diaconi sint unius uxoris viri, qui filiis suis bene praesint et suis domibus;
1TIM|3|13|qui enim bene ministraverint, gradum sibi bonum acquirent et multam fiduciam in fide, quae est in Christo Iesu.
1TIM|3|14|Haec tibi scribo sperans venire ad te cito;
1TIM|3|15|si autem tardavero, ut scias quomodo oporteat in domo Dei conversari, quae est ecclesia Dei vivi, columna et firmamentum veritatis.
1TIM|3|16|Et omnium confessione magnum est pietatis mysterium:Qui manifestatus est in carne,iustificatus est in Spiritu,apparuit angelis,praedicatus est in gentibus,creditus est in mumdo,assumptus est in gloria.
1TIM|4|1|Spiritus autem manifeste dicit, quia in novissimis temporibus discedent quidam a fide, attendentes spiritibus seductoribus et doctrinis daemoniorum,
1TIM|4|2|in hypocrisi loquentium mendacium et cauteriatam habentium suam conscientiam,
1TIM|4|3|prohibentium nubere, abstinere a cibis, quos Deus creavit ad percipiendum cum gratiarum actione fidelibus et his, qui cognoverunt veritatem.
1TIM|4|4|Quia omnis creatura Dei bona, et nihil reiciendum, quod cum gratiarum actione percipitur;
1TIM|4|5|sanctificatur enim per verbum Dei et orationem.
1TIM|4|6|Haec proponens fratribus bonus eris minister Christi Iesu, enutritus verbis fidei et bonae doctrinae, quam assecutus es;
1TIM|4|7|profanas autem et aniles fabulas devita.Exerce teipsum ad pietatem;
1TIM|4|8|nam corporalis exercitatio ad modicum utilis est, pietas autem ad omnia utilis est promissionem habens vitae, quae nunc est, et futurae.
1TIM|4|9|Fidelis sermo et omni acceptione dignus:
1TIM|4|10|in hoc enim laboramus et certamus, quia sperantes sumus in Deum vivum, qui est salvator omnium hominum, maxime fidelium.
1TIM|4|11|Praecipe haec et doce.
1TIM|4|12|Nemo adulescentiam tuam contemnat; sed exemplum esto fidelium in verbo, in conversatione, in caritate, in fide, in castitate.
1TIM|4|13|Dum venio, attende lectioni, exhortationi, doctrinae.
1TIM|4|14|Noli neglegere donationem, quae in te est, quae data est tibi per prophetiam cum impositione manuum presbyterii.
1TIM|4|15|Haec meditare, in his esto, ut profectus tuus manifestus sit omnibus.
1TIM|4|16|Attende tibi et doctrinae; insta in illis; hoc enim faciens et teipsum salvum facies et eos, qui te audiunt.
1TIM|5|1|Seniorem ne increpaveris, sed obsecra ut patrem, iuvenes ut fratres,
1TIM|5|2|anus ut matres, iuvenculas ut sorores in omni castitate.
1TIM|5|3|Viduas honora, quae vere viduae sunt.
1TIM|5|4|Si qua autem vidua filios aut nepotes habet, discant primum domum suam pie regere et mutuam vicem reddere parentibus; hoc enim acceptum est coram Deo.
1TIM|5|5|Quae autem vere vidua est et desolata, sperat in Deum et instat obsecrationibus et orationibus nocte ac die;
1TIM|5|6|nam quae in deliciis est vivens, mortua est.
1TIM|5|7|Et haec praecipe, ut irreprehensibiles sint.
1TIM|5|8|Si quis autem suorum et maxime domesticorum curam non habet, fidem negavit et est infideli deterior.
1TIM|5|9|Vidua adscribatur non minus sexaginta annorum, quae fuerit unius viri uxor,
1TIM|5|10|in operibus bonis testimonium habens: si filios educavit, si hospitio recepit, si sanctorum pedes lavit, si tribulationem patientibus subministravit, si omne opus bonum subsecuta est.
1TIM|5|11|Adulescentiores autem viduas devita; cum enim luxuriatae fuerint adversus Christum, nubere volunt,
1TIM|5|12|habentes damnationem, quia primam fidem irritam fecerunt;
1TIM|5|13|simul autem et otiosae discunt circumire domos, non solum otiosae sed et verbosae et curiosae, loquentes quae non oportet.
1TIM|5|14|Volo ergo iuniores nubere, filios procreare, dominas domus esse, nullam occasionem dare adversario maledicti gratia;
1TIM|5|15|iam enim quaedam conversae sunt retro Satanam.
1TIM|5|16|Si qua fidelis habet viduas, subministret illis, et non gravetur ecclesia, ut his, quae vere viduae sunt, sufficiat.
1TIM|5|17|Qui bene praesunt presbyteri, duplici honore digni habeantur, maxime qui laborant in verbo et doctrina;
1TIM|5|18|dicit enim Scriptura: " Non infrenabis os bovi trituranti " et: " Dignus operarius mercede sua ".
1TIM|5|19|Adversus presbyterum accusationem noli recipere, nisi sub duobus vel tribus testibus.
1TIM|5|20|Peccantes coram omnibus argue, ut et ceteri timorem habeant.
1TIM|5|21|Testificor coram Deo et Christo Iesu et electis angelis, ut haec custodias sine praeiudicio nihil faciens in aliquam partem declinando.
1TIM|5|22|Manus cito nemini imposueris neque communicaveris peccatis alienis; teipsum castum custodi.
1TIM|5|23|Noli adhuc aquam bibere, sed vino modico utere propter stomachum et frequentes tuas infirmitates.
1TIM|5|24|Quorundam hominum peccata manifesta sunt praecedentia ad iudicium, quosdam autem et subsequuntur;
1TIM|5|25|similiter et facta bona manifesta sunt, et, quae aliter se habent, abscondi non possunt.
1TIM|6|1|Quicumque sunt sub iugo, servi dominos suos omni honore di gnos arbitrentur, ne nomen Dei et doctrina blasphemetur.
1TIM|6|2|Qui autem fideles habent dominos, non contemnant, quia fratres sunt, sed magis serviant, quia fideles sunt et dilecti, qui beneficii participes sunt. Haec doce et exhortare.
1TIM|6|3|Si quis aliter docet et non accedit sanis sermonibus Domini nostri Iesu Christi et ei, quae secundum pietatem est, doctrinae,
1TIM|6|4|superbus est, nihil sciens, sed languens circa quaestiones et pugnas verborum, ex quibus oriuntur invidiae, contentiones, blasphemiae, suspiciones malae,
1TIM|6|5|conflictationes hominum mente corruptorum et qui veritate privati sunt, existimantium quaestum esse pietatem.
1TIM|6|6|Est autem quaestus magnus pietas cum sufficientia.
1TIM|6|7|Nihil enim intulimus in mundum, quia nec auferre quid possumus;
1TIM|6|8|habentes autem alimenta et quibus tegamur, his contenti erimus.
1TIM|6|9|Nam qui volunt divites fieri, incidunt in tentationem et laqueum et desideria multa stulta et nociva, quae mergunt homines in interitum et perditionem;
1TIM|6|10|radix enim omnium malorum est cupiditas, quam quidam appetentes erraverunt a fide et inseruerunt se doloribus multis.
1TIM|6|11|Tu autem, o homo Dei, haec fuge; sectare vero iustitiam, pietatem, fidem, caritatem, patientiam, mansuetudinem.
1TIM|6|12|Certa bonum certamen fidei, apprehende vitam aeternam, ad quam vocatus es, et confessus es bonam confessionem coram multis testibus.
1TIM|6|13|Praecipio tibi coram Deo, qui vivificat omnia, et Christo Iesu, qui testimonium reddidit sub Pontio Pilato bonam confessionem,
1TIM|6|14|ut serves mandatum sine macula irreprehensibile usque in adventum Domini nostri Iesu Christi,
1TIM|6|15|quem suis temporibus ostendet beatus et solus potens, Rex regnantium et Dominus dominantium,
1TIM|6|16|qui solus habet immortalitatem, lucem habitans inaccessibilem, quem vidit nullus hominum nec videre potest; cui honor et imperium sempiternum. Amen.
1TIM|6|17|Divitibus huius saeculi praecipe non superbe sapere neque sperare in incerto divitiarum sed in Deo, qui praestat nobis omnia abunde ad fruendum,
1TIM|6|18|bene agere, divites fieri in operibus bonis, facile tribuere, communicare,
1TIM|6|19|thesaurizare sibi fundamentum bonum in futurum, ut apprehendant veram vitam.
1TIM|6|20|O Timothee, depositum custodi, devitans profanas vocum novitates et oppositiones falsi nominis scientiae,
1TIM|6|21|quam quidam profitentes circa fidem aberraverunt.Gratia vobiscum.
2TIM|1|1|Paulus, apostolus Christi Iesu per voluntatem Dei secundum promissionem vitae, quae est in Christo Iesu,
2TIM|1|2|Timotheo carissimo filio: gratia, misericordia, pax a Deo Patre et Christo Iesu Domino nostro.
2TIM|1|3|Gratias ago Deo, cui servio a progenitoribus in conscientia pura, quod sine intermissione habeo tui memoriam in orationibus meis nocte ac die
2TIM|1|4|desiderans te videre, memor lacrimarum tuarum, ut gaudio implear,
2TIM|1|5|recordationem accipiens eius fidei, quae est in te non ficta, quae et habitavit primum in avia tua Loide et matre tua Eunice, certus sum autem quod et in te.
2TIM|1|6|Propter quam causam admoneo te, ut resuscites donationem Dei, quae est in te per impositionem manuum mearum;
2TIM|1|7|non enim dedit nobis Deus Spiritum timoris sed virtutis et dilectionis et sobrietatis.
2TIM|1|8|Noli itaque erubescere testimonium Domini nostri neque me vinctum eius, sed collabora evangelio secundum virtutem Dei,
2TIM|1|9|qui nos salvos fecit et vocavit vocatione sancta, non secundum opera nostra sed secundum propositum suum et gratiam, quae data est nobis in Christo Iesu ante tempora saecularia;
2TIM|1|10|manifestata autem nunc per illustrationem salvatoris nostri Iesu Christi, qui destruxit quidem mortem, illuminavit autem vitam et incorruptionem per evangelium,
2TIM|1|11|in quo positus sum ego praedicator et apostolus et doctor.
2TIM|1|12|Ob quam causam etiam haec patior, sed non confundor; scio enim, cui credidi, et certus sum quia potens est depositum meum servare in illum diem.
2TIM|1|13|Formam habe sanorum verborum, quae a me audisti, in fide et dilectione, quae sunt in Christo Iesu;
2TIM|1|14|bonum depositum custodi per Spiritum Sanctum, qui habitat in nobis.
2TIM|1|15|Scis hoc, quod aversi sunt a me omnes, qui in Asia sunt, ex quibus est Phygelus et Hermogenes.
2TIM|1|16|Det misericordiam Dominus Onesiphori domui, quia saepe me refrigeravit et catenam meam non erubuit;
2TIM|1|17|sed cum Romam venisset, sollicite me quaesivit et invenit
2TIM|1|18|det illi Dominus invenire misericordiam a Domino in illa die et quanta Ephesi ministravit, melius tu nosti.
2TIM|2|1|Tu ergo, fili mi, confortare in gratia, quae est in Christo Iesu;
2TIM|2|2|et quae audisti a me per multos testes, haec commenda fidelibus hominibus, qui idonei erunt et alios docere.
2TIM|2|3|Collabora sicut bonus miles Christi Iesu.
2TIM|2|4|Nemo militans implicat se saeculi negotiis, ut ei placeat, qui eum elegit;
2TIM|2|5|si autem certat quis agone, non coronatur nisi legitime certaverit.
2TIM|2|6|Laborantem agricolam oportet primum de fructibus accipere.
2TIM|2|7|Intellege, quae dico; dabit enim tibi Dominus in omnibus intellectum.
2TIM|2|8|Memor esto Iesum Christum resuscitatum esse a mortuis, ex semine David, secundum evangelium meum,
2TIM|2|9|in quo laboro usque ad vincula quasi male operans; sed verbum Dei non est alligatum!
2TIM|2|10|Ideo omnia sustineo propter electos, ut et ipsi salutem consequantur, quae est in Christo Iesu cum gloria aeterna.
2TIM|2|11|Fidelis sermo, Nam, si commortui sumus, et convivemus;
2TIM|2|12|si sustinemus, et conregnabimus; si negabimus, et ille negabit nos;
2TIM|2|13|si non credimus, ille fidelis manet, negare enim seipsum non potest.
2TIM|2|14|Haec commone testificans coram Deo verbis non contendere: in nihil utile est, nisi ad subversionem audientium.
2TIM|2|15|Sollicite cura teipsum probabilem exhibere Deo, operarium inconfusibilem, recte tractantem verbum veritatis.
2TIM|2|16|Profana autem inaniloquia devita, magis enim proficient ad impietatem,
2TIM|2|17|et sermo eorum ut cancer serpit; ex quibus est Hymenaeus et Philetus,
2TIM|2|18|qui circa veritatem aberraverunt dicentes resurrectionem iam factam, et subvertunt quorundam fidem.
2TIM|2|19|Sed firmum fundamentum Dei stat habens signaculum hoc: Cognovit Dominus, qui sunt eius, et: Discedat ab iniquitate omnis, qui nominat nomen Domini.
2TIM|2|20|In magna autem domo non solum sunt vasa aurea et argentea sed et lignea et fictilia, et quaedam quidem in honorem, quaedam autem in ignominiam;
2TIM|2|21|si quis ergo emundaverit se ab istis, erit vas in honorem, sanctificatum, utile Domino, ad omne opus bonum paratum.
2TIM|2|22|Iuvenilia autem desideria fuge, sectare vero iustitiam, fidem, caritatem, pacem cum his, qui invocant Dominum de corde puro.
2TIM|2|23|Stultas autem et sine disciplina quaestiones devita, sciens quia generant lites;
2TIM|2|24|servum autem Domini non oportet litigare, sed mansuetum esse ad omnes, aptum ad docendum, patientem,
2TIM|2|25|cum mansuetudine corripientem eos, qui resistunt, si quando det illis Deus paenitentiam ad cognoscendam veritatem,
2TIM|2|26|et resipiscant a Diaboli laqueo, a quo capti tenentur ad ipsius voluntatem.
2TIM|3|1|Hoc autem scito, quod in no vissimis diebus instabunt tem pora periculosa.
2TIM|3|2|Erunt enim homines seipsos amantes, cupidi, elati, superbi, blasphemi, parentibus inoboedientes, ingrati, scelesti,
2TIM|3|3|sine affectione, sine foedere, criminatores, incontinentes, immites, sine benignitate,
2TIM|3|4|proditores, protervi, tumidi, voluptatum amatores magis quam Dei,
2TIM|3|5|habentes speciem quidem pietatis, virtutem autem eius abnegantes; et hos devita.
2TIM|3|6|Ex his enim sunt, qui penetrant domos et captivas ducunt mulierculas oneratas peccatis, quae ducuntur variis concupiscentiis,
2TIM|3|7|semper discentes et numquam ad scientiam veritatis pervenire valentes.
2TIM|3|8|Quemadmodum autem Iannes et Iambres restiterunt Moysi, ita et hi resistunt veritati, homines corrupti mente, reprobi circa fidem;
2TIM|3|9|sed ultra non proficient, insipientia enim eorum manifesta erit omnibus, sicut et illorum fuit.
2TIM|3|10|Tu autem assecutus es meam doctrinam, institutionem, propositum, fidem, longanimitatem, dilectionem, patientiam,
2TIM|3|11|persecutiones, passiones, qualia mihi facta sunt Antiochiae, Iconii, Lystris, quales persecutiones sustinui; et ex omnibus me eripuit Dominus.
2TIM|3|12|Et omnes, qui volunt pie vivere in Christo Iesu, persecutionem patientur;
2TIM|3|13|mali autem homines et seductores proficient in peius, in errorem mittentes et errantes.
2TIM|3|14|Tu vero permane in his, quae didicisti et credita sunt tibi, sciens a quibus didiceris,
2TIM|3|15|et quia ab infantia Sacras Litteras nosti, quae te possunt instruere ad salutem per fidem, quae est in Christo Iesu.
2TIM|3|16|Omnis Scriptura divinitus inspirata est et utilis ad docendum, ad arguendum, ad corrigendum, ad erudiendum in iustitia,
2TIM|3|17|ut perfectus sit homo Dei, ad omne opus bonum instructus.
2TIM|4|1|Testificor coram Deo et Christo Iesu, qui iudicaturus est vivos ac mortuos, per adventum ipsius et regnum eius:
2TIM|4|2|praedica verbum, insta opportune, importune, argue, increpa, obsecra in omni longanimitate et doctrina.
2TIM|4|3|Erit enim tempus, cum sanam doctrinam non sustinebunt, sed ad sua desideria coacervabunt sibi magistros prurientes auribus,
2TIM|4|4|et a veritate quidem auditum avertent, ad fabulas autem convertentur.
2TIM|4|5|Tu vero vigila in omnibus, labora, opus fac evangelistae, ministerium tuum imple.
2TIM|4|6|Ego enim iam delibor, et tempus meae resolutionis instat.
2TIM|4|7|Bonum certamen certavi, cursum consummavi, fidem servavi;
2TIM|4|8|in reliquo reposita est mihi iustitiae corona, quam reddet mihi Dominus in illa die, iustus iudex, non solum autem mihi sed et omnibus, qui diligunt adventum eius.
2TIM|4|9|Festina venire ad me cito.
2TIM|4|10|Demas enim me dereliquit diligens hoc saeculum et abiit Thessalonicam, Crescens in Galatiam, Titus in Dalmatiam;
2TIM|4|11|Lucas est mecum solus. Marcum assumens adduc tecum, est enim mihi utilis in ministerium.
2TIM|4|12|Tychicum autem misi Ephesum.
2TIM|4|13|Paenulam, quam reliqui Troade apud Carpum, veniens affer, et libros, maxime autem membranas.
2TIM|4|14|Alexander aerarius multa mala mihi ostendit. Reddet ei Dominus secundum opera eius;
2TIM|4|15|quem et tu devita, valde enim restitit verbis nostris.
2TIM|4|16|In prima mea defensione nemo mihi affuit, sed omnes me dereliquerunt. Non illis reputetur;
2TIM|4|17|Dominus autem mihi astitit et confortavit me, ut per me praedicatio impleatur, et audiant omnes gentes; et liberatus sum de ore leonis.
2TIM|4|18|Liberabit me Dominus ab omni opere malo et salvum faciet in regnum suum caeleste; cui gloria in saecula saeculorum. Amen.
2TIM|4|19|Saluta Priscam et Aquilam et Onesiphori domum.
2TIM|4|20|Erastus remansit Corinthi, Trophimum autem reliqui infirmum Mileti.
2TIM|4|21|Festina ante hiemem venire.Salutat te Eubulus et Pudens et Linus et Claudia et fratres omnes.
2TIM|4|22|Dominus cum spiritu tuo. Gratia vobiscum.
TITUS|1|1|Paulus servus Dei, apostolus autem Iesu Christi secundum fi dem electorum Dei et agnitionem veritatis, quae secundum pietatem est
TITUS|1|2|in spem vitae aeternae, quam promisit, qui non mentitur, Deus ante tempora saecularia;
TITUS|1|3|manifestavit autem temporibus suis verbum suum in praedicatione, quae credita est mihi secundum praeceptum salvatoris nostri Dei,
TITUS|1|4|Tito germano filio secundum communem fidem: gratia et pax a Deo Patre et Christo Iesu salvatore nostro.
TITUS|1|5|Huius rei gratia reliqui te Cretae, ut ea, quae desunt, corrigas et constituas per civitates presbyteros, sicut ego tibi disposui,
TITUS|1|6|si quis sine crimine est, unius uxoris vir, filios habens fideles, non in accusatione luxuriae aut non subiectos.
TITUS|1|7|Oportet enim episcopum sine crimine esse sicut Dei dispensatorem, non superbum, non iracundum, non vinolentum, non percussorem, non turpis lucri cupidum,
TITUS|1|8|sed hospitalem, benignum, sobrium, iustum, sanctum, continentem,
TITUS|1|9|amplectentem eum, qui secundum doctrinam est, fidelem sermonem, ut potens sit et exhortari in doctrina sana et eos, qui contradicunt, arguere.
TITUS|1|10|Sunt enim multi et non subiecti, vaniloqui et seductores, maxime qui de circumcisione sunt,
TITUS|1|11|quibus oportet silentium imponere, quia universas domos subvertunt docentes, quae non oportet, turpis lucri gratia.
TITUS|1|12|Dixit quidam ex illis, proprius ipsorum propheta: " Cretenses semper mendaces, malae bestiae, ventres pigri ".
TITUS|1|13|Testimonium hoc verum est. Quam ob causam increpa illos dure, ut sani sint in fide,
TITUS|1|14|non intendentes Iudaicis fabulis et mandatis hominum aversantium veritatem.
TITUS|1|15|Omnia munda mundis; coinquinatis autem et infidelibus nihil mundum, sed inquinatae sunt eorum et mens et conscientia.
TITUS|1|16|Confitentur se nosse Deum, factis autem negant, cum sunt abominati et inoboedientes et ad omne opus bonum reprobi.
TITUS|2|1|Tu autem loquere, quae decent sanam doctrinam.
TITUS|2|2|Senes, ut sobrii sint, pudici, prudentes, sani fide, dilectione, patientia.
TITUS|2|3|Anus similiter in habitu sanctae, non criminatrices, non vino multo deditae, bene docentes,
TITUS|2|4|ut prudentiam doceant adulescentulas, ut viros suos ament, filios diligant,
TITUS|2|5|prudentes sint, castae, domus curam habentes, benignae, subditae suis viris, ut non blasphemetur verbum Dei.
TITUS|2|6|Iuvenes similiter hortare, ut sobrii sint.
TITUS|2|7|In omnibus teipsum praebens exemplum bonorum operum, in doctrina integritatem, gravitatem,
TITUS|2|8|in verbo sano irreprehensibilem, ut is, qui ex adverso est, vereatur, nihil habens malum dicere de nobis.
TITUS|2|9|Servos dominis suis subditos esse in omnibus, placentes esse, non contradicentes,
TITUS|2|10|non fraudantes, sed omnem fidem bonam ostendentes, ut doctrinam salutaris nostri Dei ornent in omnibus.
TITUS|2|11|Apparuit enim gratia Dei salutaris omnibus hominibus
TITUS|2|12|erudiens nos, ut abnegantes impietatem et saecularia desideria sobrie et iuste et pie vivamus in hoc saeculo,
TITUS|2|13|exspectantes beatam spem et adventum gloriae magni Dei et salvatoris nostri Iesu Christi;
TITUS|2|14|qui dedit semetipsum pro nobis, ut nos redimeret ab omni iniquitate et mundaret sibi populum peculiarem, sectatorem bonorum operum.
TITUS|2|15|Haec loquere et exhortare et argue cum omni imperio. Nemo te contemnat!
TITUS|3|1|Admone illos principibus, pote statibus subditos esse, dicto oboedire, ad omne opus bonum paratos esse,
TITUS|3|2|neminem blasphemare, non litigiosos esse, modestos, omnem ostendentes mansuetudinem ad omnes homines.
TITUS|3|3|Eramus enim et nos aliquando insipientes, inoboedientes, errantes, servientes concupiscentiis et voluptatibus variis, in malitia et invidia agentes, odibiles, odientes invicem.
TITUS|3|4|Cum autem benignitas et humanitas apparuit salvatoris nostri Dei,
TITUS|3|5|non ex operibus iustitiae, quae fecimus nos, sed secundum suam misericordiam salvos nos fecit per lavacrum regenerationis et renovationis Spiritus Sancti,
TITUS|3|6|quem effudit super nos abunde per Iesum Christum salvatorem nostrum,
TITUS|3|7|ut iustificati gratia ipsius heredes simus secundum spem vitae aeternae.
TITUS|3|8|Fidelis sermo, et volo te de his confirmare, ut curent bonis operibus praeesse, qui crediderunt Deo. Haec sunt bona et utilia hominibus;
TITUS|3|9|stultas autem quaestiones et genealogias et contentiones et pugnas circa legem devita, sunt enim inutiles et vanae.
TITUS|3|10|Haereticum hominem post unam et secundam correptionem devita,
TITUS|3|11|sciens quia subversus est, qui eiusmodi est, et delinquit, proprio iudicio condemnatus.
TITUS|3|12|Cum misero ad te Artemam aut Tychicum, festina ad me venire Nicopolim; ibi enim statui hiemare.
TITUS|3|13|Zenam legis peritum et Apollo sollicite instrue, ut nihil illis desit.
TITUS|3|14|Discant autem et nostri bonis operibus praeesse ad usus necessarios, ut non sint infructuosi.
TITUS|3|15|Salutant te, qui mecum sunt, omnes. Saluta, qui nos amant in fide.Gratia cum omnibus vobis.
PHLM|1|1|Paulus vinctus Christi Iesu et Timotheus frater Philemoni dilecto et adiutori nostro
PHLM|1|2|et Apphiae sorori et Archippo commilitoni nostro et ecclesiae, quae in domo tua est:
PHLM|1|3|gratia vobis et pax a Deo Patre nostro et Domino Iesu Christo.
PHLM|1|4|Gratias ago Deo meo semper memoriam tui faciens in orationibus meis,
PHLM|1|5|audiens caritatem tuam et fidem, quam habes in Dominum Iesum et in omnes sanctos,
PHLM|1|6|ut communio fidei tuae evidens fiat in agnitione omnis boni, quod est in nobis in Christum;
PHLM|1|7|gaudium enim magnum habui et consolationem in caritate tua, quia viscera sanctorum requieverunt per te, frater.
PHLM|1|8|Propter quod multam fiduciam habens in Christo imperandi tibi, quod ad rem pertinet,
PHLM|1|9|propter caritatem magis obsecro, cum sim talis ut Paulus senex, nunc autem et vinctus Christi Iesu;
PHLM|1|10|obsecro te de meo filio, quem genui in vinculis, Onesimo,
PHLM|1|11|qui tibi aliquando inutilis fuit, nunc autem et tibi et mihi utilis,
PHLM|1|12|quem remisi tibi: eum, hoc est viscera mea;
PHLM|1|13|quem ego volueram mecum detinere, ut pro te mihi ministraret in vinculis evangelii.
PHLM|1|14|Sine consilio autem tuo nihil volui facere, uti ne velut ex necessitate bonum tuum esset sed voluntarium.
PHLM|1|15|Forsitan enim ideo discessit ad horam, ut aeternum illum reciperes,
PHLM|1|16|iam non ut servum sed plus servo, carissimum fratrem, maxime mihi, quanto autem magis tibi et in carne et in Domino.
PHLM|1|17|Si ergo habes me socium, suscipe illum sicut me.
PHLM|1|18|Si autem aliquid nocuit tibi aut debet, hoc mihi imputa.
PHLM|1|19|Ego Paulus scripsi mea manu, ego reddam; ut non dicam tibi quod et teipsum mihi debes.
PHLM|1|20|Ita, frater! Ego te fruar in Domino; refice viscera mea in Christo!
PHLM|1|21|Confidens oboedientia tua scripsi tibi, sciens quoniam et super id, quod dico, facies.
PHLM|1|22|Simul autem et para mihi hospitium, nam spero per orationes vestras donari me vobis.
PHLM|1|23|Salutat te Epaphras, concaptivus meus in Christo Iesu,
PHLM|1|24|Marcus, Aristarchus, Demas, Lucas, adiutores mei.
PHLM|1|25|Gratia Domini Iesu Christi cum spiritu vestro.
HEB|1|1|Multifariam et multis modis olim Deus locutus patribus in prophetis,
HEB|1|2|in novissimis his diebus locutus est nobis in Filio, quem constituit heredem universorum, per quem fecit et saecula;
HEB|1|3|qui, cum sit splendor gloriae et figura substantiae eius et portet omnia verbo virtutis suae, purgatione peccatorum facta, consedit ad dexteram maiestatis in excelsis,
HEB|1|4|tanto melior angelis effectus, quanto differentius prae illis nomen hereditavit.
HEB|1|5|Cui enim dixit aliquando angelorum: Filius meus es tu;ego hodie genui te "et rursum: " Ego ero illi in patrem, et ipse erit mihi in filium "?
HEB|1|6|Cum autem iterum introducit primogenitum in orbem terrae, dicit: Et adorent eum omnes angeli Dei ".
HEB|1|7|Et ad angelos quidem dicit: Qui facit angelos suos spirituset ministros suos flammam ignis ";
HEB|1|8|ad Filium autem: Thronus tuus, Deus, in saeculum saeculi,et virga aequitatis virga regni tui.
HEB|1|9|Dilexisti iustitiam et odisti iniquitatem,propterea unxit te Deus, Deus tuus,oleo exsultationis prae participibus tuis "
HEB|1|10|et: Tu in principio, Domine, terram fundasti;et opera manuum tuarum sunt caeli.
HEB|1|11|Ipsi peribunt, tu autem permanes;et omnes ut vestimentum veterascent,
HEB|1|12|et velut amictum involves eos,sicut vestimentum et mutabuntur.Tu autem idem es, et anni tui non deficient ".
HEB|1|13|Ad quem autem angelorum dixit aliquando: Sede a dextris meis,donec ponam inimicos tuos scabellum pedum tuorum "?
HEB|1|14|Nonne omnes sunt administratorii spiritus, qui in ministerium mittuntur propter eos, qui hereditatem capient salutis?
HEB|2|1|Propterea abundantius oportet observare nos ea, quae audivi mus, ne forte praeterfluamus.
HEB|2|2|Si enim, qui per angelos dictus est, sermo factus est firmus, et omnis praevaricatio et inoboedientia accepit iustam mercedis retributionem,
HEB|2|3|quomodo nos effugiemus, si tantam neglexerimus salutem? Quae, cum initium accepisset enarrari per Dominum, ab eis, qui audierunt, in nos confirmata est,
HEB|2|4|contestante Deo signis et portentis et variis virtutibus et Spiritus Sancti distributionibus secundum suam voluntatem.
HEB|2|5|Non enim angelis subiecit orbem terrae futurum, de quo loquimur.
HEB|2|6|Testatus est autem in quodam loco quis dicens: Quid est homo, quod memor es eius,aut filius hominis, quoniam visitas eum?
HEB|2|7|Minuisti eum paulo minus ab angelis,gloria et honore coronasti eum,
HEB|2|8|omnia subiecisti sub pedibus eius ".In eo enim quod ei omnia subiecit, nihil dimisit non subiectibile ei. Nunc autem necdum videmus omnia subiecta ei;
HEB|2|9|eum autem, qui paulo minus ab angelis minoratus est, videmus Iesum propter passionem mortis gloria et honore coronatum, ut gratia Dei pro omnibus gustaverit mortem.
HEB|2|10|Decebat enim eum, propter quem omnia et per quem omnia, qui multos filios in gloriam adduxit, ducem salutis eorum per passiones consummare.
HEB|2|11|Qui enim sanctificat et qui sanctificantur, ex uno omnes; propter quam causam non erubescit fratres eos vocare
HEB|2|12|dicens: Nuntiabo nomen tuum fratribus meis,in medio ecclesiae laudabo te";
HEB|2|13|et iterum: " Ego ero fidens in eum ";et iterum: " Ecce ego et pueri, quos mihi dedit Deus ".
HEB|2|14|Quia ergo pueri communicaverunt sanguini et carni, et ipse similiter participavit iisdem, ut per mortem destrueret eum, qui habebat mortis imperium, id est Diabolum,
HEB|2|15|et liberaret eos, qui timore mortis per totam vitam obnoxii erant servituti.
HEB|2|16|Nusquam enim angelos apprehendit, sed semen Abrahae apprehendit.
HEB|2|17|Unde debuit per omnia fratribus similari, ut misericors fieret et fidelis pontifex in iis,quae sunt ad Deum, ut repropitiaret delicta populi;
HEB|2|18|in quo enim passus est ipse tentatus, po tens est eis, qui tentantur, auxiliari.
HEB|3|1|Unde, fratres sancti, vocationis caelestis participes, considerate apostolum et pontificem confessionis nostrae Iesum,
HEB|3|2|qui fidelis est ei, qui fecit illum, sicut et Moyses in tota domo illius.
HEB|3|3|Amplioris enim gloriae iste prae Moyse dignus est habitus, quanto ampliorem honorem habet quam domus, qui fabricavit illam.
HEB|3|4|Omnis namque domus fabricatur ab aliquo; qui autem omnia fabricavit, Deus est.
HEB|3|5|Et Moyses quidem fidelis erat in tota domo eius tamquam famulus in testimonium eorum, quae dicenda erant,
HEB|3|6|Christus vero tamquam Filius super domum illius; cuius domus sumus nos, si fiduciam et gloriationem spei retineamus.
HEB|3|7|Quapropter, sicut dicit Spiritus Sanctus: Hodie, si vocem eius audieritis,
HEB|3|8|nolite obdurare corda vestra sicut in exacerbatione,secundum diem tentationis in deserto,
HEB|3|9|ubi tentaverunt me patres vestri in probationeet viderunt opera mea
HEB|3|10|quadraginta annos. Propter quod infensus fui generationi huic et dixi: Semper errant corde.Ipsi autem non cognoverunt vias meas;
HEB|3|11|sicut icut iuravi in ira mea:Non introibunt in requiem meam ".
HEB|3|12|Videte, fratres, ne forte sit in aliquo vestrum cor malum incredulitatis discedendi a Deo vivo,
HEB|3|13|sed adhortamini vosmetipsos per singulos dies, donec illud " hodie " vocatur, ut non obduretur quis ex vobis fallacia peccati;
HEB|3|14|participes enim Christi effecti sumus, si tamen initium substantiae usque ad finem firmum retineamus,
HEB|3|15|dum dicitur: Hodie, si vocem eius audieritis,nolite obdurare corda vestra quemadmodum in illa exacerbatione ".
HEB|3|16|Qui sunt enim qui audientes exacerbaverunt? Nonne universi, qui profecti sunt ab Aegypto per Moysen?
HEB|3|17|Quibus autem infensus fuit quadraginta annos? Nonne illis, qui peccaverunt, quorum membra ceciderunt in deserto?
HEB|3|18|Quibus autem iuravit non introire in requiem ipsius, nisi illis, qui increduli fuerunt?
HEB|3|19|Et videmus quia non potuerunt introire propter incredulitatem.
HEB|4|1|Timeamus ergo, ne forte, relicta pollicitatione introeundi in re quiem eius, existimetur aliquis ex vobis deesse;
HEB|4|2|etenim et nobis evangelizatum est quemadmodum et illis, sed non profuit illis sermo auditus, non commixtis fide cum iis, qui audierant.
HEB|4|3|Ingredimur enim in requiem, qui credidimus, quemadmodum dixit: Sicut iuravi in ira mea:Non introibunt in requiem meam ",et quidem operibus ab institutione mundi factis.
HEB|4|4|Dixit enim quodam loco de die septima sic: "Et requievit Deus die septima ab omnibus operibus suis ";
HEB|4|5|et in isto rursum: " Non introibunt in requiem meam ".
HEB|4|6|Quoniam ergo superest quosdam introire in illam, et hi, quibus prioribus evangelizatum est, non introierunt propter inoboedientiam,
HEB|4|7|iterum terminat diem quendam, " Hodie ", in David dicendo post tantum temporis, sicut supra dictum est: Hodie, si vocem eius audieritis,nolite obdurare corda vestra ".
HEB|4|8|Nam, si eis Iesus requiem praestitisset, non de alio loqueretur posthac die.
HEB|4|9|Itaque relinquitur sabbatismus populo Dei;
HEB|4|10|qui enim ingressus est in requiem eius, etiam ipse requievit ab operibus suis, sicut a suis Deus.
HEB|4|11|Festinemus ergo ingredi in illam requiem, ut ne in idipsum quis incidat inoboedientiae exemplum.
HEB|4|12|Vivus est enim Dei sermo et efficax et penetrabilior omni gladio ancipiti et pertingens usque ad divisionem animae ac spiritus, compagum quoque et medullarum, et discretor cogitationum et intentionum cordis;
HEB|4|13|et non est creatura invisibilis in conspectu eius, omnia autem nuda et aperta sunt oculis eius, ad quem nobis sermo.
HEB|4|14|Habentes ergo pontificem magnum, qui penetravit caelos, Iesum Filium Dei, teneamus confessionem.
HEB|4|15|Non enim habemus pontificem, qui non possit compati infirmitatibus nostris, tentatum autem per omnia secundum similitudinem absque peccato;
HEB|4|16|adeamus ergo cum fiducia ad thronum gratiae, ut misericordiam consequamur et gratiam inveniamus in auxilium opportunum.
HEB|5|1|Omnis namque pontifex ex hominibus assumptus pro homi nibus constituitur in his, quae sunt ad Deum, ut offerat dona et sacrificia pro peccatis;
HEB|5|2|qui aeque condolere possit his, qui ignorant et errant, quoniam et ipse circumdatus est infirmitate
HEB|5|3|et propter eam debet, quemadmodum et pro populo, ita etiam pro semetipso offerre pro peccatis.
HEB|5|4|Nec quisquam sumit sibi illum honorem, sed qui vocatur a Deo tamquam et Aaron.
HEB|5|5|Sic et Christus non semetipsum glorificavit, ut pontifex fieret, sed qui locutus est ad eum: Filius meus es tu;ego hodie genui te ";
HEB|5|6|quemadmodum et in alio dicit: Tu es sacerdos in aeternum secundum ordinem Melchisedech ".
HEB|5|7|Qui in diebus carnis suae, preces supplicationesque ad eum, qui possit salvum illum a morte facere, cum clamore valido et lacrimis offerens et exauditus pro sua reverentia,
HEB|5|8|et quidem cum esset Filius, didicit ex his, quae passus est, oboedientiam;
HEB|5|9|et, consummatus, factus est omnibus oboedientibus sibi auctor salutis aeternae,
HEB|5|10|appellatus a Deo pontifex iuxta ordinem Melchisedech.
HEB|5|11|De quo grandis nobis sermo et ininterpretabilis ad dicendum, quoniam segnes facti estis ad audiendum.
HEB|5|12|Etenim cum deberetis magistri esse propter tempus, rursum indigetis, ut vos doceat aliquis elementa exordii sermonum Dei, et facti estis, quibus lacte opus sit, non solido cibo.
HEB|5|13|Omnis enim, qui lactis est particeps, expers est sermonis iustitiae, parvulus enim est;
HEB|5|14|perfectorum autem est solidus cibus, eorum, qui pro consuetudine exercitatos habent sensus ad discretionem boni ac mali.
HEB|6|1|Quapropter praetermittentes inchoationis Christi sermonem ad perfectionem feramur, non rursum iacientes fundamentum paenitentiae ab operibus mortuis et fidei ad Deum,
HEB|6|2|baptismatum doctrinae, impositionis quoque manuum, ac resurrectionis mortuorum et iudicii aeterni.
HEB|6|3|Et hoc faciemus, si quidem permiserit Deus.
HEB|6|4|Impossibile est enim eos, qui semel sunt illuminati, gustaverunt etiam donum caeleste et participes sunt facti Spiritus Sancti
HEB|6|5|et bonum gustaverunt Dei verbum virtutesque saeculi venturi
HEB|6|6|et prolapsi sunt, rursus renovari ad paenitentiam, rursum crucifigentes sibimetipsis Filium Dei et ostentui habentes.
HEB|6|7|Terra enim saepe venientem super se bibens imbrem et generans herbam opportunam illis, propter quos et colitur, accipit benedictionem a Deo;
HEB|6|8|proferens autem spinas ac tribulos reproba est et maledicto proxima, cuius finis in combustionem.
HEB|6|9|Confidimus autem de vobis, dilectissimi, meliora et viciniora saluti, tametsi ita loquimur;
HEB|6|10|non enim iniustus Deus, ut obliviscatur operis vestri et dilectionis, quam ostendistis nomini ipsius, qui ministrastis sanctis et ministratis.
HEB|6|11|Cupimus autem unumquemque vestrum eandem ostentare sollicitudinem ad expletionem spei usque in finem,
HEB|6|12|ut non segnes efficiamini, verum imitatores eorum, qui fide et patientia hereditant promissiones.
HEB|6|13|Abrahae namque promittens Deus, quoniam neminem habuit, per quem iuraret maiorem, iuravit per semetipsum
HEB|6|14|dicens: " Utique benedicens benedicam te et multiplicans multiplicabo te ";
HEB|6|15|et sic longanimiter ferens adeptus est repromissionem.
HEB|6|16|Homines enim per maiorem sui iurant, et omnis controversiae eorum finis ad confirmationem est iuramentum;
HEB|6|17|in quo abundantius volens Deus ostendere pollicitationis heredibus immobilitatem consilii sui, se interposuit iure iurando,
HEB|6|18|ut per duas res immobiles, in quibus impossibile est mentiri Deum, fortissimum solacium habeamus, qui confugimus ad tenendam propositam spem;
HEB|6|19|quam sicut ancoram habemus animae, tutam ac firmam et incedentem usque in interiora velaminis,
HEB|6|20|ubi praecursor pro nobis introivit Iesus, secundum ordinem Melchisedech pontifex factus in aeternum.
HEB|7|1|Hic enim Melchisedech, rex Salem, sacerdos Dei summi, qui ob viavit Abrahae regresso a caede regum et benedixit ei,
HEB|7|2|cui et decimam omnium divisit Abraham, primum quidem, qui interpretatur rex iustitiae, deinde autem et rex Salem, quod est rex Pacis,
HEB|7|3|sine patre, sine matre, sine genealogia, neque initium dierum neque finem vitae habens, assimilatus autem Filio Dei, manet sacerdos in perpetuum.
HEB|7|4|Intuemini autem quantus sit hic, cui et decimam dedit de praecipuis Abraham patriarcha.
HEB|7|5|Et illi quidem, qui de filiis Levi sacerdotium accipiunt, mandatum habent decimas sumere a populo secundum legem, id est a fratribus suis, quamquam et ipsi exierunt de lumbis Abrahae;
HEB|7|6|hic autem, cuius generatio non annumeratur in eis, decimam sumpsit ab Abraham et eum, qui habebat repromissiones, benedixit.
HEB|7|7|Sine ulla autem contradictione, quod minus est, a meliore benedicitur.
HEB|7|8|Et hic quidem decimas morientes homines sumunt; ibi autem testimonium accipiens quia vivit.
HEB|7|9|Et, ut ita dictum sit, per Abraham et Levi, qui decimas accipit, decimatus est;
HEB|7|10|adhuc enim in lumbis patris erat, quando obviavit ei Melchisedech.
HEB|7|11|Si ergo consummatio per sacerdotium leviticum erat, populus enim sub ipso legem accepit, quid adhuc necessarium secundum ordinem Melchisedech alium surgere sacerdotem et non secundum ordinem Aaron dici?
HEB|7|12|Translato enim sacerdotio, necesse est, ut et legis translatio fiat.
HEB|7|13|De quo enim haec dicuntur, ex alia tribu est, ex qua nullus altari praesto fuit;
HEB|7|14|manifestum enim quod ex Iuda ortus sit Dominus noster, in quam tribum nihil de sacerdotibus Moyses locutus est.
HEB|7|15|Et amplius adhuc manifestum est, si secundum similitudinem Melchisedech exsurgit alius sacerdos,
HEB|7|16|qui non secundum legem mandati carnalis factus est sed secundum virtutem vitae insolubilis,
HEB|7|17|testimonium enim accipit: Tu es sacerdos in aeternum secundum ordinem Melchisedech ".
HEB|7|18|Reprobatio quidem fit praecedentis mandati propter infirmitatem eius et inutilitatem,
HEB|7|19|nihil enim ad perfectum adduxit lex; introductio vero melioris spei, per quam proximamus ad Deum.
HEB|7|20|Et quantum non est sine iure iurando; illi quidem sine iure iurando sacerdotes facti sunt,
HEB|7|21|hic autem cum iure iurando per eum, qui dicit ad illum: Iuravit Dominus et non paenitebit eum: Tu es sacerdos in aeternum ",
HEB|7|22|in tantum et melioris testamenti sponsor factus est Iesus.
HEB|7|23|Et illi quidem plures facti sunt sacerdotes, idcirco quod morte prohibebantur permanere;
HEB|7|24|hic autem eo quod manet in aeternum, intransgressibile habet sacerdotium;
HEB|7|25|unde et salvare in perpetuum potest accedentes per semetipsum ad Deum, semper vivens ad interpellandum pro eis.
HEB|7|26|Talis enim et decebat ut nobis esset pontifex, sanctus, innocens, impollutus, segregatus a peccatoribus et excelsior caelis factus;
HEB|7|27|qui non habet necessitatem cotidie, quemadmodum pontifices, prius pro suis delictis hostias offerre, deinde pro populi; hoc enim fecit semel semetipsum offerendo.
HEB|7|28|Lex enim homines constituit pontifices infirmitatem habentes; sermo autem iuris iurandi, quod post legem est, Filium in aeternum consummatum.
HEB|8|1|Caput autem super ea, quae dicuntur: talem habemus ponti ficem, qui consedit in dextera throni Maiestatis in caelis,
HEB|8|2|sanctorum minister et tabernaculi veri, quod fixit Dominus, non homo.
HEB|8|3|Omnis enim pontifex ad offerenda munera et hostias constituitur; unde necesse erat et hunc habere aliquid, quod offerret.
HEB|8|4|Si ergo esset super terram, nec esset sacerdos, cum sint qui offerant secundum legem munera;
HEB|8|5|qui figurae et umbrae deserviunt caelestium, sicut responsum est Moysi, cum consummaturus esset tabernaculum: " Vide enim, inquit, omnia facies secundum exemplar, quod tibi ostensum est in monte ".
HEB|8|6|Nunc autem differentius sortitus est ministerium, quanto et melioris testamenti mediator est, quod in melioribus repromissionibus sancitum est.
HEB|8|7|Nam si illud prius culpa vacasset, non secundi locus inquireretur;
HEB|8|8|vituperans enim eos dicit: " Ecce dies veniunt, dicit Dominus, et consummabo super domum Israel et super domum Iudae testamentum novum;
HEB|8|9|non secundum testamentum, quod feci patribus eorum in die, qua apprehendi manum illorum, ut educerem illos de terra Aegypti; quoniam ipsi non permanserunt in testamento meo, et ego neglexi eos, dicit Dominus.
HEB|8|10|Quia hoc est testamentum, quod testabor domui Israel post dies illos, dicit Dominus, dando leges meas in mentem eorum, et in corde eorum superscribam eas; et ero eis in Deum, et ipsi erunt mihi in populum.
HEB|8|11|Et non docebit unusquisque civem suum, et unusquisque fratrem suum dicens: "Cognosce Dominum"; quoniam omnes scient me, a minore usque ad maiorem eorum,
HEB|8|12|quia propitius ero iniquitatibus eorum et peccatorum illorum iam non memorabor ".
HEB|8|13|Dicendo " novum " veteravit prius; quod autem antiquatur et senescit, prope interitum est.
HEB|9|1|Habuit ergo et prius praecepta cultus et Sanctum huius saeculi.
HEB|9|2|Tabernaculum enim praeparatum est primum, in quo inerat candelabrum et mensa et propositio panum, quod dicitur Sancta;
HEB|9|3|post secundum autem velamentum, tabernaculum, quod dicitur Sancta Sanctorum,
HEB|9|4|aureum habens turibulum et arcam testamenti circumtectam ex omni parte auro, in qua urna aurea habens manna et virga Aaron, quae fronduerat, et tabulae testamenti,
HEB|9|5|superque eam cherubim gloriae obumbrantia propitiatorium; de quibus non est modo dicendum per singula.
HEB|9|6|His vero ita praeparatis, in prius quidem tabernaculum semper intrant sacerdotes sacrorum officia consummantes;
HEB|9|7|in secundum autem semel in anno solus pontifex, non sine sanguine, quem offert pro suis et populi ignorantiis;
HEB|9|8|hoc significante Spiritu Sancto, nondum propalatam esse sanctorum viam, adhuc priore tabernaculo habente statum;
HEB|9|9|quae parabola est temporis instantis, iuxta quam munera et hostiae offeruntur, quae non possunt iuxta conscientiam perfectum facere servientem,
HEB|9|10|solummodo in cibis et in potibus et variis baptismis, quae sunt praecepta carnis usque ad tempus correctionis imposita.
HEB|9|11|Christus autem cum advenit pontifex futurorum bonorum, per amplius et perfectius tabernaculum, non manufactum, id est non huius creationis,
HEB|9|12|neque per sanguinem hircorum et vitulorum sed per proprium sanguinem introivit semel in Sancta, aeterna redemptione inventa.
HEB|9|13|Si enim sanguis hircorum et taurorum et cinis vitulae aspersus inquinatos sanctificat ad emundationem carnis,
HEB|9|14|quanto magis sanguis Christi, qui per Spiritum aeternum semetipsum obtulit immaculatum Deo, emundabit conscientiam nostram ab operibus mortuis ad serviendum Deo viventi.
HEB|9|15|Et ideo novi testamenti mediator est, ut, morte intercedente in redemptionem earum praevaricationum, quae erant sub priore testamento, repromissionem accipiant, qui vocati sunt aeternae hereditatis.
HEB|9|16|Ubi enim testamentum, mors necesse est afferatur testatoris;
HEB|9|17|testamentum autem in mortuis est confirmatum, nondum enim valet, dum vivit, qui testatus est.
HEB|9|18|Unde ne prius quidem sine sanguine dedicatum est;
HEB|9|19|enuntiato enim omni mandato secundum legem a Moyse universo populo, accipiens sanguinem vitulorum et hircorum cum aqua et lana coccinea et hyssopo, ipsum librum et omnem populum aspersit
HEB|9|20|dicens: " Hic sanguis testamenti, quod mandavit ad vos Deus ";
HEB|9|21|etiam tabernaculum et omnia vasa ministerii sanguine similiter aspersit.
HEB|9|22|Et omnia paene in sanguine mundantur secundum legem, et sine sanguinis effusione non fit remissio.
HEB|9|23|Necesse erat ergo figuras quidem caelestium his mundari, ipsa autem caelestia melioribus hostiis quam istis.
HEB|9|24|Non enim in manufacta Sancta Christus introivit, quae sunt similitudo verorum, sed in ipsum caelum, ut appareat nunc vultui Dei pro nobis;
HEB|9|25|neque ut saepe offerat semetipsum, quemadmodum pontifex intrat in Sancta per singulos annos in sanguine alieno.
HEB|9|26|Alioquin oportebat eum frequenter pati ab origine mundi; nunc autem semel in consummatione saeculorum ad destitutionem peccati per sacrificium sui manifestatus est.
HEB|9|27|Et quemadmodum statutum est hominibus semel mori, post hoc autem iudicium,
HEB|9|28|sic et Christus, semel oblatus ad multorum auferenda peccata, secundo sine peccato apparebit exspectantibus se in salutem.
HEB|10|1|Umbram enim habens lex bonorum futurorum, non ip sam imaginem rerum, per singulos annos iisdem ipsis hostiis, quas offerunt indesinenter, numquam potest accedentes perfectos facere.
HEB|10|2|Alioquin nonne cessassent offerri, ideo quod nullam haberent ultra conscientiam peccatorum cultores semel mundati?
HEB|10|3|Sed in ipsis commemoratio peccatorum per singulos annos fit.
HEB|10|4|Impossibile enim est sanguinem taurorum et hircorum auferre peccata.
HEB|10|5|Ideo ingrediens mundum dicit: Hostiam et oblationem noluisti,corpus autem aptasti mihi;
HEB|10|6|holocautomata et sacrificia pro peccatonon tibi placuerunt.
HEB|10|7|Tunc dixi: Ecce venio,in capitulo libri scriptum est de me,ut faciam, Deus, voluntatem tuam ".
HEB|10|8|Superius dicens: " Hostias et oblationes et holocautomata et sacrificia pro peccato noluisti, nec placuerunt tibi ", quae secundum legem offeruntur,
HEB|10|9|tunc dixit: " Ecce venio, ut faciam voluntatem tuam ". Aufert primum, ut secundum statuat;
HEB|10|10|in qua voluntate sanctificati sumus per oblationem corporis Christi Iesu in semel.
HEB|10|11|Et omnis quidem sacerdos stat cotidie ministrans et easdem saepe offerens hostias, quae numquam possunt auferre peccata.
HEB|10|12|Hic autem, una pro peccatis oblata hostia, in sempiternum consedit in dextera Dei,
HEB|10|13|de cetero exspectans, donec ponantur inimici eius scabellum pedum eius;
HEB|10|14|una enim oblatione consummavit in sempiternum eos, qui sanctificantur.
HEB|10|15|Testificatur autem nobis et Spiritus Sanctus; postquam enim dixit:
HEB|10|16|" Hoc est testamentum, quod testabor ad illos post dies illos, dicit Dominus, dando leges meas in cordibus eorum, et in mente eorum superscribam eas;
HEB|10|17|et peccatorum eorum et iniquitatum eorum iam non recordabor amplius ".
HEB|10|18|Ubi autem horum remissio, iam non oblatio pro peccato.
HEB|10|19|Habentes itaque, fratres, fiduciam in introitum Sanctorum in sanguine Iesu,
HEB|10|20|quam initiavit nobis viam novam et viventem per velamen, id est carnem suam,
HEB|10|21|et sacerdotem magnum super domum Dei,
HEB|10|22|accedamus cum vero corde in plenitudine fidei, aspersi corda a conscientia mala et abluti corpus aqua munda;
HEB|10|23|teneamus spei confessionem indeclinabilem, fidelis enim est, qui repromisit;
HEB|10|24|et consideremus invicem in provocationem caritatis et bonorum operum,
HEB|10|25|non deserentes congregationem nostram, sicut est consuetudinis quibusdam, sed exhortantes, et tanto magis quanto videtis appropinquantem diem.
HEB|10|26|Voluntarie enim peccantibus nobis, post acceptam notitiam veritatis, iam non relinquitur pro peccatis hostia,
HEB|10|27|terribilis autem quaedam exspectatio iudicii, et ignis aemulatio, quae consumptura est adversarios.
HEB|10|28|Irritam quis faciens legem Moysis, sine ulla miseratione duobus vel tribus testibus moritur;
HEB|10|29|quanto deteriora putatis merebitur supplicia, qui Filium Dei conculcaverit et sanguinem testamenti communem duxerit, in quo sanctificatus est, et Spiritui gratiae contumeliam fecerit?
HEB|10|30|Scimus enim eum, qui dixit: " Mihi vindicta, ego retribuam "; et iterum: " Iudicabit Dominus populum suum ".
HEB|10|31|Horrendum est incidere in manus Dei viventis.
HEB|10|32|Rememoramini autem pristinos dies, in quibus illuminati magnum certamen sustinuistis passionum,
HEB|10|33|in altero quidem opprobriis et tribulationibus spectaculum facti, in altero autem socii taliter conversantium effecti;
HEB|10|34|nam et vinctis compassi estis et rapinam bonorum vestrorum cum gaudio suscepistis, cognoscentes vos habere meliorem substantiam et manentem.
HEB|10|35|Nolite itaque abicere confidentiam vestram, quae magnam habet remunerationem;
HEB|10|36|patientia enim vobis necessaria est, ut voluntatem Dei facientes reportetis promissionem.
HEB|10|37|Adhuc enim modicum quantulum,qui venturus est, veniet et non tardabit.
HEB|10|38|Iustus autem meus ex fide vivet;quod si subtraxerit se,non sibi complacet in eo anima mea.
HEB|10|39|Nos autem non sumus subtractionis in perditionem, sed fidei in acquisitionem animae.
HEB|11|1|Est autem fides sperando rum substantia, rerum argu mentum non apparentium.
HEB|11|2|In hac enim testimonium consecuti sunt seniores.
HEB|11|3|Fide intellegimus aptata esse saecula verbo Dei, ut ex invisibilibus visibilia facta sint.
HEB|11|4|Fide ampliorem hostiam Abel quam Cain obtulit Deo, per quam testimonium consecutus est esse iustus, testimonium perhibente muneribus eius Deo; et per illam defunctus adhuc loquitur.
HEB|11|5|Fide Henoch translatus est, ne videret mortem, et non inveniebatur, quia transtulit illum Deus; ante translationem enim testimonium accepit placuisse Deo.
HEB|11|6|Sine fide autem impossibile placere; credere enim oportet accedentem ad Deum quia est et inquirentibus se remunerator fit.
HEB|11|7|Fide Noe, responso accepto de his, quae adhuc non videbantur, reveritus aptavit arcam in salutem domus suae; per quam damnavit mundum, et iustitiae, quae secundum fidem est, heres est institutus.
HEB|11|8|Fide vocatus Abraham oboedivit in locum exire, quem accepturus erat in hereditatem; et exivit nesciens quo iret.
HEB|11|9|Fide peregrinatus est in terra promissionis tamquam in aliena, in casulis habitando cum Isaac et Iacob, coheredibus promissionis eiusdem;
HEB|11|10|exspectabat enim fundamenta habentem civitatem, cuius artifex et conditor Deus.
HEB|11|11|Fide - et ipsa Sara sterilis - virtutem in conceptionem seminis accepit etiam praeter tempus aetatis, quoniam fidelem credidit esse, qui promiserat;
HEB|11|12|propter quod et ab uno orti sunt, et hoc emortuo, tamquam sidera caeli in multitudine, et sicut arena, quae est ad oram maris, innumerabilis.
HEB|11|13|Iuxta fidem defuncti sunt omnes isti, non acceptis promissionibus, sed a longe eas aspicientes et salutantes, et confitentes quia peregrini et hospites sunt supra terram;
HEB|11|14|qui enim haec dicunt, significant se patriam inquirere.
HEB|11|15|Et si quidem illius meminissent, de qua exierant, habebant utique tempus revertendi;
HEB|11|16|nunc autem meliorem appetunt, id est caelestem. Ideo non confunditur Deus vocari Deus eorum, paravit enim illis civitatem.
HEB|11|17|Fide obtulit Abraham Isaac, cum tentaretur; et unigenitum offerebat ille, qui susceperat promissiones,
HEB|11|18|ad quem dictum erat: " In Isaac vocabitur tibi semen ",
HEB|11|19|arbitratus quia et a mortuis suscitare potens est Deus; unde eum et in parabola reportavit.
HEB|11|20|Fide et de futuris benedixit Isaac Iacob et Esau.
HEB|11|21|Fide Iacob moriens singulis filiorum Ioseph benedixit et adoravit super fastigium virgae suae.
HEB|11|22|Fide Ioseph moriens de profectione filiorum Israel memoratus est et de ossibus suis mandavit.
HEB|11|23|Fide Moyses natus occultatus est mensibus tribus a parentibus suis, eo quod vidissent formosum infantem et non timuerunt regis edictum.
HEB|11|24|Fide Moyses grandis factus negavit se dici filium filiae pharaonis,
HEB|11|25|magis eligens affligi cum populo Dei quam temporalem peccati habere iucunditatem,
HEB|11|26|maiores divitias aestimans thesauris Aegypti improperium Christi; aspiciebat enim in remunerationem.
HEB|11|27|Fide reliquit Aegyptum non veritus animositatem regis, invisibilem enim tamquam videns sustinuit.
HEB|11|28|Fide celebravit Pascha et sanguinis effusionem, ne, qui vastabat primogenita, tangeret ea.
HEB|11|29|Fide transierunt mare Rubrum tamquam per aridam terram, quod experti Aegyptii devorati sunt.
HEB|11|30|Fide muri Iericho ruerunt circuiti diebus septem.
HEB|11|31|Fide Rahab meretrix non periit cum incredulis, quia exceperat exploratores cum pace.
HEB|11|32|Et quid adhuc dicam? Deficiet enim me tempus enarrantem de Gedeon, Barac, Samson, Iephte, David et Samuel atque prophetis,
HEB|11|33|qui per fidem devicerunt regna, operati sunt iustitiam, adepti sunt repromissiones, obturaverunt ora leonum,
HEB|11|34|exstinxerunt impetum ignis, effugerunt aciem gladii, convaluerunt de infirmitate, fortes facti sunt in bello, castra verterunt exterorum;
HEB|11|35|acceperunt mulieres de resurrectione mortuos suos; alii autem distenti sunt, non suscipientes redemptionem, ut meliorem invenirent resurrectionem;
HEB|11|36|alii vero ludibria et verbera experti sunt, insuper et vincula et carcerem;
HEB|11|37|lapidati sunt, secti sunt, in occisione gladii mortui sunt, circumierunt in melotis, in pellibus caprinis, egentes, angustiati, afflicti,
HEB|11|38|quibus dignus non erat mundus, in solitudinibus errantes et montibus et speluncis et in cavernis terrae.
HEB|11|39|Et hi omnes testimonium per fidem consecuti non reportaverunt promissionem,
HEB|11|40|Deo pro nobis melius aliquid providente, ut ne sine nobis consummarentur.
HEB|12|1|Ideoque et nos tantam ha bentes circumpositam nobis nubem testium, deponentes omne pondus et circumstans nos peccatum, per patientiam curramus propositum nobis certamen,
HEB|12|2|aspicientes in ducem fidei et consummatorem Iesum, qui pro gaudio sibi proposito sustinuit crucem, confusione contempta, atque in dextera throni Dei sedet.
HEB|12|3|Recogitate enim eum, qui talem sustinuit a peccatoribus adversum semetipsum contradictionem, ut ne fatigemini animis vestris deficientes.
HEB|12|4|Nondum usque ad sanguinem restitistis adversus peccatum repugnantes;
HEB|12|5|et obliti estis exhortationis, quae vobis tamquam filiis loquitur: Fili mi, noli neglegere disciplinam Dominineque deficias, dum ab eo argueris:
HEB|12|6|quem enim diligit, Dominus castigat,flagellat autem omnem filium, quem recipit ".
HEB|12|7|Ad disciplinam suffertis; tamquam filios vos tractat Deus. Quis enim filius, quem non corripit pater?
HEB|12|8|Quod si extra disciplinam estis, cuius participes facti sunt omnes, ergo adulterini et non filii estis!
HEB|12|9|Deinde patres quidem carnis nostrae habebamus eruditores et reverebamur; non multo magis obtemperabimus Patri spirituum et vivemus?
HEB|12|10|Et illi quidem ad tempus paucorum dierum, secundum quod videbatur illis, castigabant; hic autem ad id, quod utile est ad participandam sanctitatem eius.
HEB|12|11|Omnis autem disciplina in praesenti quidem videtur non esse gaudii sed maeroris; postea autem fructum pacificum exercitatis per eam reddit iustitiae.
HEB|12|12|Propter quod remissas manus et soluta genua erigite
HEB|12|13|et gressus rectos facite pedibus vestris, ut, quod claudum est, non extorqueatur, magis autem sanetur.
HEB|12|14|Pacem sectamini cum omnibus et sanctificationem, sine qua nemo videbit Dominum,
HEB|12|15|providentes, ne quis desit gratiae Dei, ne qua radix amaritudinis sursum germinans perturbet, et per illam inquinentur multi;
HEB|12|16|ne quis fornicator aut profanus ut Esau, qui propter unam escam vendidit primogenita sua.
HEB|12|17|Scitis enim quoniam et postea cupiens hereditare benedictionem reprobatus est; non enim invenit paenitentiae locum, quamquam cum lacrimis inquisisset eam.
HEB|12|18|Non enim accessistis ad tractabilem et ardentem ignem et turbinem et caliginem et procellam
HEB|12|19|et tubae sonum et vocem verborum, quam qui audierunt, recusaverunt, ne ultra eis fieret verbum;
HEB|12|20|non enim portabant mandatum: " Et si bestia tetigerit montem, lapidabitur";
HEB|12|21|et ita terribile erat, quod videbatur, Moyses dixit: " Exterritus sum et tremebundus ".
HEB|12|22|Sed accessistis ad Sion montem et civitatem Dei viventis, Ierusalem caelestem, et multa milia angelorum, frequentiam
HEB|12|23|et ecclesiam primogenitorum, qui conscripti sunt in caelis, et iudicem Deum omnium et spiritus iustorum, qui consummati sunt,
HEB|12|24|et testamenti novi mediatorem Iesum et sanguinem aspersionis, melius loquentem quam Abel.
HEB|12|25|Videte, ne recusetis loquentem; si enim illi non effugerunt recusantes eum, qui super terram loquebatur, multo magis nos, qui de caelis loquentem avertimus;
HEB|12|26|cuius vox movit terram tunc, modo autem pronuntiavit dicens: " Adhuc semel ego movebo non solum terram sed et caelum ".
HEB|12|27|Hoc autem " adhuc semel " declarat mobilium translationem tamquam factorum, ut maneant ea, quae sunt immobilia.
HEB|12|28|Itaque, regnum immobile suscipientes, habeamus gratiam, per quam serviamus placentes Deo cum reverentia et metu;
HEB|12|29|etenim Deus noster ignis consumens est.
HEB|13|1|Caritas fraternitatis maneat.
HEB|13|2|Hospitalitatem nolite obli visci; per hanc enim quidam nescientes hospitio receperunt angelos.
HEB|13|3|Mementote vinctorum tamquam simul vincti, laborantium tamquam et ipsi in corpore morantes.
HEB|13|4|Honorabile conubium in omnibus, et torus immaculatus; fornicatores enim et adulteros iudicabit Deus.
HEB|13|5|Sint mores sine avaritia; contenti praesentibus. Ipse enim dixit: " Non te deseram neque derelinquam ",
HEB|13|6|ita ut confidenter dicamus: Dominus mihi adiutor est, non timebo; quid faciet mihi homo? ".
HEB|13|7|Mementote praepositorum vestrorum, qui vobis locuti sunt verbum Dei; quorum intuentes exitum conversationis, imitamini fidem.
HEB|13|8|Iesus Christus heri et hodie idem, et in saecula!
HEB|13|9|Doctrinis variis et peregrinis nolite abduci; optimum enim est gratia stabiliri cor, non escis, quae non profuerunt ambulantibus in eis.
HEB|13|10|Habemus altare, de quo edere non habent potestatem, qui tabernaculo deserviunt.
HEB|13|11|Quorum enim animalium infertur sanguis pro peccato in Sancta per pontificem, horum corpora cremantur extra castra.
HEB|13|12|Propter quod et Iesus, ut sanctificaret per suum sanguinem populum, extra portam passus est.
HEB|13|13|Exeamus igitur ad eum extra castra, improperium eius portantes;
HEB|13|14|non enim habemus hic manentem civitatem, sed futuram inquirimus.
HEB|13|15|Per ipsum ergo offeramus hostiam laudis semper Deo, id est fructum labiorum confitentium nomini eius.
HEB|13|16|Beneficientiae autem et communionis nolite oblivisci; talibus enim hostiis oblectatur Deus.
HEB|13|17|Oboedite praepositis vestris et subiacete eis; ipsi enim pervigilant pro animabus vestris quasi rationem reddituri, ut cum gaudio hoc faciant et non gementes; hoc enim non expedit vobis.
HEB|13|18|Orate pro nobis; confidimus enim quia bonam conscientiam habemus, in omnibus bene volentes conversari.
HEB|13|19|Amplius autem deprecor vos hoc facere, ut quo celerius restituar vobis.
HEB|13|20|Deus autem pacis, qui eduxit de mortuis pastorem magnum ovium in sanguine testamenti aeterni, Dominum nostrum Iesum,
HEB|13|21|aptet vos in omni bono, ut faciatis voluntatem eius, faciens in nobis, quod placeat coram se per Iesum Christum, cui gloria in saecula saeculorum. Amen.
HEB|13|22|Rogo autem vos, fratres, sufferte sermonem exhortationis; etenim perpaucis scripsi vobis.
HEB|13|23|Cognoscite fratrem nostrum Timotheum dimissum esse; cum quo, si celerius venerit, videbo vos.
HEB|13|24|Salutate omnes praepositos vestros et omnes sanctos. Salutant vos, qui de Italia sunt.
HEB|13|25|Gratia cum omnibus vobis.
JAS|1|1|Iacobus, Dei et Domini Iesu Christi servus, duodecim tribu bus, quae sunt in dispersione, salutem.
JAS|1|2|Omne gaudium existimate, fratres mei, cum in tentationibus variis incideritis,
JAS|1|3|scientes quod probatio fidei vestrae patientiam operatur;
JAS|1|4|patientia autem opus perfectum habeat, ut sitis perfecti et integri, in nullo deficientes.
JAS|1|5|Si quis autem vestrum indiget sapientia, postulet a Deo, qui dat omnibus affluenter et non improperat, et dabitur ei.
JAS|1|6|Postulet autem in fide nihil haesitans; qui enim haesitat, similis est fluctui maris, qui a vento movetur et circumfertur.
JAS|1|7|Non ergo aestimet homo ille quod accipiat aliquid a Domino,
JAS|1|8|vir duplex animo, inconstans in omnibus viis suis.
JAS|1|9|Glorietur autem frater humilis in exaltatione sua,
JAS|1|10|dives autem in humilitate sua, quoniam sicut flos feni transibit.
JAS|1|11|Exortus est enim sol cum ardore et arefecit fenum, et flos eius decidit, et decor vultus eius deperiit; ita et dives in itineribus suis marcescet.
JAS|1|12|Beatus vir, qui suffert tentationem, quia, cum probatus fuerit, accipiet coronam vitae, quam repromisit Deus diligentibus se.
JAS|1|13|Nemo, cum tentatur, dicat: " A Deo tentor "; Deus enim non tentatur malis, ipse autem neminem tentat.
JAS|1|14|Unusquisque vero tentatur a concupiscentia sua abstractus et illectus;
JAS|1|15|dein concupiscentia, cum conceperit, parit peccatum; peccatum vero, cum consummatum fuerit, generat mortem.
JAS|1|16|Nolite errare, fratres mei dilectissimi.
JAS|1|17|Omne datum optimum et omne donum perfectum de sursum est, descendens a Patre luminum, apud quem non est transmutatio nec vicissitudinis obumbratio.
JAS|1|18|Voluntarie genuit nos verbo veritatis, ut simus primitiae quaedam creaturae eius.
JAS|1|19|Scitis, fratres mei dilecti. Sit autem omnis homo velox ad audiendum, tardus autem ad loquendum et tardus ad iram;
JAS|1|20|ira enim viri iustitiam Dei non operatur.
JAS|1|21|Propter quod abicientes omnem immunditiam et abundantiam malitiae, in mansuetudine suscipite insitum verbum, quod potest salvare animas vestras.
JAS|1|22|Estote autem factores verbi et non auditores tantum fallentes vosmetipsos.
JAS|1|23|Quia si quis auditor est verbi et non factor, hic comparabitur viro consideranti vultum nativitatis suae in speculo;
JAS|1|24|consideravit enim se et abiit, et statim oblitus est qualis fuerit.
JAS|1|25|Qui autem perspexerit in lege perfecta libertatis et permanserit, non auditor obliviosus factus sed factor operis, hic beatus in facto suo erit.
JAS|1|26|Si quis putat se religiosum esse, non freno circumducens linguam suam sed seducens cor suum, huius vana est religio.
JAS|1|27|Religio munda et immaculata apud Deum et Patrem haec est: visitare pupillos et viduas in tribulatione eorum, immaculatum se custodire ab hoc saeculo.
JAS|2|1|Fratres mei, nolite in persona rum acceptione habere fidem Domini nostri Iesu Christi gloriae.
JAS|2|2|Etenim, si introierit in synagogam vestram vir aureum anulum habens in veste candida, introierit autem et pauper in sordido habitu,
JAS|2|3|et intendatis in eum, qui indutus est veste praeclara, et dixeritis: " Tu sede hic bene ", pauperi autem dicatis: " Tu sta illic aut sede sub scabello meo ";
JAS|2|4|nonne iudicatis apud vosmetipsos et facti estis iudices cogitationum iniquarum?
JAS|2|5|Audite, fratres mei dilectissimi. Nonne Deus elegit, qui pauperes sunt mundo, divites in fide et heredes regni, quod repromisit diligentibus se?
JAS|2|6|Vos autem exhonorastis pauperem. Nonne divites opprimunt vos et ipsi trahunt vos ad iudicia?
JAS|2|7|Nonne ipsi blasphemant bonum nomen, quod invocatum est super vos?
JAS|2|8|Si tamen legem perficitis regalem secundum Scripturam: " Diliges proximum tuum sicut teipsum ", bene facitis;
JAS|2|9|si autem personas accipitis, peccatum operamini, redarguti a lege quasi transgressores.
JAS|2|10|Quicumque autem totam legem servaverit, offendat autem in uno, factus est omnium reus.
JAS|2|11|Qui enim dixit: " Non moechaberis ", dixit et: " Non occides "; quod si non moecharis, occidis autem, factus es transgressor legis.
JAS|2|12|Sic loquimini et sic facite sicut per legem libertatis iudicandi.
JAS|2|13|Iudicium enim sine misericordia illi, qui non fecit misericordiam; superexsultat misericordia iudicio.
JAS|2|14|Quid proderit, fratres mei, si fidem quis dicat se habere, opera autem non habeat? Numquid poterit fides salvare eum?
JAS|2|15|Si frater aut soror nudi sunt et indigent victu cotidiano,
JAS|2|16|dicat autem aliquis de vobis illis: " Ite in pace, calefacimini et saturamini ", non dederitis autem eis, quae necessaria sunt corporis, quid proderit?
JAS|2|17|Sic et fides, si non habeat opera, mortua est in semetipsa.
JAS|2|18|Sed dicet quis: " Tu fidem habes, et ego opera habeo ". Ostende mihi fidem tuam sine operibus, et ego tibi ostendam ex operibus meis fidem.
JAS|2|19|Tu credis quoniam unus est Deus? Bene facis; et daemones credunt et contremiscunt!
JAS|2|20|Vis autem scire, o homo inanis, quoniam fides sine operibus otiosa est?
JAS|2|21|Abraham, pater noster, nonne ex operibus iustificatus est offerens Isaac filium suum super altare?
JAS|2|22|Vides quoniam fides cooperabatur operibus illius, et ex operibus fides consummata est;
JAS|2|23|et suppleta est Scriptura dicens: " Credidit Abraham Deo, et reputatum est illi ad iustitiam ", et amicus Dei appellatus est.
JAS|2|24|Videtis quoniam ex operibus iustificatur homo et non ex fide tantum.
JAS|2|25|Similiter autem et Rahab, meretrix nonne ex operibus iustificata est suscipiens nuntios et alia via eiciens?
JAS|2|26|Sicut enim corpus sine spiritu emortuum est, ita et fides sine operibus mortua est.
JAS|3|1|Nolite plures magistri fieri, fra tres mei, scientes quoniam maius iudicium accipiemus.
JAS|3|2|In multis enim offendimus omnes. Si quis in verbo non offendit, hic perfectus est vir, potens etiam freno circumducere totum corpus.
JAS|3|3|Si autem equorum frenos in ora mittimus ad oboediendum nobis, et omne corpus illorum circumferimus.
JAS|3|4|Ecce et naves, cum tam magnae sint et a ventis validis minentur, circumferuntur a minimo gubernaculo, ubi impetus dirigentis voluerit;
JAS|3|5|ita et lingua modicum quidem membrum est et magna exsultat. Ecce quantus ignis quam magnam silvam incendit!
JAS|3|6|Et lingua ignis est, universitas iniquitatis; lingua constituitur in membris nostris, quae maculat totum corpus et inflammat rotam nativitatis et inflammatur a gehenna.
JAS|3|7|Omnis enim natura et bestiarum et volucrum et serpentium et etiam cetorum domatur et domita est a natura humana;
JAS|3|8|linguam autem nullus hominum domare potest, inquietum malum, plena veneno mortifero.
JAS|3|9|In ipsa benedicimus Dominum et Patrem et in ipsa maledicimus homines, qui ad similitudinem Dei facti sunt;
JAS|3|10|ex ipso ore procedit benedictio et maledictio. Non oportet, fratres mei, haec ita fieri.
JAS|3|11|Numquid fons de eodem foramine emanat dulcem et amaram aquam?
JAS|3|12|Numquid potest, fratres mei, ficus olivas facere, aut vitis ficus? Neque salsa dulcem potest facere aquam.
JAS|3|13|Quis sapiens et disciplinatus inter vos? Ostendat ex bona conversatione operationem suam in mansuetudine sapientiae.
JAS|3|14|Quod si zelum amarum habetis et contentiones in cordibus vestris, nolite gloriari et mendaces esse adversus veritatem.
JAS|3|15|Non est ista sapientia desursum descendens, sed terrena, animalis, diabolica;
JAS|3|16|ubi enim zelus et contentio, ibi inconstantia et omne opus pravum.
JAS|3|17|Quae autem desursum est sapientia primum quidem pudica est, deinde pacifica, modesta, suadibilis, plena misericordia et fructibus bonis, non iudicans, sine simulatione;
JAS|3|18|fructus autem iustitiae in pace seminatur facientibus pacem.
JAS|4|1|Unde bella et unde lites in vobis? Nonne hinc, ex concupi scentiis vestris, quae militant in membris vestris?
JAS|4|2|Concupiscitis et non habetis; occiditis et zelatis et non potestis adipisci; litigatis et belligeratis. Non habetis, propter quod non postulatis;
JAS|4|3|petitis et non accipitis, eo quod male petitis, ut in concupiscentiis vestris insumatis.
JAS|4|4|Adulteri, nescitis quia amicitia huius mundi inimica est Dei?Quicumque ergo voluerit amicus esse saeculi huius, inimicus Dei constituitur.
JAS|4|5|Aut putatis quia inaniter Scriptura dicat: " Ad invidiam concupiscit Spiritus, qui inhabitat in nobis? ".
JAS|4|6|Maiorem autem dat gratiam; propter quod dicit: Deus superbis resistit,humilibus autem dat gratiam ".
JAS|4|7|Subicimini igitur Deo; resistite autem Diabolo, et fugiet a vobis.
JAS|4|8|Appropiate Deo, et appropinquabit vobis. Emundate manus, peccatores; et purificate corda, duplices animo.
JAS|4|9|Miseri estote et lugete et plorate; risus vester in luctum convertatur, et gaudium in maerorem.
JAS|4|10|Humiliamini in conspectu Domini, et exaltabit vos.
JAS|4|11|Nolite detrahere alterutrum, fratres; qui detrahit fratri, aut qui iudicat fratrem suum, detrahit legi et iudicat legem; si autem iudicas legem, non es factor legis sed iudex.
JAS|4|12|Unus est legislator et iudex, qui potest salvare et perdere; tu autem quis es, qui iudicas proximum?
JAS|4|13|Age nunc, qui dicitis: " Hodie aut crastino ibimus in illam civitatem et faciemus quidem ibi annum et mercabimur et lucrum faciemus ";
JAS|4|14|qui ignoratis, quae erit in crastinum vita vestra! Vapor enim estis ad modicum parens, deinceps exterminatur;
JAS|4|15|pro eo ut dicatis: " Si Dominus voluerit, et vivemus et faciemus hoc aut illud ".
JAS|4|16|Nunc autem gloriamini in superbiis vestris; omnis gloriatio talis maligna est.
JAS|4|17|Scienti igitur bonum facere et non facienti, peccatum est illi!
JAS|5|1|Age nunc, divites, plorate ulu lantes in miseriis, quae adve nient vobis.
JAS|5|2|Divitiae vestrae putrefactae sunt, et vestimenta vestra a tineis comesta sunt,
JAS|5|3|aurum et argentum vestrum aeruginavit, et aerugo eorum in testimonium vobis erit et manducabit carnes vestras sicut ignis: thesaurizastis in novissimis diebus.
JAS|5|4|Ecce merces operariorum, qui messuerunt regiones vestras, quae fraudata est a vobis, clamat, et clamores eorum, qui messuerunt, in aures Domini Sabaoth introierunt.
JAS|5|5|Epulati estis super terram et in luxuriis fuistis, enutristis corda vestra in die occisionis.
JAS|5|6|Addixistis, occidistis iustum. Non resistit vobis.
JAS|5|7|Patientes igitur estote, fratres, usque ad adventum Domini. Ecce agricola exspectat pretiosum fructum terrae, patienter ferens, donec accipiat imbrem temporaneum et serotinum.
JAS|5|8|Patientes estote, et vos, confirmate corda vestra, quoniam adventus Domini appropinquavit.
JAS|5|9|Nolite ingemiscere, fratres, in alterutrum, ut non iudicemini; ecce iudex ante ianuam assistit.
JAS|5|10|Exemplum accipite, fratres, laboris et patientiae prophetas, qui locuti sunt in nomine Domini.
JAS|5|11|Ecce beatificamus eos, qui sustinuerunt; sufferentiam Iob audistis et finem Domini vidistis, quoniam misericors est Dominus et miserator.
JAS|5|12|Ante omnia autem, fratres mei, nolite iurare neque per caelum neque per terram, neque aliud quodcumque iuramentum; sit autem vestrum " Est " est, et " Non " non, uti non sub iudicio decidatis.
JAS|5|13|Tristatur aliquis vestrum? Oret. Aequo animo est? Psallat.
JAS|5|14|Infirmatur quis in vobis? Advocet presbyteros ecclesiae, et orent super eum, unguentes eum oleo in nomine Domini.
JAS|5|15|Et oratio fidei salvabit infirmum, et allevabit eum Dominus; et si peccata operatus fuerit, dimittentur ei.
JAS|5|16|Confitemini ergo alterutrum peccata et orate pro invicem, ut sanemini. Multum enim valet deprecatio iusti operans.
JAS|5|17|Elias homo erat similis nobis passibilis et oratione oravit, ut non plueret, et non pluit super terram annos tres et menses sex;
JAS|5|18|et rursum oravit, et caelum dedit pluviam, et terra germinavit fructum suum.
JAS|5|19|Fratres mei, si quis ex vobis erraverit a veritate, et converterit quis eum,
JAS|5|20|scire debet quoniam, qui converti fecerit peccatorem ab errore viae eius, salvabit animam suam a morte et operiet multitudinem peccatorum.
1PET|1|1|Petrus apostolus Iesu Christi electis advenis dispersionis Pon ti, Galatiae, Cappadociae, Asiae et Bithyniae,
1PET|1|2|secundum praescientiam Dei Patris, in sanctificatione Spiritus, in oboedientiam et aspersionem sanguinis Iesu Christi: gratia vobis et pax multiplicetur.
1PET|1|3|Benedictus Deus et Pater Domini nostri Iesu Christi, qui secundum magnam misericordiam suam regeneravit nos in spem vivam per resurrectionem Iesu Christi ex mortuis,
1PET|1|4|in hereditatem incorruptibilem et incontaminatam et immarcescibilem, conservatam in caelis propter vos,
1PET|1|5|qui in virtute Dei custodimini per fidem in salutem, paratam revelari in tempore novissimo.
1PET|1|6|In quo exsultatis, modicum nunc si oportet contristati in variis tentationibus,
1PET|1|7|ut probatio vestrae fidei multo pretiosior auro, quod perit, per ignem quidem probato, inveniatur in laudem et gloriam et honorem in revelatione Iesu Christi.
1PET|1|8|Quem cum non videritis, diligitis; in quem nunc non videntes, credentes autem, exsultatis laetitia inenarrabili et glorificata,
1PET|1|9|reportantes finem fidei vestrae salutem animarum.
1PET|1|10|De qua salute exquisierunt atque scrutati sunt prophetae, qui de futura in vos gratia prophetaverunt,
1PET|1|11|scrutantes in quod vel quale tempus significaret, qui erat in eis Spiritus Christi, praenuntians eas, quae in Christo sunt, passiones et posteriores glorias;
1PET|1|12|quibus revelatum est quia non sibi ipsis, vobis autem ministrabant ea, quae nunc nuntiata sunt vobis per eos, qui evangelizaverunt vos, Spiritu Sancto misso de caelo, in quae desiderant angeli prospicere.
1PET|1|13|Propter quod succincti lumbos mentis vestrae, sobrii, perfecte sperate in eam, quae offertur vobis, gratiam in revelatione Iesu Christi.
1PET|1|14|Quasi filii oboedientiae, non configurati prioribus in ignorantia vestra desideriis,
1PET|1|15|sed secundum eum, qui vocavit vos, sanctum, et ipsi sancti in omni conversatione sitis,
1PET|1|16|quoniam scriptum est: " Sancti eritis, quia ego sanctus sum ".
1PET|1|17|Et si Patrem invocatis eum, qui sine acceptione personarum iudicat secundum uniuscuiusque opus, in timore incolatus vestri tempore conversamini,
1PET|1|18|scientes quod non corruptibilibus argento vel auro redempti estis de vana vestra conversatione a patribus tradita,
1PET|1|19|sed pretioso sanguine quasi Agni incontaminati et immaculati Christi,
1PET|1|20|praecogniti quidem ante constitutionem mundi, manifestati autem novissimis temporibus propter vos,
1PET|1|21|qui per ipsum fideles estis in Deum, qui suscitavit eum a mortuis et dedit ei gloriam, ut fides vestra et spes esset in Deum.
1PET|1|22|Animas vestras castificantes in oboedientia veritatis ad fraternitatis amorem non fictum, ex corde invicem diligite attentius,
1PET|1|23|renati non ex semine corruptibili sed incorruptibili per verbum Dei vivum et permanens:
1PET|1|24|quiaomnis caro ut fenum,et omnis gloria eius tamquam flos feni.Exaruit fenum, et flos decidit;
1PET|1|25|verbum autem Domini manet in aeternum.Hoc est autem verbum, quod evangelizatum est in vos.
1PET|2|1|Deponentes igitur omnem ma litiam et omnem dolum et simu lationes et invidias et omnes detractiones,
1PET|2|2|sicut modo geniti infantes, rationale sine dolo lac concupiscite, ut in eo crescatis in salutem,
1PET|2|3|si gustastis quoniam dulcis Dominus.
1PET|2|4|Ad quem accedentes, lapidem vivum, ab hominibus quidem reprobatum, coram Deo autem electum, pretiosum,
1PET|2|5|et ipsi tamquam lapides vivi aedificamini domus spiritalis in sacerdotium sanctum offerre spiritales hostias acceptabiles Deo per Iesum Christum.
1PET|2|6|Propter quod continet Scriptura: Ecce pono in Sion lapidem angularem, electum, pretiosum;et, qui credit in eo, non confundetur ".
1PET|2|7|Vobis igitur honor credentibus; non credentibus autem Lapis, quem reprobaverunt aedificantes, hic factus est in caput anguli "
1PET|2|8|et " lapis offensionis et petra scandali "; qui offendunt verbo non credentes, in quod et positi sunt.
1PET|2|9|Vos autem genus electum, regale sacerdotium, gens sancta, populus in acquisitionem, ut virtutes annuntietis eius, qui de tenebris vos vocavit in admirabile lumen suum:
1PET|2|10|qui aliquando non populus, nunc autem populus Dei; qui non consecuti misericordiam, nunc autem misericordiam consecuti.
1PET|2|11|Carissimi, obsecro tamquam advenas et peregrinos abstinere vos a carnalibus desideriis, quae militant adversus animam;
1PET|2|12|conversationem vestram inter gentes habentes bonam, ut in eo, quod detrectant de vobis tamquam de malefactoribus, ex bonis operibus considerantes glorificent Deum in die visitationis.
1PET|2|13|Subiecti estote omni humanae creaturae propter Dominum: sive regi quasi praecellenti
1PET|2|14|sive ducibus tamquam ab eo missis ad vindictam malefactorum, laudem vero bonorum;
1PET|2|15|quia sic est voluntas Dei, ut benefacientes obmutescere faciatis imprudentium hominum ignorantiam,
1PET|2|16|quasi liberi, et non quasi velamen habentes malitiae libertatem, sed sicut servi Dei.
1PET|2|17|Omnes honorate, fraternitatem diligite, Deum timete, regem honorificate.
1PET|2|18|Servi, subditi estote in omni timore dominis, non tantum bonis et modestis sed etiam pravis.
1PET|2|19|Haec est enim gratia, si propter conscientiam Dei sustinet quis tristitias, patiens iniuste.
1PET|2|20|Quae enim gloria est, si peccantes et colaphizati sustinetis? Sed si benefacientes et patientes sustinetis, haec est gratia apud Deum.
1PET|2|21|In hoc enim vocati estis, quiaet Christus passus est pro vobis,vobis relinquens exemplum,ut sequamini vestigia eius:
1PET|2|22|qui peccatum non fecit,nec inventus est dolus in ore ipsius;
1PET|2|23|qui cum malediceretur, non remaledicebat;cum pateretur, non comminabatur, commendabat autem iuste iudicanti;
1PET|2|24|qui peccata nostra ipse pertulitin corpore suo super lignum,ut peccatis mortui iustitiae viveremus;cuius livore sanati estis.
1PET|2|25|Eratis enim sicut oves errantes,sed conversi estis nunc ad pastorem et episcopum animarum vestrarum.
1PET|3|1|Similiter mulieres subditae sint suis viris, ut et si qui non cre dunt verbo, per mulierum conversationem sine verbo lucrifiant,
1PET|3|2|considerantes castam in timore conversationem vestram;
1PET|3|3|quarum sit non extrinsecus capillaturae aut circumdationis auri aut indumenti vestimentorum cultus,
1PET|3|4|sed qui absconditus cordis est homo, in incorruptibilitate mitis et quieti spiritus, qui est in conspectu Dei locuples.
1PET|3|5|Sic enim aliquando et sanctae mulieres sperantes in Deo ornabant se subiectae propriis viris,
1PET|3|6|sicut Sara oboediebat Abrahae dominum eum vocans: cuius estis filiae benefacientes et non timentes ullam perturbationem.
1PET|3|7|Viri similiter cohabitantes secundum scientiam quasi infirmiori vaso muliebri impertientes honorem, tamquam et coheredibus gratiae vitae, uti ne impediantur orationes vestrae.
1PET|3|8|In fine autem omnes unanimes, compatientes, fraternitatis amatores, misericordes, humiles,
1PET|3|9|non reddentes malum pro malo vel maledictum pro maledicto, sed e contrario benedicentes, quia in hoc vocati estis, ut benedictionem hereditate accipiatis.
1PET|3|10|" Qui enim vult vitam diligereet videre dies bonos,coerceat linguam suam a malo,
1PET|3|11|et labia eius ne loquantur dolum;declinet autem a malo et faciat bonum,inquirat pacem et persequatur eam.
1PET|3|12|Quia oculi Domini super iustos,et aures eius in preces eorum;vultus autem Domini super facientes mala ".
1PET|3|13|Et quis est qui vobis noceat, si boni aemulatores fueritis?
1PET|3|14|Sed et si patimini propter iustitiam, beati! Timorem autem eorum ne timueritis et non conturbemini,
1PET|3|15|Dominum autem Christum sanctificate in cordibus vestris, parati semper ad defensionem omni poscenti vos rationem de ea, quae in vobis est spe;
1PET|3|16|sed cum mansuetudine et timore, conscientiam habentes bonam, ut in quo de vobis detrectatur, confundantur, qui calumniantur vestram bonam in Christo conversationem.
1PET|3|17|Melius est enim benefacientes, si velit voluntas Dei, pati quam malefacientes.
1PET|3|18|Quia et Christus semel pro peccatis passus est, iustus pro iniustis, ut vos adduceret ad Deum, mortificatus quidem carne, vivificatus autem Spiritu:
1PET|3|19|in quo et his, qui in carcere erant, spiritibus adveniens praedicavit,
1PET|3|20|qui increduli fuerant aliquando, quando exspectabat Dei patientia in diebus Noe, cum fabricaretur arca, in qua pauci, id est octo animae, salvae factae sunt per aquam.
1PET|3|21|Cuius antitypum, baptisma, et vos nunc salvos facit, non carnis depositio sordium sed conscientiae bonae rogatio in Deum, per resurrectionem Iesu Christi,
1PET|3|22|qui est in dextera Dei, profectus in caelum, subiectis sibi angelis et potestatibus et virtutibus.
1PET|4|1|Christo igitur passo in carne, et vos eadem cogitatione armami ni, quia, qui passus est carne, desiit a peccato;
1PET|4|2|ut iam non hominum concupiscentiis sed voluntate Dei, quod reliquum est in carne vivat temporis.
1PET|4|3|Sufficit enim praeteritum tempus ad voluntatem gentium consummandam, vobis, qui ambulastis in luxuriis, concupiscentiis, vinolentiis, comissationibus, potationibus et illicitis idolorum cultibus.
1PET|4|4|In quo mirantur non concurrentibus vobis in eandem luxuriae effusionem, blasphemantes;
1PET|4|5|qui reddent rationem ei, qui paratus est iudicare vivos et mortuos.
1PET|4|6|Propter hoc enim et mortuis evangelizatum est, ut iudicentur quidem secundum homines carne, vivant autem secundum Deum Spiritu.
1PET|4|7|Omnium autem finis appropinquavit. Estote itaque prudentes et vigilate in orationibus.
1PET|4|8|Ante omnia mutuam in vosmetipsos caritatem continuam habentes, quia caritas operit multitudinem peccatorum;
1PET|4|9|hospitales invicem sine murmuratione;
1PET|4|10|unusquisque, sicut accepit donationem, in alterutrum illam administrantes, sicut boni dispensatores multiformis gratiae Dei.
1PET|4|11|Si quis loquitur, quasi sermones Dei; si quis ministrat, tamquam ex virtute, quam largitur Deus, ut in omnibus glorificetur Deus per Iesum Christum: cui est gloria et imperium in saecula saeculorum. Amen.
1PET|4|12|Carissimi, nolite mirari in fervore, qui ad tentationem vobis fit, quasi novi aliquid vobis contingat,
1PET|4|13|sed, quemadmodum communicatis Christi passionibus, gaudete, ut et in revelatione gloriae eius gaudeatis exsultantes.
1PET|4|14|Si exprobramini in nomine Christi, beati, quoniam Spiritus gloriae et Dei super vos requiescit.
1PET|4|15|Nemo enim vestrum patiatur quasi homicida aut fur aut maleficus aut alienorum speculator;
1PET|4|16|si autem ut christianus, non erubescat, glorificet autem Deum in isto nomine.
1PET|4|17|Quoniam tempus est, ut incipiat iudicium a domo Dei; si autem primum a nobis, qui finis eorum, qui non credunt Dei evangelio?
1PET|4|18|" Et si iustus vix salvatur,impius et peccator ubi parebit? ".
1PET|4|19|Itaque et hi, qui patiuntur secundum voluntatem Dei, fideli Creatori commendent animas suas in benefacto.
1PET|5|1|Seniores ergo, qui in vobis sunt, obsecro, consenior et testis Chri sti passionum, qui et eius, quae in futuro revelanda est, gloriae communicator:
1PET|5|2|Pascite, qui est in vobis, gregem Dei, providentes non coacto sed spontanee secundum Deum, neque turpis lucri gratia sed voluntarie,
1PET|5|3|neque ut dominantes in cleris sed formae facti gregis.
1PET|5|4|Et cum apparuerit Princeps pastorum, percipietis immarcescibilem gloriae coro nam.
1PET|5|5|Similiter, adulescentes, subditi estote senioribus. Omnes autem invicem humilitatem induite, quiaDeus superbis resistit,humilibus autem dat gratiam.
1PET|5|6|Humiliamini igitur sub potenti manu Dei, ut vos exaltet in tempore,
1PET|5|7|omnem sollicitudinem vestram proicientes in eum, quoniam ipsi cura est de vobis.
1PET|5|8|Sobrii estote, vigilate. Adversarius vester Diabolus tamquam leo rugiens circuit quaerens quem devoret.
1PET|5|9|Cui resistite fortes fide, scientes eadem passionum ei, quae in mundo est, vestrae fraternitati fieri.
1PET|5|10|Deus autem omnis gratiae, qui vocavit vos in aeternam suam gloriam in Christo Iesu, modicum passos ipse perficiet, confirmabit, solidabit, fundabit.
1PET|5|11|Ipsi imperium in saecula saeculorum. Amen.
1PET|5|12|Per Silvanum vobis fidelem fratrem, ut arbitror, breviter scripsi, obsecrans et contestans hanc esse veram gratiam Dei; in qua state.
1PET|5|13|Salutat vos, quae est in Babylone, coelecta et Marcus filius meus.
1PET|5|14|Salutate invicem in osculo caritatis.Pax vobis omnibus, qui estis in Christo.
2PET|1|1|Simon Petrus servus et apo stolus Iesu Christi his, qui coae qualem nobis sortiti sunt fidem in iustitia Dei nostri et salvatoris Iesu Christi:
2PET|1|2|gratia vobis et pax multiplicetur in cognitione Dei et Iesu Domini nostri.
2PET|1|3|Quomodo omnia nobis divinae virtutis suae ad vitam et pietatem donatae per cognitionem eius, qui vocavit nos propria gloria et virtute,
2PET|1|4|per quae pretiosa et maxima nobis promissa donata sunt, ut per haec efficiamini divinae consortes naturae, fugientes eam, quae in mundo est in concupiscentia, corruptionem;
2PET|1|5|et propter hoc ipsum curam omnem subinferentes ministrate in fide vestra virtutem, in virtute autem scientiam,
2PET|1|6|in scientia autem continentiam, in continentia autem patientiam, in patientia autem pietatem,
2PET|1|7|in pietate autem amorem fraternitatis, in amore autem fraternitatis caritatem.
2PET|1|8|Haec enim vobis, cum adsint et abundent, non vacuos nec sine fructu vos constituunt in Domini nostri Iesu Christi cognitionem;
2PET|1|9|cui enim non praesto sunt haec, caecus est et nihil procul cernens, oblivionem accipiens purgationis veterum suorum delictorum.
2PET|1|10|Quapropter, fratres, magis satagite, ut firmam vestram vocationem et electionem faciatis. Haec enim facientes non offendetis aliquando;
2PET|1|11|sic enim abundanter ministrabitur vobis introitus in aeternum regnum Domini nostri et salvatoris Iesu Christi.
2PET|1|12|Propter quod incipiam vos semper commonere de his, et quidem scientes et confirmatos in praesenti veritate.
2PET|1|13|Iustum autem arbitror, quamdiu sum in hoc tabernaculo, suscitare vos in commonitione,
2PET|1|14|certus quod velox est depositio tabernaculi mei, secundum quod et Dominus noster Iesus Christus significavit mihi;
2PET|1|15|dabo autem operam et frequenter habere vos post obitum meum, ut horum memoriam faciatis.
2PET|1|16|Non enim captiosas fabulas secuti notam fecimus vobis Domini nostri Iesu Christi virtutem et adventum, sed speculatores facti illius magnitudinis.
2PET|1|17|Accipiens enim a Deo Patre honorem et gloriam, voce prolata ad eum huiuscemodi a magnifica gloria: " Filius meus, dilectus meus hic est, in quo ego mihi complacui ";
2PET|1|18|et hanc vocem nos audivimus de caelo prolatam, cum essemus cum ipso in monte sancto.
2PET|1|19|Et habemus firmiorem propheticum sermonem, cui bene facitis attendentes quasi lucernae lucenti in caliginoso loco, donec dies illucescat, et lucifer oriatur in cordibus vestris,
2PET|1|20|hoc primum intellegentes quod omnis prophetia Scripturae propria interpretatione non fit;
2PET|1|21|non enim voluntate humana prolata est prophetia aliquando, sed a Spiritu Sancto ducti locuti sunt a Deo homines.
2PET|2|1|Fuerunt vero et pseudopro phetae in populo, sicut et in vo bis erunt magistri mendaces, qui introducent sectas perditionis et eum, qui emit eos, Dominatorem negantes superducent sibi celerem perditionem.
2PET|2|2|Et multi sequentur eorum luxurias, propter quos via veritatis blasphemabitur;
2PET|2|3|et in avaritia fictis verbis de vobis negotiabuntur. Quibus iudicium iam olim non cessat, et perditio eorum non dormitat.
2PET|2|4|Si enim Deus angelis peccantibus non pepercit, sed rudentibus inferni detractos in tartarum tradidit in iudicium reservatos:
2PET|2|5|et originali mundo non pepercit, sed octavum Noe iustitiae praeconem custodivit diluvium mundo impiorum inducens;
2PET|2|6|et civitates Sodomae et Gomorrae in cinerem redigens eversione damnavit, exemplum ponens eorum, quae sunt impiis futura:
2PET|2|7|et iustum Lot oppressum a nefandorum luxuria conversationis eruit:
2PET|2|8|aspectu enim et auditu iustus habitans apud eos, de die in diem animam iustam iniquis operibus cruciabat.
2PET|2|9|Novit Dominus pios de tentatione eripere, iniquos vero in diem iudicii puniendos reservare,
2PET|2|10|maxime autem eos, qui post carnem in concupiscentia immunditiae ambulant dominationemque contemnunt.Audaces, superbi, glorias non metuunt blasphemantes,
2PET|2|11|ubi angeli fortitudine et virtute cum sint maiores, non portant adversum illas coram Domino iudicium blasphemiae.
2PET|2|12|Hi vero, velut irrationabilia animalia naturaliter genita in captionem et in corruptionem, in his, quae ignorant, blasphemantes, in corruptione sua et corrumpentur
2PET|2|13|inviti percipientes mercedem iniustitiae; voluptatem existimantes diei delicias, coinquinationes et maculae deliciis affluentes, in voluptatibus suis luxuriantes vobiscum,
2PET|2|14|oculos habentes plenos adulterae et incessabiles delicti, pellicientes animas instabiles, cor exercitatum avaritiae habentes, maledictionis filii;
2PET|2|15|derelinquentes rectam viam erraverunt, secuti viam Balaam ex Bosor, qui mercedem iniquitatis amavit,
2PET|2|16|correptionem vero habuit suae praevaricationis; subiugale mutum in hominis voce loquens prohibuit prophetae insipientiam.
2PET|2|17|Hi sunt fontes sine aqua, et nebulae turbine exagitatae, quibus caligo tenebrarum reservatur.
2PET|2|18|Superba enim vanitatis loquentes pelliciunt in concupiscentiis carnis luxuriis illos, qui paululum effugiunt eos, qui in errore conversantur,
2PET|2|19|libertatem illis promittentes, cum ipsi servi sint corruptionis; a quo enim quis superatus est, huius servus est.
2PET|2|20|Si enim refugientes coinquinationes mundi in cognitione Domini nostri et Salvatoris Iesu Christi his rursus implicati superantur, facta sunt eis posteriora deteriora prioribus.
2PET|2|21|Melius enim erat illis non cognoscere viam iustitiae, quam post agnitionem retrorsum converti ab eo, quod illis traditum est, sancto mandato.
2PET|2|22|Contigit enim eis illud veri proverbii: Canis reversus ad suum vomitum ",et " Sus lota in volutabro luti ".
2PET|3|1|Hanc vobis, carissimi, iam se cundam scribo epistulam, in quibus excito vestram in commonitione sinceram mentem,
2PET|3|2|ut memores sitis eorum, quae praedicta sunt verborum a sanctis prophetis, et ab apostolis traditi vobis praecepti Domini et Salvatoris;
2PET|3|3|hoc primum scientes, quod venient in novissimis diebus in illusione illudentes, iuxta proprias concupiscentias suas ambulantes,
2PET|3|4|dicentes: " Ubi est promissio adventus eius? Ex quo enim patres dormierunt, omnia sic perseverant ab initio creaturae ".
2PET|3|5|Latet enim eos hoc volentes, quod caeli erant prius, et terra de aqua et per aquam consistens Dei verbo,
2PET|3|6|per quae ille tunc mundus aqua inundatus periit;
2PET|3|7|caeli autem, qui nunc sunt, et terra eodem verbo repositi sunt igni, servati in diem iudicii et perditionis impiorum hominum.
2PET|3|8|Unum vero hoc non lateat vos, carissimi, quia unus dies apud Dominum sicut mille anni, et mille anni sicut dies unus.
2PET|3|9|Non tardat Dominus promissionem, sicut quidam tarditatem existimant, sed patienter agit in vos nolens aliquos perire, sed omnes ad paenitentiam reverti.
2PET|3|10|Adveniet autem dies Domini ut fur, in qua caeli magno impetu transient, elementa vero calore solventur, et terra et opera, quae in ea invenientur.
2PET|3|11|Cum haec omnia ita dissolvenda sint, quales oportet esse vos in sanctis conversationibus et pietatibus,
2PET|3|12|exspectantes et properantes adventum diei Dei, propter quam caeli ardentes solventur, et elementa ignis ardore tabescent!
2PET|3|13|Novos vero caelos et terram novam secundum promissum ipsius exspectamus, in quibus iustitia habitat.
2PET|3|14|Propter quod, carissimi, haec exspectantes satagite immaculati et inviolati ei inveniri in pace;
2PET|3|15|et Domini nostri longanimitatem, salutem arbitramini, sicut et carissimus frater noster Paulus secundum datam sibi sapientiam scripsit vobis,
2PET|3|16|sicut et in omnibus epistulis loquens in eis de his; in quibus sunt quaedam difficilia intellectu, quae indocti et instabiles depravant, sicut et ceteras Scripturas, ad suam ipsorum perditionem.
2PET|3|17|Vos igitur, dilecti, praescientes custodite, ne iniquorum errore simul abducti excidatis a propria firmitate;
2PET|3|18|crescite vero in gratia et in cognitione Domini nostri et Salvatoris Iesu Christi. Ipsi gloria et nunc et in diem aeternitatis. Amen.
1JOHN|1|1|Quod fuit ab initio, quod audi vimus, quod vidimus oculis no stris, quod perspeximus, et manus nostrae contrectaverunt de verbo vitae
1JOHN|1|2|- et vita apparuit, et vidimus et testamur et annuntiamus vobis vitam aeternam, quae erat coram Patre et apparuit nobis -
1JOHN|1|3|quod vidimus et audivimus, annuntiamus et vobis, ut et vos communionem habeatis nobiscum. Communio autem nostra est cum Patre et cum Filio eius Iesu Christo.
1JOHN|1|4|Et haec scribimus nos, ut gaudium nostrum sit plenum.
1JOHN|1|5|Et haec est annuntiatio, quam audivimus ab eo et annuntiamus vobis, quoniam Deus lux est, et tenebrae in eo non sunt ullae.
1JOHN|1|6|Si dixerimus quoniam communionem habemus cum eo, et in tenebris ambulamus, mentimur et non facimus veritatem;
1JOHN|1|7|si autem in luce ambulemus, sicut ipse est in luce, communionem habemus ad invicem, et sanguis Iesu Filii eius mundat nos ab omni peccato.
1JOHN|1|8|Si dixerimus quoniam peccatum non habemus, nosmetipsos seducimus, et veritas in nobis non est.
1JOHN|1|9|Si confiteamur peccata nostra, fidelis est et iustus, ut remittat nobis peccata et emundet nos ab omni iniustitia.
1JOHN|1|10|Si dixerimus quoniam non peccavimus, mendacem facimus eum, et verbum eius non est in nobis.
1JOHN|2|1|Filioli mei, haec scribo vobis, ut non peccetis. Sed si quis pecca verit, advocatum habemus ad Patrem, Iesum Christum iustum;
1JOHN|2|2|et ipse est propitiatio pro peccatis nostris, non pro nostris autem tantum sed etiam pro totius mundi.
1JOHN|2|3|Et in hoc cognoscimus quoniam novimus eum: si mandata eius servemus.
1JOHN|2|4|Qui dicit: " Novi eum ", et mandata eius non servat, mendax est, et in isto veritas non est;
1JOHN|2|5|qui autem servat verbum eius, vere in hoc caritas Dei consummata est. In hoc cognoscimus quoniam in ipso sumus.
1JOHN|2|6|Qui dicit se in ipso manere, debet, sicut ille ambulavit, et ipse ambulare.
1JOHN|2|7|Carissimi, non mandatum novum scribo vobis sed mandatum vetus, quod habuistis ab initio: mandatum vetus est verbum, quod audistis.
1JOHN|2|8|Verumtamen mandatum novum scribo vobis, quod est verum in ipso et in vobis, quoniam tenebrae transeunt, et lumen verum iam lucet.
1JOHN|2|9|Qui dicit se in luce esse, et fratrem suum odit, in tenebris est usque adhuc.
1JOHN|2|10|Qui diligit fratrem suum, in lumine manet, et scandalum ei non est;
1JOHN|2|11|qui autem odit fratrem suum, in tenebris est et in tenebris ambulat et nescit quo vadat, quoniam tenebrae obcaecaverunt oculos eius.
1JOHN|2|12|Scribo vobis, filioli: Remissa sunt vobis peccata propter nomen eius.
1JOHN|2|13|Scribo vobis, patres: Nostis eum, qui ab initio est. Scribo vobis, adulescentes: Vicistis Malignum.
1JOHN|2|14|Scripsi vobis, parvuli: Nostis Patrem. Scripsi vobis, patres: Nostis eum, qui ab initio est. Scripsi vobis, adulescentes: Fortes estis, et verbum Dei in vobis manet, et vicistis Malignum.
1JOHN|2|15|Nolite diligere mundum neque ea, quae in mundo sunt. Si quis diligit mundum, non est caritas Patris in eo;
1JOHN|2|16|quoniam omne, quod est in mundo, concupiscentia carnis et concupiscentia oculorum et iactantia divitiarum, non est ex Patre, sed ex mundo est.
1JOHN|2|17|Et mundus transit, et concupiscentia eius; qui autem facit voluntatem Dei, manet in aeternum.
1JOHN|2|18|Filioli, novissima hora est; et sicut audistis quia antichristus venit, ita nunc antichristi multi adsunt, unde cognoscimus quoniam novissima hora est.
1JOHN|2|19|Ex nobis prodierunt, sed non erant ex nobis, nam si fuissent ex nobis, permansissent nobiscum; sed ut manifestaretur quoniam illi omnes non sunt ex nobis.
1JOHN|2|20|Sed vos unctionem habetis a Sancto et scitis omnes.
1JOHN|2|21|Non scripsi vobis quasi nescientibus veritatem sed quasi scientibus eam, et quoniam omne mendacium ex veritate non est.
1JOHN|2|22|Quis est mendax, nisi is qui negat quoniam Iesus est Christus? Hic est antichristus, qui negat Patrem et Filium.
1JOHN|2|23|Omnis, qui negat Filium, nec Patrem habet; qui confitetur Filium, et Patrem habet.
1JOHN|2|24|Vos, quod audistis ab initio, in vobis permaneat; si in vobis permanserit, quod ab initio audistis, et vos in Filio et in Patre manebitis.
1JOHN|2|25|Et haec est repromissio, quam ipse pollicitus est nobis: vitam aeternam.
1JOHN|2|26|Haec scripsi vobis de eis, qui seducunt vos.
1JOHN|2|27|Et vos, unctionem, quam accepistis ab eo, manet in vobis, et non necesse habetis, ut aliquis doceat vos; sed sicut unctio ipsius docet vos de omnibus, et verum est, et non est mendacium, et, sicut docuit vos, manetis in eo.
1JOHN|2|28|Et nunc, filioli, manete in eo, ut, cum apparuerit, habeamus fiduciam et non confundamur ab eo in adventu eius.
1JOHN|2|29|Si scitis quoniam iustus est, scitote quoniam et omnis, qui facit iustitiam, ex ipso natus est.
1JOHN|3|1|Videte qualem caritatem dedit nobis Pater, ut filii Dei nomine mur, et sumus! Propter hoc mundus non cognoscit nos, quia non cognovit eum.
1JOHN|3|2|Carissimi, nunc filii Dei sumus, et nondum manifestatum est quid erimus; scimus quoniam, cum ipse apparuerit, similes ei erimus, quoniam videbimus eum, sicuti est.
1JOHN|3|3|Et omnis, qui habet spem hanc in eo, purificat se, sicut ille purus est.
1JOHN|3|4|Omnis, qui facit peccatum, et iniquitatem facit, quia peccatum est iniquitas.
1JOHN|3|5|Et scitis quoniam ille apparuit, ut peccata tolleret, et peccatum in eo non est.
1JOHN|3|6|Omnis, qui in eo manet, non peccat; omnis, qui peccat, non vidit eum nec novit eum.
1JOHN|3|7|Filioli, nemo vos seducat. Qui facit iustitiam, iustus est, sicut ille iustus est;
1JOHN|3|8|qui facit peccatum, ex Diabolo est, quoniam a principio Diabolus peccat. Propter hoc apparuit Filius Dei, ut dissolvat opera Diaboli.
1JOHN|3|9|Omnis, qui natus est ex Deo, peccatum non facit, quoniam semen ipsius in eo manet; et non potest peccare, quoniam ex Deo natus est.
1JOHN|3|10|In hoc manifesti sunt filii Dei et filii Diaboli: omnis, qui non facit iustitiam, non est ex Deo, et qui non diligit fratrem suum.
1JOHN|3|11|Quoniam haec est annuntiatio, quam audistis ab initio, ut diligamus alterutrum.
1JOHN|3|12|Non sicut Cain: ex Maligno erat et occidit fratrem suum. Et propter quid occidit eum? Quoniam opera eius maligna erant, fratris autem eius iusta.
1JOHN|3|13|Nolite mirari, fratres, si odit vos mundus.
1JOHN|3|14|Nos scimus quoniam transivimus de morte in vitam, quoniam diligimus fratres; qui non diligit, manet in morte.
1JOHN|3|15|Omnis, qui odit fratrem suum, homicida est, et scitis quoniam omnis homicida non habet vitam aeternam in semetipso manentem.
1JOHN|3|16|In hoc novimus caritatem, quoniam ille pro nobis animam suam posuit; et nos debemus pro fratribus animas ponere.
1JOHN|3|17|Qui habuerit substantiam mundi et viderit fratrem suum necesse habere et clauserit viscera sua ab eo, quomodo caritas Dei manet in eo?
1JOHN|3|18|Filioli, non diligamus verbo nec lingua sed in opere et veritate.
1JOHN|3|19|In hoc cognoscemus quoniam ex veritate sumus, et in conspectu eius placabimus corda nostra,
1JOHN|3|20|quoniam si reprehenderit nos cor, maior est Deus corde nostro et cognoscit omnia.
1JOHN|3|21|Carissimi, si cor nostrum non reprehenderit nos, fiduciam habemus ad Deum
1JOHN|3|22|et, quodcumque petierimus, accipimus ab eo, quoniam mandata eius custodimus et ea, quae sunt placita coram eo, facimus.
1JOHN|3|23|Et hoc est mandatum eius, ut credamus nomini Filii eius Iesu Christi et diligamus alterutrum, sicut dedit mandatum nobis.
1JOHN|3|24|Et, qui servat mandata eius, in ipso manet, et ipse in eo; et in hoc cognoscimus quoniam manet in nobis, ex Spiritu, quem nobis dedit.
1JOHN|4|1|Carissimi, nolite omni spiritui credere, sed probate spiritus si ex Deo sint, quoniam multi pseudoprophetae prodierunt in mundum.
1JOHN|4|2|In hoc cognoscitis Spiritum Dei: omnis spiritus, qui confitetur Iesum Christum in carne venisse, ex Deo est.
1JOHN|4|3|Et omnis spiritus, qui non confitetur Iesum, ex Deo non est; et hoc est antichristi, quod audistis quoniam venit, et nunc iam in mundo est.
1JOHN|4|4|Vos ex Deo estis, filioli, et vicistis eos, quoniam maior est, qui in vobis est, quam qui in mundo.
1JOHN|4|5|Ipsi ex mundo sunt; ideo ex mundo loquuntur, et mundus eos audit.
1JOHN|4|6|Nos ex Deo sumus. Qui cognoscit Deum, audit nos; qui non est ex Deo, non audit nos. Ex hoc cognoscimus Spiritum veritatis et spiritum erroris.
1JOHN|4|7|Carissimi, diligamus invicem, quoniam caritas ex Deo est; et omnis, qui diligit, ex Deo natus est et cognoscit Deum.
1JOHN|4|8|Qui non diligit, non cognovit Deum, quoniam Deus caritas est.
1JOHN|4|9|In hoc apparuit caritas Dei in nobis, quoniam Filium suum unigenitum misit Deus in mundum, ut vivamus per eum.
1JOHN|4|10|In hoc est caritas, non quasi nos dilexerimus Deum, sed quoniam ipse dilexit nos et misit Filium suum propitiationem pro peccatis nostris.
1JOHN|4|11|Carissimi, si sic Deus dilexit nos, et nos debemus alterutrum diligere.
1JOHN|4|12|Deum nemo vidit umquam; si diligamus invicem, Deus in nobis manet, et caritas eius in nobis consummata est.
1JOHN|4|13|In hoc cognoscimus quoniam in ipso manemus, et ipse in nobis, quoniam de Spiritu suo dedit nobis.
1JOHN|4|14|Et nos vidimus et testificamur quoniam Pater misit Filium salvatorem mundi.
1JOHN|4|15|Quisque confessus fuerit: " Iesus est Filius Dei ", Deus in ipso manet, et ipse in Deo.
1JOHN|4|16|Et nos, qui credidimus, novimus caritatem, quam habet Deus in nobis. Deus caritas est; et, qui manet in caritate, in Deo manet, et Deus in eo manet.
1JOHN|4|17|In hoc consummata est caritas nobiscum, ut fiduciam habeamus in die iudicii; quia sicut ille est, et nos sumus in hoc mundo.
1JOHN|4|18|Timor non est in caritate, sed perfecta caritas foras mittit timorem, quoniam timor poenam habet; qui autem timet, non est consummatus in caritate.
1JOHN|4|19|Nos diligimus, quoniam ipse prior dilexit nos.
1JOHN|4|20|Si quis dixerit: " Diligo Deum ", et fratrem suum oderit, mendax est; qui enim non diligit fratrem suum, quem videt, Deum, quem non videt, non potest diligere.
1JOHN|4|21|Et hoc mandatum habemus ab eo, ut, qui diligit Deum, diligat et fratrem suum.
1JOHN|5|1|Omnis, qui credit quoniam Iesus est Christus, ex Deo natus est; et omnis, qui diligit Deum, qui genuit, diligit et eum, qui natus est ex eo.
1JOHN|5|2|In hoc cognoscimus quoniam diligimus natos Dei, cum Deum diligamus et mandata eius faciamus.
1JOHN|5|3|Haec est enim caritas Dei, ut mandata eius servemus; et mandata eius gravia non sunt,
1JOHN|5|4|quoniam omne, quod natum est ex Deo, vincit mundum; et haec est victoria, quae vicit mundum: fides nostra.
1JOHN|5|5|Quis est qui vincit mundum, nisi qui credit quoniam Iesus est Filius Dei?
1JOHN|5|6|Hic est, qui venit per aquam et sanguinem, Iesus Christus; non in aqua solum sed in aqua et in sanguine. Et Spiritus est, qui testificatur, quoniam Spiritus est veritas.
1JOHN|5|7|Quia tres sunt, qui testificantur:
1JOHN|5|8|Spiritus et aqua et sanguis; et hi tres in unum sunt.
1JOHN|5|9|Si testimonium hominum accipimus, testimonium Dei maius est, quoniam hoc est testimonium Dei, quia testificatus est de Filio suo.
1JOHN|5|10|Qui credit in Filium Dei, habet testimonium in se. Qui non credit Deo, mendacem facit eum, quoniam non credidit in testimonium, quod testificatus est Deus de Filio suo.
1JOHN|5|11|Et hoc est testimonium, quoniam vitam aeternam dedit nobis Deus, et haec vita in Filio eius est.
1JOHN|5|12|Qui habet Filium, habet vitam; qui non habet Filium Dei, vitam non habet.
1JOHN|5|13|Haec scripsi vobis, ut sciatis quoniam vitam habetis aeternam, qui creditis in nomen Filii Dei.
1JOHN|5|14|Et haec est fiducia, quam habemus ad eum, quia si quid petierimus secundum voluntatem eius, audit nos.
1JOHN|5|15|Et si scimus quoniam audit nos, quidquid petierimus, scimus quoniam habemus petitiones, quas postulavimus ab eo.
1JOHN|5|16|Si quis videt fratrem suum peccare peccatum non ad mortem, petet, et dabit ei Deus vitam, peccantibus non ad mortem. Est peccatum ad mortem; non pro illo dico, ut roget.
1JOHN|5|17|Omnis iniustitia peccatum est, et est peccatum non ad mortem.
1JOHN|5|18|Scimus quoniam omnis, qui natus est ex Deo, non peccat, sed ille, qui genitus est ex Deo, conservat eum, et Malignus non tangit eum.
1JOHN|5|19|Scimus quoniam ex Deo sumus, et mundus totus in Maligno positus est.
1JOHN|5|20|Et scimus quoniam Filius Dei venit et dedit nobis sensum, ut cognoscamus eum, qui verus est; et sumus in eo, qui verus est, in Filio eius Iesu Christo. Hic est qui verus est, Deus et vita aeterna.
1JOHN|5|21|Filioli, custodite vos a simulacris!
2JOHN|1|1|Presbyter electae dominae et filiis eius, quos ego diligo in veritate, et non ego solus, sed et omnes, qui noverunt veritatem,
2JOHN|1|2|propter veritatem, quae permanet in nobis et nobiscum erit in sempiternum.
2JOHN|1|3|Erit nobiscum gratia, misericordia, pax a Deo Patre et a Iesu Christo, Filio Patris, in veritate et caritate.
2JOHN|1|4|Gavisus sum valde, quoniam inveni de filiis tuis ambulantes in veritate, sicut mandatum accepimus a Patre.
2JOHN|1|5|Et nunc rogo te, domina, non tamquam mandatum novum scribens tibi, sed quod habuimus ab initio, ut diligamus alterutrum.
2JOHN|1|6|Et haec est caritas, ut ambulemus secundum mandata eius; hoc mandatum est, quemadmodum audistis ab initio, ut in eo ambuletis.
2JOHN|1|7|Quoniam multi seductores prodierunt in mundum, qui non confitentur Iesum Christum venientem in carne; hic est seductor et antichristus.
2JOHN|1|8|Videte vosmetipsos, ne perdatis, quae operati estis, sed ut mercedem plenam accipiatis.
2JOHN|1|9|Omnis, qui ultra procedit et non manet in doctrina Christi, Deum non habet; qui permanet in doctri na, hic et Patrem et Filium habet.
2JOHN|1|10|Si quis venit ad vos et hanc doctrinam non affert, nolite accipere eum in domum nec " Ave " ei dixeritis;
2JOHN|1|11|qui enim dicit illi: " Ave ", communicat operibus illius malignis.
2JOHN|1|12|Plura habens vobis scribere, nolui per chartam et atramentum; spero enim me futurum apud vos, et os ad os loqui, ut gaudium nostrum plenum sit.
2JOHN|1|13|Salutant te filii sororis tuae electae.
3JOHN|1|1|Presbyter Gaio carissimo, quem ego diligo in veritate.
3JOHN|1|2|Carissime, in omnibus exopto prospere te agere et valere, sicut prospere agit anima tua.
3JOHN|1|3|Nam gavisus sum valde, venientibus fratribus et testimonium perhibentibus veritati tuae, quomodo tu in veritate ambules.
3JOHN|1|4|Maius horum non habeo gaudium, quam ut audiam filios meos in veritate ambulare.
3JOHN|1|5|Carissime, fideliter facis, quidquid operaris in fratres et hoc in peregrinos,
3JOHN|1|6|qui testimonium reddiderunt caritati tuae in conspectu ecclesiae. Bene facies subveniens illis in via digne Deo;
3JOHN|1|7|pro nomine enim profecti sunt, nihil accipientes a gentilibus.
3JOHN|1|8|Nos ergo debemus sublevare huiusmodi, ut cooperatores simus veritatis.
3JOHN|1|9|Scripsi aliquid ecclesiae; sed is qui amat primatum gerere in eis, Diotrephes, non recipit nos.
3JOHN|1|10|Propter hoc, si venero, commonebo eius opera, quae facit verbis malignis garriens in nos; et quasi non ei ista sufficiant, nec ipse suscipit fratres et eos, qui cu piunt, prohibet et de ecclesia eicit.
3JOHN|1|11|Carissime, noli imitari malum, sed quod bonum est. Qui benefacit, ex Deo est; qui malefacit, non vidit Deum.
3JOHN|1|12|Demetrio testimonium redditur ab omnibus et ab ipsa veritate; sed et nos testimonium perhibemus, et scis quoniam testimonium nostrum verum est.
3JOHN|1|13|Multa habui scribere tibi, sed nolo per atramentum et calamum scribere tibi;
3JOHN|1|14|spero autem protinus te videre, et os ad os loquemur.
3JOHN|1|15|Pax tibi. Salutant te amici. Saluta amicos nominatim.
JUDE|1|1|Iudas Iesu Christi servus, frater autem Iacobi, his qui sunt vocati, in Deo Patre dilecti et Christo Iesu conservati:
JUDE|1|2|misericordia vobis et pax et caritas adimpleatur.
JUDE|1|3|Carissimi, omnem sollicitudinem faciens scribendi vobis de communi nostra salute, necesse habui scribere vobis, deprecans certare pro semel tradita sanctis fide.
JUDE|1|4|Subintroierunt enim quidam homines, qui olim praescripti sunt in hoc iudicium, impii, Dei nostri gratiam transferentes in luxuriam, et solum Dominatorem et Dominum nostrum Iesum Christum negantes.
JUDE|1|5|Commonere autem vos volo, scientes vos omnia, quoniam Dominus semel populum de terra Aegypti salvans, secundo eos, qui non crediderunt, perdidit;
JUDE|1|6|angelos vero, qui non servaverunt suum principatum, sed dereliquerunt suum domicilium, in iudicium magni diei vinculis aeternis sub caligine reservavit.
JUDE|1|7|Sicut Sodoma et Gomorra et finitimae civitates, simili modo exfornicatae et abeuntes post carnem alteram, factae sunt exemplum, ignis aeterni poenam sustinentes.
JUDE|1|8|Similiter vero et hi somniantes carnem quidem maculant, dominationem autem spernunt, glorias autem blasphemant.
JUDE|1|9|Cum Michael archangelus cum Diabolo disputans altercaretur de Moysis corpore, non est ausus iudicium inferre blasphemiae, sed dixit: " Increpet te Dominus! ".
JUDE|1|10|Hi autem, quaecumque quidem ignorant, blasphemant; quaecumque autem naturaliter tamquam muta animalia norunt, in his corrumpuntur.
JUDE|1|11|Vae illis, quia via Cain abierunt et errore Balaam mercede effusi sunt et contradictione Core perierunt!
JUDE|1|12|Hi sunt in agapis vestris maculae, convivantes sine timore, semetipsos pascentes; nubes sine aqua, quae a ventis circumferuntur; arbores autumnales infructuosae bis mortuae, eradicatae;
JUDE|1|13|fluctus feri maris despumantes suas confusiones; sidera errantia, quibus procella tenebrarum in aeternum servata est.
JUDE|1|14|Prophetavit autem et his septimus ab Adam Henoch dicens: " Ecce venit Dominus in sanctis milibus suis
JUDE|1|15|facere iudicium contra omnes et arguere omnem animam de omnibus operibus impietatis eorum, quibus impie egerunt, et de omnibus duris, quae locuti sunt contra eum peccatores impii ".
JUDE|1|16|Hi sunt murmuratores, querelosi, secundum concupiscentias suas ambulantes, et os illorum loquitur superba, mirantes personas quaestus causa.
JUDE|1|17|Vos autem, carissimi, memores estote verborum, quae praedicta sunt ab apostolis Domini nostri Iesu Christi,
JUDE|1|18|quoniam dicebant vobis: " In novissimo tempore venient illusores, secundum suas concupiscentias ambulantes impietatum".
JUDE|1|19|Hi sunt qui segregant, animales, Spiritum non habentes.
JUDE|1|20|Vos autem, carissimi, superaedificantes vosmetipsos sanctissimae vestrae fidei, in Spiritu Sancto orantes,
JUDE|1|21|ipsos vos in dilectione Dei servate, exspectantes misericordiam Domini nostri Iesu Christi in vitam aeternam.
JUDE|1|22|Et his quidem miseremini disputantibus;
JUDE|1|23|illos vero salvate de igne rapientes; aliis autem miseremini in timore, odientes et eam, quae carnalis est, maculatam tunicam.
JUDE|1|24|Ei autem, qui potest vos conservare sine peccato et constituere ante conspectum gloriae suae immaculatos in exsultatione,
JUDE|1|25|soli Deo salvatori nostro per Iesum Christum Dominum nostrum gloria, magnificentia, imperium et potestas ante omne saeculum et nunc et in omnia saecula. Amen.
REV|1|1|Apocalypsis Iesu Christi, quam dedit illi Deus palam facere ser vis suis, quae oportet fieri cito, et significavit mittens per angelum suum servo suo Ioanni,
REV|1|2|qui testificatus est verbum Dei et testimonium Iesu Christi, quaecumque vidit.
REV|1|3|Beatus, qui legit et qui audiunt verba prophetiae et servant ea, quae in ea scripta sunt; tempus enim prope est.
REV|1|4|Ioannes septem ecclesiis, quae sunt in Asia: Gratia vobis et pax ab eo, qui est et qui erat et qui venturus est, et a septem spiritibus, qui in conspectu throni eius sunt,
REV|1|5|et ab Iesu Christo, qui est testis fidelis, primogenitus mortuorum et princeps regum terrae.Ei, qui diligit nos et solvit nos a peccatis nostris in sanguine suo
REV|1|6|et fecit nos regnum, sacerdotes Deo et Patri suo, ipsi gloria et imperium in saecula saeculorum. Amen.
REV|1|7|Ecce venit cum nubibus, et videbit eum omnis oculus et qui eum pupugerunt, et plangent se super eum omnes tribus terrae. Etiam, amen.
REV|1|8|Ego sum Alpha et Omega, dicit Dominus Deus, qui est et qui erat et qui venturus est, Omnipotens.
REV|1|9|Ego Ioannes, frater vester et particeps in tribulatione et regno et patientia in Iesu, fui in insula, quae appellatur Patmos, propter verbum Dei et testimonium Iesu.
REV|1|10|Fui in spiritu in dominica die et audivi post me vocem magnam tamquam tubae
REV|1|11|dicentis: " Quod vides, scribe in libro et mitte septem ecclesiis: Ephesum et Smyrnam et Pergamum et Thyatiram et Sardis et Philadelphiam et Laodiciam ".
REV|1|12|Et conversus sum, ut viderem vocem, quae loquebatur mecum; et conversus vidi septem candelabra aurea
REV|1|13|et in medio candelabrorum quasi Filium hominis, vestitum podere et praecinctum ad mamillas zonam auream;
REV|1|14|caput autem eius et capilli erant candidi tamquam lana alba, tamquam nix, et oculi eius velut flamma ignis,
REV|1|15|et pedes eius similes orichalco sicut in camino ardenti, et vox illius tamquam vox aquarum multarum,
REV|1|16|et habebat in dextera manu sua stellas septem, et de ore eius gladius anceps acutus exibat, et facies eius sicut sol lucet in virtute sua.
REV|1|17|Et cum vidissem eum, cecidi ad pedes eius tamquam mortuus; et posuit dexteram suam super me dicens: " Noli timere! Ego sum primus et novissimus,
REV|1|18|et vivens et fui mortuus et ecce sum vivens in saecula saeculorum et habeo claves mortis et inferni.
REV|1|19|Scribe ergo, quae vidisti et quae sunt et quae oportet fieri post haec.
REV|1|20|Mysterium septem stellarum, quas vidisti ad dexteram meam, et septem candelabra aurea: septem stellae, angeli sunt septem ecclesiarum; et candelabra septem, septem ecclesiae sunt.
REV|2|1|Angelo ecclesiae, quae est Ephesi, scribe:Haec dicit, qui tenet septem stellas in dextera sua, qui ambulat in medio septem candelabrorum aureorum:
REV|2|2|Scio opera tua et laborem et patientiam tuam, et quia non potes sustinere malos et tentasti eos, qui se dicunt apostolos et non sunt, et invenisti eos mendaces;
REV|2|3|et patientiam habes et sustinuisti propter nomen meum et non defecisti.
REV|2|4|Sed habeo adversus te quod caritatem tuam primam reliquisti.
REV|2|5|Memor esto itaque unde excideris, et age paenitentiam et prima opera fac; sin autem, venio tibi et movebo candelabrum tuum de loco suo, nisi paenitentiam egeris.
REV|2|6|Sed hoc habes, quia odisti facta Nicolaitarum, quae et ego odi.
REV|2|7|Qui habet aurem, audiat quid Spiritus dicat ecclesiis. Vincenti dabo ei edere de ligno vitae, quod est in paradiso Dei.
REV|2|8|Et angelo ecclesiae, quae est Smyrnae, scribe:Haec dicit Primus et Novissimus, qui fuit mortuus et vixit:
REV|2|9|Scio tribulationem tuam et paupertatem tuam - sed dives es - et blasphemiam ab his, qui se dicunt Iudaeos esse et non sunt, sed sunt synagoga Satanae.
REV|2|10|Nihil horum timeas, quae passurus es. Ecce missurus est Diabolus ex vobis in carcerem, ut tentemini, et habebitis tribulationem diebus decem. Esto fidelis usque ad mortem, et dabo tibi coronam vitae.
REV|2|11|Qui habet aurem, audiat quid Spiritus dicat ecclesiis. Qui vicerit, non laedetur a morte secunda.
REV|2|12|Et angelo ecclesiae, quae est Pergami, scribe:Haec dicit, qui habet romphaeam ancipitem acutam:
REV|2|13|Scio, ubi habitas, ubi thronus est Satanae, et tenes nomen meum et non negasti fidem meam et in diebus Antipas, testis meus fidelis, qui occisus est apud vos, ubi Satanas habitat.
REV|2|14|Sed habeo adversus te pauca, quia habes illic tenentes doctrinam Balaam, qui docebat Balac mittere scandalum coram filiis Israel, edere idolothyta et fornicari;
REV|2|15|ita habes et tu tenentes doctrinam Nicolaitarum similiter.
REV|2|16|Ergo paenitentiam age; si quo minus, venio tibi cito et pugnabo cum illis in gladio oris mei.
REV|2|17|Qui habet aurem, audiat quid Spiritus dicat ecclesiis. Vincenti dabo ei de manna abscondito et dabo illi calculum candidum, et in calculo nomen novum scriptum, quod nemo scit, nisi qui accipit.
REV|2|18|Et angelo ecclesiae, quae est Thyatirae, scribe: Haec dicit Filius Dei, qui habet oculos ut flammam ignis, et pedes eius similes orichalco:
REV|2|19|Novi opera tua et caritatem et fidem et ministerium et patientiam tuam et opera tua novissima plura prioribus.
REV|2|20|Sed habeo adversus te, quia permittis mulierem Iezabel, quae se dicit prophetissam, et docet et seducit servos meos fornicari et manducare idolothyta.
REV|2|21|Et dedi illi tempus, ut paenitentiam ageret, et non vult paeniteri a fornicatione sua.
REV|2|22|Ecce mitto eam in lectum et, qui moechantur cum ea, in tribulationem magnam, nisi paenitentiam egerint ab operibus eius.
REV|2|23|Et filios eius interficiam in morte, et scient omnes ecclesiae quia ego sum scrutans renes et corda, et dabo unicuique vestrum secundum opera vestra.
REV|2|24|Vobis autem dico ceteris, qui Thyatirae estis, quicumque non habent doctrinam hanc, qui non cognoverunt altitudines Satanae, quemadmodum dicunt, non mittam super vos aliud pondus;
REV|2|25|tamen id quod habetis, tenete, donec veniam.
REV|2|26|Et, qui vicerit et qui custodierit usque in finem opera mea, dabo illi potestatem super gentes,
REV|2|27|et reget illas in virga ferrea,tamquam vasa fictilia confringentur,
REV|2|28|sicut et ego accepi a Patre meo, et dabo illi stellam matutinam.
REV|2|29|Qui habet aurem, audiat quid Spiritus dicat ecclesiis.
REV|3|1|Et angelo ecclesiae, quae est Sardis, scribe:Haec dicit, qui habet septem spiritus Dei et septem stellas: Scio opera tua, quia nomen habes quod vivas, et mortuus es.
REV|3|2|Esto vigilans et confirma cetera, quae moritura erant, non enim invenio opera tua plena coram Deo meo;
REV|3|3|in mente ergo habe qualiter acceperis et audieris, et serva et paenitentiam age. Si ergo non vigilaveris, veniam tamquam fur, et nescies qua hora veniam ad te.
REV|3|4|Sed habes pauca nomina in Sardis, qui non inquinaverunt vestimenta sua et ambulabunt mecum in albis, quia digni sunt.
REV|3|5|Qui vicerit, sic vestietur vestimentis albis, et non delebo nomen eius de libro vitae et confitebor nomen eius coram Patre meo et coram angelis eius.
REV|3|6|Qui habet aurem, audiat quid Spiritus dicat ecclesiis.
REV|3|7|Et angelo ecclesiae, quae est Philadelphiae, scribe:Haec dicit Sanctus, Verus, qui habet clavem David, qui aperit, et nemo claudet; et claudit, et nemo aperit:
REV|3|8|Scio opera tua - ecce dedi coram te ostium apertum, quod nemo potest claudere - quia modicam habes virtutem, et servasti verbum meum et non negasti nomen meum.
REV|3|9|Ecce dabo de synagoga Satanae, qui dicunt se Iudaeos esse et non sunt, sed mentiuntur; ecce faciam illos, ut veniant et adorent ante pedes tuos et scient quia ego dilexi te.
REV|3|10|Quoniam servasti verbum patientiae meae, et ego te servabo ab hora tentationis, quae ventura est super orbem universum tentare habitantes in terra.
REV|3|11|Venio cito; tene quod habes, ut nemo accipiat coronam tuam.
REV|3|12|Qui vicerit, faciam illum columnam in templo Dei mei, et foras non egredietur amplius; et scribam super eum nomen Dei mei et nomen civitatis Dei mei, novae Ierusalem, quae descendit de caelo a Deo meo, et nomen meum novum.
REV|3|13|Qui habet aurem, audiat quid Spiritus dicat ecclesiis.
REV|3|14|Et angelo ecclesiae, quae est Laodiciae, scribe:Haec dicit Amen, testis fidelis et verus, principium creaturae Dei:
REV|3|15|Scio opera tua, quia neque frigidus es neque calidus. Utinam frigidus esses aut calidus!
REV|3|16|Sic quia tepidus es et nec calidus nec frigidus, incipiam te evomere ex ore meo.
REV|3|17|Quia dicis: "Dives sum et locupletatus et nullius egeo", et nescis quia tu es miser et miserabilis et pauper et caecus et nudus,
REV|3|18|suadeo tibi emere a me aurum igne probatum, ut locuples fias et vestimentis albis induaris, et non appareat confusio nuditatis tuae, et collyrium ad inunguendum oculos tuos, ut videas.
REV|3|19|Ego, quos amo, arguo et castigo. Aemulare ergo et paenitentiam age.
REV|3|20|Ecce sto ad ostium et pulso. Si quis audierit vocem meam et aperuerit ianuam, introibo ad illum et cenabo cum illo, et ipse mecum.
REV|3|21|Qui vicerit, dabo ei sedere mecum in throno meo, sicut et ego vici et sedi cum Patre meo in throno eius.
REV|3|22|Qui habet aurem, audiat quid Spiritus dicat ecclesiis ".
REV|4|1|Post haec vidi: et ecce ostium apertum in caelo, et vox prima, quam audivi, tamquam tubae loquentis mecum dicens: " Ascende huc, et ostendam tibi, quae oportet fieri post haec ".
REV|4|2|Statim fui in spiritu: et ecce thronus positus erat in caelo; et supra thronum sedens;
REV|4|3|et, qui sedebat, similis erat aspectu lapidi iaspidi et sardino; et iris erat in circuitu throni, aspectu similis smaragdo.
REV|4|4|Et in circuitu throni, viginti quattuor thronos, et super thronos viginti quattuor seniores sedentes, circumamictos vestimentis albis, et super capita eorum coronas aureas.
REV|4|5|Et de throno procedunt fulgura et voces et tonitrua; et septem lampades ignis ardentes ante thronum, quae sunt septem spiritus Dei;
REV|4|6|et in conspectu throni tamquam mare vitreum simile crystallo. Et in medio throni et in circuitu throni quattuor animalia, plena oculis ante et retro:
REV|4|7|et animal primum simile leoni, et secundum animal simile vitulo, et tertium animal habens faciem quasi hominis, et quartum animal simile aquilae volanti.
REV|4|8|Et quattuor animalia singula eorum habebant alas senas, in circuitu et intus plenae sunt oculis; et requiem non habent die et nocte dicentia: " Sanctus, sanctus, sanctus Dominus, Deus omnipotens, qui erat et qui est et qui venturus est! ".
REV|4|9|Et cum darent illa animalia gloriam et honorem et gratiarum actionem sedenti super thronum, viventi in saecula saeculorum,
REV|4|10|procidebant viginti quattuor seniores ante sedentem in throno et adorabant viventem in saecula saeculorum et mittebant coronas suas ante thronum dicentes:
REV|4|11|" Dignus es, Domine et Deus noster,accipere gloriam et honorem et virtutem,quia tu creasti omnia,et propter voluntatem tuam erant et creata sunt ".
REV|5|1|Et vidi in dextera sedentis super thronum librum scriptum intus et foris, signatum sigillis septem.
REV|5|2|Et vidi angelum fortem praedicantem voce magna: " Quis est dignus aperire librum et solvere signacula eius? ".
REV|5|3|Et nemo poterat in caelo neque in terra neque subtus terram aperire librum neque respicere illum.
REV|5|4|Et ego flebam multum, quoniam nemo dignus inventus est aperire librum nec respicere eum.
REV|5|5|Et unus de senioribus dicit mihi: " Ne fleveris; ecce vicit leo de tribu Iudae, radix David, aperire librum et septem signacula eius ".
REV|5|6|Et vidi in medio throni et quattuor animalium et in medio seniorum Agnum stantem tamquam occisum, habentem cornua septem et oculos septem, qui sunt septem spiritus Dei missi in omnem terram.
REV|5|7|Et venit et accepit de dextera sedentis in throno.
REV|5|8|Et cum accepisset librum, quattuor animalia et viginti quattuor seniores ceciderunt coram Agno, habentes singuli citharas et phialas aureas plenas incensorum, quae sunt orationes sanctorum.
REV|5|9|Et cantant novum canticum dicentes: Dignus es accipere librumet aperire signacula eius,quoniam occisus es et redemisti Deo in sanguine tuoex omni tribu et lingua et populo et natione;
REV|5|10|et fecisti eos Deo nostro regnum et sacerdotes,et regnabunt super terram ".
REV|5|11|Et vidi et audivi vocem angelorum multorum in circuitu throni et animalium et seniorum, et erat numerus eorum myriades myriadum et milia milium,
REV|5|12|dicentium voce magna: Dignus est Agnus, qui occisus est, accipere virtutem et divitias et sapientiamet fortitudinem et honorem et gloriam et benedictionem ".
REV|5|13|Et omnem creaturam, quae in caelo est et super terram et sub terra et super mare et quae in eis omnia, audivi dicentes: "Sedenti super thronum et Agno benedictio et honor et gloria et potestas in saecula saeculorum ".
REV|5|14|Et quattuor animalia dicebant: " Amen "; et seniores ceciderunt et adoraverunt.
REV|6|1|Et vidi, cum aperuisset Agnus unum de septem sigillis, et audi vi unum de quattuor animalibus dicens tamquam voce tonitrui: " Veni ".
REV|6|2|Et vidi: et ecce equus albus; et, qui sedebat super illum, habebat arcum, et data est ei corona, et exivit vincens et ut vinceret.
REV|6|3|Et cum aperuisset sigillum secundum, audivi secundum animal dicens: " Veni ".
REV|6|4|Et exivit alius equus rufus; et, qui sedebat super illum, datum est ei, ut sumeret pacem de terra, et ut invicem se interficiant; et datus est illi gladius magnus.
REV|6|5|Et cum aperuisset sigillum tertium, audivi tertium animal dicens: " Veni. Et vidi: et ecce equus niger; et, qui sedebat super eum, habebat stateram in manu sua.
REV|6|6|Et audivi tamquam vocem in medio quattuor animalium dicentem: " Bilibris tritici denario, et tres bilibres hordei denario; et oleum et vinum ne laeseris ".
REV|6|7|Et cum aperuisset sigillum quartum, audivi vocem quarti animalis dicentis: " Veni ".
REV|6|8|Et vidi: et ecce equus pallidus; et, qui sedebat desuper, nomen illi Mors, et Infernus sequebatur eum; et data est illis potestas super quartam partem terrae interficere gladio et fame et morte et a bestiis terrae.
REV|6|9|Et cum aperuisset quintum sigillum, vidi subtus altare animas interfectorum propter verbum Dei et propter testimonium, quod habebant.
REV|6|10|Et clamaverunt voce magna dicentes: " Usquequo, Domine, sanctus et verus, non iudicas et vindicas sanguinem nostrum de his, qui habitant in terra? ".
REV|6|11|Et datae sunt illis singulae stolae albae; et dictum est illis, ut requiescant tempus adhuc modicum, donec impleantur et conservi eorum et fratres eorum, qui interficiendi sunt sicut et illi.
REV|6|12|Et vidi, cum aperuisset sigillum sextum, et terraemotus factus est magnus, et sol factus est niger tamquam saccus cilicinus, et luna tota facta est sicut sanguis,
REV|6|13|et stellae caeli ceciderunt in terram, sicut ficus mittit grossos suos, cum vento magno movetur,
REV|6|14|et caelum recessit sicut liber involutus, et omnis mons et insula de locis suis motae sunt.
REV|6|15|Et reges terrae et magnates et tribuni et divites et fortes et omnis servus et liber absconderunt se in speluncis et in petris montium;
REV|6|16|et dicunt montibus et petris: " Cadite super nos et abscondite nos a facie sedentis super thronum et ab ira Agni,
REV|6|17|quoniam venit dies magnus irae ipsorum, et quis poterit stare? ".
REV|7|1|Post haec vidi quattuor angelos stantes super quattuor angulos terrae tenentes quattuor ventos terrae, ne flaret ventus super terram neque super mare neque in ullam arborem.
REV|7|2|Et vidi alterum angelum ascendentem ab ortu solis, habentem sigillum Dei vivi; et clamavit voce magna quattuor angelis, quibus datum est nocere terrae et mari,
REV|7|3|dicens: " Nolite nocere terrae neque mari neque arboribus, quoadusque signemus servos Dei nostri in frontibus eorum ".
REV|7|4|Et audivi numerum signatorum, centum quadraginta quattuor milia signati ex omni tribu filiorum Israel:
REV|7|5|ex tribu Iudae duodecim milia signati, ex tribu Ruben duodecim milia, ex tribu Gad duodecim milia,
REV|7|6|ex tribu Aser duodecim milia, ex tribu Nephthali duodecim milia, ex tribu Manasse duodecim milia,
REV|7|7|ex tribu Simeon duodecim milia, ex tribu Levi duodecim milia, ex tribu Issachar duodecim milia,
REV|7|8|ex tribu Zabulon duodecim milia, ex tribu Ioseph duodecim milia, ex tribu Beniamin duodecim milia signati.
REV|7|9|Post haec vidi: et ecce turba magna, quam dinumerare nemo poterat, ex omnibus gentibus et tribubus et populis et linguis stantes ante thronum et in conspectu Agni, amicti stolis albis, et palmae in manibus eorum;
REV|7|10|et clamant voce magna dicentes: " Salus Deo nostro, qui sedet super thronum, et Agno ".
REV|7|11|Et omnes angeli stabant in circuitu throni et seniorum et quattuor animalium, et ceciderunt in conspectu throni in facies suas et adoraverunt Deum
REV|7|12|dicentes: Amen! Benedictio et gloria et sapientia et gratiarum actio et honor et virtus et fortitudo Deo nostro in saecula saeculorum. Amen ".
REV|7|13|Et respondit unus de senioribus dicens mihi: " Hi, qui amicti sunt stolis albis, qui sunt et unde venerunt? ".
REV|7|14|Et dixi illi: " Domine mi, tu scis ". Et dixit mihi: " Hi sunt qui veniunt de tribulatione magna et laverunt stolas suas et dealbaverunt eas in sanguine Agni.
REV|7|15|Ideo sunt ante thronum Dei et serviunt ei die ac nocte in templo eius; et, qui sedet in throno, habitabit super illos.
REV|7|16|Non esurient amplius neque sitient amplius, neque cadet super illos sol neque ullus aestus,
REV|7|17|quoniam Agnus, qui in medio throni est, pascet illos et deducet eos ad vitae fontes aquarum, et absterget Deus omnem lacrimam ex oculis eorum ".
REV|8|1|Et cum aperuisset sigillum septimum, factum est silentium in caelo quasi media hora.
REV|8|2|Et vidi septem angelos, qui stant in conspectu Dei, et datae sunt illis septem tubae.
REV|8|3|Et alius angelus venit et stetit ante altare habens turibulum aureum, et data sunt illi incensa multa, ut daret orationibus sanctorum omnium super altare aureum, quod est ante thronum.
REV|8|4|Et ascendit fumus incensorum de orationibus sanctorum de manu angeli coram Deo.
REV|8|5|Et accepit angelus turibulum et implevit illud de igne altaris et misit in terram; et facta sunt tonitrua et voces et fulgura et terraemotus.
REV|8|6|Et septem angeli, qui habebant septem tubas, paraverunt se, ut tuba canerent.
REV|8|7|Et primus tuba cecinit. Et facta est grando et ignis mixta in sanguine, et missum est in terram: et tertia pars terrae combusta est, et tertia pars arborum combusta est, et omne fenum viride combustum est.
REV|8|8|Et secundus angelus tuba cecinit. Et tamquam mons magnus igne ardens missus est in mare: et facta est tertia pars maris sanguis,
REV|8|9|et mortua est tertia pars creaturarum, quae in mari sunt, quae habent animas, et tertia pars navium interiit.
REV|8|10|Et tertius angelus tuba cecinit. Et cecidit de caelo stella magna ardens tamquam facula et cecidit super tertiam partem fluminum et super fontes aquarum.
REV|8|11|Et nomen stellae dicitur Absinthius. Et facta est tertia pars aquarum in absinthium, et multi hominum mortui sunt de aquis, quia amarae factae sunt.
REV|8|12|Et quartus angelus tuba cecinit. Et percussa est tertia pars solis et tertia pars lunae et tertia pars stellarum, ut obscuraretur tertia pars eorum, et diei non luceret pars tertia, et nox similiter.
REV|8|13|Et vidi et audivi unam aquilam volantem per medium caelum dicentem voce magna: " Vae, vae, vae habitantibus in terra de ceteris vocibus tubae trium angelorum, qui tuba canituri sunt!".
REV|9|1|Et quintus angelus tuba cecinit. Et vidi stellam de caelo cecidis se in terram, et data est illi clavis putei abyssi.
REV|9|2|Et aperuit puteum abyssi, et ascendit fumus ex puteo sicut fumus fornacis magnae; et obscuratus est sol et aer de fumo putei.
REV|9|3|Et de fumo exierunt locustae in terram, et data est illis potestas, sicut habent potestatem scorpiones terrae.
REV|9|4|Et dictum est illis, ne laederent fenum terrae neque omne viride neque omnem arborem, nisi tantum homines, qui non habent signum Dei in frontibus.
REV|9|5|Et datum est illis, ne occiderent eos, sed ut cruciarentur mensibus quinque; et cruciatus eorum ut cruciatus scorpii, cum percutit hominem.
REV|9|6|Et in diebus illis quaerent homines mortem et non invenient eam; et desiderabunt mori, et fugit mors ab ipsis.
REV|9|7|Et similitudines locustarum similes equis paratis in proelium, et super capita earum tamquam coronae similes auro, et facies earum sicut facies hominum;
REV|9|8|et habebant capillos sicut capillos mulierum, et dentes earum sicut leonum erant,
REV|9|9|et habebant loricas sicut loricas ferreas, et vox alarum earum sicut vox curruum equorum multorum currentium in bellum.
REV|9|10|Et habent caudas similes scorpionibus et aculeos, et in caudis earum potestas earum nocere hominibus mensibus quinque.
REV|9|11|Habent super se regem angelum abyssi, cui nomen Hebraice Abaddon et Graece nomen habet Apollyon.
REV|9|12|Vae unum abiit. Ecce veniunt adhuc duo vae post haec.
REV|9|13|Et sextus angelus tuba cecinit. Et audivi vocem unam ex cornibus altaris aurei, quod est ante Deum,
REV|9|14|dicentem sexto angelo, qui habebat tubam: " Solve quattuor angelos, qui alligati sunt super flumen magnum Euphraten ".
REV|9|15|Et soluti sunt quattuor angeli, qui parati erant in horam et diem et mensem et annum, ut occiderent tertiam partem hominum.
REV|9|16|Et numerus equestris exercitus vicies milies dena milia; audivi numerum eorum.
REV|9|17|Et ita vidi equos in visione et, qui sedebant super eos, habentes loricas igneas et hyacinthinas et sulphureas; et capita equorum erant tamquam capita leonum, et de ore ipsorum procedit ignis et fumus et sulphur.
REV|9|18|Ab his tribus plagis occisa est tertia pars hominum, de igne et fumo et sulphure, quod procedebat ex ore ipsorum.
REV|9|19|Potestas enim equorum in ore eorum est et in caudis eorum; nam caudae illorum similes serpentibus habentes capita, et in his nocent.
REV|9|20|Et ceteri homines, qui non sunt occisi in his plagis neque paenitentiam egerunt de operibus manuum suarum, ut non adorarent daemonia et simulacra aurea et argentea et aerea et lapidea et lignea, quae neque videre possunt neque audire neque ambulare,
REV|9|21|et non egerunt paenitentiam ab homicidiis suis neque a veneficiis suis neque a fornicatione sua neque a furtis suis.
REV|10|1|Et vidi alium angelum for tem descendentem de caelo amictum nube, et iris super caput, et facies eius erat ut sol, et pedes eius tamquam columnae ignis;
REV|10|2|et habebat in manu sua libellum apertum. Et posuit pedem suum dexterum supra mare, sinistrum autem super terram,
REV|10|3|et clamavit voce magna, quemadmodum cum leo rugit. Et cum clamasset, locuta sunt septem tonitrua voces suas.
REV|10|4|Et cum locuta fuissent septem tonitrua, scripturus eram; et audivi vocem de caelo dicentem: " Signa, quae locuta sunt septem tonitrua, et noli ea scribere ".
REV|10|5|Et angelus, quem vidi stantem supra mare et supra terram, levavit manum suam dexteram ad caelum
REV|10|6|et iuravit per Viventem in saecula saeculorum, qui creavit caelum et ea, quae in illo sunt, et terram et ea, quae in ea sunt, et mare et ea, quae in eo sunt: " Tempus amplius non erit,
REV|10|7|sed in diebus vocis septimi angeli, cum coeperit tuba canere, et consummatum est mysterium Dei, sicut evangelizavit servis suis prophetis.
REV|10|8|Et vox, quam audivi de caelo, iterum loquentem mecum et dicentem: " Vade, accipe librum apertum de manu angeli stantis supra mare et supra terram ".
REV|10|9|Et abii ad angelum dicens ei, ut daret mihi libellum. Et dicit mihi: " Accipe et devora illum; et faciet amaricare ventrem tuum, sed in ore tuo erit dulcis tamquam mel ".
REV|10|10|Et accepi libellum de manu angeli et devoravi eum, et erat in ore meo tamquam mel dulcis; et cum devorassem eum, amaricatus est venter meus.
REV|10|11|Et dicunt mihi: " Oportet te iterum prophetare super populis et gentibus et linguis et regibus multis ".
REV|11|1|Et datus est mihi calamus similis virgae dicens: " Surge et metire templum Dei et altare et adorantes in eo.
REV|11|2|Atrium autem, quod est foris templum, eice foras et ne metiaris illud, quoniam datum est gentibus, et civitatem sanctam calcabunt mensibus quadraginta duobus.
REV|11|3|Et dabo duobus testibus meis, et prophetabunt diebus mille ducentis sexaginta amicti saccis ".
REV|11|4|Hi sunt duae olivae et duo candelabra in conspectu Domini terrae stantes.
REV|11|5|Et si quis eis vult nocere, ignis exit de ore illorum et devorat inimicos eorum; et si quis voluerit eos laedere, sic oportet eum occidi.
REV|11|6|Hi habent potestatem claudendi caelum, ne pluat pluvia diebus prophetiae ipsorum; et potestatem habent super aquas convertendi eas in sanguinem et percutere terram omni plaga, quotienscumque voluerint.
REV|11|7|Et cum finierint testimonium suum, bestia, quae ascendit de abysso, faciet adversus illos bellum et vincet eos et occidet illos.
REV|11|8|Et corpus eorum in platea civitatis magnae, quae vocatur spiritaliter Sodoma et Aegyptus, ubi et Dominus eorum crucifixus est;
REV|11|9|et vident de populis et tribubus et linguis et gentibus corpus eorum per tres dies et dimidium, et corpora eorum non sinunt poni in monumento.
REV|11|10|Et inhabitantes terram gaudent super illis et iucundantur et munera mittent invicem, quoniam hi duo prophetae cruciaverunt eos, qui inhabitant super terram.
REV|11|11|Et post dies tres et dimidium spiritus vitae a Deo intravit in eos, et steterunt super pedes suos; et timor magnus cecidit super eos, qui videbant eos.
REV|11|12|Et audierunt vocem magnam de caelo dicentem illis: " Ascendite huc "; et ascenderunt in caelum in nube, et viderunt illos inimici eorum.
REV|11|13|Et in illa hora factus est terraemotus magnus, et decima pars civitatis cecidit, et occisi sunt in terraemotu nomina hominum septem milia, et reliqui in timorem sunt missi et dederunt gloriam Deo caeli.
REV|11|14|Vae secundum abiit; ecce vae tertium venit cito.
REV|11|15|Et septimus angelus tuba cecinit, et factae sunt voces magnae in caelo dicentes: " Factum est regnum huius mundi Domini nostri et Christi eius, et regnabit in saecula saeculorum ".
REV|11|16|Et viginti quattuor seniores, qui in conspectu Dei sedent in thronis suis, ceciderunt super facies suas et adoraverunt Deum
REV|11|17|dicentes: Gratias agimus tibi,Domine, Deus omnipotens,qui es et qui eras,quia accepisti virtutem tuam magnam et regnasti.
REV|11|18|Et iratae sunt gentes,et advenit ira tua, et tempus mortuorum iudicariet reddere mercedem servis tuis prophetis et sanctiset timentibus nomen tuum, pusillis et magnis,et exterminare eos, qui exterminant terram ".
REV|11|19|Et apertum est templum Dei in caelo, et visa est arca testamenti eius in templo eius; et facta sunt fulgura et voces et terraemotus et grando magna.
REV|12|1|Et signum magnum appa ruit in caelo: mulier amicta sole, et luna sub pedibus eius, et super caput eius corona stellarum duodecim;
REV|12|2|et in utero habens, et clamat parturiens et cruciatur, ut pariat.
REV|12|3|Et visum est aliud signum in caelo: et ecce draco rufus magnus, habens capita septem et cornua decem, et super capita sua septem diademata;
REV|12|4|et cauda eius trahit tertiam partem stellarum caeli et misit eas in terram. Et draco stetit ante mulierem, quae erat paritura, ut, cum peperisset, filium eius devoraret.
REV|12|5|Et peperit filium, masculum, qui recturus est omnes gentes in virga ferrea; et raptus est filius eius ad Deum et ad thronum eius.
REV|12|6|Et mulier fugit in desertum, ubi habet locum paratum a Deo, ut ibi pascant illam diebus mille ducentis sexaginta.
REV|12|7|Et factum est proelium in caelo, Michael et angeli eius, ut proeliarentur cum dracone. Et draco pugnavit et angeli eius,
REV|12|8|et non valuit, neque locus inventus est eorum amplius in caelo.
REV|12|9|Et proiectus est draco ille magnus, serpens antiquus, qui vocatur Diabolus et Satanas, qui seducit universum orbem; proiectus est in terram, et angeli eius cum illo proiecti sunt.
REV|12|10|Et audivi vocem magnam in caelo dicentem: Nunc facta est salus et virtus et regnum Dei nostriet potestas Christi eius,quia proiectus est accusator fratrum nostrorum,qui accusabat illos ante conspectum Dei nostri die ac nocte.
REV|12|11|Et ipsi vicerunt illum propter sanguinem Agniet propter verbum testimonii sui;et non dilexerunt animam suamusque ad mortem.
REV|12|12|Propterea laetamini, caeliet qui habitatis in eis.Vae terrae et mari, quia descendit Diabolus ad vos habens iram magnam, sciens quod modicum tempus habet! ".
REV|12|13|Et postquam vidit draco quod proiectus est in terram, persecutus est mulierem, quae peperit masculum.
REV|12|14|Et datae sunt mulieri duae alae aquilae magnae, ut volaret in desertum in locum suum, ubi alitur per tempus et tempora et dimidium temporis a facie serpentis.
REV|12|15|Et misit serpens ex ore suo post mulierem aquam tamquam flumen, ut eam faceret trahi a flumine.
REV|12|16|Et adiuvit terra mulierem, et aperuit terra os suum et absorbuit flumen, quod misit draco de ore suo.
REV|12|17|Et iratus est draco in mulierem et abiit facere proelium cum reliquis de semine eius, qui custodiunt mandata Dei et habent testimonium Iesu.
REV|12|18|Et stetit super arenam maris.
REV|13|1|Et vidi de mari bestiam ascendentem, habentem cor nua decem et capita septem, et super cornua eius decem diademata, et super capita eius nomina blasphemiae.
REV|13|2|Et bestia, quam vidi, similis erat pardo, et pedes eius sicut ursi, et os eius sicut os leonis. Et dedit illi draco virtutem suam et thronum suum et potestatem magnam.
REV|13|3|Et unum de capitibus suis quasi occisum in mortem, et plaga mortis eius curata est.Et admirata est universa terra post bestiam,
REV|13|4|et adoraverunt draconem, quia dedit potestatem bestiae, et adoraverunt bestiam dicentes: " Quis similis bestiae, et quis potest pugnare cum ea?.
REV|13|5|Et datum est ei os loquens magna et blasphemias, et data est illi potestas facere menses quadraginta duos.
REV|13|6|Et aperuit os suum in blasphemias ad Deum, blasphemare nomen eius et tabernaculum eius, eos, qui in caelo habitant.
REV|13|7|Et datum est illi bellum facere cum sanctis et vincere illos, et data est ei potestas super omnem tribum et populum et linguam et gentem.
REV|13|8|Et adorabunt eum omnes, qui inhabitant terram, cuiuscumque non est scriptum nomen in libro vitae Agni, qui occisus est, ab origine mundi.
REV|13|9|Si quis habet aurem, audiat:
REV|13|10|Si quis in captivitatem,in captivitatem vadit;si quis in gladio debet occidi,oportet eum in gladio occidi.Hic est patientia et fides sanctorum.
REV|13|11|Et vidi aliam bestiam ascendentem de terra, et habebat cornua duo similia agni, et loquebatur sicut draco.
REV|13|12|Et potestatem prioris bestiae omnem facit in conspectu eius. Et facit terram et inhabitantes in ea adorare bestiam primam, cuius curata est plaga mortis.
REV|13|13|Et facit signa magna, ut etiam ignem faciat de caelo descendere in terram in conspectu hominum.
REV|13|14|Et seducit habitantes terram propter signa, quae data sunt illi facere in conspectu bestiae, dicens habitantibus in terra, ut faciant imaginem bestiae, quae habet plagam gladii et vixit.
REV|13|15|Et datum est illi, ut daret spiritum imagini bestiae, ut et loquatur imago bestiae; et faciat, ut quicumque non adoraverint imaginem bestiae, occidantur.
REV|13|16|Et facit omnes pusillos et magnos et divites et pauperes et liberos et servos accipere characterem in dextera manu sua aut in frontibus suis,
REV|13|17|et ne quis possit emere aut vendere, nisi qui habet characterem, nomen bestiae aut numerum nominis eius.
REV|13|18|Hic sapientia est: qui habet intellectum, computet numerum bestiae; numerus enim hominis est: et numerus eius est sescenti sexaginta sex.
REV|14|1|Et vidi: et ecce Agnus stans supra montem Sion, et cum illo centum quadraginta quattuor milia, habentes nomen eius et nomen Patris eius scriptum in frontibus suis.
REV|14|2|Et audivi vocem de caelo tamquam vocem aquarum multarum et tamquam vocem tonitrui magni; et vox, quam audivi, sicut citharoedorum citharizantium in citharis suis.
REV|14|3|Et cantant quasi canticum novum ante thronum et ante quattuor animalia et seniores. Et nemo poterat discere canticum, nisi illa centum quadraginta quattuor milia, qui empti sunt de terra.
REV|14|4|Hi sunt qui cum mulieribus non sunt coinquinati, virgines enim sunt. Hi qui sequuntur Agnum, quocumque abierit. Hi empti sunt ex hominibus primitiae Deo et Agno;
REV|14|5|et in ore ipsorum non est inventum mendacium: sine macula sunt.
REV|14|6|Et vidi alterum angelum volantem per medium caelum, habentem evangelium aeternum, ut evangelizaret super sedentes in terra et super omnem gentem et tribum et linguam et populum;
REV|14|7|dicens magna voce: " Timete Deum et date illi gloriam, quia venit hora iudicii eius; et adorate eum, qui fecit caelum et terram et mare et fontes aquarum ".
REV|14|8|Et alius angelus secutus est dicens: " Cecidit, cecidit Babylon illa magna, quae a vino irae fornicationis suae potionavit omnes gentes! ".
REV|14|9|Et alius angelus tertius secutus est illos dicens voce magna: " Si quis adoraverit bestiam et imaginem eius et acceperit characterem in fronte sua aut in manu sua,
REV|14|10|et hic bibet de vino irae Dei, quod mixtum est mero in calice irae ipsius, et cruciabitur igne et sulphure in conspectu angelorum sanctorum et ante conspectum Agni.
REV|14|11|Et fumus tormentorum eorum in saecula saeculorum ascendit, nec habent requiem die ac nocte, qui adoraverunt bestiam et imaginem eius, et si quis acceperit characterem nominis eius ".
REV|14|12|Hic patientia sanctorum est, qui custodiunt mandata Dei et fidem Iesu.
REV|14|13|Et audivi vocem de caelo dicentem: " Scribe: Beati mortui, qui in Domino moriuntur amodo. Etiam, dicit Spiritus, ut requiescant a laboribus suis; opera enim illorum sequuntur illos ".
REV|14|14|Et vidi: et ecce nubem candidam, et supra nubem sedentem quasi Filium hominis, habentem super caput suum coronam auream et in manu sua falcem acutam.
REV|14|15|Et alter angelus exivit de templo clamans voce magna ad sedentem super nubem: " Mitte falcem tuam et mete, quia venit hora, ut metatur, quoniam aruit messis terrae ".
REV|14|16|Et misit, qui sedebat supra nubem, falcem suam in terram, et messa est terra.
REV|14|17|Et alius angelus exivit de templo, quod est in caelo, habens et ipse falcem acutam.
REV|14|18|Et alius angelus de altari, habens potestatem supra ignem, et clamavit voce magna ad eum, qui habebat falcem acutam, dicens: " Mitte falcem tuam acutam et vindemia botros vineae terrae, quoniam maturae sunt uvae eius ".
REV|14|19|Et misit angelus falcem suam in terram et vindemiavit vineam terrae et misit in lacum irae Dei magnum.
REV|14|20|Et calcatus est lacus extra civitatem, et exivit sanguis de lacu usque ad frenos equorum per stadia mille sescenta.
REV|15|1|Et vidi aliud signum in caelo magnum et mirabile: angelos septem habentes plagas septem novissimas, quoniam in illis consummata est ira Dei.
REV|15|2|Et vidi tamquam mare vitreum mixtum igne; et eos, qui vicerunt bestiam et imaginem illius et numerum nominis eius, stantes supra mare vitreum, habentes citharas Dei.
REV|15|3|Et cantant canticum Moysis servi Dei et canticum Agni dicentes: Magna et mirabilia opera tua,Domine, Deus omnipotens;iustae et verae viae tuae,Rex gentium!
REV|15|4|Quis non timebit, Domine,et glorificabit nomen tuum?Quia solus Sanctus,quoniam omnes gentes venientet adorabunt in conspectu tuo,quoniam iudicia tua manifestata sunt ".
REV|15|5|Et post haec vidi: et apertum est templum tabernaculi testimonii in caelo,
REV|15|6|et exierunt septem angeli habentes septem plagas de templo, vestiti lino mundo candido et praecincti circa pectora zonis aureis.
REV|15|7|Et unum ex quattuor animalibus dedit septem angelis septem phialas aureas plenas iracundiae Dei viventis in saecula saeculorum.
REV|15|8|Et impletum est templum fumo de gloria Dei et de virtute eius; et nemo poterat introire in templum, donec consummarentur septem plagae septem angelorum.
REV|16|1|Et audivi vocem magnam de templo dicentem septem an gelis: " Ite et effundite septem phialas irae Dei in terram ".
REV|16|2|Et abiit primus et effudit phialam suam in terram; et factum est vulnus saevum ac pessimum in homines, qui habebant characterem bestiae, et eos, qui adorabant imaginem eius.
REV|16|3|Et secundus effudit phialam suam in mare; et factus est sanguis tamquam mortui, et omnis anima vivens mortua est, quae est in mari.
REV|16|4|Et tertius effudit phialam suam in flumina et in fontes aquarum; et factus est sanguis.
REV|16|5|Et audivi angelum aquarum dicentem: " Iustus es, qui es et qui eras, Sanctus, quia haec iudicasti;
REV|16|6|quia sanguinem sanctorum et prophetarum fuderunt, et sanguinem eis dedisti bibere: digni sunt! ".
REV|16|7|Et audivi altare dicens: " Etiam, Domine, Deus omnipotens, vera et iusta iudicia tua! ".
REV|16|8|Et quartus effudit phialam suam in solem; et datum est illi aestu afficere homines in igne.
REV|16|9|Et aestuaverunt homines aestu magno; et blasphemaverunt nomen Dei habentis potestatem super has plagas et non egerunt paenitentiam, ut darent illi gloriam.
REV|16|10|Et quintus effudit phialam suam super thronum bestiae; et factum est regnum eius tenebrosum, et commanducaverunt linguas suas prae dolore
REV|16|11|et blasphemaverunt Deum caeli prae doloribus suis et vulneribus suis et non egerunt paenitentiam ex operibus suis.
REV|16|12|Et sextus effudit phialam suam super flumen illud magnum Euphraten; et exsiccata est aqua eius, ut praepararetur via regibus, qui sunt ab ortu solis.
REV|16|13|Et vidi de ore draconis et de ore bestiae et de ore pseudoprophetae spiritus tres immundos velut ranas;
REV|16|14|sunt enim spiritus daemoniorum facientes signa, qui procedunt ad reges universi orbis congregare illos in proelium diei magni Dei omnipotentis.
REV|16|15|Ecce venio sicut fur. Beatus, qui vigilat et custodit vestimenta sua, ne nudus ambulet, et videant turpitudinem eius.
REV|16|16|Et congregavit illos in locum, qui vocatur Hebraice Harmagedon.
REV|16|17|Et septimus effudit phialam suam in aerem; et exivit vox magna de templo a throno dicens: " Factum est! ".
REV|16|18|Et facta sunt fulgura et voces et tonitrua, et terraemotus factus est magnus, qualis numquam fuit, ex quo homo fuit super terram, talis terraemotus sic magnus.
REV|16|19|Et facta est civitas magna in tres partes, et civitates gentium ceciderunt. Et Babylon magna venit in memoriam ante Deum dare ei calicem vini indignationis irae eius.
REV|16|20|Et omnis insula fugit, et montes non sunt inventi.
REV|16|21|Et grando magna sicut talentum descendit de caelo in homines; et blasphemaverunt homines Deum propter plagam grandinis, quoniam magna est plaga eius nimis.
REV|17|1|Et venit unus de septem angelis, qui habebant septem phialas, et locutus est mecum dicens: " Veni, ostendam tibi damnationem meretricis magnae, quae sedet super aquas multas,
REV|17|2|cum qua fornicati sunt reges terrae, et inebriati sunt, qui inhabitant terram, de vino prostitutionis eius ".
REV|17|3|Et abstulit me in desertum in spiritu. Et vidi mulierem sedentem super bestiam coccineam, plenam nominibus blasphemiae, habentem capita septem et cornua decem.
REV|17|4|Et mulier erat circumdata purpura et coccino, et inaurata auro et lapide pretioso et margaritis, habens poculum aureum in manu sua plenum abominationibus et immunditiis fornicationis eius;
REV|17|5|et in fronte eius nomen scriptum, mysterium: " Babylon magna, mater fornicationum et abominationum terrae ".
REV|17|6|Et vidi mulierem ebriam de sanguine sanctorum et de sanguine martyrum Iesu. Et miratus sum, cum vidissem illam, admiratione magna.
REV|17|7|Et dixit mihi angelus. " Quare miraris? Ego tibi dicam mysterium mulieris et bestiae, quae portat eam, quae habet capita septem et decem cornua:
REV|17|8|bestia, quam vidisti, fuit et non est, et ascensura est de abysso et in interitum ibit. Et mirabuntur inhabitantes terram, quorum non sunt scripta nomina in libro vitae a constitutione mundi, videntes bestiam, quia erat et non est et aderit.
REV|17|9|Hic est sensus, qui habet sapientiam. Septem capita, septem montes sunt, super quos mulier sedet. Et reges septem sunt:
REV|17|10|quinque ceciderunt, unus est, alius nondum venit; et, cum venerit, oportet illum breve tempus manere.
REV|17|11|Et bestia, quae erat et non est, et is octavus est et de septem est et in interitum vadit.
REV|17|12|Et decem cornua, quae vidisti, decem reges sunt, qui regnum nondum acceperunt, sed potestatem tamquam reges una hora accipiunt cum bestia.
REV|17|13|Hi unum consilium habent et virtutem et potestatem suam bestiae tradunt.
REV|17|14|Hi cum Agno pugnabunt; et Agnus vincet illos, quoniam Dominus dominorum est et Rex regum, et qui cum illo sunt vocati et electi et fideles ".
REV|17|15|Et dicit mihi: " Aquae, quas vidisti, ubi meretrix sedet, populi et turbae sunt et gentes et linguae.
REV|17|16|Et decem cornua, quae vidisti, et bestia, hi odient fornicariam et desolatam facient illam et nudam, et carnes eius manducabunt et ipsam igne concremabunt;
REV|17|17|Deus enim dedit in corda eorum, ut faciant, quod illi placitum est, et faciant unum consilium et dent regnum suum bestiae, donec consummentur verba Dei.
REV|17|18|Et mulier, quam vidisti, est civitas magna, quae habet regnum super reges terrae ".
REV|18|1|Post haec vidi alium ange lum descendentem de caelo, habentem potestatem magnam; et terra illuminata est a claritate eius.
REV|18|2|Et clamavit in forti voce dicens: " Cecidit, cecidit Babylon magna et facta est habitatio daemoniorum et custodia omnis spiritus immundi et custodia omnis bestiae immundae et odibilis;
REV|18|3|quia de vino irae fornicationis eius biberunt omnes gentes, et reges terrae cum illa fornicati sunt, et mercatores terrae de virtute deliciarum eius divites facti sunt! ".
REV|18|4|Et audivi aliam vocem de caelo dicentem: " Exite de illa, populus meus, ut ne comparticipes sitis peccatorum eius et de plagis eius non accipiatis,
REV|18|5|quoniam pervenerunt peccata eius usque ad caelum, et recordatus est Deus iniquitatum eius.
REV|18|6|Reddite illi, sicut et ipsa reddidit, et duplicate duplicia secundum opera eius; in poculo, quo miscuit, miscete illi duplum.
REV|18|7|Quantum glorificavit se et in deliciis fuit, tantum date illi tormentum et luctum. Quia in corde suo dicit: "Sedeo regina et vidua non sum et luctum non videbo",
REV|18|8|ideo in una die venient plagae eius, mors et luctus et fames, et igne comburetur, quia fortis est Dominus Deus, qui iudicavit illam ".
REV|18|9|Et flebunt et plangent se super illam reges terrae, qui cum illa fornicati sunt et in deliciis vixerunt, cum viderint fumum incendii eius,
REV|18|10|longe stantes propter timorem tormentorum eius, dicentes: " Vae, vae, civitas illa magna, Babylon, civitas illa fortis, quoniam una hora venit iudicium tuum! ".
REV|18|11|Et negotiatores terrae flent et lugent super illam, quoniam mercem eorum nemo emit amplius:
REV|18|12|mercem auri et argenti et lapidis pretiosi et margaritarum, et byssi et purpurae et serici et cocci, et omne lignum thyinum et omnia vasa eboris et omnia vasa de ligno pretiosissimo et aeramento et ferro et marmore,
REV|18|13|et cinnamomum et amomum et odoramenta et unguenta et tus, et vinum et oleum et similam et triticum, et iumenta et oves et equorum et raedarum, et mancipiorum et animas hominum.
REV|18|14|Et fructus tui, desiderium animae, discesserunt a te, et omnia pinguia et clara perierunt a te, et amplius illa iam non invenient.
REV|18|15|Mercatores horum, qui divites facti sunt ab ea, longe stabunt propter timorem tormentorum eius flentes ac lugentes,
REV|18|16|dicentes: " Vae, vae, civitas illa magna, quae amicta erat byssino et purpura et cocco, et deaurata auro et lapide pretioso et margarita,
REV|18|17|quoniam una hora desolatae sunt tantae divitiae! ".Et omnis gubernator et omnis, qui in locum navigat, et nautae et, quotquot maria operantur, longe steterunt
REV|18|18|et clamabant, videntes fumum incendii eius, dicentes: " Quae similis civitati huic magnae? ".
REV|18|19|Et miserunt pulverem super capita sua et clamabant, flentes et lugentes, dicentes: " Vae, vae, civitas illa magna, in qua divites facti sunt omnes, qui habent naves in mari, de opibus eius, quoniam una hora desolata est!
REV|18|20|Exsulta super eam, caelum, et sancti et apostoli et prophetae, quoniam iudicavit Deus iudicium vestrum de illa! ".
REV|18|21|Et sustulit unus angelus fortis lapidem quasi molarem magnum et misit in mare dicens: "Impetu sic mittetur Babylon magna illa civitas et ultra iam non invenietur.
REV|18|22|Et vox citharoedorum et musicorum et tibia canentium et tuba non audietur in te amplius, et omnis artifex omnis artis non invenietur in te amplius, et vox molae non audietur in te amplius,
REV|18|23|et lux lucernae non lucebit tibi amplius, et vox sponsi et sponsae non audietur in te amplius; quia mercatores tui erant magnates terrae, quia in veneficiis tuis erraverunt omnes gentes,
REV|18|24|et in ea sanguis prophetarum et sanctorum inventus est et omnium, qui interfecti sunt in terra! ".
REV|19|1|Post haec audivi quasi vo cem magnam turbae multae in caelo dicentium: Alleluia!Salus et gloria et virtus Deo nostro,
REV|19|2|quia vera et iusta iudicia eius;quia iudicavit de meretrice magna, quae corrupit terram in prostitutione sua, et vindicavit sanguinem servorum suorum de manibus eius! ".
REV|19|3|Et iterum dixerunt: " Alleluia! Et fumus eius ascendit in saecula saeculorum! ".
REV|19|4|Et ceciderunt seniores viginti quattuor et quattuor animalia et adoraverunt Deum sedentem super thronum dicentes: " Amen. Alleluia ".
REV|19|5|Et vox de throno exivit dicens: Laudem dicite Deo nostro, omnes servi eiuset qui timetis eum, pusilli et magni! ".
REV|19|6|Et audivi quasi vocem turbae magnae et sicut vocem aquarum multarum et sicut vocem tonitruum magnorum dicentium: Alleluia,quoniam regnavit Dominus, Deus noster omnipotens.
REV|19|7|Gaudeamus et exsultemus et demus gloriam ei,quia venerunt nuptiae Agni,et uxor eius praeparavit se.
REV|19|8|Et datum est illi, ut cooperiat se byssino splendenti mundo: byssinum enim iustificationes sunt sanctorum ".
REV|19|9|Et dicit mihi: " Scribe: Beati, qui ad cenam nuptiarum Agni vocati sunt!. Et dicit mihi: " Haec verba Dei vera sunt ".
REV|19|10|Et cecidi ante pedes eius, ut adorarem eum. Et dicit mihi: " Vide, ne feceris! Conservus tuus sum et fratrum tuorum habentium testimonium Iesu. Deum adora. Testimonium enim Iesu est spiritus prophetiae ".
REV|19|11|Et vidi caelum apertum: et ecce equus albus; et, qui sedebat super eum, vocabatur Fidelis et Verax, et in iustitia iudicat et pugnat.
REV|19|12|Oculi autem eius sicut flamma ignis, et in capite eius diademata multa, habens nomen scriptum, quod nemo novit nisi ipse;
REV|19|13|et vestitus veste aspersa sanguine, et vocatur nomen eius Verbum Dei.
REV|19|14|Et exercitus, qui sunt in caelo, sequebantur eum in equis albis, vestiti byssino albo mundo.
REV|19|15|Et de ore ipsius procedit gladius acutus, ut in ipso percutiat gentes, et ipse reget eos in virga ferrea; et ipse calcat torcular vini furoris irae Dei omnipotentis.
REV|19|16|Et habet super vestimentum et super femur suum nomen scriptum: Rex regum et Dominus dominorum.
REV|19|17|Et vidi unum angelum stantem in sole, et clamavit voce magna dicens omnibus avibus, quae volabant per medium caeli: "Venite, congregamini ad cenam magnam Dei,
REV|19|18|ut manducetis carnes regum et carnes tribunorum et carnes fortium et carnes equorum et sedentium in ipsis et carnes omnium liberorum ac servorum et pusillorum ac magnorum ".
REV|19|19|Et vidi bestiam et reges terrae et exercitus eorum congregatos ad faciendum proelium cum illo, qui sedebat super equum, et cum exercitu eius.
REV|19|20|Et apprehensa est bestia et cum illa pseudopropheta, qui fecit signa coram ipsa, quibus seduxit eos, qui acceperunt characterem bestiae et qui adorant imaginem eius; vivi missi sunt hi duo in stagnum ignis ardentis sulphure.
REV|19|21|Et ceteri occisi sunt in gladio sedentis super equum, qui procedit de ore ipsius, et omnes aves saturatae sunt carnibus eorum.
REV|20|1|Et vidi angelum descen dentem de caelo habentem clavem abyssi et catenam magnam in manu sua.
REV|20|2|Et apprehendit draconem, serpentem antiquum, qui est Diabolus et Satanas, et ligavit eum per annos mille;
REV|20|3|et misit eum in abyssum et clausit et signavit super illum, ut non seducat amplius gentes, donec consummentur mille anni; post haec oportet illum solvi modico tempore.
REV|20|4|Et vidi thronos, et sederunt super eos, et iudicium datum est illis; et animas decollatorum propter testimonium Iesu et propter verbum Dei, et qui non adoraverunt bestiam neque imaginem eius nec acceperunt characterem in frontibus et in manibus suis; et vixerunt et regnaverunt cum Christo mille annis.
REV|20|5|Ceteri mortuorum non vixerunt, donec consummentur mille anni. Haec est resurrectio prima.
REV|20|6|Beatus et sanctus, qui habet partem in resurrectione prima! In his secunda mors non habet potestatem, sed erunt sacerdotes Dei et Christi et regnabunt cum illo mille annis.
REV|20|7|Et cum consummati fuerint mille anni, solvetur Satanas de carcere suo
REV|20|8|et exibit seducere gentes, quae sunt in quattuor angulis terrae, Gog et Magog; congregare eos in proelium, quorum numerus est sicut arena maris.
REV|20|9|Et ascenderunt super latitudinem terrae et circumierunt castra sanctorum et civitatem dilectam. Et descendit ignis de caelo et devoravit eos;
REV|20|10|et Diabolus, qui seducebat eos, missus est in stagnum ignis et sulphuris, ubi et bestia et pseudopropheta, et cruciabuntur die ac nocte in saecula saeculorum.
REV|20|11|Et vidi thronum magnum candidum et sedentem super eum, a cuius aspectu fugit terra et caelum, et locus non est inventus eis.
REV|20|12|Et vidi mortuos, magnos et pusillos, stantes in conspectu throni; et libri aperti sunt. Et alius liber apertus est, qui est vitae; et iudicati sunt mortui ex his, quae scripta erant in libris, secundum opera ipsorum.
REV|20|13|Et dedit mare mortuos, qui in eo erant, et mors et infernus dederunt mortuos, qui in ipsis erant; et iudicati sunt singuli secundum opera ipsorum.
REV|20|14|Et mors et infernus missi sunt in stagnum ignis. Haec mors secunda est, stagnum ignis.
REV|20|15|Et si quis non est inventus in libro vitae scriptus, missus est in stagnum ignis.
REV|21|1|Et vidi caelum novum et ter ram novam; primum enim caelum et prima terra abierunt, et mare iam non est.
REV|21|2|Et civitatem sanctam Ierusalem novam vidi descendentem de caelo a Deo, paratam sicut sponsam ornatam viro suo.
REV|21|3|Et audivi vocem magnam de throno dicentem: "Ecce tabernaculum Dei cum hominibus! Et habitabit cum eis, et ipsi populi eius erunt, et ipse Deus cum eis erit eorum Deus;
REV|21|4|et absterget omnem lacrimam ab oculis eorum, et mors ultra non erit, neque luctus neque clamor neque dolor erit ultra, quia prima abierunt ".
REV|21|5|Et dixit, qui sedebat super throno: " Ecce nova facio omnia ". Et dicit: Scribe: Haec verba fidelia sunt et vera ".
REV|21|6|Et dixit mihi: " Facta sunt! Ego sum Alpha et Omega, principium et finis. Ego sitienti dabo de fonte aquae vivae gratis.
REV|21|7|Qui vicerit, hereditabit haec, et ero illi Deus, et ille erit mihi filius.
REV|21|8|Timidis autem et incredulis et exsecratis et homicidis et fornicatoribus et veneficis et idololatris et omnibus mendacibus, pars illorum erit in stagno ardenti igne et sulphure, quod est mors secunda ".
REV|21|9|Et venit unus de septem angelis habentibus septem phialas plenas septem plagis novissimis et locutus est mecum dicens: " Veni, ostendam tibi sponsam uxorem Agni ".
REV|21|10|Et sustulit me in spiritu super montem magnum et altum et ostendit mihi civitatem sanctam Ierusalem descendentem de caelo a Deo,
REV|21|11|habentem claritatem Dei; lumen eius simile lapidi pretiosissimo, tamquam lapidi iaspidi, in modum crystalli;
REV|21|12|et habebat murum magnum et altum et habebat portas duodecim et super portas angelos duodecim et nomina inscripta, quae sunt duodecim tribuum filiorum Israel.
REV|21|13|Ab oriente portae tres, et ab aquilone portae tres, et ab austro portae tres, et ab occasu portae tres;
REV|21|14|et murus civitatis habens fundamenta duodecim, et super ipsis duodecim nomina duodecim apostolorum Agni.
REV|21|15|Et, qui loquebatur mecum, habebat mensuram arundinem auream, ut metiretur civitatem et portas eius et murum eius.
REV|21|16|Et civitas in quadro posita est, et longitudo eius tanta est quanta et latitudo. Et mensus est civitatem arundine per stadia duodecim milia; longitudo et latitudo et altitudo eius aequales sunt.
REV|21|17|Et mensus est murum eius centum quadraginta quattuor cubitorum, mensura hominis, quae est angeli.
REV|21|18|Et erat structura muri eius ex iaspide, ipsa vero civitas aurum mundum simile vitro mundo.
REV|21|19|Fundamenta muri civitatis omni lapide pretioso ornata: fundamentum primum iaspis, secundus sapphirus, tertius chalcedonius, quartus smaragdus,
REV|21|20|quintus sardonyx, sextus sardinus, septimus chrysolithus, octavus beryllus, nonus topazius, decimus chrysoprasus, undecimus hyacinthus, duodecimus amethystus.
REV|21|21|Et duodecim portae duodecim margaritae sunt, et singulae portae erant ex singulis margaritis. Et platea civitatis aurum mundum tamquam vitrum perlucidum.
REV|21|22|Et templum non vidi in ea: Dominus enim, Deus omnipotens, templum illius est, et Agnus.
REV|21|23|Et civitas non eget sole neque luna, ut luceant ei, nam claritas Dei illuminavit eam, et lucerna eius est Agnus.
REV|21|24|Et ambulabunt gentes per lumen eius, et reges terrae afferunt gloriam suam in illam;
REV|21|25|et portae eius non claudentur per diem, nox enim non erit illic;
REV|21|26|et afferent gloriam et divitias gentium in illam.
REV|21|27|Nec intrabit in ea aliquid coinquinatum et faciens abominationem et mendacium, nisi qui scripti sunt in libro vitae Agni.
REV|22|1|Et ostendit mihi fluvium aquae vitae splendidum tamquam crystallum, procedentem de throno Dei et Agni.
REV|22|2|In medio plateae eius et fluminis ex utraque parte lignum vitae afferens fructus duodecim, per menses singulos reddens fructum suum; et folia ligni ad sanitatem gentium.
REV|22|3|Et omne maledictum non erit amplius. Et thronus Dei et Agni in illa erit; et servi eius servient illi
REV|22|4|et videbunt faciem eius, et nomen eius in frontibus eorum.
REV|22|5|Et nox ultra non erit, et non egent lumine lucernae neque lumine solis, quoniam Dominus Deus illuminabit super illos, et regnabunt in saecula saeculorum.
REV|22|6|Et dixit mihi: " Haec verba fidelissima et vera sunt, et Dominus, Deus spirituum prophetarum, misit angelum suum ostendere servis suis, quae oportet fieri cito.
REV|22|7|Et ecce venio velociter. Beatus, qui servat verba prophetiae libri huius.
REV|22|8|Et ego Ioannes, qui audivi et vidi haec. Et postquam audissem et vidissem, cecidi, ut adorarem ante pedes angeli, qui mihi haec ostendebat.
REV|22|9|Et dicit mihi: " Vide, ne feceris. Conservus tuus sum et fratrum tuorum prophetarum et eorum, qui servant verba libri huius; Deum adora! ".
REV|22|10|Et dicit mihi: " Ne signaveris verba prophetiae libri huius; tempus enim prope est!
REV|22|11|Qui nocet, noceat adhuc; et, qui sordidus est, sordescat adhuc; et iustus iustitiam faciat adhuc; et sanctus sanctificetur adhuc.
REV|22|12|Ecce venio cito, et merces mea mecum est, reddere unicuique sicut opus eius est.
REV|22|13|Ego Alpha et Omega, primus et novissimus, principium et finis.
REV|22|14|Beati, qui lavant stolas suas, ut sit potestas eorum super lignum vitae, et per portas intrent in civitatem.
REV|22|15|Foris canes et venefici et impudici et homicidae et idolis servientes et omnis, qui amat et facit mendacium!
REV|22|16|Ego Iesus misi angelum meum testificari vobis haec super ecclesiis. Ego sum radix et genus David, stella splendida matutina ".
REV|22|17|Et Spiritus et sponsa dicunt: " Veni! ". Et, qui audit, dicat: " Veni!. Et, qui sitit, veniat; qui vult, accipiat aquam vitae gratis.
REV|22|18|Contestor ego omni audienti verba prophetiae libri huius: Si quis apposuerit ad haec, apponet Deus super illum plagas scriptas in libro isto;
REV|22|19|et si quis abstulerit de verbis libri prophetiae huius, auferet Deus partem eius de ligno vitae et de civitate sancta, de his, quae scripta sunt in libro isto.
REV|22|20|Dicit, qui testimonium perhibet istorum: " Etiam, venio cito ". Amen. Veni, Domine Iesu! ".
REV|22|21|Gratia Domini Iesu cum omnibus.
