2THESS|1|1|Paulus et Silvanus et Timo theus ecclesiae Thessalonicen sium in Deo Patre nostro et Domino Iesu Christo:
2THESS|1|2|gratia vobis et pax a Deo Patre nostro et Domino Iesu Christo.
2THESS|1|3|Gratias agere debemus Deo semper pro vobis, fratres, sicut dignum est, quoniam supercrescit fides vestra, et abundat caritas uniuscuiusque omnium vestrum in invicem,
2THESS|1|4|ita ut et nos ipsi in vobis gloriemur in ecclesiis Dei pro patientia vestra et fide in omnibus persecutionibus vestris et tribulationibus, quas sustinetis,
2THESS|1|5|indicium iusti iudicii Dei, ut digni habeamini regno Dei, pro quo et patimini;
2THESS|1|6|si quidem iustum est apud Deum retribuere tribulationem his, qui vos tribulant,
2THESS|1|7|et vobis, qui tribulamini, requiem nobiscum in revelatione Domini Iesu de caelo cum angelis virtutis eius,
2THESS|1|8|in igne flammae, dantis vindictam his, qui non noverunt Deum et qui non oboediunt evangelio Domini nostri Iesu;
2THESS|1|9|qui poenas dabunt interitu aeterno a facie Domini et a gloria virtutis eius,
2THESS|1|10|cum venerit glorificari in sanctis suis et admirabilis fieri in omnibus, qui crediderunt; quia creditum est testimonium nostrum super vos in die illo.
2THESS|1|11|Ad quod etiam oramus semper pro vobis, ut dignetur vos vocatione sua Deus noster et impleat omnem voluntatem bonitatis et opus fidei in virtute;
2THESS|1|12|ut glorificetur nomen Domini nostri Iesu Christi in vobis, et vos in illo, secundum gratiam Dei nostri et Domini Iesu Christi.
2THESS|2|1|Rogamus autem vos, fratres, circa adventum Domini nostri Iesu Christi et nostram congregationem in ipsum,
2THESS|2|2|ut non cito moveamini a sensu neque terreamini, neque per spiritum neque per verbum neque per epistulam tamquam per nos, quasi instet dies Domini.
2THESS|2|3|Ne quis vos seducat ullo modo; quoniam, nisi venerit discessio primum, et revelatus fuerit homo iniquitatis, filius perditionis,
2THESS|2|4|qui adversatur et extollitur supra omne, quod dicitur Deus aut quod colitur, ita ut in templo Dei sedeat, ostendens se quia sit Deus.
2THESS|2|5|Non retinetis quod, cum adhuc essem apud vos, haec dicebam vobis?
2THESS|2|6|Et nunc quid detineat scitis, ut ipse reveletur in suo tempore.
2THESS|2|7|Nam mysterium iam operatur iniquitatis; tantum qui tenet nunc, donec de medio fiat.
2THESS|2|8|Et tunc revelabitur ille iniquus, quem Dominus Iesus interficiet spiritu oris sui et destruet illustratione adventus sui,
2THESS|2|9|eum, cuius est adventus secundum operationem Satanae in omni virtute et signis et prodigiis mendacibus
2THESS|2|10|et in omni seductione iniquitatis his, qui pereunt, eo quod caritatem veritatis non receperunt, ut salvi fierent.
2THESS|2|11|Et ideo mittit illis Deus operationem erroris, ut credant mendacio,
2THESS|2|12|ut iudicentur omnes, qui non crediderunt veritati, sed consenserunt iniquitati.
2THESS|2|13|Nos autem debemus gratias agere Deo semper pro vobis, fratres, dilecti a Domino, quod elegerit vos Deus primitias in salutem, in sanctificatione Spiritus et fide veritatis;
2THESS|2|14|ad quod et vocavit vos per evangelium nostrum in acquisitionem gloriae Domini nostri Iesu Christi.
2THESS|2|15|Itaque, fratres, state et tenete traditiones, quas didicistis sive per sermonem sive per epistulam nostram.
2THESS|2|16|Ipse autem Dominus noster Iesus Christus et Deus Pater noster, qui dilexit nos et dedit consolationem aeternam et spem bonam in gratia,
2THESS|2|17|consoletur corda vestra et confirmet in omni opere et sermone bono.
2THESS|3|1|De cetero, fratres, orate pro nobis, ut sermo Domini currat et glorificetur sicut et apud vos,
2THESS|3|2|et ut liberemur ab importunis et malis hominibus; non enim omnium est fides.
2THESS|3|3|Fidelis autem Dominus est, qui confirmabit vos et custodiet a Malo.
2THESS|3|4|Confidimus autem de vobis in Domino, quoniam, quae praecipimus, et facitis et facietis.
2THESS|3|5|Dominus autem dirigat corda vestra in caritatem Dei et patientiam Christi.
2THESS|3|6|Praecipimus autem vobis, fratres, in nomine Domini nostri Iesu Christi, ut subtrahatis vos ab omni fratre ambulante inordinate et non secundum traditionem, quam acceperunt a nobis.
2THESS|3|7|Ipsi enim scitis quemadmodum oporteat imitari nos, quoniam non inordinati fuimus inter vos
2THESS|3|8|neque gratìs panem manducavimus ab aliquo sed in labore et fatigatione, nocte et die operantes, ne quem vestrum gravaremus;
2THESS|3|9|non quasi non habuerimus potestatem, sed ut nosmetipsos formam daremus vobis ad imitandum nos.
2THESS|3|10|Nam et cum essemus apud vos, hoc praecipiebamus vobis: Si quis non vult operari, nec manducet.
2THESS|3|11|Audimus enim inter vos quosdam ambulare inordinate, nihil operantes sed curiose agentes;
2THESS|3|12|his autem, qui eiusmodi sunt, praecipimus et obsecramus in Domino Iesu Christo, ut cum quiete operantes suum panem manducent.
2THESS|3|13|Vos autem, fratres, nolite deficere benefacientes.
2THESS|3|14|Quod si quis non oboedit verbo nostro per epistulam, hunc notate, non commisceamini cum illo, ut confundatur;
2THESS|3|15|et nolite quasi inimicum existimare, sed corripite ut fratrem.
2THESS|3|16|Ipse autem Dominus pacis det vobis pacem sempiternam in omni modo. Dominus cum omnibus vobis.
2THESS|3|17|Salutatio mea manu Pauli, quod est signum in omni epistula; ita scribo.
2THESS|3|18|Gratia Domini nostri Iesu Christi cum omnibus vobis.
