TITUS|1|1|Павло, раб Божий, а апостол Ісуса Христа, по вірі вибраних Божих і пізнанні правди, що за благочестям,
TITUS|1|2|в надії вічного життя, яке обіцяв був від вічних часів необманливий Бог,
TITUS|1|3|і часу свого з'явив Слово Своє в проповіданні, що доручене було мені з наказу Спасителя нашого Бога,
TITUS|1|4|до Тита, щирого сина за спільною вірою: благодать, милість та мир від Бога Отця й Христа Ісуса, Спасителя нашого!
TITUS|1|5|Я для того тебе полишив був у Кріті, щоб ти впорядкував недокінчене та пресвітерів настановив по містах, як тобі я звелів,
TITUS|1|6|коли хто бездоганний, муж єдиної дружини, має вірних дітей, недокорених за блуд або неслухняність.
TITUS|1|7|Бо єпископ мусить бути бездоганний, як Божий доморядник, не самолюбний, не гнівливий, не п'яниця, не заводіяка, не корисливий,
TITUS|1|8|але гостинний до приходнів, добролюбець, поміркований, справедливий, побожний, стриманий,
TITUS|1|9|що тримається вірного слова згідно з наукою, щоб мав силу й навчати в здоровій науці, і переконувати противних.
TITUS|1|10|Багато бо є неслухняних, марнословців, зводників, особливо ж з обрізаних,
TITUS|1|11|їм треба уста затуляти: вони цілі доми баламутять, навчаючи, чого не належить, для зиску брудного.
TITUS|1|12|Сказав один з них, їхній власний пророк: Крітяни завжди брехливі, люті звірі, черевані ліниві!...
TITUS|1|13|Це свідоцтво правдиве. Ради цієї причини докоряй їм суворо, щоб у вірі здорові були,
TITUS|1|14|і на юдейські байки не вважали, ані на накази людей, що від правди відвертаються.
TITUS|1|15|Для чистих все чисте, а для занечищених та для невірних не чисте ніщо, але занечистилися і розум їхній, і сумління.
TITUS|1|16|Вони твердять, немов знають Бога, але відкидаються вчинками, бувши бридкі й неслухняні, і до всякого доброго діла нездатні.
TITUS|2|1|А ти говори, що відповідає здоровій науці.
TITUS|2|2|Щоб старі чоловіки тверезі були, поважні, помірковані, здорові у вірі, у любові, у терпеливості.
TITUS|2|3|Щоб старі жінки в своїм стані так само були, як належить святим, не обмовниці, не віддані п'янству, навчали добра,
TITUS|2|4|щоб навчали жінок молодих любити своїх чоловіків, любити дітей,
TITUS|2|5|щоб були помірковані, чисті, господарні, добрі, слухняні своїм чоловікам, щоб не зневажалося Боже Слово.
TITUS|2|6|Так само благай юнаків, щоб були помірковані.
TITUS|2|7|У всім сам себе подавай за зразка добрих діл, у навчанні непорушеність, повагу,
TITUS|2|8|слово здорове, неосудливе, щоб противник був засоромлений, не мавши нічого лихого казати про нас.
TITUS|2|9|Раби щоб корилися панам своїм, щоб догоджали, не перечили,
TITUS|2|10|не крали, але виявляли всяку добру вірність, щоб у всьому вони прикрашали науку Спасителя нашого Бога.
TITUS|2|11|Бо з'явилася Божа благодать, що спасає всіх людей,
TITUS|2|12|і навчає нас, щоб ми, відцуравшись безбожности та світських пожадливостей, жили помірковано та праведно, і побожно в теперішнім віці,
TITUS|2|13|і чекали блаженної надії та з'явлення слави великого Бога й Спаса нашого Христа Ісуса,
TITUS|2|14|що Самого Себе дав за нас, щоб нас визволити від усякого беззаконства та очистити Собі людей вибраних, у добрих ділах запопадливих.
TITUS|2|15|Оце говори та нагадуй, та з усяким наказом картай. Хай тобою ніхто не погордує!
TITUS|3|1|Нагадуй їм, щоб слухали влади верховної та корилися їй, і до всякого доброго діла готові були,
TITUS|3|2|щоб не зневажали нікого, щоб були не сварливі, а тихі, виявляючи повну лагідність усім людям.
TITUS|3|3|Бо колись були й ми нерозсудні, неслухняні, зведені, служили різним пожадливостям та розкошам, жили в злобі та в заздрощах, бридкими були, ненавиділи один одного.
TITUS|3|4|А коли з'явилась благодать та людинолюбство Спасителя, нашого Бога,
TITUS|3|5|Він нас спас не з діл праведности, що ми їх учинили були, а з Своєї милости через купіль відродження й обновлення Духом Святим,
TITUS|3|6|Якого Він щедро вилив на нас через Христа Ісуса, Спасителя нашого,
TITUS|3|7|щоб ми виправдались Його благодаттю, і стали спадкоємцями за надією на вічне життя.
TITUS|3|8|Вірне слово, і я хочу, щоб ти і про це впевняв, щоб ті, хто ввірував у Бога, дбали про добрі діла пильнувати. Для людей оце добре й корисне!
TITUS|3|9|Вистерігайсь нерозумних змагань, і родоводів, і спорів, і суперечок про Закон, бо вони некорисні й марні.
TITUS|3|10|Людини єретика, по першім та другім наставленні, відрікайся,
TITUS|3|11|знавши, що зіпсувся такий та грішить, і він сам себе засудив.
TITUS|3|12|Як пришлю я до тебе Артема або Тихика, поквапся прибути до мене в Нікополь, бо думаю там перезимувати.
TITUS|3|13|Законника Зину та Аполлоса вишли квапливо вперед, щоб для них не забракло нічого.
TITUS|3|14|Нехай же навчаються й наші дбати про добрі діла при конечних потребах, щоб безплодні вони не були.
TITUS|3|15|Вітають тебе всі, хто зо мною. Вітай тих, хто любить нас у вірі. Благодать з вами всіма! Амінь.
