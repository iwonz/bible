1KGS|1|1|Когда царь Давид состарился, вошел в [преклонные] лета, то покрывали его одеждами, но не мог он согреться.
1KGS|1|2|И сказали ему слуги его: пусть поищут для господина нашего царя молодую девицу, чтоб она предстояла царю и ходила за ним и лежала с ним, – и будет тепло господину нашему, царю.
1KGS|1|3|И искали красивой девицы во всех пределах Израильских, и нашли Ависагу Сунамитянку, и привели ее к царю.
1KGS|1|4|Девица была очень красива, и ходила она за царем и прислуживала ему; но царь не познал ее.
1KGS|1|5|Адония, сын Аггифы, возгордившись говорил: я буду царем. И завел себе колесницы и всадников и пятьдесят человек скороходов.
1KGS|1|6|Отец же никогда не стеснял его вопросом: для чего ты это делаешь? Он же был очень красив и родился ему после Авессалома.
1KGS|1|7|И советовался он с Иоавом, сыном Саруиным, и с Авиафаром священником, и они помогали Адонии.
1KGS|1|8|Но священник Садок и Ванея, сын Иодаев, и пророк Нафан, и Семей, и Рисий, и сильные Давидовы не были на стороне Адонии.
1KGS|1|9|И заколол Адония овец и волов и тельцов у камня Зохелет, что у источника Рогель, и пригласил всех братьев своих, сыновей царя, со всеми Иудеянами, служившими у царя.
1KGS|1|10|Пророка же Нафана и Ванею, и тех сильных, и Соломона, брата своего, не пригласил.
1KGS|1|11|Тогда Нафан сказал Вирсавии, матери Соломона, говоря: слышала ли ты, что Адония, сын Аггифин, сделался царем, а господин наш Давид не знает [о том]?
1KGS|1|12|Теперь, вот, я советую тебе: спасай жизнь твою и жизнь сына твоего Соломона.
1KGS|1|13|Иди и войди к царю Давиду и скажи ему: не клялся ли ты, господин мой царь, рабе твоей, говоря: "сын твой Соломон будет царем после меня и он сядет на престоле моем"? Почему же воцарился Адония?
1KGS|1|14|И вот, когда ты еще будешь говорить там с царем, войду и я вслед за тобою и дополню слова твои.
1KGS|1|15|Вирсавия пошла к царю в спальню; царь был очень стар, и Ависага Сунамитянка прислуживала царю;
1KGS|1|16|и наклонилась Вирсавия и поклонилась царю; и сказал царь: что тебе?
1KGS|1|17|Она сказала ему: господин мой царь! ты клялся рабе твоей Господом Богом твоим: "сын твой Соломон будет царствовать после меня и он сядет на престоле моем".
1KGS|1|18|А теперь, вот, Адония [воцарился], и ты, господин мой царь, не знаешь [о том].
1KGS|1|19|И заколол он множество волов, тельцов и овец, и пригласил всех сыновей царских и священника Авиафара, и военачальника Иоава; Соломона же, раба твоего, не пригласил.
1KGS|1|20|Но ты, господин мой, – царь, и глаза всех Израильтян [устремлены] на тебя, чтобы ты объявил им, кто сядет на престоле господина моего царя после него;
1KGS|1|21|иначе, когда господин мой царь почиет с отцами своими, падет обвинение на меня и на сына моего Соломона.
1KGS|1|22|Когда она еще говорила с царем, пришел и пророк Нафан.
1KGS|1|23|И сказали царю, говоря: вот Нафан пророк. И вошел он к царю и поклонился царю лицем до земли.
1KGS|1|24|И сказал Нафан: господин мой царь! сказал ли ты: "Адония будет царствовать после меня и он сядет на престоле моем"?
1KGS|1|25|Потому что он ныне сошел и заколол множество волов, тельцов и овец, и пригласил всех сыновей царских и военачальников и священника Авиафара, и вот, они едят и пьют у него и говорят: да живет царь Адония!
1KGS|1|26|А меня, раба твоего, и священника Садока, и Ванею, сына Иодаева, и Соломона, раба твоего, не пригласил.
1KGS|1|27|Не сталось ли это по [воле] господина моего царя, и для чего ты не открыл рабу твоему, кто сядет на престоле господина моего царя после него?
1KGS|1|28|И отвечал царь Давид и сказал: позовите ко мне Вирсавию. И вошла она и стала пред царем.
1KGS|1|29|И клялся царь и сказал: жив Господь, избавлявший душу мою от всякой беды!
1KGS|1|30|Как я клялся тебе Господом Богом Израилевым, говоря, что Соломон, сын твой, будет царствовать после меня и он сядет на престоле моем вместо меня, так я и сделаю это сегодня.
1KGS|1|31|И наклонилась Вирсавия лицем до земли, и поклонилась царю, и сказала: да живет господин мой царь Давид во веки!
1KGS|1|32|И сказал царь Давид: позовите ко мне священника Садока и пророка Нафана и Ванею, сына Иодаева. И вошли они к царю.
1KGS|1|33|И сказал им царь: возьмите с собою слуг господина вашего и посадите Соломона, сына моего, на мула моего, и сведите его к Гиону,
1KGS|1|34|и да помажет его там Садок священник и Нафан пророк в царя над Израилем, и затрубите трубою и возгласите: да живет царь Соломон!
1KGS|1|35|Потом проводите его назад, и он придет и сядет на престоле моем; он будет царствовать вместо меня; ему завещал я быть вождем Израиля и Иуды.
1KGS|1|36|И отвечал Ванея, сын Иодаев, царю и сказал: аминь, – да скажет так Господь Бог господина моего царя!
1KGS|1|37|Как был Господь Бог с господином моим царем, так да будет Он с Соломоном и да возвеличит престол его более престола господина моего царя Давида!
1KGS|1|38|И пошли Садок священник и Нафан пророк и Ванея, сын Иодая, и Хелефеи и Фелефеи, и посадили Соломона на мула царя Давида, и повели его к Гиону.
1KGS|1|39|И взял Садок священник рог с елеем из скинии и помазал Соломона. И затрубили трубою, и весь народ восклицал: да живет царь Соломон!
1KGS|1|40|И весь народ провожал Соломона, и играл народ на свирелях, и весьма радовался, так что земля расседалась от криков его.
1KGS|1|41|И услышал Адония и все приглашенные им, как только перестали есть; а Иоав, услышав звук трубы, сказал: отчего этот шум волнующегося города?
1KGS|1|42|Еще он говорил, как пришел Ионафан, сын священника Авиафара. И сказал Адония: войди; ты – честный человек и несешь добрую весть.
1KGS|1|43|И отвечал Ионафан и сказал Адонии: да, господин наш царь Давид поставил Соломона царем;
1KGS|1|44|и послал царь с ним Садока священника и Нафана пророка, и Ванею, сына Иодая, и Хелефеев и Фелефеев, и они посадили его на мула царского;
1KGS|1|45|и помазали его Садок священник и Нафан пророк в царя в Гионе, и оттуда отправились с радостью, и пришел в движение город. Вот отчего шум, который вы слышите.
1KGS|1|46|И Соломон уже сел на царском престоле.
1KGS|1|47|И слуги царя приходили поздравить господина нашего царя Давида, говоря: Бог твой да прославит имя Соломона более твоего имени и да возвеличит престол его более твоего престола. И поклонился царь на ложе своем,
1KGS|1|48|и сказал царь так: "благословен Господь Бог Израилев, Который сегодня дал сидящего на престоле моем, и очи мои видят это!"
1KGS|1|49|[Тогда] испугались и встали все приглашенные, которые были у Адонии, и пошли каждый своею дорогою.
1KGS|1|50|Адония же, боясь Соломона, встал и пошел и ухватился за роги жертвенника.
1KGS|1|51|И донесли Соломону, говоря: вот, Адония боится царя Соломона, и вот, он держится за роги жертвенника, говоря: пусть поклянется мне теперь царь Соломон, что он не умертвит раба своего мечом.
1KGS|1|52|И сказал Соломон: если он будет человеком честным, то ни один волос его не упадет на землю; если же найдется в нем лукавство, то умрет.
1KGS|1|53|И послал царь Соломон, и привели его от жертвенника. И он пришел и поклонился царю Соломону; и сказал ему Соломон: иди в дом свой.
1KGS|2|1|Приблизилось время умереть Давиду, и завещал он сыну своему Соломону, говоря:
1KGS|2|2|вот, я отхожу в путь всей земли, ты же будь тверд и будь мужествен
1KGS|2|3|и храни завет Господа Бога твоего, ходя путями Его и соблюдая уставы Его и заповеди Его, и определения Его и постановления Его, как написано в законе Моисеевом, чтобы быть тебе благоразумным во всем, что ни будешь делать, и везде, куда ни обратишься;
1KGS|2|4|чтобы Господь исполнил слово Свое, которое Он сказал обо мне, говоря: "если сыны твои будут наблюдать за путями своими, чтобы ходить предо Мною в истине от всего сердца своего и от всей души своей, то не прекратится муж от тебя на престоле Израилевом".
1KGS|2|5|Еще: ты знаешь, что сделал мне Иоав, сын Саруин, как поступил он с двумя вождями войска Израильского, с Авениром, сыном Нировым, и Амессаем, сыном Иеферовым, как он умертвил их и пролил кровь бранную во время мира, обагрив кровью бранною пояс на чреслах своих и обувь на ногах своих:
1KGS|2|6|поступи по мудрости твоей, чтобы не отпустить седины его мирно в преисподнюю.
1KGS|2|7|А сынам Верзеллия Галаадитянина окажи милость, чтоб они были между питающимися твоим столом, ибо они пришли ко мне, когда я бежал от Авессалома, брата твоего.
1KGS|2|8|Вот еще у тебя Семей, сын Геры Вениамитянина из Бахурима; он злословил меня тяжким злословием, когда я шел в Маханаим; но он вышел навстречу мне у Иордана, и я поклялся ему Господом, говоря: "я не умерщвлю тебя мечом".
1KGS|2|9|Ты же не оставь его безнаказанным; ибо ты человек мудрый и знаешь, что тебе сделать с ним, чтобы низвести седину его в крови в преисподнюю.
1KGS|2|10|И почил Давид с отцами своими и погребен был в городе Давидовом.
1KGS|2|11|Времени царствования Давида над Израилем было сорок лет: в Хевроне царствовал он семь лет и тридцать три года царствовал в Иерусалиме.
1KGS|2|12|И сел Соломон на престоле Давида, отца своего, и царствование его было очень твердо.
1KGS|2|13|И пришел Адония, сын Аггифы, к Вирсавии, матери Соломона. Она сказала: с миром ли приход твой? И сказал он: с миром.
1KGS|2|14|И сказал он: у меня есть слово к тебе. Она сказала: говори.
1KGS|2|15|И сказал он: ты знаешь, что царство принадлежало мне, и весь Израиль обращал на меня взоры свои, как на будущего царя; но царство отошло от меня и досталось брату моему, ибо от Господа это было ему;
1KGS|2|16|теперь я прошу тебя об одном, не откажи мне. Она сказала ему: говори.
1KGS|2|17|И сказал он: прошу тебя, поговори царю Соломону, ибо он не откажет тебе, чтоб он дал мне Ависагу Сунамитянку в жену.
1KGS|2|18|И сказала Вирсавия: хорошо, я поговорю о тебе царю.
1KGS|2|19|И вошла Вирсавия к царю Соломону говорить ему об Адонии. Царь встал перед нею, и поклонился ей, и сел на престоле своем. Поставили престол и для матери царя, и она села по правую руку его
1KGS|2|20|и сказала: я имею к тебе одну небольшую просьбу, не откажи мне. И сказал ей царь: проси, мать моя; я не откажу тебе.
1KGS|2|21|И сказала она: дай Ависагу Сунамитянку Адонии, брату твоему, в жену.
1KGS|2|22|И отвечал царь Соломон и сказал матери своей: а зачем ты просишь Ависагу Сунамитянку для Адонии? проси ему [также] и царства; ибо он мой старший брат, и ему священник Авиафар и Иоав, сын Саруин, [друг].
1KGS|2|23|И поклялся царь Соломон Господом, говоря: то и то пусть сделает со мною Бог и еще больше сделает, если не на свою душу сказал Адония такое слово;
1KGS|2|24|ныне же, – жив Господь, укрепивший меня и посадивший меня на престоле Давида, отца моего, и устроивший мне дом, как говорил Он, – ныне же Адония должен умереть.
1KGS|2|25|И послал царь Соломон Ванею, сына Иодаева, который поразил его, и он умер.
1KGS|2|26|А священнику Авиафару царь сказал: ступай в Анафоф на твое поле; ты достоин смерти, но в настоящее время я не умерщвлю тебя, ибо ты носил ковчег Владыки Господа пред Давидом, отцом моим, и терпел все, что терпел отец мой.
1KGS|2|27|И удалил Соломон Авиафара от священства Господня, и исполнилось слово Господа, которое сказал Он о доме Илия в Силоме.
1KGS|2|28|Слух [об этом] дошел до Иоава, – так как Иоав склонялся на сторону Адонии, а на сторону Соломона не склонялся, – и убежал Иоав в скинию Господню и ухватился за роги жертвенника.
1KGS|2|29|И донесли царю Соломону, что Иоав убежал в скинию Господню и что он у жертвенника. И послал Соломон Ванею, сына Иодаева, говоря: пойди, умертви его.
1KGS|2|30|И пришел Ванея в скинию Господню и сказал ему: так сказал царь: выходи. И сказал тот: нет, я хочу умереть здесь. Ванея передал это царю, говоря: так сказал Иоав, и так отвечал мне.
1KGS|2|31|Царь сказал ему: сделай, как он сказал, и умертви его и похорони его, и сними невинную кровь, пролитую Иоавом, с меня и с дома отца моего;
1KGS|2|32|да обратит Господь кровь его на голову его за то, что он убил двух мужей невинных и лучших его: поразил мечом, без ведома отца моего Давида, Авенира, сына Нирова, военачальника Израильского, и Амессая, сына Иеферова, военачальника Иудейского;
1KGS|2|33|да обратится кровь их на голову Иоава и на голову потомства его на веки, а Давиду и потомству его, и дому его и престолу его да будет мир на веки от Господа!
1KGS|2|34|И пошел Ванея, сын Иодаев, и поразил Иоава, и умертвил его, и он был похоронен в доме своем в пустыне.
1KGS|2|35|И поставил царь Соломон Ванею, сына Иодаева, вместо его над войском; а Садока священника поставил царь вместо Авиафара.
1KGS|2|36|И послав царь призвал Семея и сказал ему: построй себе дом в Иерусалиме и живи здесь, и никуда не выходи отсюда;
1KGS|2|37|и знай, что в тот день, в который ты выйдешь и перейдешь поток Кедрон, непременно умрешь; кровь твоя будет на голове твоей.
1KGS|2|38|И сказал Семей царю: хорошо; как приказал господин мой царь, так сделает раб твой. И жил Семей в Иерусалиме долгое время.
1KGS|2|39|Но через три года случилось, что у Семея двое рабов убежали к Анхусу, сыну Маахи, царю Гефскому. И сказали Семею, говоря: вот, рабы твои в Гефе.
1KGS|2|40|И встал Семей, и оседлал осла своего, и отправился в Геф к Анхусу искать рабов своих. И возвратился Семей и привел рабов своих из Гефа.
1KGS|2|41|И донесли Соломону, что Семей ходил из Иерусалима в Геф и возвратился.
1KGS|2|42|И послав призвал царь Семея и сказал ему: не клялся ли я тебе Господом и не объявлял ли тебе, говоря: "знай, что в тот день, в который ты выйдешь и пойдешь куда–нибудь, непременно умрешь"? и ты сказал мне: "хорошо";
1KGS|2|43|зачем же ты не соблюл приказания, которое я дал тебе пред Господом с клятвою?
1KGS|2|44|И сказал царь Семею: ты знаешь и знает сердце твое все зло, какое ты сделал отцу моему Давиду; да обратит же Господь злобу твою на голову твою!
1KGS|2|45|а царь Соломон да будет благословен, и престол Давида да будет непоколебим пред Господом во веки!
1KGS|2|46|и повелел царь Ванее, сыну Иодаеву, и он пошел и поразил Семея, и тот умер.
1KGS|3|1|Соломон породнился с фараоном, царем Египетским, и взял за себя дочь фараона и ввел ее в город Давидов, доколе не построил дома своего и дома Господня и стены вокруг Иерусалима.
1KGS|3|2|Народ еще приносил жертвы на высотах, ибо не был построен дом имени Господа до того времени.
1KGS|3|3|И возлюбил Соломон Господа, ходя по уставу Давида, отца своего; но и он приносил жертвы и курения на высотах.
1KGS|3|4|И пошел царь в Гаваон, чтобы принести там жертву, ибо там был главный жертвенник. Тысячу всесожжений вознес Соломон на том жертвеннике.
1KGS|3|5|В Гаваоне явился Господь Соломону во сне ночью, и сказал Бог: проси, что дать тебе.
1KGS|3|6|И сказал Соломон: Ты сделал рабу Твоему Давиду, отцу моему, великую милость; и за то, что он ходил пред Тобою в истине и правде и с искренним сердцем пред Тобою, Ты сохранил ему эту великую милость и даровал ему сына, который сидел бы на престоле его, как это и есть ныне;
1KGS|3|7|и ныне, Господи Боже мой, Ты поставил раба Твоего царем вместо Давида, отца моего; но я отрок малый, не знаю ни моего выхода, ни входа;
1KGS|3|8|и раб Твой – среди народа Твоего, который избрал Ты, народа столь многочисленного, что по множеству его нельзя ни исчислить его, ни обозреть;
1KGS|3|9|даруй же рабу Твоему сердце разумное, чтобы судить народ Твой и различать, что добро и что зло; ибо кто может управлять этим многочисленным народом Твоим?
1KGS|3|10|И благоугодно было Господу, что Соломон просил этого.
1KGS|3|11|И сказал ему Бог: за то, что ты просил этого и не просил себе долгой жизни, не просил себе богатства, не просил себе душ врагов твоих, но просил себе разума, чтоб уметь судить, –
1KGS|3|12|вот, Я сделаю по слову твоему: вот, Я даю тебе сердце мудрое и разумное, так что подобного тебе не было прежде тебя, и после тебя не восстанет подобный тебе;
1KGS|3|13|и то, чего ты не просил, Я даю тебе, и богатство и славу, так что не будет подобного тебе между царями во все дни твои;
1KGS|3|14|и если будешь ходить путем Моим, сохраняя уставы Мои и заповеди Мои, как ходил отец твой Давид, Я продолжу и дни твои.
1KGS|3|15|И пробудился Соломон, и вот, [это было] сновидение. И пошел он в Иерусалим и стал пред ковчегом завета Господня, и принес всесожжения и совершил [жертвы] мирные, и сделал большой пир для всех слуг своих.
1KGS|3|16|Тогда пришли две женщины блудницы к царю и стали пред ним.
1KGS|3|17|И сказала одна женщина: о, господин мой! я и эта женщина живем в одном доме; и я родила при ней в этом доме;
1KGS|3|18|на третий день после того, как я родила, родила и эта женщина; и были мы вместе, и в доме никого постороннего с нами не было; только мы две были в доме;
1KGS|3|19|и умер сын этой женщины ночью, ибо она заспала его;
1KGS|3|20|и встала она ночью, и взяла сына моего от меня, когда я, раба твоя, спала, и положила его к своей груди, а своего мертвого сына положила к моей груди;
1KGS|3|21|утром я встала, чтобы покормить сына моего, и вот, он был мертвый; а когда я всмотрелась в него утром, то это был не мой сын, которого я родила.
1KGS|3|22|И сказала другая женщина: нет, мой сын живой, а твой сын мертвый. А та говорила ей: нет, твой сын мертвый, а мой живой. И говорили они так пред царем.
1KGS|3|23|И сказал царь: эта говорит: мой сын живой, а твой сын мертвый; а та говорит: нет, твой сын мертвый, а мой сын живой.
1KGS|3|24|И сказал царь: подайте мне меч. И принесли меч к царю.
1KGS|3|25|И сказал царь: рассеките живое дитя надвое и отдайте половину одной и половину другой.
1KGS|3|26|И отвечала та женщина, которой сын был живой, царю, ибо взволновалась вся внутренность ее от жалости к сыну своему: о, господин мой! отдайте ей этого ребенка живого и не умерщвляйте его. А другая говорила: пусть же не будет ни мне, ни тебе, рубите.
1KGS|3|27|И отвечал царь и сказал: отдайте этой живое дитя, и не умерщвляйте его: она – его мать.
1KGS|3|28|И услышал весь Израиль о суде, как рассудил царь; и стали бояться царя, ибо увидели, что мудрость Божия в нем, чтобы производить суд.
1KGS|4|1|И был царь Соломон царем над всем Израилем.
1KGS|4|2|И вот начальники, которые [были] у него: Азария, сын Садока священника;
1KGS|4|3|Елихореф и Ахия, сыновья Сивы, писцы; Иосафат, сын Ахилуда, дееписатель;
1KGS|4|4|Ванея, сын Иодая, военачальник; Садок и Авиафар – священники;
1KGS|4|5|Азария, сын Нафана, начальник над приставниками, и Завуф, сын Нафана священника – друг царя;
1KGS|4|6|Ахисар – начальник над домом [царским], и Адонирам, сын Авды, – над податями.
1KGS|4|7|И было у Соломона двенадцать приставников над всем Израилем, и они доставляли продовольствие царю и дому его; каждый должен был доставлять продовольствие на один месяц в году.
1KGS|4|8|Вот имена их: Бен–Хур – на горе Ефремовой;
1KGS|4|9|Бен–Декер– в Макаце и в Шаалбиме, в Вефсамисе и в Елоне и в Беф–Ханане;
1KGS|4|10|Бен–Хесед – в Арюбофе; ему же принадлежал Соко и вся земля Хефер;
1KGS|4|11|Бен–Авинадав – [над] всем Нафаф–Дором; Тафафь, дочь Соломона, была его женою;
1KGS|4|12|Ваана, сын Ахилуда, в Фаанахе и Мегиддо и во всем Беф–Сане, что близ Цартана ниже Иезрееля, от Беф–Сана до Абел–Мехола, и даже за Иокмеам;
1KGS|4|13|Бен–Гевер – в Рамофе Галаадском; у него были селения Иаира, сына Манассиина, что в Галааде; у него также область Аргов, что в Васане, шестьдесят больших городов со стенами и медными затворами;
1KGS|4|14|Ахинадав, сын Гиддо, в Маханаиме;
1KGS|4|15|Ахимаас – в [земле] Неффалимовой; он взял себе в жену Васемафу, дочь Соломона;
1KGS|4|16|Ваана, сын Хушая, в [земле] Асировой и в Баалофе;
1KGS|4|17|Иосафат, сын Паруаха, в [земле] Иссахаровой;
1KGS|4|18|Шимей, сын Елы, в [земле] Вениаминовой;
1KGS|4|19|Гевер, сын Урия, в земле Галаадской, в земле Сигона, царя Аморрейского, и Ога, царя Васанского. Он был приставник в этой земле.
1KGS|4|20|Иуда и Израиль, многочисленные как песок у моря, ели, пили и веселились.
1KGS|4|21|Соломон владел всеми царствами от реки [Евфрата] до земли Филистимской и до пределов Египта. Они приносили дары и служили Соломону во все дни жизни его.
1KGS|4|22|Продовольствие Соломона на каждый день составляли: тридцать коров муки пшеничной и шестьдесят коров прочей муки,
1KGS|4|23|десять волов откормленных и двадцать волов с пастбища, и сто овец, кроме оленей, и серн, и сайгаков, и откормленных птиц;
1KGS|4|24|ибо он владычествовал над всею землею по эту сторону реки, от Типсаха до Газы, над всеми царями по эту сторону реки, и был у него мир со всеми окрестными странами.
1KGS|4|25|И жили Иуда и Израиль спокойно, каждый под виноградником своим и под смоковницею своею, от Дана до Вирсавии, во все дни Соломона.
1KGS|4|26|И было у Соломона сорок тысяч стойл для коней колесничных и двенадцать тысяч для конницы.
1KGS|4|27|И те приставники доставляли царю Соломону все принадлежащее к столу царя, каждый в свой месяц, и не допускали недостатка ни в чем.
1KGS|4|28|И ячмень и солому для коней и для мулов доставляли каждый в свою очередь на место, где находился царь.
1KGS|4|29|И дал Бог Соломону мудрость и весьма великий разум, и обширный ум, как песок на берегу моря.
1KGS|4|30|И была мудрость Соломона выше мудрости всех сынов востока и всей мудрости Египтян.
1KGS|4|31|Он был мудрее всех людей, мудрее и Ефана Езрахитянина, и Емана, и Халкола, и Дарды, сыновей Махола, и имя его было в славе у всех окрестных народов.
1KGS|4|32|И изрек он три тысячи притчей, и песней его было тысяча и пять;
1KGS|4|33|и говорил он о деревах, от кедра, что в Ливане, до иссопа, вырастающего из стены; говорил и о животных, и о птицах, и о пресмыкающихся, и о рыбах.
1KGS|4|34|И приходили от всех народов послушать мудрости Соломона, от всех царей земных, которые слышали о мудрости его.
1KGS|5|1|И послал Хирам, царь Тирский, слуг своих к Соломону, когда услышал, что его помазали в царя на место отца его; ибо Хирам был другом Давида во всю жизнь.
1KGS|5|2|И послал также и Соломон к Хираму сказать:
1KGS|5|3|ты знаешь, что Давид, отец мой, не мог построить дом имени Господа Бога своего по причине войн с окрестными народами, доколе Господь не покорил их под стопы ног его;
1KGS|5|4|ныне же Господь Бог мой даровал мне покой отовсюду: нет противника и нет более препон;
1KGS|5|5|и вот, я намерен построить дом имени Господа Бога моего, как сказал Господь отцу моему Давиду, говоря: "сын твой, которого Я посажу вместо тебя на престоле твоем, он построит дом имени Моему";
1KGS|5|6|итак прикажи нарубить для меня кедров с Ливана; и вот, рабы мои будут вместе с твоими рабами, и я буду давать тебе плату за рабов твоих, какую ты назначишь; ибо ты знаешь, что у нас нет людей, которые умели бы рубить дерева так, как Сидоняне.
1KGS|5|7|Когда услышал Хирам слова Соломона, очень обрадовался и сказал: благословен ныне Господь, Который дал Давиду сына мудрого [для] [управления] этим многочисленным народом!
1KGS|5|8|И послал Хирам к Соломону сказать: я выслушал то, за чем ты посылал ко мне, и исполню все желание твое о деревах кедровых и деревах кипарисовых;
1KGS|5|9|рабы мои свезут их с Ливана к морю, и я плотами доставлю их морем к месту, которое ты назначишь мне, и там сложу их, и ты возьмешь; но и ты исполни мое желание, чтобы доставлять хлеб для моего дома.
1KGS|5|10|И давал Хирам Соломону дерева кедровые и дерева кипарисовые, вполне по его желанию.
1KGS|5|11|А Соломон давал Хираму двадцать тысяч коров пшеницы для продовольствия дома его и двадцать коров оливкового выбитого масла: столько давал Соломон Хираму каждый год.
1KGS|5|12|Господь дал мудрость Соломону, как обещал ему. И был мир между Хирамом и Соломоном, и они заключили между собою союз.
1KGS|5|13|И обложил царь Соломон повинностью весь Израиль; повинность же состояла в тридцати тысячах человек.
1KGS|5|14|И посылал их на Ливан, по десяти тысяч на месяц, попеременно; месяц они были на Ливане, а два месяца в доме своем. Адонирам же начальствовал над ними.
1KGS|5|15|Еще у Соломона было семьдесят тысяч носящих тяжести и восемьдесят тысяч каменосеков в горах,
1KGS|5|16|кроме трех тысяч трехсот начальников, поставленных Соломоном над работою для надзора за народом, который производил работу.
1KGS|5|17|И повелел царь привозить камни большие, камни дорогие, для основания дома, камни обделанные.
1KGS|5|18|Обтесывали же их работники Соломоновы и работники Хирамовы и Гивлитяне, и приготовляли дерева и камни для строения дома.
1KGS|6|1|В четыреста восьмидесятом году по исшествии сынов Израилевых из земли Египетской, в четвертый год царствования Соломонова над Израилем, в месяц Зиф, который есть второй месяц, начал он строить храм Господу.
1KGS|6|2|Храм, который построил царь Соломон Господу, длиною был в шестьдесят локтей, шириною в двадцать и вышиною в тридцать локтей,
1KGS|6|3|и притвор пред храмом в двадцать локтей длины, соответственно ширине храма, и в десять локтей ширины пред храмом.
1KGS|6|4|И сделал он в доме окна решетчатые, глухие с откосами.
1KGS|6|5|И сделал пристройку вокруг стен храма, вокруг храма и давира; и сделал боковые комнаты кругом.
1KGS|6|6|Нижний [ярус] пристройки шириною был в пять локтей, средний шириною в шесть локтей, а третий шириною в семь локтей; ибо вокруг храма извне сделаны были уступы, дабы пристройка не прикасалась к стенам храма.
1KGS|6|7|Когда строился храм, на строение употребляемы были обтесанные камни; ни молота, ни тесла, ни всякого другого железного орудия не было слышно в храме при строении его.
1KGS|6|8|Вход в средний ярус был с правой стороны храма. По круглым лестницам всходили в средний [ярус], а от среднего в третий.
1KGS|6|9|И построил он храм, и кончил его, и обшил храм кедровыми досками.
1KGS|6|10|И пристроил ко всему храму боковые комнаты вышиною в пять локтей; они прикреплены были к храму посредством кедровых бревен.
1KGS|6|11|И было слово Господа к Соломону, и сказано ему:
1KGS|6|12|вот, ты строишь храм; если ты будешь ходить по уставам Моим, и поступать по определениям Моим и соблюдать все заповеди Мои, поступая по ним, то Я исполню на тебе слово Мое, которое Я сказал Давиду, отцу твоему,
1KGS|6|13|и буду жить среди сынов Израилевых, и не оставлю народа Моего Израиля.
1KGS|6|14|И построил Соломон храм и кончил его.
1KGS|6|15|И обложил стены храма внутри кедровыми досками; от пола храма до потолка внутри обложил деревом и покрыл пол храма кипарисовыми досками.
1KGS|6|16|И устроил в задней стороне храма, в двадцати локтях от края, стену, и обложил стены и потолок кедровыми досками, и устроил давир для Святаго–святых.
1KGS|6|17|Сорока локтей [был] храм, то есть передняя часть храма.
1KGS|6|18|На кедрах внутри храма были вырезаны [подобия] огурцов и распускающихся цветов; все было покрыто кедром, камня не видно было.
1KGS|6|19|Давир же внутри храма он приготовил для того, чтобы поставить там ковчег завета Господня.
1KGS|6|20|И давир был длиною в двадцать локтей, шириною в двадцать локтей и вышиною в двадцать локтей; он обложил его чистым золотом; обложил также и кедровый жертвенник.
1KGS|6|21|И обложил Соломон храм внутри чистым золотом, и протянул золотые цепи пред давиром, и обложил его золотом.
1KGS|6|22|Весь храм он обложил золотом, весь храм до конца, и весь жертвенник, который пред давиром, обложил золотом.
1KGS|6|23|И сделал в давире двух херувимов из масличного дерева, вышиною в десять локтей.
1KGS|6|24|Одно крыло херувима было в пять локтей и другое крыло херувима в пять локтей; десять локтей было от одного конца крыльев его до другого конца крыльев его.
1KGS|6|25|В десять локтей [был] и другой херувим; одинаковой меры и одинакового вида [были] оба херувима.
1KGS|6|26|Высота одного херувима [была] десять локтей, также и другого херувима.
1KGS|6|27|И поставил он херувимов среди внутренней части храма. Крылья же херувимов были распростерты, и касалось крыло одного [одной] стены, а крыло другого херувима касалось другой стены; другие же крылья их среди храма сходились крыло с крылом.
1KGS|6|28|И обложил он херувимов золотом.
1KGS|6|29|И на всех стенах храма кругом сделал резные изображения херувимов и пальмовых дерев и распускающихся цветов, внутри и вне.
1KGS|6|30|И пол в храме обложил золотом во внутренней и передней части.
1KGS|6|31|Для входа в давир сделал двери из масличного дерева, с пятиугольными косяками.
1KGS|6|32|На двух половинах дверей из масличного дерева он сделал резных херувимов и пальмы и распускающиеся цветы и обложил золотом; покрыл золотом и херувимов и пальмы.
1KGS|6|33|И у входа в храм сделал косяки из масличного дерева четырехугольные,
1KGS|6|34|и две двери из кипарисового дерева; обе половинки одной двери были подвижные, и обе половинки другой двери были подвижные.
1KGS|6|35|И вырезал [на них] херувимов и пальмы и распускающиеся цветы и обложил золотом по резьбе.
1KGS|6|36|И построил внутренний двор из трех рядов обтесанного камня и из ряда кедровых брусьев.
1KGS|6|37|В четвертый год, в месяц Зиф, положил он основание храму Господа,
1KGS|6|38|а на одиннадцатом году, в месяце Буле, – это месяц восьмой, – он окончил храм со всеми принадлежностями его и по всем предначертаниям его; строил его семь лет.
1KGS|7|1|А свой дом Соломон строил тринадцать лет и окончил весь дом свой.
1KGS|7|2|И построил он дом из дерева Ливанского, длиною во сто локтей, шириною в пятьдесят локтей, а вышиною в тридцать локтей, на четырех рядах кедровых столбов; и кедровые бревна [положены были] на столбах.
1KGS|7|3|И настлан был помост из кедра над бревнами на сорока пяти столбах, по пятнадцати в ряд.
1KGS|7|4|Оконных косяков [было] три ряда; и три ряда [окон], окно против окна.
1KGS|7|5|И все двери и дверные косяки были четырехугольные, и окно против окна, в три ряда.
1KGS|7|6|И притвор из столбов сделал он длиною в пятьдесят локтей, шириною в тридцать локтей, и пред ними крыльцо, и столбы, и порог пред ними.
1KGS|7|7|Еще притвор с престолом, с которого он судил, притвор для судилища сделал он и покрыл все полы кедром.
1KGS|7|8|В доме, где он жил, другой двор позади притвора был такого же устройства. И в доме дочери фараоновой, которую взял за себя Соломон, он сделал такой же притвор.
1KGS|7|9|Все это сделано было из дорогих камней, обтесанных по размеру, обрезанных пилою, с внутренней и наружной стороны, от основания до выступов, и с наружной стороны до большого двора.
1KGS|7|10|И в основание положены были камни дорогие, камни большие, камни в десять локтей и камни в восемь локтей,
1KGS|7|11|и сверху дорогие камни, обтесанные по размеру, и кедр.
1KGS|7|12|Большой двор огорожен был кругом тремя рядами тесаных камней и одним рядом кедровых бревен; также и внутренний двор храма Господа и притвор храма.
1KGS|7|13|И послал царь Соломон и взял из Тира Хирама,
1KGS|7|14|сына одной вдовы, из колена Неффалимова. Отец его Тирянин был медник; он владел способностью, искусством и уменьем выделывать всякие вещи из меди. И пришел он к царю Соломону и производил у него всякие работы:
1KGS|7|15|и сделал он два медных столба, каждый в восемнадцать локтей вышиною, и снурок в двенадцать локтей обнимал [окружность] того и другого столба;
1KGS|7|16|и два венца, вылитых из меди, он сделал, чтобы положить на верху столбов: пять локтей вышины в одном венце и пять локтей вышины в другом венце;
1KGS|7|17|сетки плетеной работы и снурки в виде цепочек для венцов, которые были на верху столбов: семь на одном венце и семь на другом венце.
1KGS|7|18|Так сделал он столбы и два ряда гранатовых яблок вокруг сетки, чтобы покрыть венцы, которые на верху столбов; то же сделал и для другого венца.
1KGS|7|19|А в притворе венцы на верху столбов сделаны [на подобие лилии], в четыре локтя,
1KGS|7|20|и венцы на обоих столбах вверху, прямо над выпуклостью, которая подле сетки; и на другом венце, рядами кругом, двести гранатовых яблок.
1KGS|7|21|И поставил столбы к притвору храма; поставил столб направой стороне и дал ему имя Иахин, и поставил столб на левой стороне и дал ему имя Воаз.
1KGS|7|22|И над столбами поставил [венцы], сделанные [наподобие] лилии; так окончена работа над столбами.
1KGS|7|23|И сделал литое [из меди] море, – от края его до края его десять локтей, – совсем круглое, вышиною в пять локтей, и снурок в тридцать локтей обнимал его кругом.
1KGS|7|24|[Подобия] огурцов под краями его окружали его по десяти на локоть, окружали море со всех сторон в два ряда; [подобия] огурцов были вылиты с ним одним литьем.
1KGS|7|25|Оно стояло на двенадцати волах: три глядели к северу, три глядели к западу, три глядели к югу и три глядели к востоку; море лежало на них, и зады их [обращены были] внутрь под него.
1KGS|7|26|Толщиною оно было в ладонь, и края его, сделанные подобно краям чаши, [походили] на распустившуюся лилию. Оно вмещало две тысячи батов.
1KGS|7|27|И сделал он десять медных подстав; длина каждой подставы – четыре локтя, ширина – четыре локтя и три локтя – вышина.
1KGS|7|28|И вот устройство подстав: у них стенки, стенки между наугольными пластинками;
1KGS|7|29|на стенках, которые между наугольниками, [изображены] были львы, волы и херувимы; также и на наугольниках, а выше и ниже львов и волов – развесистые венки;
1KGS|7|30|у каждой подставы по четыре медных колеса и оси медные. На четырех углах выступы на подобие плеч, выступы литые внизу, под чашею, подле каждого венка.
1KGS|7|31|Отверстие от внутреннего венка до верха в один локоть; отверстие его круглое, подобно подножию столбов, в полтора локтя, и при отверстии его изваяния; но боковые стенки четырехугольные, не круглые.
1KGS|7|32|Под стенками было четыре колеса, и оси колес в подставах; вышина каждого колеса – полтора локтя.
1KGS|7|33|Устройство колес такое же, как устройство колес в колеснице; оси их, и ободья их, и спицы их, и ступицы их, все было литое.
1KGS|7|34|Четыре выступа на четырех углах каждой подставы; из подставы [выходили] выступы ее.
1KGS|7|35|И на верху подставы круглое возвышение на поллоктя вышины; и на верху подставы рукоятки ее и стенки ее из одной с нею массы.
1KGS|7|36|И изваял он на дощечках ее рукоятки и на стенках ее херувимов, львов и пальмы, сколько где позволяло место, и вокруг развесистые венки.
1KGS|7|37|Так сделал он десять подстав: у всех их одно литье, одна мера, один вид.
1KGS|7|38|И сделал десять медных умывальниц: каждая умывальница вмещала сорок батов, каждая умывальница была в четыре локтя, каждая умывальница стояла на одной из десяти подстав.
1KGS|7|39|И расставил подставы – пять на правой стороне храма и пять на левой стороне храма, а море поставил на правой стороне храма, на восточно–южной стороне.
1KGS|7|40|И сделал Хирам умывальницы и лопатки и чаши. И кончил Хирам всю работу, которую производил у царя Соломона для храма Господня:
1KGS|7|41|два столба и две опояски венцов, которые на верху столбов, и две сетки для покрытия двух опоясок венцов, которые на верху столбов;
1KGS|7|42|и четыреста гранатовых яблок на двух сетках; два ряда гранатовых яблок для каждой сетки, для покрытия двух опоясок венцов, которые на столбах;
1KGS|7|43|и десять подстав и десять умывальниц на подставах;
1KGS|7|44|одно море и двенадцать волов под морем;
1KGS|7|45|и тазы, и лопатки, и чаши. Все вещи, которые сделал Хирам царю Соломону для храма Господа, [были] из полированной меди.
1KGS|7|46|Царь выливал их в глинистой земле, в окрестности Иордана, между Сокхофом и Цартаном.
1KGS|7|47|И поставил Соломон все сии вещи [на место]. По причине чрезвычайного их множества, вес меди не определен.
1KGS|7|48|И сделал Соломон все вещи, которые в храме Господа: золотой жертвенник и золотой стол, на котором хлебы предложения;
1KGS|7|49|и светильники – пять по правую сторону и пять по левую сторону, пред задним отделением храма, из чистого золота, и цветы, и лампадки, и щипцы из золота;
1KGS|7|50|и блюда, и ножи, и чаши, и лотки, и кадильницы из чистого золота, и петли у дверей внутреннего храма во Святом Святых и у дверей в храме из золота же.
1KGS|7|51|Так совершена вся работа, которую производил царь Соломон для храма Господа. И принес Соломон посвященное Давидом, отцом его; серебро и золото и вещи отдал в сокровищницы храма Господня.
1KGS|8|1|Тогда созвал Соломон старейшин Израилевых и всех начальников колен, глав поколений сынов Израилевых, к царю Соломону в Иерусалим, чтобы перенести ковчег завета Господня из города Давидова, то есть Сиона.
1KGS|8|2|И собрались к царю Соломону на праздник все Израильтяне в месяце Афаниме, который есть седьмой месяц.
1KGS|8|3|И пришли все старейшины Израилевы; и подняли священники ковчег,
1KGS|8|4|и понесли ковчег Господень и скинию собрания и все священные вещи, которые были в скинии; и несли их священники и левиты.
1KGS|8|5|А царь Соломон и с ним все общество Израилево, собравшееся к нему, шли пред ковчегом, принося жертвы из мелкого и крупного скота, которых невозможно исчислить и определить, по множеству их.
1KGS|8|6|И внесли священники ковчег завета Господня на место его, в давир храма, во Святое Святых, под крылья херувимов.
1KGS|8|7|Ибо херувимы простирали крылья над местом ковчега, и покрывали херувимы сверху ковчег и шесты его.
1KGS|8|8|И выдвинулись шесты так, что головки шестов видны были из святилища пред давиром, но не выказывались наружу; они там и до сего дня.
1KGS|8|9|В ковчеге ничего не было, кроме двух каменных скрижалей, которые положил туда Моисей на Хориве, когда Господь заключил завет с сынами Израилевыми, по исшествии их из земли Египетской.
1KGS|8|10|Когда священники вышли из святилища, облако наполнило дом Господень;
1KGS|8|11|и не могли священники стоять на служении, по причине облака, ибо слава Господня наполнила храм Господень.
1KGS|8|12|Тогда сказал Соломон: Господь сказал, что Он благоволит обитать во мгле;
1KGS|8|13|я построил храм в жилище Тебе, место, чтобы пребывать Тебе во веки.
1KGS|8|14|И обратился царь лицем своим, и благословил все собрание Израильтян; все собрание Израильтян стояло, –
1KGS|8|15|и сказал: благословен Господь Бог Израилев, Который сказал Своими устами Давиду, отцу моему, и ныне исполнил рукою Своею! Он говорил:
1KGS|8|16|"с того дня, как Я вывел народ Мой Израиля из Египта, Я не избрал города ни в одном из колен Израилевых, чтобы построен был дом, в котором пребывало бы имя Мое; и избрал Давида, чтобы быть ему над народом Моим Израилем".
1KGS|8|17|У Давида, отца моего, было на сердце построить храм имени Господа Бога Израилева;
1KGS|8|18|но Господь сказал Давиду, отцу моему: "у тебя есть на сердце построить храм имени Моему; хорошо, что это у тебя лежит на сердце;
1KGS|8|19|однако не ты построишь храм, а сын твой, исшедший из чресл твоих, он построит храм имени Моему".
1KGS|8|20|И исполнил Господь слово Свое, которое изрек. Я вступил на место отца моего Давида и сел на престоле Израилевом, как сказал Господь, и построил храм имени Господа Бога Израилева;
1KGS|8|21|и приготовил там место для ковчега, в котором завет Господа, заключенный Им с отцами нашими, когда Он вывел их из земли Египетской.
1KGS|8|22|И стал Соломон пред жертвенником Господним впереди всего собрания Израильтян, и воздвиг руки свои к небу,
1KGS|8|23|и сказал: Господи Боже Израилев! нет подобного Тебе Бога на небесах вверху и на земле внизу; Ты хранишь завет и милость к рабам Твоим, ходящим пред Тобою всем сердцем своим.
1KGS|8|24|Ты исполнил рабу Твоему Давиду, отцу моему, что говорил ему; что изрек Ты устами Твоими, то в сей день совершил рукою Твоею.
1KGS|8|25|И ныне, Господи Боже Израилев, исполни рабу Твоему Давиду, отцу моему, то, что говорил Ты ему, сказав: "не прекратится у тебя пред лицем Моим сидящий на престоле Израилевом, если только сыновья твои будут держаться пути своего, ходя предо Мною так, как ты ходил предо Мною".
1KGS|8|26|И ныне, Боже Израилев, да будет верно слово Твое, которое Ты изрек рабу Твоему Давиду, отцу моему!
1KGS|8|27|Поистине, Богу ли жить на земле? Небо и небо небес не вмещают Тебя, тем менее сей храм, который я построил.
1KGS|8|28|но призри на молитву раба Твоего и на прошение его, Господи Боже мой; услышь воззвание и молитву, которою раб Твой умоляет Тебя ныне.
1KGS|8|29|Да будут очи Твои отверсты на храм сей день и ночь, на сие место, о котором Ты сказал: "Мое имя будет там"; услышь молитву, которою будет молиться раб Твой на месте сем.
1KGS|8|30|Услышь моление раба Твоего и народа Твоего Израиля, когда они будут молиться на месте сем; услышь на месте обитания Твоего, на небесах, услышь и помилуй.
1KGS|8|31|Когда кто согрешит против ближнего своего, и потребует от него клятвы, чтобы он поклялся, и для клятвы придут пред жертвенник Твой в храм сей,
1KGS|8|32|тогда Ты услышь с неба и произведи суд над рабами Твоими, обвини виновного, возложив поступок его на голову его, и оправдай правого, воздав ему по правде его.
1KGS|8|33|Когда народ Твой Израиль будет поражен неприятелем за то, что согрешил пред Тобою, и когда они обратятся к Тебе, и исповедают имя Твое, и будут просить и умолять Тебя в сем храме,
1KGS|8|34|тогда Ты услышь с неба и прости грех народа Твоего Израиля, и возврати их в землю, которую Ты дал отцам их.
1KGS|8|35|Когда заключится небо и не будет дождя за то, что они согрешат пред Тобою, и когда помолятся на месте сем и исповедают имя Твое и обратятся от греха своего, ибо Ты смирил их,
1KGS|8|36|тогда услышь с неба и прости грех рабов Твоих и народа Твоего Израиля, указав им добрый путь, по которому идти, и пошли дождь на землю Твою, которую Ты дал народу Твоему в наследие.
1KGS|8|37|Будет ли на земле голод, будет ли моровая язва, будет ли палящий ветер, ржавчина, саранча, червь, неприятель ли будет теснить его в земле его, [будет ли] какое бедствие, какая болезнь, –
1KGS|8|38|при всякой молитве, при всяком прошении, какое будет от какого–либо человека во всем народе Твоем Израиле, когда они почувствуют бедствие в сердце своем и прострут руки свои к храму сему,
1KGS|8|39|Ты услышь с неба, с места обитания Твоего, и помилуй; соделай и воздай каждому по путям его, как Ты усмотришь сердце его, ибо Ты один знаешь сердце всех сынов человеческих:
1KGS|8|40|чтобы они боялись Тебя во все дни, доколе живут на земле, которую Ты дал отцам нашим.
1KGS|8|41|Если и иноплеменник, который не от Твоего народа Израиля, придет из земли далекой ради имени Твоего, –
1KGS|8|42|ибо и они услышат о Твоем имени великом и о Твоей руке сильной и о Твоей мышце простертой, – и придет он и помолится у храма сего,
1KGS|8|43|услышь с неба, с места обитания Твоего, и сделай все, о чем будет взывать к Тебе иноплеменник, чтобы все народы земли знали имя Твое, чтобы боялись Тебя, как народ Твой Израиль, чтобы знали, что именем Твоим называется храм сей, который я построил.
1KGS|8|44|Когда выйдет народ Твой на войну против врага своего путем, которым Ты пошлешь его, и будет молиться Господу, обратившись к городу, который Ты избрал, и к храму, который я построил имени Твоему,
1KGS|8|45|тогда услышь с неба молитву их и прошение их и сделай, что потребно для них.
1KGS|8|46|Когда они согрешат пред Тобою, – ибо нет человека, который не грешил бы, – и Ты прогневаешься на них и предашь их врагам, и пленившие их отведут их в неприятельскую землю, далекую или близкую;
1KGS|8|47|и когда они в земле, в которой будут находиться в плену, войдут в себя и обратятся и будут молиться Тебе в земле пленивших их, говоря: "мы согрешили, сделали беззаконие, мы виновны";
1KGS|8|48|и когда обратятся к Тебе всем сердцем своим и всею душею своею в земле врагов, которые пленили их, и будут молиться Тебе, обратившись к земле своей, которую Ты дал отцам их, к городу, который Ты избрал, и к храму, который я построил имени Твоему,
1KGS|8|49|тогда услышь с неба, с места обитания Твоего, молитву и прошение их и сделай, что потребно для них;
1KGS|8|50|и прости народу Твоему, в чем он согрешил пред Тобою, и все проступки его, которые он сделал пред Тобою, и возбуди сострадание к ним в пленивших их, чтобы они были милостивы к ним:
1KGS|8|51|ибо они Твой народ и Твой удел, который Ты вывел из Египта, из железной печи.
1KGS|8|52|Да будут очи Твои отверсты на молитву раба Твоего и на молитву народа Твоего Израиля, чтобы слышать их всегда, когда они будут призывать Тебя,
1KGS|8|53|ибо Ты отделил их Себе в удел из всех народов земли, как Ты изрек чрез Моисея, раба Твоего, когда вывел отцов наших из Египта, Владыка Господи!
1KGS|8|54|Когда Соломон произнес все сие моление и прошение к Господу, тогда встал с колен от жертвенника Господня, [руки же] его были распростерты к небу.
1KGS|8|55|И стоя благословил все собрание Израильтян, громким голосом говоря:
1KGS|8|56|благословен Господь, Который дал покой народу Своему Израилю, как говорил! не осталось неисполненным ни одного слова из всех благих слов Его, которые Он изрек чрез раба Своего Моисея;
1KGS|8|57|да будет с нами Господь Бог наш, как был Он с отцами нашими, да не оставит нас, да не покинет нас,
1KGS|8|58|наклоняя к Себе сердце наше, чтобы мы ходили по всем путям Его и соблюдали заповеди Его и уставы Его и законы Его, которые Он заповедал отцам нашим;
1KGS|8|59|и да будут слова сии, которыми я молился пред Господом, близки к Господу Богу нашему день и ночь, дабы Он делал, что потребно для раба Своего, и что потребно для народа Своего Израиля, изо дня в день,
1KGS|8|60|чтобы все народы познали, что Господь есть Бог и нет кроме Его;
1KGS|8|61|да будет сердце ваше вполне предано Господу Богу нашему, чтобы ходить по уставам Его и соблюдать заповеди Его, как ныне.
1KGS|8|62|И царь и все Израильтяне с ним принесли жертву Господу.
1KGS|8|63|И принес Соломон в мирную жертву, которую принес он Господу, двадцать две тысячи крупного скота и сто двадцать тысяч мелкого скота. Так освятили храм Господу царь и все сыны Израилевы.
1KGS|8|64|В тот же день освятил царь среднюю часть двора, который пред храмом Господним, совершив там всесожжение и хлебное приношение и [вознеся] тук мирных жертв, потому что медный жертвенник, который пред Господом, был мал для помещения всесожжения и хлебного приношения и тука мирных жертв.
1KGS|8|65|И сделал Соломон в это время праздник, и весь Израиль с ним, – большое собрание, [сошедшееся] от входа в Емаф до реки Египетской пред Господом Богом нашим; – семь дней и еще семь дней, четырнадцать дней.
1KGS|8|66|В восьмой день Соломон отпустил народ. И благословили царя и пошли в шатры свои, радуясь и веселясь в сердце о всем добром, что сделал Господь рабу Своему Давиду и народу Своему Израилю.
1KGS|9|1|После того, как Соломон кончил строение храма Господня и дома царского и все, что Соломон желал сделать,
1KGS|9|2|явился Соломону Господь во второй раз, как явился ему в Гаваоне.
1KGS|9|3|И сказал ему Господь: Я услышал молитву твою и прошение твое, о чем ты просил Меня. Я освятил сей храм, который ты построил, чтобы пребывать имени Моему там вовек; и будут очи Мои и сердце Мое там во все дни.
1KGS|9|4|И если ты будешь ходить пред лицем Моим, как ходил отец твой Давид, в чистоте сердца и в правоте, исполняя все, что Я заповедал тебе, и если будешь хранить уставы Мои и законы Мои,
1KGS|9|5|то Я поставлю царский престол твой над Израилем вовек, как Я сказал отцу твоему Давиду, говоря: "не прекратится у тебя сидящий на престоле Израилевом".
1KGS|9|6|Если же вы и сыновья ваши отступите от Меня и не будете соблюдать заповедей Моих и уставов Моих, которые Я дал вам, и пойдете и станете служить иным богам и поклоняться им,
1KGS|9|7|то Я истреблю Израиля с лица земли, которую Я дал ему, и храм, который Я освятил имени Моему, отвергну от лица Моего, и будет Израиль притчею и посмешищем у всех народов.
1KGS|9|8|И о храме сем высоком всякий, проходящий мимо его, ужаснется и свистнет, и скажет: "за что Господь поступил так с сею землею и с сим храмом?"
1KGS|9|9|И скажут: "за то, что они оставили Господа Бога своего, Который вывел отцов их из земли Египетской, и приняли других богов, и поклонялись им и служили им, – за это навел на них Господь все сие бедствие".
1KGS|9|10|По окончании двадцати лет, в которые Соломон построил два дома, – дом Господень и дом царский, –
1KGS|9|11|на что Хирам, царь Тирский, доставлял Соломону дерева кедровые и дерева кипарисовые и золото, по его желанию, – царь Соломон дал Хираму двадцать городов в земле Галилейской.
1KGS|9|12|И вышел Хирам из Тира посмотреть города, которые дал ему Соломон, и они не понравились ему.
1KGS|9|13|И сказал он: что это за города, которые ты, брат мой, дал мне? И назвал их землею Кавул, [как называются они] до сего дня.
1KGS|9|14|И послал Хирам царю сто двадцать талантов золота.
1KGS|9|15|Вот распоряжение о подати, которую наложил царь Соломон, чтобы построить храм Господень и дом свой, и Милло, и стену Иерусалимскую, Гацор, и Мегиддо, и Газер.
1KGS|9|16|Фараон, царь Египетский, пришел и взял Газер, и сжег его огнем, и Хананеев, живших в городе, побил, и отдал его в приданое дочери своей, жене Соломоновой.
1KGS|9|17|И построил Соломон Газер и нижний Бефорон,
1KGS|9|18|и Ваалаф и Фадмор в пустыне,
1KGS|9|19|и все города для запасов, которые были у Соломона, и города для колесниц, и города для конницы и все то, что Соломон хотел построить в Иерусалиме и на Ливане и во всей земле своего владения.
1KGS|9|20|Весь народ, оставшийся от Аморреев, Хеттеев, Ферезеев, Евеев, и Иевусеев, которые были не из сынов Израилевых,
1KGS|9|21|детей их, оставшихся после них на земле, которых сыны Израилевы не могли истребить, Соломон сделал оброчными работниками до сего дня.
1KGS|9|22|Сынов же Израилевых Соломон не делал работниками, но они были его воинами, его слугами, его вельможами, его военачальниками и вождями его колесниц и его всадников.
1KGS|9|23|Вот главные приставники над работами Соломоновыми: управлявших народом, который производил работы, было пятьсот пятьдесят.
1KGS|9|24|Дочь фараонова перешла из города Давидова в свой дом, который построил для нее Соломон; потом построил он Милло.
1KGS|9|25|И приносил Соломон три раза в год всесожжения и мирные жертвы на жертвеннике, который он построил Господу, и курение на нем совершал пред Господом. И окончил он [строение] дома.
1KGS|9|26|Царь Соломон также сделал корабль в Ецион–Гавере, что при Елафе, на берегу Чермного моря, в земле Идумейской.
1KGS|9|27|И послал Хирам на корабле своих подданных корабельщиков, знающих море, с подданными Соломоновыми;
1KGS|9|28|и отправились они в Офир, и взяли оттуда золота четыреста двадцать талантов, и привезли царю Соломону.
1KGS|10|1|Царица Савская, услышав о славе Соломона во имя Господа, пришла испытать его загадками.
1KGS|10|2|И пришла она в Иерусалим с весьма большим богатством: верблюды навьючены [были] благовониями и великим множеством золота и драгоценными камнями; и пришла к Соломону и беседовала с ним обо всем, что было у нее на сердце.
1KGS|10|3|И объяснил ей Соломон все слова ее, и не было ничего незнакомого царю, чего бы он не изъяснил ей.
1KGS|10|4|И увидела царица Савская всю мудрость Соломона и дом, который он построил,
1KGS|10|5|и пищу за столом его, и жилище рабов его, и стройность слуг его, и одежду их, и виночерпиев его, и всесожжения его, которые он приносил в храме Господнем. И не могла она более удержаться
1KGS|10|6|и сказала царю: верно то, что я слышала в земле своей о делах твоих и о мудрости твоей;
1KGS|10|7|но я не верила словам, доколе не пришла, и не увидели глаза мои: и вот, мне и в половину не сказано; мудрости и богатства у тебя больше, нежели как я слышала.
1KGS|10|8|Блаженны люди твои и блаженны сии слуги твои, которые всегда предстоят пред тобою и слышат мудрость твою!
1KGS|10|9|Да будет благословен Господь Бог твой, Который благоволил посадить тебя на престол Израилев! Господь, по вечной любви Своей к Израилю, поставил тебя царем, творить суд и правду.
1KGS|10|10|И подарила она царю сто двадцать талантов золота и великое множество благовоний и драгоценные камни; никогда еще не приходило такого множества благовоний, какое подарила царица Савская царю Соломону.
1KGS|10|11|И корабль Хирамов, который привозил золото из Офира, привез из Офира великое множество красного дерева и драгоценных камней.
1KGS|10|12|И сделал царь из сего красного дерева перила для храма Господня и для дома царского, и гусли и псалтири для певцов; никогда не приходило столько красного дерева и не видано было до сего дня.
1KGS|10|13|И царь Соломон дал царице Савской все, чего она желала и чего просила, сверх того, что подарил ей царь Соломон своими руками. И отправилась она обратно в свою землю, она и все слуги ее.
1KGS|10|14|В золоте, которое приходило Соломону в каждый год, весу было шестьсот шестьдесят шесть талантов золотых,
1KGS|10|15|сверх того, что [получаемо было] от разносчиков товара и от торговли купцов, и от всех царей Аравийских и от областных начальников.
1KGS|10|16|И сделал царь Соломон двести больших щитов из кованого золота, по шестисот [сиклей] пошло на каждый щит;
1KGS|10|17|и триста меньших щитов из кованого золота, по три мины золота пошло на каждый щит; и поставил их царь в доме из Ливанского дерева.
1KGS|10|18|И сделал царь большой престол из слоновой кости и обложил его чистым золотом;
1KGS|10|19|к престолу было шесть ступеней; верх сзади у престола был круглый, и были с обеих сторон у места сиденья локотники, и два льва стояли у локотников;
1KGS|10|20|и еще двенадцать львов стояли там на шести ступенях по обе стороны. Подобного сему не бывало ни в одном царстве.
1KGS|10|21|И все сосуды для питья у царя Соломона [были] золотые, и все сосуды в доме из Ливанского дерева были из чистого золота; из серебра ничего не было, потому что серебро во дни Соломоновы считалось ни за что;
1KGS|10|22|ибо у царя был на море Фарсисский корабль с кораблем Хирамовым; в три года раз приходил Фарсисский корабль, привозивший золото и серебро, и слоновую кость, и обезьян, и павлинов.
1KGS|10|23|Царь Соломон превосходил всех царей земли богатством и мудростью.
1KGS|10|24|И все [цари] на земле искали видеть Соломона, чтобы послушать мудрости его, которую вложил Бог в сердце его.
1KGS|10|25|И они подносили ему, каждый от себя, в дар: сосуды серебряные и сосуды золотые, и одежды, и оружие, и благовония, коней и мулов, каждый год.
1KGS|10|26|И набрал Соломон колесниц и всадников; у него было тысяча четыреста колесниц и двенадцать тысяч всадников; и разместил он их по колесничным городам и при царе в Иерусалиме.
1KGS|10|27|И сделал царь серебро в Иерусалиме равноценным с простыми камнями, а кедры, по их множеству, сделал равноценными с сикоморами, [растущими] на низких местах.
1KGS|10|28|Коней же царю Соломону приводили из Египта и из Кувы; царские купцы покупали их из Кувы за деньги.
1KGS|10|29|Колесница из Египта получаема и доставляема была за шестьсот [сиклей] серебра, а конь за сто пятьдесят. Таким же образом они руками своими доставляли [все это] царям Хеттейским и царям Арамейским.
1KGS|11|1|И полюбил царь Соломон многих чужестранных женщин, кроме дочери фараоновой, Моавитянок, Аммонитянок, Идумеянок, Сидонянок, Хеттеянок,
1KGS|11|2|из тех народов, о которых Господь сказал сынам Израилевым: "не входите к ним, и они пусть не входят к вам, чтобы они не склонили сердца вашего к своим богам"; к ним прилепился Соломон любовью.
1KGS|11|3|И было у него семьсот жен и триста наложниц; и развратили жены его сердце его.
1KGS|11|4|Во время старости Соломона жены его склонили сердце его к иным богам, и сердце его не было вполне предано Господу Богу своему, как сердце Давида, отца его.
1KGS|11|5|И стал Соломон служить Астарте, божеству Сидонскому, и Милхому, мерзости Аммонитской.
1KGS|11|6|И делал Соломон неугодное пред очами Господа и не вполне последовал Господу, как Давид, отец его.
1KGS|11|7|Тогда построил Соломон капище Хамосу, мерзости Моавитской, на горе, которая пред Иерусалимом, и Молоху, мерзости Аммонитской.
1KGS|11|8|Так сделал он для всех своих чужестранных жен, которые кадили и приносили жертвы своим богам.
1KGS|11|9|И разгневался Господь на Соломона за то, что он уклонил сердце свое от Господа Бога Израилева, Который два раза являлся ему
1KGS|11|10|и заповедал ему, чтобы он не следовал иным богам; но он не исполнил того, что заповедал ему Господь.
1KGS|11|11|И сказал Господь Соломону: за то, что так у тебя делается, и ты не сохранил завета Моего и уставов Моих, которые Я заповедал тебе, Я отторгну от тебя царство и отдам его рабу твоему;
1KGS|11|12|но во дни твои Я не сделаю сего ради Давида, отца твоего; из руки сына твоего исторгну его;
1KGS|11|13|и не все царство исторгну; одно колено дам сыну твоему ради Давида, раба Моего, и ради Иерусалима, который Я избрал.
1KGS|11|14|И воздвиг Господь противника на Соломона, Адера Идумеянина, из царского Идумейского рода.
1KGS|11|15|Когда Давид был в Идумее, и военачальник Иоав пришел для погребения убитых и избил весь мужеский пол в Идумее, –
1KGS|11|16|ибо шесть месяцев прожил там Иоав и все Израильтяне, доколе не истребили всего мужеского пола в Идумее, –
1KGS|11|17|тогда сей Адер убежал в Египет и с ним несколько Идумеян, служивших при отце его; Адер [был тогда] малым ребенком.
1KGS|11|18|Отправившись из Мадиама, они пришли в Фаран и взяли с собою людей из Фарана и пришли в Египет к фараону, царю Египетскому. он дал ему дом, и назначил ему содержание, и дал ему землю.
1KGS|11|19|Адер снискал у фараона большую милость, так что он дал ему в жену сестру своей жены, сестру царицы Тахпенесы.
1KGS|11|20|И родила ему сестра Тахпенесы сына Генувата. Тахпенеса воспитывала его в доме фараоновом; и жил Генуват в доме фараоновом вместе с сыновьями фараоновыми.
1KGS|11|21|Когда Адер услышал, что Давид почил с отцами своими и что военачальник Иоав умер, то сказал фараону: отпусти меня, я пойду в свою землю.
1KGS|11|22|И сказал ему фараон: разве ты нуждаешься в чем у меня, что хочешь идти в свою землю? Он отвечал: нет, но отпусти меня.
1KGS|11|23|И воздвиг Бог против Соломона еще противника, Разона, сына Елиады, который убежал от государя своего Адраазара, царя Сувского,
1KGS|11|24|и, собрав около себя людей, сделался начальником шайки, после того, как Давид разбил [Адраазара]; и пошли они в Дамаск, и водворились там, и владычествовали в Дамаске.
1KGS|11|25|И был он противником Израиля во все дни Соломона. Кроме зла, [причиненного] Адером, он всегда вредил Израилю и сделался царем Сирии.
1KGS|11|26|И Иеровоам, сын Наватов, Ефремлянин из Цареды, – имя матери его вдовы: Церуа, – раб Соломонов, поднял руку на царя.
1KGS|11|27|И вот обстоятельство, по которому он поднял руку на царя: Соломон строил Милло, починивал повреждения в городе Давида, отца своего.
1KGS|11|28|Иеровоам был человек мужественный. Соломон, заметив, что этот молодой человек умеет делать дело, поставил его смотрителем над оброчными из дома Иосифова.
1KGS|11|29|В то время случилось Иеровоаму выйти из Иерусалима; и встретил его на дороге пророк Ахия Силомлянин, и на нем была новая одежда. На поле их было только двое.
1KGS|11|30|И взял Ахия новую одежду, которая была на нем, и разодрал ее на двенадцать частей,
1KGS|11|31|и сказал Иеровоаму: возьми себе десять частей, ибо так говорит Господь Бог Израилев: вот, Я исторгаю царство из руки Соломоновой и даю тебе десять колен,
1KGS|11|32|а одно колено останется за ним ради раба Моего Давида и ради города Иерусалима, который Я избрал из всех колен Израилевых.
1KGS|11|33|Это за то, что они оставили Меня и стали поклоняться Астарте, божеству Сидонскому, и Хамосу, богу Моавитскому, и Милхому, богу Аммонитскому, и не пошли путями Моими, чтобы делать угодное пред очами Моими и [соблюдать] уставы Мои и заповеди Мои, подобно Давиду, отцу его.
1KGS|11|34|Я не беру всего царства из руки его, но Я оставлю его владыкою на все дни жизни его ради Давида, раба Моего, которого Я избрал, который соблюдал заповеди Мои и уставы Мои;
1KGS|11|35|но возьму царство из руки сына его и дам тебе из него десять колен;
1KGS|11|36|а сыну его дам одно колено, дабы оставался светильник Давида, раба Моего, во все дни пред лицем Моим, в городе Иерусалиме, который Я избрал Себе для пребывания там имени Моего.
1KGS|11|37|Тебя Я избираю, и ты будешь владычествовать над всем, чего пожелает душа твоя, и будешь царем над Израилем;
1KGS|11|38|и если будешь соблюдать все, что Я заповедую тебе, и будешь ходить путями Моими и делать угодное пред очами Моими, соблюдая уставы Мои и заповеди Мои, как делал раб Мой Давид, то Я буду с тобою и устрою тебе дом твердый, как Я устроил Давиду, и отдам тебе Израиля;
1KGS|11|39|и смирю Я род Давидов за сие, но не на все дни.
1KGS|11|40|Соломон же хотел умертвить Иеровоама; но Иеровоам встал и убежал в Египет к Сусакиму, царю Египетскому, и жил в Египте до смерти Соломоновой.
1KGS|11|41|Прочие события Соломоновы и все, что он делал, и мудрость его описаны в книге дел Соломоновых.
1KGS|11|42|Времени царствования Соломонова в Иерусалиме над всем Израилем [было] сорок лет.
1KGS|11|43|И почил Соломон с отцами своими и погребен был в городе Давида, отца своего, и воцарился вместо него сын его Ровоам.
1KGS|12|1|И пошел Ровоам в Сихем, ибо в Сихем пришли все Израильтяне, чтобы воцарить его.
1KGS|12|2|И услышал о том Иеровоам, сын Наватов, когда находился еще в Египте, куда убежал от царя Соломона, и возвратился Иеровоам из Египта;
1KGS|12|3|и послали за ним и призвали его. Тогда Иеровоам и все собрание Израильтян пришли и говорили Ровоаму и сказали:
1KGS|12|4|отец твой наложил на нас тяжкое иго, ты же облегчи нам жестокую работу отца твоего и тяжкое иго, которое он наложил на нас, и тогда мы будем служить тебе.
1KGS|12|5|И сказал он им: пойдите и чрез три дня опять придите ко мне. И пошел народ.
1KGS|12|6|Царь Ровоам советовался со старцами, которые предстояли пред Соломоном, отцом его, при жизни его, и говорил: как посоветуете вы мне отвечать сему народу?
1KGS|12|7|Они говорили ему и сказали: если ты на сей день будешь слугою народу сему и услужишь ему, и удовлетворишь им и будешь говорить им ласково, то они будут твоими рабами на все дни.
1KGS|12|8|Но он пренебрег совет старцев, что они советовали ему, и советовался с молодыми людьми, которые выросли вместе с ним и которые предстояли пред ним,
1KGS|12|9|и сказал им: что вы посоветуете мне отвечать народу сему, который говорил мне и сказал: "облегчи иго, которое наложил на нас отец твой"?
1KGS|12|10|И говорили ему молодые люди, которые выросли вместе с ним, и сказали: так скажи народу сему, который говорил тебе и сказал: "отец твой наложил на нас тяжкое иго, ты же облегчи нас"; так скажи им: "мой мизинец толще чресл отца моего;
1KGS|12|11|итак, если отец мой обременял вас тяжким игом, то я увеличу иго ваше; отец мой наказывал вас бичами, а я буду наказывать вас скорпионами".
1KGS|12|12|Иеровоам и весь народ пришли к Ровоаму на третий день, как приказал царь, сказав: придите ко мне на третий день.
1KGS|12|13|И отвечал царь народу сурово и пренебрег совет старцев, что они советовали ему;
1KGS|12|14|и говорил он по совету молодых людей и сказал: отец мой наложил на вас тяжкое иго, а я увеличу иго ваше; отец мой наказывал вас бичами, а я буду наказывать вас скорпионами.
1KGS|12|15|И не послушал царь народа, ибо так суждено было Господом, чтобы исполнилось слово Его, которое изрек Господь чрез Ахию Силомлянина Иеровоаму, сыну Наватову.
1KGS|12|16|И увидели все Израильтяне, что царь не послушал их. И отвечал народ царю и сказал: какая нам часть в Давиде? нет нам доли в сыне Иессеевом; по шатрам своим, Израиль! теперь знай свой дом, Давид! И разошелся Израиль по шатрам своим.
1KGS|12|17|Только над сынами Израилевыми, жившими в городах Иудиных, царствовал Ровоам.
1KGS|12|18|И послал царь Ровоам Адонирама, начальника над податью; но все Израильтяне забросали его каменьями, и он умер; царь же Ровоам поспешно взошел на колесницу, чтоб убежать в Иерусалим.
1KGS|12|19|И отложился Израиль от дома Давидова до сего дня.
1KGS|12|20|Когда услышали все Израильтяне, что Иеровоам возвратился, то послали и призвали его в собрание, и воцарили его над всеми Израильтянами. За домом Давидовым не осталось никого, кроме колена Иудина [и Вениаминова].
1KGS|12|21|Ровоам, прибыв в Иерусалим, собрал из всего дома Иудина и из колена Вениаминова сто восемьдесят тысяч отборных воинов, дабы воевать с домом Израилевым для того, чтобы возвратить царство Ровоаму, сыну Соломонову.
1KGS|12|22|И было слово Божие к Самею, человеку Божию, и сказано:
1KGS|12|23|скажи Ровоаму, сыну Соломонову, царю Иудейскому, и всему дому Иудину и Вениаминову и прочему народу:
1KGS|12|24|так говорит Господь: не ходите и не начинайте войны с братьями вашими, сынами Израилевыми; возвратитесь каждый в дом свой, ибо от Меня это было. И послушались они слова Господня и пошли назад по слову Господню.
1KGS|12|25|И обстроил Иеровоам Сихем на горе Ефремовой и поселился в нем; оттуда пошел и построил Пенуил.
1KGS|12|26|И говорил Иеровоам в сердце своем: царство может опять перейти к дому Давидову;
1KGS|12|27|если народ сей будет ходить в Иерусалим для жертвоприношения в доме Господнем, то сердце народа сего обратится к государю своему, к Ровоаму, царю Иудейскому, и убьют они меня и возвратятся к Ровоаму, царю Иудейскому.
1KGS|12|28|И посоветовавшись царь сделал двух золотых тельцов и сказал [народу]: не нужно вам ходить в Иерусалим; вот боги твои, Израиль, которые вывели тебя из земли Египетской.
1KGS|12|29|И поставил одного в Вефиле, а другого в Дане.
1KGS|12|30|И повело это ко греху, ибо народ стал ходить к одному [из] [них], даже в Дан.
1KGS|12|31|И построил он капище на высоте и поставил из народа священников, которые не были из сынов Левииных.
1KGS|12|32|И установил Иеровоам праздник в восьмой месяц, в пятнадцатый день месяца, подобный тому празднику, какой был в Иудее, и приносил жертвы на жертвеннике; то же сделал он в Вефиле, чтобы приносить жертву тельцам, которых сделал. И поставил в Вефиле священников высот, которые устроил,
1KGS|12|33|и принес жертвы на жертвеннике, который он сделал в Вефиле, в пятнадцатый день восьмого месяца, месяца, который он произвольно назначил; и установил праздник для сынов Израилевых, и подошел к жертвеннику, чтобы совершить курение.
1KGS|13|1|И вот, человек Божий пришел из Иудеи по слову Господню в Вефиль, в то время, как Иеровоам стоял у жертвенника, чтобы совершить курение.
1KGS|13|2|И произнес к жертвеннику слово Господне и сказал: жертвенник, жертвенник! так говорит Господь: вот, родится сын дому Давидову, имя ему Иосия, и принесет на тебе в жертву священников высот, совершающих на тебе курение, и человеческие кости сожжет на тебе.
1KGS|13|3|И дал в тот день знамение, сказав: вот знамение того, что это изрек Господь: вот, этот жертвенник распадется, и пепел, который на нем, рассыплется.
1KGS|13|4|Когда царь услышал слово человека Божия, произнесенное к жертвеннику в Вефиле, то простер Иеровоам руку свою от жертвенника, говоря: возьмите его. И одеревенела рука его, которую он простер на него, и не мог он поворотить ее к себе.
1KGS|13|5|И жертвенник распался, и пепел с жертвенника рассыпался, по знамению, которое дал человек Божий словом Господним.
1KGS|13|6|И сказал царь человеку Божию: умилостиви лице Господа Бога твоего и помолись обо мне, чтобы рука моя могла поворотиться ко мне. И умилостивил человек Божий лице Господа, и рука царя поворотилась к нему и стала, как прежде.
1KGS|13|7|И сказал царь человеку Божию: зайди со мною в дом и подкрепи себя пищею, и я дам тебе подарок.
1KGS|13|8|Но человек Божий сказал царю: хотя бы ты давал мне полдома твоего, я не пойду с тобою и не буду есть хлеба и не буду пить воды в этом месте,
1KGS|13|9|ибо так заповедано мне словом Господним: "не ешь там хлеба и не пей воды и не возвращайся тою дорогою, которою ты шел".
1KGS|13|10|И пошел он другою дорогою и не пошел обратно тою дорогою, которою пришел в Вефиль.
1KGS|13|11|В Вефиле жил один пророк–старец. Сын его пришел и рассказал ему все, что сделал сегодня человек Божий в Вефиле; и слова, какие он говорил царю, пересказали [сыновья] отцу своему.
1KGS|13|12|И спросил их отец их: какою дорогою он пошел? И показали сыновья его, какою дорогою пошел человек Божий, приходивший из Иудеи.
1KGS|13|13|И сказал он сыновьям своим: оседлайте мне осла. И оседлали ему осла, и он сел на него.
1KGS|13|14|И поехал за человеком Божиим, и нашел его сидящего под дубом, и сказал ему: ты ли человек Божий, пришедший из Иудеи? И сказал тот: я.
1KGS|13|15|И сказал ему: зайди ко мне в дом и поешь хлеба.
1KGS|13|16|Тот сказал: я не могу возвратиться с тобою и пойти к тебе; не буду есть хлеба и не буду пить у тебя воды в сем месте,
1KGS|13|17|ибо словом Господним сказано мне: "не ешь хлеба и не пей там воды и не возвращайся тою дорогою, которою ты шел".
1KGS|13|18|И сказал он ему: и я пророк такой же, как ты, и Ангел говорил мне словом Господним, и сказал: "вороти его к себе в дом; пусть поест он хлеба и напьется воды". – Он солгал ему.
1KGS|13|19|И тот воротился с ним, и поел хлеба в его доме, и напился воды.
1KGS|13|20|Когда они еще сидели за столом, слово Господне было к пророку, воротившему его.
1KGS|13|21|И произнес он к человеку Божию, пришедшему из Иудеи, и сказал: так говорит Господь: за то, что ты не повиновался устам Господа и не соблюл повеления, которое заповедал тебе Господь Бог твой,
1KGS|13|22|но воротился, ел хлеб и пил воду в том месте, о котором Он сказал тебе: "не ешь хлеба и не пей воды", тело твое не войдет в гробницу отцов твоих.
1KGS|13|23|После того, как тот поел хлеба и напился, он оседлал осла для пророка, которого он воротил.
1KGS|13|24|И отправился тот. И встретил его на дороге лев и умертвил его. И лежало тело его, брошенное на дороге; осел же стоял подле него, и лев стоял подле тела.
1KGS|13|25|И вот, проходившие мимо люди увидели тело, брошенное на дороге, и льва, стоящего подле тела, и пошли и рассказали в городе, в котором жил пророк–старец.
1KGS|13|26|Пророк, воротивший его с дороги, услышав [это], сказал: это тот человек Божий, который не повиновался устам Господа; Господь предал его льву, который изломал его и умертвил его, по слову Господа, которое Он изрек ему.
1KGS|13|27|И сказал сыновьям своим: оседлайте мне осла. И оседлали они.
1KGS|13|28|Он отправился и нашел тело его, брошенное на дороге; осел же и лев стояли подле тела; лев не съел тела и не изломал осла.
1KGS|13|29|И поднял пророк тело человека Божия, и положил его на осла, и повез его обратно. И пошел пророк–старец в город [свой], чтобы оплакать и похоронить его.
1KGS|13|30|И положил тело его в своей гробнице и плакал по нем: увы, брат мой!
1KGS|13|31|После погребения его он сказал сыновьям своим: когда я умру, похороните меня в гробнице, в которой погребен человек Божий; подле костей его положите кости мои;
1KGS|13|32|ибо сбудется слово, которое он по повелению Господню произнес о жертвеннике в Вефиле и о всех капищах на высотах, в городах Самарийских.
1KGS|13|33|И после сего события Иеровоам не сошел со своей худой дороги, но продолжал ставить из народа священников высот; кто хотел, того он посвящал, и тот становился священником высот.
1KGS|13|34|Это вело дом Иеровоамов ко греху и к погибели и к истреблению его с лица земли.
1KGS|14|1|В то время заболел Авия, сын Иеровоамов.
1KGS|14|2|И сказал Иеровоам жене своей: встань и переоденься, чтобы не узнали, что ты жена Иеровоамова, и пойди в Силом. Там есть пророк Ахия; он предсказал мне, что я буду царем сего народа.
1KGS|14|3|И возьми с собою десять хлебов, и лепешек, и кувшин меду, и пойди к нему: он скажет тебе, что будет с отроком.
1KGS|14|4|Жена Иеровоама так и сделала: встала, пошла в Силом и пришла в дом Ахии. Ахия уже не мог видеть, ибо глаза его сделались неподвижны от старости.
1KGS|14|5|И сказал Господь Ахии: вот, идет жена Иеровоамова спросить тебя о сыне своем, ибо он болен; так и так говори ей; она придет переодетая.
1KGS|14|6|Ахия, услышав шорох от ног ее, когда она вошла в дверь, сказал: войди, жена Иеровоамова; для чего было тебе переодеваться? Я грозный посланник к тебе.
1KGS|14|7|Пойди, скажи Иеровоаму: так говорит Господь Бог Израилев: Я возвысил тебя из среды простого народа и поставил вождем народа Моего Израиля,
1KGS|14|8|и отторг царство от дома Давидова и дал его тебе; а ты не таков, как раб Мой Давид, который соблюдал заповеди Мои и который последовал Мне всем сердцем своим, делая только угодное пред очами Моими;
1KGS|14|9|ты поступал хуже всех, которые были прежде тебя, и пошел, и сделал себе иных богов и истуканов, чтобы раздражить Меня, Меня же отбросил назад;
1KGS|14|10|за это Я наведу беды на дом Иеровоамов и истреблю у Иеровоама [до] мочащегося к стене, заключенного и оставшегося в Израиле, и вымету дом Иеровоамов, как выметают сор, дочиста;
1KGS|14|11|кто умрет у Иеровоама в городе, того съедят псы, а кто умрет на поле, того склюют птицы небесные; так Господь сказал.
1KGS|14|12|Встань и иди в дом твой; и как скоро нога твоя ступит в город, умрет дитя;
1KGS|14|13|и оплачут его все Израильтяне и похоронят его, ибо он один у Иеровоама войдет в гробницу, так как в нем, из дома Иеровоамова, нашлось нечто доброе пред Господом Богом Израилевым.
1KGS|14|14|И восставит Себе Господь над Израилем царя, который истребит дом Иеровоамов в тот день; и что? даже теперь.
1KGS|14|15|И поразит Господь Израиля, и [будет он], как тростник, колеблемый в воде, и извергнет Израильтян из этой доброй земли, которую дал отцам их, и развеет их за реку, за то, что они сделали у себя идолов, раздражая Господа;
1KGS|14|16|и предаст [Господь] Израиля за грехи Иеровоама, которые он сам сделал и которыми ввел в грех Израиля.
1KGS|14|17|И встала жена Иеровоамова, и пошла, и пришла в Фирцу; и лишь только переступила чрез порог дома, дитя умерло.
1KGS|14|18|И похоронили его, и оплакали его все Израильтяне, по слову Господа, которое Он изрек чрез раба Своего Ахию пророка.
1KGS|14|19|Прочие дела Иеровоама, как он воевал и как царствовал, описаны в летописи царей Израильских.
1KGS|14|20|Времени царствования Иеровоамова было двадцать два года; и почил он с отцами своими, и воцарился Нават, сын его, вместо него.
1KGS|14|21|Ровоам, сын Соломонов, царствовал в Иудее. Сорок один год было Ровоаму, когда он воцарился, и семнадцать лет царствовал в Иерусалиме, в городе, который избрал Господь из всех колен Израилевых, чтобы пребывало там имя Его. Имя матери его Наама Аммонитянка.
1KGS|14|22|И делал Иуда неугодное пред очами Господа, и раздражали Его более всего того, что сделали отцы их своими грехами, какими они грешили.
1KGS|14|23|И устроили они у себя высоты и статуи и капища на всяком высоком холме и под всяким тенистым деревом.
1KGS|14|24|И блудники были также в этой земле и делали все мерзости тех народов, которых Господь прогнал от лица сынов Израилевых.
1KGS|14|25|На пятом году царствования Ровоамова, Сусаким, царь Египетский, вышел против Иерусалима
1KGS|14|26|и взял сокровища дома Господня и сокровища дома царского, – Все взял; взял и все золотые щиты, которые сделал Соломон.
1KGS|14|27|И сделал царь Ровоам вместо них медные щиты и отдал их на руки начальникам телохранителей, которые охраняли вход в дом царя.
1KGS|14|28|Когда царь выходил в дом Господень, телохранители несли их, и потом опять относили их в палату телохранителей.
1KGS|14|29|Прочее о Ровоаме и обо всем, что он делал, описано в летописи царей Иудейских.
1KGS|14|30|Между Ровоамом и Иеровоамом была война во все дни [жизни их].
1KGS|14|31|И почил Ровоам с отцами своими и погребен с отцами своими в городе Давидовом. Имя матери его Наама Аммонитянка. И воцарился Авия, сын его, вместо него.
1KGS|15|1|В восемнадцатый год царствования Иеровоама, сына Наватова, Авия воцарился над Иудеями.
1KGS|15|2|Три года он царствовал в Иерусалиме; имя матери его Мааха, дочь Авессалома.
1KGS|15|3|Он ходил во всех грехах отца своего, которые тот делал прежде него, и сердце его не было предано Господу Богу его, как сердце Давида, отца его.
1KGS|15|4|Но ради Давида Господь Бог его дал ему светильник в Иерусалиме, восставив по нем сына его и утвердив Иерусалим,
1KGS|15|5|потому что Давид делал угодное пред очами Господа и не отступал от всего того, что Он заповедал ему, во все дни жизни своей, кроме поступка с Уриею Хеттеянином.
1KGS|15|6|И война была между Ровоамом и Иеровоамом во все дни жизни их.
1KGS|15|7|Прочие дела Авии, все, что он сделал, описано в летописи царей Иудейских. И была война между Авиею и Иеровоамом.
1KGS|15|8|И почил Авия с отцами своими, и похоронили его в городе Давидовом. И воцарился Аса, сын его, вместо него.
1KGS|15|9|В двадцатый год [царствования] Иеровоама, царя Израильского, воцарился Аса над Иудеями
1KGS|15|10|и сорок один год царствовал в Иерусалиме; имя матери его Ана, дочь Авессалома.
1KGS|15|11|Аса делал угодное пред очами Господа, как Давид, отец его.
1KGS|15|12|Он изгнал блудников из земли и отверг всех идолов, которых сделали отцы его,
1KGS|15|13|и даже мать свою Ану лишил звания царицы за то, что она сделала истукан Астарты; и изрубил Аса истукан ее и сжег у потока Кедрона.
1KGS|15|14|Высоты же не были уничтожены. Но сердце Асы было предано Господу во все дни его.
1KGS|15|15|И внес он в дом Господень вещи, посвященные отцом его, и вещи, посвященные им: серебро и золото и сосуды.
1KGS|15|16|И война была между Асою и Ваасою, царем Израильским, во все дни их.
1KGS|15|17|И вышел Вааса, царь Израильский, против Иудеи и начал строить Раму, чтобы никто не выходил и не уходил к Асе, царю Иудейскому.
1KGS|15|18|И взял Аса все серебро и золото, остававшееся в сокровищницах дома Господня и в сокровищницах дома царского, и дал его в руки слуг своих, и послал их царь Аса к Венададу, сыну Тавримона, сына Хезионова, царю Сирийскому, жившему в Дамаске, и сказал:
1KGS|15|19|союз да будет между мною и между тобою, [как был] между отцом моим и между отцом твоим; вот, я посылаю тебе в дар серебро и золото; расторгни союз твой с Ваасою, царем Израильским, чтобы он отошел от меня.
1KGS|15|20|И послушался Венадад царя Асы, и послал военачальников своих против городов Израильских, и поразил Аин и Дан и Авел–Беф–Мааху и весь Киннероф, по всей земле Неффалима.
1KGS|15|21|Услышав [о сем], Вааса перестал строить Раму и возвратился в Фирцу.
1KGS|15|22|Царь же Аса созвал всех Иудеев, никого не исключая, и вынесли они из Рамы камни и дерева, которые Вааса употреблял для строения. И выстроил из них царь Аса Гиву Вениаминову и Мицпу.
1KGS|15|23|Все прочие дела Асы и все подвиги его, и все, что он сделал, и города, которые он построил, описаны в летописи царей Иудейских, кроме того, что в старости своей он был болен ногами.
1KGS|15|24|И почил Аса с отцами своими и погребен с отцами своими в городе Давида, отца своего. И воцарился Иосафат, сын его, вместо него.
1KGS|15|25|Нават же, сын Иеровоамов, воцарился над Израилем во второй год Асы, царя Иудейского, и царствовал над Израилем два года.
1KGS|15|26|И делал он неугодное пред очами Господа, ходил путем отца своего и во грехах его, которыми тот ввел Израиля в грех.
1KGS|15|27|И сделал против него заговор Вааса, сын Ахии, из дома Иссахарова, и убил его Вааса при Гавафоне Филистимском, когда Нават и все Израильтяне осаждали Гавафон:
1KGS|15|28|и умертвил его Вааса в третий год Асы, царя Иудейского, и воцарился вместо него.
1KGS|15|29|Когда он воцарился, то избил весь дом Иеровоамов, не оставил ни души у Иеровоама, доколе не истребил его, по слову Господа, которое Он изрек чрез раба Своего Ахию Силомлянина,
1KGS|15|30|за грехи Иеровоама, которые он сам делал и которыми ввел в грех Израиля, за оскорбление, которым он прогневал Господа Бога Израилева.
1KGS|15|31|Прочие дела Навата, все, что он сделал, описано в летописи царей Израильских.
1KGS|15|32|И война была между Асою и Ваасою, царем Израильским, во все дни их.
1KGS|15|33|В третий год Асы, царя Иудейского, воцарился Вааса, сын Ахии, над всеми Израильтянами в Фирце [и царствовал] двадцать четыре года.
1KGS|15|34|И делал неугодное пред очами Господними и ходил путем Иеровоама и во грехах его, которыми тот ввел в грех Израиля.
1KGS|16|1|И было слово Господне к Иую, сыну Ананиеву, о Ваасе:
1KGS|16|2|за то, что Я поднял тебя из праха и сделал тебя вождем народа Моего Израиля, ты же пошел путем Иеровоама и ввел в грех народ Мой Израильтян, чтобы он прогневлял Меня грехами своими,
1KGS|16|3|вот, Я отвергну дом Ваасы и дом потомства его и сделаю с домом твоим то же, что с домом Иеровоама, сына Наватова;
1KGS|16|4|кто умрет у Ваасы в городе, того съедят псы; а кто умрет у него на поле, того склюют птицы небесные.
1KGS|16|5|Прочие дела Ваасы, все, что он сделал, и подвиги его описаны в летописи царей Израильских.
1KGS|16|6|И почил Вааса с отцами своими, и погребен в Фирце. И воцарился Ила, сын его, вместо него.
1KGS|16|7|Но чрез Иуя, сына Ананиева, уже было [сказано] слово Господне о Ваасе и о доме его и о всем зле, какое он делал пред очами Господа, раздражая Его делами рук своих, подражая дому Иеровоамову, за что он истреблен был.
1KGS|16|8|В двадцать шестой год Асы, царя Иудейского, воцарился Ила, сын Ваасы, над Израилем в Фирце, [и царствовал] два года.
1KGS|16|9|И составил против него заговор раб его Замврий, начальствовавший над половиною колесниц. Когда он в Фирце напился допьяна в доме Арсы, начальствующего над дворцом в Фирце,
1KGS|16|10|тогда вошел Замврий, поразил его и умертвил его, в двадцать седьмой год Асы, царя Иудейского, и воцарился вместо него.
1KGS|16|11|Когда он воцарился и сел на престоле его, то истребил весь дом Ваасы, не оставив ему мочащегося к стене, ни родственников его, ни друзей его.
1KGS|16|12|И истребил Замврий весь дом Ваасы, по слову Господа, которое Он изрек о Ваасе чрез Иуя пророка,
1KGS|16|13|за все грехи Ваасы и за грехи Илы, сына его, которые они сами делали и которыми вводили Израиля в грех, раздражая Господа Бога Израилева своими идолами.
1KGS|16|14|Прочие дела Илы, все, что он сделал, описано в летописи царей Израильских.
1KGS|16|15|В двадцать седьмой год Асы, царя Иудейского, воцарился Замврий и царствовал семь дней в Фирце, когда народ осаждал Гавафон Филистимский.
1KGS|16|16|Когда народ осаждавший услышал, что Замврий сделал заговор и умертвил царя, то все Израильтяне воцарили Амврия, военачальника, над Израилем в тот же день, в стане.
1KGS|16|17|И отступили Амврий и все Израильтяне с ним от Гавафона и осадили Фирцу.
1KGS|16|18|Когда увидел Замврий, что город взят, вошел во внутреннюю комнату царского дома и зажег за собою царский дом огнем и погиб
1KGS|16|19|за свои грехи, в чем он согрешил, делая неугодное пред очами Господними, ходя путем Иеровоама и во грехах его, которые тот сделал, чтобы ввести Израиля в грех.
1KGS|16|20|Прочие дела Замврия и заговор его, который он составил, описаны в летописи царей Израильских.
1KGS|16|21|Тогда разделился народ Израильский надвое: половина народа стояла за Фамния, сына Гонафова, чтобы воцарить его, а половина за Амврия.
1KGS|16|22|И одержал верх народ, который за Амврия, над народом, который за Фамния, сына Гонафова, и умер Фамний, и воцарился Амврий.
1KGS|16|23|В тридцать первый год Асы, царя Иудейского, воцарился Амврий над Израилем [и царствовал] двенадцать лет. В Фирце он царствовал шесть лет.
1KGS|16|24|И купил Амврий гору Семерон у Семира за два таланта серебра, и застроил гору, и назвал построенный им город Самариею, по имени Семира, владельца горы.
1KGS|16|25|И делал Амврий неугодное пред очами Господа и поступал хуже всех бывших перед ним.
1KGS|16|26|Он во всем ходил путем Иеровоама, сына Наватова, и во грехах его, которыми тот ввел в грех Израильтян, чтобы прогневлять Господа Бога Израилева идолами своими.
1KGS|16|27|Прочие дела Амврия, которые он сделал, и мужество, которое он показал, описаны в летописи царей Израильских.
1KGS|16|28|И почил Амврий с отцами своими и погребен в Самарии. И воцарился Ахав, сын его, вместо него.
1KGS|16|29|Ахав, сын Амвриев, воцарился над Израилем в тридцать восьмой год Асы, царя Иудейского, и царствовал Ахав, сын Амврия, над Израилем в Самарии двадцать два года.
1KGS|16|30|И делал Ахав, сын Амврия, неугодное пред очами Господа более всех бывших прежде него.
1KGS|16|31|Мало было для него впадать в грехи Иеровоама, сына Наватова; он взял себе в жену Иезавель, дочь Ефваала царя Сидонского, и стал служить Ваалу и поклоняться ему.
1KGS|16|32|И поставил он Ваалу жертвенник в капище Ваала, который построил в Самарии.
1KGS|16|33|И сделал Ахав дубраву, и более всех царей Израильских, которые были прежде него, Ахав делал то, что раздражает Господа Бога Израилева.
1KGS|16|34|В его дни Ахиил Вефилянин построил Иерихон: на первенце своем Авираме он положил основание его и на младшем своем [сыне] Сегубе поставил ворота его, по слову Господа, которое Он изрек чрез Иисуса, сына Навина.
1KGS|17|1|И сказал Илия Фесвитянин, из жителей Галаадских, Ахаву: жив Господь Бог Израилев, пред Которым я стою! в сии годы не будет ни росы, ни дождя, разве только по моему слову.
1KGS|17|2|И было к нему слово Господне:
1KGS|17|3|пойди отсюда и обратись на восток и скройся у потока Хорафа, что против Иордана;
1KGS|17|4|из этого потока ты будешь пить, а воронам Я повелел кормить тебя там.
1KGS|17|5|И пошел он и сделал по слову Господню; пошел и остался у потока Хорафа, что против Иордана.
1KGS|17|6|И вороны приносили ему хлеб и мясо поутру, и хлеб и мясо по вечеру, а из потока он пил.
1KGS|17|7|По прошествии некоторого времени этот поток высох, ибо не было дождя на землю.
1KGS|17|8|И было к нему слово Господне:
1KGS|17|9|встань и пойди в Сарепту Сидонскую, и оставайся там; Я повелел там женщине вдове кормить тебя.
1KGS|17|10|И встал он и пошел в Сарепту; и когда пришел к воротам города, вот, там женщина вдова собирает дрова. И подозвал он ее и сказал: дай мне немного воды в сосуде напиться.
1KGS|17|11|И пошла она, чтобы взять; а он закричал вслед ей и сказал: возьми для меня и кусок хлеба в руки свои.
1KGS|17|12|Она сказала: жив Господь Бог твой! у меня ничего нет печеного, а только есть горсть муки в кадке и немного масла в кувшине; и вот, я наберу полена два дров, и пойду, и приготовлю это для себя и для сына моего; съедим это и умрем.
1KGS|17|13|И сказал ей Илия: не бойся, пойди, сделай, что ты сказала; но прежде из этого сделай небольшой опреснок для меня и принеси мне; а для себя и для своего сына сделаешь после;
1KGS|17|14|ибо так говорит Господь Бог Израилев: мука в кадке не истощится, и масло в кувшине не убудет до того дня, когда Господь даст дождь на землю.
1KGS|17|15|И пошла она и сделала так, как сказал Илия; и кормилась она, и он, и дом ее несколько времени.
1KGS|17|16|Мука в кадке не истощалась, и масло в кувшине не убывало, по слову Господа, которое Он изрек чрез Илию.
1KGS|17|17|После этого заболел сын этой женщины, хозяйки дома, и болезнь его была так сильна, что не осталось в нем дыхания.
1KGS|17|18|И сказала она Илии: что мне и тебе, человек Божий? ты пришел ко мне напомнить грехи мои и умертвить сына моего.
1KGS|17|19|И сказал он ей: дай мне сына твоего. И взял его с рук ее, и понес его в горницу, где он жил, и положил его на свою постель,
1KGS|17|20|и воззвал к Господу и сказал: Господи Боже мой! неужели Ты и вдове, у которой я пребываю, сделаешь зло, умертвив сына ее?
1KGS|17|21|И простершись над отроком трижды, он воззвал к Господу и сказал: Господи Боже мой! да возвратится душа отрока сего в него!
1KGS|17|22|И услышал Господь голос Илии, и возвратилась душа отрока сего в него, и он ожил.
1KGS|17|23|И взял Илия отрока, и свел его из горницы в дом, и отдал его матери его, и сказал Илия: смотри, сын твой жив.
1KGS|17|24|И сказала та женщина Илии: теперь–то я узнала, что ты человек Божий, и что слово Господне в устах твоих истинно.
1KGS|18|1|По прошествии многих дней было слово Господне к Илии в третий год: пойди и покажись Ахаву, и Я дам дождь на землю.
1KGS|18|2|И пошел Илия, чтобы показаться Ахаву. Голод же сильный был в Самарии.
1KGS|18|3|И призвал Ахав Авдия, начальствовавшего над дворцом. Авдий же был человек весьма богобоязненный,
1KGS|18|4|и когда Иезавель истребляла пророков Господних, Авдий взял сто пророков, и скрывал их, по пятидесяти человек, в пещерах, и питал их хлебом и водою.
1KGS|18|5|И сказал Ахав Авдию: пойди по земле ко всем источникам водным и ко всем потокам на земле, не найдем ли где травы, чтобы нам прокормить коней и лошаков и не лишиться скота.
1KGS|18|6|И разделили они между собою землю, чтобы обойти ее: Ахав особо пошел одною дорогою, и Авдий особо пошел другою дорогою.
1KGS|18|7|Когда Авдий шел дорогою, вот, навстречу ему идет Илия. Он узнал его и пал на лице свое и сказал: ты ли это, господин мой Илия?
1KGS|18|8|Тот сказал ему: я; пойди, скажи господину твоему: "Илия здесь".
1KGS|18|9|Он сказал: чем я провинился, что ты предаешь раба твоего в руки Ахава, чтоб умертвить меня?
1KGS|18|10|Жив Господь Бог твой! нет ни одного народа и царства, куда бы не посылал государь мой искать тебя; и когда ему говорили, [что тебя] нет, он брал клятву с того царства и народа, что не могли отыскать тебя;
1KGS|18|11|а ты теперь говоришь: "пойди, скажи господину твоему: Илия здесь".
1KGS|18|12|Когда я пойду от тебя, тогда Дух Господень унесет тебя, не знаю, куда; и если я пойду уведомить Ахава, и он не найдет тебя, то он убьет меня; а раб твой богобоязнен от юности своей.
1KGS|18|13|Разве не сказано господину моему, что я сделал, когда Иезавель убивала пророков Господних, как я скрывал сто человек пророков Господних, по пятидесяти человек, в пещерах и питал их хлебом и водою?
1KGS|18|14|А ты теперь говоришь: "пойди, скажи господину твоему: Илия здесь"; он убьет меня.
1KGS|18|15|И сказал Илия: жив Господь Саваоф, пред Которым я стою! сегодня я покажусь ему.
1KGS|18|16|И пошел Авдий навстречу Ахаву и донес ему. И пошел Ахав навстречу Илии.
1KGS|18|17|Когда Ахав увидел Илию, то сказал Ахав ему: ты ли это, смущающий Израиля?
1KGS|18|18|И сказал Илия: не я смущаю Израиля, а ты и дом отца твоего, тем, что вы презрели повеления Господни и идете вслед Ваалам;
1KGS|18|19|теперь пошли и собери ко мне всего Израиля на гору Кармил, и четыреста пятьдесят пророков Вааловых, и четыреста пророков дубравных, питающихся от стола Иезавели.
1KGS|18|20|И послал Ахав ко всем сынам Израилевым и собрал всех пророков на гору Кармил.
1KGS|18|21|И подошел Илия ко всему народу и сказал: долго ли вам хромать на оба колена? если Господь есть Бог, то последуйте Ему; а если Ваал, то ему последуйте. И не отвечал народ ему ни слова.
1KGS|18|22|И сказал Илия народу: я один остался пророк Господень, а пророков Вааловых четыреста пятьдесят человек.
1KGS|18|23|пусть дадут нам двух тельцов, и пусть они выберут себе одного тельца, и рассекут его, и положат на дрова, но огня пусть не подкладывают; а я приготовлю другого тельца и положу на дрова, а огня не подложу;
1KGS|18|24|и призовите вы имя бога вашего, а я призову имя Господа Бога моего. Тот Бог, Который даст ответ посредством огня, есть Бог. И отвечал весь народ и сказал: хорошо.
1KGS|18|25|И сказал Илия пророкам Вааловым: выберите себе одного тельца и приготовьте вы прежде, ибо вас много; и призовите имя бога вашего, но огня не подкладывайте.
1KGS|18|26|И взяли они тельца, который дан был им, и приготовили, и призывали имя Ваала от утра до полудня, говоря: Ваале, услышь нас! Но не было ни голоса, ни ответа. И скакали они у жертвенника, который сделали.
1KGS|18|27|В полдень Илия стал смеяться над ними и говорил: кричите громким голосом, ибо он бог; может быть, он задумался, или занят чем–либо, или в дороге, а может быть, и спит, так он проснется!
1KGS|18|28|И стали они кричать громким голосом, и кололи себя по своему обыкновению ножами и копьями, так что кровь лилась по ним.
1KGS|18|29|Прошел полдень, а они все еще бесновались до самого времени вечернего жертвоприношения; но не было ни голоса, ни ответа, ни слуха.
1KGS|18|30|Тогда Илия сказал всему народу: подойдите ко мне. И подошел весь народ к нему. Он восстановил разрушенный жертвенник Господень.
1KGS|18|31|И взял Илия двенадцать камней, по числу колен сынов Иакова, которому Господь сказал так: Израиль будет имя твое.
1KGS|18|32|И построил из сих камней жертвенник во имя Господа, и сделал вокруг жертвенника ров, вместимостью в две саты зерен,
1KGS|18|33|и положил дрова, и рассек тельца, и возложил его на дрова,
1KGS|18|34|и сказал: наполните четыре ведра воды и выливайте на всесожигаемую жертву и на дрова. Потом сказал: повторите. И они повторили. И сказал: сделайте [то же] в третий раз. И сделали в третий раз,
1KGS|18|35|и вода полилась вокруг жертвенника, и ров наполнился водою.
1KGS|18|36|Во время приношения вечерней жертвы подошел Илия пророк и сказал: Господи, Боже Авраамов, Исааков и Израилев! Да познают в сей день, что Ты один Бог в Израиле, и что я раб Твой и сделал все по слову Твоему.
1KGS|18|37|Услышь меня, Господи, услышь меня! Да познает народ сей, что Ты, Господи, Бог, и Ты обратишь сердце их [к Тебе].
1KGS|18|38|И ниспал огонь Господень и пожрал всесожжение, и дрова, и камни, и прах, и поглотил воду, которая во рве.
1KGS|18|39|Увидев [это], весь народ пал на лице свое и сказал: Господь есть Бог, Господь есть Бог!
1KGS|18|40|И сказал им Илия: схватите пророков Вааловых, чтобы ни один из них не укрылся. И схватили их, и отвел их Илия к потоку Киссону и заколол их там.
1KGS|18|41|И сказал Илия Ахаву: пойди, ешь и пей, ибо слышен шум дождя.
1KGS|18|42|И пошел Ахав есть и пить, а Илия взошел на верх Кармила и наклонился к земле, и положил лице свое между коленами своими,
1KGS|18|43|и сказал отроку своему: пойди, посмотри к морю. Тот пошел и посмотрел, и сказал: ничего нет. Он сказал: продолжай [это] до семи раз.
1KGS|18|44|В седьмой раз тот сказал: вот, небольшое облако поднимается от моря, величиною в ладонь человеческую. Он сказал: пойди, скажи Ахаву: "запрягай [колесницу твою] и поезжай, чтобы не застал тебя дождь".
1KGS|18|45|Между тем небо сделалось мрачно от туч и от ветра, и пошел большой дождь. Ахав же сел в колесницу, и поехал в Изреель.
1KGS|18|46|И была на Илии рука Господня. Он опоясал чресла свои и бежал пред Ахавом до самого Изрееля.
1KGS|19|1|И пересказал Ахав Иезавели все, что сделал Илия, и то, что он убил всех пророков мечом.
1KGS|19|2|И послала Иезавель посланца к Илии сказать: пусть то и то сделают мне боги, и еще больше сделают, если я завтра к этому времени не сделаю с твоею душею того, что [сделано] с душею каждого из них.
1KGS|19|3|Увидев это, он встал и пошел, чтобы спасти жизнь свою, и пришел в Вирсавию, которая в Иудее, и оставил отрока своего там.
1KGS|19|4|А сам отошел в пустыню на день пути и, придя, сел под можжевеловым кустом, и просил смерти себе и сказал: довольно уже, Господи; возьми душу мою, ибо я не лучше отцов моих.
1KGS|19|5|И лег и заснул под можжевеловым кустом. И вот, Ангел коснулся его и сказал ему: встань, ешь.
1KGS|19|6|И взглянул Илия, и вот, у изголовья его печеная лепешка и кувшин воды. Он поел и напился и опять заснул.
1KGS|19|7|И возвратился Ангел Господень во второй раз, коснулся его и сказал: встань, ешь; ибо дальняя дорога пред тобою.
1KGS|19|8|И встал он, поел и напился, и, подкрепившись тою пищею, шел сорок дней и сорок ночей до горы Божией Хорива.
1KGS|19|9|И вошел он там в пещеру и ночевал в ней. И вот, было к нему слово Господне, и сказал ему [Господь]: что ты здесь, Илия?
1KGS|19|10|Он сказал: возревновал я о Господе Боге Саваофе, ибо сыны Израилевы оставили завет Твой, разрушили Твои жертвенники и пророков Твоих убили мечом; остался я один, но и моей души ищут, чтобы отнять ее.
1KGS|19|11|И сказал: выйди и стань на горе пред лицем Господним, и вот, Господь пройдет, и большой и сильный ветер, раздирающий горы и сокрушающий скалы пред Господом, но не в ветре Господь; после ветра землетрясение, но не в землетрясении Господь;
1KGS|19|12|после землетрясения огонь, но не в огне Господь; после огня веяние тихого ветра.
1KGS|19|13|Услышав [сие], Илия закрыл лице свое милотью своею, и вышел, и стал у входа в пещеру. И был к нему голос и сказал ему: что ты здесь, Илия?
1KGS|19|14|Он сказал: возревновал я о Господе Боге Саваофе, ибо сыны Израилевы оставили завет Твой, разрушили жертвенники Твои и пророков Твоих убили мечом; остался я один, но и моей души ищут, чтоб отнять ее.
1KGS|19|15|И сказал ему Господь: пойди обратно своею дорогою чрез пустыню в Дамаск, и когда придешь, то помажь Азаила в царя над Сириею,
1KGS|19|16|а Ииуя, сына Намессиина, помажь в царя над Израилем; Елисея же, сына Сафатова, из Авел–Мехолы, помажь в пророка вместо себя;
1KGS|19|17|кто убежит от меча Азаилова, того умертвит Ииуй; а кто спасется от меча Ииуева, того умертвит Елисей.
1KGS|19|18|Впрочем, Я оставил между Израильтянами семь тысяч [мужей]; всех сих колени не преклонялись пред Ваалом, и всех сих уста не лобызали его.
1KGS|19|19|И пошел он оттуда, и нашел Елисея, сына Сафатова, когда он орал; двенадцать пар [волов] было у него, и сам он был при двенадцатой. Илия, проходя мимо него, бросил на него милоть свою.
1KGS|19|20|И оставил [Елисей] волов, и побежал за Илиею, и сказал: позволь мне поцеловать отца моего и мать мою, и я пойду за тобою. Он сказал ему: пойди и приходи назад, ибо что сделал я тебе?
1KGS|19|21|Он, отойдя от него, взял пару волов и заколол их и, зажегши плуг волов, изжарил мясо их, и роздал людям, и они ели. А сам встал и пошел за Илиею, и стал служить ему.
1KGS|20|1|Венадад, царь Сирийский, собрал все свое войско, и с ним были тридцать два царя, и кони и колесницы, и пошел, осадил Самарию и воевал против нее.
1KGS|20|2|И послал послов к Ахаву, царю Израильскому, в город,
1KGS|20|3|и сказал ему: так говорит Венадад: серебро твое и золото твое – мои, и жены твои и лучшие сыновья твои – мои.
1KGS|20|4|И отвечал царь Израильский и сказал: да будет по слову твоему, господин мой царь: я и все мое – твое.
1KGS|20|5|И опять пришли послы и сказали: так говорит Венадад: я послал к тебе сказать: "серебро твое, и золото твое, и жен твоих, и сыновей твоих отдай мне";
1KGS|20|6|поэтому я завтра, к этому времени, пришлю к тебе рабов моих, чтобы они осмотрели твой дом и домы служащих при тебе, и все дорогое для глаз твоих взяли в свои руки и унесли.
1KGS|20|7|И созвал царь Израильский всех старейшин земли и сказал: замечайте и смотрите, он замышляет зло; когда он присылал ко мне за женами моими, и сыновьями моими, и серебром моим, и золотом моим, я ему не отказал.
1KGS|20|8|И сказали ему все старейшины и весь народ: не слушай и не соглашайся.
1KGS|20|9|И сказал он послам Венадада: скажите господину моему царю: все, о чем ты присылал в первый раз к рабу твоему, я готов сделать, а этого не могу сделать. И пошли послы и отнесли ему ответ.
1KGS|20|10|И прислал к нему Венадад сказать: пусть то и то сделают мне боги, и еще больше сделают, если праха Самарийского достанет по горсти для всех людей, идущих за мною.
1KGS|20|11|И отвечал царь Израильский и сказал: скажите: пусть не хвалится подпоясывающийся, как распоясывающийся.
1KGS|20|12|Услышав это слово, Венадад, который пил вместе с царями в палатках, сказал рабам своим: осаждайте город. И они осадили город.
1KGS|20|13|И вот, один пророк подошел к Ахаву, царю Израильскому, и сказал: так говорит Господь: видишь ли все это большое полчище? вот, Я сегодня предам его в руку твою, чтобы ты знал, что Я Господь.
1KGS|20|14|И сказал Ахав: чрез кого? Он сказал: так говорит Господь: чрез слуг областных начальников. И сказал [Ахав]: кто начнет сражение? Он сказал: ты.
1KGS|20|15|[Ахав] счел слуг областных начальников, и нашлось их двести тридцать два; после них счел весь народ, всех сынов Израилевых, семь тысяч.
1KGS|20|16|И они выступили в полдень. Венадад же напился допьяна в палатках вместе с царями, с тридцатью двумя царями, помогавшими ему.
1KGS|20|17|И выступили прежде слуги областных начальников. И послал Венадад, и донесли ему, что люди вышли из Самарии.
1KGS|20|18|Он сказал: если за миром вышли они, то схватите их живыми, и если на войну вышли, также схватите их живыми.
1KGS|20|19|Вышли из города слуги областных начальников, и войско за ними.
1KGS|20|20|И поражал каждый противника своего; и побежали Сирияне, а Израильтяне погнались за ними. Венадад же, царь Сирийский, спасся на коне с всадниками.
1KGS|20|21|И вышел царь Израильский, и взял коней и колесниц, и произвел большое поражение у Сириян.
1KGS|20|22|И подошел пророк к царю Израильскому и сказал ему: пойди, укрепись, и знай и смотри, что тебе делать, ибо по прошествии года царь Сирийский опять пойдет против тебя.
1KGS|20|23|Слуги царя Сирийского сказали ему: Бог их есть Бог гор, поэтому они одолели нас; если же мы сразимся с ними на равнине, то верно одолеем их.
1KGS|20|24|Итак вот что сделай: удали царей, каждого с места его, и вместо них поставь областеначальников;
1KGS|20|25|и набери себе войска столько, сколько пало у тебя, и коней, сколько было коней, и колесниц, сколько было колесниц; и сразимся с ними на равнине, и тогда верно одолеем их. И послушался он голоса их и сделал так.
1KGS|20|26|По прошествии года Венадад собрал Сириян и выступил к Афеку, чтобы сразиться с Израилем.
1KGS|20|27|Собраны были и сыны Израилевы и, взяв продовольствие, пошли навстречу им. И расположились сыны Израилевы станом пред ними, как бы два небольшие стада коз, а Сирияне наполнили землю.
1KGS|20|28|И подошел человек Божий, и сказал царю Израильскому: так говорит Господь: за то, что Сирияне говорят: "Господь есть Бог гор, а не Бог долин", Я все это большое полчище предам в руку твою, чтобы вы знали, что Я – Господь.
1KGS|20|29|И стояли станом одни против других семь дней. В седьмой день началась битва, и сыны Израилевы поразили сто тысяч пеших Сириян в один день.
1KGS|20|30|Остальные убежали в город Афек; [там] упала стена на остальных двадцать семь тысяч человек. А Венадад ушел в город и бегал из одной внутренней комнаты в другую.
1KGS|20|31|И сказали ему слуги его: мы слышали, что цари дома Израилева цари милостивые; позволь нам возложить вретища на чресла свои и веревки на головы свои и пойти к царю Израильскому; может быть, он пощадит жизнь твою.
1KGS|20|32|И опоясали они вретищами чресла свои и возложили веревки на головы свои, и пришли к царю Израильскому и сказали: раб твой Венадад говорит: "пощади жизнь мою". Тот сказал: разве он жив? он брат мой.
1KGS|20|33|Люди сии приняли это за [хороший] знак и поспешно подхватили слово из уст его и сказали: брат твой Венадад. И сказал он: пойдите, приведите его. И вышел к нему Венадад, и он посадил его [с собою] на колесницу.
1KGS|20|34|И сказал ему [Венадад]: города, которые взял мой отец у твоего отца, я возвращу, и площади ты можешь иметь для себя в Дамаске, как отец мой имел в Самарии. [Ахав сказал]: после договора я отпущу тебя. И, заключив с ним договор, отпустил его.
1KGS|20|35|Тогда один человек из сынов пророческих сказал другому, по слову Господа: бей меня. Но этот человек не согласился бить его.
1KGS|20|36|И сказал ему: за то, что ты не слушаешь гласа Господня, убьет тебя лев, когда пойдешь от меня. Он пошел от него, и лев, встретив его, убил его.
1KGS|20|37|И нашел он другого человека, и сказал: бей меня. Этот человек бил его до того, что изранил побоями.
1KGS|20|38|И пошел пророк и предстал пред царя на дороге, прикрыв покрывалом глаза свои.
1KGS|20|39|Когда царь проезжал мимо, он закричал царю и сказал: раб твой ходил на сражение, и вот, один человек, отошедший в сторону, подвел ко мне человека и сказал: "стереги этого человека; если его не станет, то твоя душа будет за его душу, или ты должен будешь отвесить талант серебра".
1KGS|20|40|Когда раб твой занялся теми и другими делами, его не стало. – И сказал ему царь Израильский: таков тебе и приговор, ты сам решил.
1KGS|20|41|Он тотчас снял покрывало с глаз своих, и узнал его царь, что он из пророков.
1KGS|20|42|И сказал ему: так говорит Господь: за то, что ты выпустил из рук твоих человека, заклятого Мною, душа твоя будет вместо его души, народ твой вместо его народа.
1KGS|20|43|И отправился царь Израильский домой встревоженный и огорченный, и прибыл в Самарию.
1KGS|21|1|И было после сих происшествий: у Навуфея Изреелитянина в Изреели был виноградник подле дворца Ахава, царя Самарийского.
1KGS|21|2|И сказал Ахав Навуфею, говоря: отдай мне свой виноградник; из него будет у меня овощной сад, ибо он близко к моему дому; а вместо него я дам тебе виноградник лучше этого, или, если угодно тебе, дам тебе серебра, сколько он стоит.
1KGS|21|3|Но Навуфей сказал Ахаву: сохрани меня Господь, чтоб я отдал тебе наследство отцов моих!
1KGS|21|4|И пришел Ахав домой встревоженный и огорченный тем словом, которое сказал ему Навуфей Изреелитянин, говоря: не отдам тебе наследства отцов моих. И лег на постель свою, и отворотил лице свое, и хлеба не ел.
1KGS|21|5|И вошла к нему жена его Иезавель и сказала ему: отчего встревожен дух твой, что ты и хлеба не ешь?
1KGS|21|6|Он сказал ей: когда я стал говорить Навуфею Изреелитянину и сказал ему: "отдай мне виноградник твой за серебро, или, если хочешь, я дам тебе [другой] виноградник вместо него", тогда он сказал: "не отдам тебе виноградника моего".
1KGS|21|7|И сказала ему Иезавель, жена его: что за царство было бы в Израиле, если бы ты так поступал? встань, ешь хлеб и будь спокоен; я доставлю тебе виноградник Навуфея Изреелитянина.
1KGS|21|8|И написала она от имени Ахава письма, и запечатала их его печатью, и послала эти письма к старейшинам и знатным в его городе, живущим с Навуфеем.
1KGS|21|9|В письмах она писала так: объявите пост и посадите Навуфея на первое место в народе;
1KGS|21|10|и против него посадите двух негодных людей, которые свидетельствовали бы на него и сказали: "ты хулил Бога и царя"; и потом выведите его, и побейте его камнями, чтоб он умер.
1KGS|21|11|И сделали мужи города его, старейшины и знатные, жившие в городе его, как приказала им Иезавель, так, как писано в письмах, которые она послала к ним.
1KGS|21|12|Объявили пост и посадили Навуфея во главе народа;
1KGS|21|13|и выступили два негодных человека и сели против него, и свидетельствовали на него эти недобрые люди пред народом, и говорили: Навуфей хулил Бога и царя. И вывели его за город, и побили его камнями, и он умер.
1KGS|21|14|И послали к Иезавели сказать: Навуфей побит камнями и умер.
1KGS|21|15|Услышав, что Навуфей побит камнями и умер, Иезавель сказала Ахаву: встань, возьми во владение виноградник Навуфея Изреелитянина, который не хотел отдать тебе за серебро; ибо Навуфея нет в живых, он умер.
1KGS|21|16|Когда услышал Ахав, что Навуфей был убит, встал Ахав, чтобы пойти в виноградник Навуфея Изреелитянина и взять его во владение.
1KGS|21|17|И было слово Господне к Илии Фесвитянину:
1KGS|21|18|встань, пойди навстречу Ахаву, царю Израильскому, который в Самарии, вот, он теперь в винограднике Навуфея, куда пришел, чтобы взять [его] во владение;
1KGS|21|19|и скажи ему: "так говорит Господь: ты убил, и еще вступаешь в наследство?" и скажи ему: "так говорит Господь: на том месте, где псы лизали кровь Навуфея, псы будут лизать и твою кровь".
1KGS|21|20|И сказал Ахав Илии: нашел ты меня, враг мой! Он сказал: нашел, ибо ты предался тому, чтобы делать неугодное пред очами Господа.
1KGS|21|21|[Так говорит Господь]: вот, Я наведу на тебя беды и вымету за тобою и истреблю у Ахава мочащегося к стене и заключенного и оставшегося в Израиле.
1KGS|21|22|И поступлю с домом твоим так, как поступил Я с домом Иеровоама, сына Наватова, и с домом Ваасы, сына Ахиина, за оскорбление, которым ты раздражил [Меня] и ввел Израиля в грех.
1KGS|21|23|Также и о Иезавели сказал Господь: псы съедят Иезавель за стеною Изрееля.
1KGS|21|24|Кто умрет у Ахава в городе, того съедят псы, а кто умрет на поле, того расклюют птицы небесные;
1KGS|21|25|не было еще такого, как Ахав, который предался бы тому, чтобы делать неугодное пред очами Господа, к чему подущала его жена его Иезавель;
1KGS|21|26|он поступал весьма гнусно, последуя идолам, как делали Аморреи, которых Господь прогнал от лица сынов Израилевых.
1KGS|21|27|Выслушав все слова сии, Ахав разодрал одежды свои, и возложил на тело свое вретище, и постился, и спал во вретище, и ходил печально.
1KGS|21|28|И было слово Господне к Илии Фесвитянину, и сказал Господь:
1KGS|21|29|видишь, как смирился предо Мною Ахав? За то, что он смирился предо Мною, Я не наведу бед в его дни; во дни сына его наведу беды на дом его.
1KGS|22|1|Прожили три года, и не было войны между Сириею и Израилем.
1KGS|22|2|На третий год Иосафат, царь Иудейский, пошел к царю Израильскому.
1KGS|22|3|И сказал царь Израильский слугам своим: знаете ли, что Рамоф Галаадский наш? А мы так долго молчим, и не берем его из руки царя Сирийского.
1KGS|22|4|И сказал он Иосафату: пойдешь ли ты со мною на войну против Рамофа Галаадского? И сказал Иосафат царю Израильскому: как ты, так и я; как твой народ, так и мой народ; как твои кони, так и мои кони.
1KGS|22|5|И сказал Иосафат царю Израильскому: спроси сегодня, что скажет Господь.
1KGS|22|6|И собрал царь Израильский пророков, около четырехсот человек и сказал им: идти ли мне войною на Рамоф Галаадский, или нет? Они сказали: иди, Господь предаст [его] в руки царя.
1KGS|22|7|И сказал Иосафат: нет ли здесь еще пророка Господня, чтобы нам вопросить чрез него Господа?
1KGS|22|8|И сказал царь Израильский Иосафату: есть еще один человек, чрез которого можно вопросить Господа, но я не люблю его, ибо он не пророчествует о мне доброго, а только худое, – это Михей, сын Иемвлая. И сказал Иосафат: не говори, царь, так.
1KGS|22|9|И позвал царь Израильский одного евнуха и сказал: сходи поскорее за Михеем, сыном Иемвлая.
1KGS|22|10|Царь Израильский и Иосафат, царь Иудейский, сидели каждый на седалище своем, одетые в [царские] одежды, на площади у ворот Самарии, и все пророки пророчествовали пред ними.
1KGS|22|11|И сделал себе Седекия, сын Хенааны, железные рога, и сказал: так говорит Господь: сими избодешь Сириян до истребления их.
1KGS|22|12|И все пророки пророчествовали то же, говоря: иди на Рамоф Галаадский, будет успех, Господь предаст [его] в руку царя.
1KGS|22|13|Посланный, который пошел позвать Михея, говорил ему: вот, речи пророков единогласно [предвещают] царю доброе; пусть бы и твое слово было согласно с словом каждого из них; изреки и ты доброе.
1KGS|22|14|И сказал Михей: жив Господь! я изреку то, что скажет мне Господь.
1KGS|22|15|И пришел он к царю. Царь сказал ему: Михей! идти ли нам войною на Рамоф Галаадский, или нет? И сказал тот ему: иди, будет успех, Господь предаст [его] в руку царя.
1KGS|22|16|И сказал ему царь: еще и еще заклинаю тебя, чтобы ты не говорил мне ничего, кроме истины во имя Господа.
1KGS|22|17|И сказал он: я вижу всех Израильтян, рассеянных по горам, как овец, у которых нет пастыря. И сказал Господь: нет у них начальника, пусть возвращаются с миром каждый в свой дом.
1KGS|22|18|И сказал царь Израильский Иосафату: не говорил ли я тебе, что он не пророчествует о мне доброго, а только худое?
1KGS|22|19|И сказал [Михей]: выслушай слово Господне: я видел Господа, сидящего на престоле Своем, и все воинство небесное стояло при Нем, по правую и по левую руку Его;
1KGS|22|20|и сказал Господь: кто склонил бы Ахава, чтобы он пошел и пал в Рамофе Галаадском? И один говорил так, другой говорил иначе;
1KGS|22|21|и выступил один дух, стал пред лицем Господа и сказал: я склоню его. И сказал ему Господь: чем?
1KGS|22|22|Он сказал: я выйду и сделаюсь духом лживым в устах всех пророков его. [Господь] сказал: ты склонишь его и выполнишь это; пойди и сделай так.
1KGS|22|23|И вот, теперь попустил Господь духа лживого в уста всех сих пророков твоих; но Господь изрек о тебе недоброе.
1KGS|22|24|И подошел Седекия, сын Хенааны, и, ударив Михея по щеке, сказал: как, неужели от меня отошел Дух Господень, чтобы говорить в тебе?
1KGS|22|25|И сказал Михей: вот, ты увидишь [это] в тот день, когда будешь бегать из одной комнаты в другую, чтоб укрыться,
1KGS|22|26|и сказал царь Израильский: возьмите Михея и отведите его к Амону градоначальнику и к Иоасу, сыну царя,
1KGS|22|27|и скажите: так говорит царь: посадите этого в темницу и кормите его скудно хлебом и скудно водою, доколе я не возвращусь в мире.
1KGS|22|28|И сказал Михей: если возвратишься в мире, то не Господь говорил чрез меня. И сказал: слушай, весь народ!
1KGS|22|29|И пошел царь Израильский и Иосафат, царь Иудейский, к Рамофу Галаадскому.
1KGS|22|30|И сказал царь Израильский Иосафату: я переоденусь и вступлю в сражение, а ты надень твои [царские] одежды. И переоделся царь Израильский и вступил в сражение.
1KGS|22|31|Сирийский царь повелел начальникам колесниц, которых у него было тридцать два, сказав: не сражайтесь ни с малым, ни с великим, а только с одним царем Израильским.
1KGS|22|32|Начальники колесниц, увидев Иосафата, подумали: "верно это царь Израильский", и поворотили на него, чтобы сразиться [с ним]. И закричал Иосафат.
1KGS|22|33|Начальники колесниц, видя, что это не Израильский царь, поворотили от него.
1KGS|22|34|А один человек случайно натянул лук и ранил царя Израильского сквозь швы лат. И сказал он своему вознице: повороти назад и вывези меня из войска, ибо я ранен.
1KGS|22|35|Но сражение в тот день усилилось, и царь стоял на колеснице против Сириян, и вечером умер, и кровь из раны лилась в колесницу.
1KGS|22|36|И провозглашено было по всему стану при захождении солнца: каждый иди в свой город, каждый в свою землю!
1KGS|22|37|И умер царь, и привезен был в Самарию, и похоронили царя в Самарии.
1KGS|22|38|И обмыли колесницу на пруде Самарийском, и псы лизали кровь его, и омывали блудницы, по слову Господа, которое Он изрек.
1KGS|22|39|Прочие дела Ахава, все, что он делал, и дом из слоновой кости, который он построил, и все города, которые он строил, описаны в летописи царей Израильских.
1KGS|22|40|И почил Ахав с отцами своими, и воцарился Охозия, сын его, вместо него.
1KGS|22|41|Иосафат, сын Асы, воцарился над Иудеею в четвертый год Ахава, царя Израильского.
1KGS|22|42|Тридцати пяти лет был Иосафат, когда воцарился, и двадцать пять лет царствовал в Иерусалиме. Имя матери его Азува, дочь Салаиля.
1KGS|22|43|Он ходил во всем путем отца своего Асы, не сходил с него, делая угодное пред очами Господними.
1KGS|22|44|Только высоты не были отменены; народ еще совершал жертвы и курения на высотах.
1KGS|22|45|Иосафат заключил мир с царем Израильским.
1KGS|22|46|Прочие дела Иосафата и подвиги его, какие он совершил, и как он воевал, описаны в летописи царей Иудейских.
1KGS|22|47|И остатки блудников, которые остались во дни отца его Асы, он истребил с земли.
1KGS|22|48|В Идумее тогда не было царя; [был] наместник царский.
1KGS|22|49|Иосафат сделал корабли на море, чтобы ходить в Офир за золотом; но они не дошли, ибо разбились в Ецион–Гавере.
1KGS|22|50|Тогда сказал Охозия, сын Ахава, Иосафату: пусть мои слуги пойдут с твоими слугами на кораблях. Но Иосафат не согласился.
1KGS|22|51|И почил Иосафат с отцами своими и был погребен с отцами своими в городе Давида, отца своего. И воцарился Иорам, сын его, вместо него.
1KGS|22|52|Охозия, сын Ахава, воцарился над Израилем в Самарии, в семнадцатый год Иосафата, царя Иудейского, и царствовал над Израилем два года,
1KGS|22|53|и делал неугодное пред очами Господа, и ходил путем отца своего и путем матери своей и путем Иеровоама, сына Наватова, который ввел Израиля в грех:
1KGS|22|54|он служил Ваалу и поклонялся ему и прогневал Господа Бога Израилева всем тем, что делал отец его.
