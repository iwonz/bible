RUTH|1|1|士师统治的时候，国中有饥荒。在 犹大 的 伯利恒 ，有一个人带着妻子和两个儿子往 摩押 地去寄居。
RUTH|1|2|这人名叫 以利米勒 ，他的妻子名叫 拿娥米 ；他两个儿子，一个名叫 玛伦 ，一个名叫 基连 ，都是 犹大伯利恒 的 以法他 人。他们到了 摩押 地，就住在那里。
RUTH|1|3|后来 拿娥米 的丈夫 以利米勒 死了，剩下她和两个儿子。
RUTH|1|4|两个儿子娶了 摩押 女子，一个名叫 俄珥巴 ，第二个名叫 路得 ，在那里住了约有十年。
RUTH|1|5|玛伦 和 基连 二人也死了，剩下 拿娥米 ，没有丈夫，也没有儿子。
RUTH|1|6|拿娥米 与两个媳妇起身，要从 摩押 地回去，因为她在 摩押 地听见耶和华眷顾自己的百姓，赐粮食给他们。
RUTH|1|7|她和两个媳妇就起行，离开所住的地方，上路回 犹大 地去。
RUTH|1|8|拿娥米 对两个媳妇说：“你们各自回娘家去吧！愿耶和华恩待你们，像你们待已故的人和我一样。
RUTH|1|9|愿耶和华使你们各自在新的丈夫家中得归宿！”于是 拿娥米 与她们亲吻，她们就放声大哭，
RUTH|1|10|对她说：“不，我们要与你一同回你的百姓那里去。”
RUTH|1|11|拿娥米 说：“我的女儿啊，回去吧！为何要跟我去呢？我还能生儿子作你们的丈夫吗？
RUTH|1|12|我的女儿啊，回去吧！我年纪老了，不能再有丈夫。就算我还有希望，今夜有丈夫，而且也生了儿子，
RUTH|1|13|你们岂能等着他们长大呢？你们能守住自己不嫁人吗？我的女儿啊，不要这样。我比你们更苦，因为耶和华伸手击打我。”
RUTH|1|14|两个媳妇又放声大哭， 俄珥巴 与婆婆吻别，但是 路得 却紧跟着 拿娥米 。
RUTH|1|15|拿娥米 说：“看哪，你嫂嫂已经回她的百姓和她的神明那里去了，你也跟你嫂嫂回去吧！”
RUTH|1|16|路得 说： “不要劝我离开你， 转去不跟随你。 你往哪里去， 我也往哪里去； 你在哪里住， 我也在哪里住； 你的百姓就是我的百姓； 你的上帝就是我的上帝。
RUTH|1|17|你死在哪里， 我也死在哪里，葬在哪里。 只有死能使你我分离； 不然，愿耶和华重重惩罚我！”
RUTH|1|18|拿娥米 见 路得 决意要跟自己去，就不再对她说什么了。
RUTH|1|19|于是二人同行，来到 伯利恒 。她们到了 伯利恒 ，全城因她们骚动起来。妇女们说：“这是 拿娥米 吗？”
RUTH|1|20|拿娥米 对她们说： “不要叫我 拿娥米 ， 要叫我 玛拉 ， 因为全能者使我受尽了苦。
RUTH|1|21|我满满地出去， 耶和华使我空空地回来。 耶和华使我受苦， 全能者降祸于我。 你们为何还叫我 拿娥米 呢？”
RUTH|1|22|拿娥米 从 摩押 地回来了，她的媳妇 摩押 女子 路得 跟她在一起。她们到了 伯利恒 ，正是开始收割大麦的时候。
RUTH|2|1|拿娥米 有一个亲戚，是她丈夫 以利米勒 本族的人，名叫 波阿斯 ，是个大财主。
RUTH|2|2|摩押 女子 路得 对 拿娥米 说：“让我到田里去拾取麦穗，我在谁的眼中蒙恩，就跟在谁的身后。” 拿娥米 说：“女儿啊，你去吧。”
RUTH|2|3|路得 就去了。她来到田间，在收割的人身后拾取麦穗。她恰巧来到 以利米勒 本族的人 波阿斯 那块田里。
RUTH|2|4|看哪， 波阿斯 正从 伯利恒 来，对收割的人说：“愿耶和华与你们同在！”他们对他说：“愿耶和华赐福给你！”
RUTH|2|5|波阿斯 对监督收割的仆人说：“那是谁家的女子？”
RUTH|2|6|监督收割的仆人回答说：“她是 摩押 女子，跟随 拿娥米 从 摩押 地回来的。
RUTH|2|7|她说：‘请你容许我拾取麦穗，在收割的人身后捡禾捆中掉落的麦穗。’她就来了，从早晨直到如今，除了在屋子里坐一会儿，她都留在这里。”
RUTH|2|8|波阿斯 对 路得 说：“女儿啊，听我说，不要到别人田里去拾取麦穗，也不要离开这里，要紧跟着我的女仆们。
RUTH|2|9|你要看好我的仆人正在哪块田收割，就跟着女仆们去。我已经吩咐仆人不可侵犯你。你渴了，可以到水缸那里喝仆人打来的水。”　
RUTH|2|10|路得 就脸伏于地叩拜，对他说：“我既是外邦女子，怎么会在你眼中蒙恩，使你这样照顾我呢？”
RUTH|2|11|波阿斯 回答她说：“自从你丈夫死后，凡你向婆婆所行的，以及你离开父母和你的出生地，到素不相识的百姓中，这些事人都告诉我了。
RUTH|2|12|愿耶和华照你所行的报偿你。你来投靠在耶和华－ 以色列 上帝的翅膀下，愿你满得他的报偿。”
RUTH|2|13|路得 说：“我主啊，愿我在你眼前蒙恩。我虽然不及你的一个婢女，你还安慰我，对你的婢女说关心的话。”
RUTH|2|14|吃饭的时候， 波阿斯 对 路得 说：“你到这里来吃些饼，把你的一块蘸在醋里。” 路得 就在收割的人旁边坐下。 波阿斯 把烘了的穗子递给她。她吃饱了，还有剩余的。
RUTH|2|15|她又起来拾取麦穗， 波阿斯 吩咐仆人说：“她即使在禾捆中拾取麦穗，也不可羞辱她。
RUTH|2|16|你们还要从捆里抽一些出来，留给她拾取，不可责备她。”
RUTH|2|17|这样， 路得 在田间拾取麦穗，直到晚上。她把所拾取的麦穗打了约有一伊法的大麦。
RUTH|2|18|路得 把所拾取的带进城去给婆婆看，又把她吃饱所剩的拿出来，给了婆婆。
RUTH|2|19|婆婆问她说：“你今日在哪里拾取麦穗？在哪里做工呢？愿那照顾你的得福。” 路得 告诉婆婆，她在谁那里做工，说：“我今日在一个名叫 波阿斯 的人那里做工。”
RUTH|2|20|拿娥米 对媳妇说：“愿那人蒙耶和华赐福，因为他不断地恩待活人死人。” 拿娥米 又对她说：“那人是我们本族的人，是一个可以赎我们产业的至亲。”
RUTH|2|21|摩押 女子 路得 说：“他还对我说：‘你要紧跟着我的仆人拾取麦穗，直到他们把我所有的庄稼收割完毕。’”
RUTH|2|22|拿娥米 对媳妇 路得 说：“女儿啊，你要跟着他的女仆出去，免得你在别人的田间受人骚扰。”
RUTH|2|23|于是 路得 紧跟着 波阿斯 的女仆拾取麦穗，直到大麦和小麦收割完毕。 路得 仍与婆婆同住。
RUTH|3|1|路得 的婆婆 拿娥米 对她说：“女儿啊，我不该为你找个归宿，使你享福吗？
RUTH|3|2|你与 波阿斯 的女仆常在一处，现在， 波阿斯 不是我们的亲人吗？看哪，他今夜将在禾场簸大麦。
RUTH|3|3|你要沐浴抹膏，穿上外衣，下到禾场，一直到那人吃喝完了，都不要让他认出你来。
RUTH|3|4|他躺下的时候，你看准他躺卧的地方，就进去掀露他的脚，躺卧在那里，他必告诉你所当做的事。”
RUTH|3|5|路得 说：“凡你所吩咐我的，我必遵行。”
RUTH|3|6|路得 就下到禾场，照她婆婆吩咐她的一切去做。
RUTH|3|7|波阿斯 吃喝完了，心情畅快，就去躺卧在麦堆旁边。 路得 悄悄走来，掀露他的脚，躺卧在那里。
RUTH|3|8|到了半夜，那人惊醒，翻过身来，看哪，有个女子躺在他的脚旁。
RUTH|3|9|他就说：“你是谁？” 路得 说：“我是你的使女 路得 。请你用你衣服的边来遮盖你的使女，因为你是可以赎我产业的至亲。”
RUTH|3|10|波阿斯 说：“女儿啊，愿你蒙耶和华赐福。你后来的忠诚比先前的更美，因为无论贫富的年轻人，你都没有跟从。
RUTH|3|11|女儿啊，现在不要惧怕，凡你所说的，我必为你做，因为我城里的百姓都知道你是个贤德的女子。
RUTH|3|12|现在，我的确是一个可以赎你产业的至亲，可是还有一个人比我更亲。
RUTH|3|13|你今夜在这里住宿，明早他若肯为你尽至亲的本分，很好，就由他吧！倘若他不肯，我指着永生的耶和华起誓，我必为你尽上至亲的本分。你只管躺到早晨。”
RUTH|3|14|路得 就在他脚旁躺到早晨，在人还无法彼此辨认的时候就起来了。 波阿斯 说：“不可让人知道有女子到禾场来。”　
RUTH|3|15|他又对 路得 说：“把你所披的外衣拿来，握紧它。”她就握紧外衣， 波阿斯 量了六簸箕的大麦，帮 路得 扛上，他就进城去了 。”
RUTH|3|16|路得 回到婆婆那里，婆婆说：“女儿啊，怎么样了 ？” 路得 就把那人向她所做的一切都告诉了婆婆，
RUTH|3|17|又说：“那人给了我这六簸箕的大麦，对我说：‘你不可空手回去见婆婆。’”
RUTH|3|18|婆婆说：“女儿啊，等着吧，看这事结果如何，因为那人今日不办妥这事，必不罢休。”
RUTH|4|1|波阿斯 上到城门，坐在那里，看哪， 波阿斯 所说那个可以赎产业的至亲经过。 波阿斯 说：“某某先生，请你转回来，坐在这里。”他就转回来坐下。
RUTH|4|2|波阿斯 又请了本城的十个长老来，对他们说：“请你们坐在这里。”他们就都坐下。
RUTH|4|3|波阿斯 对那至亲说：“从 摩押 地回来的 拿娥米 ，现在要卖我们弟兄 以利米勒 的那块地。
RUTH|4|4|我想我应该向你说清楚：你可以买那块地，当着在座的众人和我百姓的长老面前，你若要赎就赎吧！倘若你不赎 就告诉我，让我知道，因为除了你以外，没有人可以先赎，在你之后才轮到我。”那人说：“我要赎。”
RUTH|4|5|波阿斯 说：“你从 拿娥米 和 摩押 女子 路得 手中买这地的时候，也当买死人的妻子，使死人在产业上留名。”
RUTH|4|6|那至亲说：“这样我就不能赎了，免得对我的产业有损。你尽管去赎我所当赎的吧，我不能赎了！”
RUTH|4|7|从前，在 以色列 中要确认任何交易，无论是赎业或买卖，一方必须脱鞋给另一方。 以色列 中都以此为证。
RUTH|4|8|那至亲对 波阿斯 说：“你自己买吧！”于是把鞋脱了下来。
RUTH|4|9|波阿斯 对长老和所有在场的百姓说：“你们今日都是证人；凡属 以利米勒 ，以及 基连 和 玛伦 的，我都从 拿娥米 手中买下来了。
RUTH|4|10|我也娶 玛伦 的妻子 摩押 女子 路得 ，好让死人可以在产业上留名，免得他的名在本族本乡的城门中消失了。你们今日都是证人。”
RUTH|4|11|在城门坐着的所有百姓和长老说：“我们都是证人。愿耶和华使进你家的这女子，像建立 以色列 家的 拉结 和 利亚 二人一样。又愿你在 以法他 得亨通，在 伯利恒 有名声。
RUTH|4|12|愿耶和华从这年轻女子赐你后裔，使你的家像 她玛 从 犹大 所生 法勒斯 的家一样。”
RUTH|4|13|于是， 波阿斯 娶了 路得 为妻，与她同房。耶和华使她怀孕生了一个儿子。
RUTH|4|14|妇女们对 拿娥米 说：“耶和华是应当称颂的！因为他今日没有使你断绝可以赎产业的至亲。愿这孩子在 以色列 中得名声。
RUTH|4|15|他必振奋你的精神，奉养你的晚年，因为他是爱慕你的媳妇所生的。有这样的媳妇，比有七个儿子更好！”
RUTH|4|16|拿娥米 接过孩子来，抱在怀中抚养他。
RUTH|4|17|邻居的妇人给孩子起名，说：“ 拿娥米 得了一个孩子了！”她们就给他起名叫 俄备得 。 俄备得 是 耶西 的父亲，是 大卫 的祖父。
RUTH|4|18|这是 法勒斯 的后代： 法勒斯 生 希斯仑 ；
RUTH|4|19|希斯仑 生 兰 ； 兰 生 亚米拿达 ；
RUTH|4|20|亚米拿达 生 拿顺 ； 拿顺 生 撒门 ；
RUTH|4|21|撒门 生 波阿斯 ； 波阿斯 生 俄备得 ；
RUTH|4|22|俄备得 生 耶西 ； 耶西 生 大卫 。
