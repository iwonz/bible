1CHR|1|1|Adam, Seth, Enosh,
1CHR|1|2|Kenan, Mahalalel, Jared,
1CHR|1|3|Enoch, Methuselah, Lamech, Noah.
1CHR|1|4|The sons of Noah: Shem, Ham and Japheth. The Japhethites
1CHR|1|5|The sons of Japheth: Gomer, Magog, Madai, Javan, Tubal, Meshech and Tiras.
1CHR|1|6|The sons of Gomer: Ashkenaz, Riphath and Togarmah.
1CHR|1|7|The sons of Javan: Elishah, Tarshish, the Kittim and the Rodanim. The Hamites
1CHR|1|8|The sons of Ham: Cush, Mizraim, Put and Canaan.
1CHR|1|9|The sons of Cush: Seba, Havilah, Sabta, Raamah and Sabteca. The sons of Raamah: Sheba and Dedan.
1CHR|1|10|Cush was the father of Nimrod, who grew to be a mighty warrior on earth.
1CHR|1|11|Mizraim was the father of the Ludites, Anamites, Lehabites, Naphtuhites,
1CHR|1|12|Pathrusites, Casluhites (from whom the Philistines came) and Caphtorites.
1CHR|1|13|Canaan was the father of Sidon his firstborn, and of the Hittites,
1CHR|1|14|Jebusites, Amorites, Girgashites,
1CHR|1|15|Hivites, Arkites, Sinites,
1CHR|1|16|Arvadites, Zemarites and Hamathites. The Semites
1CHR|1|17|The sons of Shem: Elam, Asshur, Arphaxad, Lud and Aram. The sons of Aram: Uz, Hul, Gether and Meshech.
1CHR|1|18|Arphaxad was the father of Shelah, and Shelah the father of Eber.
1CHR|1|19|Two sons were born to Eber: One was named Peleg, because in his time the earth was divided; his brother was named Joktan.
1CHR|1|20|Joktan was the father of Almodad, Sheleph, Hazarmaveth, Jerah,
1CHR|1|21|Hadoram, Uzal, Diklah,
1CHR|1|22|Obal, Abimael, Sheba,
1CHR|1|23|Ophir, Havilah and Jobab. All these were sons of Joktan.
1CHR|1|24|Shem, Arphaxad, Shelah,
1CHR|1|25|Eber, Peleg, Reu,
1CHR|1|26|Serug, Nahor, Terah
1CHR|1|27|and Abram (that is, Abraham).
1CHR|1|28|The sons of Abraham: Isaac and Ishmael. Descendants of Hagar
1CHR|1|29|These were their descendants: Nebaioth the firstborn of Ishmael, Kedar, Adbeel, Mibsam,
1CHR|1|30|Mishma, Dumah, Massa, Hadad, Tema,
1CHR|1|31|Jetur, Naphish and Kedemah. These were the sons of Ishmael. Descendants of Keturah
1CHR|1|32|The sons born to Keturah, Abraham's concubine: Zimran, Jokshan, Medan, Midian, Ishbak and Shuah. The sons of Jokshan: Sheba and Dedan.
1CHR|1|33|The sons of Midian: Ephah, Epher, Hanoch, Abida and Eldaah. All these were descendants of Keturah. Descendants of Sarah
1CHR|1|34|Abraham was the father of Isaac. The sons of Isaac: Esau and Israel.
1CHR|1|35|The sons of Esau: Eliphaz, Reuel, Jeush, Jalam and Korah.
1CHR|1|36|The sons of Eliphaz: Teman, Omar, Zepho, Gatam and Kenaz; by Timna: Amalek.
1CHR|1|37|The sons of Reuel: Nahath, Zerah, Shammah and Mizzah. The People of Seir in Edom
1CHR|1|38|The sons of Seir: Lotan, Shobal, Zibeon, Anah, Dishon, Ezer and Dishan.
1CHR|1|39|The sons of Lotan: Hori and Homam. Timna was Lotan's sister.
1CHR|1|40|The sons of Shobal: Alvan, Manahath, Ebal, Shepho and Onam. The sons of Zibeon: Aiah and Anah.
1CHR|1|41|The son of Anah: Dishon. The sons of Dishon: Hemdan, Eshban, Ithran and Keran.
1CHR|1|42|The sons of Ezer: Bilhan, Zaavan and Akan. The sons of Dishan: Uz and Aran. The Rulers of Edom
1CHR|1|43|These were the kings who reigned in Edom before any Israelite king reigned: Bela son of Beor, whose city was named Dinhabah.
1CHR|1|44|When Bela died, Jobab son of Zerah from Bozrah succeeded him as king.
1CHR|1|45|When Jobab died, Husham from the land of the Temanites succeeded him as king.
1CHR|1|46|When Husham died, Hadad son of Bedad, who defeated Midian in the country of Moab, succeeded him as king. His city was named Avith.
1CHR|1|47|When Hadad died, Samlah from Masrekah succeeded him as king.
1CHR|1|48|When Samlah died, Shaul from Rehoboth on the river succeeded him as king.
1CHR|1|49|When Shaul died, Baal-Hanan son of Acbor succeeded him as king.
1CHR|1|50|When Baal-Hanan died, Hadad succeeded him as king. His city was named Pau, and his wife's name was Mehetabel daughter of Matred, the daughter of Me-Zahab.
1CHR|1|51|Hadad also died. The chiefs of Edom were: Timna, Alvah, Jetheth,
1CHR|1|52|Oholibamah, Elah, Pinon,
1CHR|1|53|Kenaz, Teman, Mibzar,
1CHR|1|54|Magdiel and Iram. These were the chiefs of Edom.
1CHR|2|1|These were the sons of Israel: Reuben, Simeon, Levi, Judah, Issachar, Zebulun,
1CHR|2|2|Dan, Joseph, Benjamin, Naphtali, Gad and Asher.
1CHR|2|3|The sons of Judah: Er, Onan and Shelah. These three were born to him by a Canaanite woman, the daughter of Shua. Er, Judah's firstborn, was wicked in the LORD's sight; so the LORD put him to death.
1CHR|2|4|Tamar, Judah's daughter-in-law, bore him Perez and Zerah. Judah had five sons in all.
1CHR|2|5|The sons of Perez: Hezron and Hamul.
1CHR|2|6|The sons of Zerah: Zimri, Ethan, Heman, Calcol and Darda -five in all.
1CHR|2|7|The son of Carmi: Achar, who brought trouble on Israel by violating the ban on taking devoted things.
1CHR|2|8|The son of Ethan: Azariah.
1CHR|2|9|The sons born to Hezron were: Jerahmeel, Ram and Caleb. From Ram Son of Hezron
1CHR|2|10|Ram was the father of Amminadab, and Amminadab the father of Nahshon, the leader of the people of Judah.
1CHR|2|11|Nahshon was the father of Salmon, Salmon the father of Boaz,
1CHR|2|12|Boaz the father of Obed and Obed the father of Jesse.
1CHR|2|13|Jesse was the father of Eliab his firstborn; the second son was Abinadab, the third Shimea,
1CHR|2|14|the fourth Nethanel, the fifth Raddai,
1CHR|2|15|the sixth Ozem and the seventh David.
1CHR|2|16|Their sisters were Zeruiah and Abigail. Zeruiah's three sons were Abishai, Joab and Asahel.
1CHR|2|17|Abigail was the mother of Amasa, whose father was Jether the Ishmaelite. Caleb Son of Hezron
1CHR|2|18|Caleb son of Hezron had children by his wife Azubah (and by Jerioth). These were her sons: Jesher, Shobab and Ardon.
1CHR|2|19|When Azubah died, Caleb married Ephrath, who bore him Hur.
1CHR|2|20|Hur was the father of Uri, and Uri the father of Bezalel.
1CHR|2|21|Later, Hezron lay with the daughter of Makir the father of Gilead (he had married her when he was sixty years old), and she bore him Segub.
1CHR|2|22|Segub was the father of Jair, who controlled twenty-three towns in Gilead.
1CHR|2|23|(But Geshur and Aram captured Havvoth Jair, as well as Kenath with its surrounding settlements-sixty towns.) All these were descendants of Makir the father of Gilead.
1CHR|2|24|After Hezron died in Caleb Ephrathah, Abijah the wife of Hezron bore him Ashhur the father of Tekoa. Jerahmeel Son of Hezron
1CHR|2|25|The sons of Jerahmeel the firstborn of Hezron: Ram his firstborn, Bunah, Oren, Ozem and Ahijah.
1CHR|2|26|Jerahmeel had another wife, whose name was Atarah; she was the mother of Onam.
1CHR|2|27|The sons of Ram the firstborn of Jerahmeel: Maaz, Jamin and Eker.
1CHR|2|28|The sons of Onam: Shammai and Jada. The sons of Shammai: Nadab and Abishur.
1CHR|2|29|Abishur's wife was named Abihail, who bore him Ahban and Molid.
1CHR|2|30|The sons of Nadab: Seled and Appaim. Seled died without children.
1CHR|2|31|The son of Appaim: Ishi, who was the father of Sheshan. Sheshan was the father of Ahlai.
1CHR|2|32|The sons of Jada, Shammai's brother: Jether and Jonathan. Jether died without children.
1CHR|2|33|The sons of Jonathan: Peleth and Zaza. These were the descendants of Jerahmeel.
1CHR|2|34|Sheshan had no sons-only daughters. He had an Egyptian servant named Jarha.
1CHR|2|35|Sheshan gave his daughter in marriage to his servant Jarha, and she bore him Attai.
1CHR|2|36|Attai was the father of Nathan, Nathan the father of Zabad,
1CHR|2|37|Zabad the father of Ephlal, Ephlal the father of Obed,
1CHR|2|38|Obed the father of Jehu, Jehu the father of Azariah,
1CHR|2|39|Azariah the father of Helez, Helez the father of Eleasah,
1CHR|2|40|Eleasah the father of Sismai, Sismai the father of Shallum,
1CHR|2|41|Shallum the father of Jekamiah, and Jekamiah the father of Elishama. The Clans of Caleb
1CHR|2|42|The sons of Caleb the brother of Jerahmeel: Mesha his firstborn, who was the father of Ziph, and his son Mareshah, who was the father of Hebron.
1CHR|2|43|The sons of Hebron: Korah, Tappuah, Rekem and Shema.
1CHR|2|44|Shema was the father of Raham, and Raham the father of Jorkeam. Rekem was the father of Shammai.
1CHR|2|45|The son of Shammai was Maon, and Maon was the father of Beth Zur.
1CHR|2|46|Caleb's concubine Ephah was the mother of Haran, Moza and Gazez. Haran was the father of Gazez.
1CHR|2|47|The sons of Jahdai: Regem, Jotham, Geshan, Pelet, Ephah and Shaaph.
1CHR|2|48|Caleb's concubine Maacah was the mother of Sheber and Tirhanah.
1CHR|2|49|She also gave birth to Shaaph the father of Madmannah and to Sheva the father of Macbenah and Gibea. Caleb's daughter was Acsah.
1CHR|2|50|These were the descendants of Caleb. The sons of Hur the firstborn of Ephrathah: Shobal the father of Kiriath Jearim,
1CHR|2|51|Salma the father of Bethlehem, and Hareph the father of Beth Gader.
1CHR|2|52|The descendants of Shobal the father of Kiriath Jearim were: Haroeh, half the Manahathites,
1CHR|2|53|and the clans of Kiriath Jearim: the Ithrites, Puthites, Shumathites and Mishraites. From these descended the Zorathites and Eshtaolites.
1CHR|2|54|The descendants of Salma: Bethlehem, the Netophathites, Atroth Beth Joab, half the Manahathites, the Zorites,
1CHR|2|55|and the clans of scribes who lived at Jabez: the Tirathites, Shimeathites and Sucathites. These are the Kenites who came from Hammath, the father of the house of Recab.
1CHR|3|1|These were the sons of David born to him in Hebron: The firstborn was Amnon the son of Ahinoam of Jezreel; the second, Daniel the son of Abigail of Carmel;
1CHR|3|2|the third, Absalom the son of Maacah daughter of Talmai king of Geshur; the fourth, Adonijah the son of Haggith;
1CHR|3|3|the fifth, Shephatiah the son of Abital; and the sixth, Ithream, by his wife Eglah.
1CHR|3|4|These six were born to David in Hebron, where he reigned seven years and six months. David reigned in Jerusalem thirty-three years,
1CHR|3|5|and these were the children born to him there: Shammua, Shobab, Nathan and Solomon. These four were by Bathsheba daughter of Ammiel.
1CHR|3|6|There were also Ibhar, Elishua, Eliphelet,
1CHR|3|7|Nogah, Nepheg, Japhia,
1CHR|3|8|Elishama, Eliada and Eliphelet-nine in all.
1CHR|3|9|All these were the sons of David, besides his sons by his concubines. And Tamar was their sister. The Kings of Judah
1CHR|3|10|Solomon's son was Rehoboam, Abijah his son, Asa his son, Jehoshaphat his son,
1CHR|3|11|Jehoram his son, Ahaziah his son, Joash his son,
1CHR|3|12|Amaziah his son, Azariah his son, Jotham his son,
1CHR|3|13|Ahaz his son, Hezekiah his son, Manasseh his son,
1CHR|3|14|Amon his son, Josiah his son.
1CHR|3|15|The sons of Josiah: Johanan the firstborn, Jehoiakim the second son, Zedekiah the third, Shallum the fourth.
1CHR|3|16|The successors of Jehoiakim: Jehoiachin his son, and Zedekiah. The Royal Line After the Exile
1CHR|3|17|The descendants of Jehoiachin the captive: Shealtiel his son,
1CHR|3|18|Malkiram, Pedaiah, Shenazzar, Jekamiah, Hoshama and Nedabiah.
1CHR|3|19|The sons of Pedaiah: Zerubbabel and Shimei. The sons of Zerubbabel: Meshullam and Hananiah. Shelomith was their sister.
1CHR|3|20|There were also five others: Hashubah, Ohel, Berekiah, Hasadiah and Jushab-Hesed.
1CHR|3|21|The descendants of Hananiah: Pelatiah and Jeshaiah, and the sons of Rephaiah, of Arnan, of Obadiah and of Shecaniah.
1CHR|3|22|The descendants of Shecaniah: Shemaiah and his sons: Hattush, Igal, Bariah, Neariah and Shaphat-six in all.
1CHR|3|23|The sons of Neariah: Elioenai, Hizkiah and Azrikam-three in all.
1CHR|3|24|The sons of Elioenai: Hodaviah, Eliashib, Pelaiah, Akkub, Johanan, Delaiah and Anani-seven in all.
1CHR|4|1|The descendants of Judah: Perez, Hezron, Carmi, Hur and Shobal.
1CHR|4|2|Reaiah son of Shobal was the father of Jahath, and Jahath the father of Ahumai and Lahad. These were the clans of the Zorathites.
1CHR|4|3|These were the sons of Etam: Jezreel, Ishma and Idbash. Their sister was named Hazzelelponi.
1CHR|4|4|Penuel was the father of Gedor, and Ezer the father of Hushah. These were the descendants of Hur, the firstborn of Ephrathah and father of Bethlehem.
1CHR|4|5|Ashhur the father of Tekoa had two wives, Helah and Naarah.
1CHR|4|6|Naarah bore him Ahuzzam, Hepher, Temeni and Haahashtari. These were the descendants of Naarah.
1CHR|4|7|The sons of Helah: Zereth, Zohar, Ethnan,
1CHR|4|8|and Koz, who was the father of Anub and Hazzobebah and of the clans of Aharhel son of Harum.
1CHR|4|9|Jabez was more honorable than his brothers. His mother had named him Jabez, saying, "I gave birth to him in pain."
1CHR|4|10|Jabez cried out to the God of Israel, "Oh, that you would bless me and enlarge my territory! Let your hand be with me, and keep me from harm so that I will be free from pain." And God granted his request.
1CHR|4|11|Kelub, Shuhah's brother, was the father of Mehir, who was the father of Eshton.
1CHR|4|12|Eshton was the father of Beth Rapha, Paseah and Tehinnah the father of Ir Nahash. These were the men of Recah.
1CHR|4|13|The sons of Kenaz: Othniel and Seraiah. The sons of Othniel: Hathath and Meonothai.
1CHR|4|14|Meonothai was the father of Ophrah. Seraiah was the father of Joab, the father of Ge Harashim. It was called this because its people were craftsmen.
1CHR|4|15|The sons of Caleb son of Jephunneh: Iru, Elah and Naam. The son of Elah: Kenaz.
1CHR|4|16|The sons of Jehallelel: Ziph, Ziphah, Tiria and Asarel.
1CHR|4|17|The sons of Ezrah: Jether, Mered, Epher and Jalon. One of Mered's wives gave birth to Miriam, Shammai and Ishbah the father of Eshtemoa.
1CHR|4|18|(His Judean wife gave birth to Jered the father of Gedor, Heber the father of Soco, and Jekuthiel the father of Zanoah.) These were the children of Pharaoh's daughter Bithiah, whom Mered had married.
1CHR|4|19|The sons of Hodiah's wife, the sister of Naham: the father of Keilah the Garmite, and Eshtemoa the Maacathite.
1CHR|4|20|The sons of Shimon: Amnon, Rinnah, Ben-Hanan and Tilon. The descendants of Ishi: Zoheth and Ben-Zoheth.
1CHR|4|21|The sons of Shelah son of Judah: Er the father of Lecah, Laadah the father of Mareshah and the clans of the linen workers at Beth Ashbea,
1CHR|4|22|Jokim, the men of Cozeba, and Joash and Saraph, who ruled in Moab and Jashubi Lehem. (These records are from ancient times.)
1CHR|4|23|They were the potters who lived at Netaim and Gederah; they stayed there and worked for the king.
1CHR|4|24|The descendants of Simeon: Nemuel, Jamin, Jarib, Zerah and Shaul;
1CHR|4|25|Shallum was Shaul's son, Mibsam his son and Mishma his son.
1CHR|4|26|The descendants of Mishma: Hammuel his son, Zaccur his son and Shimei his son.
1CHR|4|27|Shimei had sixteen sons and six daughters, but his brothers did not have many children; so their entire clan did not become as numerous as the people of Judah.
1CHR|4|28|They lived in Beersheba, Moladah, Hazar Shual,
1CHR|4|29|Bilhah, Ezem, Tolad,
1CHR|4|30|Bethuel, Hormah, Ziklag,
1CHR|4|31|Beth Marcaboth, Hazar Susim, Beth Biri and Shaaraim. These were their towns until the reign of David.
1CHR|4|32|Their surrounding villages were Etam, Ain, Rimmon, Token and Ashan-five towns-
1CHR|4|33|and all the villages around these towns as far as Baalath. These were their settlements. And they kept a genealogical record.
1CHR|4|34|Meshobab, Jamlech, Joshah son of Amaziah,
1CHR|4|35|Joel, Jehu son of Joshibiah, the son of Seraiah, the son of Asiel,
1CHR|4|36|also Elioenai, Jaakobah, Jeshohaiah, Asaiah, Adiel, Jesimiel, Benaiah,
1CHR|4|37|and Ziza son of Shiphi, the son of Allon, the son of Jedaiah, the son of Shimri, the son of Shemaiah.
1CHR|4|38|The men listed above by name were leaders of their clans. Their families increased greatly,
1CHR|4|39|and they went to the outskirts of Gedor to the east of the valley in search of pasture for their flocks.
1CHR|4|40|They found rich, good pasture, and the land was spacious, peaceful and quiet. Some Hamites had lived there formerly.
1CHR|4|41|The men whose names were listed came in the days of Hezekiah king of Judah. They attacked the Hamites in their dwellings and also the Meunites who were there and completely destroyed them, as is evident to this day. Then they settled in their place, because there was pasture for their flocks.
1CHR|4|42|And five hundred of these Simeonites, led by Pelatiah, Neariah, Rephaiah and Uzziel, the sons of Ishi, invaded the hill country of Seir.
1CHR|4|43|They killed the remaining Amalekites who had escaped, and they have lived there to this day.
1CHR|5|1|The sons of Reuben the firstborn of Israel (he was the firstborn, but when he defiled his father's marriage bed, his rights as firstborn were given to the sons of Joseph son of Israel; so he could not be listed in the genealogical record in accordance with his birthright,
1CHR|5|2|and though Judah was the strongest of his brothers and a ruler came from him, the rights of the firstborn belonged to Joseph)-
1CHR|5|3|the sons of Reuben the firstborn of Israel: Hanoch, Pallu, Hezron and Carmi.
1CHR|5|4|The descendants of Joel: Shemaiah his son, Gog his son, Shimei his son,
1CHR|5|5|Micah his son, Reaiah his son, Baal his son,
1CHR|5|6|and Beerah his son, whom Tiglath-Pileser king of Assyria took into exile. Beerah was a leader of the Reubenites.
1CHR|5|7|Their relatives by clans, listed according to their genealogical records: Jeiel the chief, Zechariah,
1CHR|5|8|and Bela son of Azaz, the son of Shema, the son of Joel. They settled in the area from Aroer to Nebo and Baal Meon.
1CHR|5|9|To the east they occupied the land up to the edge of the desert that extends to the Euphrates River, because their livestock had increased in Gilead.
1CHR|5|10|During Saul's reign they waged war against the Hagrites, who were defeated at their hands; they occupied the dwellings of the Hagrites throughout the entire region east of Gilead.
1CHR|5|11|The Gadites lived next to them in Bashan, as far as Salecah:
1CHR|5|12|Joel was the chief, Shapham the second, then Janai and Shaphat, in Bashan.
1CHR|5|13|Their relatives, by families, were: Michael, Meshullam, Sheba, Jorai, Jacan, Zia and Eber-seven in all.
1CHR|5|14|These were the sons of Abihail son of Huri, the son of Jaroah, the son of Gilead, the son of Michael, the son of Jeshishai, the son of Jahdo, the son of Buz.
1CHR|5|15|Ahi son of Abdiel, the son of Guni, was head of their family.
1CHR|5|16|The Gadites lived in Gilead, in Bashan and its outlying villages, and on all the pasturelands of Sharon as far as they extended.
1CHR|5|17|All these were entered in the genealogical records during the reigns of Jotham king of Judah and Jeroboam king of Israel.
1CHR|5|18|The Reubenites, the Gadites and the half-tribe of Manasseh had 44,760 men ready for military service-able-bodied men who could handle shield and sword, who could use a bow, and who were trained for battle.
1CHR|5|19|They waged war against the Hagrites, Jetur, Naphish and Nodab.
1CHR|5|20|They were helped in fighting them, and God handed the Hagrites and all their allies over to them, because they cried out to him during the battle. He answered their prayers, because they trusted in him.
1CHR|5|21|They seized the livestock of the Hagrites-fifty thousand camels, two hundred fifty thousand sheep and two thousand donkeys. They also took one hundred thousand people captive,
1CHR|5|22|and many others fell slain, because the battle was God's. And they occupied the land until the exile.
1CHR|5|23|The people of the half-tribe of Manasseh were numerous; they settled in the land from Bashan to Baal Hermon, that is, to Senir (Mount Hermon).
1CHR|5|24|These were the heads of their families: Epher, Ishi, Eliel, Azriel, Jeremiah, Hodaviah and Jahdiel. They were brave warriors, famous men, and heads of their families.
1CHR|5|25|But they were unfaithful to the God of their fathers and prostituted themselves to the gods of the peoples of the land, whom God had destroyed before them.
1CHR|5|26|So the God of Israel stirred up the spirit of Pul king of Assyria (that is, Tiglath-Pileser king of Assyria), who took the Reubenites, the Gadites and the half-tribe of Manasseh into exile. He took them to Halah, Habor, Hara and the river of Gozan, where they are to this day.
1CHR|6|1|The sons of Levi: Gershon, Kohath and Merari.
1CHR|6|2|The sons of Kohath: Amram, Izhar, Hebron and Uzziel.
1CHR|6|3|The children of Amram: Aaron, Moses and Miriam. The sons of Aaron: Nadab, Abihu, Eleazar and Ithamar.
1CHR|6|4|Eleazar was the father of Phinehas, Phinehas the father of Abishua,
1CHR|6|5|Abishua the father of Bukki, Bukki the father of Uzzi,
1CHR|6|6|Uzzi the father of Zerahiah, Zerahiah the father of Meraioth,
1CHR|6|7|Meraioth the father of Amariah, Amariah the father of Ahitub,
1CHR|6|8|Ahitub the father of Zadok, Zadok the father of Ahimaaz,
1CHR|6|9|Ahimaaz the father of Azariah, Azariah the father of Johanan,
1CHR|6|10|Johanan the father of Azariah (it was he who served as priest in the temple Solomon built in Jerusalem),
1CHR|6|11|Azariah the father of Amariah, Amariah the father of Ahitub,
1CHR|6|12|Ahitub the father of Zadok, Zadok the father of Shallum,
1CHR|6|13|Shallum the father of Hilkiah, Hilkiah the father of Azariah,
1CHR|6|14|Azariah the father of Seraiah, and Seraiah the father of Jehozadak.
1CHR|6|15|Jehozadak was deported when the LORD sent Judah and Jerusalem into exile by the hand of Nebuchadnezzar.
1CHR|6|16|The sons of Levi: Gershon, Kohath and Merari.
1CHR|6|17|These are the names of the sons of Gershon: Libni and Shimei.
1CHR|6|18|The sons of Kohath: Amram, Izhar, Hebron and Uzziel.
1CHR|6|19|The sons of Merari: Mahli and Mushi. These are the clans of the Levites listed according to their fathers:
1CHR|6|20|Of Gershon: Libni his son, Jehath his son, Zimmah his son,
1CHR|6|21|Joah his son, Iddo his son, Zerah his son and Jeatherai his son.
1CHR|6|22|The descendants of Kohath: Amminadab his son, Korah his son, Assir his son,
1CHR|6|23|Elkanah his son, Ebiasaph his son, Assir his son,
1CHR|6|24|Tahath his son, Uriel his son, Uzziah his son and Shaul his son.
1CHR|6|25|The descendants of Elkanah: Amasai, Ahimoth,
1CHR|6|26|Elkanah his son, Zophai his son, Nahath his son,
1CHR|6|27|Eliab his son, Jeroham his son, Elkanah his son and Samuel his son.
1CHR|6|28|The sons of Samuel: Joel the firstborn and Abijah the second son.
1CHR|6|29|The descendants of Merari: Mahli, Libni his son, Shimei his son, Uzzah his son,
1CHR|6|30|Shimea his son, Haggiah his son and Asaiah his son. The Temple Musicians
1CHR|6|31|These are the men David put in charge of the music in the house of the LORD after the ark came to rest there.
1CHR|6|32|They ministered with music before the tabernacle, the Tent of Meeting, until Solomon built the temple of the LORD in Jerusalem. They performed their duties according to the regulations laid down for them.
1CHR|6|33|Here are the men who served, together with their sons: From the Kohathites: Heman, the musician, the son of Joel, the son of Samuel,
1CHR|6|34|the son of Elkanah, the son of Jeroham, the son of Eliel, the son of Toah,
1CHR|6|35|the son of Zuph, the son of Elkanah, the son of Mahath, the son of Amasai,
1CHR|6|36|the son of Elkanah, the son of Joel, the son of Azariah, the son of Zephaniah,
1CHR|6|37|the son of Tahath, the son of Assir, the son of Ebiasaph, the son of Korah,
1CHR|6|38|the son of Izhar, the son of Kohath, the son of Levi, the son of Israel;
1CHR|6|39|and Heman's associate Asaph, who served at his right hand: Asaph son of Berekiah, the son of Shimea,
1CHR|6|40|the son of Michael, the son of Baaseiah, the son of Malkijah,
1CHR|6|41|the son of Ethni, the son of Zerah, the son of Adaiah,
1CHR|6|42|the son of Ethan, the son of Zimmah, the son of Shimei,
1CHR|6|43|the son of Jahath, the son of Gershon, the son of Levi;
1CHR|6|44|and from their associates, the Merarites, at his left hand: Ethan son of Kishi, the son of Abdi, the son of Malluch,
1CHR|6|45|the son of Hashabiah, the son of Amaziah, the son of Hilkiah,
1CHR|6|46|the son of Amzi, the son of Bani, the son of Shemer,
1CHR|6|47|the son of Mahli, the son of Mushi, the son of Merari, the son of Levi.
1CHR|6|48|Their fellow Levites were assigned to all the other duties of the tabernacle, the house of God.
1CHR|6|49|But Aaron and his descendants were the ones who presented offerings on the altar of burnt offering and on the altar of incense in connection with all that was done in the Most Holy Place, making atonement for Israel, in accordance with all that Moses the servant of God had commanded.
1CHR|6|50|These were the descendants of Aaron: Eleazar his son, Phinehas his son, Abishua his son,
1CHR|6|51|Bukki his son, Uzzi his son, Zerahiah his son,
1CHR|6|52|Meraioth his son, Amariah his son, Ahitub his son,
1CHR|6|53|Zadok his son and Ahimaaz his son.
1CHR|6|54|These were the locations of their settlements allotted as their territory (they were assigned to the descendants of Aaron who were from the Kohathite clan, because the first lot was for them):
1CHR|6|55|They were given Hebron in Judah with its surrounding pasturelands.
1CHR|6|56|But the fields and villages around the city were given to Caleb son of Jephunneh.
1CHR|6|57|So the descendants of Aaron were given Hebron (a city of refuge), and Libnah, Jattir, Eshtemoa,
1CHR|6|58|Hilen, Debir,
1CHR|6|59|Ashan, Juttah and Beth Shemesh, together with their pasturelands.
1CHR|6|60|And from the tribe of Benjamin they were given Gibeon, Geba, Alemeth and Anathoth, together with their pasturelands. These towns, which were distributed among the Kohathite clans, were thirteen in all.
1CHR|6|61|The rest of Kohath's descendants were allotted ten towns from the clans of half the tribe of Manasseh.
1CHR|6|62|The descendants of Gershon, clan by clan, were allotted thirteen towns from the tribes of Issachar, Asher and Naphtali, and from the part of the tribe of Manasseh that is in Bashan.
1CHR|6|63|The descendants of Merari, clan by clan, were allotted twelve towns from the tribes of Reuben, Gad and Zebulun.
1CHR|6|64|So the Israelites gave the Levites these towns and their pasturelands.
1CHR|6|65|From the tribes of Judah, Simeon and Benjamin they allotted the previously named towns.
1CHR|6|66|Some of the Kohathite clans were given as their territory towns from the tribe of Ephraim.
1CHR|6|67|In the hill country of Ephraim they were given Shechem (a city of refuge), and Gezer,
1CHR|6|68|Jokmeam, Beth Horon,
1CHR|6|69|Aijalon and Gath Rimmon, together with their pasturelands.
1CHR|6|70|And from half the tribe of Manasseh the Israelites gave Aner and Bileam, together with their pasturelands, to the rest of the Kohathite clans.
1CHR|6|71|The Gershonites received the following: From the clan of the half-tribe of Manasseh they received Golan in Bashan and also Ashtaroth, together with their pasturelands;
1CHR|6|72|from the tribe of Issachar they received Kedesh, Daberath,
1CHR|6|73|Ramoth and Anem, together with their pasturelands;
1CHR|6|74|from the tribe of Asher they received Mashal, Abdon,
1CHR|6|75|Hukok and Rehob, together with their pasturelands;
1CHR|6|76|and from the tribe of Naphtali they received Kedesh in Galilee, Hammon and Kiriathaim, together with their pasturelands.
1CHR|6|77|The Merarites (the rest of the Levites) received the following: From the tribe of Zebulun they received Jokneam, Kartah, Rimmono and Tabor, together with their pasturelands;
1CHR|6|78|from the tribe of Reuben across the Jordan east of Jericho they received Bezer in the desert, Jahzah,
1CHR|6|79|Kedemoth and Mephaath, together with their pasturelands;
1CHR|6|80|and from the tribe of Gad they received Ramoth in Gilead, Mahanaim,
1CHR|6|81|Heshbon and Jazer, together with their pasturelands.
1CHR|7|1|The sons of Issachar: Tola, Puah, Jashub and Shimron-four in all.
1CHR|7|2|The sons of Tola: Uzzi, Rephaiah, Jeriel, Jahmai, Ibsam and Samuel-heads of their families. During the reign of David, the descendants of Tola listed as fighting men in their genealogy numbered 22,600.
1CHR|7|3|The son of Uzzi: Izrahiah. The sons of Izrahiah: Michael, Obadiah, Joel and Isshiah. All five of them were chiefs.
1CHR|7|4|According to their family genealogy, they had 36,000 men ready for battle, for they had many wives and children.
1CHR|7|5|The relatives who were fighting men belonging to all the clans of Issachar, as listed in their genealogy, were 87,000 in all.
1CHR|7|6|Three sons of Benjamin: Bela, Beker and Jediael.
1CHR|7|7|The sons of Bela: Ezbon, Uzzi, Uzziel, Jerimoth and Iri, heads of families-five in all. Their genealogical record listed 22,034 fighting men.
1CHR|7|8|The sons of Beker: Zemirah, Joash, Eliezer, Elioenai, Omri, Jeremoth, Abijah, Anathoth and Alemeth. All these were the sons of Beker.
1CHR|7|9|Their genealogical record listed the heads of families and 20,200 fighting men.
1CHR|7|10|The son of Jediael: Bilhan. The sons of Bilhan: Jeush, Benjamin, Ehud, Kenaanah, Zethan, Tarshish and Ahishahar.
1CHR|7|11|All these sons of Jediael were heads of families. There were 17,200 fighting men ready to go out to war.
1CHR|7|12|The Shuppites and Huppites were the descendants of Ir, and the Hushites the descendants of Aher.
1CHR|7|13|The sons of Naphtali: Jahziel, Guni, Jezer and Shillem -the descendants of Bilhah.
1CHR|7|14|The descendants of Manasseh: Asriel was his descendant through his Aramean concubine. She gave birth to Makir the father of Gilead.
1CHR|7|15|Makir took a wife from among the Huppites and Shuppites. His sister's name was Maacah. Another descendant was named Zelophehad, who had only daughters.
1CHR|7|16|Makir's wife Maacah gave birth to a son and named him Peresh. His brother was named Sheresh, and his sons were Ulam and Rakem.
1CHR|7|17|The son of Ulam: Bedan. These were the sons of Gilead son of Makir, the son of Manasseh.
1CHR|7|18|His sister Hammoleketh gave birth to Ishhod, Abiezer and Mahlah.
1CHR|7|19|The sons of Shemida were: Ahian, Shechem, Likhi and Aniam.
1CHR|7|20|The descendants of Ephraim: Shuthelah, Bered his son, Tahath his son, Eleadah his son, Tahath his son,
1CHR|7|21|Zabad his son and Shuthelah his son. Ezer and Elead were killed by the native-born men of Gath, when they went down to seize their livestock.
1CHR|7|22|Their father Ephraim mourned for them many days, and his relatives came to comfort him.
1CHR|7|23|Then he lay with his wife again, and she became pregnant and gave birth to a son. He named him Beriah, because there had been misfortune in his family.
1CHR|7|24|His daughter was Sheerah, who built Lower and Upper Beth Horon as well as Uzzen Sheerah.
1CHR|7|25|Rephah was his son, Resheph his son, Telah his son, Tahan his son,
1CHR|7|26|Ladan his son, Ammihud his son, Elishama his son,
1CHR|7|27|Nun his son and Joshua his son.
1CHR|7|28|Their lands and settlements included Bethel and its surrounding villages, Naaran to the east, Gezer and its villages to the west, and Shechem and its villages all the way to Ayyah and its villages.
1CHR|7|29|Along the borders of Manasseh were Beth Shan, Taanach, Megiddo and Dor, together with their villages. The descendants of Joseph son of Israel lived in these towns.
1CHR|7|30|The sons of Asher: Imnah, Ishvah, Ishvi and Beriah. Their sister was Serah.
1CHR|7|31|The sons of Beriah: Heber and Malkiel, who was the father of Birzaith.
1CHR|7|32|Heber was the father of Japhlet, Shomer and Hotham and of their sister Shua.
1CHR|7|33|The sons of Japhlet: Pasach, Bimhal and Ashvath. These were Japhlet's sons.
1CHR|7|34|The sons of Shomer: Ahi, Rohgah, Hubbah and Aram.
1CHR|7|35|The sons of his brother Helem: Zophah, Imna, Shelesh and Amal.
1CHR|7|36|The sons of Zophah: Suah, Harnepher, Shual, Beri, Imrah,
1CHR|7|37|Bezer, Hod, Shamma, Shilshah, Ithran and Beera.
1CHR|7|38|The sons of Jether: Jephunneh, Pispah and Ara.
1CHR|7|39|The sons of Ulla: Arah, Hanniel and Rizia.
1CHR|7|40|All these were descendants of Asher-heads of families, choice men, brave warriors and outstanding leaders. The number of men ready for battle, as listed in their genealogy, was 26,000.
1CHR|8|1|Benjamin was the father of Bela his firstborn, Ashbel the second son, Aharah the third,
1CHR|8|2|Nohah the fourth and Rapha the fifth.
1CHR|8|3|The sons of Bela were: Addar, Gera, Abihud,
1CHR|8|4|Abishua, Naaman, Ahoah,
1CHR|8|5|Gera, Shephuphan and Huram.
1CHR|8|6|These were the descendants of Ehud, who were heads of families of those living in Geba and were deported to Manahath:
1CHR|8|7|Naaman, Ahijah, and Gera, who deported them and who was the father of Uzza and Ahihud.
1CHR|8|8|Sons were born to Shaharaim in Moab after he had divorced his wives Hushim and Baara.
1CHR|8|9|By his wife Hodesh he had Jobab, Zibia, Mesha, Malcam,
1CHR|8|10|Jeuz, Sakia and Mirmah. These were his sons, heads of families.
1CHR|8|11|By Hushim he had Abitub and Elpaal.
1CHR|8|12|The sons of Elpaal: Eber, Misham, Shemed (who built Ono and Lod with its surrounding villages),
1CHR|8|13|and Beriah and Shema, who were heads of families of those living in Aijalon and who drove out the inhabitants of Gath.
1CHR|8|14|Ahio, Shashak, Jeremoth,
1CHR|8|15|Zebadiah, Arad, Eder,
1CHR|8|16|Michael, Ishpah and Joha were the sons of Beriah.
1CHR|8|17|Zebadiah, Meshullam, Hizki, Heber,
1CHR|8|18|Ishmerai, Izliah and Jobab were the sons of Elpaal.
1CHR|8|19|Jakim, Zicri, Zabdi,
1CHR|8|20|Elienai, Zillethai, Eliel,
1CHR|8|21|Adaiah, Beraiah and Shimrath were the sons of Shimei.
1CHR|8|22|Ishpan, Eber, Eliel,
1CHR|8|23|Abdon, Zicri, Hanan,
1CHR|8|24|Hananiah, Elam, Anthothijah,
1CHR|8|25|Iphdeiah and Penuel were the sons of Shashak.
1CHR|8|26|Shamsherai, Shehariah, Athaliah,
1CHR|8|27|Jaareshiah, Elijah and Zicri were the sons of Jeroham.
1CHR|8|28|All these were heads of families, chiefs as listed in their genealogy, and they lived in Jerusalem.
1CHR|8|29|Jeiel the father of Gibeon lived in Gibeon. His wife's name was Maacah,
1CHR|8|30|and his firstborn son was Abdon, followed by Zur, Kish, Baal, Ner, Nadab,
1CHR|8|31|Gedor, Ahio, Zeker
1CHR|8|32|and Mikloth, who was the father of Shimeah. They too lived near their relatives in Jerusalem.
1CHR|8|33|Ner was the father of Kish, Kish the father of Saul, and Saul the father of Jonathan, Malki-Shua, Abinadab and Esh-Baal.
1CHR|8|34|The son of Jonathan: Merib-Baal, who was the father of Micah.
1CHR|8|35|The sons of Micah: Pithon, Melech, Tarea and Ahaz.
1CHR|8|36|Ahaz was the father of Jehoaddah, Jehoaddah was the father of Alemeth, Azmaveth and Zimri, and Zimri was the father of Moza.
1CHR|8|37|Moza was the father of Binea; Raphah was his son, Eleasah his son and Azel his son.
1CHR|8|38|Azel had six sons, and these were their names: Azrikam, Bokeru, Ishmael, Sheariah, Obadiah and Hanan. All these were the sons of Azel.
1CHR|8|39|The sons of his brother Eshek: Ulam his firstborn, Jeush the second son and Eliphelet the third.
1CHR|8|40|The sons of Ulam were brave warriors who could handle the bow. They had many sons and grandsons-150 in all. All these were the descendants of Benjamin.
1CHR|9|1|All Israel was listed in the genealogies recorded in the book of the kings of Israel. The people of Judah were taken captive to Babylon because of their unfaithfulness.
1CHR|9|2|Now the first to resettle on their own property in their own towns were some Israelites, priests, Levites and temple servants.
1CHR|9|3|Those from Judah, from Benjamin, and from Ephraim and Manasseh who lived in Jerusalem were:
1CHR|9|4|Uthai son of Ammihud, the son of Omri, the son of Imri, the son of Bani, a descendant of Perez son of Judah.
1CHR|9|5|Of the Shilonites: Asaiah the firstborn and his sons.
1CHR|9|6|Of the Zerahites: Jeuel. The people from Judah numbered 690.
1CHR|9|7|Of the Benjamites: Sallu son of Meshullam, the son of Hodaviah, the son of Hassenuah;
1CHR|9|8|Ibneiah son of Jeroham; Elah son of Uzzi, the son of Micri; and Meshullam son of Shephatiah, the son of Reuel, the son of Ibnijah.
1CHR|9|9|The people from Benjamin, as listed in their genealogy, numbered 956. All these men were heads of their families.
1CHR|9|10|Of the priests: Jedaiah; Jehoiarib; Jakin;
1CHR|9|11|Azariah son of Hilkiah, the son of Meshullam, the son of Zadok, the son of Meraioth, the son of Ahitub, the official in charge of the house of God;
1CHR|9|12|Adaiah son of Jeroham, the son of Pashhur, the son of Malkijah; and Maasai son of Adiel, the son of Jahzerah, the son of Meshullam, the son of Meshillemith, the son of Immer.
1CHR|9|13|The priests, who were heads of families, numbered 1,760. They were able men, responsible for ministering in the house of God.
1CHR|9|14|Of the Levites: Shemaiah son of Hasshub, the son of Azrikam, the son of Hashabiah, a Merarite;
1CHR|9|15|Bakbakkar, Heresh, Galal and Mattaniah son of Mica, the son of Zicri, the son of Asaph;
1CHR|9|16|Obadiah son of Shemaiah, the son of Galal, the son of Jeduthun; and Berekiah son of Asa, the son of Elkanah, who lived in the villages of the Netophathites.
1CHR|9|17|The gatekeepers: Shallum, Akkub, Talmon, Ahiman and their brothers, Shallum their chief
1CHR|9|18|being stationed at the King's Gate on the east, up to the present time. These were the gatekeepers belonging to the camp of the Levites.
1CHR|9|19|Shallum son of Kore, the son of Ebiasaph, the son of Korah, and his fellow gatekeepers from his family (the Korahites) were responsible for guarding the thresholds of the Tent just as their fathers had been responsible for guarding the entrance to the dwelling of the LORD.
1CHR|9|20|In earlier times Phinehas son of Eleazar was in charge of the gatekeepers, and the LORD was with him.
1CHR|9|21|Zechariah son of Meshelemiah was the gatekeeper at the entrance to the Tent of Meeting.
1CHR|9|22|Altogether, those chosen to be gatekeepers at the thresholds numbered 212. They were registered by genealogy in their villages. The gatekeepers had been assigned to their positions of trust by David and Samuel the seer.
1CHR|9|23|They and their descendants were in charge of guarding the gates of the house of the LORD -the house called the Tent.
1CHR|9|24|The gatekeepers were on the four sides: east, west, north and south.
1CHR|9|25|Their brothers in their villages had to come from time to time and share their duties for seven-day periods.
1CHR|9|26|But the four principal gatekeepers, who were Levites, were entrusted with the responsibility for the rooms and treasuries in the house of God.
1CHR|9|27|They would spend the night stationed around the house of God, because they had to guard it; and they had charge of the key for opening it each morning.
1CHR|9|28|Some of them were in charge of the articles used in the temple service; they counted them when they were brought in and when they were taken out.
1CHR|9|29|Others were assigned to take care of the furnishings and all the other articles of the sanctuary, as well as the flour and wine, and the oil, incense and spices.
1CHR|9|30|But some of the priests took care of mixing the spices.
1CHR|9|31|A Levite named Mattithiah, the firstborn son of Shallum the Korahite, was entrusted with the responsibility for baking the offering bread.
1CHR|9|32|Some of their Kohathite brothers were in charge of preparing for every Sabbath the bread set out on the table.
1CHR|9|33|Those who were musicians, heads of Levite families, stayed in the rooms of the temple and were exempt from other duties because they were responsible for the work day and night.
1CHR|9|34|All these were heads of Levite families, chiefs as listed in their genealogy, and they lived in Jerusalem.
1CHR|9|35|Jeiel the father of Gibeon lived in Gibeon. His wife's name was Maacah,
1CHR|9|36|and his firstborn son was Abdon, followed by Zur, Kish, Baal, Ner, Nadab,
1CHR|9|37|Gedor, Ahio, Zechariah and Mikloth.
1CHR|9|38|Mikloth was the father of Shimeam. They too lived near their relatives in Jerusalem.
1CHR|9|39|Ner was the father of Kish, Kish the father of Saul, and Saul the father of Jonathan, Malki-Shua, Abinadab and Esh-Baal.
1CHR|9|40|The son of Jonathan: Merib-Baal, who was the father of Micah.
1CHR|9|41|The sons of Micah: Pithon, Melech, Tahrea and Ahaz.
1CHR|9|42|Ahaz was the father of Jadah, Jadah was the father of Alemeth, Azmaveth and Zimri, and Zimri was the father of Moza.
1CHR|9|43|Moza was the father of Binea; Rephaiah was his son, Eleasah his son and Azel his son.
1CHR|9|44|Azel had six sons, and these were their names: Azrikam, Bokeru, Ishmael, Sheariah, Obadiah and Hanan. These were the sons of Azel.
1CHR|10|1|Now the Philistines fought against Israel; the Israelites fled before them, and many fell slain on Mount Gilboa.
1CHR|10|2|The Philistines pressed hard after Saul and his sons, and they killed his sons Jonathan, Abinadab and Malki-Shua.
1CHR|10|3|The fighting grew fierce around Saul, and when the archers overtook him, they wounded him.
1CHR|10|4|Saul said to his armor-bearer, "Draw your sword and run me through, or these uncircumcised fellows will come and abuse me." But his armor-bearer was terrified and would not do it; so Saul took his own sword and fell on it.
1CHR|10|5|When the armor-bearer saw that Saul was dead, he too fell on his sword and died.
1CHR|10|6|So Saul and his three sons died, and all his house died together.
1CHR|10|7|When all the Israelites in the valley saw that the army had fled and that Saul and his sons had died, they abandoned their towns and fled. And the Philistines came and occupied them.
1CHR|10|8|The next day, when the Philistines came to strip the dead, they found Saul and his sons fallen on Mount Gilboa.
1CHR|10|9|They stripped him and took his head and his armor, and sent messengers throughout the land of the Philistines to proclaim the news among their idols and their people.
1CHR|10|10|They put his armor in the temple of their gods and hung up his head in the temple of Dagon.
1CHR|10|11|When all the inhabitants of Jabesh Gilead heard of everything the Philistines had done to Saul,
1CHR|10|12|all their valiant men went and took the bodies of Saul and his sons and brought them to Jabesh. Then they buried their bones under the great tree in Jabesh, and they fasted seven days.
1CHR|10|13|Saul died because he was unfaithful to the LORD; he did not keep the word of the LORD and even consulted a medium for guidance,
1CHR|10|14|and did not inquire of the LORD. So the LORD put him to death and turned the kingdom over to David son of Jesse.
1CHR|11|1|All Israel came together to David at Hebron and said, "We are your own flesh and blood.
1CHR|11|2|In the past, even while Saul was king, you were the one who led Israel on their military campaigns. And the LORD your God said to you, 'You will shepherd my people Israel, and you will become their ruler.'"
1CHR|11|3|When all the elders of Israel had come to King David at Hebron, he made a compact with them at Hebron before the LORD, and they anointed David king over Israel, as the LORD had promised through Samuel.
1CHR|11|4|David and all the Israelites marched to Jerusalem (that is, Jebus). The Jebusites who lived there
1CHR|11|5|said to David, "You will not get in here." Nevertheless, David captured the fortress of Zion, the City of David.
1CHR|11|6|David had said, "Whoever leads the attack on the Jebusites will become commander-in-chief." Joab son of Zeruiah went up first, and so he received the command.
1CHR|11|7|David then took up residence in the fortress, and so it was called the City of David.
1CHR|11|8|He built up the city around it, from the supporting terraces to the surrounding wall, while Joab restored the rest of the city.
1CHR|11|9|And David became more and more powerful, because the LORD Almighty was with him.
1CHR|11|10|These were the chiefs of David's mighty men-they, together with all Israel, gave his kingship strong support to extend it over the whole land, as the LORD had promised-
1CHR|11|11|this is the list of David's mighty men: Jashobeam, a Hacmonite, was chief of the officers; he raised his spear against three hundred men, whom he killed in one encounter.
1CHR|11|12|Next to him was Eleazar son of Dodai the Ahohite, one of the three mighty men.
1CHR|11|13|He was with David at Pas Dammim when the Philistines gathered there for battle. At a place where there was a field full of barley, the troops fled from the Philistines.
1CHR|11|14|But they took their stand in the middle of the field. They defended it and struck the Philistines down, and the LORD brought about a great victory.
1CHR|11|15|Three of the thirty chiefs came down to David to the rock at the cave of Adullam, while a band of Philistines was encamped in the Valley of Rephaim.
1CHR|11|16|At that time David was in the stronghold, and the Philistine garrison was at Bethlehem.
1CHR|11|17|David longed for water and said, "Oh, that someone would get me a drink of water from the well near the gate of Bethlehem!"
1CHR|11|18|So the Three broke through the Philistine lines, drew water from the well near the gate of Bethlehem and carried it back to David. But he refused to drink it; instead, he poured it out before the LORD.
1CHR|11|19|"God forbid that I should do this!" he said. "Should I drink the blood of these men who went at the risk of their lives?" Because they risked their lives to bring it back, David would not drink it. Such were the exploits of the three mighty men.
1CHR|11|20|Abishai the brother of Joab was chief of the Three. He raised his spear against three hundred men, whom he killed, and so he became as famous as the Three.
1CHR|11|21|He was doubly honored above the Three and became their commander, even though he was not included among them.
1CHR|11|22|Benaiah son of Jehoiada was a valiant fighter from Kabzeel, who performed great exploits. He struck down two of Moab's best men. He also went down into a pit on a snowy day and killed a lion.
1CHR|11|23|And he struck down an Egyptian who was seven and a half feet tall. Although the Egyptian had a spear like a weaver's rod in his hand, Benaiah went against him with a club. He snatched the spear from the Egyptian's hand and killed him with his own spear.
1CHR|11|24|Such were the exploits of Benaiah son of Jehoiada; he too was as famous as the three mighty men.
1CHR|11|25|He was held in greater honor than any of the Thirty, but he was not included among the Three. And David put him in charge of his bodyguard.
1CHR|11|26|The mighty men were: Asahel the brother of Joab, Elhanan son of Dodo from Bethlehem,
1CHR|11|27|Shammoth the Harorite, Helez the Pelonite,
1CHR|11|28|Ira son of Ikkesh from Tekoa, Abiezer from Anathoth,
1CHR|11|29|Sibbecai the Hushathite, Ilai the Ahohite,
1CHR|11|30|Maharai the Netophathite, Heled son of Baanah the Netophathite,
1CHR|11|31|Ithai son of Ribai from Gibeah in Benjamin, Benaiah the Pirathonite,
1CHR|11|32|Hurai from the ravines of Gaash, Abiel the Arbathite,
1CHR|11|33|Azmaveth the Baharumite, Eliahba the Shaalbonite,
1CHR|11|34|the sons of Hashem the Gizonite, Jonathan son of Shagee the Hararite,
1CHR|11|35|Ahiam son of Sacar the Hararite, Eliphal son of Ur,
1CHR|11|36|Hepher the Mekerathite, Ahijah the Pelonite,
1CHR|11|37|Hezro the Carmelite, Naarai son of Ezbai,
1CHR|11|38|Joel the brother of Nathan, Mibhar son of Hagri,
1CHR|11|39|Zelek the Ammonite, Naharai the Berothite, the armor-bearer of Joab son of Zeruiah,
1CHR|11|40|Ira the Ithrite, Gareb the Ithrite,
1CHR|11|41|Uriah the Hittite, Zabad son of Ahlai,
1CHR|11|42|Adina son of Shiza the Reubenite, who was chief of the Reubenites, and the thirty with him,
1CHR|11|43|Hanan son of Maacah, Joshaphat the Mithnite,
1CHR|11|44|Uzzia the Ashterathite, Shama and Jeiel the sons of Hotham the Aroerite,
1CHR|11|45|Jediael son of Shimri, his brother Joha the Tizite,
1CHR|11|46|Eliel the Mahavite, Jeribai and Joshaviah the sons of Elnaam, Ithmah the Moabite,
1CHR|11|47|Eliel, Obed and Jaasiel the Mezobaite.
1CHR|12|1|These were the men who came to David at Ziklag, while he was banished from the presence of Saul son of Kish (they were among the warriors who helped him in battle;
1CHR|12|2|they were armed with bows and were able to shoot arrows or to sling stones right-handed or left-handed; they were kinsmen of Saul from the tribe of Benjamin):
1CHR|12|3|Ahiezer their chief and Joash the sons of Shemaah the Gibeathite; Jeziel and Pelet the sons of Azmaveth; Beracah, Jehu the Anathothite,
1CHR|12|4|and Ishmaiah the Gibeonite, a mighty man among the Thirty, who was a leader of the Thirty; Jeremiah, Jahaziel, Johanan, Jozabad the Gederathite,
1CHR|12|5|Eluzai, Jerimoth, Bealiah, Shemariah and Shephatiah the Haruphite;
1CHR|12|6|Elkanah, Isshiah, Azarel, Joezer and Jashobeam the Korahites;
1CHR|12|7|and Joelah and Zebadiah the sons of Jeroham from Gedor.
1CHR|12|8|Some Gadites defected to David at his stronghold in the desert. They were brave warriors, ready for battle and able to handle the shield and spear. Their faces were the faces of lions, and they were as swift as gazelles in the mountains.
1CHR|12|9|Ezer was the chief, Obadiah the second in command, Eliab the third,
1CHR|12|10|Mishmannah the fourth, Jeremiah the fifth,
1CHR|12|11|Attai the sixth, Eliel the seventh,
1CHR|12|12|Johanan the eighth, Elzabad the ninth,
1CHR|12|13|Jeremiah the tenth and Macbannai the eleventh.
1CHR|12|14|These Gadites were army commanders; the least was a match for a hundred, and the greatest for a thousand.
1CHR|12|15|It was they who crossed the Jordan in the first month when it was overflowing all its banks, and they put to flight everyone living in the valleys, to the east and to the west.
1CHR|12|16|Other Benjamites and some men from Judah also came to David in his stronghold.
1CHR|12|17|David went out to meet them and said to them, "If you have come to me in peace, to help me, I am ready to have you unite with me. But if you have come to betray me to my enemies when my hands are free from violence, may the God of our fathers see it and judge you."
1CHR|12|18|Then the Spirit came upon Amasai, chief of the Thirty, and he said: "We are yours, O David! We are with you, O son of Jesse! Success, success to you, and success to those who help you, for your God will help you." So David received them and made them leaders of his raiding bands.
1CHR|12|19|Some of the men of Manasseh defected to David when he went with the Philistines to fight against Saul. (He and his men did not help the Philistines because, after consultation, their rulers sent him away. They said, "It will cost us our heads if he deserts to his master Saul.")
1CHR|12|20|When David went to Ziklag, these were the men of Manasseh who defected to him: Adnah, Jozabad, Jediael, Michael, Jozabad, Elihu and Zillethai, leaders of units of a thousand in Manasseh.
1CHR|12|21|They helped David against raiding bands, for all of them were brave warriors, and they were commanders in his army.
1CHR|12|22|Day after day men came to help David, until he had a great army, like the army of God.
1CHR|12|23|These are the numbers of the men armed for battle who came to David at Hebron to turn Saul's kingdom over to him, as the LORD had said:
1CHR|12|24|men of Judah, carrying shield and spear-6,800 armed for battle;
1CHR|12|25|men of Simeon, warriors ready for battle-7,100;
1CHR|12|26|men of Levi-4,600,
1CHR|12|27|including Jehoiada, leader of the family of Aaron, with 3,700 men,
1CHR|12|28|and Zadok, a brave young warrior, with 22 officers from his family;
1CHR|12|29|men of Benjamin, Saul's kinsmen-3,000, most of whom had remained loyal to Saul's house until then;
1CHR|12|30|men of Ephraim, brave warriors, famous in their own clans-20,800;
1CHR|12|31|men of half the tribe of Manasseh, designated by name to come and make David king-18,000;
1CHR|12|32|men of Issachar, who understood the times and knew what Israel should do-200 chiefs, with all their relatives under their command;
1CHR|12|33|men of Zebulun, experienced soldiers prepared for battle with every type of weapon, to help David with undivided loyalty-50,000;
1CHR|12|34|men of Naphtali-1,000 officers, together with 37,000 men carrying shields and spears;
1CHR|12|35|men of Dan, ready for battle-28,600;
1CHR|12|36|men of Asher, experienced soldiers prepared for battle-40,000;
1CHR|12|37|and from east of the Jordan, men of Reuben, Gad and the half-tribe of Manasseh, armed with every type of weapon-120,000.
1CHR|12|38|All these were fighting men who volunteered to serve in the ranks. They came to Hebron fully determined to make David king over all Israel. All the rest of the Israelites were also of one mind to make David king.
1CHR|12|39|The men spent three days there with David, eating and drinking, for their families had supplied provisions for them.
1CHR|12|40|Also, their neighbors from as far away as Issachar, Zebulun and Naphtali came bringing food on donkeys, camels, mules and oxen. There were plentiful supplies of flour, fig cakes, raisin cakes, wine, oil, cattle and sheep, for there was joy in Israel.
1CHR|13|1|David conferred with each of his officers, the commanders of thousands and commanders of hundreds.
1CHR|13|2|He then said to the whole assembly of Israel, "If it seems good to you and if it is the will of the LORD our God, let us send word far and wide to the rest of our brothers throughout the territories of Israel, and also to the priests and Levites who are with them in their towns and pasturelands, to come and join us.
1CHR|13|3|Let us bring the ark of our God back to us, for we did not inquire of it during the reign of Saul."
1CHR|13|4|The whole assembly agreed to do this, because it seemed right to all the people.
1CHR|13|5|So David assembled all the Israelites, from the Shihor River in Egypt to Lebo Hamath, to bring the ark of God from Kiriath Jearim.
1CHR|13|6|David and all the Israelites with him went to Baalah of Judah (Kiriath Jearim) to bring up from there the ark of God the LORD, who is enthroned between the cherubim-the ark that is called by the Name.
1CHR|13|7|They moved the ark of God from Abinadab's house on a new cart, with Uzzah and Ahio guiding it.
1CHR|13|8|David and all the Israelites were celebrating with all their might before God, with songs and with harps, lyres, tambourines, cymbals and trumpets.
1CHR|13|9|When they came to the threshing floor of Kidon, Uzzah reached out his hand to steady the ark, because the oxen stumbled.
1CHR|13|10|The LORD's anger burned against Uzzah, and he struck him down because he had put his hand on the ark. So he died there before God.
1CHR|13|11|Then David was angry because the LORD's wrath had broken out against Uzzah, and to this day that place is called Perez Uzzah.
1CHR|13|12|David was afraid of God that day and asked, "How can I ever bring the ark of God to me?"
1CHR|13|13|He did not take the ark to be with him in the City of David. Instead, he took it aside to the house of Obed-Edom the Gittite.
1CHR|13|14|The ark of God remained with the family of Obed-Edom in his house for three months, and the LORD blessed his household and everything he had.
1CHR|14|1|Now Hiram king of Tyre sent messengers to David, along with cedar logs, stonemasons and carpenters to build a palace for him.
1CHR|14|2|And David knew that the LORD had established him as king over Israel and that his kingdom had been highly exalted for the sake of his people Israel.
1CHR|14|3|In Jerusalem David took more wives and became the father of more sons and daughters.
1CHR|14|4|These are the names of the children born to him there: Shammua, Shobab, Nathan, Solomon,
1CHR|14|5|Ibhar, Elishua, Elpelet,
1CHR|14|6|Nogah, Nepheg, Japhia,
1CHR|14|7|Elishama, Beeliada and Eliphelet.
1CHR|14|8|When the Philistines heard that David had been anointed king over all Israel, they went up in full force to search for him, but David heard about it and went out to meet them.
1CHR|14|9|Now the Philistines had come and raided the Valley of Rephaim;
1CHR|14|10|so David inquired of God: "Shall I go and attack the Philistines? Will you hand them over to me?" The LORD answered him, "Go, I will hand them over to you."
1CHR|14|11|So David and his men went up to Baal Perazim, and there he defeated them. He said, "As waters break out, God has broken out against my enemies by my hand." So that place was called Baal Perazim.
1CHR|14|12|The Philistines had abandoned their gods there, and David gave orders to burn them in the fire.
1CHR|14|13|Once more the Philistines raided the valley;
1CHR|14|14|so David inquired of God again, and God answered him, "Do not go straight up, but circle around them and attack them in front of the balsam trees.
1CHR|14|15|As soon as you hear the sound of marching in the tops of the balsam trees, move out to battle, because that will mean God has gone out in front of you to strike the Philistine army."
1CHR|14|16|So David did as God commanded him, and they struck down the Philistine army, all the way from Gibeon to Gezer.
1CHR|14|17|So David's fame spread throughout every land, and the LORD made all the nations fear him.
1CHR|15|1|After David had constructed buildings for himself in the City of David, he prepared a place for the ark of God and pitched a tent for it.
1CHR|15|2|Then David said, "No one but the Levites may carry the ark of God, because the LORD chose them to carry the ark of the LORD and to minister before him forever."
1CHR|15|3|David assembled all Israel in Jerusalem to bring up the ark of the LORD to the place he had prepared for it.
1CHR|15|4|He called together the descendants of Aaron and the Levites:
1CHR|15|5|From the descendants of Kohath, Uriel the leader and 120 relatives;
1CHR|15|6|from the descendants of Merari, Asaiah the leader and 220 relatives;
1CHR|15|7|from the descendants of Gershon, Joel the leader and 130 relatives;
1CHR|15|8|from the descendants of Elizaphan, Shemaiah the leader and 200 relatives;
1CHR|15|9|from the descendants of Hebron, Eliel the leader and 80 relatives;
1CHR|15|10|from the descendants of Uzziel, Amminadab the leader and 112 relatives.
1CHR|15|11|Then David summoned Zadok and Abiathar the priests, and Uriel, Asaiah, Joel, Shemaiah, Eliel and Amminadab the Levites.
1CHR|15|12|He said to them, "You are the heads of the Levitical families; you and your fellow Levites are to consecrate yourselves and bring up the ark of the LORD, the God of Israel, to the place I have prepared for it.
1CHR|15|13|It was because you, the Levites, did not bring it up the first time that the LORD our God broke out in anger against us. We did not inquire of him about how to do it in the prescribed way."
1CHR|15|14|So the priests and Levites consecrated themselves in order to bring up the ark of the LORD, the God of Israel.
1CHR|15|15|And the Levites carried the ark of God with the poles on their shoulders, as Moses had commanded in accordance with the word of the LORD.
1CHR|15|16|David told the leaders of the Levites to appoint their brothers as singers to sing joyful songs, accompanied by musical instruments: lyres, harps and cymbals.
1CHR|15|17|So the Levites appointed Heman son of Joel; from his brothers, Asaph son of Berekiah; and from their brothers the Merarites, Ethan son of Kushaiah;
1CHR|15|18|and with them their brothers next in rank: Zechariah, Jaaziel, Shemiramoth, Jehiel, Unni, Eliab, Benaiah, Maaseiah, Mattithiah, Eliphelehu, Mikneiah, Obed-Edom and Jeiel, the gatekeepers.
1CHR|15|19|The musicians Heman, Asaph and Ethan were to sound the bronze cymbals;
1CHR|15|20|Zechariah, Aziel, Shemiramoth, Jehiel, Unni, Eliab, Maaseiah and Benaiah were to play the lyres according to alamoth,
1CHR|15|21|and Mattithiah, Eliphelehu, Mikneiah, Obed-Edom, Jeiel and Azaziah were to play the harps, directing according to sheminith.
1CHR|15|22|Kenaniah the head Levite was in charge of the singing; that was his responsibility because he was skillful at it.
1CHR|15|23|Berekiah and Elkanah were to be doorkeepers for the ark.
1CHR|15|24|Shebaniah, Joshaphat, Nethanel, Amasai, Zechariah, Benaiah and Eliezer the priests were to blow trumpets before the ark of God. Obed-Edom and Jehiah were also to be doorkeepers for the ark.
1CHR|15|25|So David and the elders of Israel and the commanders of units of a thousand went to bring up the ark of the covenant of the LORD from the house of Obed-Edom, with rejoicing.
1CHR|15|26|Because God had helped the Levites who were carrying the ark of the covenant of the LORD, seven bulls and seven rams were sacrificed.
1CHR|15|27|Now David was clothed in a robe of fine linen, as were all the Levites who were carrying the ark, and as were the singers, and Kenaniah, who was in charge of the singing of the choirs. David also wore a linen ephod.
1CHR|15|28|So all Israel brought up the ark of the covenant of the LORD with shouts, with the sounding of rams' horns and trumpets, and of cymbals, and the playing of lyres and harps.
1CHR|15|29|As the ark of the covenant of the LORD was entering the City of David, Michal daughter of Saul watched from a window. And when she saw King David dancing and celebrating, she despised him in her heart.
1CHR|16|1|They brought the ark of God and set it inside the tent that David had pitched for it, and they presented burnt offerings and fellowship offerings before God.
1CHR|16|2|After David had finished sacrificing the burnt offerings and fellowship offerings, he blessed the people in the name of the LORD.
1CHR|16|3|Then he gave a loaf of bread, a cake of dates and a cake of raisins to each Israelite man and woman.
1CHR|16|4|He appointed some of the Levites to minister before the ark of the LORD, to make petition, to give thanks, and to praise the LORD, the God of Israel:
1CHR|16|5|Asaph was the chief, Zechariah second, then Jeiel, Shemiramoth, Jehiel, Mattithiah, Eliab, Benaiah, Obed-Edom and Jeiel. They were to play the lyres and harps, Asaph was to sound the cymbals,
1CHR|16|6|and Benaiah and Jahaziel the priests were to blow the trumpets regularly before the ark of the covenant of God.
1CHR|16|7|That day David first committed to Asaph and his associates this psalm of thanks to the LORD:
1CHR|16|8|Give thanks to the LORD, call on his name; make known among the nations what he has done.
1CHR|16|9|Sing to him, sing praise to him; tell of all his wonderful acts.
1CHR|16|10|Glory in his holy name; let the hearts of those who seek the LORD rejoice.
1CHR|16|11|Look to the LORD and his strength; seek his face always.
1CHR|16|12|Remember the wonders he has done, his miracles, and the judgments he pronounced,
1CHR|16|13|O descendants of Israel his servant, O sons of Jacob, his chosen ones.
1CHR|16|14|He is the LORD our God; his judgments are in all the earth.
1CHR|16|15|He remembers his covenant forever, the word he commanded, for a thousand generations,
1CHR|16|16|the covenant he made with Abraham, the oath he swore to Isaac.
1CHR|16|17|He confirmed it to Jacob as a decree, to Israel as an everlasting covenant:
1CHR|16|18|"To you I will give the land of Canaan as the portion you will inherit."
1CHR|16|19|When they were but few in number, few indeed, and strangers in it,
1CHR|16|20|they wandered from nation to nation, from one kingdom to another.
1CHR|16|21|He allowed no man to oppress them; for their sake he rebuked kings:
1CHR|16|22|"Do not touch my anointed ones; do my prophets no harm."
1CHR|16|23|Sing to the LORD, all the earth; proclaim his salvation day after day.
1CHR|16|24|Declare his glory among the nations, his marvelous deeds among all peoples.
1CHR|16|25|For great is the LORD and most worthy of praise; he is to be feared above all gods.
1CHR|16|26|For all the gods of the nations are idols, but the LORD made the heavens.
1CHR|16|27|Splendor and majesty are before him; strength and joy in his dwelling place.
1CHR|16|28|Ascribe to the LORD, O families of nations, ascribe to the LORD glory and strength,
1CHR|16|29|ascribe to the LORD the glory due his name. Bring an offering and come before him; worship the LORD in the splendor of his holiness.
1CHR|16|30|Tremble before him, all the earth! The world is firmly established; it cannot be moved.
1CHR|16|31|Let the heavens rejoice, let the earth be glad; let them say among the nations, "The LORD reigns!"
1CHR|16|32|Let the sea resound, and all that is in it; let the fields be jubilant, and everything in them!
1CHR|16|33|Then the trees of the forest will sing, they will sing for joy before the LORD, for he comes to judge the earth.
1CHR|16|34|Give thanks to the LORD, for he is good; his love endures forever.
1CHR|16|35|Cry out, "Save us, O God our Savior; gather us and deliver us from the nations, that we may give thanks to your holy name, that we may glory in your praise."
1CHR|16|36|Praise be to the LORD, the God of Israel, from everlasting to everlasting. Then all the people said "Amen" and "Praise the LORD."
1CHR|16|37|David left Asaph and his associates before the ark of the covenant of the LORD to minister there regularly, according to each day's requirements.
1CHR|16|38|He also left Obed-Edom and his sixty-eight associates to minister with them. Obed-Edom son of Jeduthun, and also Hosah, were gatekeepers.
1CHR|16|39|David left Zadok the priest and his fellow priests before the tabernacle of the LORD at the high place in Gibeon
1CHR|16|40|to present burnt offerings to the LORD on the altar of burnt offering regularly, morning and evening, in accordance with everything written in the Law of the LORD, which he had given Israel.
1CHR|16|41|With them were Heman and Jeduthun and the rest of those chosen and designated by name to give thanks to the LORD, "for his love endures forever."
1CHR|16|42|Heman and Jeduthun were responsible for the sounding of the trumpets and cymbals and for the playing of the other instruments for sacred song. The sons of Jeduthun were stationed at the gate.
1CHR|16|43|Then all the people left, each for his own home, and David returned home to bless his family.
1CHR|17|1|After David was settled in his palace, he said to Nathan the prophet, "Here I am, living in a palace of cedar, while the ark of the covenant of the LORD is under a tent."
1CHR|17|2|Nathan replied to David, "Whatever you have in mind, do it, for God is with you."
1CHR|17|3|That night the word of God came to Nathan, saying:
1CHR|17|4|"Go and tell my servant David, 'This is what the LORD says: You are not the one to build me a house to dwell in.
1CHR|17|5|I have not dwelt in a house from the day I brought Israel up out of Egypt to this day. I have moved from one tent site to another, from one dwelling place to another.
1CHR|17|6|Wherever I have moved with all the Israelites, did I ever say to any of their leaders whom I commanded to shepherd my people, "Why have you not built me a house of cedar?"'
1CHR|17|7|"Now then, tell my servant David, 'This is what the LORD Almighty says: I took you from the pasture and from following the flock, to be ruler over my people Israel.
1CHR|17|8|I have been with you wherever you have gone, and I have cut off all your enemies from before you. Now I will make your name like the names of the greatest men of the earth.
1CHR|17|9|And I will provide a place for my people Israel and will plant them so that they can have a home of their own and no longer be disturbed. Wicked people will not oppress them anymore, as they did at the beginning
1CHR|17|10|and have done ever since the time I appointed leaders over my people Israel. I will also subdue all your enemies. "'I declare to you that the LORD will build a house for you:
1CHR|17|11|When your days are over and you go to be with your fathers, I will raise up your offspring to succeed you, one of your own sons, and I will establish his kingdom.
1CHR|17|12|He is the one who will build a house for me, and I will establish his throne forever.
1CHR|17|13|I will be his father, and he will be my son. I will never take my love away from him, as I took it away from your predecessor.
1CHR|17|14|I will set him over my house and my kingdom forever; his throne will be established forever.'"
1CHR|17|15|Nathan reported to David all the words of this entire revelation.
1CHR|17|16|Then King David went in and sat before the LORD, and he said: "Who am I, O LORD God, and what is my family, that you have brought me this far?
1CHR|17|17|And as if this were not enough in your sight, O God, you have spoken about the future of the house of your servant. You have looked on me as though I were the most exalted of men, O LORD God.
1CHR|17|18|"What more can David say to you for honoring your servant? For you know your servant,
1CHR|17|19|O LORD. For the sake of your servant and according to your will, you have done this great thing and made known all these great promises.
1CHR|17|20|"There is no one like you, O LORD, and there is no God but you, as we have heard with our own ears.
1CHR|17|21|And who is like your people Israel-the one nation on earth whose God went out to redeem a people for himself, and to make a name for yourself, and to perform great and awesome wonders by driving out nations from before your people, whom you redeemed from Egypt?
1CHR|17|22|You made your people Israel your very own forever, and you, O LORD, have become their God.
1CHR|17|23|"And now, LORD, let the promise you have made concerning your servant and his house be established forever. Do as you promised,
1CHR|17|24|so that it will be established and that your name will be great forever. Then men will say, 'The LORD Almighty, the God over Israel, is Israel's God!' And the house of your servant David will be established before you.
1CHR|17|25|"You, my God, have revealed to your servant that you will build a house for him. So your servant has found courage to pray to you.
1CHR|17|26|O LORD, you are God! You have promised these good things to your servant.
1CHR|17|27|Now you have been pleased to bless the house of your servant, that it may continue forever in your sight; for you, O LORD, have blessed it, and it will be blessed forever."
1CHR|18|1|In the course of time, David defeated the Philistines and subdued them, and he took Gath and its surrounding villages from the control of the Philistines.
1CHR|18|2|David also defeated the Moabites, and they became subject to him and brought tribute.
1CHR|18|3|Moreover, David fought Hadadezer king of Zobah, as far as Hamath, when he went to establish his control along the Euphrates River.
1CHR|18|4|David captured a thousand of his chariots, seven thousand charioteers and twenty thousand foot soldiers. He hamstrung all but a hundred of the chariot horses.
1CHR|18|5|When the Arameans of Damascus came to help Hadadezer king of Zobah, David struck down twenty-two thousand of them.
1CHR|18|6|He put garrisons in the Aramean kingdom of Damascus, and the Arameans became subject to him and brought tribute. The LORD gave David victory everywhere he went.
1CHR|18|7|David took the gold shields carried by the officers of Hadadezer and brought them to Jerusalem.
1CHR|18|8|From Tebah and Cun, towns that belonged to Hadadezer, David took a great quantity of bronze, which Solomon used to make the bronze Sea, the pillars and various bronze articles.
1CHR|18|9|When Tou king of Hamath heard that David had defeated the entire army of Hadadezer king of Zobah,
1CHR|18|10|he sent his son Hadoram to King David to greet him and congratulate him on his victory in battle over Hadadezer, who had been at war with Tou. Hadoram brought all kinds of articles of gold and silver and bronze.
1CHR|18|11|King David dedicated these articles to the LORD, as he had done with the silver and gold he had taken from all these nations: Edom and Moab, the Ammonites and the Philistines, and Amalek.
1CHR|18|12|Abishai son of Zeruiah struck down eighteen thousand Edomites in the Valley of Salt.
1CHR|18|13|He put garrisons in Edom, and all the Edomites became subject to David. The LORD gave David victory everywhere he went.
1CHR|18|14|David reigned over all Israel, doing what was just and right for all his people.
1CHR|18|15|Joab son of Zeruiah was over the army; Jehoshaphat son of Ahilud was recorder;
1CHR|18|16|Zadok son of Ahitub and Ahimelech son of Abiathar were priests; Shavsha was secretary;
1CHR|18|17|Benaiah son of Jehoiada was over the Kerethites and Pelethites; and David's sons were chief officials at the king's side.
1CHR|19|1|In the course of time, Nahash king of the Ammonites died, and his son succeeded him as king.
1CHR|19|2|David thought, "I will show kindness to Hanun son of Nahash, because his father showed kindness to me." So David sent a delegation to express his sympathy to Hanun concerning his father. When David's men came to Hanun in the land of the Ammonites to express sympathy to him,
1CHR|19|3|the Ammonite nobles said to Hanun, "Do you think David is honoring your father by sending men to you to express sympathy? Haven't his men come to you to explore and spy out the country and overthrow it?"
1CHR|19|4|So Hanun seized David's men, shaved them, cut off their garments in the middle at the buttocks, and sent them away.
1CHR|19|5|When someone came and told David about the men, he sent messengers to meet them, for they were greatly humiliated. The king said, "Stay at Jericho till your beards have grown, and then come back."
1CHR|19|6|When the Ammonites realized that they had become a stench in David's nostrils, Hanun and the Ammonites sent a thousand talents of silver to hire chariots and charioteers from Aram Naharaim, Aram Maacah and Zobah.
1CHR|19|7|They hired thirty-two thousand chariots and charioteers, as well as the king of Maacah with his troops, who came and camped near Medeba, while the Ammonites were mustered from their towns and moved out for battle.
1CHR|19|8|On hearing this, David sent Joab out with the entire army of fighting men.
1CHR|19|9|The Ammonites came out and drew up in battle formation at the entrance to their city, while the kings who had come were by themselves in the open country.
1CHR|19|10|Joab saw that there were battle lines in front of him and behind him; so he selected some of the best troops in Israel and deployed them against the Arameans.
1CHR|19|11|He put the rest of the men under the command of Abishai his brother, and they were deployed against the Ammonites.
1CHR|19|12|Joab said, "If the Arameans are too strong for me, then you are to rescue me; but if the Ammonites are too strong for you, then I will rescue you.
1CHR|19|13|Be strong and let us fight bravely for our people and the cities of our God. The LORD will do what is good in his sight."
1CHR|19|14|Then Joab and the troops with him advanced to fight the Arameans, and they fled before him.
1CHR|19|15|When the Ammonites saw that the Arameans were fleeing, they too fled before his brother Abishai and went inside the city. So Joab went back to Jerusalem.
1CHR|19|16|After the Arameans saw that they had been routed by Israel, they sent messengers and had Arameans brought from beyond the River, with Shophach the commander of Hadadezer's army leading them.
1CHR|19|17|When David was told of this, he gathered all Israel and crossed the Jordan; he advanced against them and formed his battle lines opposite them. David formed his lines to meet the Arameans in battle, and they fought against him.
1CHR|19|18|But they fled before Israel, and David killed seven thousand of their charioteers and forty thousand of their foot soldiers. He also killed Shophach the commander of their army.
1CHR|19|19|When the vassals of Hadadezer saw that they had been defeated by Israel, they made peace with David and became subject to him. So the Arameans were not willing to help the Ammonites anymore.
1CHR|20|1|In the spring, at the time when kings go off to war, Joab led out the armed forces. He laid waste the land of the Ammonites and went to Rabbah and besieged it, but David remained in Jerusalem. Joab attacked Rabbah and left it in ruins.
1CHR|20|2|David took the crown from the head of their king -its weight was found to be a talent of gold, and it was set with precious stones-and it was placed on David's head. He took a great quantity of plunder from the city
1CHR|20|3|and brought out the people who were there, consigning them to labor with saws and with iron picks and axes. David did this to all the Ammonite towns. Then David and his entire army returned to Jerusalem.
1CHR|20|4|In the course of time, war broke out with the Philistines, at Gezer. At that time Sibbecai the Hushathite killed Sippai, one of the descendants of the Rephaites, and the Philistines were subjugated.
1CHR|20|5|In another battle with the Philistines, Elhanan son of Jair killed Lahmi the brother of Goliath the Gittite, who had a spear with a shaft like a weaver's rod.
1CHR|20|6|In still another battle, which took place at Gath, there was a huge man with six fingers on each hand and six toes on each foot-twenty-four in all. He also was descended from Rapha.
1CHR|20|7|When he taunted Israel, Jonathan son of Shimea, David's brother, killed him.
1CHR|20|8|These were descendants of Rapha in Gath, and they fell at the hands of David and his men.
1CHR|21|1|Satan rose up against Israel and incited David to take a census of Israel.
1CHR|21|2|So David said to Joab and the commanders of the troops, "Go and count the Israelites from Beersheba to Dan. Then report back to me so that I may know how many there are."
1CHR|21|3|But Joab replied, "May the LORD multiply his troops a hundred times over. My lord the king, are they not all my lord's subjects? Why does my lord want to do this? Why should he bring guilt on Israel?"
1CHR|21|4|The king's word, however, overruled Joab; so Joab left and went throughout Israel and then came back to Jerusalem.
1CHR|21|5|Joab reported the number of the fighting men to David: In all Israel there were one million one hundred thousand men who could handle a sword, including four hundred and seventy thousand in Judah.
1CHR|21|6|But Joab did not include Levi and Benjamin in the numbering, because the king's command was repulsive to him.
1CHR|21|7|This command was also evil in the sight of God; so he punished Israel.
1CHR|21|8|Then David said to God, "I have sinned greatly by doing this. Now, I beg you, take away the guilt of your servant. I have done a very foolish thing."
1CHR|21|9|The LORD said to Gad, David's seer,
1CHR|21|10|"Go and tell David, 'This is what the LORD says: I am giving you three options. Choose one of them for me to carry out against you.'"
1CHR|21|11|So Gad went to David and said to him, "This is what the LORD says: 'Take your choice:
1CHR|21|12|three years of famine, three months of being swept away before your enemies, with their swords overtaking you, or three days of the sword of the LORD -days of plague in the land, with the angel of the LORD ravaging every part of Israel.' Now then, decide how I should answer the one who sent me."
1CHR|21|13|David said to Gad, "I am in deep distress. Let me fall into the hands of the LORD, for his mercy is very great; but do not let me fall into the hands of men."
1CHR|21|14|So the LORD sent a plague on Israel, and seventy thousand men of Israel fell dead.
1CHR|21|15|And God sent an angel to destroy Jerusalem. But as the angel was doing so, the LORD saw it and was grieved because of the calamity and said to the angel who was destroying the people, "Enough! Withdraw your hand." The angel of the LORD was then standing at the threshing floor of Araunah the Jebusite.
1CHR|21|16|David looked up and saw the angel of the LORD standing between heaven and earth, with a drawn sword in his hand extended over Jerusalem. Then David and the elders, clothed in sackcloth, fell facedown.
1CHR|21|17|David said to God, "Was it not I who ordered the fighting men to be counted? I am the one who has sinned and done wrong. These are but sheep. What have they done? O LORD my God, let your hand fall upon me and my family, but do not let this plague remain on your people."
1CHR|21|18|Then the angel of the LORD ordered Gad to tell David to go up and build an altar to the LORD on the threshing floor of Araunah the Jebusite.
1CHR|21|19|So David went up in obedience to the word that Gad had spoken in the name of the LORD.
1CHR|21|20|While Araunah was threshing wheat, he turned and saw the angel; his four sons who were with him hid themselves.
1CHR|21|21|Then David approached, and when Araunah looked and saw him, he left the threshing floor and bowed down before David with his face to the ground.
1CHR|21|22|David said to him, "Let me have the site of your threshing floor so I can build an altar to the LORD, that the plague on the people may be stopped. Sell it to me at the full price."
1CHR|21|23|Araunah said to David, "Take it! Let my lord the king do whatever pleases him. Look, I will give the oxen for the burnt offerings, the threshing sledges for the wood, and the wheat for the grain offering. I will give all this."
1CHR|21|24|But King David replied to Araunah, "No, I insist on paying the full price. I will not take for the LORD what is yours, or sacrifice a burnt offering that costs me nothing."
1CHR|21|25|So David paid Araunah six hundred shekels of gold for the site.
1CHR|21|26|David built an altar to the LORD there and sacrificed burnt offerings and fellowship offerings. He called on the LORD, and the LORD answered him with fire from heaven on the altar of burnt offering.
1CHR|21|27|Then the LORD spoke to the angel, and he put his sword back into its sheath.
1CHR|21|28|At that time, when David saw that the LORD had answered him on the threshing floor of Araunah the Jebusite, he offered sacrifices there.
1CHR|21|29|The tabernacle of the LORD, which Moses had made in the desert, and the altar of burnt offering were at that time on the high place at Gibeon.
1CHR|21|30|But David could not go before it to inquire of God, because he was afraid of the sword of the angel of the LORD.
1CHR|22|1|Then David said, "The house of the LORD God is to be here, and also the altar of burnt offering for Israel."
1CHR|22|2|So David gave orders to assemble the aliens living in Israel, and from among them he appointed stonecutters to prepare dressed stone for building the house of God.
1CHR|22|3|He provided a large amount of iron to make nails for the doors of the gateways and for the fittings, and more bronze than could be weighed.
1CHR|22|4|He also provided more cedar logs than could be counted, for the Sidonians and Tyrians had brought large numbers of them to David.
1CHR|22|5|David said, "My son Solomon is young and inexperienced, and the house to be built for the LORD should be of great magnificence and fame and splendor in the sight of all the nations. Therefore I will make preparations for it." So David made extensive preparations before his death.
1CHR|22|6|Then he called for his son Solomon and charged him to build a house for the LORD, the God of Israel.
1CHR|22|7|David said to Solomon: "My son, I had it in my heart to build a house for the Name of the LORD my God.
1CHR|22|8|But this word of the LORD came to me: 'You have shed much blood and have fought many wars. You are not to build a house for my Name, because you have shed much blood on the earth in my sight.
1CHR|22|9|But you will have a son who will be a man of peace and rest, and I will give him rest from all his enemies on every side. His name will be Solomon, and I will grant Israel peace and quiet during his reign.
1CHR|22|10|He is the one who will build a house for my Name. He will be my son, and I will be his father. And I will establish the throne of his kingdom over Israel forever.'
1CHR|22|11|"Now, my son, the LORD be with you, and may you have success and build the house of the LORD your God, as he said you would.
1CHR|22|12|May the LORD give you discretion and understanding when he puts you in command over Israel, so that you may keep the law of the LORD your God.
1CHR|22|13|Then you will have success if you are careful to observe the decrees and laws that the LORD gave Moses for Israel. Be strong and courageous. Do not be afraid or discouraged.
1CHR|22|14|"I have taken great pains to provide for the temple of the LORD a hundred thousand talents of gold, a million talents of silver, quantities of bronze and iron too great to be weighed, and wood and stone. And you may add to them.
1CHR|22|15|You have many workmen: stonecutters, masons and carpenters, as well as men skilled in every kind of work
1CHR|22|16|in gold and silver, bronze and iron-craftsmen beyond number. Now begin the work, and the LORD be with you."
1CHR|22|17|Then David ordered all the leaders of Israel to help his son Solomon.
1CHR|22|18|He said to them, "Is not the LORD your God with you? And has he not granted you rest on every side? For he has handed the inhabitants of the land over to me, and the land is subject to the LORD and to his people.
1CHR|22|19|Now devote your heart and soul to seeking the LORD your God. Begin to build the sanctuary of the LORD God, so that you may bring the ark of the covenant of the LORD and the sacred articles belonging to God into the temple that will be built for the Name of the LORD."
1CHR|23|1|When David was old and full of years, he made his son Solomon king over Israel.
1CHR|23|2|He also gathered together all the leaders of Israel, as well as the priests and Levites.
1CHR|23|3|The Levites thirty years old or more were counted, and the total number of men was thirty-eight thousand.
1CHR|23|4|David said, "Of these, twenty-four thousand are to supervise the work of the temple of the LORD and six thousand are to be officials and judges.
1CHR|23|5|Four thousand are to be gatekeepers and four thousand are to praise the LORD with the musical instruments I have provided for that purpose."
1CHR|23|6|David divided the Levites into groups corresponding to the sons of Levi: Gershon, Kohath and Merari.
1CHR|23|7|Belonging to the Gershonites: Ladan and Shimei.
1CHR|23|8|The sons of Ladan: Jehiel the first, Zetham and Joel-three in all.
1CHR|23|9|The sons of Shimei: Shelomoth, Haziel and Haran-three in all. These were the heads of the families of Ladan.
1CHR|23|10|And the sons of Shimei: Jahath, Ziza, Jeush and Beriah. These were the sons of Shimei-four in all.
1CHR|23|11|Jahath was the first and Ziza the second, but Jeush and Beriah did not have many sons; so they were counted as one family with one assignment.
1CHR|23|12|The sons of Kohath: Amram, Izhar, Hebron and Uzziel-four in all.
1CHR|23|13|The sons of Amram: Aaron and Moses. Aaron was set apart, he and his descendants forever, to consecrate the most holy things, to offer sacrifices before the LORD, to minister before him and to pronounce blessings in his name forever.
1CHR|23|14|The sons of Moses the man of God were counted as part of the tribe of Levi.
1CHR|23|15|The sons of Moses: Gershom and Eliezer.
1CHR|23|16|The descendants of Gershom: Shubael was the first.
1CHR|23|17|The descendants of Eliezer: Rehabiah was the first. Eliezer had no other sons, but the sons of Rehabiah were very numerous.
1CHR|23|18|The sons of Izhar: Shelomith was the first.
1CHR|23|19|The sons of Hebron: Jeriah the first, Amariah the second, Jahaziel the third and Jekameam the fourth.
1CHR|23|20|The sons of Uzziel: Micah the first and Isshiah the second.
1CHR|23|21|The sons of Merari: Mahli and Mushi. The sons of Mahli: Eleazar and Kish.
1CHR|23|22|Eleazar died without having sons: he had only daughters. Their cousins, the sons of Kish, married them.
1CHR|23|23|The sons of Mushi: Mahli, Eder and Jerimoth-three in all.
1CHR|23|24|These were the descendants of Levi by their families-the heads of families as they were registered under their names and counted individually, that is, the workers twenty years old or more who served in the temple of the LORD.
1CHR|23|25|For David had said, "Since the LORD, the God of Israel, has granted rest to his people and has come to dwell in Jerusalem forever,
1CHR|23|26|the Levites no longer need to carry the tabernacle or any of the articles used in its service."
1CHR|23|27|According to the last instructions of David, the Levites were counted from those twenty years old or more.
1CHR|23|28|The duty of the Levites was to help Aaron's descendants in the service of the temple of the LORD: to be in charge of the courtyards, the side rooms, the purification of all sacred things and the performance of other duties at the house of God.
1CHR|23|29|They were in charge of the bread set out on the table, the flour for the grain offerings, the unleavened wafers, the baking and the mixing, and all measurements of quantity and size.
1CHR|23|30|They were also to stand every morning to thank and praise the LORD. They were to do the same in the evening
1CHR|23|31|and whenever burnt offerings were presented to the LORD on Sabbaths and at New Moon festivals and at appointed feasts. They were to serve before the LORD regularly in the proper number and in the way prescribed for them.
1CHR|23|32|And so the Levites carried out their responsibilities for the Tent of Meeting, for the Holy Place and, under their brothers the descendants of Aaron, for the service of the temple of the LORD.
1CHR|24|1|These were the divisions of the sons of Aaron: The sons of Aaron were Nadab, Abihu, Eleazar and Ithamar.
1CHR|24|2|But Nadab and Abihu died before their father did, and they had no sons; so Eleazar and Ithamar served as the priests.
1CHR|24|3|With the help of Zadok a descendant of Eleazar and Ahimelech a descendant of Ithamar, David separated them into divisions for their appointed order of ministering.
1CHR|24|4|A larger number of leaders were found among Eleazar's descendants than among Ithamar's, and they were divided accordingly: sixteen heads of families from Eleazar's descendants and eight heads of families from Ithamar's descendants.
1CHR|24|5|They divided them impartially by drawing lots, for there were officials of the sanctuary and officials of God among the descendants of both Eleazar and Ithamar.
1CHR|24|6|The scribe Shemaiah son of Nethanel, a Levite, recorded their names in the presence of the king and of the officials: Zadok the priest, Ahimelech son of Abiathar and the heads of families of the priests and of the Levites-one family being taken from Eleazar and then one from Ithamar.
1CHR|24|7|The first lot fell to Jehoiarib, the second to Jedaiah,
1CHR|24|8|the third to Harim, the fourth to Seorim,
1CHR|24|9|the fifth to Malkijah, the sixth to Mijamin,
1CHR|24|10|the seventh to Hakkoz, the eighth to Abijah,
1CHR|24|11|the ninth to Jeshua, the tenth to Shecaniah,
1CHR|24|12|the eleventh to Eliashib, the twelfth to Jakim,
1CHR|24|13|the thirteenth to Huppah, the fourteenth to Jeshebeab,
1CHR|24|14|the fifteenth to Bilgah, the sixteenth to Immer,
1CHR|24|15|the seventeenth to Hezir, the eighteenth to Happizzez,
1CHR|24|16|the nineteenth to Pethahiah, the twentieth to Jehezkel,
1CHR|24|17|the twenty-first to Jakin, the twenty-second to Gamul,
1CHR|24|18|the twenty-third to Delaiah and the twenty-fourth to Maaziah.
1CHR|24|19|This was their appointed order of ministering when they entered the temple of the LORD, according to the regulations prescribed for them by their forefather Aaron, as the LORD, the God of Israel, had commanded him.
1CHR|24|20|As for the rest of the descendants of Levi: from the sons of Amram: Shubael; from the sons of Shubael: Jehdeiah.
1CHR|24|21|As for Rehabiah, from his sons: Isshiah was the first.
1CHR|24|22|From the Izharites: Shelomoth; from the sons of Shelomoth: Jahath.
1CHR|24|23|The sons of Hebron: Jeriah the first, Amariah the second, Jahaziel the third and Jekameam the fourth.
1CHR|24|24|The son of Uzziel: Micah; from the sons of Micah: Shamir.
1CHR|24|25|The brother of Micah: Isshiah; from the sons of Isshiah: Zechariah.
1CHR|24|26|The sons of Merari: Mahli and Mushi. The son of Jaaziah: Beno.
1CHR|24|27|The sons of Merari: from Jaaziah: Beno, Shoham, Zaccur and Ibri.
1CHR|24|28|From Mahli: Eleazar, who had no sons.
1CHR|24|29|From Kish: the son of Kish: Jerahmeel.
1CHR|24|30|And the sons of Mushi: Mahli, Eder and Jerimoth. These were the Levites, according to their families.
1CHR|24|31|They also cast lots, just as their brothers the descendants of Aaron did, in the presence of King David and of Zadok, Ahimelech, and the heads of families of the priests and of the Levites. The families of the oldest brother were treated the same as those of the youngest.
1CHR|25|1|David, together with the commanders of the army, set apart some of the sons of Asaph, Heman and Jeduthun for the ministry of prophesying, accompanied by harps, lyres and cymbals. Here is the list of the men who performed this service:
1CHR|25|2|From the sons of Asaph: Zaccur, Joseph, Nethaniah and Asarelah. The sons of Asaph were under the supervision of Asaph, who prophesied under the king's supervision.
1CHR|25|3|As for Jeduthun, from his sons: Gedaliah, Zeri, Jeshaiah, Shimei, Hashabiah and Mattithiah, six in all, under the supervision of their father Jeduthun, who prophesied, using the harp in thanking and praising the LORD.
1CHR|25|4|As for Heman, from his sons: Bukkiah, Mattaniah, Uzziel, Shubael and Jerimoth; Hananiah, Hanani, Eliathah, Giddalti and Romamti-Ezer; Joshbekashah, Mallothi, Hothir and Mahazioth.
1CHR|25|5|All these were sons of Heman the king's seer. They were given him through the promises of God to exalt him. God gave Heman fourteen sons and three daughters.
1CHR|25|6|All these men were under the supervision of their fathers for the music of the temple of the LORD, with cymbals, lyres and harps, for the ministry at the house of God. Asaph, Jeduthun and Heman were under the supervision of the king.
1CHR|25|7|Along with their relatives-all of them trained and skilled in music for the LORD -they numbered 288.
1CHR|25|8|Young and old alike, teacher as well as student, cast lots for their duties.
1CHR|25|9|The first lot, which was for Asaph, fell to Joseph, his sons and relatives, 12 the second to Gedaliah, he and his relatives and sons, 12
1CHR|25|10|the third to Zaccur, his sons and relatives, 12
1CHR|25|11|the fourth to Izri, his sons and relatives, 12
1CHR|25|12|the fifth to Nethaniah, his sons and relatives, 12
1CHR|25|13|the sixth to Bukkiah, his sons and relatives, 12
1CHR|25|14|the seventh to Jesarelah, his sons and relatives, 12
1CHR|25|15|the eighth to Jeshaiah, his sons and relatives, 12
1CHR|25|16|the ninth to Mattaniah, his sons and relatives, 12
1CHR|25|17|the tenth to Shimei, his sons and relatives, 12
1CHR|25|18|the eleventh to Azarel, his sons and relatives, 12
1CHR|25|19|the twelfth to Hashabiah, his sons and relatives, 12
1CHR|25|20|the thirteenth to Shubael, his sons and relatives, 12
1CHR|25|21|the fourteenth to Mattithiah, his sons and relatives, 12
1CHR|25|22|the fifteenth to Jerimoth, his sons and relatives, 12
1CHR|25|23|the sixteenth to Hananiah, his sons and relatives, 12
1CHR|25|24|the seventeenth to Joshbekashah, his sons and relatives, 12
1CHR|25|25|the eighteenth to Hanani, his sons and relatives, 12
1CHR|25|26|the nineteenth to Mallothi, his sons and relatives, 12
1CHR|25|27|the twentieth to Eliathah, his sons and relatives, 12
1CHR|25|28|the twenty-first to Hothir, his sons and relatives, 12
1CHR|25|29|the twenty-second to Giddalti, his sons and relatives, 12
1CHR|25|30|the twenty-third to Mahazioth, his sons and relatives, 12
1CHR|25|31|the twenty-fourth to Romamti-Ezer, his sons and relatives, 12
1CHR|26|1|The divisions of the gatekeepers: From the Korahites: Meshelemiah son of Kore, one of the sons of Asaph.
1CHR|26|2|Meshelemiah had sons: Zechariah the firstborn, Jediael the second, Zebadiah the third, Jathniel the fourth,
1CHR|26|3|Elam the fifth, Jehohanan the sixth and Eliehoenai the seventh.
1CHR|26|4|Obed-Edom also had sons: Shemaiah the firstborn, Jehozabad the second, Joah the third, Sacar the fourth, Nethanel the fifth,
1CHR|26|5|Ammiel the sixth, Issachar the seventh and Peullethai the eighth. (For God had blessed Obed-Edom.)
1CHR|26|6|His son Shemaiah also had sons, who were leaders in their father's family because they were very capable men.
1CHR|26|7|The sons of Shemaiah: Othni, Rephael, Obed and Elzabad; his relatives Elihu and Semakiah were also able men.
1CHR|26|8|All these were descendants of Obed-Edom; they and their sons and their relatives were capable men with the strength to do the work-descendants of Obed-Edom, 62 in all.
1CHR|26|9|Meshelemiah had sons and relatives, who were able men-18 in all.
1CHR|26|10|Hosah the Merarite had sons: Shimri the first (although he was not the firstborn, his father had appointed him the first),
1CHR|26|11|Hilkiah the second, Tabaliah the third and Zechariah the fourth. The sons and relatives of Hosah were 13 in all.
1CHR|26|12|These divisions of the gatekeepers, through their chief men, had duties for ministering in the temple of the LORD, just as their relatives had.
1CHR|26|13|Lots were cast for each gate, according to their families, young and old alike.
1CHR|26|14|The lot for the East Gate fell to Shelemiah. Then lots were cast for his son Zechariah, a wise counselor, and the lot for the North Gate fell to him.
1CHR|26|15|The lot for the South Gate fell to Obed-Edom, and the lot for the storehouse fell to his sons.
1CHR|26|16|The lots for the West Gate and the Shalleketh Gate on the upper road fell to Shuppim and Hosah. Guard was alongside of guard:
1CHR|26|17|There were six Levites a day on the east, four a day on the north, four a day on the south and two at a time at the storehouse.
1CHR|26|18|As for the court to the west, there were four at the road and two at the court itself.
1CHR|26|19|These were the divisions of the gatekeepers who were descendants of Korah and Merari.
1CHR|26|20|Their fellow Levites were in charge of the treasuries of the house of God and the treasuries for the dedicated things.
1CHR|26|21|The descendants of Ladan, who were Gershonites through Ladan and who were heads of families belonging to Ladan the Gershonite, were Jehieli,
1CHR|26|22|the sons of Jehieli, Zetham and his brother Joel. They were in charge of the treasuries of the temple of the LORD.
1CHR|26|23|From the Amramites, the Izharites, the Hebronites and the Uzzielites:
1CHR|26|24|Shubael, a descendant of Gershom son of Moses, was the officer in charge of the treasuries.
1CHR|26|25|His relatives through Eliezer: Rehabiah his son, Jeshaiah his son, Joram his son, Zicri his son and Shelomith his son.
1CHR|26|26|Shelomith and his relatives were in charge of all the treasuries for the things dedicated by King David, by the heads of families who were the commanders of thousands and commanders of hundreds, and by the other army commanders.
1CHR|26|27|Some of the plunder taken in battle they dedicated for the repair of the temple of the LORD.
1CHR|26|28|And everything dedicated by Samuel the seer and by Saul son of Kish, Abner son of Ner and Joab son of Zeruiah, and all the other dedicated things were in the care of Shelomith and his relatives.
1CHR|26|29|From the Izharites: Kenaniah and his sons were assigned duties away from the temple, as officials and judges over Israel.
1CHR|26|30|From the Hebronites: Hashabiah and his relatives-seventeen hundred able men-were responsible in Israel west of the Jordan for all the work of the LORD and for the king's service.
1CHR|26|31|As for the Hebronites, Jeriah was their chief according to the genealogical records of their families. In the fortieth year of David's reign a search was made in the records, and capable men among the Hebronites were found at Jazer in Gilead.
1CHR|26|32|Jeriah had twenty-seven hundred relatives, who were able men and heads of families, and King David put them in charge of the Reubenites, the Gadites and the half-tribe of Manasseh for every matter pertaining to God and for the affairs of the king.
1CHR|27|1|This is the list of the Israelites-heads of families, commanders of thousands and commanders of hundreds, and their officers, who served the king in all that concerned the army divisions that were on duty month by month throughout the year. Each division consisted of 24,000 men.
1CHR|27|2|In charge of the first division, for the first month, was Jashobeam son of Zabdiel. There were 24,000 men in his division.
1CHR|27|3|He was a descendant of Perez and chief of all the army officers for the first month.
1CHR|27|4|In charge of the division for the second month was Dodai the Ahohite; Mikloth was the leader of his division. There were 24,000 men in his division.
1CHR|27|5|The third army commander, for the third month, was Benaiah son of Jehoiada the priest. He was chief and there were 24,000 men in his division.
1CHR|27|6|This was the Benaiah who was a mighty man among the Thirty and was over the Thirty. His son Ammizabad was in charge of his division.
1CHR|27|7|The fourth, for the fourth month, was Asahel the brother of Joab; his son Zebadiah was his successor. There were 24,000 men in his division.
1CHR|27|8|The fifth, for the fifth month, was the commander Shamhuth the Izrahite. There were 24,000 men in his division.
1CHR|27|9|The sixth, for the sixth month, was Ira the son of Ikkesh the Tekoite. There were 24,000 men in his division.
1CHR|27|10|The seventh, for the seventh month, was Helez the Pelonite, an Ephraimite. There were 24,000 men in his division.
1CHR|27|11|The eighth, for the eighth month, was Sibbecai the Hushathite, a Zerahite. There were 24,000 men in his division.
1CHR|27|12|The ninth, for the ninth month, was Abiezer the Anathothite, a Benjamite. There were 24,000 men in his division.
1CHR|27|13|The tenth, for the tenth month, was Maharai the Netophathite, a Zerahite. There were 24,000 men in his division.
1CHR|27|14|The eleventh, for the eleventh month, was Benaiah the Pirathonite, an Ephraimite. There were 24,000 men in his division.
1CHR|27|15|The twelfth, for the twelfth month, was Heldai the Netophathite, from the family of Othniel. There were 24,000 men in his division.
1CHR|27|16|The officers over the tribes of Israel: over the Reubenites: Eliezer son of Zicri; over the Simeonites: Shephatiah son of Maacah;
1CHR|27|17|over Levi: Hashabiah son of Kemuel; over Aaron: Zadok;
1CHR|27|18|over Judah: Elihu, a brother of David; over Issachar: Omri son of Michael;
1CHR|27|19|over Zebulun: Ishmaiah son of Obadiah; over Naphtali: Jerimoth son of Azriel;
1CHR|27|20|over the Ephraimites: Hoshea son of Azaziah; over half the tribe of Manasseh: Joel son of Pedaiah;
1CHR|27|21|over the half-tribe of Manasseh in Gilead: Iddo son of Zechariah; over Benjamin: Jaasiel son of Abner;
1CHR|27|22|over Dan: Azarel son of Jeroham. These were the officers over the tribes of Israel.
1CHR|27|23|David did not take the number of the men twenty years old or less, because the LORD had promised to make Israel as numerous as the stars in the sky.
1CHR|27|24|Joab son of Zeruiah began to count the men but did not finish. Wrath came on Israel on account of this numbering, and the number was not entered in the book of the annals of King David.
1CHR|27|25|Azmaveth son of Adiel was in charge of the royal storehouses. Jonathan son of Uzziah was in charge of the storehouses in the outlying districts, in the towns, the villages and the watchtowers.
1CHR|27|26|Ezri son of Kelub was in charge of the field workers who farmed the land.
1CHR|27|27|Shimei the Ramathite was in charge of the vineyards. Zabdi the Shiphmite was in charge of the produce of the vineyards for the wine vats.
1CHR|27|28|Baal-Hanan the Gederite was in charge of the olive and sycamore-fig trees in the western foothills. Joash was in charge of the supplies of olive oil.
1CHR|27|29|Shitrai the Sharonite was in charge of the herds grazing in Sharon. Shaphat son of Adlai was in charge of the herds in the valleys.
1CHR|27|30|Obil the Ishmaelite was in charge of the camels. Jehdeiah the Meronothite was in charge of the donkeys.
1CHR|27|31|Jaziz the Hagrite was in charge of the flocks. All these were the officials in charge of King David's property.
1CHR|27|32|Jonathan, David's uncle, was a counselor, a man of insight and a scribe. Jehiel son of Hacmoni took care of the king's sons.
1CHR|27|33|Ahithophel was the king's counselor. Hushai the Arkite was the king's friend.
1CHR|27|34|Ahithophel was succeeded by Jehoiada son of Benaiah and by Abiathar. Joab was the commander of the royal army.
1CHR|28|1|David summoned all the officials of Israel to assemble at Jerusalem: the officers over the tribes, the commanders of the divisions in the service of the king, the commanders of thousands and commanders of hundreds, and the officials in charge of all the property and livestock belonging to the king and his sons, together with the palace officials, the mighty men and all the brave warriors.
1CHR|28|2|King David rose to his feet and said: "Listen to me, my brothers and my people. I had it in my heart to build a house as a place of rest for the ark of the covenant of the LORD, for the footstool of our God, and I made plans to build it.
1CHR|28|3|But God said to me, 'You are not to build a house for my Name, because you are a warrior and have shed blood.'
1CHR|28|4|"Yet the LORD, the God of Israel, chose me from my whole family to be king over Israel forever. He chose Judah as leader, and from the house of Judah he chose my family, and from my father's sons he was pleased to make me king over all Israel.
1CHR|28|5|Of all my sons-and the LORD has given me many-he has chosen my son Solomon to sit on the throne of the kingdom of the LORD over Israel.
1CHR|28|6|He said to me: 'Solomon your son is the one who will build my house and my courts, for I have chosen him to be my son, and I will be his father.
1CHR|28|7|I will establish his kingdom forever if he is unswerving in carrying out my commands and laws, as is being done at this time.'
1CHR|28|8|"So now I charge you in the sight of all Israel and of the assembly of the LORD, and in the hearing of our God: Be careful to follow all the commands of the LORD your God, that you may possess this good land and pass it on as an inheritance to your descendants forever.
1CHR|28|9|"And you, my son Solomon, acknowledge the God of your father, and serve him with wholehearted devotion and with a willing mind, for the LORD searches every heart and understands every motive behind the thoughts. If you seek him, he will be found by you; but if you forsake him, he will reject you forever.
1CHR|28|10|Consider now, for the LORD has chosen you to build a temple as a sanctuary. Be strong and do the work."
1CHR|28|11|Then David gave his son Solomon the plans for the portico of the temple, its buildings, its storerooms, its upper parts, its inner rooms and the place of atonement.
1CHR|28|12|He gave him the plans of all that the Spirit had put in his mind for the courts of the temple of the LORD and all the surrounding rooms, for the treasuries of the temple of God and for the treasuries for the dedicated things.
1CHR|28|13|He gave him instructions for the divisions of the priests and Levites, and for all the work of serving in the temple of the LORD, as well as for all the articles to be used in its service.
1CHR|28|14|He designated the weight of gold for all the gold articles to be used in various kinds of service, and the weight of silver for all the silver articles to be used in various kinds of service:
1CHR|28|15|the weight of gold for the gold lampstands and their lamps, with the weight for each lampstand and its lamps; and the weight of silver for each silver lampstand and its lamps, according to the use of each lampstand;
1CHR|28|16|the weight of gold for each table for consecrated bread; the weight of silver for the silver tables;
1CHR|28|17|the weight of pure gold for the forks, sprinkling bowls and pitchers; the weight of gold for each gold dish; the weight of silver for each silver dish;
1CHR|28|18|and the weight of the refined gold for the altar of incense. He also gave him the plan for the chariot, that is, the cherubim of gold that spread their wings and shelter the ark of the covenant of the LORD.
1CHR|28|19|"All this," David said, "I have in writing from the hand of the LORD upon me, and he gave me understanding in all the details of the plan."
1CHR|28|20|David also said to Solomon his son, "Be strong and courageous, and do the work. Do not be afraid or discouraged, for the LORD God, my God, is with you. He will not fail you or forsake you until all the work for the service of the temple of the LORD is finished.
1CHR|28|21|The divisions of the priests and Levites are ready for all the work on the temple of God, and every willing man skilled in any craft will help you in all the work. The officials and all the people will obey your every command."
1CHR|29|1|Then King David said to the whole assembly: "My son Solomon, the one whom God has chosen, is young and inexperienced. The task is great, because this palatial structure is not for man but for the LORD God.
1CHR|29|2|With all my resources I have provided for the temple of my God-gold for the gold work, silver for the silver, bronze for the bronze, iron for the iron and wood for the wood, as well as onyx for the settings, turquoise, stones of various colors, and all kinds of fine stone and marble-all of these in large quantities.
1CHR|29|3|Besides, in my devotion to the temple of my God I now give my personal treasures of gold and silver for the temple of my God, over and above everything I have provided for this holy temple:
1CHR|29|4|three thousand talents of gold (gold of Ophir) and seven thousand talents of refined silver, for the overlaying of the walls of the buildings,
1CHR|29|5|for the gold work and the silver work, and for all the work to be done by the craftsmen. Now, who is willing to consecrate himself today to the LORD?"
1CHR|29|6|Then the leaders of families, the officers of the tribes of Israel, the commanders of thousands and commanders of hundreds, and the officials in charge of the king's work gave willingly.
1CHR|29|7|They gave toward the work on the temple of God five thousand talents and ten thousand darics of gold, ten thousand talents of silver, eighteen thousand talents of bronze and a hundred thousand talents of iron.
1CHR|29|8|Any who had precious stones gave them to the treasury of the temple of the LORD in the custody of Jehiel the Gershonite.
1CHR|29|9|The people rejoiced at the willing response of their leaders, for they had given freely and wholeheartedly to the LORD. David the king also rejoiced greatly.
1CHR|29|10|David praised the LORD in the presence of the whole assembly, saying, "Praise be to you, O LORD, God of our father Israel, from everlasting to everlasting.
1CHR|29|11|Yours, O LORD, is the greatness and the power and the glory and the majesty and the splendor, for everything in heaven and earth is yours. Yours, O LORD, is the kingdom; you are exalted as head over all.
1CHR|29|12|Wealth and honor come from you; you are the ruler of all things. In your hands are strength and power to exalt and give strength to all.
1CHR|29|13|Now, our God, we give you thanks, and praise your glorious name.
1CHR|29|14|"But who am I, and who are my people, that we should be able to give as generously as this? Everything comes from you, and we have given you only what comes from your hand.
1CHR|29|15|We are aliens and strangers in your sight, as were all our forefathers. Our days on earth are like a shadow, without hope.
1CHR|29|16|O LORD our God, as for all this abundance that we have provided for building you a temple for your Holy Name, it comes from your hand, and all of it belongs to you.
1CHR|29|17|I know, my God, that you test the heart and are pleased with integrity. All these things have I given willingly and with honest intent. And now I have seen with joy how willingly your people who are here have given to you.
1CHR|29|18|O LORD, God of our fathers Abraham, Isaac and Israel, keep this desire in the hearts of your people forever, and keep their hearts loyal to you.
1CHR|29|19|And give my son Solomon the wholehearted devotion to keep your commands, requirements and decrees and to do everything to build the palatial structure for which I have provided."
1CHR|29|20|Then David said to the whole assembly, "Praise the LORD your God." So they all praised the LORD, the God of their fathers; they bowed low and fell prostrate before the LORD and the king.
1CHR|29|21|The next day they made sacrifices to the LORD and presented burnt offerings to him: a thousand bulls, a thousand rams and a thousand male lambs, together with their drink offerings, and other sacrifices in abundance for all Israel.
1CHR|29|22|They ate and drank with great joy in the presence of the LORD that day. Then they acknowledged Solomon son of David as king a second time, anointing him before the LORD to be ruler and Zadok to be priest.
1CHR|29|23|So Solomon sat on the throne of the LORD as king in place of his father David. He prospered and all Israel obeyed him.
1CHR|29|24|All the officers and mighty men, as well as all of King David's sons, pledged their submission to King Solomon.
1CHR|29|25|The LORD highly exalted Solomon in the sight of all Israel and bestowed on him royal splendor such as no king over Israel ever had before.
1CHR|29|26|David son of Jesse was king over all Israel.
1CHR|29|27|He ruled over Israel forty years-seven in Hebron and thirty-three in Jerusalem.
1CHR|29|28|He died at a good old age, having enjoyed long life, wealth and honor. His son Solomon succeeded him as king.
1CHR|29|29|As for the events of King David's reign, from beginning to end, they are written in the records of Samuel the seer, the records of Nathan the prophet and the records of Gad the seer,
1CHR|29|30|together with the details of his reign and power, and the circumstances that surrounded him and Israel and the kingdoms of all the other lands.
