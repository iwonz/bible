TITUS|1|1|Paulus servus Dei apostolus autem Iesu Christi secundum fidem electorum Dei et agnitionem veritatis quae secundum pietatem est
TITUS|1|2|in spem vitae aeternae quam promisit qui non mentitur Deus ante tempora saecularia
TITUS|1|3|manifestavit autem temporibus suis verbum suum in praedicatione quae credita est mihi secundum praeceptum salvatoris nostri Dei
TITUS|1|4|Tito dilecto filio secundum communem fidem gratia et pax a Deo Patre et Christo Iesu salvatore nostro
TITUS|1|5|huius rei gratia reliqui te Cretae ut ea quae desunt corrigas et constituas per civitates presbyteros sicut ego tibi disposui
TITUS|1|6|si quis sine crimine est unius uxoris vir filios habens fideles non in accusatione luxuriae aut non subditos
TITUS|1|7|oportet enim episcopum sine crimine esse sicut Dei dispensatorem non superbum non iracundum non vinolentum non percussorem non turpilucri cupidum
TITUS|1|8|sed hospitalem benignum sobrium iustum sanctum continentem
TITUS|1|9|amplectentem eum qui secundum doctrinam est fidelem sermonem ut potens sit et exhortari in doctrina sana et eos qui contradicunt arguere
TITUS|1|10|sunt enim multi et inoboedientes vaniloqui et seductores maxime qui de circumcisione sunt
TITUS|1|11|quos oportet redargui qui universas domos subvertunt docentes quae non oportet turpis lucri gratia
TITUS|1|12|dixit quidam ex illis proprius ipsorum propheta Cretenses semper mendaces malae bestiae ventres pigri
TITUS|1|13|testimonium hoc verum est quam ob causam increpa illos dure ut sani sint in fide
TITUS|1|14|non intendentes iudaicis fabulis et mandatis hominum aversantium se a veritate
TITUS|1|15|omnia munda mundis coinquinatis autem et infidelibus nihil mundum sed inquinatae sunt eorum et mens et conscientia
TITUS|1|16|confitentur se nosse Deum factis autem negant cum sunt abominati et incredibiles et ad omne opus bonum reprobi
TITUS|2|1|tu autem loquere quae decet sanam doctrinam
TITUS|2|2|senes ut sobrii sint pudici prudentes sani fide dilectione patientia
TITUS|2|3|anus similiter in habitu sancto non criminatrices non vino multo servientes bene docentes
TITUS|2|4|ut prudentiam doceant adulescentulas ut viros suos ament filios diligant
TITUS|2|5|prudentes castas domus curam habentes benignas subditas suis viris ut non blasphemetur verbum Dei
TITUS|2|6|iuvenes similiter hortare ut sobrii sint
TITUS|2|7|in omnibus te ipsum praebe exemplum bonorum operum in doctrina integritatem gravitatem
TITUS|2|8|verbum sanum inreprehensibilem ut is qui ex adverso est vereatur nihil habens malum dicere de nobis
TITUS|2|9|servos dominis suis subditos esse in omnibus placentes non contradicentes
TITUS|2|10|non fraudantes, sed in omnibus fidem bonam ostendentes ut doctrinam salutaris nostri Dei ornent in omnibus
TITUS|2|11|apparuit enim gratia Dei salutaris omnibus hominibus
TITUS|2|12|erudiens nos ut abnegantes impietatem et saecularia desideria sobrie et iuste et pie vivamus in hoc saeculo
TITUS|2|13|expectantes beatam spem et adventum gloriae magni Dei et salvatoris nostri Iesu Christi
TITUS|2|14|qui dedit semet ipsum pro nobis ut nos redimeret ab omni iniquitate et mundaret sibi populum acceptabilem sectatorem bonorum operum
TITUS|2|15|haec loquere et exhortare et argue cum omni imperio nemo te contemnat
TITUS|3|1|admone illos principibus et potestatibus subditos esse dicto oboedire ad omne opus bonum paratos esse
TITUS|3|2|neminem blasphemare non litigiosos esse modestos omnem ostendentes mansuetudinem ad omnes homines
TITUS|3|3|eramus enim et nos aliquando insipientes increduli errantes servientes desideriis et voluptatibus variis in malitia et invidia agentes odibiles odientes invicem
TITUS|3|4|cum autem benignitas et humanitas apparuit salvatoris nostri Dei
TITUS|3|5|non ex operibus iustitiae quae fecimus nos sed secundum suam misericordiam salvos nos fecit per lavacrum regenerationis et renovationis Spiritus Sancti
TITUS|3|6|quem effudit in nos abunde per Iesum Christum salvatorem nostrum
TITUS|3|7|ut iustificati gratia ipsius heredes simus secundum spem vitae aeternae
TITUS|3|8|fidelis sermo est et de his volo te confirmare ut curent bonis operibus praeesse qui credunt Deo haec sunt bona et utilia hominibus
TITUS|3|9|stultas autem quaestiones et genealogias et contentiones et pugnas legis devita sunt enim inutiles et vanae
TITUS|3|10|hereticum hominem post unam et secundam correptionem devita
TITUS|3|11|sciens quia subversus est qui eiusmodi est et delinquit proprio iudicio condemnatus
TITUS|3|12|cum misero ad te Arteman aut Tychicum festina ad me venire Nicopolim ibi enim statui hiemare
TITUS|3|13|Zenan legis peritum et Apollo sollicite praemitte ut nihil illis desit
TITUS|3|14|discant autem et nostri bonis operibus praeesse ad usus necessarios ut non sint infructuosi
TITUS|3|15|salutant te qui mecum sunt omnes saluta qui nos amant in fide gratia Dei cum omnibus vobis amen
