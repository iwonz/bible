HOS|1|1|Verbum Domini, quod factum est ad Osee filium Beeri in die bus Oziae, Ioatham, Achaz, Ezechiae regum Iudae, et in diebus Ieroboam filii Ioas regis Israel.
HOS|1|2|Principium verbi Domini per Osee. Dixit Dominus ad Osee: Vade, sume tibi mulierem fornicationumet filios fornicationum,quia fornicans fornicatur terra a Domino ".
HOS|1|3|Et abiit et accepit Gomer filiam Debelaim, quae concepit et peperit ei filium.
HOS|1|4|Et dixit Dominus ad eum: " Voca nomen eius 'Iezrahel', quoniam adhuc modicum et visitabo sanguinem Iezrahel super domum Iehu et cessare faciam regnum domus Israel;
HOS|1|5|et in illa die conteram arcum Israel in valle Iezrahel ".
HOS|1|6|Et concepit adhuc et peperit filiam; et dixit ei: " Voca nomen eius Absque misericordia", quia non addam ultra misereri domui Israel, ut ignoscam eis.
HOS|1|7|Et domui Iudae miserebor et salvabo eos in Domino Deo suo et non salvabo eos in arcu et gladio et in bello et in equis et in equitibus ".
HOS|1|8|Et ablactavit eam, quae erat 'Absque misericordia', et concepit et peperit filium.
HOS|1|9|Et dixit: " Voca nomen eius 'Non populus meus', quia vos non populus meus, et ego 'Non sum' vobis.
HOS|2|1|Et erit numerus filiorum Israelquasi arena maris,quae sine mensura est et non numerabitur.Et erit: in loco, ubi dicebatur eis:Non populus meus vos",dicetur eis: "Filii Dei viventis".
HOS|2|2|Et congregabuntur filii Iudaeet filii Israel pariteret ponent sibimet caput unumet ascendent de terra,quia magnus dies Iezrahel.
HOS|2|3|Dicite fratribus vestris: "Populus meus"et sororibus vestris: "Misericordiam consecuta".
HOS|2|4|Contendite adversum matrem vestram; contendite,quoniam ipsa non uxor mea,et ego non vir eius;auferat fornicationes suas a facie suaet adulteria sua de medio uberum suorum,
HOS|2|5|ne forte exspoliem eam nudamet statuam eam secundum diem nativitatis suaeet ponam eam quasi solitudinemet statuam eam velut terram aridamet interficiam eam siti.
HOS|2|6|Et filiorum illius non miserebor,quoniam filii fornicationum sunt,
HOS|2|7|quia fornicata est mater eorum,turpiter egit, quae concepit eos;quia dixit: "Vadam post amatores meos,qui dant panes mihi et aquas meas,lanam meam et linum meum,oleum meum et potum meum".
HOS|2|8|Propter hoc ecce ego saepiamviam tuam spiniset saepiam eam maceria,et semitas suas non inveniet;
HOS|2|9|et sequetur amatores suoset non apprehendet eos;et quaeret eos et non invenietet dicet: "Vadam et revertarad virum meum priorem,quia bene mihi erat tunc magis quam nunc".
HOS|2|10|Et haec nescivit quia egodedi ei frumentum et vinum et oleumet argentum multiplicavi eiet aurum, quae fecerunt Baal.
HOS|2|11|Idcirco convertar et sumamfrumentum meum in tempore suoet vinum meum in tempore suo;et auferam lanam meam et linum meum,quae operiebant pudenda eius,
HOS|2|12|et nunc revelabo ignominiam eiusin oculis amatorum eius,et nullus est qui eruat eam de manu mea.
HOS|2|13|Et cessare faciam omne gaudium eius,sollemnitatem eius, neomeniam eius,sabbatum eius et omnia festa tempora eius;
HOS|2|14|et corrumpam vineam eius et ficum eius,de quibus dixit: "Mercedes hae meae sunt,quas dederunt mihi amatores mei".Et ponam eas in saltum,et comedet illas bestia agri.
HOS|2|15|Et visitabo super eam dies Baalim,quibus accendebat incensumet ornabatur inaure sua et monili suoet ibat post amatores suos,sed mei obliviscebatur,dicit Dominus.
HOS|2|16|Propter hoc ecce ego lactabo eamet ducam eam in solitudinemet loquar ad cor eius;
HOS|2|17|et dabo ei vineas eius ex eodem locoet vallem Achor, portam spei,et respondebit ibiiuxta dies iuventutis suaeet iuxta dies ascensionis suae de terra Aegypti.
HOS|2|18|Et erit: in die illa,ait Dominus,vocabis me: "Vir meus"et non vocabis me ultra: "Baal meus".
HOS|2|19|Et auferam nomina Baalim de ore eius,et non recordabitur ultra nominis eorum.
HOS|2|20|Et percutiam eis foedus in die illacum bestia agri et cum volucre caeli et cum reptili terrae;et arcum et gladium et bellumconteram de terraet cubare eos faciam confidenter.
HOS|2|21|Et sponsabo te mihi in sempiternum;et sponsabo te mihi in iustitia et iudicioet in misericordia et miserationibus.
HOS|2|22|Et sponsabo te mihi in fide,et cognosces Dominum.
HOS|2|23|Et erit: in illa die exaudiam,dicit Dominus,exaudiam caelos,et illi exaudient terram;
HOS|2|24|et terra exaudiettriticum et vinum et oleum,et haec exaudient Iezrahel.
HOS|2|25|Et seminabo eam mihi in terramet miserebor eius, quae fuit "Absque misericordia";
HOS|2|26|et dicam "Non populo meo": "Populus meus tu";et ipse dicet: "Deus meus es tu" ".
HOS|3|1|Et dixit Dominus ad me: " Adhuc vade, dilige mulierem dilectam amico et adulteram, sicut diligit Dominus filios Israel, et ipsi respectant ad deos alienos et diligunt placentas uvarum ".
HOS|3|2|Et emi eam mihi quindecim argenteis et choro hordei et dimidio choro hordei.
HOS|3|3|Et dixi ad eam: " Dies multos exspectabis me; non fornicaberis et non eris viro, neque ibo ego ad te ".
HOS|3|4|Quia dies multos sedebunt filii Israel sine rege et sine principe et sine sacrificio et sine lapide et sine ephod et sine theraphim.
HOS|3|5|Et post haec revertentur filii Israel et quaerent Dominum Deum suum et David regem suum et pavebunt ad Dominum et ad bonum eius in fine dierum.
HOS|4|1|" Audite verbum Domini,filii Israel,quia iudicium Dominocum habitatoribus terrae:non est enim veritas, et non est benignitas,et non est scientia Dei in terra;
HOS|4|2|maledictum et mendaciumet homicidium et furtum et adulterium inundaverunt,et sanguis sanguinem tetigit.
HOS|4|3|Propter hoc lugebit terra,et infirmabitur omnis, qui habitat in ea,cum bestia agri et volucre caeli,sed et pisces maris auferentur.
HOS|4|4|Verumtamen non sit qui contendatnec qui arguat,sed tecum iudicium meum, sacerdos.
HOS|4|5|Et corrues plena die,et corruet etiam propheta tecum nocte;et perdam matrem tuam.
HOS|4|6|Perit populus meus,eo quod non habuerit scientiam.Quia tu scientiam reppulisti,repellam te, ne sacerdotio fungaris mihi;et quia oblitus es legis Dei tui,obliviscar filiorum tuorum et ego.
HOS|4|7|Secundum multitudinem eorum, sic peccaverunt mihi;gloriam eorum in ignominiam commutabo.
HOS|4|8|Peccatum populi mei comeduntet ad iniquitatem eorum sublevabunt animas eorum.
HOS|4|9|Et erit sicut populus sic sacerdos;et visitabo super eum vias eiuset opera eius reddam ei.
HOS|4|10|Et comedent et non saturabuntur;fornicabuntur et non multiplicabuntur,quoniam Dominum reliqueruntin non custodiendo.
HOS|4|11|Fornicatio et vinum et ebrietas auferunt cor.
HOS|4|12|Populus meus in ligno suo interrogat,et baculus eius annuntiat ei;spiritus enim fornicationum decepit eos,et fornicantur a Deo suo.
HOS|4|13|Super capita montium sacrificantet super colles accendunt thymiama,subtus quercum et populum et terebinthum,quia bona est umbra eius;ideo fornicantur filiae vestrae,et sponsae vestrae adulterae sunt.
HOS|4|14|Non visitabo super filias vestras,cum fuerint fornicatae,et super sponsas vestras,cum adulteraverint,quoniam hi ipsi cum meretricibus seceduntet cum prostibulis delubrorum sacrificant,et populus non intellegens corruet.
HOS|4|15|Si fornicaris tu, Israel,non delinquat saltem Iuda;et nolite ingredi in Galgalaet ne ascenderitis in Bethavenneque iuraveritis: "Vivit Dominus".
HOS|4|16|Quoniam sicut vacca lasciviensIsrael contumax est;nunc pascet eos Dominusquasi agnum in latitudine?
HOS|4|17|Particeps idolorum Ephraim,dimitte eum.
HOS|4|18|Transiit convivium eorum,fornicatione fornicati sunt,diligunt vehementerignominiam impudicitiae.
HOS|4|19|Ligabit spiritus eos in alis suis,et confundentur a sacrificiis suis.
HOS|5|1|Audite hoc, sacerdotes,et attendite, domus Israel;et domus regis, auscultate,quia vobis iudicium est;quoniam laqueus facti estis pro Masphaet rete expansum super Thabor.
HOS|5|2|Et foveam Settim profundam fecerunt;ego autem castigabo vos omnes.
HOS|5|3|Ego scio Ephraim,et Israel non est absconditus a me;quia nunc fornicatus es, Ephraim,contaminatus est Israel.
HOS|5|4|Non dabunt opera sua,ut revertantur ad Deum suum,quia spiritus fornicationis in medio eorum,et Dominum non cognoverunt.
HOS|5|5|Et testatur arrogantia Israel in faciem suam,et Israel et Ephraim ruent in iniquitate sua:ruet etiam Iudas cum eis.
HOS|5|6|In gregibus suis et in armentis suisvadent ad quaerendum Dominumet non invenient;subtraxit se ab eis.
HOS|5|7|In Dominum praevaricati sunt,quia filios alienos genuerunt;nunc devorabit eos uno mense cum partibus suis.
HOS|5|8|Clangite bucina in Gabaa,tuba in Rama,conclamate in Bethaven,exterrete Beniamin.
HOS|5|9|Ephraim vastabitur in die correptionis;in tribubus Israel annuntio rem certam.
HOS|5|10|Facti sunt principes Iudaequasi transferentes terminos;super eos effundamquasi aquam iram meam.
HOS|5|11|Oppressus est Ephraim,fractum est ius,quoniam voluit abire post sordem.
HOS|5|12|Et ego quasi sanies Ephraim,et quasi putredo domui Iudae.
HOS|5|13|Et vidit Ephraim languorem suum,et Iuda ulcus suum;et abiit Ephraim ad Assyriamet misit ad regem magnum;sed et ipse non poterit sanare vosnec solvere poterit vos ab ulcere.
HOS|5|14|Quoniam ego quasi leaena Ephraimet quasi catulus leonis domui Iudae;ego, ego capiam et vadam,tollam, et non est qui eruat.
HOS|5|15|Vadens revertar ad locum meum,donec poenas solvantet quaerant faciem meam,in tribulatione sua me desiderent.
HOS|6|1|"Venite, et revertamur ad Do minum,quia ipse laceravit et sanabit nos,percussit et curabit nos.
HOS|6|2|Vivificabit nos post duos dies,in die tertia suscitabit nos,et vivemus in conspectu eius.
HOS|6|3|Sciamus sequamurque,ut cognoscamus Dominum.Quasi diluculum praeparatus est egressus eius,et veniet quasi imber nobis temporaneus,quasi imber serotinus irrigans terram".
HOS|6|4|Quid faciam tibi, Ephraim?Quid faciam tibi, Iuda?Caritas vestra quasi nubes matutinaet quasi ros mane pertransiens.
HOS|6|5|Propter hoc dolavi per prophetas,occidi eos in verbis oris mei,sed ius meum quasi lux egredietur;
HOS|6|6|quia caritatem volo et non sacrificium,et scientiam Dei plus quam holocausta.
HOS|6|7|Ipsi autem in Adam transgressi sunt pactum;ibi praevaricati sunt in me.
HOS|6|8|Galaad civitas operantium iniquitatemmaculata sanguine.
HOS|6|9|Et quasi insidiantes virum latronescaterva sacerdotum;in via interficiunt pergentes Sichem,vere scelus operantur.
HOS|6|10|In domo Israel vidi horrendum:ibi fornicationes Ephraim,contaminatus est Israel.
HOS|6|11|Sed et tibi, Iuda, parata est messis,cum convertero sortem populi mei.
HOS|7|1|Cum sanare vellem Israel,revelata est iniquitas Ephraimet malitia Samariae,quia operati sunt mendacium;et fur ingressus est,foris autem spoliat turma latronum.
HOS|7|2|Et non dicunt in cordibus suisomnem malitiam eorum me recordari.Nunc circumdederunt eos opera sua,coram facie mea facta sunt.
HOS|7|3|In malitia sua laetificaverunt regem et in mendaciis suis principes.
HOS|7|4|Omnes adulterantes;quasi clibanus succensus illi,pistor cessat excitare ignema commixtione fermenti, donec fermentetur totum.
HOS|7|5|Die regis nostriinfirmi facti sunt principes ardore vini,quod apprehendit protervos.
HOS|7|6|Quia applicuerunt quasi clibanum cor suumin insidiando;tota nocte dormivit ira eorum,mane ipsa ardet quasi ignis flammae.
HOS|7|7|Omnes calefacti sunt quasi clibanuset devorant iudices suos.Omnes reges eorum ceciderunt;non est qui clamet in eis ad me.
HOS|7|8|Ephraim in populis ipse commiscebatur;Ephraim factus est subcinericius panis, qui non reversatur.
HOS|7|9|Comederunt alieni robur eius,et ipse nescit;sed et cani effusi sunt in eo,et ipse ignorat.
HOS|7|10|Et testatur superbia Israel in faciem suam,nec reversi sunt ad Dominum Deum suumet non quaesierunt eum in omnibus his.
HOS|7|11|Et factus est Ephraim quasi columbainsipiens non habens sensum:Aegyptum invocabant,ad Assyrios abierunt.
HOS|7|12|Et cum profecti fuerint,expandam super eos rete meum;quasi volucrem caeli detraham eos, corripiam eos secundum auditionem coetus eorum.
HOS|7|13|Vae eis, quoniam recesserunt a me!Vastabuntur, quia praevaricati sunt in me.Et ego redimam eos,cum ipsi locuti sint contra me mendacia?
HOS|7|14|Et non clamaverunt ad me in corde suo,sed ululabant in cubilibus suis;super triticum et vinum se incidebant,contumaces sunt adversum me.
HOS|7|15|Et ego erudivi eos et confortavi brachia eorum,et in me cogitaverunt malitiam.
HOS|7|16|Convertuntur ad eum, qui non prodest,facti sunt quasi arcus dolosus;cadent in gladio principes eorumpropter execrationem linguae suae: ista subsannatio eorum in terra Aegypti.
HOS|8|1|In gutture tuo sit tuba!Quasi aquila super domum Do minipro eo quod transgressi sunt foedus meumet legem meam praevaricati sunt.
HOS|8|2|Me invocant: "Deus meus";cognovimus te, Israel.
HOS|8|3|Proiecit Israel bonum;inimicus persequetur eum.
HOS|8|4|Ipsi constituerunt reges, et non ex me;principes constituerunt, et non cognovi:argentum suum et aurum suumfecerunt sibi idola,ut interirent.
HOS|8|5|Proiectus est vitulus tuus, Samaria;iratus est furor meus in eos.Usquequo non poterunt emundari?
HOS|8|6|Quia ex Israel et ipse est:artifex fecit illum,et non est Deus;quoniam in scintillas eritvitulus Samariae.
HOS|8|7|Quia ventum seminabuntet turbinem metent;cum culmus non sit in eo,germen non faciet farinam:quod et si fecerit,alieni comedent eam.
HOS|8|8|Devoratus est Israel,nunc factus est in nationibusquasi vas immundum.
HOS|8|9|Quia ipsi ascenderunt ad Assyriam, onager est solitarius sibi;Ephraim autem munera dederunt amatoribus.
HOS|8|10|Sed et cum mercede conduxerint nationes,nunc compellam eos,et trement paulisper sub onere regis principum.
HOS|8|11|Cum multiplicaret Ephraim altaria pro peccato,factae sunt ei arae in peccatum.
HOS|8|12|Scribebam ei multiplices leges meas;velut alienae computatae sunt.
HOS|8|13|Hostias amant,immolant carnes et comedunt;sed Dominus non suscipiet eas.Nunc recordabitur iniquitatis eorumet visitabit peccata eorum:ipsi in Aegyptum convertentur.
HOS|8|14|Et oblitus est Israel factoris suiet aedificavit delubra;et Iudas multiplicavit urbes munitas.Et mittam ignem in civitates eius,et devorabit aedes illius.
HOS|9|1|Noli laetari, Israel;noli exsultare sicut populi,quia fornicatus es a Deo tuo,dilexisti mercedem super omnes areas tritici.
HOS|9|2|Area et torcular non pascet eos,et vinum mentietur eis.
HOS|9|3|Non manebunt in terra Domini:revertetur Ephraim in Aegyptum,et in Assyria pollutum comedent.
HOS|9|4|Non libabunt Domino vinum,et non placebunt ei sacrificia eorum;quasi panis lugentium erunt eis:omnes, qui comedent eum, contaminabuntur,quia panis eorum erit tantummodo pro vita ipsorum;non intrabit in domum Domini.
HOS|9|5|Quid facietis in die sollemni,in die festivitatis Domini?
HOS|9|6|Ecce enim profecti sunt a vastitate;Aegyptus congregabit eos,Memphis sepeliet eos:desiderabile argentum eorumurtica hereditabit,spina in tabernaculis eorum.
HOS|9|7|Venerunt dies visitationis,venerunt dies retributionis:sciat Israel!Stultus - clamet - est propheta;insanus vir spiritalis".Secundum multitudinem iniquitatis tuaemultae sunt inimicitiae tuae.
HOS|9|8|Speculatur Ephraim, populus Dei mei, prophetam;laqueus aucupis super omnes vias eius,inimicitiae in ipsa domo Dei eius.
HOS|9|9|Profunde peccaveruntsicut in diebus Gabaa;recordabitur iniquitatis eorumet visitabit peccata eorum.
HOS|9|10|Quasi uvas in desertoinveni Israel,quasi prima poma ficulneae in initio eiusvidi patres vestros;ipsi autem intraverunt ad Baalphegoret se consecraverunt Confusioniet facti sunt abominabilessicut id, quod dilexerunt.
HOS|9|11|Ephraim quasi avis avolabit gloria eorum,a partu et ab utero et a conceptu.
HOS|9|12|Quod si et enutrierint filios suos,absque liberis eos faciam, absque hominibus;sed et vae eis,cum recessero ab eis!
HOS|9|13|Ephraim, ut vidi, in venationem posuit sibi filios suos,et Ephraim educit ad interfectorem filios suos.
HOS|9|14|"Da eis, Domine! Quid dabis eis?Da eis vulvam sine liberis et ubera arentia!".
HOS|9|15|Omnes nequitiae eorum in Galgala,profecto ibi exosos habui eos.Propter malitiam operum eorumde domo mea eiciam eos.Non addam ut diligam eos;omnes principes eorum rebelles.
HOS|9|16|Percussus est Ephraim,radix eorum exsiccata est,fructum nequaquam facient;quod si et genuerint,interficiam amantissima uteri eorum ".
HOS|9|17|Abiciet eos Deus meus,quia non audierunt eum;et erunt vagi in nationibus.
HOS|10|1|Vitis frondosa Israel,fructum producens sibi;secundum multitudinem fructus sui multiplicavit altaria,iuxta ubertatem terrae suaedecoravit simulacra.
HOS|10|2|Divisum est cor eorum,nunc poenas solvent;ipse confringet aras eorum,depopulabitur simulacra eorum.
HOS|10|3|Profecto nunc dicent: Non est rex nobis;non enim timemus Dominum,et rex quid faciet nobis? ".
HOS|10|4|Loqui verba, iurare in vanum,ferire foedus;et germinabit quasi venenum iussuper sulcos agri.
HOS|10|5|De vitulo Bethaventrement habitatores Samariae;quia luget super eum populus eius;dum sacerdotes eius super eumexsultant in gloria eius;vere migrabit ab eo.
HOS|10|6|Siquidem et ipse in Assyriam delatus est,munus regi magno;confusio Ephraim capiet,et confundetur Israel in consilio suo.
HOS|10|7|Perit Samaria,rex eius quasi festuca super faciem aquae.
HOS|10|8|Et disperdentur excelsa impietatis,peccatum Israel;spina et tribulus ascendetsuper aras eorum,et dicent montibus: " Operite nos! "et collibus: " Cadite super nos! ".
HOS|10|9|Ex diebus Gabaa peccavit Israel;ibi perstiterunt.Non comprehendet eos in Gabaaproelium super filios iniquitatis?
HOS|10|10|" Iuxta desiderium meum corripiam eos;congregabuntur super eos populi,cum corripientur propter duas iniquitates suas.
HOS|10|11|Ephraim vitula docta,diligens trituram.Et ego transivi super pulchritudinem colli eius;iunxi Ephraim aratro,arabit Iudas,sarriet sibi Iacob.
HOS|10|12|Seminate vobis in iustitia,metite secundum caritatem;innovate vobis novale.Tempus est requirendi Dominum,donec veniat, ut pluat vobis iustitiam.
HOS|10|13|Arastis impietatem,iniquitatem messuistis,comedistis frugem mendacii,quia confisus es in curribus tuis,in multitudine fortium tuorum.
HOS|10|14|Consurget tumultus in populo tuo,et omnes munitiones tuae vastabuntur,sicut vastavit Salman Betharbeelin die proelii,matre super filios allisa.
HOS|10|15|Sic faciet vobis Bethelpropter maximam nequitiam vestram.Mane interibit rex Israel.
HOS|11|1|Cum puer esset Israel, dilexi eumet ex Aegypto vocavi filium meum.
HOS|11|2|Quanto magis vocabam eos,tanto recesserunt a facie mea;ipsi Baalim immolabantet simulacris sacrificabant.
HOS|11|3|Et ego dirigebam gressus Ephraim,portabam eos in brachiis meis,et nescierunt quod curarem eos.
HOS|11|4|In funiculis humanitatis trahebam eos,in vinculis caritatis;et fui eis, quasi qui elevant infantem ad maxillas suas,et declinavi ad eum, ut vesceretur.
HOS|11|5|Revertetur in terram Aegypti,et Assur ipse rex eius,quoniam noluerunt converti.
HOS|11|6|Saeviet gladius in civitatibus eiuset consumet garrulos eiuset comedet eos propter consilia eorum.
HOS|11|7|Populus meus pendet ad praevaricandum contra me;vocant eum ad altum, sed simul non erigunt eum.
HOS|11|8|Quomodo dabo te, Ephraim,tradam te, Israel?Quomodo dabo te sicut Adama,ponam te ut Seboim?Convertitur in me cor meum,simul exardescit miseratio mea.
HOS|11|9|Non faciam furorem irae meae,non convertar, ut disperdam Ephraim,quoniam Deus egoet non homo,in medio tui Sanctuset non veniam in terrore.
HOS|11|10|Post Dominum ambulabunt;quasi leo rugiet,quia ipse rugiet,et in tremore accurrent filii ab occidente.
HOS|11|11|Et avolabunt quasi avis ex Aegyptoet quasi columba de terra Assyriae;et collocabo eos in domibus suis,dicit Dominus.
HOS|12|1|Circumdedit me in fraude Ephraim,et in dolo domus Israel;C Iudas autem, dum adhuc vagatur, est cum Deoet cum Sancto fidelis " C.
HOS|12|2|Ephraim pascit ventumet sequitur aestum;tota die mendacium et violentiam multiplicatet foedus cum Assyriis initet oleum in Aegyptum fert.
HOS|12|3|Iudicium ergo Domini cum Iuda,et visitatio super Iacob;iuxta vias eius et iuxta opera eius reddet ei.
HOS|12|4|In utero supplantavit fratrem suumet in robore suo luctatus est cum Deo.
HOS|12|5|Et luctatus est cum angelo et praevaluit;flevit et deprecatus est eum.In Bethel invenit eumet ibi locutus est nobiscum
HOS|12|6|Dominus, Deus exercituum:Dominus memoriale eius.
HOS|12|7|" Et tu ad Deum tuum converteris;caritatem et iudicium custodiet spera in Deo tuo semper ".
HOS|12|8|Chanaan, in manu eius statera dolosa,fraudem diligit.
HOS|12|9|Et dixit Ephraim: " Verumtamen dives effectus sum,inveni opes mihi,omnes labores mei non invenient mihiiniquitatem, quam peccavi ".
HOS|12|10|" Ego autem Dominus, Deus tuusex terra Aegypti;adhuc sedere te faciam in tabernaculis,sicut in diebus conventus.
HOS|12|11|Et loquar ad prophetaset ego visionem multiplicaboet in manu prophetarum proponam similitudines ".
HOS|12|12|Si Galaad iniquitas fuerat,prorsus inanes facti sunt;in Galgala bobus immolantes,etiam altaria eorum erunt quasi acervisuper sulcos agri.
HOS|12|13|Fugit Iacob in regionem Aram;et servivit Israel pro uxoreet pro uxore custos fuit.
HOS|12|14|Per prophetam autem eduxit DominusIsrael de Aegypto,et per prophetam custoditus est.
HOS|12|15|Ad iracundiam provocavit Ephraim amarissime,sed sanguinem eius super eum relinquetet opprobrium eius retribuet ei Dominus suus.
HOS|13|1|Loquente Ephraim, horror factus est;dux erat in Israel.Et deliquit in Baalet mortuus est.
HOS|13|2|Et nunc addunt ad peccandumfaciuntque sibi conflatile de argento suo,secundum intellegentiam suam simulacra;factura artificum totum est. His - ipsi dicunt - immolate! ".Homines vitulos osculantur.
HOS|13|3|Idcirco erunt quasi nubes matutinaet sicut ros matutinus praeteriens,sicut palea turbine rapta ex areaet sicut fumus de fumario.
HOS|13|4|" Ego autem Dominus, Deus tuusex terra Aegypti;et Deum absque me nescies,et salvator non est praeter me.
HOS|13|5|Ego pavi te in deserto,in terra ardenti solitudinis.
HOS|13|6|Iuxta pascua sua saturati suntet saturati elevaverunt cor suum,propterea obliti sunt mei.
HOS|13|7|Et ego ero eis quasi leaena,sicut pardus iuxta viam insidiabor.
HOS|13|8|Occurram eis quasi ursa, raptis catulis,et dirumpam claustrum cordis eorum:et consumam eos ibi quasi leo;bestia agri scindet eos.
HOS|13|9|Perdo te, Israel;quis est auxiliator tuus?
HOS|13|10|Ubinam est rex tuus,ut salvet te in omnibus urbibus tuis,et iudices tui, de quibus dixisti:Da mihi regem et principes"?
HOS|13|11|Do tibi regem in furore meoet aufero in indignatione mea.
HOS|13|12|Colligata est iniquitas Ephraim,absconditum peccatum eius.
HOS|13|13|Dolores parturientis venient ei;erit filius non sapiens:suo enim tempore non stabitin ore vulvae.
HOS|13|14|De manu inferni liberabo eos,de morte redimam eos?Ubi pestilentiae tuae, o mors?Ubi pestis tua, inferne?Consolatio abscondita est ab oculis meis ".
HOS|13|15|Dum ipse inter fratres fructificat,veniet ventus urens, ventus Dominide deserto ascendens,et siccabit venas eiuset desolabit fontem eius.Ipse diripiet thesaurum,omne vas desiderabile.
HOS|14|1|Poenas solvet Samaria,quoniam rebellavit contra Deum suum:in gladio peribunt,parvuli eorum elidentur,et praegnantes discindentur.
HOS|14|2|Convertere, Israel, ad Dominum Deum tuum,quoniam corruisti in iniquitate tua.
HOS|14|3|Tollite vobiscum verbaet convertimini ad Dominum;dicite ei: " Omnem aufer iniquitatemet accipe bonum,et reddemus fructum labiorum nostrorum.
HOS|14|4|Assyria non salvabit nos;super equum non ascendemusnec vocabimus ultra: "Deos nostros!"opera manuum nostrarum,quia in te misericordiam consequetur pupillus ".
HOS|14|5|" Sanabo praevaricationem eorum,diligam eos spontanee,quia aversus est furor meus ab eis.
HOS|14|6|Ero quasi ros pro Israel;germinabit quasi liliumet mittet radices suas ut Libanus.
HOS|14|7|Expandentur rami eius;et erit quasi oliva gloria eius,et odor eius ut Libani.
HOS|14|8|Convertentur sedentes in umbra mea,colent triticumet germinabunt quasi vinea;memoriale eius sicut vinum Libani.
HOS|14|9|Ephraim, quid ei ultra idola?Ego exaudio et respicio in eum.Ego ut abies virens:ex me fructus tuus invenitur ".
HOS|14|10|Qui sapiens est, intellegat ista;intellegens sciat haec!Quia rectae viae Domini,et iusti ambulabunt in eis;praevaricatores vero corruent in eis.
