PHLM|1|1|Paulus vinctus Christi Iesu et Timotheus frater Philemoni dilecto et adiutori nostro
PHLM|1|2|et Apphiae sorori et Archippo commilitoni nostro et ecclesiae, quae in domo tua est:
PHLM|1|3|gratia vobis et pax a Deo Patre nostro et Domino Iesu Christo.
PHLM|1|4|Gratias ago Deo meo semper memoriam tui faciens in orationibus meis,
PHLM|1|5|audiens caritatem tuam et fidem, quam habes in Dominum Iesum et in omnes sanctos,
PHLM|1|6|ut communio fidei tuae evidens fiat in agnitione omnis boni, quod est in nobis in Christum;
PHLM|1|7|gaudium enim magnum habui et consolationem in caritate tua, quia viscera sanctorum requieverunt per te, frater.
PHLM|1|8|Propter quod multam fiduciam habens in Christo imperandi tibi, quod ad rem pertinet,
PHLM|1|9|propter caritatem magis obsecro, cum sim talis ut Paulus senex, nunc autem et vinctus Christi Iesu;
PHLM|1|10|obsecro te de meo filio, quem genui in vinculis, Onesimo,
PHLM|1|11|qui tibi aliquando inutilis fuit, nunc autem et tibi et mihi utilis,
PHLM|1|12|quem remisi tibi: eum, hoc est viscera mea;
PHLM|1|13|quem ego volueram mecum detinere, ut pro te mihi ministraret in vinculis evangelii.
PHLM|1|14|Sine consilio autem tuo nihil volui facere, uti ne velut ex necessitate bonum tuum esset sed voluntarium.
PHLM|1|15|Forsitan enim ideo discessit ad horam, ut aeternum illum reciperes,
PHLM|1|16|iam non ut servum sed plus servo, carissimum fratrem, maxime mihi, quanto autem magis tibi et in carne et in Domino.
PHLM|1|17|Si ergo habes me socium, suscipe illum sicut me.
PHLM|1|18|Si autem aliquid nocuit tibi aut debet, hoc mihi imputa.
PHLM|1|19|Ego Paulus scripsi mea manu, ego reddam; ut non dicam tibi quod et teipsum mihi debes.
PHLM|1|20|Ita, frater! Ego te fruar in Domino; refice viscera mea in Christo!
PHLM|1|21|Confidens oboedientia tua scripsi tibi, sciens quoniam et super id, quod dico, facies.
PHLM|1|22|Simul autem et para mihi hospitium, nam spero per orationes vestras donari me vobis.
PHLM|1|23|Salutat te Epaphras, concaptivus meus in Christo Iesu,
PHLM|1|24|Marcus, Aristarchus, Demas, Lucas, adiutores mei.
PHLM|1|25|Gratia Domini Iesu Christi cum spiritu vestro.
