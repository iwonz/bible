LAM|1|1|Як самітно сидить колись велелюдне це місто, немов удова воно стало! Могутнє посеред народів, княгиня посеред країн воно стало данницею!...
LAM|1|2|Гірко плаче по ночах вона, і сльози гарячі на щоках у неї... Нема потішителя в неї зо всіх, що кохали її, її зрадили всі її друзі, вони ворогами їй стали!
LAM|1|3|Юдея пішла на вигнання з біди та з роботи тяжкої, вона оселилася поміж поганами, спочинку собі не знайшла! Догнали її всі її переслідники серед тіснот...
LAM|1|4|Дороги сіонської доньки сумні, бо немає на свято прочан! Усі брами її попустіли, зідхає священство її, посумнілі дівчата її, а вона гірко їй!
LAM|1|5|Її грабівники взяли гору над нею, і добре ведеться її ворогам, бо їй завдав смутку Господь за численність у неї гріхів: Немовлята її до полону пішли перед ворогом...
LAM|1|6|І відійшла від сіонської доньки вся величність її... Її князі стали, немов олені ті, що паші собі не знаходять, і йдуть у безсиллі перед переслідником...
LAM|1|7|У дні лиха свого та страждання свого дочка єрусалимська спогадує всі свої скарби, що були від днів давніх, як народ її впав був у руку ворожу, і не було, хто б їй поміч подав... Вороги споглядали на неї, і сміялись з руїни її...
LAM|1|8|Дочка єрусалимська гріхом прогрішилась, тому то нечистою стала, усі, що її шанували, погорджують нею, наготу бо її вони бачили! І зідхає вона, й відвертається взад...
LAM|1|9|Нечистість її на подолках у неї. Вона не згадала свого кінця, та й упала предивно, і нікого нема, хто б потішив її... Побач, Господи, горе моє, бо звеличився ворог!
LAM|1|10|Гнобитель простяг свою руку на всі її скарби, і бачить вона, що в святиню її увіходять погани, про яких наказав Ти: Не ввійдуть вони в твої збори!
LAM|1|11|Увесь народ її стогне, шукаючи хліба, свої скарби коштовні за їжу дають, аби тільки душу свою проживити... Зглянься, Господи, і подивися, яка стала погорджена я!
LAM|1|12|Не вам кажучи, гляньте й побачте, усі, хто дорогою йде: чи є такий біль, як мій біль, що завданий мені, що Господь засмутив ним мене у день лютого гніву Свого?...
LAM|1|13|Із височини Він послав в мої кості огонь, і над ними він запанував! Розтяг сітку на ноги мої, повернув мене взад, учинив Він мене спустошілою, увесь день болящою...
LAM|1|14|Ярмо моїх прогріхів зв'язане міцно рукою Його, плетуться вони та приходять на шию мою! Він зробив, що спіткнулася сила моя, Господь передав мене в руки такого, що й звестись не можу...
LAM|1|15|Усіх моїх сильних Господь поскидав серед мене, мов на свято зібрання, Він скликав на мене, щоб моїх юнаків поторощити, як у чавилі, стоптав Господь дівчину, Юдину доньку...
LAM|1|16|За оцим плачу я, око моє, моє око слізьми запливає! бо далеко від мене втішитель, що душу мою оживив би; мої діти понехтувані, бо посилився ворог!
LAM|1|17|Сіонська дочка простягла свої руки, немає розрадника їй: Господь наказав проти Якова довкола нього його ворогам, донька єрусалимська нечистою стала між ними...
LAM|1|18|Справедливий Господь, а я слову Його неслухняна була... Послухайте но, всі народи, і побачте мій біль: дівчата мої та мої юнаки у неволю пішли!
LAM|1|19|Взивала до друзів своїх, та вони обманули мене! Священство моє й мої старші вмирають у місті, шукаючи їжі собі, щоб душу свою поживити...
LAM|1|20|Зглянься, Господи, тісно мені! Моє нутро бентежиться, перевертається серце моє у мені, бо була зовсім неслухняна... На вулиці меч осирочував, а в домі смерть...
LAM|1|21|Почули, що я ось стогну, й немає мені потішителя, вчули про лихо моє всі мої вороги, та й зраділи, що Ти це зробив... Спровадив Ти день, що його заповів, бодай сталося їм, як мені!
LAM|1|22|Бодай перед обличчя Твоє прийшло все їхнє лихо, і вчини їм, як Ти учинив ось мені за гріхи мої всі, бо численні стогнання мої, моє ж серце боляще...
LAM|2|1|Як захмарив Господь в Своїм гніві сіонську дочку! Він кинув із неба на землю пишноту Ізраїля, і не згадав у день гніву Свого про підніжка ногам Своїм,
LAM|2|2|понищив Господь, не помилував житла всі Яковові... Він позбурював у гніві Своїм у дочки Юди твердині, на землю звалив, збезчестив Він царство й князів усіх його...
LAM|2|3|В люті гніву відтяв увесь Ізраїлів ріг, правицю Свою відвернув Він від ворога, та й запалав проти Якова, мов той палючий огонь, що навколо жере!
LAM|2|4|Він нап'яв Свого лука, як ворог, противником стала правиця Його, і Він вибив усе, що для ока було пожадане, у скинії доньки сіонської вилив запеклість Свою, як огонь...
LAM|2|5|Господь став, як той ворог, понищив Ізраїля Він, всі палати його зруйнував, твердині його попустошив, і Юдиній доньці примножив зідхання та стогін!
LAM|2|6|Понищив горожу Свою, немов у садка, місце зборів Своїх попустошив, Господь учинив, що забули в Сіоні про свято й суботу, і відкинув царя та священика в лютості гніву Свого...
LAM|2|7|Покинув Господь Свого жертівника, допустив побезчестити святиню Свою, передав в руку ворога мури палаців її, вороги зашуміли в Господньому домі, немов би святкового дня!
LAM|2|8|Задумав Господь зруйнувати мур сіонської доньки, Він витягнув шнура, Своєї руки не вернув, щоб не нищити, сумними вчинив передмур'я та мур, вони разом ослабли...
LAM|2|9|Її брами запалися в землю, понищив Він та поламав її засуви... Її цар і князі її серед поганів... Немає навчання Закону, і пророки її не знаходять видіння від Господа...
LAM|2|10|Сидять на землі та мовчать старші доньки сіонської, порох посипали на свою голову, підперезались веретами, аж до землі свою голову єрусалимські дівчата схилили...
LAM|2|11|Повипливали від сліз мої очі, моє нутро клекоче, на землю печінка моя виливається через занепад дочки мого люду, коли немовля й сосунець умлівають голодні на площах міських.
LAM|2|12|Вони квилять своїм матерям: Де пожива й вино? І скулюються, як ранений, на площах міських, коли душі свої випускають на лоні своїх матерів...
LAM|2|13|Що засвідчу тобі, що вподоблю до тебе, о єрусалимськая дочко? Що вчиню тобі рівним, щоб тебе звеселити, о діво, о дочко сіонська? Бо велика, як море, руїна твоя, хто тебе полікує?
LAM|2|14|Пророки твої провіщали для тебе марноту й фальшиве, і не відкривали твого гріха, щоб долю твою відвернути, для тебе вбачали пророцтва марноти й вигнання...
LAM|2|15|Усі, що проходять дорогою, плещуть у долоні на тебе, і посвистують та головою своєю хитають над донькою Єрусалиму та кажуть: Хіба це те місто, що про нього казали: Корона пишноти, розрада всієї землі?
LAM|2|16|Усі вороги твої пащу на тебе роззявлюють, свищуть й зубами скрегочуть та кажуть: Ми пожерли її... Оце справді той день, що чекали його, знайшли ми і бачимо його!...
LAM|2|17|Учинив Господь те, що задумав, Він виповнив слово Своє, що його наказав від днів давніх: усе зруйнував, і милосердя не мав, і ворога втішив тобою, Він рога підійняв супротивних твоїх...
LAM|2|18|Їхнє серце до Господа крик підіймає, о муре, о дочко Сіону! Проливай, як потік, сльози вдень та вночі, не давай відпочинку собі, нехай не спочине зіниця твоя!
LAM|2|19|Уставай, голоси уночі на початку сторожі! Виливай своє серце, мов воду, навпроти обличчя Господнього! Підійми ти до Нього долоні свої за душу своїх немовлят, що від голоду мліють на розі всіх вулиць!...
LAM|2|20|Споглянь, Господи, і подивися, кому Ти зробив отаке? Чи конечним було, щоб жінки їли плід свій, своїх немовлят, яких виплекали? Щоб був у святині Господній забитий священик і пророк?
LAM|2|21|Лежать на землі на вулицях рядом юнак та старий... Попадали діви мої та мої парубки від меча, Ти побив їх в день гніву Свого, порізав, не мав милосердя...
LAM|2|22|Ти викликував, мов на день свята, жахоти мої із довкілля, і врятованого не було, і позостальця в день гніву Господнього, повигублював ворог мій тих, кого виплекала та зростила була...
LAM|3|1|Я той муж, який бачив біду від жезла Його гніву,
LAM|3|2|Він провадив мене й допровадив до темряви, а не до світла...
LAM|3|3|Лиш на мене все знову обертає руку Свою цілий день...
LAM|3|4|Він виснажив тіло моє й мою шкіру, мої кості сторощив,
LAM|3|5|обгородив Він мене, і мене оточив гіркотою та мукою,
LAM|3|6|у темноті мене посадив, мов померлих давно...
LAM|3|7|Обгородив Він мене і не вийду, тяжкими вчинив Він кайдани мої...
LAM|3|8|І коли я кричу й голошу, затикає Він вуха Свої на молитву мою...
LAM|3|9|Камінням обтесаним обгородив Він дороги мої, повикривлював стежки мої...
LAM|3|10|Він для мене ведмедем чатуючим став, немов лев той у сховищі!
LAM|3|11|Поплутав дороги мої та розшарпав мене, учинив Він мене опустошеним!
LAM|3|12|Натягнув Свого лука й поставив мене, наче ціль для стріли,
LAM|3|13|пустив стріли до нирок моїх з Свого сагайдака...
LAM|3|14|Для всього народу свого я став посміховиськом, глумливою піснею їхньою цілий день...
LAM|3|15|Наситив мене гіркотою, мене напоїв полином...
LAM|3|16|І стер мені зуби жорствою, до попелу кинув мене,
LAM|3|17|і душа моя спокій згубила, забув я добро...
LAM|3|18|І сказав я: Загублена сила моя, та моє сподівання на Господа...
LAM|3|19|Згадай про біду мою й муку мою, про полин та отруту,
LAM|3|20|душа моя згадує безперестанку про це, і гнеться в мені...
LAM|3|21|Оце я нагадую серцеві своєму, тому то я маю надію:
LAM|3|22|Це милість Господня, що ми не погинули, бо не покінчилось Його милосердя,
LAM|3|23|нове воно кожного ранку, велика бо вірність Твоя!
LAM|3|24|Господь це мій уділ, говорить душа моя, тому я надію на Нього складаю!
LAM|3|25|Господь добрий для тих, хто надію на Нього кладе, для душі, що шукає Його!
LAM|3|26|Добре, коли людина в мовчанні надію кладе на спасіння Господнє.
LAM|3|27|Добре для мужа, як носить ярмо в своїй молодості,
LAM|3|28|нехай він самітно сидить і мовчить, як поклав Він на нього його;
LAM|3|29|хай закриє він порохом уста свої, може є ще надія;
LAM|3|30|хай щоку тому підставляє, хто його б'є, своєю ганьбою насичується...
LAM|3|31|Бо Господь не навіки ж покине!
LAM|3|32|Бо хоч Він і засмутить кого, проте змилується за Своєю великою милістю,
LAM|3|33|бо не мучить Він з серця Свого, і не засмучує людських синів.
LAM|3|34|Щоб топтати під своїми ногами всіх в'язнів землі,
LAM|3|35|щоб перед обличчям Всевишнього право людини зігнути,
LAM|3|36|щоб гнобити людину у справі судовій його, оцього не має на оці Господь!
LAM|3|37|Хто то скаже і станеться це, як Господь того не наказав?
LAM|3|38|Хіба не виходить усе з уст Всевишнього, зле та добре?
LAM|3|39|Чого ж нарікає людина жива? Нехай скаржиться кожен на гріх свій.
LAM|3|40|Пошукаймо доріг своїх та дослідімо, і вернімось до Господа!
LAM|3|41|підіймімо своє серце та руки до Бога на небі!
LAM|3|42|Спроневірились ми й неслухняними стали, тому не пробачив Ти нам,
LAM|3|43|закрився Ти гнівом і гнав нас, убивав, не помилував,
LAM|3|44|закрив Себе хмарою, щоб до Тебе молитва моя не дійшла...
LAM|3|45|Сміттям та огидою нас Ти вчинив між народами,
LAM|3|46|наші всі вороги пороззявляли на нас свого рота,
LAM|3|47|страх та яма на нас поприходили, руїна й погибіль...
LAM|3|48|Моє око спливає потоками водними через нещастя дочки мого люду...
LAM|3|49|Виливається око моє безупинно, нема бо перерви,
LAM|3|50|аж поки не зглянеться та не побачить Господь із небес,
LAM|3|51|моє око вчиняє журбу для моєї душі через дочок усіх мого міста...
LAM|3|52|Ловлячи, ловлять мене, немов птаха, мої вороги безпричинно,
LAM|3|53|життя моє в яму замкнули вони, і каміннями кинули в мене...
LAM|3|54|Пливуть мені води на голову, я говорю: Вже погублений я!...
LAM|3|55|Кликав я, Господи, Ймення Твоє із найглибшої ями,
LAM|3|56|Ти чуєш мій голос, не заховуй же вуха Свого від зойку мого, від благання мого!
LAM|3|57|Ти близький того дня, коли кличу Тебе, Ти говориш: Не бійся!
LAM|3|58|За душу мою Ти змагався, о Господи, життя моє викупив Ти.
LAM|3|59|Ти бачиш, о Господи, кривду мою, розсуди ж Ти мій суд!
LAM|3|60|Усю їхню помсту Ти бачиш, всі задуми їхні на мене,
LAM|3|61|Ти чуєш, о Господи, їхні наруги, всі задуми їхні на мене,
LAM|3|62|мову повстанців на мене та їхнє буркотіння на мене ввесь день...
LAM|3|63|Побач їхнє сидіння та їхнє вставання, як завжди глумлива їхня пісня!
LAM|3|64|Заплати їм, о Господи, згідно з чином їхніх рук!
LAM|3|65|Подай їм темноту на серце, прокляття Твоє нехай буде на них!
LAM|3|66|Своїм гнівом жени їх, і вигуби їх з-під Господніх небес!
LAM|4|1|Як потемніло золото, як відмінилося щире те золото добре, як на розі всіх вулиць каміння святе порозкидане!
LAM|4|2|Коштовні сіонські сини, щирим золотом важені, як тепер ось за глиняний посуд полічені, за чин рук ганчарських!
LAM|4|3|Навіть шакали витягують перса, годують своїх молодят, а доня народу мого жорстока, мов струсі в пустині:
LAM|4|4|язик сосунця до його піднебіння від спраги прилип... Хліба жадають собі немовлята, й немає нікого, хто б їм відломив...
LAM|4|5|Ті, що їли присмаки, на вулицях з голоду мліють; ті, що виплекані на пурпурі, тепер смітники обіймають...
LAM|4|6|І більшою стала вина доньки люду мого за прогріх Содому, що був перевернений вмить, і не торкалися руки до нього...
LAM|4|7|Її можновладці чистіші від снігу були, біліші від молока, їхнє тіло червоне, мов перли, їхній вигляд сапфір,
LAM|4|8|а тепер їхній вигляд чорніший за сажу, не розпізнають їх на вулицях, їхня шкіра стягнулась на їхній кості, зробилась сухою, як дерево...
LAM|4|9|Забитим мечем стало ліпше, ніж повбиваним голодом, що гинуть проколені, за браком плодів польових...
LAM|4|10|Руки жінок милосердних варили своїх діточок, які стали поживою їм під час руйнування дочки мого люду...
LAM|4|11|Закінчив Господь лютість Свою, вилив жар Свого гніву, і запалив на Сіоні огонь, і пожер він основи його!
LAM|4|12|Не вірили земні царі та всі мешканці цілого світу, що ввійде противник та ворог до брам Єрусалиму...
LAM|4|13|Усе сталося це за провини пророків його, за неправду священства його, що кров праведників серед нього лили...
LAM|4|14|По вулицях бродять, немов ті сліпці, поплямовані кров'ю, так що люди не можуть діткнутись до одягу їхнього.
LAM|4|15|Уступіться, нечисті! кричали до них, уступіться, збочуйте, не доторкуйтеся!... І повтікали вони й мандрували, і казали між людьми: Мешкати в нас більш не будуть!
LAM|4|16|Господнє лице розпорошило їх, не дивиться більше на них, бо вони не звертали уваги на обличчя священиків, до старих вони ласки не мали...
LAM|4|17|Уже прогляділи ми очі свої, даремно чекавши на поміч собі, на варті своїй ми чекали народу, який нас не спас...
LAM|4|18|Чатують вони наші кроки, щоб ходити не могли ми по площах своїх. Кінець наш наблизився, сповнилися наші дні, бо прийшов нам кінець...
LAM|4|19|Гнобителі наші скоріші були за орлів піднебесних, вони уганялись за нами по горах, на нас чатували в пустині...
LAM|4|20|Попав в ями живущий наш дух, Господній помазанець, що ми говорили про нього: Ми будемо жити в тіні його серед народів.
LAM|4|21|Веселися та тішся, о дочко Едому, що сидиш в краю Уц, також над тобою перейде злий келіх, уп'єшся й оголишся й ти!
LAM|4|22|Скінчилася кара твоя, дочко Сіону, не буде Він більше тебе виганяти, та твоє беззаконня скарає Він, дочко Едому, відкриє провини твої!
LAM|5|1|Згадай, Господи, що з нами сталося, зглянься й побач нашу ганьбу,
LAM|5|2|наша спадщина дісталась чужим, доми наші чужинцям!
LAM|5|3|Поставали ми сиротами: нема батька, а матінки наші неначе ті вдови!...
LAM|5|4|Свою воду за срібло ми п'ємо, наші дрова за гроші одержуємо...
LAM|5|5|У потилицю нас поганяють, помучені ми, і спокою не маємо!
LAM|5|6|До Єгипту й Асирії руку витягуємо, щоб насититись хлібом!
LAM|5|7|Батьки наші грішили, але їх нема, а ми двигаємо їхні провини!
LAM|5|8|Раби запанували над нами, і немає нікого, хто б вирятував з їхньої руки...
LAM|5|9|Наражуючи свою душу на меч у пустині, достаємо свій хліб...
LAM|5|10|Шкіра наша, мов піч, попалилась з пекучого голоду...
LAM|5|11|Жінок на Сіоні безчестили, дівчат по Юдейських містах...
LAM|5|12|Князі їхньою рукою повішені, лиця старих не пошановані...
LAM|5|13|Юнаки носять камінь млиновий, а хлопці під ношею дров спотикаються...
LAM|5|14|Перестали сидіти старші в брамі, юнаки свою пісню співати,
LAM|5|15|втіха нашого серця спинилась, наш танець змінивсь на жалобу...
LAM|5|16|Спала корона у нас з голови, о горе, бо ми прогрішились,
LAM|5|17|тому наше серце боляще, тому наші очі потемніли,
LAM|5|18|через гору Сіон, що спустошена, бродять лисиці по ній...
LAM|5|19|Пробуваєш Ти, Господи, вічно, Твій престол з роду в рід:
LAM|5|20|Нащо ж нас забуваєш навік, покидаєш на довгі дні нас?
LAM|5|21|Приверни нас до Себе, о Господи, і вернемось ми, віднови наші дні, як давніше було!
LAM|5|22|Хіба Ти цілком нас відкинув, прогнівавсь занадто на нас?...
