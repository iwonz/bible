DEUT|1|1|Haec sunt verba, quae locutus est Moyses ad omnem Israel trans Iordanem in solitudine, in Araba contra Suph, inter Pharan et Thophel et Laban et Aseroth et Dizahab.
DEUT|1|2|Undecim dies de Horeb per viam montis Seir usque Cadesbarne.
DEUT|1|3|Quadragesimo anno, undecimo mense, prima die mensis locutus est Moyses ad filios Israel omnia, quae praeceperat illi Dominus ut diceret eis.
DEUT|1|4|Postquam percussit Sehon regem Amorraeorum, qui habitavit in Hesebon, et Og regem Basan, qui mansit in Astharoth et in Edrai,
DEUT|1|5|trans Iordanem in terra Moab coepitque Moyses explanare legem hanc et dicere:
DEUT|1|6|" Dominus Deus noster locutus est ad nos in Horeb dicens: "Sufficit vobis quod in hoc monte mansistis;
DEUT|1|7|convertimini et proficiscimini et venite ad montem Amorraeorum et ad omnes vicinos eius: in Araba atque montanis et in Sephela et in Nageb et iuxta litus maris, in terram Chananaeorum et in Libanum usque ad flumen magnum Euphraten.
DEUT|1|8|En, inquit, tradidi vobis terram: ingredimini et possidete eam, super qua iuravit Dominus patribus vestris, Abraham, Isaac et Iacob, ut daret illam eis et semini eorum post eos".
DEUT|1|9|Dixique vobis illo in tempore: Non possum solus sustinere vos;
DEUT|1|10|Dominus Deus vester multiplicavit vos, et estis hodie sicut stellae caeli plurimi.
DEUT|1|11|Dominus, Deus patrum vestrorum, addat ad hunc numerum multa milia et benedicat vobis, sicut locutus est vobis.
DEUT|1|12|Non valeo solus vestra negotia sustinere et pondus ac iurgia;
DEUT|1|13|date vobis viros sapientes et gnaros, et quorum conversatio sit probata in tribubus vestris, ut ponam eos vobis principes.
DEUT|1|14|Tunc respondistis mihi: "Bona res est, quam vis facere".
DEUT|1|15|Tulique principes de tribubus vestris viros sapientes et probatos et constitui eos principes super vos: tribunos et centuriones et quinquagenarios ac decanos et praefectos operum pro tribubus vestris.
DEUT|1|16|Praecepique iudicibus vestris in tempore illo: Audite causam fratrum vestrorum et, quod iustum est, iudicate, sive civis sit ille sive peregrinus.
DEUT|1|17|Non accipietis personam in iudicio; ita parvum audietis ut magnum nec timebitis cuiusquam personam, quia Dei iudicium est. Quod si difficile vobis aliquid visum fuerit, referte ad me, et ego audiam.
DEUT|1|18|Praecepique vobis in tempore illo omnia, quae facere deberetis.
DEUT|1|19|Profecti autem de Horeb transivimus per totam illam eremum maximam et terribilem, quam vidistis, per viam montis Amorraei, sicut praeceperat Dominus Deus noster nobis. Cumque venissemus in Cadesbarne,
DEUT|1|20|dixi vobis: Venistis ad montem Amorraei, quem Dominus Deus noster daturus est nobis.
DEUT|1|21|Vide terram, quam Dominus Deus tuus dat tibi: ascende et posside eam, sicut locutus est tibi Dominus, Deus patrum tuorum; noli metuere nec quidquam paveas.
DEUT|1|22|Et accessistis ad me vos omnes atque dixistis: "Mittamus viros ante nos, qui considerent terram et renuntient de itinere, per quod debeamus ascendere, et de civitatibus, ad quas pergere".
DEUT|1|23|Cumque mihi sermo placuisset, misi ex vobis duodecim viros singulos de tribubus suis.
DEUT|1|24|Qui cum perrexissent et ascendissent in montana, venerunt usque ad Nehelescol et, considerata terra,
DEUT|1|25|sumentes de fructibus eius attulerunt ad nos atque dixerunt: "Bona est terra, quam Dominus Deus noster daturus est nobis".
DEUT|1|26|Et noluistis ascendere, sed increduli ad sermonem Domini Dei vestri
DEUT|1|27|murmurastis in tabernaculis vestris atque dixistis: "Odit nos Dominus et idcirco eduxit nos de terra Aegypti, ut traderet nos in manu Amorraei atque deleret.
DEUT|1|28|Quo ascendemus? Fratres nostri terruerunt cor nostrum dicentes: Maxima multitudo est et nobis in statura procerior; urbes magnae et ad caelum usque munitae; etiam filios Enacim vidimus ibi".
DEUT|1|29|Et dixi vobis: Nolite metuere nec timeatis eos.
DEUT|1|30|Dominus Deus, qui ductor est vester, ipse pro vobis pugnabit, sicut fecit in Aegypto, vobis videntibus.
DEUT|1|31|Et in solitudine - ipse vidisti - portavit te Dominus Deus tuus, ut solet homo gestare parvulum filium suum, in omni via, per quam ambulastis, donec veniretis ad locum istum.
DEUT|1|32|Et nec sic quidem credidistis Domino Deo vestro,
DEUT|1|33|qui praecessit vos in via, et metatus est locum, in quo tentoria figere deberetis, nocte ostendens vobis iter per ignem et die per columnam nubis.
DEUT|1|34|Cumque audisset Dominus vocem sermonum vestrorum, iratus iuravit et ait:
DEUT|1|35|"Non videbit quispiam de viris generationis huius pessimae terram bonam, quam sub iuramento pollicitus sum patribus vestris,
DEUT|1|36|praeter Chaleb filium Iephonne: ipse enim videbit eam, et ipsi dabo terram, quam calcavit, et filiis eius, quia adimplevit ut sequeretur Dominum".
DEUT|1|37|Mihi quoque iratus Dominus propter vos dixit: "Nec tu ingredieris illuc;
DEUT|1|38|sed Iosue filius Nun minister tuus ipse intrabit illuc. Hunc robora, et ipse terram sorte dividat Israeli.
DEUT|1|39|Parvuli vestri, de quibus dixistis quod captivi ducerentur, et filii, qui hodie boni ac mali ignorant distantiam, ipsi ingredientur; et ipsis dabo terram, et possidebunt eam.
DEUT|1|40|Vos autem revertimini et abite in solitudinem per viam maris Rubri".
DEUT|1|41|Et respondistis mihi: "Peccavimus Domino; nos ascendemus atque pugnabimus, sicut praecepit nobis Dominus Deus noster". Cumque instructi armis pergeretis in montem,
DEUT|1|42|ait mihi Dominus: "Dic ad eos: Nolite ascendere neque pugnetis, non enim sum vobiscum, ne cadatis coram inimicis vestris".
DEUT|1|43|Locutus sum, et non audistis, sed adversantes imperio Domini et tumentes superbia ascendistis in montem.
DEUT|1|44|Itaque egressus Amorraeus, qui habitat in monte illo, obviam vobis, persecutus est vos, sicut solent apes persequi, et cecidit vos de Seir usque Horma.
DEUT|1|45|Cumque reversi ploraretis coram Domino, non audivit vos nec voci vestrae voluit acquiescere.
DEUT|1|46|Sedistis ergo in Cades multo illo tempore, dum ibi mansistis.
DEUT|2|1|Profectique inde venimus in solitudinem per viam maris Ru bri, sicut mihi dixerat Dominus; et circuivimus montem Seir longo tempore.
DEUT|2|2|Dixitque Dominus ad me:
DEUT|2|3|"Sufficit vobis circuire montem istum; ite contra aquilonem.
DEUT|2|4|Et populo praecipe dicens: Transibitis per terminos fratrum vestrorum filiorum Esau, qui habitant in Seir, et timebunt vos.
DEUT|2|5|Cavete ergo diligenter, ne moveamini contra eos; neque enim dabo vobis de terra eorum, quantum potest unius pedis calcare vestigium, quia in possessionem Esau dedi montem Seir.
DEUT|2|6|Cibos emetis ab eis pecunia et comedetis; etiam aquam emptam haurietis et bibetis.
DEUT|2|7|Dominus Deus tuus benedixit tibi in omni opere manuum tuarum; novit iter tuum, quomodo transieris solitudinem hanc magnam per quadraginta annos habitans tecum Dominus Deus tuus, et nihil tibi defuit".
DEUT|2|8|Cumque transissemus fratres nostros filios Esau, qui habitabant in Seir, per viam Arabae de Ailath et de Asiongaber, vertimus nos et venimus per iter, quod ducit in desertum Moab.
DEUT|2|9|Dixitque Dominus ad me: "Non pugnes contra Moabitas nec ineas adversus eos proelium; non enim dabo tibi quidquam de terra eorum, quia filiis Lot tradidi Ar in possessionem.
DEUT|2|10|- Emim primi fuerunt habitatores eius, populus magnus et multus et tam excelsus ut Enacim;
DEUT|2|11|ipsi quoque Raphaim reputabantur sicut Enacim; denique Moabitae appellant eos Emim.
DEUT|2|12|In Seir autem prius habitaverunt Horim; quibus expulsis atque deletis, habitaverunt filii Esau pro eis, sicut fecit Israel in terra possessionis suae, quam dedit eis Dominus C.
DEUT|2|13|Surgite ergo et transite torrentem Zared". Et transivimus torrentem Zared.
DEUT|2|14|Tempus autem, quo ambulavimus de Cadesbarne usque ad transitum torrentis Zared, triginta octo annorum fuit, donec consumeretur omnis generatio hominum bellatorum de castris, sicut iuraverat eis Dominus,
DEUT|2|15|cuius manus fuit adversum eos, ut interirent de castrorum medio.
DEUT|2|16|Postquam autem universi ceciderunt pugnatores de medio populi,
DEUT|2|17|locutus est Dominus ad me dicens:
DEUT|2|18|"Tu transibis hodie terminos Moab, urbem nomine Ar;
DEUT|2|19|et accedens in vicina filiorum Ammon, cave, ne pugnes contra eos nec movearis ad proelium; non enim dabo tibi de terra filiorum Ammon, quia filiis Lot dedi eam in possessionem.
DEUT|2|20|- Terra Raphaim reputata est et ipsa olim habitaverunt Raphaim in ea, quos Ammonitae vocant Zomzommim,
DEUT|2|21|populus magnus et multus et procerae longitudinis sicut Enacim, quos delevit Dominus a facie eorum et fecit illos habitare pro eis,
DEUT|2|22|sicut fecerat filiis Esau, qui habitant in Seir, delens Horim et terram eorum illis tradens, quam possident usque in praesens.
DEUT|2|23|Hevaeos quoque, qui habitabant in villis usque Gazam, Caphtorim, qui egressi de Caphtor deleverunt eos et habitaverunt pro illis C.
DEUT|2|24|Surgite! Proficiscimini et transite torrentem Arnon: ecce tradidi in manu tua Sehon regem Hesebon Amorraeum; et terram eius incipe possidere et committe adversus eum proelium.
DEUT|2|25|Hodie incipiam mittere terrorem atque formidinem tuam in populos, qui habitant sub omni caelo, ut, audito nomine tuo, paveant et contremiscant coram te".
DEUT|2|26|Misi ergo nuntios de solitudine Cademoth ad Sehon regem Hesebon verbis pacificis dicens:
DEUT|2|27|Transibo per terram tuam, publica gradiar via, non declinabo neque ad dexteram neque ad sinistram;
DEUT|2|28|alimenta pretio vende mihi, ut vescar, aquam pecunia tribue mihi, et sic bibam; tantum est ut mihi concedas transitum,
DEUT|2|29|sicut fecerunt mihi filii Esau, qui habitant in Seir, et Moabitae, qui morantur in Ar, donec veniam ad Iordanem et transeam in terram, quam Dominus Deus noster daturus est nobis.
DEUT|2|30|Noluitque Sehon rex Hesebon dare nobis transitum, quia induraverat Dominus Deus tuus spiritum eius et obfirmaverat cor illius, ut traderetur in manus tuas, sicut est in praesenti die.
DEUT|2|31|Dixitque Dominus ad me: "Ecce coepi tradere tibi Sehon et terram eius. Incipe possidere eam!".
DEUT|2|32|Egressusque est Sehon obviam nobis cum omni populo suo ad proelium in Iasa,
DEUT|2|33|et tradidit eum Dominus Deus noster nobis; percussimusque eum cum filiis suis et omni populo suo.
DEUT|2|34|Cunctasque urbes eius in tempore illo cepimus et percussimus anathemate singulas civitates cum viris ac mulieribus et parvulis; neminem reliquimus in eis superstitem,
DEUT|2|35|absque iumentis, quae in partem venere praedantium, et spoliis urbium, quas cepimus.
DEUT|2|36|Ab Aroer, quae est super ripam torrentis Arnon, et oppido, quod in valle situm est, usque Galaad non fuit civitas, quae nostras effugeret manus: omnia tradidit Dominus Deus noster nobis,
DEUT|2|37|absque terra filiorum Ammon, ad quam non accessisti, cunctis, quae adiacent torrenti Iaboc, et urbibus montanis universisque locis, a quibus nos prohibuit Dominus Deus noster.
DEUT|3|1|Itaque conversi ascendimus per iter Basan; egressusque est Og rex Basan in occursum nobis cum omni populo suo ad bellandum in Edrai.
DEUT|3|2|Dixitque Dominus ad me: "Ne timeas eum, quia in manu tua tradidi eum cum omni populo ac terra sua; faciesque ei, sicut fecisti Sehon regi Amorraeorum, qui habitavit in Hesebon".
DEUT|3|3|Tradidit ergo Dominus Deus noster in manibus nostris etiam Og regem Basan et universum populum eius; percussimusque eos usque ad internecionem.
DEUT|3|4|Et cepimus cunctas civitates eius in illo tempore. Non fuit oppidum, quod nos effugeret: sexaginta urbes, omnem regionem Argob, regnum Og in Basan.
DEUT|3|5|Cunctae urbes erant munitae muris altissimis portisque et vectibus, absque oppidis innumeris, quae non habebant muros.
DEUT|3|6|Et percussimus eos anathemate, sicut feceramus Sehon regi Hesebon, disperdentes omnem civitatem virosque ac mulieres et parvulos;
DEUT|3|7|iumenta autem et spolia urbium diripuimus.
DEUT|3|8|Tulimusque illo in tempore terram de manu duorum regum Amorraeorum, qui erant trans Iordanem, a torrente Arnon usque ad montem Hermon
DEUT|3|9|- Sidonii vocant Hermon Sarion et Amorraei Sanir -
DEUT|3|10|omnes civitates, quae sitae sunt in planitie, et universam terram Galaad et Basan usque Salcha et Edrai, civitates regni Og in Basan.
DEUT|3|11|- Solus quippe Og rex Basan remanserat de residuis Raphaim. Monstratur lectus eius ferreus. Nonne est in Rabba filiorum Ammon? Novem cubitos habet longitudinis et quattuor latitudinis ad mensuram cubiti virilis manus C.
DEUT|3|12|Terramque hanc possedimus in tempore illo ab Aroer, quae est super ripam torrentis Arnon, usque ad mediam partem montis Galaad; et civitates illius dedi Ruben et Gad.
DEUT|3|13|Reliquam autem partem Galaad et omnem Basan, regnum Og, tradidi mediae tribui Manasse, omnem regionem Argob. Cuncta Basan vocatur terra Raphaim.
DEUT|3|14|Iair filius Manasse possedit omnem regionem Argob usque ad terminos Gesuri et Maachathi; vocavitque ea ex nomine suo Basan Havoth Iair (id est villas Iair) usque in praesentem diem.
DEUT|3|15|Machir quoque dedi Galaad.
DEUT|3|16|Et tribubus Ruben et Gad dedi de terra Galaad usque ad torrentem Arnon, medium torrentis et confinium usque ad torrentem Iaboc, qui est terminus filiorum Ammon;
DEUT|3|17|et Arabam atque Iordanem et terminos a Chenereth usque ad mare Arabae, quod est mare Salis, ad radices montis Phasga contra orientem.
DEUT|3|18|Praecepique vobis in tempore illo dicens: Dominus Deus vester dedit vobis terram hanc in hereditatem; expediti praecedite fratres vestros filios Israel, omnes viri robusti,
DEUT|3|19|absque uxoribus et parvulis ac iumentis. Novi enim quod plura habeatis pecora, et in urbibus remanere debebunt, quas tradidi vobis,
DEUT|3|20|donec requiem tribuat Dominus fratribus vestris, sicut vobis tribuit, et possideant etiam ipsi terram, quam Dominus Deus vester daturus est eis trans Iordanem; tunc revertetur unusquisque in possessionem suam, quam dedi vobis.
DEUT|3|21|Iosue quoque in tempore illo praecepi dicens: Oculi tui viderunt, quae fecit Dominus Deus vester duobus his regibus; sic faciet omnibus regnis, ad quae transiturus es.
DEUT|3|22|Ne timeas eos: Dominus enim Deus vester pugnabit pro vobis.
DEUT|3|23|Precatusque sum Dominum in tempore illo dicens:
DEUT|3|24|Domine Deus, tu coepisti ostendere servo tuo magnitudinem tuam manumque fortissimam; neque enim est alius Deus vel in caelo vel in terra, qui possit facere opera tua et comparari fortitudini tuae.
DEUT|3|25|Transeam igitur et videam terram hanc optimam trans Iordanem et montem istum egregium et Libanum.
DEUT|3|26|Iratusque est Dominus mihi propter vos nec exaudivit me, sed dixit mihi: "Sufficit tibi; nequaquam ultra loquaris de hac re ad me.
DEUT|3|27|Ascende cacumen Phasgae et oculos tuos circumfer ad occidentem et aquilonem austrumque et orientem et aspice; nec enim transibis Iordanem istum.
DEUT|3|28|Praecipe Iosue et corrobora eum atque conforta, quia ipse praecedet populum istum et dividet eis terram, quam visurus es".
DEUT|3|29|Mansimusque in valle contra Bethphegor.
DEUT|4|1|Et nunc, Israel, audi praecepta et iudicia, quae ego doceo vos, ut facientes ea vivatis et ingredientes possideatis terram, quam Dominus, Deus patrum vestrorum, daturus est vobis.
DEUT|4|2|Non addetis ad verbum, quod vobis loquor, neque auferetis ex eo; custodite mandata Domini Dei vestri, quae ego praecipio vobis.
DEUT|4|3|Oculi vestri viderunt omnia, quae fecit Dominus contra Baalphegor, quomodo contriverit omnes cultores eius de medio vestri;
DEUT|4|4|vos autem, qui adhaeretis Domino Deo vestro, vivitis universi usque in praesentem diem.
DEUT|4|5|En docui vos praecepta atque iudicia, sicut mandavit mihi Dominus Deus meus, ut faceretis ea in terra, quam possessuri estis,
DEUT|4|6|et observaretis et impleretis opere. Haec est enim vestra sapientia et intellectus coram populis, ut audientes universa praecepta haec dicant: En populus sapiens et intellegens, gens magna haec!".
DEUT|4|7|Quae est enim alia natio tam grandis, quae habeat deos appropinquantes sibi, sicut Dominus Deus noster adest cunctis obsecrationibus nostris?
DEUT|4|8|Et quae est alia gens sic inclita, ut habeat praecepta iustaque iudicia, sicut est universa lex haec, quam ego proponam hodie ante oculos vestros?
DEUT|4|9|Custodi igitur temetipsum et animam tuam sollicite, ne obliviscaris verborum, quae viderunt oculi tui, et ne excidant de corde tuo cunctis diebus vitae tuae. Docebis ea filios ac nepotes tuos
DEUT|4|10|die, in quo stetisti coram Domino Deo tuo in Horeb, quando Dominus locutus est mihi: "Congrega ad me populum, ut audiant sermones meos et discant timere me omni tempore, quo vivunt in terra, doceantque filios suos".
DEUT|4|11|Et accessistis et stetistis ad radices montis, qui ardebat usque ad caelum, erantque in eo tenebrae, nubes et caligo.
DEUT|4|12|Locutusque est Dominus ad vos de medio ignis; vocem verborum audistis et formam penitus non vidistis.
DEUT|4|13|Et ostendit vobis pactum suum, quod praecepit, ut faceretis, et decem verba, quae scripsit in duabus tabulis lapideis.
DEUT|4|14|Mihique mandavit in illo tempore, ut docerem vos praecepta et iudicia, quae facere deberetis in terra, quam possessuri estis.
DEUT|4|15|Custodite igitur sollicite animas vestras. Non vidistis aliquam similitudinem in die, qua locutus est vobis Dominus in Horeb de medio ignis;
DEUT|4|16|ne forte corrupti faciatis vobis sculptam similitudinem, imaginem masculi vel feminae,
DEUT|4|17|similitudinem omnium iumentorum, quae sunt super terram, vel avium sub caelo volantium
DEUT|4|18|atque reptilium, quae moventur in terra, sive piscium, qui sub terra morantur in aquis;
DEUT|4|19|et ne forte oculis elevatis ad caelum videas solem et lunam et astra, omnem exercitum caeli, et errore deceptus adores ea et colas, quae attribuit Dominus Deus tuus cunctis gentibus, quae sub caelo sunt.
DEUT|4|20|Vos autem tulit Dominus et eduxit de fornace ferrea Aegypti, ut haberet populum hereditarium, sicut est in praesenti die.
DEUT|4|21|Iratusque est Dominus contra me propter sermones vestros et iuravit, ut non transirem Iordanem nec ingrederer terram optimam, quam Dominus Deus tuus daturus est tibi in haereditatem.
DEUT|4|22|Ecce morior in hac humo, non transibo Iordanem; vos transibitis et possidebitis terram egregiam hanc.
DEUT|4|23|Cavete, ne quando obliviscamini pacti Domini Dei vestri, quod pepigit vobiscum, et faciatis vobis sculptam similitudinem omnium, quae fieri Dominus Deus tuus prohibuit;
DEUT|4|24|quia Dominus Deus tuus ignis consumens est, Deus aemulator.
DEUT|4|25|Si genueris filios ac nepotes, et morati fueritis in terra corruptique feceritis aliquam similitudinem sculptam patrantes malum coram Domino Deo tuo, ut eum ad iracundiam provocetis,
DEUT|4|26|testes invoco contra vos hodie caelum et terram, cito perituros vos esse de terra, quam, transito Iordane, possessuri estis: non habitabitis in ea longo tempore, sed delebit vos Dominus
DEUT|4|27|atque disperget in gentes, et remanebitis pauci in nationibus, ad quas vos ducturus est Dominus.
DEUT|4|28|Ibique servietis diis, qui hominum manu fabricati sunt, ligno et lapidi, qui non vident nec audiunt nec comedunt nec odorantur.
DEUT|4|29|Cumque quaesieris ibi Dominum Deum tuum, invenies eum, si tamen toto corde quaesieris eum et tota anima tua.
DEUT|4|30|Postquam in tribulatione tua te invenerint omnia, quae praedicta sunt, novissimo tempore reverteris ad Dominum Deum tuum et audies vocem eius;
DEUT|4|31|quia Deus misericors Dominus Deus tuus est, non dimittet te nec omnino delebit neque obliviscetur pacti, in quo iuravit patribus tuis.
DEUT|4|32|Interroga de diebus antiquis, qui fuerunt ante te ex die, quo creavit Deus hominem super terram, et a summo caeli usque ad summum eius, si facta est aliquando huiuscemodi res magna, aut umquam cognitum est,
DEUT|4|33|num audivit populus vocem Dei loquentis de medio ignis, sicut tu audisti et vixisti?
DEUT|4|34|Aut tentavit Deus, ut ingrederetur et tolleret sibi gentem de medio nationis per tentationes, signa atque portenta, per pugnam et robustam manum extentumque brachium et terrores magnos, iuxta omnia, quae fecit pro vobis Dominus Deus vester in Aegypto, videntibus oculis tuis?
DEUT|4|35|Tibi monstratum est, ut scires quoniam Dominus ipse est Deus, et non est alius praeter eum.
DEUT|4|36|De caelo te fecit audire vocem suam, ut doceret te, et in terra ostendit tibi ignem suum maximum; et audisti verba illius de medio ignis,
DEUT|4|37|quia dilexit patres tuos et elegit semen eorum post eos. Eduxitque te vultu suo in virtute sua magna ex Aegypto,
DEUT|4|38|ut expelleret nationes maiores et fortiores te in introitu tuo et introduceret te daretque tibi terram earum in possessionem, sicut cernis in praesenti die.
DEUT|4|39|Scito ergo hodie et cogitato in corde tuo quod Dominus ipse sit Deus in caelo sursum et in terra deorsum, et non sit alius.
DEUT|4|40|Custodi praecepta eius atque mandata, quae ego praecipio tibi hodie, ut bene sit tibi et filiis tuis post te, et permaneas multo tempore super terram, quam Dominus Deus tuus daturus est tibi ".
DEUT|4|41|Tunc separavit Moyses tres civitates trans Iordanem ad orientalem plagam,
DEUT|4|42|ut confugiat ad eas, qui occiderit nolens proximum suum, nec fuerit inimicus ante unum et alterum diem, et ad harum aliquam urbium possit evadere et vivat:
DEUT|4|43|Bosor in solitudine, quae sita est in terra campestri, pro tribu Ruben, et Ramoth in Galaad pro tribu Gad et Golan in Basan pro tribu Manasse.
DEUT|4|44|Ista est lex, quam proposuit Moyses coram filiis Israel;
DEUT|4|45|haec testimonia et praecepta atque iudicia, quae locutus est ad filios Israel, quando egressi sunt de Aegypto,
DEUT|4|46|trans Iordanem in valle contra Bethphegor, in terra Sehon regis Amorraei, qui habitavit in Hesebon, quem percussit Moyses et filii Israel egressi ex Aegypto.
DEUT|4|47|Et possederunt terram eius et terram Og regis Basan, duorum regum Amorraeorum, qui erant trans Iordanem ad solis ortum,
DEUT|4|48|ab Aroer, quae sita est super ripam torrentis Arnon, usque ad montem Sion, qui est Hermon,
DEUT|4|49|omnem Arabam trans Iordanem ad orientalem plagam usque ad mare Arabae et usque ad radices montis Phasga.
DEUT|5|1|Vocavitque Moyses omnem Israelem et dixit ad eos: " Audi, Israel, praecepta atque iudicia, quae ego loquor in auribus vestris hodie; discite ea et opere complete.
DEUT|5|2|Dominus Deus noster pepigit nobiscum foedus in Horeb.
DEUT|5|3|Non cum patribus nostris iniit pactum hoc sed nobiscum, qui in praesentiarum hic sumus, omnibus nobis, qui vivimus.
DEUT|5|4|Facie ad faciem locutus est vobis in monte de medio ignis;
DEUT|5|5|ego sequester et medius fui inter Dominum et vos in tempore illo, ut annuntiarem vobis verba eius; timuistis enim ignem et non ascendistis in montem. Et ait:
DEUT|5|6|"Ego Dominus Deus tuus, qui eduxi te de terra Aegypti, de domo servitutis.
DEUT|5|7|Non habebis deos alienos in conspectu meo.
DEUT|5|8|Non facies tibi sculptile nec similitudinem omnium, quae in caelo sunt desuper et quae in terra deorsum et quae versantur in aquis sub terra.
DEUT|5|9|Non adorabis ea et non coles: Ego enim sum Dominus Deus tuus, Deus aemulator, reddens iniquitatem patrum super filios in tertiam et quartam generationem his, qui oderunt me,
DEUT|5|10|et faciens misericordiam in multa milia diligentibus me et custodientibus praecepta mea.
DEUT|5|11|Non usurpabis nomen Domini Dei tui frustra, quia non erit impunitus, qui super re vana nomen eius assumpserit.
DEUT|5|12|Observa diem sabbati, ut sanctifices eum, sicut praecepit tibi Dominus Deus tuus.
DEUT|5|13|Sex diebus operaberis et facies omnia opera tua.
DEUT|5|14|Septimus dies sabbatum est Domino Deo tuo. Non facies in eo quidquam operis tu et filius tuus et filia, servus et ancilla et bos et asinus et omne iumentum tuum et peregrinus tuus, qui est intra portas tuas, ut requiescat servus tuus et ancilla tua sicut et tu.
DEUT|5|15|Memento quod et ipse servieris in Aegypto, et eduxerit te inde Dominus Deus tuus in manu forti et brachio extento: idcirco praecepit tibi, ut observares diem sabbati.
DEUT|5|16|Honora patrem tuum et matrem, sicut praecepit tibi Dominus Deus tuus, ut longo vivas tempore et bene sit tibi in terra, quam Dominus Deus tuus daturus est tibi.
DEUT|5|17|Non occides.
DEUT|5|18|Neque moechaberis.
DEUT|5|19|Furtumque non facies.
DEUT|5|20|Nec loqueris contra proximum tuum falsum testimonium.
DEUT|5|21|Nec concupisces uxorem proximi tui. Nec desiderabis domum proximi tui, non agrum, non servum, non ancillam, non bovem, non asinum et universa, quae illius sunt".
DEUT|5|22|Haec verba locutus est Dominus ad omnem multitudinem vestram in monte, de medio ignis et nubis et caliginis voce magna nihil addens amplius; et scripsit ea in duabus tabulis lapideis, quas tradidit mihi.
DEUT|5|23|Vos autem, postquam audistis vocem de medio tenebrarum et montem ardere vidistis, accessistis ad me omnes principes tribuum et maiores natu
DEUT|5|24|atque dixistis: "Ecce ostendit nobis Dominus Deus noster maiestatem et magnitudinem suam; vocem eius audivimus de medio ignis et probavimus hodie quod, loquente Deo cum homine, vixerit homo.
DEUT|5|25|Nunc autem cur moriemur, et devorabit nos ignis hic maximus? Si enim audierimus ultra vocem Domini Dei nostri, moriemur.
DEUT|5|26|Quid est omnis caro, ut audiat vocem Dei viventis, qui de medio ignis loquitur, sicut nos audivimus, et possit vivere?
DEUT|5|27|Tu magis accede et audi cuncta, quae dixerit Dominus Deus noster, et tu loqueris ad nos cuncta, quae dixerit Dominus Deus noster tibi, et nos audientes faciemus ea".
DEUT|5|28|Quod cum audisset Dominus, ait ad me: "Audivi vocem verborum populi huius, quae locuti sunt tibi: bene omnia sunt locuti.
DEUT|5|29|Quis det talem eos habere mentem, ut timeant me et custodiant universa mandata mea in omni tempore, ut bene sit eis et filiis eorum in sempiternum?
DEUT|5|30|Vade et dic eis: Revertimini in tentoria vestra.
DEUT|5|31|Tu vero, hic sta mecum, et loquar tibi omnia mandata et praecepta atque iudicia, quae docebis eos, ut faciant ea in terra, quam dabo illis in possessionem".
DEUT|5|32|Custodite igitur et facite, quae praecepit Dominus Deus vester vobis; non declinabitis neque ad dexteram neque ad sinistram,
DEUT|5|33|sed per totam viam, quam praecepit Dominus Deus vester, ambulabitis, ut vivatis, et bene sit vobis, et protelentur dies in terra possessionis vestrae.
DEUT|6|1|Haec sunt mandata et praecep ta atque iudicia, quae mandavit Dominus Deus vester, ut docerem vos, et faciatis ea in terra, ad quam transgredimini possidendam;
DEUT|6|2|ut timeas Dominum Deum tuum et custodias omnia praecepta et mandata eius, quae ego praecipio tibi et filiis ac nepotibus tuis, cunctis diebus vitae tuae, ut prolongentur dies tui.
DEUT|6|3|Audi, Israel, et observa, ut facias, et bene sit tibi, et multipliceris amplius, sicut pollicitus est Dominus, Deus patrum tuorum, tibi terram lacte et melle manantem.
DEUT|6|4|Audi, Israel: Dominus Deus noster Dominus unus est.
DEUT|6|5|Diliges Dominum Deum tuum ex toto corde tuo et ex tota anima tua et ex tota fortitudine tua.
DEUT|6|6|Eruntque verba haec, quae ego praecipio tibi hodie, in corde tuo,
DEUT|6|7|et inculcabis ea filiis tuis et loqueris ea sedens in domo tua et ambulans in itinere, decumbens atque consurgens;
DEUT|6|8|et ligabis ea quasi signum in manu tua, eruntque quasi appensum quid inter oculos tuos,
DEUT|6|9|scribesque ea in postibus domus tuae et in portis tuis.
DEUT|6|10|Cumque introduxerit te Dominus Deus tuus in terram, pro qua iuravit patribus tuis Abraham, Isaac et Iacob, ut daret tibi, civitates magnas et optimas, quas non aedificasti,
DEUT|6|11|domos plenas cunctarum opum, quas non implevisti, cisternas, quas non fodisti, vineta et oliveta, quae non plantasti, et comederis et saturatus fueris,
DEUT|6|12|cave diligenter, ne obliviscaris Domini, qui eduxit te de terra Aegypti, de domo servitutis:
DEUT|6|13|Dominum Deum tuum timebis et ipsi servies ac per nomen illius iurabis.
DEUT|6|14|Non ibitis post deos alienos, de diis gentium, quae in circuitu vestro sunt,
DEUT|6|15|quoniam Deus aemulator Dominus Deus tuus in medio tui; ne quando irascatur furor Domini Dei tui contra te et auferat te de superficie terrae.
DEUT|6|16|Non tentabitis Dominum Deum vestrum, sicut tentastis in Massa.
DEUT|6|17|Custodite mandata Domini Dei vestri ac testimonia et praecepta, quae praecepit tibi;
DEUT|6|18|et fac, quod rectum est et bonum in conspectu Domini, ut bene sit tibi, et ingressus possideas terram optimam, de qua iuravit Dominus patribus tuis,
DEUT|6|19|ut deleret omnes inimicos tuos coram te, sicut locutus est Dominus.
DEUT|6|20|Cumque interrogaverit te filius tuus cras dicens: "Quid sibi volunt testimonia haec et praecepta atque iudicia, quae praecepit Dominus Deus noster vobis?",
DEUT|6|21|dices ei: "Servi eramus pharaonis in Aegypto, et eduxit nos Dominus de Aegypto in manu forti
DEUT|6|22|fecitque signa atque prodigia magna et pessima in Aegypto contra pharaonem et omnem domum illius in conspectu nostro;
DEUT|6|23|et eduxit nos inde, ut introductis daret terram, super qua iuravit patribus nostris.
DEUT|6|24|Praecepitque nobis Dominus, ut faciamus omnia praecepta haec et timeamus Dominum Deum nostrum, et bene sit nobis cunctis diebus vitae nostrae, sicut est hodie.
DEUT|6|25|Eritque iustitia nobis, si custodierimus et fecerimus omnia mandata haec coram Domino Deo nostro, sicut mandavit nobis".
DEUT|7|1|Cum introduxerit te Dominus Deus tuus in terram, quam pos sessurus ingredieris, et deleverit gentes multas coram te, Hetthaeum et Gergesaeum et Amorraeum, Chananaeum et Pherezaeum et Hevaeum et Iebusaeum, septem gentes multo maioris numeri quam tu es et robustiores te,
DEUT|7|2|tradideritque eas Dominus Deus tuus tibi, percuties eas usque ad internecionem. Non inibis cum eis foedus nec misereberis earum
DEUT|7|3|neque sociabis cum eis coniugia; filiam tuam non dabis filio eius nec filiam illius accipies filio tuo,
DEUT|7|4|quia seducet filium tuum, ne sequatur me et ut serviat diis alienis, irasceturque furor Domini contra vos et delebit te cito.
DEUT|7|5|Quin potius haec facietis eis: aras eorum subvertite et confringite lapides et palos lucosque succidite et sculptilia comburite;
DEUT|7|6|quia populus sanctus es Domino Deo tuo. Te elegit Dominus Deus tuus, ut sis ei populus peculiaris de cunctis populis, qui sunt super terram.
DEUT|7|7|Non quia cunctas gentes numero vincebatis, vobis iunctus est Dominus et elegit vos, cum omnibus sitis populis pauciores,
DEUT|7|8|sed quia dilexit vos Dominus et custodivit iuramentum, quod iuravit patribus vestris, eduxit vos in manu forti et redemit te de domo servitutis, de manu pharaonis regis Aegypti.
DEUT|7|9|Et scies quia Dominus Deus tuus ipse est Deus, Deus fidelis, custodiens pactum et misericordiam diligentibus se et his, qui custodiunt mandata eius, in mille generationes
DEUT|7|10|et reddens odientibus se protinus, ita ut disperdat eos et ultra non differat, protinus eis restituens, quod merentur.
DEUT|7|11|Custodi ergo mandata et praecepta atque iudicia, quae ego mando tibi hodie, ut facias.
DEUT|7|12|Si audieritis haec iudicia et custodieritis ea et feceritis, custodiet et Dominus Deus tuus tibi pactum et misericordiam, quam iuravit patribus tuis,
DEUT|7|13|et diliget te et benedicet tibi ac multiplicabit te benedicetque fructui ventris tui et fructui terrae tuae, frumento tuo atque vindemiae, oleo et partui armentorum et incremento ovium tuarum super terram, pro qua iuravit patribus tuis, ut daret eam tibi.
DEUT|7|14|Benedictus eris prae omnibus populis. Non erit apud te sterilis utriusque sexus, tam in hominibus quam in gregibus tuis.
DEUT|7|15|Auferet Dominus a te omnem languorem; et infirmitates Aegypti pessimas, quas novisti, non inferet tibi, sed cunctis hostibus tuis.
DEUT|7|16|Devorabis omnes populos, quos Dominus Deus tuus daturus est tibi; non parcet eis oculus tuus, nec servies diis eorum, ne sint in ruinam tui.
DEUT|7|17|Si dixeris in corde tuo: "Plures sunt gentes istae quam ego; quomodo potero delere eas?",
DEUT|7|18|noli metuere eas, sed recordare, quae fecerit Dominus Deus tuus pharaoni et cunctis Aegyptiis,
DEUT|7|19|plagas maximas, quas viderunt oculi tui, et signa atque portenta manumque robustam et extentum brachium, ut educeret te Dominus Deus tuus; sic faciet cunctis populis, quos metuis.
DEUT|7|20|Insuper et crabrones mittet Dominus Deus tuus in eos, donec deleat omnes atque disperdat, qui te fugerint et latere potuerint.
DEUT|7|21|Non timebis eos, quia Dominus Deus tuus in medio tui est, Deus magnus et terribilis.
DEUT|7|22|Ipse consumet nationes has in conspectu tuo paulatim atque per partes. Non poteris delere eas cito, ne multiplicentur contra te bestiae terrae.
DEUT|7|23|Dabitque eos Dominus Deus tuus in conspectu tuo et conturbabit illos conturbatione magna, donec penitus deleantur.
DEUT|7|24|Tradetque reges eorum in manus tuas, et disperdes nomina eorum sub caelo; nullus poterit resistere tibi, donec conteras eos.
DEUT|7|25|Sculptilia eorum igne combures; non concupisces argentum et aurum, quibus vestita sunt, neque assumes ex eis tibi quidquam, ne offendas propterea, quia abominatio est Domini Dei tui.
DEUT|7|26|Nec inferes abominationem in domum tuam, ne fias anathema sicut et illa est; quasi spurcitiam detestaberis et velut inquinamentum ac sordes abominationi habebis, quia anathema est.
DEUT|8|1|Omne mandatum, quod ego praecipio tibi hodie, cave dili genter ut facias, ut possitis vivere et multiplicemini ingressique possideatis terram, pro qua iuravit Dominus patribus vestris.
DEUT|8|2|Et recordaberis cuncti itineris, per quod adduxit te Dominus Deus tuus his quadraginta annis per desertum, ut affligeret te atque tentaret, et nota fierent, quae in tuo animo versabantur, utrum custodires mandata illius an non.
DEUT|8|3|Afflixit te penuria et dedit tibi cibum manna, quem ignorabas tu et patres tui, ut ostenderet tibi quod non in solo pane vivat homo, sed in omni verbo, quod egreditur de ore Domini.
DEUT|8|4|Vestimentum tuum, quo operiebaris, nequaquam defecit, et pes tuus non intumuit his quadraginta annis.
DEUT|8|5|Recogites ergo in corde tuo quia, sicut erudit homo filium suum, sic Dominus Deus tuus erudivit te,
DEUT|8|6|ut custodias mandata Domini Dei tui et ambules in viis eius et timeas eum.
DEUT|8|7|Dominus enim Deus tuus introducet te in terram bonam, terram rivorum aquarum et fontium, in cuius campis et montibus erumpunt fluviorum abyssi,
DEUT|8|8|terram frumenti, hordei ac vinearum, in qua ficus et malogranata et oliveta nascuntur, terram olei ac mellis,
DEUT|8|9|ubi absque ulla penuria comedes panem tuum et rerum omnium abundantia perfrueris; cuius lapides ferrum sunt, et de montibus eius aeris metalla fodiuntur;
DEUT|8|10|ut, cum comederis et satiatus fueris, benedicas Domino Deo tuo pro terra optima, quam dedit tibi.
DEUT|8|11|Observa et cave, ne quando obliviscaris Domini Dei tui et neglegas mandata eius atque iudicia et praecepta, quae ego praecipio tibi hodie;
DEUT|8|12|ne, postquam comederis et satiatus fueris, domos pulchras aedificaveris et habitaveris in eis
DEUT|8|13|habuerisque armenta et ovium greges multos, argenti et auri cunctarumque rerum copiam,
DEUT|8|14|elevetur cor tuum, et obliviscaris Domini Dei tui, qui eduxit te de terra Aegypti, de domo servitutis,
DEUT|8|15|et ductor tuus fuit in solitudine magna atque terribili, in qua erat serpens adurens et scorpio ac terra arida et nullae omnino aquae; qui eduxit tibi rivos de petra durissima
DEUT|8|16|et cibavit te manna in solitudine, quod nescierunt patres tui, et, postquam afflixit ac probavit te, ad extremum misertus est tui,
DEUT|8|17|ne diceres in corde tuo: "Fortitudo mea et robur manus meae haec mihi omnia praestiterunt";
DEUT|8|18|sed recorderis Domini Dei tui, quod ipse vires tibi praebuerit, ut consequereris prosperitatem, ut impleret pactum suum, super quo iuravit patribus tuis, sicut praesens indicat dies.
DEUT|8|19|Sin autem oblitus Domini Dei tui secutus fueris deos alienos coluerisque illos et adoraveris, ecce nunc testificor vobis quod omnino dispereatis:
DEUT|8|20|sicut gentes, quas delevit Dominus in introitu vestro, ita et vos peribitis, si inoboedientes fueritis voci Domini Dei vestri.
DEUT|9|1|Audi, Israel: Tu transgredieris hodie Iordanem, ut possideas nationes maximas et fortiores te, civitates ingentes et ad caelum usque muratas,
DEUT|9|2|populum magnum atque sublimem, filios Enacim, quos ipse nosti et audisti, quibus nullus potest ex adverso resistere.
DEUT|9|3|Scies ergo hodie quod Dominus Deus tuus ipse transibit ante te ignis devorans, qui conteret eos atque subiciet ante faciem tuam, ut velociter expellas et deleas eos, sicut locutus est tibi.
DEUT|9|4|Ne dicas in corde tuo, cum deleverit eos Dominus Deus tuus in conspectu tuo: "Propter iustitiam meam introduxit me Dominus, ut terram hanc possiderem", cum propter impietates nationum istarum expellat eas Dominus ante te.
DEUT|9|5|Neque enim propter iustitiam tuam et aequitatem cordis tui ingredieris, ut possideas terras earum, sed quia illae egerunt impie, introeunte te, Dominus Deus tuus expellet eos ante te, et ut compleat verbum suum Dominus, quod sub iuramento pollicitus est patribus tuis, Abraham, Isaac et Iacob.
DEUT|9|6|Scito igitur quod non propter iustitiam tuam Dominus Deus tuus dederit tibi terram hanc optimam in possessionem, cum durissimae cervicis sis populus.
DEUT|9|7|Memento et ne obliviscaris quomodo ad iracundiam provocaveris Dominum Deum tuum in solitudine; ex eo die, quo egressus es ex Aegypto, usque ad locum istum adversum Dominum contendistis.
DEUT|9|8|Nam et in Horeb provocastis eum, et iratus delere vos voluit,
DEUT|9|9|quando ascendi in montem, ut acciperem tabulas lapideas, tabulas pacti, quod pepigit vobiscum Dominus, et perseveravi in monte quadraginta diebus ac noctibus panem non comedens et aquam non bibens.
DEUT|9|10|Deditque mihi Dominus duas tabulas lapideas scriptas digito Dei et continentes omnia verba, quae vobis locutus est in monte de medio ignis, quando contio populi congregata est.
DEUT|9|11|Cumque transissent quadraginta dies et totidem noctes, dedit mihi Dominus duas tabulas lapideas, tabulas foederis,
DEUT|9|12|dixitque mihi: "Surge et descende hinc cito, quia peccavit populus tuus, quem eduxisti de Aegypto: deseruerunt velociter viam, quam praecepi eis, feceruntque sibi conflatile".
DEUT|9|13|Rursumque ait Dominus ad me: "Cerno quod populus iste durae cervicis sit;
DEUT|9|14|dimitte me, ut conteram eos et deleam nomen eorum sub caelo et faciam te in gentem, quae hac fortior et maior sit".
DEUT|9|15|Cumque reversus de monte ardente descenderem et duas tabulas foederis utraque tenerem manu
DEUT|9|16|vidissemque vos peccasse Domino Deo vestro et fecisse vobis vitulum conflatilem ac deseruisse velociter viam eius, quam Dominus vobis praeceperat,
DEUT|9|17|arripui duas tabulas et proieci eas de manibus meis confregique eas in conspectu vestro;
DEUT|9|18|et procidi ante Dominum, sicut prius quadraginta diebus et noctibus panem non comedens et aquam non bibens propter omnia peccata vestra, quae gessistis contra Dominum et eum ad iracundiam provocastis;
DEUT|9|19|timui enim indignationem et iram illius, qua adversum vos concitatus delere vos voluit. Et exaudivit me Dominus etiam hac vice.
DEUT|9|20|Adversum Aaron quoque vehementer iratus voluit eum conterere; et pro illo similiter tunc deprecatus sum.
DEUT|9|21|Peccatum autem vestrum, quod feceratis, id est vitulum, arripiens igne combussi et in frusta comminuens omninoque in pulverem redigens proieci in torrentem, qui de monte descendit.
DEUT|9|22|In Tabera quoque et in Massa et in Cibrottaava provocastis Dominum;
DEUT|9|23|et quando misit Dominus vos de Cadesbarne dicens: "Ascendite et possidete terram, quam dedi vobis", contempsistis imperium Domini Dei vestri et non credidistis ei neque vocem eius audire voluistis;
DEUT|9|24|semper fuistis rebelles contra Dominum a die, qua nosse vos coepi.
DEUT|9|25|Et iacui coram Domino quadraginta diebus ac noctibus, quibus eum suppliciter deprecabar, ne deleret vos, ut fuerat comminatus.
DEUT|9|26|Et orans dixi: Domine Deus, ne disperdas populum tuum et hereditatem tuam, quam redemisti in magnitudine tua, quos eduxisti de Aegypto in manu forti.
DEUT|9|27|Recordare servorum tuorum Abraham, Isaac et Iacob; ne aspicias duritiam populi huius et impietatem atque peccatum,
DEUT|9|28|ne forte dicant habitatores terrae, de qua eduxisti nos: "Non poterat Dominus introducere eos in terram, quam pollicitus est eis, et oderat illos; idcirco eduxit, ut interficeret eos in solitudine".
DEUT|9|29|Attamen ipsi sunt populus tuus et hereditas tua, quos eduxisti in fortitudine tua magna et in brachio tuo extento.
DEUT|10|1|In tempore illo dixit Dominus ad me: "Dola tibi duas tabulas lapideas, sicut priores fuerunt, et ascende ad me in montem faciesque tibi arcam ligneam.
DEUT|10|2|Et scribam in tabulis verba, quae fuerunt in his, quas ante confregisti, ponesque eas in arca".
DEUT|10|3|Feci igitur arcam de lignis acaciae; cumque dolassem duas tabulas lapideas instar priorum, ascendi in montem habens eas in manibus.
DEUT|10|4|Scripsitque in tabulis iuxta id quod prius scripserat, verba decem, quae locutus est Dominus ad vos in monte de medio ignis, quando populus congregatus est, et dedit eas mihi.
DEUT|10|5|Reversusque de monte descendi et posui tabulas in arcam, quam feceram; quae hucusque ibi sunt, sicut mihi praecepit Dominus.
DEUT|10|6|Filii autem Israel castra moverunt ex Berothbeneiacan in Mosera, ubi Aaron mortuus ac sepultus est; pro quo sacerdotio functus est Eleazar filius eius.
DEUT|10|7|Inde venerunt in Gadgad; de quo loco profecti castrametati sunt in Ietebatha, in terra torrentium aquarum.
DEUT|10|8|Eo tempore separavit Dominus tribum Levi, ut portaret arcam foederis Domini et staret coram eo in ministerio ac benediceret in nomine illius usque in praesentem diem.
DEUT|10|9|Quam ob rem non habuit Levi partem neque hereditatem cum fratribus suis, quia ipse Dominus hereditas eius est, sicut promisit ei Dominus Deus tuus.
DEUT|10|10|Ego autem steti in monte sicut prius quadraginta diebus ac noctibus, exaudivitque me Dominus etiam hac vice et te perdere noluit.
DEUT|10|11|Dixitque mihi: "Surge, vade et praecede populum, ut ingrediatur et possideat terram, quam iuravi patribus eorum, ut traderem eis".
DEUT|10|12|Et nunc, Israel, quid Dominus Deus tuus petit a te, nisi ut timeas Dominum Deum tuum et ambules in viis eius et diligas eum ac servias Domino Deo tuo in toto corde tuo et in tota anima tua
DEUT|10|13|custodiasque mandata Domini et praecepta eius, quae ego hodie praecipio, ut bene sit tibi?
DEUT|10|14|En Domini Dei tui caelum est et caelum caeli, terra et omnia, quae in ea sunt;
DEUT|10|15|et tamen patribus tuis conglutinatus est Dominus et amavit eos elegitque semen eorum post eos, id est vos, de cunctis gentibus, sicut hodie comprobatur.
DEUT|10|16|Circumcidite igitur praeputium cordis vestri et cervicem vestram, ne induretis amplius,
DEUT|10|17|quia Dominus Deus vester ipse est Deus deorum et Dominus dominantium, Deus magnus, potens et terribilis, qui personam non accipit nec munera,
DEUT|10|18|facit iudicium pupillo et viduae, amat peregrinum et dat ei victum atque vestitum.
DEUT|10|19|Et vos ergo, amate peregrinos, quia et ipsi fuistis advenae in terra Aegypti.
DEUT|10|20|Dominum Deum tuum timebis et ei servies, ipsi adhaerebis iurabisque in nomine illius.
DEUT|10|21|Ipse est laus tua et Deus tuus, qui fecit tibi haec magnalia et terribilia, quae viderunt oculi tui.
DEUT|10|22|In septuaginta animabus descenderunt patres tui in Aegyptum; et ecce nunc multiplicavit te Dominus Deus tuus sicut astra caeli.
DEUT|11|1|Ama itaque Dominum Deum tuum et custodi obser vationem eius et praecepta, iudicia atque mandata omni tempore.
DEUT|11|2|Cognoscite hodie, quae ignorant filii vestri, qui non viderunt disciplinam Domini Dei vestri, magnalia eius et robustam manum extentumque brachium,
DEUT|11|3|signa et opera, quae fecit in medio Aegypti pharaoni regi et universae terrae eius
DEUT|11|4|omnique exercitui Aegyptiorum et equis ac curribus; quomodo operuerint eos aquae maris Rubri, cum vos persequerentur, et deleverit eos Dominus usque in praesentem diem;
DEUT|11|5|vobisque, quae fecerit in solitudine, donec veniretis ad hunc locum;
DEUT|11|6|et Dathan atque Abiram filiis Eliab, qui fuit filius Ruben, quos aperto ore suo terra absorbuit cum domibus et tabernaculis et universa substantia eorum, quam habebant in medio Israel.
DEUT|11|7|Oculi vestri viderunt omnia opera Domini magna, quae fecit,
DEUT|11|8|ut custodiatis universa mandata, quae ego hodie praecipio vobis, ut roboremini et possitis introire et possidere terram, ad quam ingredimini,
DEUT|11|9|multoque in ea vivatis tempore, quam sub iuramento pollicitus est Dominus patribus vestris et semini eorum, lacte et melle manantem.
DEUT|11|10|Terra enim, ad quam ingredieris possidendam, non est sicut terra Aegypti, de qua existis, ubi, iacto semine, in hortorum morem aquae pede ducuntur irriguae;
DEUT|11|11|sed montuosa est et campestris, de caelo exspectans pluvias,
DEUT|11|12|quam Dominus Deus tuus semper invisit, et oculi illius in ea sunt a principio anni usque ad finem eius.
DEUT|11|13|Si ergo oboedieritis mandatis meis, quae hodie praecipio vobis, ut diligatis Dominum Deum vestrum et serviatis ei in toto corde vestro et in tota anima vestra,
DEUT|11|14|dabo pluviam terrae vestrae temporaneam et serotinam in tempore suo, ut colligas frumentum et vinum et oleum,
DEUT|11|15|et dabit fenum ex agris ad pascenda iumenta, et ut ipse comedas ac satureris.
DEUT|11|16|Cavete, ne decipiatur cor vestrum, et recedatis a Domino serviatisque diis alienis et adoretis eos,
DEUT|11|17|iratusque Dominus contra vos claudat caelum, et pluviae non descendant, nec terra det fructum suum, pereatisque velociter de terra optima, quam Dominus daturus est vobis.
DEUT|11|18|Ponite haec verba mea in cordibus et in animis vestris et ligate ea pro signo in manibus et inter oculos vestros collocate quasi appensum quid.
DEUT|11|19|Docete ea filios vestros, de illis loquendo, quando sederis in domo tua et ambulaveris in via et accubueris atque surrexeris.
DEUT|11|20|Scribes ea super postes domus tuae et portas tuas,
DEUT|11|21|ut multiplicentur dies tui et filiorum tuorum in terra, quam iuravit Dominus patribus tuis, ut daret eis, quamdiu caelum imminet terrae.
DEUT|11|22|Si enim custodieritis omnia mandata haec, quae ego praecipio vobis, et feceritis ea, ut diligatis Dominum Deum vestrum et ambuletis in omnibus viis eius adhaerentes ei,
DEUT|11|23|disperdet Dominus omnes gentes istas ante faciem vestram, et possidebitis eas, quae maiores et fortiores vobis sunt;
DEUT|11|24|omnis locus, quem calcaverit pes vester, vester erit. A deserto et a Libano, a flumine magno Euphrate usque ad mare occidentale erunt termini vestri.
DEUT|11|25|Nullus stabit contra vos; terrorem vestrum et formidinem dabit Dominus Deus vester super omnem terram, quam calcaturi estis, sicut locutus est vobis.
DEUT|11|26|En propono in conspectu vestro hodie benedictionem et maledictionem:
DEUT|11|27|benedictionem, si oboedieritis mandatis Domini Dei vestri, quae ego hodie praecipio vobis;
DEUT|11|28|maledictionem, si non oboedieritis mandatis Domini Dei vestri, sed recesseritis de via, quam ego nunc ostendo vobis, et ambulaveritis post deos alienos, quos ignoratis.
DEUT|11|29|Cum introduxerit te Dominus Deus tuus in terram, ad quam pergis habitandam, pones benedictionem super montem Garizim, maledictionem super montem Hebal,
DEUT|11|30|qui sunt trans Iordanem, post viam quae vergit ad solis occubitum in terra Chananaei, qui habitat in Araba contra Galgalam, quae est iuxta Quercus Moreh.
DEUT|11|31|Vos enim transibitis Iordanem, ut possideatis terram, quam Dominus Deus vester daturus est vobis, et habitetis in illa.
DEUT|11|32|Videte ergo ut impleatis omnia praecepta atque iudicia, quae ego hodie ponam in conspectu vestro.
DEUT|12|1|Haec sunt praecepta atque iudicia, quae facere debetis in terra, quam Dominus, Deus patrum tuorum, daturus est tibi, ut possideas eam cunctis diebus, quibus super humum gradieris.
DEUT|12|2|Subvertite omnia loca, in quibus coluerunt gentes, quas possessuri estis, deos suos super montes excelsos et colles et subter omne lignum frondosum.
DEUT|12|3|Dissipate aras eorum et confringite lapides, palos igne comburite et idola comminuite, disperdite nomina eorum de locis illis.
DEUT|12|4|Non facietis ita Domino Deo vestro.
DEUT|12|5|Sed ad locum, quem elegerit Dominus Deus vester de cunctis tribubus vestris, ut ponat nomen suum ibi et habitet in eo, venietis
DEUT|12|6|et offeretis in illo loco holocausta et victimas vestras, decimas et donaria manuum vestrarum et vota atque dona, primogenita boum et ovium.
DEUT|12|7|Et comedetis ibi in conspectu Domini Dei vestri ac laetabimini in cunctis, ad quae miseritis manum vos et domus vestrae, in quibus benedixerit vobis Dominus Deus vester.
DEUT|12|8|Non facietis secundum omnia, quae nos hic facimus hodie, singuli, quod sibi rectum videtur;
DEUT|12|9|neque enim usque in praesens tempus venistis ad requiem et possessionem, quam Dominus Deus vester daturus est vobis.
DEUT|12|10|Transibitis Iordanem et habitabitis in terra, quam Dominus Deus vester daturus est vobis, ut requiescatis a cunctis hostibus per circuitum et absque ullo timore habitetis
DEUT|12|11|in loco, quem elegerit Dominus Deus vester, ut habitet nomen eius in eo. Illuc omnia, quae praecipio, conferetis: holocausta et hostias ac decimas et donaria manuum vestrarum et, quidquid praecipuum est in muneribus, quae vovebitis Domino.
DEUT|12|12|Ibi laetabimini coram Domino Deo vestro vos, filii ac filiae vestrae, famuli et famulae atque Levites, qui in urbibus vestris commoratur; neque enim habet partem et possessionem inter vos.
DEUT|12|13|Cave, ne offeras holocausta tua in omni loco, quem videris,
DEUT|12|14|sed in eo, quem elegerit Dominus in una tribuum tuarum, offeres holocausta et ibi facies quaecumque praecipio tibi.
DEUT|12|15|Sin autem comedere volueris, et te esus carnium delectaverit, occide et comede carnem iuxta benedictionem Domini Dei tui, quam dedit tibi in omnibus urbibus tuis; sive immundus sive mundus comedet illam, sicut capream et cervum,
DEUT|12|16|absque esu dumtaxat sanguinis, quem super terram quasi aquam effundes.
DEUT|12|17|Non poteris comedere in oppidis tuis decimam frumenti et vini et olei tui, primogenita armentorum et pecorum et omnia, quae voveris et sponte offerre volueris, et primitiva manuum tuarum.
DEUT|12|18|Sed coram Domino Deo tuo comedes ea in loco, quem elegerit Dominus Deus tuus, tu et filius tuus ac filia tua, servus et famula atque Levites, qui manet in urbibus tuis; et laetaberis coram Domino Deo tuo in cunctis, ad quae extenderis manum tuam.
DEUT|12|19|Cave, ne derelinquas Levitem omni tempore, quo versaris in terra tua.
DEUT|12|20|Quando dilataverit Dominus Deus tuus terminos tuos, sicut locutus est tibi, et volueris vesci carnibus, quas desiderat anima tua, comedes carnem secundum omne desiderium animae tuae;
DEUT|12|21|locus autem, quem elegerit Dominus Deus tuus, ut sit nomen eius ibi, si procul fuerit, occides de armentis et pecoribus, quae dederit tibi Dominus, sicut praecepi tibi, et comedes in oppidis tuis, ut tibi placet.
DEUT|12|22|Sicut comeditur caprea et cervus, ita vesceris eis; et mundus et immundus in commune vescentur.
DEUT|12|23|Hoc solum cave, ne sanguinem comedas; sanguis enim eorum anima est, et idcirco non debes animam comedere cum carnibus.
DEUT|12|24|Non comedes eum, sed super terram fundes quasi aquam;
DEUT|12|25|non comedes eum, ut bene sit tibi et filiis tuis post te, cum feceris, quod placet in conspectu Domini.
DEUT|12|26|Quae autem sanctificaveris et voveris Domino, tolles et venies ad locum, quem elegerit Dominus,
DEUT|12|27|et offeres holocausta tua, carnem et sanguinem super altare Domini Dei tui; sanguis hostiarum tuarum fundetur in altari, carnibus autem ipse vesceris.
DEUT|12|28|Observa et audi omnia, quae ego praecipio tibi, ut bene sit tibi et filiis tuis post te in sempiternum, cum feceris, quod bonum est et placitum in conspectu Domini Dei tui.
DEUT|12|29|Quando disperdiderit Dominus Deus tuus ante faciem tuam gentes, ad quas ingredieris possidendas, et possederis eas atque habitaveris in terra earum,
DEUT|12|30|cave, ne irretiaris per eas, postquam te fuerint introeunte subversae, et requiras caeremonias earum dicens: "Sicut coluerunt gentes istae deos suos, ita et ego colam".
DEUT|12|31|Non facies similiter Domino Deo tuo; omnes enim abominationes, quas aversatur Dominus, fecerunt diis suis offerentes etiam filios et filias et comburentes igne.
DEUT|13|1|Quod praecipio vobis, hoc custodite et facite, nec addas quidquam nec minuas.
DEUT|13|2|Si surrexerit in medio tui prophetes aut, qui somnium vidisse se dicat, et dederit tibi signum vel portentum,
DEUT|13|3|et evenerit, quod locutus est, et dixerit tibi: "Eamus et sequamur deos alienos, quos ignoras, et serviamus eis",
DEUT|13|4|non audies verba prophetae illius aut somniatoris, quia tentat vos Dominus Deus vester, ut sciat utrum diligatis eum an non in toto corde et in tota anima vestra.
DEUT|13|5|Dominum Deum vestrum sequimini et ipsum timete et mandata illius custodite et audite vocem eius; ipsi servietis et ipsi adhaerebitis.
DEUT|13|6|Propheta autem ille aut fictor somniorum interficietur, quia locutus est, ut vos averteret a Domino Deo vestro, qui eduxit vos de terra Aegypti et redemit te de domo servitutis; ut errare te faceret de via, quam tibi praecepit Dominus Deus tuus; et auferes malum de medio tui.
DEUT|13|7|Si tibi voluerit persuadere frater tuus filius matris tuae aut filius tuus vel filia sive uxor, quae est in sinu tuo, aut amicus, quem diligis ut animam tuam, clam dicens: "Eamus et serviamus diis alienis", quos ignorasti tu et patres tui,
DEUT|13|8|de diis cunctarum in circuitu gentium, quae iuxta vel procul sunt ab initio usque ad finem terrae,
DEUT|13|9|non acquiescas ei nec audias, neque parcat ei oculus tuus, ut miserearis et occultes eum,
DEUT|13|10|sed interficies. Sit primum manus tua super eum, et postea omnis populus mittat manum:
DEUT|13|11|lapidibus obrutus necabitur, quia voluit te abstrahere a Domino Deo tuo, qui eduxit te de terra Aegypti, de domo servitutis,
DEUT|13|12|ut omnis Israel audiens timeat, et nequaquam ultra faciat quippiam huius rei simile in medio tui.
DEUT|13|13|Si audieris in una urbium tuarum, quas Dominus Deus tuus dabit tibi ad habitandum, dicentes aliquos:
DEUT|13|14|"Egressi sunt filii Belial de medio tui et averterunt habitatores urbis suae atque dixerunt: Eamus et serviamus diis alienis", quos ignorastis,
DEUT|13|15|quaere sollicite et, diligenter rei veritate perspecta, si inveneris certum esse, quod dicitur, et abominationem hanc opere perpetratam in medio tui,
DEUT|13|16|percuties habitatores urbis illius in ore gladii et delebis eam ac omnia, quae in illa sunt.
DEUT|13|17|Quidquid etiam supellectilis fuerit, congregabis in medio platearum eius et cum ipsa civitate succendes, ita ut universa consumas Domino Deo tuo, et sit tumulus sempiternus: non aedificabitur amplius.
DEUT|13|18|Et non adhaerebit de illo anathemate quidquam in manu tua, ut avertatur Dominus ab ira furoris sui et misereatur tui multiplicetque te, sicut iuravit patribus tuis,
DEUT|13|19|quando audieris vocem Domini Dei tui custodiens omnia mandata eius, quae ego praecipio tibi hodie, ut facias quod placitum est in conspectu Domini Dei tui.
DEUT|14|1|Filii estote Domini Dei ve stri; non vos incidetis nec fa cietis calvitium inter oculos vestros super mortuo,
DEUT|14|2|quoniam populus sanctus es Domino Deo tuo, et te elegit, ut sis ei in populum peculiarem de cunctis gentibus, quae sunt super terram.
DEUT|14|3|Ne comedatis quidquid abominabile est.
DEUT|14|4|Hoc est animal, quod comedere potestis: bovem et ovem et capram,
DEUT|14|5|cervum et capream, bubalum, tragelaphum, pygargum, orygem, rupicapram.
DEUT|14|6|Omne animal inter pecora, quod findit ungulam plene in duas partes et ruminat, comedetis;
DEUT|14|7|de his autem, quae ruminant et ungulam non findunt, haec comedere non debetis: camelum, leporem, hyracem, quia ruminant et non dividunt ungulam, immunda erunt vobis.
DEUT|14|8|Sus quoque, quoniam dividit ungulam et non ruminat, immunda erit vobis: carnibus eorum non vescemini et cadavera non tangetis.
DEUT|14|9|Haec comedetis ex omnibus, quae morantur in aquis: quae habent pinnulas et squamas comedite;
DEUT|14|10|quae absque pinnulis et squamis sunt, ne comedatis, quia immunda sunt vobis.
DEUT|14|11|Omnes aves mundas comedite;
DEUT|14|12|has autem ne comedatis: aquilam scilicet et grypem et alietum,
DEUT|14|13|ixon et vulturem ac milvum iuxta genus suum
DEUT|14|14|et omne corvini generis,
DEUT|14|15|struthionem ac noctuam et larum atque accipitrem iuxta genus suum,
DEUT|14|16|bubonem ac cycnum et ibin
DEUT|14|17|ac mergulum, porphyrionem et nycticoracem,
DEUT|14|18|erodium et charadrium, singula in genere suo, upupam quoque et vespertilionem.
DEUT|14|19|Et omne, quod reptat et pinnulas habet, immundum erit vobis, nec comedetur.
DEUT|14|20|Omne volatile, quod mundum est, comedite.
DEUT|14|21|Quidquid morticinum est, ne vescamini ex eo; advenae, qui intra portas tuas est, da, ut comedat, aut vende peregrino: quia tu populus sanctus es Domino Deo tuo.Non coques haedum in lacte matris suae.
DEUT|14|22|Decimam partem separabis de cunctis frugibus seminis tui, quae nascuntur in terra per annos singulos;
DEUT|14|23|et comedes in conspectu Domini Dei tui in loco, quem elegerit, ut in eo nomen illius habitet, decimam frumenti tui et vini et olei et primogenita de armentis et ovibus tuis, ut discas timere Dominum Deum tuum omni tempore.
DEUT|14|24|Cum autem longior fuerit tibi via et locus, quem elegerit Dominus Deus tuus, ut ponat nomen suum ibi tibique benedixerit, nec potueris ad eum haec cuncta portare,
DEUT|14|25|vendes omnia et in pretium rediges; portabisque manu tua et proficisceris ad locum, quem elegerit Dominus Deus tuus,
DEUT|14|26|et emes ex eadem pecunia, quidquid tibi placuerit, sive ex armentis sive ex ovibus, vinum quoque et siceram et omne, quod desiderat anima tua; et comedes ibi coram Domino Deo tuo et epulaberis tu et domus tua
DEUT|14|27|et Levites, qui intra portas tuas est: cave, ne derelinquas eum, quia non habet partem nec possessionem tecum.
DEUT|14|28|Anno tertio separabis aliam decimam ex omnibus, quae nascuntur tibi eo tempore, et repones intra portas tuas;
DEUT|14|29|venietque Levites, qui non habet partem nec possessionem tecum, et peregrinus ac pupillus ac vidua, qui intra portas tuas sunt, et comedent et saturabuntur, ut benedicat tibi Dominus Deus tuus in cunctis operibus manuum tuarum, quae feceris.
DEUT|15|1|Septimo anno facies remis sionem,
DEUT|15|2|quae hoc ordine ce lebrabitur: cui debetur aliquid a proximo ac fratre suo, repetere non poterit, quia annus remissionis est Domino.
DEUT|15|3|A peregrino exiges; civem et propinquum repetendi, quod tuum est, non habebis potestatem.
DEUT|15|4|Sed omnino indigens non erit apud te, quia benedicet tibi Dominus Deus tuus in terra, quam traditurus est tibi in possessionem,
DEUT|15|5|si tamen audieris vocem Domini Dei tui et custodieris universum mandatum hoc, quod ego hodie praecipio tibi,
DEUT|15|6|quia Dominus Deus tuus benedicet tibi, ut pollicitus est. Fenerabis gentibus multis et ipse a nullo accipies mutuum; dominaberis nationibus plurimis, et tui nemo dominabitur.
DEUT|15|7|Si unus de fratribus tuis, qui morantur in una civitatum tuarum in terra, quam Dominus Deus tuus daturus est tibi, ad paupertatem venerit, non obdurabis cor tuum nec contrahes manum;
DEUT|15|8|sed aperies eam pauperi fratri tuo et dabis mutuum, quod eum indigere perspexeris.
DEUT|15|9|Cave, ne forte subrepat tibi impia cogitatio, et dicas in corde tuo: Appropinquat septimus annus remissionis", et avertas oculos tuos a paupere fratre tuo nolens ei, quod postulat, mutuum commodare, ne clamet contra te ad Dominum, et fiat tibi in peccatum.
DEUT|15|10|Sed dabis ei, nec contristabitur cor tuum in eius necessitatibus sublevandis, nam propter hoc benedicet tibi Dominus Deus tuus in omni opere tuo et in cunctis, ad quae manum miseris.
DEUT|15|11|Non deerunt pauperes in terra habitationis tuae; idcirco ego praecipio tibi, ut aperias manum fratri tuo egeno et pauperi, qui tecum versatur in terra tua.
DEUT|15|12|Cum tibi venditus fuerit frater tuus Hebraeus aut Hebraea et sex annis servierit tibi, in septimo anno dimittes eum liberum;
DEUT|15|13|et quem libertate donaveris, nequaquam vacuum abire patieris.
DEUT|15|14|Sed dabis ei viaticum de gregibus et de area et torculari tuo, quibus Dominus Deus tuus benedixerit tibi.
DEUT|15|15|Memento quod et ipse servieris in terra Aegypti, et liberaverit te Dominus Deus tuus; idcirco ego nunc hoc praecipio tibi.
DEUT|15|16|Sin autem dixerit: "Nolo egredi", eo quod diligat te et domum tuam et bene sibi apud te esse sentiat,
DEUT|15|17|assumes subulam et perforabis aurem eius in ianua domus tuae, et serviet tibi usque in aeternum. Ancillae quoque similiter facies.
DEUT|15|18|Non sit durum in oculis tuis dimittere eum liberum, quoniam iuxta mercedem mercennarii per sex annos servivit tibi, et benedicet tibi Dominus Deus tuus in cunctis operibus, quae egeris.
DEUT|15|19|De primogenitis, quae nascuntur in armentis et ovibus tuis, quidquid sexus est masculini, sanctificabis Domino Deo tuo; non operaberis in primogenito bovis et non tondebis primogenita ovium.
DEUT|15|20|In conspectu Domini Dei tui comedes ea per annos singulos in loco, quem elegerit Dominus, tu et domus tua.
DEUT|15|21|Sin autem habuerit maculam et vel claudum fuerit vel caecum aut in aliqua parte deforme vel debile, non immolabis illud Domino Deo tuo,
DEUT|15|22|sed intra portas tuas comedes illud; tam mundus quam immundus similiter vescentur eis, quasi caprea et cervo.
DEUT|15|23|Solum sanguinem eorum non comedes, sed effundes in terram quasi aquam.
DEUT|16|1|Observa mensem Abib, ut facias Pascha Domino Deo tuo; quoniam in isto mense Abib eduxit te Dominus Deus tuus de Aegypto nocte.
DEUT|16|2|Immolabisque Pascha Domino Deo tuo de ovibus et de bobus in loco, quem elegerit Dominus Deus tuus, ut habitet nomen eius ibi.
DEUT|16|3|Non comedes cum eo panem fermentatum; septem diebus comedes absque fermento afflictionis panem, quoniam festinanter egressus es de Aegypto, ut memineris diei egressionis tuae de Aegypto omnibus diebus vitae tuae.
DEUT|16|4|Non apparebit fermentum in omnibus terminis tuis septem diebus; et non manebit de carnibus eius, quod immolatum est vespere in die primo, usque mane.
DEUT|16|5|Non poteris immolare Pascha in qualibet urbium tuarum, quas Dominus Deus tuus daturus est tibi,
DEUT|16|6|sed in loco, quem elegerit Dominus Deus tuus, ut habitet nomen eius ibi, immolabis Pascha vespere ad solis occasum, quando egressus es de Aegypto.
DEUT|16|7|Et coques et comedes in loco, quem elegerit Dominus Deus tuus, maneque consurgens vades in tabernacula tua.
DEUT|16|8|Sex diebus comedes azyma et in die septimo, quia collecta est Domino Deo tuo, non facies opus.
DEUT|16|9|Septem hebdomadas numerabis tibi ab ea die, qua falcem in segetem miseris,
DEUT|16|10|et celebrabis diem festum Hebdomadarum Domino Deo tuo, oblationem spontaneam manus tuae, quam offeres iuxta benedictionem Domini Dei tui.
DEUT|16|11|Et epulaberis coram Domino Deo tuo tu, filius tuus et filia tua, servus tuus et ancilla tua et Levites, qui est intra portas tuas, advena ac pupillus et vidua, qui morantur tecum in loco, quem elegerit Dominus Deus tuus, ut habitet nomen eius ibi;
DEUT|16|12|et recordaberis quoniam servus fueris in Aegypto custodiesque ac facies, quae praecepta sunt.
DEUT|16|13|Sollemnitatem quoque Tabernaculorum celebrabis per septem dies, quando collegeris de area et torculari fruges tuas;
DEUT|16|14|et epulaberis in festivitate tua tu, filius tuus et filia, servus tuus et ancilla, Levites quoque et advena, pupillus ac vidua, qui intra portas tuas sunt.
DEUT|16|15|Septem diebus Domino Deo tuo festa celebrabis in loco, quem elegerit Dominus, quia benedicet tibi Dominus Deus tuus in cunctis frugibus tuis et in omni opere manuum tuarum, erisque totus in laetitia.
DEUT|16|16|Tribus vicibus per annum apparebit omne masculinum tuum in conspectu Domini Dei tui in loco, quem elegerit: in sollemnitate Azymorum et in sollemnitate Hebdomadarum et in sollemnitate Tabernaculorum. Non apparebit ante Dominum vacuus,
DEUT|16|17|sed offeret unusquisque secundum quod habuerit, iuxta benedictionem Domini Dei tui, quam dederit tibi.
DEUT|16|18|Iudices et praefectos operum constitues in omnibus portis tuis, quas Dominus Deus tuus dederit tibi per singulas tribus tuas, ut iudicent populum iusto iudicio.
DEUT|16|19|Non declinabis iudicium. Non accipies personam nec munera, quia munera excaecant oculos sapientum et mutant causas iustorum.
DEUT|16|20|Iustitiam, iustitiam persequeris, ut vivas et possideas terram, quam Dominus Deus tuus dederit tibi.
DEUT|16|21|Non plantabis tibi palum, omnem arborem iuxta altare Domini Dei tui, quod feceris tibi.
DEUT|16|22|Neque constitues lapidem, quem odit Dominus Deus tuus.
DEUT|17|1|Non immolabis Domino Deo tuo ovem et bovem, in quo est macula aut quippiam vitii, quia abominatio est Domino Deo tuo.
DEUT|17|2|Cum reperti fuerint apud te intra unam portarum tuarum, quas Dominus Deus tuus dabit tibi, vir aut mulier, qui faciant, quod malum est in conspectu Domini Dei tui, et transgrediantur pactum illius,
DEUT|17|3|ut vadant et serviant diis alienis et adorent eos, solem vel lunam vel omnem militiam caeli, quae non praecepi,
DEUT|17|4|et hoc tibi fuerit nuntiatum, audiensque inquisieris diligenter et verum esse reppereris, et abominatio haec facta est in Israel,
DEUT|17|5|educes virum vel mulierem, qui hanc rem sceleratissimam perpetrarunt, ad portas civitatis tuae, et lapidibus obruentur.
DEUT|17|6|In ore duorum aut trium testium peribit, qui interficietur; nemo occidatur uno contra se dicente testimonium.
DEUT|17|7|Manus testium prima erit ad interficiendum eum, et manus reliqui populi extrema mittetur, ut auferas malum de medio tui.
DEUT|17|8|Si intra portas tuas in litibus difficile et ambiguum apud te iudicium esse perspexeris inter sanguinem et sanguinem, causam et causam, plagam et plagam, surge et ascende ad locum, quem elegerit Dominus Deus tuus,
DEUT|17|9|veniesque ad sacerdotes levitici generis et ad iudicem, qui fuerit illo tempore; quaeresque ab eis, qui indicabunt tibi iudicii sententiam.
DEUT|17|10|Et facies quodcumque dixerint tibi de loco, quem elegerit Dominus, et observabis, ut facias omnia quae docuerint te
DEUT|17|11|iuxta mandatum, quod mandaverunt, et iuxta sententiam, quam dixerint tibi. Nec declinabis ad dexteram vel ad sinistram.
DEUT|17|12|Qui autem superbierit nolens oboedire sacerdotis imperio, qui eo tempore ministrat Domino Deo tuo, aut decreto iudicis, morietur homo ille, et auferes malum de Israel;
DEUT|17|13|cunctusque populus audiens timebit, ut nullus deinceps intumescat superbia.
DEUT|17|14|Cum ingressus fueris terram, quam Dominus Deus tuus dabit tibi, et possederis eam habitaverisque in illa et dixeris: "Constituam super me regem, sicut habent omnes per circuitum nationes",
DEUT|17|15|eum constitues super te regem, quem Dominus Deus tuus elegerit de numero fratrum tuorum. Non poteris alterius gentis hominem regem facere, qui non sit frater tuus.
DEUT|17|16|Tantummodo non multiplicabit sibi equos nec reducet populum in Aegyptum, ut equitatus numerum augeat, praesertim cum Dominus praeceperit vobis, ut nequaquam amplius per hanc viam revertamini.
DEUT|17|17|Neque habebit uxores plurimas, ne declinet cor eius, neque argenti et auri immensa pondera.
DEUT|17|18|Postquam autem sederit in solio regni sui, describet sibi exemplar legis huius in volumine accipiens illam a sacerdotibus leviticae tribus;
DEUT|17|19|et habebit secum legetque illud omnibus diebus vitae suae, ut discat timere Dominum Deum suum. et custodire verba legis huius et praecepta ista et quae in lege praecepta sunt.
DEUT|17|20|Nec elevetur cor eius in superbiam super fratres suos neque declinet a mandatis in partem dexteram vel sinistram, ut longo tempore regnet ipse et filii eius in medio Israel.
DEUT|18|1|Non habebunt sacerdotes le vitae, omnis tribus Levi, par tem et hereditatem cum reliquo Israel; de sacrificiis Domini et hereditate eius comedent
DEUT|18|2|et nihil accipient de possessione fratrum suorum: Dominus enim ipse est hereditas eorum, sicut locutus est illis.
DEUT|18|3|Hoc erit ius sacerdotum a populo, ab his qui offerunt victimas: sive bovem sive ovem immolaverint, dabunt sacerdoti armum et duas maxillas ac ventriculum,
DEUT|18|4|primitias frumenti, vini et olei et lanarum ex ovium tonsione.
DEUT|18|5|Ipsum enim elegit Dominus Deus tuus de cunctis tribubus tuis, ut stet et ministret in nomine Domini ipse et filii eius in sempiternum.
DEUT|18|6|Si exierit Levites de una urbium tuarum ex omni Israel, in qua ut advena habitat, et voluerit venire desiderans locum, quem elegerit Dominus,
DEUT|18|7|ministrabit in nomine Domini Dei sui, sicut omnes fratres eius levitae, qui stabunt ibi coram Domino.
DEUT|18|8|Partem ciborum eandem accipiet quam et ceteri, excepto eo, quod ex paterna ei successione debetur.
DEUT|18|9|Quando ingressus fueris terram, quam Dominus Deus tuus dabit tibi, cave, ne imitari velis abominationes illarum gentium.
DEUT|18|10|Nec inveniatur in te, qui filium suum aut filiam traducat per ignem, aut qui sortes sciscitetur et observet nubes atque auguria, nec sit maleficus
DEUT|18|11|nec incantator, nec qui pythones consulat nec divinos, aut quaerat a mortuis veritatem;
DEUT|18|12|omnia enim haec abominatur Dominus et propter istiusmodi scelera expellet eos in introitu tuo.
DEUT|18|13|Perfectus eris et absque macula cum Domino Deo tuo.
DEUT|18|14|Gentes istae, quarum possidebis terram, augures et divinos audiunt; tu autem a Domino Deo tuo aliter institutus es.
DEUT|18|15|Prophetam de gente tua et de fratribus tuis sicut me suscitabit tibi Dominus Deus tuus; ipsum audietis,
DEUT|18|16|ut petiisti a Domino Deo tuo in Horeb, quando contio congregata est, atque dixisti: "Ultra non audiam vocem Domini Dei mei et ignem hunc maximum amplius non videbo, ne moriar".
DEUT|18|17|Et ait Dominus mihi: "Bene omnia sunt locuti;
DEUT|18|18|prophetam suscitabo eis de medio fratrum suorum similem tui et ponam verba mea in ore eius, loqueturque ad eos omnia, quae praecepero illi.
DEUT|18|19|Qui autem verba mea, quae loquetur in nomine meo, audire noluerit, ego ultor exsistam.
DEUT|18|20|Propheta autem qui, arrogantia depravatus, voluerit loqui in nomine meo, quae ego non praecepi illi ut diceret, aut ex nomine alienorum deorum, interficietur".
DEUT|18|21|Quod si tacita cogitatione responderis: "Quomodo possum intellegere verbum, quod Dominus non est locutus?",
DEUT|18|22|hoc habebis signum: quod in nomine Domini propheta ille praedixerit, et non evenerit, hoc Dominus non est locutus, sed per tumorem animi sui propheta confinxit; et idcirco non timebis eum.
DEUT|19|1|Cum disperderit Dominus Deus tuus gentes, quarum ti bi traditurus est terram, et possederis eam habitaverisque in urbibus eius et in aedibus,
DEUT|19|2|tres civitates separabis tibi in medio terrae, quam Dominus Deus tuus dabit tibi in possessionem
DEUT|19|3|sternens diligenter viam; et in tres aequaliter partes totam terrae tuae provinciam divides, ut habeat e vicino, qui propter homicidium profugus est, quo possit evadere.
DEUT|19|4|Haec erit lex homicidae fugientis, cuius vita servanda est: qui percusserit proximum suum nesciens et qui heri et nudiustertius nullum contra eum habuisse odium comprobatur,
DEUT|19|5|sed abiisse cum eo simpliciter in silvam ad ligna caedenda, et in succisione lignorum securis fugerit manu, ferrumque lapsum de manubrio amicum eius percusserit et occiderit, hic ad unam supradictarum urbium confugiet et vivet;
DEUT|19|6|ne forsitan ultor sanguinis cordis calore stimulatus persequatur et apprehendat eum, si longior via fuerit, et percutiat eum, et moriatur, qui non est reus mortis, quia nullum contra eum, qui occisus est, odium prius habuisse monstratur.
DEUT|19|7|Idcirco praecipio tibi, ut tres civitates aequalis inter se spatii dividas.
DEUT|19|8|Cum autem dilataverit Dominus Deus tuus terminos tuos, sicut iuravit patribus tuis, et dederit tibi cunctam terram, quam eis pollicitus est
DEUT|19|9|- si tamen custodieris omne mandatum hoc et feceris, quae hodie praecipio tibi, ut diligas Dominum Deum tuum et ambules in viis eius omni tempore - addes tibi tres alias civitates et supradictarum trium urbium numerum duplicabis,
DEUT|19|10|ut non effundatur sanguis innoxius in medio terrae, quam Dominus Deus tuus dabit tibi possidendam, nec sis sanguinis reus.
DEUT|19|11|Si quis autem odio habens proximum suum insidiatus fuerit vitae eius surgensque percusserit illum, et mortuus fuerit, fugeritque ad unam de supradictis urbibus,
DEUT|19|12|mittent seniores civitatis eius et arripient eum de loco effugii tradentque in manu ultoris sanguinis, et morietur:
DEUT|19|13|non misereberis eius et auferes innoxium sanguinem de Israel, ut bene sit tibi.
DEUT|19|14|Non transferes terminos proximi tui, quos fixerunt priores in possessione tua, quam acceperis in terra, quam Dominus Deus tuus dabit tibi possidendam.
DEUT|19|15|Non stabit testis unus contra aliquem, quidquid illius peccatum vel facinus fuerit; sed in ore duorum aut trium testium stabit omne verbum.
DEUT|19|16|Si steterit testis mendax contra hominem accusans eum praevaricationis,
DEUT|19|17|stabunt ambo, quorum causa est, ante Dominum in conspectu sacerdotum et iudicum, qui fuerint in diebus illis.
DEUT|19|18|Cumque diligentissime perscrutantes iudices invenerint falsum testem dixisse contra fratrem suum mendacium,
DEUT|19|19|reddent ei, sicut fratri suo facere cogitavit, et auferes malum de medio tui,
DEUT|19|20|ut audientes ceteri timorem habeant et nequaquam ultra talia audeant facere in medio tui.
DEUT|19|21|Non misereberis eius, sed animam pro anima, oculum pro oculo, dentem pro dente, manum pro manu, pedem pro pede exiges.
DEUT|20|1|Si exieris ad bellum contra hostes tuos et videris equita tus et currus et maiorem, quam tu habes, adversarii exercitus multitudinem, non timebis eos, quia Dominus Deus tuus tecum est, qui eduxit te de terra Aegypti.
DEUT|20|2|Appropinquante autem iam proelio, stabit sacerdos ante aciem et sic loquetur ad populum:
DEUT|20|3|"Audi, Israel: Vos hodie contra inimicos vestros pugnam committitis; non pertimescat cor vestrum, nolite metuere, nolite cedere nec formidetis eos,
DEUT|20|4|quia Dominus Deus vester incedit vobiscum et pro vobis contra adversarios vestros dimicabit, ut eruat vos de periculo".
DEUT|20|5|Praefecti quoque per singulas turmas, audiente exercitu, proclamabunt: Quis est homo, qui aedificavit domum novam et non dedicavit eam? Vadat et revertatur in domum suam, ne forte moriatur in bello, et alius dedicet illam.
DEUT|20|6|Quis est homo, qui plantavit vineam et necdum vindemiavit eam? Vadat et revertatur in domum suam, ne forte moriatur in bello, et alius homo vindemiet illam.
DEUT|20|7|Quis est homo, qui despondit uxorem et non accepit eam? Vadat et revertatur in domum suam, ne forte moriatur in bello, et alius homo accipiat eam".
DEUT|20|8|His dictis, addent reliqua et loquentur ad populum: "Quis est homo formidulosus et corde pavido? Vadat et revertatur in domum suam, ne pavere faciat corda fratrum suorum, sicut ipse timore perterritus est".
DEUT|20|9|Cumque praefecti finem loquendi ad populum fecerint, constituantur duces exercitus in capite populi.
DEUT|20|10|Si quando accesseris ad expugnandam civitatem, offeres ei primum pacem;
DEUT|20|11|si receperit et aperuerit tibi portas, cunctus populus, qui in ea est, serviet tibi sub tributo.
DEUT|20|12|Sin autem foedus inire noluerit et coeperit contra te bellum, oppugnabis eam.
DEUT|20|13|Cumque tradiderit Dominus Deus tuus illam in manu tua, percuties omne, quod in ea generis masculini est, in ore gladii
DEUT|20|14|absque mulieribus et infantibus, iumentis et ceteris, quae in civitate sunt. Omnem praedam hanc diripies tibi et comedes de spoliis hostium tuorum, quae Dominus Deus tuus dederit tibi.
DEUT|20|15|Sic facies cunctis civitatibus, quae a te procul valde sunt et non sunt de gentium istarum urbibus, quas in possessionem accepturus es.
DEUT|20|16|De his autem civitatibus, quae dabuntur tibi, nullum omnino permittes vivere,
DEUT|20|17|sed interficies in ore gladii, Hetthaeum videlicet et Amorraeum et Chananaeum, Pherezaeum et Hevaeum et Iebusaeum, sicut praecepit tibi Dominus Deus tuus,
DEUT|20|18|ne forte doceant vos facere cunctas abominationes, quas ipsi operati sunt diis suis, et peccetis in Dominum Deum vestrum.
DEUT|20|19|Quando obsederis civitatem multo tempore et munitionibus circumdederis, ut expugnes eam, non immittes securim in arbores eius, de quibus vesci potes, nec succidas eas. Numquid homo est arbor campi, ut eam obsideas?
DEUT|20|20|Si qua autem ligna non sunt pomifera, succide illa et exstrue machinas, donec capias civitatem, quae contra te dimicat.
DEUT|21|1|Quando inventum fuerit in terra, quam Dominus Deus tuus daturus est tibi, hominis cadaver occisi, et ignoratur caedis reus,
DEUT|21|2|egredientur maiores natu et iudices tui et metientur a loco cadaveris singularum per circuitum spatia civitatum
DEUT|21|3|et, quam viciniorem ceteris esse perspexerint, seniores civitatis illius tollent vitulam de armento, quae non traxit iugum nec terram scidit vomere,
DEUT|21|4|et ducent eam ad torrentem perennem, ubi numquam aratum est nec seminatum, et caedent apud eum cervices vitulae;
DEUT|21|5|accedentque sacerdotes filii Levi, quos elegerit Dominus Deus tuus, ut ministrent ei et benedicant in nomine eius, et ad verbum eorum omnis causa et omnis percussio iudicetur.
DEUT|21|6|Et omnes maiores natu civitatis illius, qui prope interfectum sunt, lavabunt manus suas super vitulam, quae apud torrentem percussa est,
DEUT|21|7|et dicent: "Manus nostrae non effuderunt hunc sanguinem, nec oculi nostri viderunt;
DEUT|21|8|propitius esto populo tuo Israel, quem redemisti, Domine, et non reputes sanguinem innocentem in medio populi tui Israel". Et auferetur ab eis reatus sanguinis.
DEUT|21|9|Tu autem removebis innocentem cruorem, cum feceris, quod rectum est in oculis Domini.
DEUT|21|10|Si egressus fueris ad pugnam contra inimicos tuos, et tradiderit eos Dominus Deus tuus in manu tua, captivosque duxeris
DEUT|21|11|et videris in numero captivorum mulierem pulchram et adamaveris eam voluerisque habere uxorem,
DEUT|21|12|introduces eam in domum tuam. Quae radet caesariem et circumcidet ungues
DEUT|21|13|et deponet vestem captivitatis sedensque in domo tua flebit patrem et matrem suam uno mense; et postea intrabis ad eam sociaberisque illi, et erit uxor tua.
DEUT|21|14|Sin autem postea non sederit animo tuo, dimittes eam liberam; nec vendere poteris pecunia nec opprimere per potentiam, quia humiliasti eam.
DEUT|21|15|Si habuerit homo uxores duas, unam dilectam et alteram odiosam, genuerintque ei liberos, et fuerit filius odiosae primogenitus,
DEUT|21|16|volueritque substantiam inter filios suos dividere, non poterit filium dilectae facere primogenitum et praeferre filio odiosae,
DEUT|21|17|sed filium odiosae agnoscet primogenitum dabitque ei de cunctis, quae habuerit, duplicia; iste est enim principium roboris eius, et huic debentur primogenita.
DEUT|21|18|Si genuerit homo filium contumacem et protervum, qui non audiat patris aut matris imperium et coercitus oboedire contempserit,
DEUT|21|19|apprehendent eum et ducent ad seniores civitatis suae et ad portam iudicii
DEUT|21|20|dicentque ad eos: "Filius noster iste protervus et contumax est: monita nostra audire contemnit, comissationibus vacat et luxuriae atque conviviis potatorum".
DEUT|21|21|Lapidibus eum obruent viri civitatis, et morietur, ut auferatis malum de medio vestri, et universus Israel audiens pertimescat.
DEUT|21|22|Quando peccaverit homo, quod morte plectendum est, et occisum appenderis in patibulo,
DEUT|21|23|non permanebit cadaver eius in ligno; sed in eadem die sepelietur, quia maledictus a Deo est, qui pendet in ligno; et nequaquam contaminabis terram tuam, quam Dominus Deus tuus dederit tibi in possessionem.
DEUT|22|1|Non videbis bovem fratris tui aut ovem errantem et praeteribis, sed reduces fratri tuo;
DEUT|22|2|si autem non est prope frater tuus nec nosti eum, duces in domum tuam, et erunt apud te quamdiu quaerat ea frater tuus et recipiat.
DEUT|22|3|Similiter facies de asino et de vestimento et de omni re fratris tui, quae perierit: si inveneris eam, ne subtrahas te.
DEUT|22|4|Si videris asinum fratris tui aut bovem cecidisse in via, non subtrahes te, sed sublevabis cum eo.
DEUT|22|5|Non induetur mulier veste virili, nec vir utetur veste feminea: abominabilis enim apud Dominum Deum tuum est omnis, qui facit haec.
DEUT|22|6|Si ambulans per viam, in arbore vel in terra nidum avis inveneris et matrem pullis vel ovis desuper incubantem, non sumes eam de filiis,
DEUT|22|7|sed abire patieris matrem tenens filios, ut bene sit tibi, et longo vivas tempore.
DEUT|22|8|Cum aedificaveris domum novam, facies murum tecto tuo per circuitum, ne adducas sanguinem super domum tuam et sis reus, labente aliquo in praeceps ruente.
DEUT|22|9|Non seres vineam tuam altero semine, ne et sementis, quam sevisti, et quae nascuntur ex vinea, pariter sanctificentur.
DEUT|22|10|Non arabis in bove simul et asino.
DEUT|22|11|Non indueris vestimento, quod ex lana linoque contextum est.
DEUT|22|12|Funiculos facies per quattuor angulos pallii tui, quo operieris.
DEUT|22|13|Si duxerit vir uxorem et intraverit ad eam et postea odio habuerit eam
DEUT|22|14|imputaveritque ei obiciens ei nomen pessimum et dixerit: "Uxorem hanc accepi et ingressus ad eam non inveni virginem",
DEUT|22|15|tollent pater et mater eius et ferent secum signa virginitatis eius ad seniores urbis, qui in porta sunt,
DEUT|22|16|et dicet pater: "Filiam meam dedi huic uxorem, quam, quia odit,
DEUT|22|17|imponit ei nomen pessimum, ut dicat: Non inveni filiam tuam virginem; et ecce haec sunt signa virginitatis filiae meae". Expandent vestimentum coram se nioribus civitatis.
DEUT|22|18|Apprehendentque senes urbis illius virum et verberabunt illum
DEUT|22|19|condemnantes insuper centum siclis argenti, quos dabunt patri puellae, quoniam diffamavit nomen pessimum super virginem Israel; habebitque eam uxorem et non poterit dimittere eam omnibus diebus vitae suae.
DEUT|22|20|Quod si verum est, quod obicit, et non est in puella inventa virginitas,
DEUT|22|21|educent eam ad fores domus patris sui, et lapidibus obruent viri civitatis eius, et morietur, quoniam fecit nefas in Israel, ut fornicaretur in domo patris sui; et auferes malum de medio tui.
DEUT|22|22|Si inventus fuerit vir dormiens cum uxore alterius, uterque morietur, id est adulter et adultera; et auferes malum de Israel.
DEUT|22|23|Si puellam virginem desponsatam viro invenerit aliquis in civitate et concubuerit cum illa,
DEUT|22|24|educetis utrumque ad portam civitatis illius et lapidibus obruetis, et morientur: puella quia non clamavit, cum esset in civitate, vir quia humiliavit uxorem proximi sui; et auferes malum de medio tui.
DEUT|22|25|Sin autem in agro reppererit vir puellam, quae desponsata est, et apprehendens concubuerit cum illa, ipse morietur solus;
DEUT|22|26|puella nihil patietur nec est rea mortis, quoniam sicut vir consurgit contra fratrem suum et occidit eum, ita et puella perpessa est:
DEUT|22|27|sola erat in agro, clamavit puella desponsata, et nullus affuit, qui liberaret eam.
DEUT|22|28|Si invenerit vir puellam virginem, quae non habet sponsum, et apprehendens concubuerit cum ea, et res ad iudicium venerit,
DEUT|22|29|dabit, qui dormivit cum ea, patri puellae quinquaginta siclos argenti et habebit eam uxorem, quia humiliavit illam: non poterit dimittere eam cunctis diebus vitae suae.
DEUT|23|1|Non accipiet homo uxorem patris sui nec revelabit operi mentum eius.
DEUT|23|2|Non intrabit eunuchus, attritis vel amputatis testiculis et absciso veretro, ecclesiam Domini.
DEUT|23|3|Non ingredietur mamzer in ecclesiam Domini neque decima generatione.
DEUT|23|4|Ammonites et Moabites etiam in decima generatione non intrabunt ecclesiam Domini in aeternum,
DEUT|23|5|quia noluerunt vobis occurrere cum pane et aqua in via, quando egressi estis de Aegypto, et quia conduxerunt contra te Balaam filium Beor de Phethor in Aramnaharaim, ut malediceret tibi;
DEUT|23|6|et noluit Dominus Deus tuus audire Balaam vertitque tibi maledictionem eius in benedictionem, eo quod diligeret te.
DEUT|23|7|Non facies cum eis pacem nec quaeres eis bona cunctis diebus vitae tuae in sempiternum.
DEUT|23|8|Non abominaberis Idumaeum, quia frater tuus est, nec Aegyptium, quia advena fuisti in terra eius:
DEUT|23|9|qui nati fuerint ex eis tertia generatione, intrabunt ecclesiam Domini.
DEUT|23|10|Quando egressus fueris adversus hostes tuos in pugnam, custodies te ab omni re mala.
DEUT|23|11|Si fuerit apud te homo, qui nocturno pollutus sit somnio, egredietur extra castra et non revertetur,
DEUT|23|12|priusquam ad vesperam lavetur aqua; et ad solis occasum regredietur in castra.
DEUT|23|13|Habebis locum extra castra, ad quem egrediaris ad requisita naturae
DEUT|23|14|gerens paxillum in balteo; cumque sederis foris, fodies foveam et egesta humo operies.
DEUT|23|15|Dominus enim Deus tuus ambulat in medio castrorum tuorum, ut eruat te et tradat tibi inimicos tuos; sint castra tua sancta, et nihil in eis videat foeditatis nec derelinquat te.
DEUT|23|16|Non trades servum domino suo, qui ad te confugerit:
DEUT|23|17|habitabit tecum in medio tui in loco, quem elegerit in una urbium tuarum, quae placuerit ei, nec contristes eum.
DEUT|23|18|Non erit prostibulum sacrum de filiabus Israel, nec scortator sacer de filiis Israel.
DEUT|23|19|Non offeres mercedem prostibuli nec pretium canis in domo Domini Dei tui, quidquid illud est, quod voveris, quia abominatio est utrumque apud Dominum Deum tuum.
DEUT|23|20|Non fenerabis fratri tuo ad usuram pecuniam nec alimenta nec quamlibet aliam rem,
DEUT|23|21|sed alieno fenerabis. Fratri autem tuo absque usura id, quo indiget, commodabis, ut benedicat tibi Dominus Deus tuus in omni opere tuo in terra, ad quam ingredieris possidendam.
DEUT|23|22|Cum voveris votum Domino Deo tuo, non tardabis reddere; quia requiret illud Dominus Deus tuus a te, et reputabitur tibi in peccatum.
DEUT|23|23|Si nolueris polliceri, absque peccato eris;
DEUT|23|24|quod autem egressum est de labiis tuis, observabis et facies, sicut promisisti Domino Deo tuo: propria voluntate et ore tuo locutus es.
DEUT|23|25|Ingressus vineam proximi tui comede uvas, quantum tibi placuerit; in sporta autem ne efferas tecum.
DEUT|23|26|Si intraveris in segetem amici tui, franges spicas manu; falce autem non metes.
DEUT|24|1|Si acceperit homo uxorem et habuerit eam, et non invene rit gratiam ante oculos eius propter aliquam foeditatem, et scripserit libellum repudii dederitque in manu illius et dimiserit eam de domo sua,
DEUT|24|2|cumque egressa alterius uxor facta fuerit,
DEUT|24|3|et ille quoque oderit eam dederitque ei libellum repudii et dimiserit de domo sua, vel mortuus fuerit,
DEUT|24|4|non poterit prior maritus recipere eam in uxorem, quia polluta est; hoc esset abominatio coram Domino. Ne peccare facias terram tuam, quam Dominus Deus tuus tradiderit tibi possidendam.
DEUT|24|5|Cum acceperit homo nuper uxorem, non procedet ad bellum, nec ei quippiam necessitatis iniungetur publicae, sed vacabit liber domui suae, ut uno anno laetetur cum uxore sua.
DEUT|24|6|Non accipies loco pignoris molam vel superiorem lapidem molarem, quia animam suam apposuit tibi.
DEUT|24|7|Si deprehensus fuerit homo rapiens unum de fratribus suis de filiis Israel et, vendito eo, accipiens pretium, interficietur; et auferes malum de medio tui.
DEUT|24|8|Observa diligenter, si incurras plagam leprae, quaecumque docuerint vos sacerdotes levitici generis; quod praecepi eis, implete sollicite.
DEUT|24|9|Memento, quae fecerit Dominus Deus tuus Mariae in via, cum egrederemini de Aegypto.
DEUT|24|10|Cum mutuam dabis proximo tuo rem aliquam, non ingredieris domum eius, ut pignus auferas,
DEUT|24|11|sed stabis foris, et ille tibi pignus proferet, quod habuerit.
DEUT|24|12|Sin autem pauper est, non pernoctabit apud te pignus,
DEUT|24|13|sed statim reddes ei ad solis occasum, ut dormiens in vestimento suo benedicat tibi, et habeas iustitiam coram Domino Deo tuo.
DEUT|24|14|Non negabis mercedem indigentis et pauperis ex fratribus tuis sive advenis, qui tecum morantur in terra intra portas tuas,
DEUT|24|15|sed eadem die reddes ei pretium laboris sui ante solis occasum, quia pauper est, et illud desiderat anima sua; ne clamet contra te ad Dominum, et reputetur tibi in peccatum.
DEUT|24|16|Non occidentur patres pro filiis, nec filii pro patribus, sed unusquisque pro peccato suo morietur.
DEUT|24|17|Non pervertes iudicium advenae et pupilli nec auferes pignoris loco viduae vestimentum.
DEUT|24|18|Memento quod servieris in Aegypto, et eruerit te Dominus Deus tuus inde; idcirco praecipio tibi, ut facias hanc rem.
DEUT|24|19|Quando messueris segetem in agro tuo et oblitus manipulum reliqueris, non reverteris, ut tollas eum, sed advenam et pupillum et viduam auferre patieris, ut benedicat tibi Dominus Deus tuus in omni opere manuum tuarum.
DEUT|24|20|Si fruges collegeris olivarum, quidquid remanserit in arboribus, non reverteris, ut colligas, sed relinques advenae, pupillo ac viduae.
DEUT|24|21|Si vindemiaveris vineam tuam, non colliges remanentes racemos, sed cedent in usus advenae, pupilli ac viduae.
DEUT|24|22|Memento quod et tu servieris in Aegypto; et idcirco praecipio tibi, ut facias hanc rem.
DEUT|25|1|Si fuerit causa inter aliquos, et interpellaverint iudices, quem iustum esse perspexerint, illi iustitiae palmam dabunt; quem impium, condemnabunt impietatis.
DEUT|25|2|Sin autem iudex eum, qui peccavit, dignum viderit plagis, prosternet et coram se faciet verberari; pro mensura peccati erit et plagarum modus,
DEUT|25|3|ita dumtaxat, ut quadragenarium numerum non excedant, ne ultra percussus plagis multis et foede laceratus ante oculos tuos abeat frater tuus.
DEUT|25|4|Non ligabis os bovis terentis in area fruges tuas.
DEUT|25|5|Quando habitaverint fratres simul, et unus ex eis absque filio mortuus fuerit, uxor defuncti non nubet foras alteri, sed accipiet eam frater eius uxorem et suscitabit semen fratris sui;
DEUT|25|6|et primogenitum ex ea filium nomine illius appellabit, ut non deleatur nomen eius ex Israel.
DEUT|25|7|Sin autem noluerit accipere uxorem fratris sui, quae ei lege debetur, perget mulier ad portam civitatis et interpellabit maiores natu dicetque: Non vult frater viri mei suscitare nomen fratris sui in Israel nec me in coniugium sumere";
DEUT|25|8|statimque accersiri eum facient et interrogabunt. Si responderit: "Nolo eam uxorem accipere",
DEUT|25|9|accedet mulier ad eum coram senioribus et tollet calceamentum de pede eius spuetque in faciem illius et dicet: "Sic fit homini, qui non aedificat domum fratris sui".
DEUT|25|10|Et vocabitur nomen illius in Israel: "Domus discalceati".
DEUT|25|11|Si habuerint inter se iurgium viri, et unus contra alterum rixari coeperit, volensque uxor alterius eruere virum suum de manu fortioris, miserit manum et apprehenderit verenda eius,
DEUT|25|12|abscides manum illius nec flecteris super eam ulla misericordia.
DEUT|25|13|Non habebis in sacculo tuo diversa pondera maius et minus;
DEUT|25|14|nec erit in domo tua ephi maius et minus.
DEUT|25|15|Pondus habebis iustum et verum, et ephi iustum et verum erit tibi, ut multo vivas tempore super terram, quam Dominus Deus tuus dederit tibi.
DEUT|25|16|Abominatur enim Dominus tuus eum, qui facit haec, et aversatur omnem iniustitiam.
DEUT|25|17|Memento quae fecerit tibi Amalec in via, quando egrediebaris ex Aegypto;
DEUT|25|18|quomodo occurrerit tibi et omnes extremos agminis tui, qui lassi residebant, ceciderit, quando tu eras fame et labore confectus, et non timuerit Deum.
DEUT|25|19|Cum ergo Dominus Deus tuus dederit tibi requiem a cunctis per circuitum inimicis tuis in terra, quam tibi daturus est, delebis nomen Amalec sub caelo: cave, ne obliviscaris!
DEUT|26|1|Cumque intraveris terram, quam Dominus Deus tuus ti bi daturus est possidendam, et obtinueris eam atque habitaveris in illa,
DEUT|26|2|tolles primitias de cunctis frugibus agri, quas collegeris de terra tua, quam Dominus Deus tuus dabit tibi, et pones in cartallo pergesque ad locum, quem Dominus Deus tuus elegerit, ut ibi habitet nomen eius,
DEUT|26|3|accedesque ad sacerdotem, qui fuerit in diebus illis, et dices ad eum: Profiteor hodie coram Domino Deo tuo quod ingressus sim terram, pro qua iuravit patribus nostris, ut daret eam nobis".
DEUT|26|4|Suscipiensque sacerdos cartallum de manu tua ponet ante altare Domini Dei tui,
DEUT|26|5|et loqueris in conspectu Domini Dei tui: "Syrus vagus erat pater meus et descendit in Aegyptum et ibi peregrinatus est in paucissimo numero; crevitque in gentem magnam ac robustam et infinitae multitudinis.
DEUT|26|6|Afflixeruntque nos Aegyptii et persecuti sunt imponentes onera gravissima.
DEUT|26|7|Et clamavimus ad Dominum, Deum patrum nostrorum, qui exaudivit nos et respexit humilitatem nostram et laborem atque angustias,
DEUT|26|8|et eduxit nos Dominus de Aegypto in manu forti et brachio extento, in ingenti pavore, in signis atque portentis,
DEUT|26|9|et introduxit ad locum istum et tradidit nobis terram hanc lacte et melle manantem.
DEUT|26|10|Et ecce nunc attuli primitias frugum terrae, quam dedisti mihi, Domine". Et dimittes eas in conspectu Domini Dei tui et adorato Domino Deo tuo.
DEUT|26|11|Et epulaberis in omnibus bonis, quae Dominus Deus tuus dederit tibi et domui tuae, tu et Levites et advena, qui tecum est.
DEUT|26|12|Quando compleveris decimam cunctarum frugum tuarum, anno tertio, anno decimarum, et dederis Levitae et advenae et pupillo et viduae, ut comedant intra portas tuas et saturentur,
DEUT|26|13|loqueris in conspectu Domini Dei tui: "Abstuli, quod sanctificatum est, de domo mea et dedi illud Levitae et advenae, pupillo ac viduae, sicut iussisti mihi; non praeterivi mandata tua nec sum oblitus imperii tui,
DEUT|26|14|non comedi ex eis in luctu meo nec separavi ex eis in qualibet immunditia nec expendi ex his quidquam mortuo: oboedivi voci Domini Dei mei et feci omnia, sicut praecepisti mihi.
DEUT|26|15|Respice de habitaculo sancto tuo, de caelo, et benedic populo tuo Israel et terrae, quam dedisti nobis, sicut iurasti patribus nostris, terrae lacte et melle mananti".
DEUT|26|16|Hodie Dominus Deus tuus mandavit tibi, ut facias praecepta haec atque iudicia et custodias et impleas illa ex toto corde tuo et ex tota anima tua.
DEUT|26|17|Dominum elegisti hodie, ut sit tibi Deus, et ambules in viis eius et custodias praecepta illius et mandata atque iudicia et oboedias eius imperio;
DEUT|26|18|et Dominus elegit te hodie, ut sis ei populus peculiaris, sicut locutus est tibi, et custodias omnia mandata illius,
DEUT|26|19|et faciat te excelsiorem cunctis gentibus, quas creavit in laudem et nomen et gloriam suam, ut sis populus sanctus Domini Dei tui, sicut locutus est ".
DEUT|27|1|Praecepit autem Moyses et seniores Israel populo dicen tes: " Custodite omne mandatum, quod praecipio vobis hodie.
DEUT|27|2|Cumque transieritis Iordanem in terram, quam Dominus Deus tuus dabit tibi, eriges ingentes lapides et calce obduces eos,
DEUT|27|3|ut possis in eis scribere omnia verba legis huius, Iordane transmisso, ut introeas terram, quam Dominus Deus tuus dabit tibi, terram lacte et melle manantem, sicut locutus est Dominus, Deus patrum tuorum, tibi.
DEUT|27|4|Quando ergo transieritis Iordanem, erigite istos lapides, sicut ego hodie praecipio vobis, in monte Hebal, et obduces eos calce;
DEUT|27|5|et aedificabis ibi altare Domino Deo tuo de lapidibus, quos ferrum non tetigit,
DEUT|27|6|de saxis impolitis, et offeres super eo holocausta Domino Deo tuo.
DEUT|27|7|Et immolabis hostias pacificas comedesque ibi et epulaberis coram Domino Deo tuo;
DEUT|27|8|et scribes super lapides omnia verba legis huius plane et lucide ".
DEUT|27|9|Dixeruntque Moyses et sacerdotes levitici generis ad omnem Israelem: " Attende et audi, Israel: hodie factus es populus Domino Deo tuo;
DEUT|27|10|audies vocem eius et facies mandata atque praecepta, quae ego praecipio tibi ".
DEUT|27|11|Praecepitque Moyses populo in die illo dicens:
DEUT|27|12|" Hi stabunt ad benedicendum populo super montem Garizim, Iordane transmisso: Simeon, Levi, Iudas, Issachar, Ioseph et Beniamin.
DEUT|27|13|Et e regione isti stabunt ad maledicendum in monte Hebal: Ruben, Gad et Aser et Zabulon, Dan et Nephthali.
DEUT|27|14|Et pronunciabunt Levitae dicentque ad omnes viros Israel excelsa voce:
DEUT|27|15|"Maledictus homo, qui facit sculptile et conflatile, abominationem Domini, opus manuum artificum, ponetque illud in abscondito". Et respondebit omnis populus et dicet: "Amen".
DEUT|27|16|"Maledictus, qui contemnit patrem suum et matrem". Et dicet omnis populus: "Amen".
DEUT|27|17|"Maledictus, qui transfert terminos proximi sui". Et dicet omnis populus: "Amen".
DEUT|27|18|"Maledictus, qui errare facit caecum in itinere". Et dicet omnis populus: "Amen".
DEUT|27|19|"Maledictus, qui pervertit iudicium advenae, pupilli et viduae". Et dicet omnis populus: "Amen".
DEUT|27|20|"Maledictus, qui dormit cum uxore patris sui, quia revelat operimentum lectuli eius". Et dicet omnis populus: "Amen".
DEUT|27|21|"Maledictus, qui dormit cum omni iumento". Et dicet omnis populus: Amen".
DEUT|27|22|"Maledictus, qui dormit cum sorore sua, filia patris sui sive matris suae". Et dicet omnis populus: "Amen".
DEUT|27|23|"Maledictus, qui dormit cum socru sua". Et dicet omnis populus: "Amen".
DEUT|27|24|"Maledictus, qui clam percusserit proximum suum". Et dicet omnis populus: "Amen".
DEUT|27|25|"Maledictus, qui accipit munera, ut percutiat sanguinem innocentem". Et dicet omnis populus: "Amen".
DEUT|27|26|"Maledictus, qui non permanet in sermonibus legis huius nec eos opere perficit". Et dicet omnis populus: "Amen".
DEUT|28|1|Sin audieris vocem Domini Dei tui, ut facias atque custo dias omnia mandata eius, quae ego praecipio tibi hodie, faciet te Dominus Deus tuus excelsiorem cunctis gentibus, quae versantur in terra,
DEUT|28|2|venientque super te universae benedictiones istae et apprehendent te, si tamen vocem Domini Dei tui audieris.
DEUT|28|3|Benedictus tu in civitate et benedictus in agro.
DEUT|28|4|Benedictus fructus ventris tui et fructus terrae tuae fructusque iumentorum tuorum, partus armentorum tuorum et incrementum ovium tuarum.
DEUT|28|5|Benedictum canistrum et pistrinum tuum.
DEUT|28|6|Benedictus eris et ingrediens et egrediens.
DEUT|28|7|Dabit Dominus inimicos tuos, qui consurgunt adversum te, corruentes in conspectu tuo; per unam viam venient contra te et per septem fugient a facie tua.
DEUT|28|8|Emittet Dominus benedictionem super cellaria tua et super omnia opera manuum tuarum; benedicetque tibi in terra, quam Dominus Deus tuus dabit tibi.
DEUT|28|9|Suscitabit te Dominus sibi in populum sanctum, sicut iuravit tibi, si custodieris mandata Domini Dei tui et ambulaveris in viis eius.
DEUT|28|10|Videbuntque omnes terrarum populi quod nomen Domini invocatum sit super te, et timebunt te.
DEUT|28|11|Abundare te faciet Dominus omnibus bonis, fructu uteri tui et fructu iumentorum tuorum, fructu terrae tuae, quam iuravit Dominus patribus tuis, ut daret tibi.
DEUT|28|12|Aperiet Dominus tibi thesaurum suum optimum, caelum, ut tribuat pluviam terrae tuae in tempore suo; benedicatque cunctis operibus manuum tuarum; et fenerabis gentibus multis et ipse a nullo fenus accipies.
DEUT|28|13|Constituet te Dominus in caput et non in caudam, et eris semper supra et non subter, si audieris mandata Domini Dei tui, quae ego praecipio tibi hodie, et custodieris et feceris
DEUT|28|14|ac non declinaveris a verbis, quae ego praecipio vobis hodie, nec ad dexteram nec ad sinistram, nec secutus fueris deos alienos neque colueris eos.
DEUT|28|15|Quod si audire nolueris vocem Domini Dei tui, ut custodias et facias omnia mandata eius et praecepta, quae ego praecipio tibi hodie, venient super te omnes maledictiones istae et apprehendent te:
DEUT|28|16|Maledictus eris in civitate, maledictus in agro.
DEUT|28|17|Maledictum canistrum et pistrinum tuum.
DEUT|28|18|Maledictus fructus ventris tui et fructus terrae tuae, partus armentorum tuorum et incrementum ovium tuarum.
DEUT|28|19|Maledictus eris ingrediens et maledictus egrediens.
DEUT|28|20|Mittet Dominus super te maledictionem et conturbationem et increpationem in omnia opera tua, quae facies, donec conterat te et perdat velociter propter adinventiones tuas pessimas, in quibus reliquisti me.
DEUT|28|21|Adiunget Dominus tibi pestilentiam, donec consumat te de terra, ad quam ingredieris possidendam.
DEUT|28|22|Percutiet te Dominus consumptione, febri et inflammatione, ardore et aestu, uredine ac aurugine, et persequentur te, donec pereas.
DEUT|28|23|Et erit caelum, quod est supra caput tuum, aeneum, et terra, quam calcas, ferrea.
DEUT|28|24|Convertet Dominus imbrem terrae tuae in pulverem, et de caelo descendet super te cinis, donec conteraris.
DEUT|28|25|Tradet te Dominus corruentem ante hostes tuos: per unam viam egredieris contra eos et per septem fugies et eris in terrorem omnibus regnis terrae.
DEUT|28|26|Eritque cadaver tuum in escam cunctis volatilibus caeli et bestiis terrae, et non erit qui abigat.
DEUT|28|27|Percutiet te Dominus ulcere Aegypti et tumore, scabie quoque et prurigine, ita ut curari nequeas.
DEUT|28|28|Percutiet te Dominus amentia et caecitate ac stupore mentis;
DEUT|28|29|et palpabis in meridie, sicut palpare solet caecus in tenebris, et non diriges vias tuas. Omnique tempore eris oppressus et exspoliatus nec habebis, qui liberet te.
DEUT|28|30|Uxorem accipies, et alius dormiet cum ea. Domum aedificabis et non habitabis in ea. Plantabis vineam et non vindemiabis eam.
DEUT|28|31|Bos tuus mactabitur coram te, et non comedes ex eo. Asinus tuus rapietur in conspectu tuo et non reddetur tibi. Oves tuae dabuntur inimicis tuis, et non erit qui te adiuvet.
DEUT|28|32|Filii tui et filiae tuae tradentur alteri populo, videntibus oculis tuis et deficientibus ad conspectum eorum tota die, et non erit fortitudo in manu tua.
DEUT|28|33|Fructus terrae tuae et omnes labores tuos comedet populus, quem ignoras, et eris semper oppressus et confractus cunctis diebus
DEUT|28|34|et insanies in aspectu eorum, quae videbunt oculi tui.
DEUT|28|35|Percutiet te Dominus ulcere pessimo in genibus et in suris, sanarique non poteris a planta pedis usque ad verticem tuum.
DEUT|28|36|Ducet te Dominus et regem tuum, quem constitueris super te, in gentem, quam ignorasti tu et patres tui, et servies ibi diis alienis, ligno et lapidi;
DEUT|28|37|et eris in stuporem et in proverbium ac fabulam omnibus populis, ad quos te introduxerit Dominus.
DEUT|28|38|Sementem multam iacies in terram et modicum congregabis, quia locustae devorabunt omnia.
DEUT|28|39|Vineas plantabis et coles et vinum non bibes nec colliges ex ea quippiam, quoniam vastabitur vermibus.
DEUT|28|40|Olivas habebis in omnibus terminis tuis et non ungeris oleo, quia defluent et peribunt.
DEUT|28|41|Filios generabis et filias et non frueris eis, quoniam ducentur in captivitatem.
DEUT|28|42|Omnes arbores tuas et fruges terrae tuae locusta consumet.
DEUT|28|43|Advena, qui tecum versatur in terra, ascendet super te eritque sublimior; tu autem descendes et eris inferior.
DEUT|28|44|Ipse fenerabit tibi, et tu non fenerabis ei; ipse erit in caput, et tu eris in caudam.
DEUT|28|45|Et venient super te omnes maledictiones istae et persequentes apprehendent te, donec intereas, quia non audisti vocem Domini Dei tui nec servasti mandata eius et praecepta, quae praecepit tibi.
DEUT|28|46|Et erunt in te signa atque prodigia et in semine tuo usque in sempiternum.
DEUT|28|47|Eo quod non servieris Domino Deo tuo in gaudio cordisque laetitia propter rerum omnium abundantiam,
DEUT|28|48|servies inimico tuo, quem immittet Dominus tibi, in fame et siti et nuditate et omnium penuria, et ponet iugum ferreum super cervicem tuam, donec te conterat.
DEUT|28|49|Adducet Dominus super te gentem de longinquo et de extremis finibus terrae in similitudinem aquilae volantis cum impetu, cuius linguam intellegere non possis:
DEUT|28|50|gentem procacissimam, quae non deferat seni nec misereatur parvulo;
DEUT|28|51|et devoret fructum iumentorum tuorum ac fruges terrae tuae, donec intereas, et non relinquat tibi triticum, vinum et oleum, partum armentorum et incrementum ovium, donec te disperdat
DEUT|28|52|et obsideat te in cunctis urbibus tuis, donec destruantur muri tui firmi atque sublimes, in quibus habebas fiduciam in omni terra tua. Obsideberis intra portas tuas in omni terra tua, quam dabit tibi Dominus Deus tuus,
DEUT|28|53|et comedes fructum uteri tui, carnes filiorum tuorum et filiarum tuarum, quas dederit tibi Dominus Deus tuus, in obsidione et angustia, qua opprimet te hostis tuus.
DEUT|28|54|Homo tener in te et delicatus valde invidebit fratri suo et uxori, quae cubat in sinu suo, et residuis filiis suis, quos reservaverit,
DEUT|28|55|ne det uni ex eis de carnibus filiorum suorum, quas comedet, eo quod nihil aliud habeat in obsidione et angustia, qua oppresserit te inimicus tuus intra omnes portas tuas.
DEUT|28|56|Tenera mulier in te et delicata, quae non tentabat pedis vestigium figere in terram propter mollitiem et teneritudinem nimiam, invidebit viro suo, qui cubat in sinu eius, filio et filiae
DEUT|28|57|et illuviei secundarum, quae egrediuntur de medio feminum eius, et liberis, qui eadem hora nati sunt; comedet enim eos clam propter rerum omnium penuriam in obsidione et angustia, qua opprimet te inimicus tuus intra portas tuas.
DEUT|28|58|Nisi custodieris et feceris omnia verba legis huius, quae scripta sunt in hoc volumine, et timueris nomen gloriosum et terribile hoc, Dominum Deum tuum,
DEUT|28|59|augebit ultra modum Dominus plagas tuas et plagas seminis tui, plagas magnas et perseverantes, infirmitates pessimas et perpetuas,
DEUT|28|60|et convertet in te omnes afflictiones Aegypti, quas timuisti, et adhaerebunt tibi.
DEUT|28|61|Insuper universos languores et plagas, quae non sunt scriptae in volumine legis huius, inducet Dominus super te, donec te conterat;
DEUT|28|62|et remanebitis pauci numero, qui prius eratis sicut astra caeli prae multitudine, quoniam non audisti vocem Domini Dei tui.
DEUT|28|63|Et sicut ante laetatus est Dominus super vos bene vobis faciens vosque multiplicans, sic laetabitur super vos disperdens vos atque subvertens, ut auferamini de terra, ad quam ingredieris possidendam.
DEUT|28|64|Disperget te Dominus in omnes populos a summitate terrae usque ad terminos eius, et servies ibi diis alienis, quos et tu ignorasti et patres tui, lignis et lapidibus.
DEUT|28|65|In gentibus quoque illis non quiesces, neque erit requies vestigio pedis tui; dabit enim tibi Dominus ibi cor pavidum et deficientes oculos et animam consumptam maerore.
DEUT|28|66|Et erit vita tua quasi pendens ante te; timebis nocte et die et non credes vitae tuae.
DEUT|28|67|Mane dices: "Quis mihi det vesperum?"; et vespere: "Quis mihi det mane?", propter cordis tui formidinem, qua terreberis, et propter ea, quae tuis videbis oculis.
DEUT|28|68|Reducet te Dominus classibus in Aegyptum per viam, de qua dixi tibi, ut eam amplius non videres; ibi vendetis vos inimicis vestris in servos et ancillas, et non erit qui emat ".
DEUT|28|69|Haec sunt verba foederis, quod praecepit Dominus Moysi, ut feriret cum filiis Israel in terra Moab, praeter illud foedus, quod cum eis pepigit in Horeb.
DEUT|29|1|Vocavitque Moyses omnem Israel et dixit ad eos: " Vos vidistis universa, quae fecit Dominus coram vobis in terra Aegypti pharaoni et omnibus servis eius universaeque terrae illius,
DEUT|29|2|tentationes magnas, quas viderunt oculi tui, signa illa portentaque ingentia;
DEUT|29|3|et non dedit Dominus vobis cor intellegens et oculos videntes et aures, quae possint audire, usque in praesentem diem.
DEUT|29|4|Adduxi vos quadraginta annis per desertum; non sunt attrita vestimenta vestra, nec calceamenta pedum tuorum vetustate consumpta sunt,
DEUT|29|5|panem non comedistis, vinum et siceram non bibistis, ut sciretis quia ego sum Dominus Deus vester.
DEUT|29|6|Et venistis ad hunc locum, egressusque est Sehon rex Hesebon et Og rex Basan occurrentes nobis ad pugnam, et percussimus eos.
DEUT|29|7|Et tulimus terram eorum ac tradidimus possidendam Ruben et Gad et dimidiae tribui Manasse.
DEUT|29|8|Custodite ergo verba pacti huius et implete ea, ut prosperemini in universis, quae facitis.
DEUT|29|9|Vos statis hodie cuncti coram Domino Deo vestro, principes vestri ac tribus et maiores natu atque praefecti, omnis vir Israel,
DEUT|29|10|liberi et uxores vestrae et advena tuus, qui tecum moratur in castris, a lignorum caesoribus usque ad hos, qui hauriunt aquas tuas,
DEUT|29|11|ut transeas in foedere Domini Dei tui et in iure iurando, quod hodie Dominus Deus tuus percutit tecum,
DEUT|29|12|ut suscitet te sibi hodie in populum, et ipse sit Deus tuus, sicut locutus est tibi et sicut iuravit patribus tuis, Abraham, Isaac et Iacob.
DEUT|29|13|Nec vobis solis ego hoc foedus ferio et haec iuramenta confirmo,
DEUT|29|14|sed cunctis hic nobiscum hodie praesentibus coram Domino Deo nostro et illis, qui hodie hic nobiscum non adsunt.
DEUT|29|15|Vos enim nostis quomodo habitaverimus in terra Aegypti et quomodo transierimus per medium nationum, quas transeuntes
DEUT|29|16|vidistis abominationes et idola eorum, lignum et lapidem, argentum et aurum, quae colebant.
DEUT|29|17|Ne forte sit inter vos vir aut mulier, familia aut tribus, cuius cor aversum est hodie a Domino Deo nostro, ut vadat et serviat diis illarum gentium, et sit inter vos radix germinans fel et absinthium;
DEUT|29|18|cumque audierit verba iuramenti huius, benedicat sibi in corde suo dicens: "Pax erit mihi, etsi ambulabo in pravitate cordis mei", et absumat terram irriguam et sitientem.
DEUT|29|19|Dominus non ignoscet ei, sed tunc quam maxime furor eius fumabit et zelus contra hominem illum, et sedebunt super eum omnia maledicta, quae scripta sunt in hoc volumine, et delebit Dominus nomen eius sub caelo
DEUT|29|20|et consumet eum in perditionem ex omnibus tribubus Israel, iuxta maledictiones foederis, quae in hoc libro legis scriptae sunt.
DEUT|29|21|Dicetque sequens generatio, filii vestri, qui nascentur deinceps, et peregrini, qui de longe venerint, videntes plagas terrae illius et infirmitates, quibus eam afflixerit Dominus,
DEUT|29|22|sulphur et salem: combusta est omnis humus eius, ita ut ultra non seratur, nec virens quippiam germinet in exemplum subversionis Sodomae et Gomorrae, Adamae et Seboim, quas subvertit Dominus in ira et furore suo.
DEUT|29|23|Et dicent omnes gentes: "Quare sic fecit Dominus terrae huic? Quae est haec ira furoris immensa?".
DEUT|29|24|Et respondebunt: "Quia dereliquerunt pactum Domini, Dei patrum suorum, quod pepigit cum eis, quando eduxit eos de terra Aegypti,
DEUT|29|25|et servierunt diis alienis et adoraverunt eos, quos nesciebant et quibus non fuerant attributi;
DEUT|29|26|idcirco iratus est furor Domini contra terram istam, ut induceret super eam omnia maledicta, quae in hoc volumine scripta sunt,
DEUT|29|27|et eiecit eos de terra eorum in ira et furore et indignatione maxima proiecitque in terram alienam, sicut hodie comprobatur".
DEUT|29|28|Abscondita Domino Deo nostro, manifesta autem nobis et filiis nostris usque in sempiternum, ut faciamus universa verba legis huius.
DEUT|30|1|Cum ergo venerint super te omnes sermones isti, benedic tio et maledictio, quas proposui in conspectu tuo, et ductus paenitudine cordis tui in universis gentibus, in quas disperserit te Dominus Deus tuus,
DEUT|30|2|et reversus fueris ad eum et oboedieris eius imperiis secundum omnia, quae ego hodie praecipio tibi, cum filiis tuis in toto corde tuo et in tota anima tua,
DEUT|30|3|reducet Dominus Deus tuus captivitatem tuam ac miserebitur tui et rursum congregabit te de cunctis populis, in quos te ante dispersit.
DEUT|30|4|Si ad cardines caeli fueris dissipatus, inde te retrahet Dominus Deus tuus et assumet
DEUT|30|5|atque introducet in terram, quam possederunt patres tui, et obtinebis eam; et feliciorem et maioris numeri esse te faciet quam fuerunt patres tui.
DEUT|30|6|Circumcidet Dominus Deus tuus cor tuum et cor seminis tui, ut diligas Dominum Deum tuum in toto corde tuo et in tota anima tua, ut possis vivere.
DEUT|30|7|Omnes autem maledictiones has convertet super inimicos tuos et eos, qui oderunt te et persequuntur.
DEUT|30|8|Tu autem reverteris et audies vocem Domini faciesque universa mandata, quae ego praecipio tibi hodie;
DEUT|30|9|et abundare te faciet Dominus Deus tuus in cunctis operibus manuum tuarum, in subole uteri tui et in fructu iumentorum tuorum et in ubertate terrae tuae, in rerum omnium largitate; revertetur enim Dominus, ut gaudeat super te in omnibus bonis, sicut gavisus est in patribus tuis.
DEUT|30|10|Si tamen audieris vocem Domini Dei tui et custodieris mandata eius et praecepta, quae in hac lege conscripta sunt, et revertaris ad Dominum Deum tuum in toto corde tuo et in tota anima tua.
DEUT|30|11|Mandatum hoc, quod ego praecipio tibi hodie, non supra te est neque procul positum
DEUT|30|12|nec in caelo situm, ut possis dicere: "Quis nobis ad caelum valet ascendere, ut deferat illud ad nos, et audiamus atque opere compleamus?".
DEUT|30|13|Neque trans mare positum, ut causeris et dicas: "Quis nobis transfretare poterit mare et illud ad nos usque deferre, ut possimus audire et facere quod praeceptum est?".
DEUT|30|14|Sed iuxta te est sermo valde in ore tuo et in corde tuo, ut facias illum.
DEUT|30|15|Considera quod hodie proposuerim in conspectu tuo vitam et bonum, et e contrario mortem et malum.
DEUT|30|16|Si oboedieris mandatis Domini Dei tui, quae ego praecipio tibi hodie, ut diligas Dominum Deum tuum et ambules in viis eius et custodias mandata illius et praecepta atque iudicia, vives; ac multiplicabit te benedicetque tibi in terra, ad quam ingredieris possidendam.
DEUT|30|17|Sin autem aversum fuerit cor tuum, et audire nolueris atque errore deceptus adoraveris deos alienos et servieris eis,
DEUT|30|18|praedico vobis hodie quod pereatis et parvo tempore moremini in terra, ad quam, Iordane transmisso, ingredieris possidendam.
DEUT|30|19|Testes invoco hodie contra vos caelum et terram quod proposuerim vobis vitam et mortem, benedictionem et maledictionem. Elige ergo vitam, ut et tu vivas et semen tuum
DEUT|30|20|et diligas Dominum Deum tuum atque oboedias voci eius et illi adhaereas ipse est enim vita tua et longitudo dierum tuorum - ut habites in terra, pro qua iuravit Dominus patribus tuis, Abraham, Isaac et Iacob, ut daret eam illis ".
DEUT|31|1|Abiit itaque Moyses et locu tus est omnia verba haec ad universum Israel
DEUT|31|2|et dixit ad eos: " Centum viginti annorum sum hodie, non possum ultra egredi et ingredi, praesertim cum et Dominus dixerit mihi: "Non transibis Iordanem istum".
DEUT|31|3|Dominus Deus tuus ipse transibit ante te; ipse delebit gentes has in conspectu tuo, et possidebis eas, et Iosue transibit ante te, sicut locutus est Dominus.
DEUT|31|4|Facietque Dominus eis, sicut fecit Sehon et Og regibus Amorraeorum et terrae eorum delevitque eos.
DEUT|31|5|Cum ergo et hos tradiderit vobis, similiter facietis eis, sicut praecepi vobis.
DEUT|31|6|Viriliter agite et confortamini; nolite timere nec paveatis a conspectu eorum, quia Dominus Deus tuus ipse est ductor tuus et non dimittet nec derelinquet te ".
DEUT|31|7|Vocavitque Moyses Iosue et dixit ei coram omni Israel: " Confortare et esto robustus; tu enim introduces populum istum in terram, quam daturum se patribus eorum iuravit Dominus, et tu eam sorte divides eis.
DEUT|31|8|Et Dominus, qui ductor tuus est, ipse erit tecum, non dimittet nec derelinquet te; noli timere nec paveas ".
DEUT|31|9|Et scripsit Moyses legem hanc et tradidit eam sacerdotibus filiis Levi, qui portabant arcam foederis Domini, et cunctis senioribus Israel;
DEUT|31|10|praecepitque eis dicens: " Post septem annos, anno remissionis, in sollemnitate Tabernaculorum,
DEUT|31|11|convenientibus cunctis ex Israel, ut appareant in conspectu Domini Dei tui in loco, quem elegerit, leges verba legis huius coram omni Israel, audientibus eis;
DEUT|31|12|congrega populum tam viros quam mulieres, parvulos et advenas, qui sunt intra portas tuas, ut audientes discant et timeant Dominum Deum vestrum et custodiant impleantque omnes sermones legis huius;
DEUT|31|13|filii quoque eorum, qui nunc ignorant, audiant et discant timere Dominum Deum vestrum cunctis diebus, quibus versamini in terra, ad quam vos, Iordane transmisso, pergitis obtinendam ".
DEUT|31|14|Et ait Dominus ad Moysen: " Ecce prope sunt dies mortis tuae; voca Iosue, et state in tabernaculo conventus, ut praecipiam ei ". Abierunt ergo Moyses et Iosue et steterunt in tabernaculo conventus;
DEUT|31|15|apparuitque Dominus ibi in columna nubis, quae stetit in introitu tabernaculi.
DEUT|31|16|Dixitque Dominus ad Moysen: " Ecce tu dormies cum patribus tuis, et populus iste consurgens fornicabitur post deos alienos terrae, ad quam ingredietur; ibi derelinquet me et irritum faciet foedus, quod pepigi cum eo.
DEUT|31|17|Et irascetur furor meus contra eum in die illo, et derelinquam eos et abscondam faciem meam ab eis, et erit in devorationem; invenient eum mala multa et afflictiones, ita ut dicat in illo die: "Vere, quia non est Deus mecum, invenerunt me haec mala".
DEUT|31|18|Ego autem abscondam et celabo faciem meam in die illo, propter omnia mala, quae fecit, quia secutus est deos alienos.
DEUT|31|19|Nunc itaque scribite vobis canticum istud, et doce filios Israel, ut memoriter teneant et ore decantent, ut sit mihi carmen istud pro testimonio inter filios Israel.
DEUT|31|20|Introducam enim eum in terram, pro qua iuravi patribus eius, lacte et melle manantem. Cumque comederit et saturatus crassusque fuerit, avertetur ad deos alienos, et servient eis detrahentque mihi et irritum facient pactum meum.
DEUT|31|21|Postquam invenerint eum mala multa et afflictiones, respondebit ei canticum istud pro testimonio, quod nulla delebit oblivio ex ore seminis sui; scio enim cogitationes eius, quae facit hodie, antequam introducam eum in terram, quam ei pollicitus sum ".
DEUT|31|22|Scripsit ergo Moyses canticum istud in die illo et docuit filios Israel.
DEUT|31|23|Praecepitque Dominus Iosue filio Nun et ait: " Confortare et esto robustus; tu enim introduces filios Israel in terram, quam eis pollicitus sum, et ego ero tecum ".
DEUT|31|24|Postquam ergo scripsit Moyses verba legis huius in volumine atque complevit,
DEUT|31|25|praecepit Levitis, qui portabant arcam foederis Domini, dicens:
DEUT|31|26|" Tollite librum legis istum et ponite eum in latere arcae foederis Domini Dei vestri, ut sit ibi contra te in testimonium.
DEUT|31|27|Ego enim scio contentionem tuam et cervicem tuam durissimam. Adhuc vivente me vobiscum, semper contentiose egistis contra Dominum; quanto magis cum mortuus fuero?
DEUT|31|28|Congregate ad me omnes maiores natu per tribus vestras atque praefectos vestros, et loquar audientibus eis sermones istos et invocabo contra eos caelum et terram.
DEUT|31|29|Novi enim quod post mortem meam inique agetis et declinabitis de via, quam praecepi vobis, et occurrent vobis mala in extremo tempore, quando feceritis malum in conspectu Domini, ut irritetis eum per opera manuum vestrarum ".
DEUT|31|30|Locutus est ergo Moyses, audiente universo coetu Israel, verba carminis huius et ad finem usque complevit:
DEUT|32|1|" Audite, caeli, quae loquor; audiat terra verba oris mei!
DEUT|32|2|Stillet ut pluvia doctrina mea, fluat ut ros eloquium meumquasi imber super herbamet quasi stillae super gramina.
DEUT|32|3|Quia nomen Domini invocabo:date magnificentiam Deo nostro!
DEUT|32|4|Petra, perfecta sunt opera eius,quia omnes viae eius iustitia.Deus fidelis et absque ulla iniquitate,iustus et rectus.
DEUT|32|5|Peccaverunt ei non filii eius in sordibus suis,generatio prava atque perversa.
DEUT|32|6|Haeccine redditis Domino,popule stulte et insipiens?Numquid non ipse est pater tuus, qui possedit te,ipse fecit et stabilivit te?
DEUT|32|7|Memento dierum antiquorum,cogita generationes singulas;interroga patrem tuum, et annuntiabit tibi,maiores tuos, et dicent tibi.
DEUT|32|8|Quando dividebat Altissimus gentes,quando separabat filios Adam,constituit terminos populorumiuxta numerum filiorum Israel;
DEUT|32|9|pars autem Domini populus eius,Iacob funiculus hereditatis eius.
DEUT|32|10|Invenit eum in terra deserta,in loco horroris et ululatu solitudinis;circumdedit eum et attenditet custodivit quasi pupillam oculi sui.
DEUT|32|11|Sicut aquila provocans ad volandum pullos suoset super eos volitans expandit alas suaset assumpsit eumatque portavit super pennas suas.
DEUT|32|12|Dominus solus dux eius fuit,et non erat cum eo deus alienus.
DEUT|32|13|Constituit eum super excelsam terram,ut comederet fructus agrorum,ut sugeret mel de petraoleumque de saxo durissimo,
DEUT|32|14|butyrum de armento et lac de ovibus,cum adipe agnorum et arietumfiliorum Basan et hircorum,cum medulla tritici,et sanguinem uvae biberet meracissimum.
DEUT|32|15|Incrassatus est dilectus et recalcitravit;incrassatus, impinguatus, dilatatus dereliquit Deum factorem suumet recessit a Petra salutari suo.
DEUT|32|16|Provocaverunt eum in diis alieniset in abominationibus ad iracundiam concitaverunt.
DEUT|32|17|Immolaverunt daemonibus et non Deo,diis, quos ignorabant;novi recentesque venerunt,quos non coluerunt patres vestri.
DEUT|32|18|Petram, quae te genuit, dereliquisti,et oblitus es Domini creatoris tui.
DEUT|32|19|Vidit Dominus et sprevit,quia provocaverunt eum filii sui et filiae.
DEUT|32|20|Et ait: "Abscondam faciem meam ab eiset considerabo novissima eorum;generatio enim perversa est,et infideles filii.
DEUT|32|21|Ipsi me provocaverunt in eo, qui non erat Deus,et irritaverunt in vanitatibus suis;et ego provocabo eos in eo, qui non est populus,et in gente stulta irritabo illos.
DEUT|32|22|Ignis succensus est in furore meoet ardebit usque ad inferni profundissima;devorabitque terram cum germine suoet montium fundamenta comburet.
DEUT|32|23|Congregabo super eos malaet sagittas meas complebo in eis.
DEUT|32|24|Consumentur fame et devorabuntur febriet peste amarissima;dentes bestiarum immittam in eos, cum veneno serpentium in pulvere.
DEUT|32|25|Foris vastabit eos gladius,et intus pavor:iuvenem simul ac virginem,lactantem cum homine sene.
DEUT|32|26|Dixi: Disperdam eos,cessare faciam ex hominibus memoriam eorum!,
DEUT|32|27|sed arrogantiam inimicorum timui,ne superbirent hostes eorumet dicerent: >Manus nostra excelsa, et non Dominus fecit haec omnia!'.
DEUT|32|28|Gens enim absque consilio estet sine prudentia.
DEUT|32|29|Utinam saperent et intellegerent haecac novissima sua providerent!
DEUT|32|30|Quomodo persequatur unus mille,et duo fugent decem milia?Nonne ideo, quia Petra eorum vendidit eos,et Dominus tradidit illos?".
DEUT|32|31|Non enim est petra eorum ut Petra nostra,et inimici nostri sunt iudices.
DEUT|32|32|Vere de vinea Sodomorum vinea eorumet de suburbanis Gomorrae;uva eorum uva felliset botri amarissimi;
DEUT|32|33|fel draconum vinum eorumet venenum aspidum insanabile.
DEUT|32|34|Nonne haec condita sunt apud meet signata in thesauris meis?
DEUT|32|35|Mea est ultio, et ego retribuam in tempore,in quo labetur pes eorum!Iuxta est dies perditionis,et adesse festinat sors eorum.
DEUT|32|36|Iudicabit Dominus populum suumet in servis suis miserebitur;videbit quod infirmata sit manus,et defecerint clausi ac liberati.
DEUT|32|37|Et dicet: "Ubi sunt dii eorum,petra, in qua habebant fiduciam,
DEUT|32|38|de quorum victimis comedebant adipeset bibebant vinum libaminum?Surgant et opitulentur vobiset in necessitate vos protegant!
DEUT|32|39|Videte nunc quod ego sim solus,et non sit Deus praeter me.Ego occidam et ego vivere faciam;percutiam et ego sanabo;et non est qui de manu mea possit eruere.
DEUT|32|40|Levabo ad caelum manum meamet dicam: Vivo ego in aeternum!
DEUT|32|41|Si acuero ut fulgur gladium meum,et arripuerit iudicium manus mea,reddam ultionem hostibus meiset his, qui oderunt me, retribuam.
DEUT|32|42|Inebriabo sagittas meas sanguine,et gladius meus devorabit carnes:de cruore occisorum et captivorum,de capite ducum inimici!".
DEUT|32|43|Laudate, gentes, populum eius,quia sanguinem servorum suorum ulcisceturet vindictam retribuet in hostes suoset propitius erit terrae populi sui ".
DEUT|32|44|Venit ergo Moyses et locutus est omnia verba cantici huius in auribus populi, ipse et Iosue filius Nun;
DEUT|32|45|complevitque omnes sermones istos loquens ad universum Israel.
DEUT|32|46|Et dixit ad eos: " Ponite corda vestra in omnia verba, quae ego testificor vobis hodie, ut mandetis ea filiis vestris custodire et facere et implere universa verba legis huius;
DEUT|32|47|quia verbum non incassum vobis, sed est vita vestra: et in verbo hoc longo perseverabitis tempore in terra, ad quam, Iordane transmisso, ingredimini possidendam ".
DEUT|32|48|Locutusque est Dominus ad Moysen in eadem die dicens:
DEUT|32|49|" Ascende in montem istum Abarim, in montem Nabo, qui est in terra Moab contra Iericho, et vide terram Chanaan, quam ego tradam filiis Israel obtinendam.
DEUT|32|50|Et morere in monte, quem conscendens iungeris populo tuo, sicut mortuus est Aaron frater tuus in monte Hor et appositus populo suo.
DEUT|32|51|Quia praevaricati estis contra me in medio filiorum Israel ad aquas Meribathcades deserti Sin, quia non sanctificastis me inter filios Israel.
DEUT|32|52|E contra videbis terram et non ingredieris in eam, quam ego dabo filiis Israel ".
DEUT|33|1|Haec est benedictio, qua be nedixit Moyses homo Dei fi liis Israel ante mortem suam.
DEUT|33|2|Et ait: Dominus de Sinai venitet de Seir ortus est eis;apparuit de monte Pharanet venit in Meribathcadesde meridie eius in Asedoth.
DEUT|33|3|Vere diligit populos;omnes sancti eius in manu illius sunt;et, qui appropinquant pedibus tuis,accipient de doctrina tua.
DEUT|33|4|Legem praecepit nobis Moyses,hereditatem multitudinis Iacob.
DEUT|33|5|Et factus est apud dilectum rex,congregatis principibus populicum tribubus Israel ".
DEUT|33|6|" Vivat Ruben et non moriaturet sit parvus in numero ".
DEUT|33|7|Haec est Iudae benedictio: Audi, Domine, vocem Iudaeet ad populum suum introduc eum.Manus eius pugnabunt pro eo,et adiutor illius contra adversarios eius eris ".
DEUT|33|8|De Levi quoque ait: Tummim et Urim tuiviro sancto tuo,quem probasti in Massaet cum quo litigasti ad aquas Meriba.
DEUT|33|9|Qui dixit de patre suo et matre sua:Nescio vos";et fratres suos ignoravitet filios suos nescivit.Quia custodierunt eloquium tuumet pactum tuum servaverunt.
DEUT|33|10|Docebunt iudicia tua Iacobet legem tuam Israel;ponent thymiama in naribus tuiset holocaustum super altare tuum.
DEUT|33|11|Benedic, Domine, fortitudini eiuset opera manuum illius suscipe.Percute lumbos inimicorum eius;et, qui oderunt eum, non consurgant ".
DEUT|33|12|De Beniamin ait: Amantissimus Dominihabitabit confidenter in eo;Altissimus proteget eum tota dieet inter umeros illius requiescet ".
DEUT|33|13|De Ioseph quoque ait: Benedicta a Domino terra eius:donis caeli, roreatque abysso subiacente,
DEUT|33|14|fructibus soliset donis mensium,
DEUT|33|15|primitiis antiquorum montiumet donis collium aeternorum,
DEUT|33|16|frugibus terrae et plenitudine eius.Benedictio illius, qui apparuit in rubo,veniat super caput Iosephet super verticem nazaraei inter fratres suos;
DEUT|33|17|quasi primogeniti tauri pulchritudo eius,cornua unicornis cornua illius,in ipsis ventilabit gentesusque ad terminos terrae.Hae sunt multitudines Ephraim,et hae milia Manasse ".
DEUT|33|18|De Zabulon ait: Laetare, Zabulon, in exitu tuo,et Issachar, in tabernaculis tuis!
DEUT|33|19|Populos ad montem vocabunt,ibi immolabunt victimas iustitiae.Qui inundationem maris, quasi lac, sugentet thesauros absconditos arenarum ".
DEUT|33|20|De Gad ait: Benedictus, qui dilatat Gad!Quasi leo requiescitdilaceratque brachium et verticem.
DEUT|33|21|Et vidit primitias sibi,quia ibi pars ducis erat reposita;qui fuit cum principibus populiet fecit iustitiam Dominiet iudicia sua cum Israel ".
DEUT|33|22|De Dan quoque ait: Dan catulus leonisprosiliet largiter de Basan ".
DEUT|33|23|De Nephthali dixit: Nephthali satiabatur beneplacitoet plenus erit benedictione Domini:mare et meridiem possidebit ".
DEUT|33|24|De Aser quoque ait: Benedictus prae filiis Aser!Sit placens fratribus suiset tingat in oleo pedem suum.
DEUT|33|25|Ferrum et aes serae tuae,sicut dies tui robur tuum ".
DEUT|33|26|" Non est ut Deus Iesurun,qui ascendit super caelos ad auxilium tuumet in magnificentia sua super nubes.
DEUT|33|27|Habitaculum Deus antiquus,et subter brachia sempiterna.Eiciet a facie tua inimicumdicetque: "Conterere!".
DEUT|33|28|Habitabit Israel confidenter,et fons Iacob solus;stillabunt in terra frumenti et vini,caelique rorem.
DEUT|33|29|Beatus tu, Israel! Quis similis tui,popule, qui salvaris in Domino?Ipse est scutum auxilii tuiet gladius gloriae tuae.Blandientur tibi inimici tui,et tu eorum altitudines calcabis ".
DEUT|34|1|Ascendit ergo Moyses de campestribus Moab super montem Nabo in verticem Phasga contra Iericho; ostenditque ei Dominus omnem terram Galaad usque Dan
DEUT|34|2|et universum Nephthali terramque Ephraim et Manasse et omnem terram Iudae usque ad mare occidentale
DEUT|34|3|et Nageb et latitudinem campi Iericho civitatis palmarum usque Segor.
DEUT|34|4|Dixitque Dominus ad eum: " Haec est terra, pro qua iuravi Abraham, Isaac et Iacob, dicens: Semini tuo dabo eam. Vidisti eam oculis tuis et non transibis ad illam ".
DEUT|34|5|Mortuusque est ibi Moyses servus Domini in terra Moab, iubente Domino.
DEUT|34|6|Et sepelivit eum in valle in terra Moab contra Bethphegor; et non cognovit homo sepulcrum eius usque in praesentem diem.
DEUT|34|7|Moyses centum et viginti annorum erat, quando mortuus est; non caligavit oculus eius, nec robur illius defecit.
DEUT|34|8|Fleveruntque eum filii Israel in campestribus Moab triginta diebus; et completi sunt dies planctus lugentium Moysen.
DEUT|34|9|Iosue vero filius Nun repletus est spiritu sapientiae, quia Moyses posuit super eum manus suas; et oboedierunt ei filii Israel feceruntque, sicut praecepit Dominus Moysi.
DEUT|34|10|Et non surrexit ultra propheta in Israel sicut Moyses, quem nosset Dominus facie ad faciem,
DEUT|34|11|in omnibus signis atque portentis, quae misit per eum, ut faceret in terra Aegypti pharaoni et omnibus servis eius universaeque terrae illius,
DEUT|34|12|et in cuncta manu robusta magnisque mirabilibus, quae fecit Moyses coram universo Israel.
