SONG|1|1|Canticum Canticorum Salomonis.
SONG|1|2|Osculetur me osculo oris sui!Nam meliores sunt amores tui vino:
SONG|1|3|in fragrantiam unguentorum tuorum optimorum.Oleum effusum nomen tuum;ideo adulescentulae dilexerunt te.
SONG|1|4|Trahe me post te. Curramus!Introducat me rex in cellaria sua;exsultemus et laetemur in tememores amorum tuorum super vinum;recte diligunt te.
SONG|1|5|Nigra sum sed formosa,filiae Ierusalem,sicut tabernacula Cedar,sicut pelles Salma.
SONG|1|6|Nolite me considerare quod fusca sim,quia decoloravit me sol.Filii matris meae irati sunt mihi;posuerunt me custodem in vineis,vineam meam non custodivi.
SONG|1|7|Indica mihi, tu, quem diligit anima mea,ubi pascas,ubi cubes in meridie,ne vagari incipiampost greges sodalium tuorum.
SONG|1|8|Si ignoras,o pulcherrima inter mulieres,egredere et abi post vestigia gregumet pasce haedos tuosiuxta tabernacula pastorum.
SONG|1|9|Equae in curribus pharaonisassimilavi te, amica mea.
SONG|1|10|Pulchrae sunt genae tuae inter inaures,collum tuum inter monilia.
SONG|1|11|Inaures aureas faciemus tibivermiculatas argento.
SONG|1|12|Dum esset rex in accubitu suo,nardus mea dedit odorem suum.
SONG|1|13|Fasciculus myrrhae dilectus meus mihi,qui inter ubera mea commoratur.
SONG|1|14|Botrus cypri dilectus meus mihiin vineis Engaddi.
SONG|1|15|Ecce tu pulchra es, amica mea,ecce tu pulchra es:oculi tui columbarum.
SONG|1|16|Ecce tu pulcher es, dilecte mi,et decorus.Lectulus noster floridus,
SONG|1|17|tigna domorum nostrarum cedrina,laquearia nostra cupressina.
SONG|2|1|Ego flos campiet lilium convallium.
SONG|2|2|Sicut lilium inter spinas,sic amica mea inter filias.
SONG|2|3|Sicut malus inter ligna silvarum,sic dilectus meus inter filios.Sub umbra illius, quem desideraveram, sedi,et fructus eius dulcis gutturi meo.
SONG|2|4|Introduxit me in cellam vinariam,et vexillum eius super me est caritas.
SONG|2|5|Fulcite me uvarum placentis,stipate me malis,quia amore langueo.
SONG|2|6|Laeva eius sub capite meo,et dextera illius amplexatur me.
SONG|2|7|Adiuro vos, filiae Ierusalem,per capreas cervasque camporum,ne suscitetis neque evigilare faciatis dilectam,quoadusque ipsa velit.
SONG|2|8|Vox dilecti mei!Ecce iste venitsaliens in montibus,transiliens colles.
SONG|2|9|Similis est dilectus meus capreaehinnuloque cervorum.En ipse statpost parietem nostrumrespiciens per fenestras,prospiciens per cancellos.
SONG|2|10|En dilectus meus loquitur mihi: Surge, amica mea,columba mea, formosa mea, et veni.
SONG|2|11|Iam enim hiems transiit,imber abiit et recessit.
SONG|2|12|Flores apparuerunt in terra,tempus putationis advenit;vox turturis audita estin terra nostra,
SONG|2|13|ficus protulit grossos suos,vineae florentes dederunt odorem suum;surge, amica mea,speciosa mea, et veni,
SONG|2|14|columba mea, in foraminibus petrae,in caverna abrupta.Ostende mihi faciem tuam,sonet vox tua in auribus meis;vox enim tua dulcis,et facies tua decora ".
SONG|2|15|Capite nobis vulpes, vulpes parvulas,quae demoliuntur vineas,nam vineae nostrae florescunt.
SONG|2|16|Dilectus meus mihi, et ego illi,qui pascitur inter lilia,
SONG|2|17|antequam aspiret dies,et festinent umbrae.Revertere; similis esto,dilecte mi, capreaehinnuloque cervorum super montes Bether.
SONG|3|1|In lectulo meo per noctesquaesivi, quem diligit anima mea;quaesivi illum et non inveni.
SONG|3|2|" Surgam et circuibo civitatem;per vicos et plateasquaeram, quem diligit anima mea".Quaesivi illum et non inveni.
SONG|3|3|Invenerunt me vigiles,qui circumeunt civitatem: Num, quem diligit anima mea, vidistis? ".
SONG|3|4|Paululum cum pertransissem eos,inveni, quem diligit anima mea;tenui eum nec dimittam,donec introducam illum in domum matris meaeet in cubiculum genetricis meae.
SONG|3|5|Adiuro vos, filiae Ierusalem,per capreas cervasque camporum,ne suscitetis neque evigilare faciatis dilectam,donec ipsa velit.
SONG|3|6|Quid hoc, quod ascendit per desertumsicut virgula fumi,aromatizans tus et myrrhamet universum pulverem pigmentarii?
SONG|3|7|En lectulum Salomonis.Sexaginta fortes ambiunt illumex fortissimis Israel,
SONG|3|8|omnes tenentes gladioset ad bella doctissimi,uniuscuiusque ensis super femur suumpropter timores nocturnos.
SONG|3|9|Ferculum fecit sibi rex Salomonde lignis Libani;
SONG|3|10|columnas eius fecit argenteas,reclinatorium aureum,sedile purpureum:medium eius stratum ebeneum.Filiae Ierusalem,
SONG|3|11|egredimini et videte,filiae Sion,regem Salomonemin diademate, quo coronavit illum mater suain die desponsationis illiuset in die laetitiae cordis eius.
SONG|4|1|Quam pulchra es, amica mea,quam pulchra es:oculi tui columbarumper velamen tuum.Capilli tui sicut grex caprarum,quae descenderunt de monte Galaad;
SONG|4|2|dentes tui sicut grex tonsarum,quae ascenderunt de lavacro:omnes gemellis fetibus,et sterilis non est inter eas.
SONG|4|3|Sicut vitta coccinea labia tua,et eloquium tuum dulce;sicut fragmen mali punici, ita genae tuaeper velamen tuum.
SONG|4|4|Sicut turris David collum tuum,quae aedificata est cum propugnaculis:mille clipei pendent ex ea,omnis armatura fortium.
SONG|4|5|Duo ubera tua sicut duo hinnuli,capreae gemelli,qui pascuntur in liliis.
SONG|4|6|Antequam aspiret dies,et festinent umbrae,vadam ad montem myrrhaeet ad collem turis.
SONG|4|7|Tota pulchra es, amica mea,et macula non est in te.
SONG|4|8|Veni de Libano, sponsa,veni de Libano,ingredere;respice de capite Amana,de vertice Sanir et Hermon,de cubilibus leonum,de montibus pardorum.
SONG|4|9|Vulnerasti cor meum, soror mea, sponsa,vulnerasti cor meum in uno oculorum tuorumet in uno monili torquis tui.
SONG|4|10|Quam pulchri sunt amores tui, soror, mea sponsa;meliores sunt amores tui vino,et odor unguentorum tuorum super omnia aromata.
SONG|4|11|Favus distillans labia tua, sponsa;mel et lac sub lingua tua,et odor vestimentorum tuorumsicut odor Libani.
SONG|4|12|Hortus conclusus, soror mea, sponsa,hortus conclusus, fons signatus;
SONG|4|13|propagines tuae paradisus malorum punicorumcum optimis fructibus,cypri cum nardo.
SONG|4|14|Nardus et crocus,fistula et cinnamomumcum universis lignis turiferis,myrrha et aloecum omnibus primis unguentis.
SONG|4|15|Fons hortorum,puteus aquarum viventium,quae fluunt impetu de Libano.
SONG|4|16|Surge, aquilo,et veni, auster;perfla hortum meum,et fluant aromata illius.
SONG|5|1|Veniat dilectus meus in hortum suumet comedat fructus eius optimos.Veni in hortum meum, soror mea, sponsa;messui myrrham meam cum aromatibus meis,comedi favum cum melle,bibi vinum cum lacte meo.Comedite, amici, et bibiteet inebriamini, carissimi.
SONG|5|2|Ego dormio, et cor meum vigilat.Vox dilecti mei pulsantis: Aperi mihi, soror mea, amica mea,columba mea, immaculata mea,quia caput meum plenum est rore, et cincinni mei guttis noctium ".
SONG|5|3|" Exspoliavi me tunica mea,quomodo induar illa?Lavi pedes meos,quomodo inquinabo illos?".
SONG|5|4|Dilectus meus misit manum suam per foramen,et venter meus ilico intremuit.
SONG|5|5|Surrexi, ut aperirem dilecto meo;manus meae stillaverunt myrrham,et digiti mei pleni myrrha probatissimasuper ansam pessuli.
SONG|5|6|Aperui dilecto meo;at ille declinaverat atque transierat.Anima mea liquefacta est, quia discesserat.Quaesivi et non inveni illum;vocavi, et non respondit mihi.
SONG|5|7|Invenerunt me custodes,qui circumeunt civitatem;percusserunt me et vulneraverunt me,tulerunt pallium meum mihicustodes murorum.
SONG|5|8|Adiuro vos, filiae Ierusalem:si inveneritis dilectum meum,quid nuntietis ei? Quia amore langueo ".
SONG|5|9|Quid est dilecto tuo prae ceteris,o pulcherrima mulierum?Quid est dilecto tuo prae ceteris,quia sic adiurasti nos?
SONG|5|10|Dilectus meus candidus et rubicundusdignoscitur ex milibus.
SONG|5|11|Caput eius aurum optimum,cincinni eius sicut racemi palmarum,nigri quasi corvus.
SONG|5|12|Oculi eius sicut columbaesuper rivulos aquarum,quae lacte sunt lotaeet resident iuxta fluenta plenissima.
SONG|5|13|Genae illius sicut areolae aromatum,turriculae unguentorum;labia eius liliadistillantia myrrham primam.
SONG|5|14|Manus illius tornatiles aureae,plenae hyacinthis;venter eius opus eburneumdistinctum sapphiris.
SONG|5|15|Crura illius columnae marmoreae,quae fundatae sunt super bases aureas;species eius ut Libani,electus ut cedri.
SONG|5|16|Guttur illius suavissimum,et totus desiderabilis.Talis est dilectus meus, et ipse est amicus meus,filiae Ierusalem.
SONG|6|1|Quo abiit dilectus tuus,o pulcherrima mulierum?Quo declinavit dilectus tuus,et quaeremus eum tecum?
SONG|6|2|Dilectus meus descendit in hortum suumad areolam aromatum,ut pascatur in hortiset lilia colligat.
SONG|6|3|Ego dilecto meo, et dilectus meus mihi,qui pascitur inter lilia.
SONG|6|4|Pulchra es, amica mea, sicut Thersa,decora sicut Ierusalem,terribilis ut castrorum acies ordinata.
SONG|6|5|Averte oculos tuos a me,quia ipsi me conturbant.Capilli tui sicut grex caprarum,quae descenderunt de Galaad.
SONG|6|6|Dentes tui sicut grex ovium,quae ascenderunt de lavacro:omnes gemellis fetibus,et sterilis non est in eis.
SONG|6|7|Sicut fragmen mali punici, sic genae tuaeper velamen tuum.
SONG|6|8|Sexaginta sunt reginae,et octoginta concubinae,et adulescentularum non est numerus;
SONG|6|9|una est columba mea, perfecta mea,una est matri suae,electa genetrici suae.Viderunt eam filiae et beatissimam praedicaverunt;reginae et concubinae, et laudaverunt eam:
SONG|6|10|" Quae est ista, quae progreditur quasi aurora consurgens,pulchra ut luna,electa ut sol,terribilis ut castrorum acies ordinata? ".
SONG|6|11|Descendi in hortum nucum,ut viderem poma convalliumet inspicerem, si floruisset vinea,et germinassent mala punica.
SONG|6|12|Non advertit animus meus,cum posuit me in quadrigas principis populi mei.
SONG|7|1|Convertere, convertere, Sula mitis;convertere, convertere, ut intueamur te.Quid aspicitis in Sulamitem,cum saltat inter binos choros?
SONG|7|2|Quam pulchri sunt pedes tui in calceamentis,filia principis!Flexurae femorum tuorum sicut monilia,quae fabricata sunt manu artificis.
SONG|7|3|Gremium tuum crater tornatilis:numquam indigeat vino mixto;venter tuus sicut acervus triticivallatus liliis.
SONG|7|4|Duo ubera tua sicut duo hinnuli,gemelli capreae,
SONG|7|5|collum tuum sicut turris eburnea.Oculi tui sicut piscinae in Hesebon,quae sunt ad portam Bathrabbim;nasus tuus sicut turris Libani,quae respicit contra Damascum.
SONG|7|6|Caput tuum ut Carmelus,et comae capitis tui sicut purpura;rex vincitur cincinnis.
SONG|7|7|Quam pulchra es et quam decora,carissima, in deliciis!
SONG|7|8|Statura tua assimilata est palmae,et ubera tua botris.
SONG|7|9|Dixi: " Ascendam in palmamet apprehendam fructus eius ".Et erunt ubera tua sicut botri vineae,et odor oris tui sicut malorum.
SONG|7|10|Guttur tuum sicut vinum optimum,dignum dilecto meo ad potandum,labiisque et dentibus illius ad ruminandum.
SONG|7|11|Ego dilecto meo,et ad me appetitus eius.
SONG|7|12|Veni, dilecte mi, egrediamur in agrum,commoremur in villis;
SONG|7|13|mane properabimus ad vineas,videbimus; si floruit vinea,si flores aperiuntur,si floruerunt mala punica;ibi dabo tibi amores meos.
SONG|7|14|Mandragorae dederunt odorem;in portis nostris omnia poma optima,nova et vetera,dilecte mi, servavi tibi.
SONG|8|1|Quis mihi det te fratrem meum,sugentem ubera matris meae,ut inveniam te foris et deosculer te,et iam me nemo despiciat?
SONG|8|2|Apprehenderem te et ducerem in domum matris meae;ibi me doceres,et darem tibi poculum ex vino conditoet mustum malorum granatorum meorum.
SONG|8|3|Laeva eius sub capite meo,et dextera illius amplexatur me.
SONG|8|4|Adiuro vos, filiae Ierusalem,ne suscitetis neque evigilare faciatis dilectam,donec ipsa velit.
SONG|8|5|Quae est ista, quae ascendit de desertoinnixa super dilectum suum?Sub arbore malo suscitavi te;ibi parturivit te mater tua,ibi parturivit te genetrix tua.
SONG|8|6|Pone me ut signaculum super cor tuum,ut signaculum super brachium tuum,quia fortis est ut mors dilectio,dura sicut infernus aemulatio;lampades eius lampades ignisatque flammae divinae.
SONG|8|7|Aquae multae non potuerunt exstinguere caritatem,nec flumina obruent illam;si dederit homo omnem substantiam domus suae pro dilectione,quasi nihil despicient eum.
SONG|8|8|Soror nostra parvaet ubera non habet;quid faciemus sorori nostraein die, quando alloquenda est?
SONG|8|9|Si murus est,aedificemus super eum propugnacula argentea;si ostium est,compingamus illud tabulis cedrinis.
SONG|8|10|Ego murus,et ubera mea sicut turris;ex quo facta sum coram eoquasi pacem reperiens.
SONG|8|11|Vinea fuit Salomoniin Baalhamon.Tradidit eam custodibus;vir affert pro fructu eiusmille argenteos.
SONG|8|12|Vinea mea coram me est;mille tibi, Salomon,et ducenti his, qui custodiunt fructus eius.
SONG|8|13|Quae habitas in hortis,amici auscultant,fac me audire vocem tuam.
SONG|8|14|Fuge, dilecte mi,et assimilare capreaehinnuloque cervorumsuper montes aromatum.
