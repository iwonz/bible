HAG|1|1|In the second year of Darius the king, in the sixth month, in the first day of the month, came the word of the LORD by Haggai the prophet unto Zerubbabel the son of Shealtiel, governor of Judah, and to Joshua the son of Josedech, the high priest, saying,
HAG|1|2|Thus speaketh the LORD of hosts, saying, This people say, The time is not come, the time that the LORD's house should be built.
HAG|1|3|Then came the word of the LORD by Haggai the prophet, saying,
HAG|1|4|Is it time for you, O ye, to dwell in your cieled houses, and this house lie waste?
HAG|1|5|Now therefore thus saith the LORD of hosts; Consider your ways.
HAG|1|6|Ye have sown much, and bring in little; ye eat, but ye have not enough; ye drink, but ye are not filled with drink; ye clothe you, but there is none warm; and he that earneth wages earneth wages to put it into a bag with holes.
HAG|1|7|Thus saith the LORD of hosts; Consider your ways.
HAG|1|8|Go up to the mountain, and bring wood, and build the house; and I will take pleasure in it, and I will be glorified, saith the LORD.
HAG|1|9|Ye looked for much, and, lo it came to little; and when ye brought it home, I did blow upon it. Why? saith the LORD of hosts. Because of mine house that is waste, and ye run every man unto his own house.
HAG|1|10|Therefore the heaven over you is stayed from dew, and the earth is stayed from her fruit.
HAG|1|11|And I called for a drought upon the land, and upon the mountains, and upon the corn, and upon the new wine, and upon the oil, and upon that which the ground bringeth forth, and upon men, and upon cattle, and upon all the labour of the hands.
HAG|1|12|Then Zerubbabel the son of Shealtiel, and Joshua the son of Josedech, the high priest, with all the remnant of the people, obeyed the voice of the LORD their God, and the words of Haggai the prophet, as the LORD their God had sent him, and the people did fear before the LORD.
HAG|1|13|Then spake Haggai the LORD's messenger in the LORD's message unto the people, saying, I am with you, saith the LORD.
HAG|1|14|And the LORD stirred up the spirit of Zerubbabel the son of Shealtiel, governor of Judah, and the spirit of Joshua the son of Josedech, the high priest, and the spirit of all the remnant of the people; and they came and did work in the house of the LORD of hosts, their God,
HAG|1|15|In the four and twentieth day of the sixth month, in the second year of Darius the king.
HAG|2|1|In the seventh month, in the one and twentieth day of the month, came the word of the LORD by the prophet Haggai, saying,
HAG|2|2|Speak now to Zerubbabel the son of Shealtiel, governor of Judah, and to Joshua the son of Josedech, the high priest, and to the residue of the people, saying,
HAG|2|3|Who is left among you that saw this house in her first glory? and how do ye see it now? is it not in your eyes in comparison of it as nothing?
HAG|2|4|Yet now be strong, O Zerubbabel, saith the LORD; and be strong, O Joshua, son of Josedech, the high priest; and be strong, all ye people of the land, saith the LORD, and work: for I am with you, saith the LORD of hosts:
HAG|2|5|According to the word that I covenanted with you when ye came out of Egypt, so my spirit remaineth among you: fear ye not.
HAG|2|6|For thus saith the LORD of hosts; Yet once, it is a little while, and I will shake the heavens, and the earth, and the sea, and the dry land;
HAG|2|7|And I will shake all nations, and the desire of all nations shall come: and I will fill this house with glory, saith the LORD of hosts.
HAG|2|8|The silver is mine, and the gold is mine, saith the LORD of hosts.
HAG|2|9|The glory of this latter house shall be greater than of the former, saith the LORD of hosts: and in this place will I give peace, saith the LORD of hosts.
HAG|2|10|In the four and twentieth day of the ninth month, in the second year of Darius, came the word of the LORD by Haggai the prophet, saying,
HAG|2|11|Thus saith the LORD of hosts; Ask now the priests concerning the law, saying,
HAG|2|12|If one bear holy flesh in the skirt of his garment, and with his skirt do touch bread, or pottage, or wine, or oil, or any meat, shall it be holy? And the priests answered and said, No.
HAG|2|13|Then said Haggai, If one that is unclean by a dead body touch any of these, shall it be unclean? And the priests answered and said, It shall be unclean.
HAG|2|14|Then answered Haggai, and said, So is this people, and so is this nation before me, saith the LORD; and so is every work of their hands; and that which they offer there is unclean.
HAG|2|15|And now, I pray you, consider from this day and upward, from before a stone was laid upon a stone in the temple of the LORD:
HAG|2|16|Since those days were, when one came to an heap of twenty measures, there were but ten: when one came to the pressfat for to draw out fifty vessels out of the press, there were but twenty.
HAG|2|17|I smote you with blasting and with mildew and with hail in all the labours of your hands; yet ye turned not to me, saith the LORD.
HAG|2|18|Consider now from this day and upward, from the four and twentieth day of the ninth month, even from the day that the foundation of the LORD's temple was laid, consider it.
HAG|2|19|Is the seed yet in the barn? yea, as yet the vine, and the fig tree, and the pomegranate, and the olive tree, hath not brought forth: from this day will I bless you.
HAG|2|20|And again the word of the LORD came unto Haggai in the four and twentieth day of the month, saying,
HAG|2|21|Speak to Zerubbabel, governor of Judah, saying, I will shake the heavens and the earth;
HAG|2|22|And I will overthrow the throne of kingdoms, and I will destroy the strength of the kingdoms of the heathen; and I will overthrow the chariots, and those that ride in them; and the horses and their riders shall come down, every one by the sword of his brother.
HAG|2|23|In that day, saith the LORD of hosts, will I take thee, O Zerubbabel, my servant, the son of Shealtiel, saith the LORD, and will make thee as a signet: for I have chosen thee, saith the LORD of hosts.
