1JOHN|1|1|That which was from the beginning, which we have heard, which we have seen with our eyes, which we have looked upon, and our hands have handled, of the Word of life;
1JOHN|1|2|(For the life was manifested, and we have seen it, and bear witness, and shew unto you that eternal life, which was with the Father, and was manifested unto us;)
1JOHN|1|3|That which we have seen and heard declare we unto you, that ye also may have fellowship with us: and truly our fellowship is with the Father, and with his Son Jesus Christ.
1JOHN|1|4|And these things write we unto you, that your joy may be full.
1JOHN|1|5|This then is the message which we have heard of him, and declare unto you, that God is light, and in him is no darkness at all.
1JOHN|1|6|If we say that we have fellowship with him, and walk in darkness, we lie, and do not the truth:
1JOHN|1|7|But if we walk in the light, as he is in the light, we have fellowship one with another, and the blood of Jesus Christ his Son cleanseth us from all sin.
1JOHN|1|8|If we say that we have no sin, we deceive ourselves, and the truth is not in us.
1JOHN|1|9|If we confess our sins, he is faithful and just to forgive us our sins, and to cleanse us from all unrighteousness.
1JOHN|1|10|If we say that we have not sinned, we make him a liar, and his word is not in us.
1JOHN|2|1|My little children, these things write I unto you, that ye sin not. And if any man sin, we have an advocate with the Father, Jesus Christ the righteous:
1JOHN|2|2|And he is the propitiation for our sins: and not for our's only, but also for the sins of the whole world.
1JOHN|2|3|And hereby we do know that we know him, if we keep his commandments.
1JOHN|2|4|He that saith, I know him, and keepeth not his commandments, is a liar, and the truth is not in him.
1JOHN|2|5|But whoso keepeth his word, in him verily is the love of God perfected: hereby know we that we are in him.
1JOHN|2|6|He that saith he abideth in him ought himself also so to walk, even as he walked.
1JOHN|2|7|Brethren, I write no new commandment unto you, but an old commandment which ye had from the beginning. The old commandment is the word which ye have heard from the beginning.
1JOHN|2|8|Again, a new commandment I write unto you, which thing is true in him and in you: because the darkness is past, and the true light now shineth.
1JOHN|2|9|He that saith he is in the light, and hateth his brother, is in darkness even until now.
1JOHN|2|10|He that loveth his brother abideth in the light, and there is none occasion of stumbling in him.
1JOHN|2|11|But he that hateth his brother is in darkness, and walketh in darkness, and knoweth not whither he goeth, because that darkness hath blinded his eyes.
1JOHN|2|12|I write unto you, little children, because your sins are forgiven you for his name's sake.
1JOHN|2|13|I write unto you, fathers, because ye have known him that is from the beginning. I write unto you, young men, because ye have overcome the wicked one. I write unto you, little children, because ye have known the Father.
1JOHN|2|14|I have written unto you, fathers, because ye have known him that is from the beginning. I have written unto you, young men, because ye are strong, and the word of God abideth in you, and ye have overcome the wicked one.
1JOHN|2|15|Love not the world, neither the things that are in the world. If any man love the world, the love of the Father is not in him.
1JOHN|2|16|For all that is in the world, the lust of the flesh, and the lust of the eyes, and the pride of life, is not of the Father, but is of the world.
1JOHN|2|17|And the world passeth away, and the lust thereof: but he that doeth the will of God abideth for ever.
1JOHN|2|18|Little children, it is the last time: and as ye have heard that antichrist shall come, even now are there many antichrists; whereby we know that it is the last time.
1JOHN|2|19|They went out from us, but they were not of us; for if they had been of us, they would no doubt have continued with us: but they went out, that they might be made manifest that they were not all of us.
1JOHN|2|20|But ye have an unction from the Holy One, and ye know all things.
1JOHN|2|21|I have not written unto you because ye know not the truth, but because ye know it, and that no lie is of the truth.
1JOHN|2|22|Who is a liar but he that denieth that Jesus is the Christ? He is antichrist, that denieth the Father and the Son.
1JOHN|2|23|Whosoever denieth the Son, the same hath not the Father: he that acknowledgeth the Son hath the Father also.
1JOHN|2|24|Let that therefore abide in you, which ye have heard from the beginning. If that which ye have heard from the beginning shall remain in you, ye also shall continue in the Son, and in the Father.
1JOHN|2|25|And this is the promise that he hath promised us, even eternal life.
1JOHN|2|26|These things have I written unto you concerning them that seduce you.
1JOHN|2|27|But the anointing which ye have received of him abideth in you, and ye need not that any man teach you: but as the same anointing teacheth you of all things, and is truth, and is no lie, and even as it hath taught you, ye shall abide in him.
1JOHN|2|28|And now, little children, abide in him; that, when he shall appear, we may have confidence, and not be ashamed before him at his coming.
1JOHN|2|29|If ye know that he is righteous, ye know that every one that doeth righteousness is born of him.
1JOHN|3|1|Behold, what manner of love the Father hath bestowed upon us, that we should be called the sons of God: therefore the world knoweth us not, because it knew him not.
1JOHN|3|2|Beloved, now are we the sons of God, and it doth not yet appear what we shall be: but we know that, when he shall appear, we shall be like him; for we shall see him as he is.
1JOHN|3|3|And every man that hath this hope in him purifieth himself, even as he is pure.
1JOHN|3|4|Whosoever committeth sin transgresseth also the law: for sin is the transgression of the law.
1JOHN|3|5|And ye know that he was manifested to take away our sins; and in him is no sin.
1JOHN|3|6|Whosoever abideth in him sinneth not: whosoever sinneth hath not seen him, neither known him.
1JOHN|3|7|Little children, let no man deceive you: he that doeth righteousness is righteous, even as he is righteous.
1JOHN|3|8|He that committeth sin is of the devil; for the devil sinneth from the beginning. For this purpose the Son of God was manifested, that he might destroy the works of the devil.
1JOHN|3|9|Whosoever is born of God doth not commit sin; for his seed remaineth in him: and he cannot sin, because he is born of God.
1JOHN|3|10|In this the children of God are manifest, and the children of the devil: whosoever doeth not righteousness is not of God, neither he that loveth not his brother.
1JOHN|3|11|For this is the message that ye heard from the beginning, that we should love one another.
1JOHN|3|12|Not as Cain, who was of that wicked one, and slew his brother. And wherefore slew he him? Because his own works were evil, and his brother's righteous.
1JOHN|3|13|Marvel not, my brethren, if the world hate you.
1JOHN|3|14|We know that we have passed from death unto life, because we love the brethren. He that loveth not his brother abideth in death.
1JOHN|3|15|Whosoever hateth his brother is a murderer: and ye know that no murderer hath eternal life abiding in him.
1JOHN|3|16|Hereby perceive we the love of God, because he laid down his life for us: and we ought to lay down our lives for the brethren.
1JOHN|3|17|But whoso hath this world's good, and seeth his brother have need, and shutteth up his bowels of compassion from him, how dwelleth the love of God in him?
1JOHN|3|18|My little children, let us not love in word, neither in tongue; but in deed and in truth.
1JOHN|3|19|And hereby we know that we are of the truth, and shall assure our hearts before him.
1JOHN|3|20|For if our heart condemn us, God is greater than our heart, and knoweth all things.
1JOHN|3|21|Beloved, if our heart condemn us not, then have we confidence toward God.
1JOHN|3|22|And whatsoever we ask, we receive of him, because we keep his commandments, and do those things that are pleasing in his sight.
1JOHN|3|23|And this is his commandment, That we should believe on the name of his Son Jesus Christ, and love one another, as he gave us commandment.
1JOHN|3|24|And he that keepeth his commandments dwelleth in him, and he in him. And hereby we know that he abideth in us, by the Spirit which he hath given us.
1JOHN|4|1|Beloved, believe not every spirit, but try the spirits whether they are of God: because many false prophets are gone out into the world.
1JOHN|4|2|Hereby know ye the Spirit of God: Every spirit that confesseth that Jesus Christ is come in the flesh is of God:
1JOHN|4|3|And every spirit that confesseth not that Jesus Christ is come in the flesh is not of God: and this is that spirit of antichrist, whereof ye have heard that it should come; and even now already is it in the world.
1JOHN|4|4|Ye are of God, little children, and have overcome them: because greater is he that is in you, than he that is in the world.
1JOHN|4|5|They are of the world: therefore speak they of the world, and the world heareth them.
1JOHN|4|6|We are of God: he that knoweth God heareth us; he that is not of God heareth not us. Hereby know we the spirit of truth, and the spirit of error.
1JOHN|4|7|Beloved, let us love one another: for love is of God; and every one that loveth is born of God, and knoweth God.
1JOHN|4|8|He that loveth not knoweth not God; for God is love.
1JOHN|4|9|In this was manifested the love of God toward us, because that God sent his only begotten Son into the world, that we might live through him.
1JOHN|4|10|Herein is love, not that we loved God, but that he loved us, and sent his Son to be the propitiation for our sins.
1JOHN|4|11|Beloved, if God so loved us, we ought also to love one another.
1JOHN|4|12|No man hath seen God at any time. If we love one another, God dwelleth in us, and his love is perfected in us.
1JOHN|4|13|Hereby know we that we dwell in him, and he in us, because he hath given us of his Spirit.
1JOHN|4|14|And we have seen and do testify that the Father sent the Son to be the Saviour of the world.
1JOHN|4|15|Whosoever shall confess that Jesus is the Son of God, God dwelleth in him, and he in God.
1JOHN|4|16|And we have known and believed the love that God hath to us. God is love; and he that dwelleth in love dwelleth in God, and God in him.
1JOHN|4|17|Herein is our love made perfect, that we may have boldness in the day of judgment: because as he is, so are we in this world.
1JOHN|4|18|There is no fear in love; but perfect love casteth out fear: because fear hath torment. He that feareth is not made perfect in love.
1JOHN|4|19|We love him, because he first loved us.
1JOHN|4|20|If a man say, I love God, and hateth his brother, he is a liar: for he that loveth not his brother whom he hath seen, how can he love God whom he hath not seen?
1JOHN|4|21|And this commandment have we from him, That he who loveth God love his brother also.
1JOHN|5|1|Whosoever believeth that Jesus is the Christ is born of God: and every one that loveth him that begat loveth him also that is begotten of him.
1JOHN|5|2|By this we know that we love the children of God, when we love God, and keep his commandments.
1JOHN|5|3|For this is the love of God, that we keep his commandments: and his commandments are not grievous.
1JOHN|5|4|For whatsoever is born of God overcometh the world: and this is the victory that overcometh the world, even our faith.
1JOHN|5|5|Who is he that overcometh the world, but he that believeth that Jesus is the Son of God?
1JOHN|5|6|This is he that came by water and blood, even Jesus Christ; not by water only, but by water and blood. And it is the Spirit that beareth witness, because the Spirit is truth.
1JOHN|5|7|For there are three that bear record in heaven, the Father, the Word, and the Holy Ghost: and these three are one.
1JOHN|5|8|And there are three that bear witness in earth, the Spirit, and the water, and the blood: and these three agree in one.
1JOHN|5|9|If we receive the witness of men, the witness of God is greater: for this is the witness of God which he hath testified of his Son.
1JOHN|5|10|He that believeth on the Son of God hath the witness in himself: he that believeth not God hath made him a liar; because he believeth not the record that God gave of his Son.
1JOHN|5|11|And this is the record, that God hath given to us eternal life, and this life is in his Son.
1JOHN|5|12|He that hath the Son hath life; and he that hath not the Son of God hath not life.
1JOHN|5|13|These things have I written unto you that believe on the name of the Son of God; that ye may know that ye have eternal life, and that ye may believe on the name of the Son of God.
1JOHN|5|14|And this is the confidence that we have in him, that, if we ask any thing according to his will, he heareth us:
1JOHN|5|15|And if we know that he hear us, whatsoever we ask, we know that we have the petitions that we desired of him.
1JOHN|5|16|If any man see his brother sin a sin which is not unto death, he shall ask, and he shall give him life for them that sin not unto death. There is a sin unto death: I do not say that he shall pray for it.
1JOHN|5|17|All unrighteousness is sin: and there is a sin not unto death.
1JOHN|5|18|We know that whosoever is born of God sinneth not; but he that is begotten of God keepeth himself, and that wicked one toucheth him not.
1JOHN|5|19|And we know that we are of God, and the whole world lieth in wickedness.
1JOHN|5|20|And we know that the Son of God is come, and hath given us an understanding, that we may know him that is true, and we are in him that is true, even in his Son Jesus Christ. This is the true God, and eternal life.
1JOHN|5|21|Little children, keep yourselves from idols. Amen.
