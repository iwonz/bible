MATT|1|1|The book of the genealogy of Jesus Christ, the son of David, the son of Abraham.
MATT|1|2|Abraham was the father of Isaac, and Isaac the father of Jacob, and Jacob the father of Judah and his brothers,
MATT|1|3|and Judah the father of Perez and Zerah by Tamar, and Perez the father of Hezron, and Hezron the father of Ram,
MATT|1|4|and Ram the father of Amminadab, and Amminadab the father of Nahshon, and Nahshon the father of Salmon,
MATT|1|5|and Salmon the father of Boaz by Rahab, and Boaz the father of Obed by Ruth, and Obed the father of Jesse,
MATT|1|6|and Jesse the father of David the king. And David was the father of Solomon by the wife of Uriah,
MATT|1|7|and Solomon the father of Rehoboam, and Rehoboam the father of Abijah, and Abijah the father of Asaph,
MATT|1|8|and Asaph the father of Jehoshaphat, and Jehoshaphat the father of Joram, and Joram the father of Uzziah,
MATT|1|9|and Uzziah the father of Jotham, and Jotham the father of Ahaz, and Ahaz the father of Hezekiah,
MATT|1|10|and Hezekiah the father of Manasseh, and Manasseh the father of Amos, and Amos the father of Josiah,
MATT|1|11|and Josiah the father of Jechoniah and his brothers, at the time of the deportation to Babylon.
MATT|1|12|And after the deportation to Babylon: Jechoniah was the father of Shealtiel, and Shealtiel the father of Zerubbabel,
MATT|1|13|and Zerubbabel the father of Abiud, and Abiud the father of Eliakim, and Eliakim the father of Azor,
MATT|1|14|and Azor the father of Zadok, and Zadok the father of Achim, and Achim the father of Eliud,
MATT|1|15|and Eliud the father of Eleazar, and Eleazar the father of Matthan, and Matthan the father of Jacob,
MATT|1|16|and Jacob the father of Joseph the husband of Mary, of whom Jesus was born, who is called Christ.
MATT|1|17|So all the generations from Abraham to David were fourteen generations, and from David to the deportation to Babylon fourteen generations, and from the deportation to Babylon to the Christ fourteen generations.
MATT|1|18|Now the birth of Jesus Christ took place in this way. When his mother Mary had been betrothed to Joseph, before they came together she was found to be with child from the Holy Spirit.
MATT|1|19|And her husband Joseph, being a just man and unwilling to put her to shame, resolved to divorce her quietly.
MATT|1|20|But as he considered these things, behold, an angel of the Lord appeared to him in a dream, saying, "Joseph, son of David, do not fear to take Mary as your wife, for that which is conceived in her is from the Holy Spirit.
MATT|1|21|She will bear a son, and you shall call his name Jesus, for he will save his people from their sins."
MATT|1|22|All this took place to fulfill what the Lord had spoken by the prophet:
MATT|1|23|"Behold, the virgin shall conceive and bear a son, and they shall call his name Immanuel" (which means, God with us).
MATT|1|24|When Joseph woke from sleep, he did as the angel of the Lord commanded him: he took his wife,
MATT|1|25|but knew her not until she had given birth to a son. And he called his name Jesus.
MATT|2|1|Now after Jesus was born in Bethlehem of Judea in the days of Herod the king, behold, wise men from the east came to Jerusalem,
MATT|2|2|saying, "Where is he who has been born king of the Jews? For we saw his star when it rose and have come to worship him."
MATT|2|3|When Herod the king heard this, he was troubled, and all Jerusalem with him;
MATT|2|4|and assembling all the chief priests and scribes of the people, he inquired of them where the Christ was to be born.
MATT|2|5|They told him, "In Bethlehem of Judea, for so it is written by the prophet:
MATT|2|6|"' And you, O Bethlehem, in the land of Judah, are by no means least among the rulers of Judah; for from you shall come a ruler who will shepherd my people Israel.'"
MATT|2|7|Then Herod summoned the wise men secretly and ascertained from them what time the star had appeared.
MATT|2|8|And he sent them to Bethlehem, saying, "Go and search diligently for the child, and when you have found him, bring me word, that I too may come and worship him."
MATT|2|9|After listening to the king, they went on their way. And behold, the star that they had seen when it rose went before them until it came to rest over the place where the child was.
MATT|2|10|When they saw the star, they rejoiced exceedingly with great joy.
MATT|2|11|And going into the house they saw the child with Mary his mother, and they fell down and worshiped him. Then, opening their treasures, they offered him gifts, gold and frankincense and myrrh.
MATT|2|12|And being warned in a dream not to return to Herod, they departed to their own country by another way.
MATT|2|13|Now when they had departed, behold, an angel of the Lord appeared to Joseph in a dream and said, "Rise, take the child and his mother, and flee to Egypt, and remain there until I tell you, for Herod is about to search for the child, to destroy him."
MATT|2|14|And he rose and took the child and his mother by night and departed to Egypt
MATT|2|15|and remained there until the death of Herod. This was to fulfill what the Lord had spoken by the prophet, "Out of Egypt I called my son."
MATT|2|16|Then Herod, when he saw that he had been tricked by the wise men, became furious, and he sent and killed all the male children in Bethlehem and in all that region who were two years old or under, according to the time that he had ascertained from the wise men.
MATT|2|17|Then was fulfilled what was spoken by the prophet Jeremiah:
MATT|2|18|"A voice was heard in Ramah, weeping and loud lamentation, Rachel weeping for her children; she refused to be comforted, because they are no more."
MATT|2|19|But when Herod died, behold, an angel of the Lord appeared in a dream to Joseph in Egypt,
MATT|2|20|saying, "Rise, take the child and his mother and go to the land of Israel, for those who sought the child's life are dead."
MATT|2|21|And he rose and took the child and his mother and went to the land of Israel.
MATT|2|22|But when he heard that Archelaus was reigning over Judea in place of his father Herod, he was afraid to go there, and being warned in a dream he withdrew to the district of Galilee.
MATT|2|23|And he went and lived in a city called Nazareth, that what was spoken by the prophets might be fulfilled: "He shall be called a Nazarene."
MATT|3|1|In those days John the Baptist came preaching in the wilderness of Judea,
MATT|3|2|"Repent, for the kingdom of heaven is at hand."
MATT|3|3|For this is he who was spoken of by the prophet Isaiah when he said, "The voice of one crying in the wilderness: Prepare the way of the Lord; make his paths straight."
MATT|3|4|Now John wore a garment of camel's hair and a leather belt around his waist, and his food was locusts and wild honey.
MATT|3|5|Then Jerusalem and all Judea and all the region about the Jordan were going out to him,
MATT|3|6|and they were baptized by him in the river Jordan, confessing their sins.
MATT|3|7|But when he saw many of the Pharisees and Sadducees coming for baptism, he said to them, "You brood of vipers! Who warned you to flee from the wrath to come?
MATT|3|8|Bear fruit in keeping with repentance.
MATT|3|9|And do not presume to say to yourselves, 'We have Abraham as our father,' for I tell you, God is able from these stones to raise up children for Abraham.
MATT|3|10|Even now the axe is laid to the root of the trees. Every tree therefore that does not bear good fruit is cut down and thrown into the fire.
MATT|3|11|"I baptize you with water for repentance, but he who is coming after me is mightier than I, whose sandals I am not worthy to carry. He will baptize you with the Holy Spirit and with fire.
MATT|3|12|His winnowing fork is in his hand, and he will clear his threshing floor and gather his wheat into the barn, but the chaff he will burn with unquenchable fire."
MATT|3|13|Then Jesus came from Galilee to the Jordan to John, to be baptized by him.
MATT|3|14|John would have prevented him, saying, "I need to be baptized by you, and do you come to me?"
MATT|3|15|But Jesus answered him, "Let it be so now, for thus it is fitting for us to fulfill all righteousness." Then he consented.
MATT|3|16|And when Jesus was baptized, immediately he went up from the water, and behold, the heavens were opened to him, and he saw the Spirit of God descending like a dove and coming to rest on him;
MATT|3|17|and behold, a voice from heaven said, "This is my beloved Son, with whom I am well pleased."
MATT|4|1|Then Jesus was led up by the Spirit into the wilderness to be tempted by the devil.
MATT|4|2|And after fasting forty days and forty nights, he was hungry.
MATT|4|3|And the tempter came and said to him, "If you are the Son of God, command these stones to become loaves of bread."
MATT|4|4|But he answered, "It is written, "' Man shall not live by bread alone, but by every word that comes from the mouth of God.'"
MATT|4|5|Then the devil took him to the holy city and set him on the pinnacle of the temple
MATT|4|6|and said to him, "If you are the Son of God, throw yourself down, for it is written, "' He will command his angels concerning you,' and "'On their hands they will bear you up, lest you strike your foot against a stone.'"
MATT|4|7|Jesus said to him, "Again it is written, 'You shall not put the Lord your God to the test.'"
MATT|4|8|Again, the devil took him to a very high mountain and showed him all the kingdoms of the world and their glory.
MATT|4|9|And he said to him, "All these I will give you, if you will fall down and worship me."
MATT|4|10|Then Jesus said to him, "Be gone, Satan! For it is written, "' You shall worship the Lord your God and him only shall you serve.'"
MATT|4|11|Then the devil left him, and behold, angels came and were ministering to him.
MATT|4|12|Now when he heard that John had been arrested, he withdrew into Galilee.
MATT|4|13|And leaving Nazareth he went and lived in Capernaum by the sea, in the territory of Zebulun and Naphtali,
MATT|4|14|so that what was spoken by the prophet Isaiah might be fulfilled:
MATT|4|15|"The land of Zebulun and the land of Naphtali, the way of the sea, beyond the Jordan, Galilee of the Gentiles-
MATT|4|16|the people dwelling in darkness have seen a great light, and for those dwelling in the region and shadow of death, on them a light has dawned."
MATT|4|17|From that time Jesus began to preach, saying, "Repent, for the kingdom of heaven is at hand."
MATT|4|18|While walking by the Sea of Galilee, he saw two brothers, Simon (who is called Peter) and Andrew his brother, casting a net into the sea, for they were fishermen.
MATT|4|19|And he said to them, "Follow me, and I will make you fishers of men."
MATT|4|20|Immediately they left their nets and followed him.
MATT|4|21|And going on from there he saw two other brothers, James the son of Zebedee and John his brother, in the boat with Zebedee their father, mending their nets, and he called them.
MATT|4|22|Immediately they left the boat and their father and followed him.
MATT|4|23|And he went throughout all Galilee, teaching in their synagogues and proclaiming the gospel of the kingdom and healing every disease and every affliction among the people.
MATT|4|24|So his fame spread throughout all Syria, and they brought him all the sick, those afflicted with various diseases and pains, those oppressed by demons, epileptics, and paralytics, and he healed them.
MATT|4|25|And great crowds followed him from Galilee and the Decapolis, and from Jerusalem and Judea, and from beyond the Jordan.
MATT|5|1|Seeing the crowds, he went up on the mountain, and when he sat down, his disciples came to him.
MATT|5|2|And he opened his mouth and taught them, saying:
MATT|5|3|"Blessed are the poor in spirit, for theirs is the kingdom of heaven.
MATT|5|4|"Blessed are those who mourn, for they shall be comforted.
MATT|5|5|"Blessed are the meek, for they shall inherit the earth.
MATT|5|6|"Blessed are those who hunger and thirst for righteousness, for they shall be satisfied.
MATT|5|7|"Blessed are the merciful, for they shall receive mercy.
MATT|5|8|"Blessed are the pure in heart, for they shall see God.
MATT|5|9|"Blessed are the peacemakers, for they shall be called sons of God.
MATT|5|10|"Blessed are those who are persecuted for righteousness' sake, for theirs is the kingdom of heaven.
MATT|5|11|"Blessed are you when others revile you and persecute you and utter all kinds of evil against you falsely on my account.
MATT|5|12|Rejoice and be glad, for your reward is great in heaven, for so they persecuted the prophets who were before you.
MATT|5|13|"You are the salt of the earth, but if salt has lost its taste, how shall its saltiness be restored? It is no longer good for anything except to be thrown out and trampled under people's feet.
MATT|5|14|"You are the light of the world. A city set on a hill cannot be hidden.
MATT|5|15|Nor do people light a lamp and put it under a basket, but on a stand, and it gives light to all in the house.
MATT|5|16|In the same way, let your light shine before others, so that they may see your good works and give glory to your Father who is in heaven.
MATT|5|17|"Do not think that I have come to abolish the Law or the Prophets; I have not come to abolish them but to fulfill them.
MATT|5|18|For truly, I say to you, until heaven and earth pass away, not an iota, not a dot, will pass from the Law until all is accomplished.
MATT|5|19|Therefore whoever relaxes one of the least of these commandments and teaches others to do the same will be called least in the kingdom of heaven, but whoever does them and teaches them will be called great in the kingdom of heaven.
MATT|5|20|For I tell you, unless your righteousness exceeds that of the scribes and Pharisees, you will never enter the kingdom of heaven.
MATT|5|21|"You have heard that it was said to those of old, 'You shall not murder; and whoever murders will be liable to judgment.'
MATT|5|22|But I say to you that everyone who is angry with his brother will be liable to judgment; whoever insults his brother will be liable to the council; and whoever says, 'You fool!' will be liable to the hell of fire.
MATT|5|23|So if you are offering your gift at the altar and there remember that your brother has something against you,
MATT|5|24|leave your gift there before the altar and go. First be reconciled to your brother, and then come and offer your gift.
MATT|5|25|Come to terms quickly with your accuser while you are going with him to court, lest your accuser hand you over to the judge, and the judge to the guard, and you be put in prison.
MATT|5|26|Truly, I say to you, you will never get out until you have paid the last penny.
MATT|5|27|"You have heard that it was said, 'You shall not commit adultery.'
MATT|5|28|But I say to you that everyone who looks at a woman with lustful intent has already committed adultery with her in his heart.
MATT|5|29|If your right eye causes you to sin, tear it out and throw it away. For it is better that you lose one of your members than that your whole body be thrown into hell.
MATT|5|30|And if your right hand causes you to sin, cut it off and throw it away. For it is better that you lose one of your members than that your whole body go into hell.
MATT|5|31|"It was also said, 'Whoever divorces his wife, let him give her a certificate of divorce.'
MATT|5|32|But I say to you that everyone who divorces his wife, except on the ground of sexual immorality, makes her commit adultery. And whoever marries a divorced woman commits adultery.
MATT|5|33|"Again you have heard that it was said to those of old, 'You shall not swear falsely, but shall perform to the Lord what you have sworn.'
MATT|5|34|But I say to you, Do not take an oath at all, either by heaven, for it is the throne of God,
MATT|5|35|or by the earth, for it is his footstool, or by Jerusalem, for it is the city of the great King.
MATT|5|36|And do not take an oath by your head, for you cannot make one hair white or black.
MATT|5|37|Let what you say be simply 'Yes' or 'No'; anything more than this comes from evil.
MATT|5|38|"You have heard that it was said, 'An eye for an eye and a tooth for a tooth.'
MATT|5|39|But I say to you, Do not resist the one who is evil. But if anyone slaps you on the right cheek, turn to him the other also.
MATT|5|40|And if anyone would sue you and take your tunic, let him have your cloak as well.
MATT|5|41|And if anyone forces you to go one mile, go with him two miles.
MATT|5|42|Give to the one who begs from you, and do not refuse the one who would borrow from you.
MATT|5|43|"You have heard that it was said, 'You shall love your neighbor and hate your enemy.'
MATT|5|44|But I say to you, Love your enemies and pray for those who persecute you,
MATT|5|45|so that you may be sons of your Father who is in heaven. For he makes his sun rise on the evil and on the good, and sends rain on the just and on the unjust.
MATT|5|46|For if you love those who love you, what reward do you have? Do not even the tax collectors do the same?
MATT|5|47|And if you greet only your brothers, what more are you doing than others? Do not even the Gentiles do the same?
MATT|5|48|You therefore must be perfect, as your heavenly Father is perfect.
MATT|6|1|"Beware of practicing your righteousness before other people in order to be seen by them, for then you will have no reward from your Father who is in heaven.
MATT|6|2|"Thus, when you give to the needy, sound no trumpet before you, as the hypocrites do in the synagogues and in the streets, that they may be praised by others. Truly, I say to you, they have received their reward.
MATT|6|3|But when you give to the needy, do not let your left hand know what your right hand is doing,
MATT|6|4|so that your giving may be in secret. And your Father who sees in secret will reward you.
MATT|6|5|"And when you pray, you must not be like the hypocrites. For they love to stand and pray in the synagogues and at the street corners, that they may be seen by others. Truly, I say to you, they have received their reward.
MATT|6|6|But when you pray, go into your room and shut the door and pray to your Father who is in secret. And your Father who sees in secret will reward you.
MATT|6|7|"And when you pray, do not heap up empty phrases as the Gentiles do, for they think that they will be heard for their many words.
MATT|6|8|Do not be like them, for your Father knows what you need before you ask him.
MATT|6|9|Pray then like this: "Our Father in heaven, hallowed be your name.
MATT|6|10|Your kingdom come, your will be done, on earth as it is in heaven.
MATT|6|11|Give us this day our daily bread,
MATT|6|12|and forgive us our debts, as we also have forgiven our debtors.
MATT|6|13|And lead us not into temptation, but deliver us from evil.
MATT|6|14|For if you forgive others their trespasses, your heavenly Father will also forgive you,
MATT|6|15|but if you do not forgive others their trespasses, neither will your Father forgive your trespasses.
MATT|6|16|"And when you fast, do not look gloomy like the hypocrites, for they disfigure their faces that their fasting may be seen by others. Truly, I say to you, they have received their reward.
MATT|6|17|But when you fast, anoint your head and wash your face,
MATT|6|18|that your fasting may not be seen by others but by your Father who is in secret. And your Father who sees in secret will reward you.
MATT|6|19|"Do not lay up for yourselves treasures on earth, where moth and rust destroy and where thieves break in and steal,
MATT|6|20|but lay up for yourselves treasures in heaven, where neither moth nor rust destroys and where thieves do not break in and steal.
MATT|6|21|For where your treasure is, there your heart will be also.
MATT|6|22|"The eye is the lamp of the body. So, if your eye is healthy, your whole body will be full of light,
MATT|6|23|but if your eye is bad, your whole body will be full of darkness. If then the light in you is darkness, how great is the darkness!
MATT|6|24|"No one can serve two masters, for either he will hate the one and love the other, or he will be devoted to the one and despise the other. You cannot serve God and money.
MATT|6|25|"Therefore I tell you, do not be anxious about your life, what you will eat or what you will drink, nor about your body, what you will put on. Is not life more than food, and the body more than clothing?
MATT|6|26|Look at the birds of the air: they neither sow nor reap nor gather into barns, and yet your heavenly Father feeds them. Are you not of more value than they?
MATT|6|27|And which of you by being anxious can add a single hour to his span of life?
MATT|6|28|And why are you anxious about clothing? Consider the lilies of the field, how they grow: they neither toil nor spin,
MATT|6|29|yet I tell you, even Solomon in all his glory was not arrayed like one of these.
MATT|6|30|But if God so clothes the grass of the field, which today is alive and tomorrow is thrown into the oven, will he not much more clothe you, O you of little faith?
MATT|6|31|Therefore do not be anxious, saying, 'What shall we eat?' or 'What shall we drink?' or 'What shall we wear?'
MATT|6|32|For the Gentiles seek after all these things, and your heavenly Father knows that you need them all.
MATT|6|33|But seek first the kingdom of God and his righteousness, and all these things will be added to you.
MATT|6|34|"Therefore do not be anxious about tomorrow, for tomorrow will be anxious for itself. Sufficient for the day is its own trouble.
MATT|7|1|"Judge not, that you be not judged.
MATT|7|2|For with the judgment you pronounce you will be judged, and with the measure you use it will be measured to you.
MATT|7|3|Why do you see the speck that is in your brother's eye, but do not notice the log that is in your own eye?
MATT|7|4|Or how can you say to your brother, 'Let me take the speck out of your eye,' when there is the log in your own eye?
MATT|7|5|You hypocrite, first take the log out of your own eye, and then you will see clearly to take the speck out of your brother's eye.
MATT|7|6|"Do not give dogs what is holy, and do not throw your pearls before pigs, lest they trample them underfoot and turn to attack you.
MATT|7|7|"Ask, and it will be given to you; seek, and you will find; knock, and it will be opened to you.
MATT|7|8|For everyone who asks receives, and the one who seeks finds, and to the one who knocks it will be opened.
MATT|7|9|Or which one of you, if his son asks him for bread, will give him a stone?
MATT|7|10|Or if he asks for a fish, will give him a serpent?
MATT|7|11|If you then, who are evil, know how to give good gifts to your children, how much more will your Father who is in heaven give good things to those who ask him!
MATT|7|12|"So whatever you wish that others would do to you, do also to them, for this is the Law and the Prophets.
MATT|7|13|"Enter by the narrow gate. For the gate is wide and the way is easy that leads to destruction, and those who enter by it are many.
MATT|7|14|For the gate is narrow and the way is hard that leads to life, and those who find it are few.
MATT|7|15|"Beware of false prophets, who come to you in sheep's clothing but inwardly are ravenous wolves.
MATT|7|16|You will recognize them by their fruits. Are grapes gathered from thornbushes, or figs from thistles?
MATT|7|17|So, every healthy tree bears good fruit, but the diseased tree bears bad fruit.
MATT|7|18|A healthy tree cannot bear bad fruit, nor can a diseased tree bear good fruit.
MATT|7|19|Every tree that does not bear good fruit is cut down and thrown into the fire.
MATT|7|20|Thus you will recognize them by their fruits.
MATT|7|21|"Not everyone who says to me, 'Lord, Lord,' will enter the kingdom of heaven, but the one who does the will of my Father who is in heaven.
MATT|7|22|On that day many will say to me, 'Lord, Lord, did we not prophesy in your name, and cast out demons in your name, and do many mighty works in your name?'
MATT|7|23|And then will I declare to them, 'I never knew you; depart from me, you workers of lawlessness.'
MATT|7|24|"Everyone then who hears these words of mine and does them will be like a wise man who built his house on the rock.
MATT|7|25|And the rain fell, and the floods came, and the winds blew and beat on that house, but it did not fall, because it had been founded on the rock.
MATT|7|26|And everyone who hears these words of mine and does not do them will be like a foolish man who built his house on the sand.
MATT|7|27|And the rain fell, and the floods came, and the winds blew and beat against that house, and it fell, and great was the fall of it."
MATT|7|28|And when Jesus finished these sayings, the crowds were astonished at his teaching,
MATT|7|29|for he was teaching them as one who had authority, and not as their scribes.
MATT|8|1|When he came down from the mountain, great crowds followed him.
MATT|8|2|And behold, a leper came to him and knelt before him, saying, "Lord, if you will, you can make me clean."
MATT|8|3|And Jesus stretched out his hand and touched him, saying, "I will; be clean." And immediately his leprosy was cleansed.
MATT|8|4|And Jesus said to him, "See that you say nothing to anyone, but go, show yourself to the priest and offer the gift that Moses commanded, for a proof to them."
MATT|8|5|When he entered Capernaum, a centurion came forward to him, appealing to him,
MATT|8|6|"Lord, my servant is lying paralyzed at home, suffering terribly."
MATT|8|7|And he said to him, "I will come and heal him."
MATT|8|8|But the centurion replied, "Lord, I am not worthy to have you come under my roof, but only say the word, and my servant will be healed.
MATT|8|9|For I too am a man under authority, with soldiers under me. And I say to one, 'Go,' and he goes, and to another, 'Come,' and he comes, and to my servant, 'Do this,' and he does it."
MATT|8|10|When Jesus heard this, he marveled and said to those who followed him, "Truly, I tell you, with no one in Israel have I found such faith.
MATT|8|11|I tell you, many will come from east and west and recline at table with Abraham, Isaac, and Jacob in the kingdom of heaven,
MATT|8|12|while the sons of the kingdom will be thrown into the outer darkness. In that place there will be weeping and gnashing of teeth."
MATT|8|13|And to the centurion Jesus said, "Go; let it be done for you as you have believed." And the servant was healed at that very moment.
MATT|8|14|And when Jesus entered Peter's house, he saw his mother-in-law lying sick with a fever.
MATT|8|15|He touched her hand, and the fever left her, and she rose and began to serve him.
MATT|8|16|That evening they brought to him many who were oppressed by demons, and he cast out the spirits with a word and healed all who were sick.
MATT|8|17|This was to fulfill what was spoken by the prophet Isaiah: "He took our illnesses and bore our diseases."
MATT|8|18|Now when Jesus saw a great crowd around him, he gave orders to go over to the other side.
MATT|8|19|And a scribe came up and said to him, "Teacher, I will follow you wherever you go."
MATT|8|20|And Jesus said to him, "Foxes have holes, and birds of the air have nests, but the Son of Man has nowhere to lay his head."
MATT|8|21|Another of the disciples said to him, "Lord, let me first go and bury my father."
MATT|8|22|And Jesus said to him, "Follow me, and leave the dead to bury their own dead."
MATT|8|23|And when he got into the boat, his disciples followed him.
MATT|8|24|And behold, there arose a great storm on the sea, so that the boat was being swamped by the waves; but he was asleep.
MATT|8|25|And they went and woke him, saying, "Save us, Lord; we are perishing."
MATT|8|26|And he said to them, "Why are you afraid, O you of little faith?" Then he rose and rebuked the winds and the sea, and there was a great calm.
MATT|8|27|And the men marveled, saying, "What sort of man is this, that even winds and sea obey him?"
MATT|8|28|And when he came to the other side, to the country of the Gadarenes, two demon-possessed men met him, coming out of the tombs, so fierce that no one could pass that way.
MATT|8|29|And behold, they cried out, "What have you to do with us, O Son of God? Have you come here to torment us before the time?"
MATT|8|30|Now a herd of many pigs was feeding at some distance from them.
MATT|8|31|And the demons begged him, saying, "If you cast us out, send us away into the herd of pigs."
MATT|8|32|And he said to them, "Go." So they came out and went into the pigs, and behold, the whole herd rushed down the steep bank into the sea and drowned in the waters.
MATT|8|33|The herdsmen fled, and going into the city they told everything, especially what had happened to the demon-possessed men.
MATT|8|34|And behold, all the city came out to meet Jesus, and when they saw him, they begged him to leave their region.
MATT|9|1|And getting into a boat he crossed over and came to his own city.
MATT|9|2|And behold, some people brought to him a paralytic, lying on a bed. And when Jesus saw their faith, he said to the paralytic, "Take heart, my son; your sins are forgiven."
MATT|9|3|And behold, some of the scribes said to themselves, "This man is blaspheming."
MATT|9|4|But Jesus, knowing their thoughts, said, "Why do you think evil in your hearts?
MATT|9|5|For which is easier, to say, 'Your sins are forgiven,' or to say, 'Rise and walk'?
MATT|9|6|But that you may know that the Son of Man has authority on earth to forgive sins"- he then said to the paralytic- "Rise, pick up your bed and go home."
MATT|9|7|And he rose and went home.
MATT|9|8|When the crowds saw it, they were afraid, and they glorified God, who had given such authority to men.
MATT|9|9|As Jesus passed on from there, he saw a man called Matthew sitting at the tax booth, and he said to him, "Follow me." And he rose and followed him.
MATT|9|10|And as Jesus reclined at table in the house, behold, many tax collectors and sinners came and were reclining with Jesus and his disciples.
MATT|9|11|And when the Pharisees saw this, they said to his disciples, "Why does your teacher eat with tax collectors and sinners?"
MATT|9|12|But when he heard it, he said, "Those who are well have no need of a physician, but those who are sick.
MATT|9|13|Go and learn what this means, 'I desire mercy, and not sacrifice.' For I came not to call the righteous, but sinners."
MATT|9|14|Then the disciples of John came to him, saying, "Why do we and the Pharisees fast, but your disciples do not fast?"
MATT|9|15|And Jesus said to them, "Can the wedding guests mourn as long as the bridegroom is with them? The days will come when the bridegroom is taken away from them, and then they will fast.
MATT|9|16|No one puts a piece of unshrunk cloth on an old garment, for the patch tears away from the garment, and a worse tear is made.
MATT|9|17|Neither is new wine put into old wineskins. If it is, the skins burst and the wine is spilled and the skins are destroyed. But new wine is put into fresh wineskins, and so both are preserved."
MATT|9|18|While he was saying these things to them, behold, a ruler came in and knelt before him, saying, "My daughter has just died, but come and lay your hand on her, and she will live."
MATT|9|19|And Jesus rose and followed him, with his disciples.
MATT|9|20|And behold, a woman who had suffered from a discharge of blood for twelve years came up behind him and touched the fringe of his garment,
MATT|9|21|for she said to herself, "If I only touch his garment, I will be made well."
MATT|9|22|Jesus turned, and seeing her he said, "Take heart, daughter; your faith has made you well." And instantly the woman was made well.
MATT|9|23|And when Jesus came to the ruler's house and saw the flute players and the crowd making a commotion,
MATT|9|24|he said, "Go away, for the girl is not dead but sleeping." And they laughed at him.
MATT|9|25|But when the crowd had been put outside, he went in and took her by the hand, and the girl arose.
MATT|9|26|And the report of this went through all that district.
MATT|9|27|And as Jesus passed on from there, two blind men followed him, crying aloud, "Have mercy on us, Son of David."
MATT|9|28|When he entered the house, the blind men came to him, and Jesus said to them, "Do you believe that I am able to do this?" They said to him, "Yes, Lord."
MATT|9|29|Then he touched their eyes, saying, "According to your faith be it done to you."
MATT|9|30|And their eyes were opened. And Jesus sternly warned them, "See that no one knows about it."
MATT|9|31|But they went away and spread his fame through all that district.
MATT|9|32|As they were going away, behold, a demon-oppressed man who was mute was brought to him.
MATT|9|33|And when the demon had been cast out, the mute man spoke. And the crowds marveled, saying, "Never was anything like this seen in Israel."
MATT|9|34|But the Pharisees said, "He casts out demons by the prince of demons."
MATT|9|35|And Jesus went throughout all the cities and villages, teaching in their synagogues and proclaiming the gospel of the kingdom and healing every disease and every affliction.
MATT|9|36|When he saw the crowds, he had compassion for them, because they were harassed and helpless, like sheep without a shepherd.
MATT|9|37|Then he said to his disciples, "The harvest is plentiful, but the laborers are few;
MATT|9|38|therefore pray earnestly to the Lord of the harvest to send out laborers into his harvest."
MATT|10|1|And he called to him his twelve disciples and gave them authority over unclean spirits, to cast them out, and to heal every disease and every affliction.
MATT|10|2|The names of the twelve apostles are these: first, Simon, who is called Peter, and Andrew his brother; James the son of Zebedee, and John his brother;
MATT|10|3|Philip and Bartholomew; Thomas and Matthew the tax collector; James the son of Alphaeus, and Thaddaeus;
MATT|10|4|Simon the Cananaean, and Judas Iscariot, who betrayed him.
MATT|10|5|These twelve Jesus sent out, instructing them, "Go nowhere among the Gentiles and enter no town of the Samaritans,
MATT|10|6|but go rather to the lost sheep of the house of Israel.
MATT|10|7|And proclaim as you go, saying, 'The kingdom of heaven is at hand.'
MATT|10|8|Heal the sick, raise the dead, cleanse lepers, cast out demons. You received without paying; give without pay.
MATT|10|9|Acquire no gold nor silver nor copper for your belts,
MATT|10|10|no bag for your journey, nor two tunics nor sandals nor a staff, for the laborer deserves his food.
MATT|10|11|And whatever town or village you enter, find out who is worthy in it and stay there until you depart.
MATT|10|12|As you enter the house, greet it.
MATT|10|13|And if the house is worthy, let your peace come upon it, but if it is not worthy, let your peace return to you.
MATT|10|14|And if anyone will not receive you or listen to your words, shake off the dust from your feet when you leave that house or town.
MATT|10|15|Truly, I say to you, it will be more bearable on the day of judgment for the land of Sodom and Gomorrah than for that town.
MATT|10|16|"Behold, I am sending you out as sheep in the midst of wolves, so be wise as serpents and innocent as doves.
MATT|10|17|Beware of men, for they will deliver you over to courts and flog you in their synagogues,
MATT|10|18|and you will be dragged before governors and kings for my sake, to bear witness before them and the Gentiles.
MATT|10|19|When they deliver you over, do not be anxious how you are to speak or what you are to say, for what you are to say will be given to you in that hour.
MATT|10|20|For it is not you who speak, but the Spirit of your Father speaking through you.
MATT|10|21|Brother will deliver brother over to death, and the father his child, and children will rise against parents and have them put to death,
MATT|10|22|and you will be hated by all for my name's sake. But the one who endures to the end will be saved.
MATT|10|23|When they persecute you in one town, flee to the next, for truly, I say to you, you will not have gone through all the towns of Israel before the Son of Man comes.
MATT|10|24|"A disciple is not above his teacher, nor a servant above his master.
MATT|10|25|It is enough for the disciple to be like his teacher, and the servant like his master. If they have called the master of the house Beelzebul, how much more will they malign those of his household.
MATT|10|26|"So have no fear of them, for nothing is covered that will not be revealed, or hidden that will not be known.
MATT|10|27|What I tell you in the dark, say in the light, and what you hear whispered, proclaim on the housetops.
MATT|10|28|And do not fear those who kill the body but cannot kill the soul. Rather fear him who can destroy both soul and body in hell.
MATT|10|29|Are not two sparrows sold for a penny? And not one of them will fall to the ground apart from your Father.
MATT|10|30|But even the hairs of your head are all numbered.
MATT|10|31|Fear not, therefore; you are of more value than many sparrows.
MATT|10|32|So everyone who acknowledges me before men, I also will acknowledge before my Father who is in heaven,
MATT|10|33|but whoever denies me before men, I also will deny before my Father who is in heaven.
MATT|10|34|"Do not think that I have come to bring peace to the earth. I have not come to bring peace, but a sword.
MATT|10|35|For I have come to set a man against his father, and a daughter against her mother, and a daughter-in-law against her mother-in-law.
MATT|10|36|And a person's enemies will be those of his own household.
MATT|10|37|Whoever loves father or mother more than me is not worthy of me, and whoever loves son or daughter more than me is not worthy of me.
MATT|10|38|And whoever does not take his cross and follow me is not worthy of me.
MATT|10|39|Whoever finds his life will lose it, and whoever loses his life for my sake will find it.
MATT|10|40|"Whoever receives you receives me, and whoever receives me receives him who sent me.
MATT|10|41|The one who receives a prophet because he is a prophet will receive a prophet's reward, and the one who receives a righteous person because he is a righteous person will receive a righteous person's reward.
MATT|10|42|And whoever gives one of these little ones even a cup of cold water because he is a disciple, truly, I say to you, he will by no means lose his reward."
MATT|11|1|When Jesus had finished instructing his twelve disciples, he went on from there to teach and preach in their cities.
MATT|11|2|Now when John heard in prison about the deeds of the Christ, he sent word by his disciples
MATT|11|3|and said to him, "Are you the one who is to come, or shall we look for another?"
MATT|11|4|And Jesus answered them, "Go and tell John what you hear and see:
MATT|11|5|the blind receive their sight and the lame walk, lepers are cleansed and the deaf hear, and the dead are raised up, and the poor have good news preached to them.
MATT|11|6|And blessed is the one who is not offended by me."
MATT|11|7|As they went away, Jesus began to speak to the crowds concerning John: "What did you go out into the wilderness to see? A reed shaken by the wind?
MATT|11|8|What then did you go out to see? A man dressed in soft clothing? Behold, those who wear soft clothing are in kings' houses.
MATT|11|9|What then did you go out to see? A prophet? Yes, I tell you, and more than a prophet.
MATT|11|10|This is he of whom it is written, "' Behold, I send my messenger before your face, who will prepare your way before you.'
MATT|11|11|Truly, I say to you, among those born of women there has arisen no one greater than John the Baptist. Yet the one who is least in the kingdom of heaven is greater than he.
MATT|11|12|From the days of John the Baptist until now the kingdom of heaven has suffered violence, and the violent take it by force.
MATT|11|13|For all the Prophets and the Law prophesied until John,
MATT|11|14|and if you are willing to accept it, he is Elijah who is to come.
MATT|11|15|He who has ears to hear, let him hear.
MATT|11|16|"But to what shall I compare this generation? It is like children sitting in the marketplaces and calling to their playmates,
MATT|11|17|"'We played the flute for you, and you did not dance; we sang a dirge, and you did not mourn.'
MATT|11|18|For John came neither eating nor drinking, and they say, 'He has a demon.'
MATT|11|19|The Son of Man came eating and drinking, and they say, 'Look at him! A glutton and a drunkard, a friend of tax collectors and sinners!' Yet wisdom is justified by her deeds."
MATT|11|20|Then he began to denounce the cities where most of his mighty works had been done, because they did not repent.
MATT|11|21|"Woe to you, Chorazin! Woe to you, Bethsaida! For if the mighty works done in you had been done in Tyre and Sidon, they would have repented long ago in sackcloth and ashes.
MATT|11|22|But I tell you, it will be more bearable on the day of judgment for Tyre and Sidon than for you.
MATT|11|23|And you, Capernaum, will you be exalted to heaven? You will be brought down to Hades. For if the mighty works done in you had been done in Sodom, it would have remained until this day.
MATT|11|24|But I tell you that it will be more tolerable on the day of judgment for the land of Sodom than for you."
MATT|11|25|At that time Jesus declared, "I thank you, Father, Lord of heaven and earth, that you have hidden these things from the wise and understanding and revealed them to little children;
MATT|11|26|yes, Father, for such was your gracious will.
MATT|11|27|All things have been handed over to me by my Father, and no one knows the Son except the Father, and no one knows the Father except the Son and anyone to whom the Son chooses to reveal him.
MATT|11|28|Come to me, all who labor and are heavy laden, and I will give you rest.
MATT|11|29|Take my yoke upon you, and learn from me, for I am gentle and lowly in heart, and you will find rest for your souls.
MATT|11|30|For my yoke is easy, and my burden is light."
MATT|12|1|At that time Jesus went through the grainfields on the Sabbath. His disciples were hungry, and they began to pluck heads of grain and to eat.
MATT|12|2|But when the Pharisees saw it, they said to him, "Look, your disciples are doing what is not lawful to do on the Sabbath."
MATT|12|3|He said to them, "Have you not read what David did when he was hungry, and those who were with him:
MATT|12|4|how he entered the house of God and ate the bread of the Presence, which it was not lawful for him to eat nor for those who were with him, but only for the priests?
MATT|12|5|Or have you not read in the Law how on the Sabbath the priests in the temple profane the Sabbath and are guiltless?
MATT|12|6|I tell you, something greater than the temple is here.
MATT|12|7|And if you had known what this means, 'I desire mercy, and not sacrifice,' you would not have condemned the guiltless.
MATT|12|8|For the Son of Man is lord of the Sabbath."
MATT|12|9|He went on from there and entered their synagogue.
MATT|12|10|And a man was there with a withered hand. And they asked him, "Is it lawful to heal on the Sabbath?"- so that they might accuse him.
MATT|12|11|He said to them, "Which one of you who has a sheep, if it falls into a pit on the Sabbath, will not take hold of it and lift it out?
MATT|12|12|Of how much more value is a man than a sheep! So it is lawful to do good on the Sabbath."
MATT|12|13|Then he said to the man, "Stretch out your hand." And the man stretched it out, and it was restored, healthy like the other.
MATT|12|14|But the Pharisees went out and conspired against him, how to destroy him.
MATT|12|15|Jesus, aware of this, withdrew from there. And many followed him, and he healed them all
MATT|12|16|and ordered them not to make him known.
MATT|12|17|This was to fulfill what was spoken by the prophet Isaiah:
MATT|12|18|"Behold, my servant whom I have chosen, my beloved with whom my soul is well pleased. I will put my Spirit upon him, and he will proclaim justice to the Gentiles.
MATT|12|19|He will not quarrel or cry aloud, nor will anyone hear his voice in the streets;
MATT|12|20|a bruised reed he will not break, and a smoldering wick he will not quench, until he brings justice to victory;
MATT|12|21|and in his name the Gentiles will hope."
MATT|12|22|Then a demon-oppressed man who was blind and mute was brought to him, and he healed him, so that the man spoke and saw.
MATT|12|23|And all the people were amazed, and said, "Can this be the Son of David?"
MATT|12|24|But when the Pharisees heard it, they said, "It is only by Beelzebul, the prince of demons, that this man casts out demons."
MATT|12|25|Knowing their thoughts, he said to them, "Every kingdom divided against itself is laid waste, and no city or house divided against itself will stand.
MATT|12|26|And if Satan casts out Satan, he is divided against himself. How then will his kingdom stand?
MATT|12|27|And if I cast out demons by Beelzebul, by whom do your sons cast them out? Therefore they will be your judges.
MATT|12|28|But if it is by the Spirit of God that I cast out demons, then the kingdom of God has come upon you.
MATT|12|29|Or how can someone enter a strong man's house and plunder his goods, unless he first binds the strong man? Then indeed he may plunder his house.
MATT|12|30|Whoever is not with me is against me, and whoever does not gather with me scatters.
MATT|12|31|Therefore I tell you, every sin and blasphemy will be forgiven people, but the blasphemy against the Spirit will not be forgiven.
MATT|12|32|And whoever speaks a word against the Son of Man will be forgiven, but whoever speaks against the Holy Spirit will not be forgiven, either in this age or in the age to come.
MATT|12|33|"Either make the tree good and its fruit good, or make the tree bad and its fruit bad, for the tree is known by its fruit.
MATT|12|34|You brood of vipers! How can you speak good, when you are evil? For out of the abundance of the heart the mouth speaks.
MATT|12|35|The good person out of his good treasure brings forth good, and the evil person out of his evil treasure brings forth evil.
MATT|12|36|I tell you, on the day of judgment people will give account for every careless word they speak,
MATT|12|37|for by your words you will be justified, and by your words you will be condemned."
MATT|12|38|Then some of the scribes and Pharisees answered him, saying, "Teacher, we wish to see a sign from you."
MATT|12|39|But he answered them, "An evil and adulterous generation seeks for a sign, but no sign will be given to it except the sign of the prophet Jonah.
MATT|12|40|For just as Jonah was three days and three nights in the belly of the great fish, so will the Son of Man be three days and three nights in the heart of the earth.
MATT|12|41|The men of Nineveh will rise up at the judgment with this generation and condemn it, for they repented at the preaching of Jonah, and behold, something greater than Jonah is here.
MATT|12|42|The queen of the South will rise up at the judgment with this generation and condemn it, for she came from the ends of the earth to hear the wisdom of Solomon, and behold, something greater than Solomon is here.
MATT|12|43|"When the unclean spirit has gone out of a person, it passes through waterless places seeking rest, but finds none.
MATT|12|44|Then it says, 'I will return to my house from which I came.' And when it comes, it finds the house empty, swept, and put in order.
MATT|12|45|Then it goes and brings with it seven other spirits more evil than itself, and they enter and dwell there, and the last state of that person is worse than the first. So also will it be with this evil generation."
MATT|12|46|While he was still speaking to the people, behold, his mother and his brothers stood outside, asking to speak to him.
MATT|12|47|***
MATT|12|48|But he replied to the man who told him, "Who is my mother, and who are my brothers?"
MATT|12|49|And stretching out his hand toward his disciples, he said, "Here are my mother and my brothers!
MATT|12|50|For whoever does the will of my Father in heaven is my brother and sister and mother."
MATT|13|1|That same day Jesus went out of the house and sat beside the sea.
MATT|13|2|And great crowds gathered about him, so that he got into a boat and sat down. And the whole crowd stood on the beach.
MATT|13|3|And he told them many things in parables, saying: "A sower went out to sow.
MATT|13|4|And as he sowed, some seeds fell along the path, and the birds came and devoured them.
MATT|13|5|Other seeds fell on rocky ground, where they did not have much soil, and immediately they sprang up, since they had no depth of soil,
MATT|13|6|but when the sun rose they were scorched. And since they had no root, they withered away.
MATT|13|7|Other seeds fell among thorns, and the thorns grew up and choked them.
MATT|13|8|Other seeds fell on good soil and produced grain, some a hundredfold, some sixty, some thirty.
MATT|13|9|He who has ears, let him hear."
MATT|13|10|Then the disciples came and said to him, "Why do you speak to them in parables?"
MATT|13|11|And he answered them, "To you it has been given to know the secrets of the kingdom of heaven, but to them it has not been given.
MATT|13|12|For to the one who has, more will be given, and he will have an abundance, but from the one who has not, even what he has will be taken away.
MATT|13|13|This is why I speak to them in parables, because seeing they do not see, and hearing they do not hear, nor do they understand.
MATT|13|14|Indeed, in their case the prophecy of Isaiah is fulfilled that says: "' You will indeed hear but never understand, and you will indeed see but never perceive.
MATT|13|15|For this people's heart has grown dull, and with their ears they can barely hear, and their eyes they have closed, lest they should see with their eyes and hear with their ears and understand with their heart and turn, and I would heal them.'
MATT|13|16|But blessed are your eyes, for they see, and your ears, for they hear.
MATT|13|17|Truly, I say to you, many prophets and righteous people longed to see what you see, and did not see it, and to hear what you hear, and did not hear it.
MATT|13|18|"Hear then the parable of the sower:
MATT|13|19|When anyone hears the word of the kingdom and does not understand it, the evil one comes and snatches away what has been sown in his heart. This is what was sown along the path.
MATT|13|20|As for what was sown on rocky ground, this is the one who hears the word and immediately receives it with joy,
MATT|13|21|yet he has no root in himself, but endures for a while, and when tribulation or persecution arises on account of the word, immediately he falls away.
MATT|13|22|As for what was sown among thorns, this is the one who hears the word, but the cares of the world and the deceitfulness of riches choke the word, and it proves unfruitful.
MATT|13|23|As for what was sown on good soil, this is the one who hears the word and understands it. He indeed bears fruit and yields, in one case a hundredfold, in another sixty, and in another thirty."
MATT|13|24|He put another parable before them, saying, "The kingdom of heaven may be compared to a man who sowed good seed in his field,
MATT|13|25|but while his men were sleeping, his enemy came and sowed weeds among the wheat and went away.
MATT|13|26|So when the plants came up and bore grain, then the weeds appeared also.
MATT|13|27|And the servants of the master of the house came and said to him, 'Master, did you not sow good seed in your field? How then does it have weeds?'
MATT|13|28|He said to them, 'An enemy has done this.' So the servants said to him, 'Then do you want us to go and gather them?'
MATT|13|29|But he said, 'No, lest in gathering the weeds you root up the wheat along with them.
MATT|13|30|Let both grow together until the harvest, and at harvest time I will tell the reapers, Gather the weeds first and bind them in bundles to be burned, but gather the wheat into my barn.'"
MATT|13|31|He put another parable before them, saying, "The kingdom of heaven is like a grain of mustard seed that a man took and sowed in his field.
MATT|13|32|It is the smallest of all seeds, but when it has grown it is larger than all the garden plants and becomes a tree, so that the birds of the air come and make nests in its branches."
MATT|13|33|He told them another parable. "The kingdom of heaven is like leaven that a woman took and hid in three measures of flour, till it was all leavened."
MATT|13|34|All these things Jesus said to the crowds in parables; indeed, he said nothing to them without a parable.
MATT|13|35|This was to fulfill what was spoken by the prophet: "I will open my mouth in parables; I will utter what has been hidden since the foundation of the world."
MATT|13|36|Then he left the crowds and went into the house. And his disciples came to him, saying, "Explain to us the parable of the weeds of the field."
MATT|13|37|He answered, "The one who sows the good seed is the Son of Man.
MATT|13|38|The field is the world, and the good seed is the children of the kingdom. The weeds are the sons of the evil one,
MATT|13|39|and the enemy who sowed them is the devil. The harvest is the close of the age, and the reapers are angels.
MATT|13|40|Just as the weeds are gathered and burned with fire, so will it be at the close of the age.
MATT|13|41|The Son of Man will send his angels, and they will gather out of his kingdom all causes of sin and all law-breakers,
MATT|13|42|and throw them into the fiery furnace. In that place there will be weeping and gnashing of teeth.
MATT|13|43|Then the righteous will shine like the sun in the kingdom of their Father. He who has ears, let him hear.
MATT|13|44|"The kingdom of heaven is like treasure hidden in a field, which a man found and covered up. Then in his joy he goes and sells all that he has and buys that field.
MATT|13|45|"Again, the kingdom of heaven is like a merchant in search of fine pearls,
MATT|13|46|who, on finding one pearl of great value, went and sold all that he had and bought it.
MATT|13|47|"Again, the kingdom of heaven is like a net that was thrown into the sea and gathered fish of every kind.
MATT|13|48|When it was full, men drew it ashore and sat down and sorted the good into containers but threw away the bad.
MATT|13|49|So it will be at the close of the age. The angels will come out and separate the evil from the righteous
MATT|13|50|and throw them into the fiery furnace. In that place there will be weeping and gnashing of teeth.
MATT|13|51|"Have you understood all these things?" They said to him, "Yes."
MATT|13|52|And he said to them, "Therefore every scribe who has been trained for the kingdom of heaven is like a master of a house, who brings out of his treasure what is new and what is old."
MATT|13|53|And when Jesus had finished these parables, he went away from there,
MATT|13|54|and coming to his hometown he taught them in their synagogue, so that they were astonished, and said, "Where did this man get this wisdom and these mighty works?
MATT|13|55|Is not this the carpenter's son? Is not his mother called Mary? And are not his brothers James and Joseph and Simon and Judas?
MATT|13|56|And are not all his sisters with us? Where then did this man get all these things?"
MATT|13|57|And they took offense at him. But Jesus said to them, "A prophet is not without honor except in his hometown and in his own household."
MATT|13|58|And he did not do many mighty works there, because of their unbelief.
MATT|14|1|At that time Herod the tetrarch heard about the fame of Jesus,
MATT|14|2|and he said to his servants, "This is John the Baptist. He has been raised from the dead; that is why these miraculous powers are at work in him."
MATT|14|3|For Herod had seized John and bound him and put him in prison for the sake of Herodias, his brother Philip's wife,
MATT|14|4|because John had been saying to him, "It is not lawful for you to have her."
MATT|14|5|And though he wanted to put him to death, he feared the people, because they held him to be a prophet.
MATT|14|6|But when Herod's birthday came, the daughter of Herodias danced before the company and pleased Herod,
MATT|14|7|so that he promised with an oath to give her whatever she might ask.
MATT|14|8|Prompted by her mother, she said, "Give me the head of John the Baptist here on a platter."
MATT|14|9|And the king was sorry, but because of his oaths and his guests he commanded it to be given.
MATT|14|10|He sent and had John beheaded in the prison,
MATT|14|11|and his head was brought on a platter and given to the girl, and she brought it to her mother.
MATT|14|12|And his disciples came and took the body and buried it, and they went and told Jesus.
MATT|14|13|Now when Jesus heard this, he withdrew from there in a boat to a desolate place by himself. But when the crowds heard it, they followed him on foot from the towns.
MATT|14|14|When he went ashore he saw a great crowd, and he had compassion on them and healed their sick.
MATT|14|15|Now when it was evening, the disciples came to him and said, "This is a desolate place, and the day is now over; send the crowds away to go into the villages and buy food for themselves."
MATT|14|16|But Jesus said, "They need not go away; you give them something to eat."
MATT|14|17|They said to him, "We have only five loaves here and two fish."
MATT|14|18|And he said, "Bring them here to me."
MATT|14|19|Then he ordered the crowds to sit down on the grass, and taking the five loaves and the two fish, he looked up to heaven and said a blessing. Then he broke the loaves and gave them to the disciples, and the disciples gave them to the crowds.
MATT|14|20|And they all ate and were satisfied. And they took up twelve baskets full of the broken pieces left over.
MATT|14|21|And those who ate were about five thousand men, besides women and children.
MATT|14|22|Immediately he made the disciples get into the boat and go before him to the other side, while he dismissed the crowds.
MATT|14|23|And after he had dismissed the crowds, he went up on the mountain by himself to pray. When evening came, he was there alone,
MATT|14|24|but the boat by this time was a long way from the land, beaten by the waves, for the wind was against them.
MATT|14|25|And in the fourth watch of the night he came to them, walking on the sea.
MATT|14|26|But when the disciples saw him walking on the sea, they were terrified, and said, "It is a ghost!" and they cried out in fear.
MATT|14|27|But immediately Jesus spoke to them, saying, "Take heart; it is I. Do not be afraid."
MATT|14|28|And Peter answered him, "Lord, if it is you, command me to come to you on the water."
MATT|14|29|He said, "Come." So Peter got out of the boat and walked on the water and came to Jesus.
MATT|14|30|But when he saw the wind, he was afraid, and beginning to sink he cried out, "Lord, save me."
MATT|14|31|Jesus immediately reached out his hand and took hold of him, saying to him, "O you of little faith, why did you doubt?"
MATT|14|32|And when they got into the boat, the wind ceased.
MATT|14|33|And those in the boat worshiped him, saying, "Truly you are the Son of God."
MATT|14|34|And when they had crossed over, they came to land at Gennesaret.
MATT|14|35|And when the men of that place recognized him, they sent around to all that region and brought to him all who were sick
MATT|14|36|and implored him that they might only touch the fringe of his garment. And as many as touched it were made well.
MATT|15|1|Then Pharisees and scribes came to Jesus from Jerusalem and said,
MATT|15|2|"Why do your disciples break the tradition of the elders? For they do not wash their hands when they eat."
MATT|15|3|He answered them, "And why do you break the commandment of God for the sake of your tradition?
MATT|15|4|For God commanded, 'Honor your father and your mother,' and, 'Whoever reviles father or mother must surely die.'
MATT|15|5|But you say, 'If anyone tells his father or his mother, What you would have gained from me is given to God,
MATT|15|6|he need not honor his father.' So for the sake of your tradition you have made void the word of God.
MATT|15|7|You hypocrites! Well did Isaiah prophesy of you, when he said:
MATT|15|8|"'This people honors me with their lips, but their heart is far from me;
MATT|15|9|in vain do they worship me, teaching as doctrines the commandments of men.'"
MATT|15|10|And he called the people to him and said to them, "Hear and understand:
MATT|15|11|it is not what goes into the mouth that defiles a person, but what comes out of the mouth; this defiles a person."
MATT|15|12|Then the disciples came and said to him, "Do you know that the Pharisees were offended when they heard this saying?"
MATT|15|13|He answered, "Every plant that my heavenly Father has not planted will be rooted up.
MATT|15|14|Let them alone; they are blind guides. And if the blind lead the blind, both will fall into a pit."
MATT|15|15|But Peter said to him, "Explain the parable to us."
MATT|15|16|And he said, "Are you also still without understanding?
MATT|15|17|Do you not see that whatever goes into the mouth passes into the stomach and is expelled?
MATT|15|18|But what comes out of the mouth proceeds from the heart, and this defiles a person.
MATT|15|19|For out of the heart come evil thoughts, murder, adultery, sexual immorality, theft, false witness, slander.
MATT|15|20|These are what defile a person. But to eat with unwashed hands does not defile anyone."
MATT|15|21|And Jesus went away from there and withdrew to the district of Tyre and Sidon.
MATT|15|22|And behold, a Canaanite woman from that region came out and was crying, "Have mercy on me, O Lord, Son of David; my daughter is severely oppressed by a demon."
MATT|15|23|But he did not answer her a word. And his disciples came and begged him, saying, "Send her away, for she is crying out after us."
MATT|15|24|He answered, "I was sent only to the lost sheep of the house of Israel."
MATT|15|25|But she came and knelt before him, saying, "Lord, help me."
MATT|15|26|And he answered, "It is not right to take the children's bread and throw it to the dogs."
MATT|15|27|She said, "Yes, Lord, yet even the dogs eat the crumbs that fall from their masters' table."
MATT|15|28|Then Jesus answered her, "O woman, great is your faith! Be it done for you as you desire." And her daughter was healed instantly.
MATT|15|29|Jesus went on from there and walked beside the Sea of Galilee. And he went up on the mountain and sat down there.
MATT|15|30|And great crowds came to him, bringing with them the lame, the blind, the crippled, the mute, and many others, and they put them at his feet, and he healed them,
MATT|15|31|so that the crowd wondered, when they saw the mute speaking, the crippled healthy, the lame walking, and the blind seeing. And they glorified the God of Israel.
MATT|15|32|Then Jesus called his disciples to him and said, "I have compassion on the crowd because they have been with me now three days and have nothing to eat. And I am unwilling to send them away hungry, lest they faint on the way."
MATT|15|33|And the disciples said to him, "Where are we to get enough bread in such a desolate place to feed so great a crowd?"
MATT|15|34|And Jesus said to them, "How many loaves do you have?" They said, "Seven, and a few small fish."
MATT|15|35|And directing the crowd to sit down on the ground,
MATT|15|36|he took the seven loaves and the fish, and having given thanks he broke them and gave them to the disciples, and the disciples gave them to the crowds.
MATT|15|37|And they all ate and were satisfied. And they took up seven baskets full of the broken pieces left over.
MATT|15|38|Those who ate were four thousand men, besides women and children.
MATT|15|39|And after sending away the crowds, he got into the boat and went to the region of Magadan.
MATT|16|1|And the Pharisees and Sadducees came, and to test him they asked him to show them a sign from heaven.
MATT|16|2|He answered them, "When it is evening, you say, 'It will be fair weather, for the sky is red.'
MATT|16|3|And in the morning, 'It will be stormy today, for the sky is red and threatening.' You know how to interpret the appearance of the sky, but you cannot interpret the signs of the times.
MATT|16|4|An evil and adulterous generation seeks for a sign, but no sign will be given to it except the sign of Jonah." So he left them and departed.
MATT|16|5|When the disciples reached the other side, they had forgotten to bring any bread.
MATT|16|6|Jesus said to them, "Watch and beware of the leaven of the Pharisees and Sadducees."
MATT|16|7|And they began discussing it among themselves, saying, "We brought no bread."
MATT|16|8|But Jesus, aware of this, said, "O you of little faith, why are you discussing among yourselves the fact that you have no bread?
MATT|16|9|Do you not yet perceive? Do you not remember the five loaves for the five thousand, and how many baskets you gathered?
MATT|16|10|Or the seven loaves for the four thousand, and how many baskets you gathered?
MATT|16|11|How is it that you fail to understand that I did not speak about bread? Beware of the leaven of the Pharisees and Sadducees."
MATT|16|12|Then they understood that he did not tell them to beware of the leaven of bread, but of the teaching of the Pharisees and Sadducees.
MATT|16|13|Now when Jesus came into the district of Caesarea Philippi, he asked his disciples, "Who do people say that the Son of Man is?"
MATT|16|14|And they said, "Some say John the Baptist, others say Elijah, and others Jeremiah or one of the prophets."
MATT|16|15|He said to them, "But who do you say that I am?"
MATT|16|16|Simon Peter replied, "You are the Christ, the Son of the living God."
MATT|16|17|And Jesus answered him, "Blessed are you, Simon Bar-Jonah! For flesh and blood has not revealed this to you, but my Father who is in heaven.
MATT|16|18|And I tell you, you are Peter, and on this rock I will build my church, and the gates of hell shall not prevail against it.
MATT|16|19|I will give you the keys of the kingdom of heaven, and whatever you bind on earth shall be bound in heaven, and whatever you loose on earth shall be loosed in heaven."
MATT|16|20|Then he strictly charged the disciples to tell no one that he was the Christ.
MATT|16|21|From that time Jesus began to show his disciples that he must go to Jerusalem and suffer many things from the elders and chief priests and scribes, and be killed, and on the third day be raised.
MATT|16|22|And Peter took him aside and began to rebuke him, saying, "Far be it from you, Lord! This shall never happen to you."
MATT|16|23|But he turned and said to Peter, "Get behind me, Satan! You are a hindrance to me. For you are not setting your mind on the things of God, but on the things of man."
MATT|16|24|Then Jesus told his disciples, "If anyone would come after me, let him deny himself and take up his cross and follow me.
MATT|16|25|For whoever would save his life will lose it, but whoever loses his life for my sake will find it.
MATT|16|26|For what will it profit a man if he gains the whole world and forfeits his life? Or what shall a man give in return for his life?
MATT|16|27|For the Son of Man is going to come with his angels in the glory of his Father, and then he will repay each person according to what he has done.
MATT|16|28|Truly, I say to you, there are some standing here who will not taste death until they see the Son of Man coming in his kingdom."
MATT|17|1|And after six days Jesus took with him Peter and James, and John his brother, and led them up a high mountain by themselves.
MATT|17|2|And he was transfigured before them, and his face shone like the sun, and his clothes became white as light.
MATT|17|3|And behold, there appeared to them Moses and Elijah, talking with him.
MATT|17|4|And Peter said to Jesus, "Lord, it is good that we are here. If you wish, I will make three tents here, one for you and one for Moses and one for Elijah."
MATT|17|5|He was still speaking when, behold, a bright cloud overshadowed them, and a voice from the cloud said, "This is my beloved Son, with whom I am well pleased; listen to him."
MATT|17|6|When the disciples heard this, they fell on their faces and were terrified.
MATT|17|7|But Jesus came and touched them, saying, "Rise, and have no fear."
MATT|17|8|And when they lifted up their eyes, they saw no one but Jesus only.
MATT|17|9|And as they were coming down the mountain, Jesus commanded them, "Tell no one the vision, until the Son of Man is raised from the dead."
MATT|17|10|And the disciples asked him, "Then why do the scribes say that first Elijah must come?"
MATT|17|11|He answered, "Elijah does come, and he will restore all things.
MATT|17|12|But I tell you that Elijah has already come, and they did not recognize him, but did to him whatever they pleased. So also the Son of Man will certainly suffer at their hands."
MATT|17|13|Then the disciples understood that he was speaking to them of John the Baptist.
MATT|17|14|And when they came to the crowd, a man came up to him and, kneeling before him,
MATT|17|15|said, "Lord, have mercy on my son, for he is an epileptic and he suffers terribly. For often he falls into the fire, and often into the water.
MATT|17|16|And I brought him to your disciples, and they could not heal him."
MATT|17|17|And Jesus answered, "O faithless and twisted generation, how long am I to be with you? How long am I to bear with you? Bring him here to me."
MATT|17|18|And Jesus rebuked him, and the demon came out of him, and the boy was healed instantly.
MATT|17|19|Then the disciples came to Jesus privately and said, "Why could we not cast it out?"
MATT|17|20|He said to them, "Because of your little faith. For truly, I say to you, if you have faith like a grain of mustard seed, you will say to this mountain, 'Move from here to there,' and it will move, and nothing will be impossible for you."
MATT|17|21|***
MATT|17|22|As they were gathering in Galilee, Jesus said to them, "The Son of Man is about to be delivered into the hands of men,
MATT|17|23|and they will kill him, and he will be raised on the third day." And they were greatly distressed.
MATT|17|24|When they came to Capernaum, the collectors of the half-shekel tax went up to Peter and said, "Does your teacher not pay the tax?"
MATT|17|25|He said, "Yes." And when he came into the house, Jesus spoke to him first, saying, "What do you think, Simon? From whom do kings of the earth take toll or tax? From their sons or from others?"
MATT|17|26|And when he said, "From others," Jesus said to him, "Then the sons are free.
MATT|17|27|However, not to give offense to them, go to the sea and cast a hook and take the first fish that comes up, and when you open its mouth you will find a shekel. Take that and give it to them for me and for yourself."
MATT|18|1|At that time the disciples came to Jesus, saying, "Who is the greatest in the kingdom of heaven?"
MATT|18|2|And calling to him a child, he put him in the midst of them
MATT|18|3|and said, "Truly, I say to you, unless you turn and become like children, you will never enter the kingdom of heaven.
MATT|18|4|Whoever humbles himself like this child is the greatest in the kingdom of heaven.
MATT|18|5|"Whoever receives one such child in my name receives me,
MATT|18|6|but whoever causes one of these little ones who believe in me to sin, it would be better for him to have a great millstone fastened around his neck and to be drowned in the depth of the sea.
MATT|18|7|"Woe to the world for temptations to sin! For it is necessary that temptations come, but woe to the one by whom the temptation comes!
MATT|18|8|And if your hand or your foot causes you to sin, cut it off and throw it away. It is better for you to enter life crippled or lame than with two hands or two feet to be thrown into the eternal fire.
MATT|18|9|And if your eye causes you to sin, tear it out and throw it away. It is better for you to enter life with one eye than with two eyes to be thrown into the hell of fire.
MATT|18|10|"See that you do not despise one of these little ones. For I tell you that in heaven their angels always see the face of my Father who is in heaven.
MATT|18|11|***
MATT|18|12|What do you think? If a man has a hundred sheep and one of them has gone astray, does he not leave the ninety-nine on the mountains and go in search of the one that went astray?
MATT|18|13|And if he finds it, truly, I say to you, he rejoices over it more than over the ninety-nine that never went astray.
MATT|18|14|So it is not the will of my Father who is in heaven that one of these little ones should perish.
MATT|18|15|"If your brother sins against you, go and tell him his fault, between you and him alone. If he listens to you, you have gained your brother.
MATT|18|16|But if he does not listen, take one or two others along with you, that every charge may be established by the evidence of two or three witnesses.
MATT|18|17|If he refuses to listen to them, tell it to the church. And if he refuses to listen even to the church, let him be to you as a Gentile and a tax collector.
MATT|18|18|Truly, I say to you, whatever you bind on earth shall be bound in heaven, and whatever you loose on earth shall be loosed in heaven.
MATT|18|19|Again I say to you, if two of you agree on earth about anything they ask, it will be done for them by my Father in heaven.
MATT|18|20|For where two or three are gathered in my name, there am I among them."
MATT|18|21|Then Peter came up and said to him, "Lord, how often will my brother sin against me, and I forgive him? As many as seven times?"
MATT|18|22|Jesus said to him, "I do not say to you seven times, but seventy times seven.
MATT|18|23|"Therefore the kingdom of heaven may be compared to a king who wished to settle accounts with his servants.
MATT|18|24|When he began to settle, one was brought to him who owed him ten thousand talents.
MATT|18|25|And since he could not pay, his master ordered him to be sold, with his wife and children and all that he had, and payment to be made.
MATT|18|26|So the servant fell on his knees, imploring him, 'Have patience with me, and I will pay you everything.'
MATT|18|27|And out of pity for him, the master of that servant released him and forgave him the debt.
MATT|18|28|But when that same servant went out, he found one of his fellow servants who owed him a hundred denarii, and seizing him, he began to choke him, saying, 'Pay what you owe.'
MATT|18|29|So his fellow servant fell down and pleaded with him, 'Have patience with me, and I will pay you.'
MATT|18|30|He refused and went and put him in prison until he should pay the debt.
MATT|18|31|When his fellow servants saw what had taken place, they were greatly distressed, and they went and reported to their master all that had taken place.
MATT|18|32|Then his master summoned him and said to him, 'You wicked servant! I forgave you all that debt because you pleaded with me.
MATT|18|33|And should not you have had mercy on your fellow servant, as I had mercy on you?'
MATT|18|34|And in anger his master delivered him to the jailers, until he should pay all his debt.
MATT|18|35|So also my heavenly Father will do to every one of you, if you do not forgive your brother from your heart."
MATT|19|1|Now when Jesus had finished these sayings, he went away from Galilee and entered the region of Judea beyond the Jordan.
MATT|19|2|And large crowds followed him, and he healed them there.
MATT|19|3|And Pharisees came up to him and tested him by asking, "Is it lawful to divorce one's wife for any cause?"
MATT|19|4|He answered, "Have you not read that he who created them from the beginning made them male and female,
MATT|19|5|and said, 'Therefore a man shall leave his father and his mother and hold fast to his wife, and they shall become one flesh'?
MATT|19|6|So they are no longer two but one flesh. What therefore God has joined together, let not man separate."
MATT|19|7|They said to him, "Why then did Moses command one to give a certificate of divorce and to send her away?"
MATT|19|8|He said to them, "Because of your hardness of heart Moses allowed you to divorce your wives, but from the beginning it was not so.
MATT|19|9|And I say to you: whoever divorces his wife, except for sexual immorality, and marries another, commits adultery."
MATT|19|10|The disciples said to him, "If such is the case of a man with his wife, it is better not to marry."
MATT|19|11|But he said to them, "Not everyone can receive this saying, but only those to whom it is given.
MATT|19|12|For there are eunuchs who have been so from birth, and there are eunuchs who have been made eunuchs by men, and there are eunuchs who have made themselves eunuchs for the sake of the kingdom of heaven. Let the one who is able to receive this receive it."
MATT|19|13|Then children were brought to him that he might lay his hands on them and pray. The disciples rebuked the people,
MATT|19|14|but Jesus said, "Let the little children come to me and do not hinder them, for to such belongs the kingdom of heaven."
MATT|19|15|And he laid his hands on them and went away.
MATT|19|16|And behold, a man came up to him, saying, "Teacher, what good deed must I do to have eternal life?"
MATT|19|17|And he said to him, "Why do you ask me about what is good? There is only one who is good. If you would enter life, keep the commandments."
MATT|19|18|He said to him, "Which ones?" And Jesus said, "You shall not murder, You shall not commit adultery, You shall not steal, You shall not bear false witness,
MATT|19|19|Honor your father and mother, and, You shall love your neighbor as yourself."
MATT|19|20|The young man said to him, "All these I have kept. What do I still lack?"
MATT|19|21|Jesus said to him, "If you would be perfect, go, sell what you possess and give to the poor, and you will have treasure in heaven; and come, follow me."
MATT|19|22|When the young man heard this he went away sorrowful, for he had great possessions.
MATT|19|23|And Jesus said to his disciples, "Truly, I say to you, only with difficulty will a rich person enter the kingdom of heaven.
MATT|19|24|Again I tell you, it is easier for a camel to go through the eye of a needle than for a rich person to enter the kingdom of God."
MATT|19|25|When the disciples heard this, they were greatly astonished, saying, "Who then can be saved?"
MATT|19|26|But Jesus looked at them and said, "With man this is impossible, but with God all things are possible."
MATT|19|27|Then Peter said in reply, "See, we have left everything and followed you. What then will we have?"
MATT|19|28|Jesus said to them, "Truly, I say to you, in the new world, when the Son of Man will sit on his glorious throne, you who have followed me will also sit on twelve thrones, judging the twelve tribes of Israel.
MATT|19|29|And everyone who has left houses or brothers or sisters or father or mother or children or lands, for my name's sake, will receive a hundredfold and will inherit eternal life.
MATT|19|30|But many who are first will be last, and the last first.
MATT|20|1|"For the kingdom of heaven is like a master of a house who went out early in the morning to hire laborers for his vineyard.
MATT|20|2|After agreeing with the laborers for a denarius a day, he sent them into his vineyard.
MATT|20|3|And going out about the third hour he saw others standing idle in the marketplace,
MATT|20|4|and to them he said, 'You go into the vineyard too, and whatever is right I will give you.'
MATT|20|5|So they went. Going out again about the sixth hour and the ninth hour, he did the same.
MATT|20|6|And about the eleventh hour he went out and found others standing. And he said to them, 'Why do you stand here idle all day?'
MATT|20|7|They said to him, 'Because no one has hired us.' He said to them, 'You go into the vineyard too.'
MATT|20|8|And when evening came, the owner of the vineyard said to his foreman, 'Call the laborers and pay them their wages, beginning with the last, up to the first.'
MATT|20|9|And when those hired about the eleventh hour came, each of them received a denarius.
MATT|20|10|Now when those hired first came, they thought they would receive more, but each of them also received a denarius.
MATT|20|11|And on receiving it they grumbled at the master of the house,
MATT|20|12|saying, 'These last worked only one hour, and you have made them equal to us who have borne the burden of the day and the scorching heat.'
MATT|20|13|But he replied to one of them, 'Friend, I am doing you no wrong. Did you not agree with me for a denarius?
MATT|20|14|Take what belongs to you and go. I choose to give to this last worker as I give to you.
MATT|20|15|Am I not allowed to do what I choose with what belongs to me? Or do you begrudge my generosity?'
MATT|20|16|So the last will be first, and the first last."
MATT|20|17|And as Jesus was going up to Jerusalem, he took the twelve disciples aside, and on the way he said to them,
MATT|20|18|"See, we are going up to Jerusalem. And the Son of Man will be delivered over to the chief priests and scribes, and they will condemn him to death
MATT|20|19|and deliver him over to the Gentiles to be mocked and flogged and crucified, and he will be raised on the third day."
MATT|20|20|Then the mother of the sons of Zebedee came up to him with her sons, and kneeling before him she asked him for something.
MATT|20|21|And he said to her, "What do you want?" She said to him, "Say that these two sons of mine are to sit, one at your right hand and one at your left, in your kingdom."
MATT|20|22|Jesus answered, "You do not know what you are asking. Are you able to drink the cup that I am to drink?" They said to him, "We are able."
MATT|20|23|He said to them, "You will drink my cup, but to sit at my right hand and at my left is not mine to grant, but it is for those for whom it has been prepared by my Father."
MATT|20|24|And when the ten heard it, they were indignant at the two brothers.
MATT|20|25|But Jesus called them to him and said, "You know that the rulers of the Gentiles lord it over them, and their great ones exercise authority over them.
MATT|20|26|It shall not be so among you. But whoever would be great among you must be your servant,
MATT|20|27|and whoever would be first among you must be your slave,
MATT|20|28|even as the Son of Man came not to be served but to serve, and to give his life as a ransom for many."
MATT|20|29|And as they went out of Jericho, a great crowd followed him.
MATT|20|30|And behold, there were two blind men sitting by the roadside, and when they heard that Jesus was passing by, they cried out, "Lord, have mercy on us, Son of David!"
MATT|20|31|The crowd rebuked them, telling them to be silent, but they cried out all the more, "Lord, have mercy on us, Son of David!"
MATT|20|32|And stopping, Jesus called them and said, "What do you want me to do for you?"
MATT|20|33|They said to him, "Lord, let our eyes be opened."
MATT|20|34|And Jesus in pity touched their eyes, and immediately they recovered their sight and followed him.
MATT|21|1|Now when they drew near to Jerusalem and came to Bethphage, to the Mount of Olives, then Jesus sent two disciples,
MATT|21|2|saying to them, "Go into the village in front of you, and immediately you will find a donkey tied, and a colt with her. Untie them and bring them to me.
MATT|21|3|If anyone says anything to you, you shall say, 'The Lord needs them,' and he will send them at once."
MATT|21|4|This took place to fulfill what was spoken by the prophet, saying,
MATT|21|5|"Say to the daughter of Zion, 'Behold, your king is coming to you, humble, and mounted on a donkey, and on a colt, the foal of a beast of burden.'"
MATT|21|6|The disciples went and did as Jesus had directed them.
MATT|21|7|They brought the donkey and the colt and put on them their cloaks, and he sat on them.
MATT|21|8|Most of the crowd spread their cloaks on the road, and others cut branches from the trees and spread them on the road.
MATT|21|9|And the crowds that went before him and that followed him were shouting, "Hosanna to the Son of David! Blessed is he who comes in the name of the Lord! Hosanna in the highest!"
MATT|21|10|And when he entered Jerusalem, the whole city was stirred up, saying, "Who is this?"
MATT|21|11|And the crowds said, "This is the prophet Jesus, from Nazareth of Galilee."
MATT|21|12|And Jesus entered the temple and drove out all who sold and bought in the temple, and he overturned the tables of the money-changers and the seats of those who sold pigeons.
MATT|21|13|He said to them, "It is written, 'My house shall be called a house of prayer,' but you make it a den of robbers."
MATT|21|14|And the blind and the lame came to him in the temple, and he healed them.
MATT|21|15|But when the chief priests and the scribes saw the wonderful things that he did, and the children crying out in the temple, "Hosanna to the Son of David!" they were indignant,
MATT|21|16|and they said to him, "Do you hear what these are saying?" And Jesus said to them, "Yes; have you never read, "' Out of the mouth of infants and nursing babies you have prepared praise'?"
MATT|21|17|And leaving them, he went out of the city to Bethany and lodged there.
MATT|21|18|In the morning, as he was returning to the city, he became hungry.
MATT|21|19|And seeing a fig tree by the wayside, he went to it and found nothing on it but only leaves. And he said to it, "May no fruit ever come from you again!" And the fig tree withered at once.
MATT|21|20|When the disciples saw it, they marveled, saying, "How did the fig tree wither at once?"
MATT|21|21|And Jesus answered them, "Truly, I say to you, if you have faith and do not doubt, you will not only do what has been done to the fig tree, but even if you say to this mountain, 'Be taken up and thrown into the sea,' it will happen.
MATT|21|22|And whatever you ask in prayer, you will receive, if you have faith."
MATT|21|23|And when he entered the temple, the chief priests and the elders of the people came up to him as he was teaching, and said, "By what authority are you doing these things, and who gave you this authority?"
MATT|21|24|Jesus answered them, "I also will ask you one question, and if you tell me the answer, then I also will tell you by what authority I do these things.
MATT|21|25|The baptism of John, from where did it come? From heaven or from man?" And they discussed it among themselves, saying, "If we say, 'From heaven,' he will say to us, 'Why then did you not believe him?'
MATT|21|26|But if we say, 'From man,' we are afraid of the crowd, for they all hold that John was a prophet."
MATT|21|27|So they answered Jesus, "We do not know." And he said to them, "Neither will I tell you by what authority I do these things.
MATT|21|28|"What do you think? A man had two sons. And he went to the first and said, 'Son, go and work in the vineyard today.'
MATT|21|29|And he answered, 'I will not,' but afterward he changed his mind and went.
MATT|21|30|And he went to the other son and said the same. And he answered, 'I go, sir,' but did not go.
MATT|21|31|Which of the two did the will of his father?" They said, "The first." Jesus said to them, "Truly, I say to you, the tax collectors and the prostitutes go into the kingdom of God before you.
MATT|21|32|For John came to you in the way of righteousness, and you did not believe him, but the tax collectors and the prostitutes believed him. And even when you saw it, you did not afterward change your minds and believe him.
MATT|21|33|"Hear another parable. There was a master of a house who planted a vineyard and put a fence around it and dug a winepress in it and built a tower and leased it to tenants, and went into another country.
MATT|21|34|When the season for fruit drew near, he sent his servants to the tenants to get his fruit.
MATT|21|35|And the tenants took his servants and beat one, killed another, and stoned another.
MATT|21|36|Again he sent other servants, more than the first. And they did the same to them.
MATT|21|37|Finally he sent his son to them, saying, 'They will respect my son.'
MATT|21|38|But when the tenants saw the son, they said to themselves, 'This is the heir. Come, let us kill him and have his inheritance.'
MATT|21|39|And they took him and threw him out of the vineyard and killed him.
MATT|21|40|When therefore the owner of the vineyard comes, what will he do to those tenants?"
MATT|21|41|They said to him, "He will put those wretches to a miserable death and let out the vineyard to other tenants who will give him the fruits in their seasons."
MATT|21|42|Jesus said to them, "Have you never read in the Scriptures: "' The stone that the builders rejected has become the cornerstone; this was the Lord's doing, and it is marvelous in our eyes'?
MATT|21|43|Therefore I tell you, the kingdom of God will be taken away from you and given to a people producing its fruits.
MATT|21|44|And the one who falls on this stone will be broken to pieces; and when it falls on anyone, it will crush him."
MATT|21|45|When the chief priests and the Pharisees heard his parables, they perceived that he was speaking about them.
MATT|21|46|And although they were seeking to arrest him, they feared the crowds, because they held him to be a prophet.
MATT|22|1|And again Jesus spoke to them in parables, saying,
MATT|22|2|"The kingdom of heaven may be compared to a king who gave a wedding feast for his son,
MATT|22|3|and sent his servants to call those who were invited to the wedding feast, but they would not come.
MATT|22|4|Again he sent other servants, saying, 'Tell those who are invited, See, I have prepared my dinner, my oxen and my fat calves have been slaughtered, and everything is ready. Come to the wedding feast.'
MATT|22|5|But they paid no attention and went off, one to his farm, another to his business,
MATT|22|6|while the rest seized his servants, treated them shamefully, and killed them.
MATT|22|7|The king was angry, and he sent his troops and destroyed those murderers and burned their city.
MATT|22|8|Then he said to his servants, 'The wedding feast is ready, but those invited were not worthy.
MATT|22|9|Go therefore to the main roads and invite to the wedding feast as many as you find.'
MATT|22|10|And those servants went out into the roads and gathered all whom they found, both bad and good. So the wedding hall was filled with guests.
MATT|22|11|"But when the king came in to look at the guests, he saw there a man who had no wedding garment.
MATT|22|12|And he said to him, 'Friend, how did you get in here without a wedding garment?' And he was speechless.
MATT|22|13|Then the king said to the attendants, 'Bind him hand and foot and cast him into the outer darkness. In that place there will be weeping and gnashing of teeth.'
MATT|22|14|For many are called, but few are chosen."
MATT|22|15|Then the Pharisees went and plotted how to entangle him in his talk.
MATT|22|16|And they sent their disciples to him, along with the Herodians, saying, "Teacher, we know that you are true and teach the way of God truthfully, and you do not care about anyone's opinion, for you are not swayed by appearances.
MATT|22|17|Tell us, then, what you think. Is it lawful to pay taxes to Caesar, or not?"
MATT|22|18|But Jesus, aware of their malice, said, "Why put me to the test, you hypocrites?
MATT|22|19|Show me the coin for the tax." And they brought him a denarius.
MATT|22|20|And Jesus said to them, "Whose likeness and inscription is this?"
MATT|22|21|They said, "Caesar's." Then he said to them, "Therefore render to Caesar the things that are Caesar's, and to God the things that are God's."
MATT|22|22|When they heard it, they marveled. And they left him and went away.
MATT|22|23|The same day Sadducees came to him, who say that there is no resurrection, and they asked him a question,
MATT|22|24|saying, "Teacher, Moses said, 'If a man dies having no children, his brother must marry the widow and raise up children for his brother.'
MATT|22|25|Now there were seven brothers among us. The first married and died, and having no children left his wife to his brother.
MATT|22|26|So too the second and third, down to the seventh.
MATT|22|27|After them all, the woman died.
MATT|22|28|In the resurrection, therefore, of the seven, whose wife will she be? For they all had her."
MATT|22|29|But Jesus answered them, "You are wrong, because you know neither the Scriptures nor the power of God.
MATT|22|30|For in the resurrection they neither marry nor are given in marriage, but are like angels in heaven.
MATT|22|31|And as for the resurrection of the dead, have you not read what was said to you by God:
MATT|22|32|'I am the God of Abraham, and the God of Isaac, and the God of Jacob'? He is not God of the dead, but of the living."
MATT|22|33|And when the crowd heard it, they were astonished at his teaching.
MATT|22|34|But when the Pharisees heard that he had silenced the Sadducees, they gathered together.
MATT|22|35|And one of them, a lawyer, asked him a question to test him.
MATT|22|36|"Teacher, which is the great commandment in the Law?"
MATT|22|37|And he said to him, "You shall love the Lord your God with all your heart and with all your soul and with all your mind.
MATT|22|38|This is the great and first commandment.
MATT|22|39|And a second is like it: You shall love your neighbor as yourself.
MATT|22|40|On these two commandments depend all the Law and the Prophets."
MATT|22|41|Now while the Pharisees were gathered together, Jesus asked them a question,
MATT|22|42|saying, "What do you think about the Christ? Whose son is he?" They said to him, "The son of David."
MATT|22|43|He said to them, "How is it then that David, in the Spirit, calls him Lord, saying,
MATT|22|44|"'The Lord said to my Lord, Sit at my right hand, until I put your enemies under your feet'?
MATT|22|45|If then David calls him Lord, how is he his son?"
MATT|22|46|And no one was able to answer him a word, nor from that day did anyone dare to ask him any more questions.
MATT|23|1|Then Jesus said to the crowds and to his disciples,
MATT|23|2|"The scribes and the Pharisees sit on Moses' seat,
MATT|23|3|so practice and observe whatever they tell you- but not what they do. For they preach, but do not practice.
MATT|23|4|They tie up heavy burdens, hard to bear, and lay them on people's shoulders, but they themselves are not willing to move them with their finger.
MATT|23|5|They do all their deeds to be seen by others. For they make their phylacteries broad and their fringes long,
MATT|23|6|and they love the place of honor at feasts and the best seats in the synagogues
MATT|23|7|and greetings in the marketplaces and being called rabbi by others.
MATT|23|8|But you are not to be called rabbi, for you have one teacher, and you are all brothers.
MATT|23|9|And call no man your father on earth, for you have one Father, who is in heaven.
MATT|23|10|Neither be called instructors, for you have one instructor, the Christ.
MATT|23|11|The greatest among you shall be your servant.
MATT|23|12|Whoever exalts himself will be humbled, and whoever humbles himself will be exalted.
MATT|23|13|"But woe to you, scribes and Pharisees, hypocrites! For you shut the kingdom of heaven in people's faces. For you neither enter yourselves nor allow those who would enter to go in.
MATT|23|14|***
MATT|23|15|Woe to you, scribes and Pharisees, hypocrites! For you travel across sea and land to make a single proselyte, and when he becomes a proselyte, you make him twice as much a child of hell as yourselves.
MATT|23|16|"Woe to you, blind guides, who say, 'If anyone swears by the temple, it is nothing, but if anyone swears by the gold of the temple, he is bound by his oath.'
MATT|23|17|You blind fools! For which is greater, the gold or the temple that has made the gold sacred?
MATT|23|18|And you say, 'If anyone swears by the altar, it is nothing, but if anyone swears by the gift that is on the altar, he is bound by his oath.'
MATT|23|19|You blind men! For which is greater, the gift or the altar that makes the gift sacred?
MATT|23|20|So whoever swears by the altar swears by it and by everything on it.
MATT|23|21|And whoever swears by the temple swears by it and by him who dwells in it.
MATT|23|22|And whoever swears by heaven swears by the throne of God and by him who sits upon it.
MATT|23|23|"Woe to you, scribes and Pharisees, hypocrites! For you tithe mint and dill and cumin, and have neglected the weightier matters of the law: justice and mercy and faithfulness. These you ought to have done, without neglecting the others.
MATT|23|24|You blind guides, straining out a gnat and swallowing a camel!
MATT|23|25|"Woe to you, scribes and Pharisees, hypocrites! For you clean the outside of the cup and the plate, but inside they are full of greed and self-indulgence.
MATT|23|26|You blind Pharisee! First clean the inside of the cup and the plate, that the outside also may be clean.
MATT|23|27|"Woe to you, scribes and Pharisees, hypocrites! For you are like whitewashed tombs, which outwardly appear beautiful, but within are full of dead people's bones and all uncleanness.
MATT|23|28|So you also outwardly appear righteous to others, but within you are full of hypocrisy and lawlessness.
MATT|23|29|"Woe to you, scribes and Pharisees, hypocrites! For you build the tombs of the prophets and decorate the monuments of the righteous,
MATT|23|30|saying, 'If we had lived in the days of our fathers, we would not have taken part with them in shedding the blood of the prophets.'
MATT|23|31|Thus you witness against yourselves that you are sons of those who murdered the prophets.
MATT|23|32|Fill up, then, the measure of your fathers.
MATT|23|33|You serpents, you brood of vipers, how are you to escape being sentenced to hell?
MATT|23|34|Therefore I send you prophets and wise men and scribes, some of whom you will kill and crucify, and some you will flog in your synagogues and persecute from town to town,
MATT|23|35|so that on you may come all the righteous blood shed on earth, from the blood of innocent Abel to the blood of Zechariah the son of Barachiah, whom you murdered between the sanctuary and the altar.
MATT|23|36|Truly, I say to you, all these things will come upon this generation.
MATT|23|37|"O Jerusalem, Jerusalem, the city that kills the prophets and stones those who are sent to it! How often would I have gathered your children together as a hen gathers her brood under her wings, and you would not!
MATT|23|38|See, your house is left to you desolate.
MATT|23|39|For I tell you, you will not see me again, until you say, 'Blessed is he who comes in the name of the Lord.'"
MATT|24|1|Jesus left the temple and was going away, when his disciples came to point out to him the buildings of the temple.
MATT|24|2|But he answered them, "You see all these, do you not? Truly, I say to you, there will not be left here one stone upon another that will not be thrown down."
MATT|24|3|As he sat on the Mount of Olives, the disciples came to him privately, saying, "Tell us, when will these things be, and what will be the sign of your coming and of the close of the age?"
MATT|24|4|And Jesus answered them, "See that no one leads you astray.
MATT|24|5|For many will come in my name, saying, 'I am the Christ,' and they will lead many astray.
MATT|24|6|And you will hear of wars and rumors of wars. See that you are not alarmed, for this must take place, but the end is not yet.
MATT|24|7|For nation will rise against nation, and kingdom against kingdom, and there will be famines and earthquakes in various places.
MATT|24|8|All these are but the beginning of the birth pains.
MATT|24|9|"Then they will deliver you up to tribulation and put you to death, and you will be hated by all nations for my name's sake.
MATT|24|10|And then many will fall away and betray one another and hate one another.
MATT|24|11|And many false prophets will arise and lead many astray.
MATT|24|12|And because lawlessness will be increased, the love of many will grow cold.
MATT|24|13|But the one who endures to the end will be saved.
MATT|24|14|And this gospel of the kingdom will be proclaimed throughout the whole world as a testimony to all nations, and then the end will come.
MATT|24|15|"So when you see the abomination of desolation spoken of by the prophet Daniel, standing in the holy place (let the reader understand),
MATT|24|16|then let those who are in Judea flee to the mountains.
MATT|24|17|Let the one who is on the housetop not go down to take what is in his house,
MATT|24|18|and let the one who is in the field not turn back to take his cloak.
MATT|24|19|And alas for women who are pregnant and for those who are nursing infants in those days!
MATT|24|20|Pray that your flight may not be in winter or on a Sabbath.
MATT|24|21|For then there will be great tribulation, such as has not been from the beginning of the world until now, no, and never will be.
MATT|24|22|And if those days had not been cut short, no human being would be saved. But for the sake of the elect those days will be cut short.
MATT|24|23|Then if anyone says to you, 'Look, here is the Christ!' or 'There he is!' do not believe it.
MATT|24|24|For false christs and false prophets will arise and perform great signs and wonders, so as to lead astray, if possible, even the elect.
MATT|24|25|See, I have told you beforehand.
MATT|24|26|So, if they say to you, 'Look, he is in the wilderness,' do not go out. If they say, 'Look, he is in the inner rooms,' do not believe it.
MATT|24|27|For as the lightning comes from the east and shines as far as the west, so will be the coming of the Son of Man.
MATT|24|28|Wherever the corpse is, there the vultures will gather.
MATT|24|29|"Immediately after the tribulation of those days the sun will be darkened, and the moon will not give its light, and the stars will fall from heaven, and the powers of the heavens will be shaken.
MATT|24|30|Then will appear in heaven the sign of the Son of Man, and then all the tribes of the earth will mourn, and they will see the Son of Man coming on the clouds of heaven with power and great glory.
MATT|24|31|And he will send out his angels with a loud trumpet call, and they will gather his elect from the four winds, from one end of heaven to the other.
MATT|24|32|"From the fig tree learn its lesson: as soon as its branch becomes tender and puts out its leaves, you know that summer is near.
MATT|24|33|So also, when you see all these things, you know that he is near, at the very gates.
MATT|24|34|Truly, I say to you, this generation will not pass away until all these things take place.
MATT|24|35|Heaven and earth will pass away, but my words will not pass away.
MATT|24|36|"But concerning that day and hour no one knows, not even the angels of heaven, nor the Son, but the Father only.
MATT|24|37|As were the days of Noah, so will be the coming of the Son of Man.
MATT|24|38|For as in those days before the flood they were eating and drinking, marrying and giving in marriage, until the day when Noah entered the ark,
MATT|24|39|and they were unaware until the flood came and swept them all away, so will be the coming of the Son of Man.
MATT|24|40|Then two men will be in the field; one will be taken and one left.
MATT|24|41|Two women will be grinding at the mill; one will be taken and one left.
MATT|24|42|Therefore, stay awake, for you do not know on what day your Lord is coming.
MATT|24|43|But know this, that if the master of the house had known in what part of the night the thief was coming, he would have stayed awake and would not have let his house be broken into.
MATT|24|44|Therefore you also must be ready, for the Son of Man is coming at an hour you do not expect.
MATT|24|45|"Who then is the faithful and wise servant, whom his master has set over his household, to give them their food at the proper time?
MATT|24|46|Blessed is that servant whom his master will find so doing when he comes.
MATT|24|47|Truly, I say to you, he will set him over all his possessions.
MATT|24|48|But if that wicked servant says to himself, 'My master is delayed,'
MATT|24|49|and begins to beat his fellow servants and eats and drinks with drunkards,
MATT|24|50|the master of that servant will come on a day when he does not expect him and at an hour he does not know
MATT|24|51|and will cut him in pieces and put him with the hypocrites. In that place there will be weeping and gnashing of teeth.
MATT|25|1|"Then the kingdom of heaven will be like ten virgins who took their lamps and went to meet the bridegroom.
MATT|25|2|Five of them were foolish, and five were wise.
MATT|25|3|For when the foolish took their lamps, they took no oil with them,
MATT|25|4|but the wise took flasks of oil with their lamps.
MATT|25|5|As the bridegroom was delayed, they all became drowsy and slept.
MATT|25|6|But at midnight there was a cry, 'Here is the bridegroom! Come out to meet him.'
MATT|25|7|Then all those virgins rose and trimmed their lamps.
MATT|25|8|And the foolish said to the wise, 'Give us some of your oil, for our lamps are going out.'
MATT|25|9|But the wise answered, saying, 'Since there will not be enough for us and for you, go rather to the dealers and buy for yourselves.'
MATT|25|10|And while they were going to buy, the bridegroom came, and those who were ready went in with him to the marriage feast, and the door was shut.
MATT|25|11|Afterward the other virgins came also, saying, 'Lord, lord, open to us.'
MATT|25|12|But he answered, 'Truly, I say to you, I do not know you.'
MATT|25|13|Watch therefore, for you know neither the day nor the hour.
MATT|25|14|"For it will be like a man going on a journey, who called his servants and entrusted to them his property.
MATT|25|15|To one he gave five talents, to another two, to another one, to each according to his ability. Then he went away.
MATT|25|16|He who had received the five talents went at once and traded with them, and he made five talents more.
MATT|25|17|So also he who had the two talents made two talents more.
MATT|25|18|But he who had received the one talent went and dug in the ground and hid his master's money.
MATT|25|19|Now after a long time the master of those servants came and settled accounts with them.
MATT|25|20|And he who had received the five talents came forward, bringing five talents more, saying, 'Master, you delivered to me five talents; here I have made five talents more.'
MATT|25|21|His master said to him, 'Well done, good and faithful servant. You have been faithful over a little; I will set you over much. Enter into the joy of your master.'
MATT|25|22|And he also who had the two talents came forward, saying, 'Master, you delivered to me two talents; here I have made two talents more.'
MATT|25|23|His master said to him, 'Well done, good and faithful servant. You have been faithful over a little; I will set you over much. Enter into the joy of your master.'
MATT|25|24|He also who had received the one talent came forward, saying, 'Master, I knew you to be a hard man, reaping where you did not sow, and gathering where you scattered no seed,
MATT|25|25|so I was afraid, and I went and hid your talent in the ground. Here you have what is yours.'
MATT|25|26|But his master answered him, 'You wicked and slothful servant! You knew that I reap where I have not sowed and gather where I scattered no seed?
MATT|25|27|Then you ought to have invested my money with the bankers, and at my coming I should have received what was my own with interest.
MATT|25|28|So take the talent from him and give it to him who has the ten talents.
MATT|25|29|For to everyone who has will more be given, and he will have an abundance. But from the one who has not, even what he has will be taken away.
MATT|25|30|And cast the worthless servant into the outer darkness. In that place there will be weeping and gnashing of teeth.'
MATT|25|31|"When the Son of Man comes in his glory, and all the angels with him, then he will sit on his glorious throne.
MATT|25|32|Before him will be gathered all the nations, and he will separate people one from another as a shepherd separates the sheep from the goats.
MATT|25|33|And he will place the sheep on his right, but the goats on the left.
MATT|25|34|Then the King will say to those on his right, 'Come, you who are blessed by my Father, inherit the kingdom prepared for you from the foundation of the world.
MATT|25|35|For I was hungry and you gave me food, I was thirsty and you gave me drink, I was a stranger and you welcomed me,
MATT|25|36|I was naked and you clothed me, I was sick and you visited me, I was in prison and you came to me.'
MATT|25|37|Then the righteous will answer him, saying, 'Lord, when did we see you hungry and feed you, or thirsty and give you drink?
MATT|25|38|And when did we see you a stranger and welcome you, or naked and clothe you?
MATT|25|39|And when did we see you sick or in prison and visit you?'
MATT|25|40|And the King will answer them, 'Truly, I say to you, as you did it to one of the least of these my brothers, you did it to me.'
MATT|25|41|"Then he will say to those on his left, 'Depart from me, you cursed, into the eternal fire prepared for the devil and his angels.
MATT|25|42|For I was hungry and you gave me no food, I was thirsty and you gave me no drink,
MATT|25|43|I was a stranger and you did not welcome me, naked and you did not clothe me, sick and in prison and you did not visit me.'
MATT|25|44|Then they also will answer, saying, 'Lord, when did we see you hungry or thirsty or a stranger or naked or sick or in prison, and did not minister to you?'
MATT|25|45|Then he will answer them, saying, 'Truly, I say to you, as you did not do it to one of the least of these, you did not do it to me.'
MATT|25|46|And these will go away into eternal punishment, but the righteous into eternal life."
MATT|26|1|When Jesus had finished all these sayings, he said to his disciples,
MATT|26|2|"You know that after two days the Passover is coming, and the Son of Man will be delivered up to be crucified."
MATT|26|3|Then the chief priests and the elders of the people gathered in the palace of the high priest, whose name was Caiaphas,
MATT|26|4|and plotted together in order to arrest Jesus by stealth and kill him.
MATT|26|5|But they said, "Not during the feast, lest there be an uproar among the people."
MATT|26|6|Now when Jesus was at Bethany in the house of Simon the leper,
MATT|26|7|a woman came up to him with an alabaster flask of very expensive ointment, and she poured it on his head as he reclined at table.
MATT|26|8|And when the disciples saw it, they were indignant, saying, "Why this waste?
MATT|26|9|For this could have been sold for a large sum and given to the poor."
MATT|26|10|But Jesus, aware of this, said to them, "Why do you trouble the woman? For she has done a beautiful thing to me.
MATT|26|11|For you always have the poor with you, but you will not always have me.
MATT|26|12|In pouring this ointment on my body, she has done it to prepare me for burial.
MATT|26|13|Truly, I say to you, wherever this gospel is proclaimed in the whole world, what she has done will also be told in memory of her."
MATT|26|14|Then one of the twelve, whose name was Judas Iscariot, went to the chief priests
MATT|26|15|and said, "What will you give me if I deliver him over to you?" And they paid him thirty pieces of silver.
MATT|26|16|And from that moment he sought an opportunity to betray him.
MATT|26|17|Now on the first day of Unleavened Bread the disciples came to Jesus, saying, "Where will you have us prepare for you to eat the Passover?"
MATT|26|18|He said, "Go into the city to a certain man and say to him, 'The Teacher says, My time is at hand. I will keep the Passover at your house with my disciples.'"
MATT|26|19|And the disciples did as Jesus had directed them, and they prepared the Passover.
MATT|26|20|When it was evening, he reclined at table with the twelve.
MATT|26|21|And as they were eating, he said, "Truly, I say to you, one of you will betray me."
MATT|26|22|And they were very sorrowful and began to say to him one after another, "Is it I, Lord?"
MATT|26|23|He answered, "He who has dipped his hand in the dish with me will betray me.
MATT|26|24|The Son of Man goes as it is written of him, but woe to that man by whom the Son of Man is betrayed! It would have been better for that man if he had not been born."
MATT|26|25|Judas, who would betray him, answered, "Is it I, Rabbi?" He said to him, "You have said so."
MATT|26|26|Now as they were eating, Jesus took bread, and after blessing it broke it and gave it to the disciples, and said, "Take, eat; this is my body."
MATT|26|27|And he took a cup, and when he had given thanks he gave it to them, saying, "Drink of it, all of you,
MATT|26|28|for this is my blood of the covenant, which is poured out for many for the forgiveness of sins.
MATT|26|29|I tell you I will not drink again of this fruit of the vine until that day when I drink it new with you in my Father's kingdom."
MATT|26|30|And when they had sung a hymn, they went out to the Mount of Olives.
MATT|26|31|Then Jesus said to them, "You will all fall away because of me this night. For it is written, 'I will strike the shepherd, and the sheep of the flock will be scattered.'
MATT|26|32|But after I am raised up, I will go before you to Galilee."
MATT|26|33|Peter answered him, "Though they all fall away because of you, I will never fall away."
MATT|26|34|Jesus said to him, "Truly, I tell you, this very night, before the rooster crows, you will deny me three times."
MATT|26|35|Peter said to him, "Even if I must die with you, I will not deny you!" And all the disciples said the same.
MATT|26|36|Then Jesus went with them to a place called Gethsemane, and he said to his disciples, "Sit here, while I go over there and pray."
MATT|26|37|And taking with him Peter and the two sons of Zebedee, he began to be sorrowful and troubled.
MATT|26|38|Then he said to them, "My soul is very sorrowful, even to death; remain here, and watch with me."
MATT|26|39|And going a little farther he fell on his face and prayed, saying, "My Father, if it be possible, let this cup pass from me; nevertheless, not as I will, but as you will."
MATT|26|40|And he came to the disciples and found them sleeping. And he said to Peter, "So, could you not watch with me one hour?
MATT|26|41|Watch and pray that you may not enter into temptation. The spirit indeed is willing, but the flesh is weak."
MATT|26|42|Again, for the second time, he went away and prayed, "My Father, if this cannot pass unless I drink it, your will be done."
MATT|26|43|And again he came and found them sleeping, for their eyes were heavy.
MATT|26|44|So, leaving them again, he went away and prayed for the third time, saying the same words again.
MATT|26|45|Then he came to the disciples and said to them, "Sleep and take your rest later on. See, the hour is at hand, and the Son of Man is betrayed into the hands of sinners.
MATT|26|46|Rise, let us be going; see, my betrayer is at hand."
MATT|26|47|While he was still speaking, Judas came, one of the twelve, and with him a great crowd with swords and clubs, from the chief priests and the elders of the people.
MATT|26|48|Now the betrayer had given them a sign, saying, "The one I will kiss is the man; seize him."
MATT|26|49|And he came up to Jesus at once and said, "Greetings, Rabbi!" And he kissed him.
MATT|26|50|Jesus said to him, "Friend, do what you came to do." Then they came up and laid hands on Jesus and seized him.
MATT|26|51|And behold, one of those who were with Jesus stretched out his hand and drew his sword and struck the servant of the high priest and cut off his ear.
MATT|26|52|Then Jesus said to him, "Put your sword back into its place. For all who take the sword will perish by the sword.
MATT|26|53|Do you think that I cannot appeal to my Father, and he will at once send me more than twelve legions of angels?
MATT|26|54|But how then should the Scriptures be fulfilled, that it must be so?"
MATT|26|55|At that hour Jesus said to the crowds, "Have you come out as against a robber, with swords and clubs to capture me? Day after day I sat in the temple teaching, and you did not seize me.
MATT|26|56|But all this has taken place that the Scriptures of the prophets might be fulfilled." Then all the disciples left him and fled.
MATT|26|57|Then those who had seized Jesus led him to Caiaphas the high priest, where the scribes and the elders had gathered.
MATT|26|58|And Peter was following him at a distance, as far as the courtyard of the high priest, and going inside he sat with the guards to see the end.
MATT|26|59|Now the chief priests and the whole Council were seeking false testimony against Jesus that they might put him to death,
MATT|26|60|but they found none, though many false witnesses came forward. At last two came forward
MATT|26|61|and said, "This man said, 'I am able to destroy the temple of God, and to rebuild it in three days.'"
MATT|26|62|And the high priest stood up and said, "Have you no answer to make? What is it that these men testify against you?"
MATT|26|63|But Jesus remained silent. And the high priest said to him, "I adjure you by the living God, tell us if you are the Christ, the Son of God."
MATT|26|64|Jesus said to him, "You have said so. But I tell you, from now on you will see the Son of Man seated at the right hand of Power and coming on the clouds of heaven."
MATT|26|65|Then the high priest tore his robes and said, "He has uttered blasphemy. What further witnesses do we need? You have now heard his blasphemy.
MATT|26|66|What is your judgment?" They answered, "He deserves death."
MATT|26|67|Then they spit in his face and struck him. And some slapped him,
MATT|26|68|saying, "Prophesy to us, you Christ! Who is it that struck you?"
MATT|26|69|Now Peter was sitting outside in the courtyard. And a servant girl came up to him and said, "You also were with Jesus the Galilean."
MATT|26|70|But he denied it before them all, saying, "I do not know what you mean."
MATT|26|71|And when he went out to the entrance, another servant girl saw him, and she said to the bystanders, "This man was with Jesus of Nazareth."
MATT|26|72|And again he denied it with an oath: "I do not know the man."
MATT|26|73|After a little while the bystanders came up and said to Peter, "Certainly you too are one of them, for your accent betrays you."
MATT|26|74|Then he began to invoke a curse on himself and to swear, "I do not know the man." And immediately the rooster crowed.
MATT|26|75|And Peter remembered the saying of Jesus, "Before the rooster crows, you will deny me three times." And he went out and wept bitterly.
MATT|27|1|When morning came, all the chief priests and the elders of the people took counsel against Jesus to put him to death.
MATT|27|2|And they bound him and led him away and delivered him over to Pilate the governor.
MATT|27|3|Then when Judas, his betrayer, saw that Jesus was condemned, he changed his mind and brought back the thirty pieces of silver to the chief priests and the elders,
MATT|27|4|saying, "I have sinned by betraying innocent blood." They said, "What is that to us? See to it yourself."
MATT|27|5|And throwing down the pieces of silver into the temple, he departed, and he went and hanged himself.
MATT|27|6|But the chief priests, taking the pieces of silver, said, "It is not lawful to put them into the treasury, since it is blood money."
MATT|27|7|So they took counsel and bought with them the potter's field as a burial place for strangers.
MATT|27|8|Therefore that field has been called the Field of Blood to this day.
MATT|27|9|Then was fulfilled what had been spoken by the prophet Jeremiah, saying, "And they took the thirty pieces of silver, the price of him on whom a price had been set by some of the sons of Israel,
MATT|27|10|and they gave them for the potter's field, as the Lord directed me."
MATT|27|11|Now Jesus stood before the governor, and the governor asked him, "Are you the King of the Jews?" Jesus said, "You have said so."
MATT|27|12|But when he was accused by the chief priests and elders, he gave no answer.
MATT|27|13|Then Pilate said to him, "Do you not hear how many things they testify against you?"
MATT|27|14|But he gave him no answer, not even to a single charge, so that the governor was greatly amazed.
MATT|27|15|Now at the feast the governor was accustomed to release for the crowd any one prisoner whom they wanted.
MATT|27|16|And they had then a notorious prisoner called Barabbas.
MATT|27|17|So when they had gathered, Pilate said to them, "Whom do you want me to release for you: Barabbas, or Jesus who is called Christ?"
MATT|27|18|For he knew that it was out of envy that they had delivered him up.
MATT|27|19|Besides, while he was sitting on the judgment seat, his wife sent word to him, "Have nothing to do with that righteous man, for I have suffered much because of him today in a dream."
MATT|27|20|Now the chief priests and the elders persuaded the crowd to ask for Barabbas and destroy Jesus.
MATT|27|21|The governor again said to them, "Which of the two do you want me to release for you?" And they said, "Barabbas."
MATT|27|22|Pilate said to them, "Then what shall I do with Jesus who is called Christ?" They all said, "Let him be crucified!"
MATT|27|23|And he said, "Why, what evil has he done?" But they shouted all the more, "Let him be crucified!"
MATT|27|24|So when Pilate saw that he was gaining nothing, but rather that a riot was beginning, he took water and washed his hands before the crowd, saying, "I am innocent of this man's blood; see to it yourselves."
MATT|27|25|And all the people answered, "His blood be on us and on our children!"
MATT|27|26|Then he released for them Barabbas, and having scourged Jesus, delivered him to be crucified.
MATT|27|27|Then the soldiers of the governor took Jesus into the governor's headquarters, and they gathered the whole battalion before him.
MATT|27|28|And they stripped him and put a scarlet robe on him,
MATT|27|29|and twisting together a crown of thorns, they put it on his head and put a reed in his right hand. And kneeling before him, they mocked him, saying, "Hail, King of the Jews!"
MATT|27|30|And they spit on him and took the reed and struck him on the head.
MATT|27|31|And when they had mocked him, they stripped him of the robe and put his own clothes on him and led him away to crucify him.
MATT|27|32|As they went out, they found a man of Cyrene, Simon by name. They compelled this man to carry his cross.
MATT|27|33|And when they came to a place called Golgotha (which means Place of a Skull),
MATT|27|34|they offered him wine to drink, mixed with gall, but when he tasted it, he would not drink it.
MATT|27|35|And when they had crucified him, they divided his garments among them by casting lots.
MATT|27|36|Then they sat down and kept watch over him there.
MATT|27|37|And over his head they put the charge against him, which read, "This is Jesus, the King of the Jews."
MATT|27|38|Then two robbers were crucified with him, one on the right and one on the left.
MATT|27|39|And those who passed by derided him, wagging their heads
MATT|27|40|and saying, "You who would destroy the temple and rebuild it in three days, save yourself! If you are the Son of God, come down from the cross."
MATT|27|41|So also the chief priests, with the scribes and elders, mocked him, saying,
MATT|27|42|"He saved others; he cannot save himself. He is the King of Israel; let him come down now from the cross, and we will believe in him.
MATT|27|43|He trusts in God; let God deliver him now, if he desires him. For he said, 'I am the Son of God.'"
MATT|27|44|And the robbers who were crucified with him also reviled him in the same way.
MATT|27|45|Now from the sixth hour there was darkness over all the land until the ninth hour.
MATT|27|46|And about the ninth hour Jesus cried out with a loud voice, saying, "Eli, Eli, lema sabachthani?" that is, "My God, my God, why have you forsaken me?"
MATT|27|47|And some of the bystanders, hearing it, said, "This man is calling Elijah."
MATT|27|48|And one of them at once ran and took a sponge, filled it with sour wine, and put it on a reed and gave it to him to drink.
MATT|27|49|But the others said, "Wait, let us see whether Elijah will come to save him."
MATT|27|50|And Jesus cried out again with a loud voice and yielded up his spirit.
MATT|27|51|And behold, the curtain of the temple was torn in two, from top to bottom. And the earth shook, and the rocks were split.
MATT|27|52|The tombs also were opened. And many bodies of the saints who had fallen asleep were raised,
MATT|27|53|and coming out of the tombs after his resurrection they went into the holy city and appeared to many.
MATT|27|54|When the centurion and those who were with him, keeping watch over Jesus, saw the earthquake and what took place, they were filled with awe and said, "Truly this was the Son of God!"
MATT|27|55|There were also many women there, looking on from a distance, who had followed Jesus from Galilee, ministering to him,
MATT|27|56|among whom were Mary Magdalene and Mary the mother of James and Joseph and the mother of the sons of Zebedee.
MATT|27|57|When it was evening, there came a rich man from Arimathea, named Joseph, who also was a disciple of Jesus.
MATT|27|58|He went to Pilate and asked for the body of Jesus. Then Pilate ordered it to be given to him.
MATT|27|59|And Joseph took the body and wrapped it in a clean linen shroud
MATT|27|60|and laid it in his own new tomb, which he had cut in the rock. And he rolled a great stone to the entrance of the tomb and went away.
MATT|27|61|Mary Magdalene and the other Mary were there, sitting opposite the tomb.
MATT|27|62|Next day, that is, after the day of Preparation, the chief priests and the Pharisees gathered before Pilate
MATT|27|63|and said, "Sir, we remember how that impostor said, while he was still alive, 'After three days I will rise.'
MATT|27|64|Therefore order the tomb to be made secure until the third day, lest his disciples go and steal him away and tell the people, 'He has risen from the dead,' and the last fraud will be worse than the first."
MATT|27|65|Pilate said to them, "You have a guard of soldiers. Go, make it as secure as you can."
MATT|27|66|So they went and made the tomb secure by sealing the stone and setting a guard.
MATT|28|1|Now after the Sabbath, toward the dawn of the first day of the week, Mary Magdalene and the other Mary went to see the tomb.
MATT|28|2|And behold, there was a great earthquake, for an angel of the Lord descended from heaven and came and rolled back the stone and sat on it.
MATT|28|3|His appearance was like lightning, and his clothing white as snow.
MATT|28|4|And for fear of him the guards trembled and became like dead men.
MATT|28|5|But the angel said to the women, "Do not be afraid, for I know that you seek Jesus who was crucified.
MATT|28|6|He is not here, for he has risen, as he said. Come, see the place where he lay.
MATT|28|7|Then go quickly and tell his disciples that he has risen from the dead, and behold, he is going before you to Galilee; there you will see him. See, I have told you."
MATT|28|8|So they departed quickly from the tomb with fear and great joy, and ran to tell his disciples.
MATT|28|9|And behold, Jesus met them and said, "Greetings!" And they came up and took hold of his feet and worshiped him.
MATT|28|10|Then Jesus said to them, "Do not be afraid; go and tell my brothers to go to Galilee, and there they will see me."
MATT|28|11|While they were going, behold, some of the guard went into the city and told the chief priests all that had taken place.
MATT|28|12|And when they had assembled with the elders and taken counsel, they gave a sufficient sum of money to the soldiers
MATT|28|13|and said, "Tell people, 'His disciples came by night and stole him away while we were asleep.'
MATT|28|14|And if this comes to the governor's ears, we will satisfy him and keep you out of trouble."
MATT|28|15|So they took the money and did as they were directed. And this story has been spread among the Jews to this day.
MATT|28|16|Now the eleven disciples went to Galilee, to the mountain to which Jesus had directed them.
MATT|28|17|And when they saw him they worshiped him, but some doubted.
MATT|28|18|And Jesus came and said to them, "All authority in heaven and on earth has been given to me.
MATT|28|19|Go therefore and make disciples of all nations, baptizing them in the name of the Father and of the Son and of the Holy Spirit,
MATT|28|20|teaching them to observe all that I have commanded you. And behold, I am with you always, to the end of the age."
