PROV|1|1|Parabolae Salomonis filii David regis Israel
PROV|1|2|ad sciendam sapientiam et disciplinam,ad intellegenda verba prudentiae;
PROV|1|3|ad suscipiendam eruditionem doctrinae,iustitiam et iudicium et aequitatem,
PROV|1|4|ut detur parvulis astutia,adulescenti scientia et recogitatio.
PROV|1|5|Audiat sapiens et addet doctrinam,et intellegens dispositiones possidebit:
PROV|1|6|animadvertet parabolam et allegoriam,verba sapientium et aenigmata eorum.
PROV|1|7|Timor Domini principium scientiae.Sapientiam atque doctrinam stulti despiciunt.
PROV|1|8|Audi, fili mi, disciplinam patris tuiet ne reicias legem matris tuae,
PROV|1|9|quia diadema gratiae sunt capiti tuo,et torques collo tuo.
PROV|1|10|Fili mi, si te lactaverint peccatores,ne acquiescas eis.
PROV|1|11|Si dixerint: " Veni nobiscum, insidiemur sanguini,abscondamus tendiculas contra insontem frustra;
PROV|1|12|deglutiamus eos sicut infernus viventeset integros quasi descendentes in lacum:
PROV|1|13|omnem pretiosam substantiam reperiemus,implebimus domos nostras spoliis;
PROV|1|14|sortem mitte nobiscum,marsupium unum sit omnium nostrum ";
PROV|1|15|fili mi, ne ambules cum eis,prohibe pedem tuum a semitis eorum.
PROV|1|16|Pedes enim illorum ad malum curruntet festinant, ut effundant sanguinem.
PROV|1|17|Frustra autem iacitur rete ante oculos pinnatorum.
PROV|1|18|Ipsique contra sanguinem suum insidianturet moliuntur fraudes contra animas suas.
PROV|1|19|Sic semitae omnis ad rapinam intenti:animam ipsius possidentis rapiunt.
PROV|1|20|Sapientia foris praedicat,in plateis dat vocem suam,
PROV|1|21|in capite viarum frequentium clamitat,in foribus portarum urbis profert verba sua:
PROV|1|22|" Usquequo, parvuli, diligitis infantiam,et derisores sibi derisionem cupient,et imprudentes odibunt scientiam?
PROV|1|23|Convertimini ad correptionem meam;en proferam vobis spiritum meumet ostendam vobis verba mea.
PROV|1|24|Quia vocavi, et renuistis,extendi manum meam, et non fuit qui aspiceret;
PROV|1|25|despexistis omne consilium meumet increpationes meas neglexistis.
PROV|1|26|Ego quoque in interitu vestro rideboet subsannabo, cum terror vobis advenerit,
PROV|1|27|cum irruerit ut procella terror,et interitus quasi tempestas ingruerit,quando venerit super vos tribulatio et angustia ".
PROV|1|28|Tunc invocabunt me, et non exaudiam,instanter quaerent me et non invenient me,
PROV|1|29|eo quod exosam habuerint disciplinamet timorem Domini non elegerint
PROV|1|30|nec acquieverint consilio meoet despexerint universam correptionem meam.
PROV|1|31|Comedent igitur fructus viae suaesuisque consiliis saturabuntur.
PROV|1|32|Aversio parvulorum interficiet eos,et securitas stultorum perdet illos.
PROV|1|33|Qui autem me audierit, absque terrore requiescetet tranquillus erit timore malorum sublato.
PROV|2|1|Fili mi, si susceperis sermones meoset mandata mea absconderis penes te,
PROV|2|2|intendens ad sapientiam aurem tuam,inclinans cor tuum ad cognoscendam prudentiam;
PROV|2|3|si enim sapientiam invocaveriset dederis vocem tuam prudentiae,
PROV|2|4|si quaesieris eam quasi pecuniamet sicut thesauros conquisieris illam,
PROV|2|5|tunc intelleges timorem Dominiet scientiam Dei invenies.
PROV|2|6|Quia Dominus dat sapientiam,et ex ore eius scientia et prudentia.
PROV|2|7|Thesaurizabit rectis sollertiamet clipeus erit gradientibus simpliciter
PROV|2|8|servans semitas iustitiaeet vias sanctorum custodiens.
PROV|2|9|Tunc intelleges iustitiam et iudiciumet aequitatem et omnem semitam bonam,
PROV|2|10|quia intrabit sapientia cor tuum,et scientia animae tuae placebit.
PROV|2|11|Consilium custodiet te,et prudentia servabit te,
PROV|2|12|ut eruaris a via malaet ab homine, qui perversa loquitur;
PROV|2|13|qui relinquunt iter rectum,ut ambulent per vias tenebrosas;
PROV|2|14|qui laetantur, cum malefecerint,et exsultant in rebus pessimis:
PROV|2|15|quorum viae perversae sunt,et pravi gressus eorum.
PROV|2|16|Ut eruaris a muliere alienaet ab extranea, quae mollit sermones suos
PROV|2|17|et relinquit ducem pubertatis suaeet pacti Dei sui oblita est.
PROV|2|18|Inclinata est enim ad mortem domus eius,et ad inferos semitae ipsius;
PROV|2|19|omnes, qui ingrediuntur ad eam, non revertenturnec apprehendent semitas vitae.
PROV|2|20|Ut ambules in via bonorumet calles iustorum custodias:
PROV|2|21|qui enim recti sunt, habitabunt in terra,et simplices permanebunt in ea;
PROV|2|22|impii vero de terra perdentur,et, qui inique agunt, auferentur ex ea.
PROV|3|1|Fili mi, ne obliviscaris legis meae,et praecepta mea cor tuum custodiat;
PROV|3|2|longitudinem enim dierum et annos vitaeet pacem apponent tibi.
PROV|3|3|Misericordia et veritas te non deserant;circumda eas gutturi tuoet describe in tabulis cordis tui,
PROV|3|4|et invenies gratiam et successum bonumcoram Deo et hominibus.
PROV|3|5|Habe fiduciam in Domino ex toto corde tuoet ne innitaris prudentiae tuae.
PROV|3|6|In omnibus viis tuis cogita illum,et ipse diriget gressus tuos.
PROV|3|7|Ne sis sapiens apud temetipsum;time Dominum et recede a malo.
PROV|3|8|Sanitas quippe erit umbilico tuo,et irrigatio ossibus tuis.
PROV|3|9|Honora Dominum de tua substantiaet de primitiis omnium frugum tuarum,
PROV|3|10|et implebuntur horrea tua frumento,et vino torcularia tua redundabunt.
PROV|3|11|Disciplinam Domini, fili mi, ne abiciasnec asperneris, cum ab eo corriperis:
PROV|3|12|quem enim diligit, Dominus corripitet quasi pater in filio complacet sibi.
PROV|3|13|Beatus homo, qui invenit sapientiamet qui affluit prudentia:
PROV|3|14|melior est acquisitio eius negotiatione argenti,et auro primo fructus eius.
PROV|3|15|Pretiosior est cunctis gemmis,et omnia pretiosa tua huic non valent comparari;
PROV|3|16|longitudo dierum in dextera eius,et in sinistra illius divitiae et gloria.
PROV|3|17|Viae eius viae pulchrae,et omnes semitae illius pacificae.
PROV|3|18|Lignum vitae est his, qui apprehenderint eam;et, qui tenuerit eam, beatus.
PROV|3|19|Dominus sapientia fundavit terram,stabilivit caelos prudentia;
PROV|3|20|sapientia illius eruperunt abyssi,et nubes rorem stillant.
PROV|3|21|Fili mi, ne effluant haec ab oculis tuis;custodi prudentiam atque consilium,
PROV|3|22|et erit vita animae tuae,et gratia collo tuo;
PROV|3|23|tunc ambulabis fiducialiter in via tua,et pes tuus non impinget.
PROV|3|24|Si dormieris, non timebis;quiesces, et suavis erit somnus tuus.
PROV|3|25|Ne paveas repentino terroreet irruentem tibi turbinem impiorum, cum venerit.
PROV|3|26|Dominus enim erit in latere tuoet custodiet pedem tuum, ne capiaris.
PROV|3|27|Noli prohibere beneficium ab eo, cui debetur,si in potestate manus tuae est, ut facias.
PROV|3|28|Ne dicas amico tuo: " Vade et revertere,cras dabo tibi ", cum statim possis dare.
PROV|3|29|Ne moliaris amico tuo malum,cum ille apud te sedeat cum fiducia.
PROV|3|30|Ne contendas adversus hominem frustra,cum ipse tibi nihil mali fecerit.
PROV|3|31|Ne aemuleris hominem iniustumnec imiteris omnes vias eius,
PROV|3|32|quia abominatio Domini est omnis pravus,et cum simplicibus societas eius.
PROV|3|33|Maledictio a Domino in domo impii,habitacula autem iustorum benedicentur.
PROV|3|34|Ipse deludet illusoreset mansuetis dabit gratiam;
PROV|3|35|gloriam sapientes possidebunt,stultorum exaltatio ignominia.
PROV|4|1|Audite, filii, disciplinam patriset attendite, ut sciatis prudentiam;
PROV|4|2|quoniam doctrinam bonam tribuam vobis,legem meam ne derelinquatis.
PROV|4|3|Nam et ego filius fui patris mei,tenellus et unigenitus coram matre mea;
PROV|4|4|et docebat me atque dicebat: Suscipiat verba mea cor tuum,custodi praecepta mea et vives.
PROV|4|5|Posside sapientiam, posside prudentiam,ne obliviscaris neque declines a verbis oris mei.
PROV|4|6|Ne dimittas eam, et custodiet te,dilige eam, et servabit te.
PROV|4|7|Principium sapientiae: posside sapientiamet in omni possessione tua acquire prudentiam.
PROV|4|8|Arripe illam, et exaltabit te,glorificaberis ab ea, cum eam fueris amplexatus.
PROV|4|9|Dabit capiti tuo diadema gratiae,et corona inclita proteget te ".
PROV|4|10|Audi, fili mi, et suscipe verba mea,ut multiplicentur tibi anni vitae.
PROV|4|11|Viam sapientiae monstravi tibi;duxi te per semitas aequitatis,
PROV|4|12|quas cum ingressus fueris, non arctabuntur gressus tui,et currens non habebis offendiculum.
PROV|4|13|Tene disciplinam nec laxes;custodi illam, quia ipsa est vita tua.
PROV|4|14|Ne ingrediaris in semitas impiorumnec procedas in malorum via.
PROV|4|15|Fuge ab ea nec transeas per illam;declina et desere eam.
PROV|4|16|Non enim dormiunt, nisi malefecerint,et rapitur somnus ab eis, nisi supplantaverint.
PROV|4|17|Comedunt enim panem impietatiset vinum iniquitatis bibunt.
PROV|4|18|Iustorum autem semita quasi lux splendensprocedit et crescit usque ad perfectam diem.
PROV|4|19|Via impiorum tenebrosa;nesciunt, ubi corruant.
PROV|4|20|Fili mi, ausculta sermones meoset ad eloquia mea inclina aurem tuam;
PROV|4|21|ne recedant ab oculis tuis,custodi ea in medio cordis tui:
PROV|4|22|vita enim sunt invenientibus ea,et universae carni sanitas.
PROV|4|23|Omni custodia serva cor tuum,quia ex ipso vita procedit.
PROV|4|24|Remove a te os pravum,et detrahentia labia sint procul a te.
PROV|4|25|Oculi tui recta videant,et palpebrae tuae dirigantur coram te.
PROV|4|26|Observa semitam pedum tuorum,et omnes viae tuae stabilientur.
PROV|4|27|Ne declines ad dexteram neque ad sinistram,averte pedem tuum a malo.
PROV|5|1|Fili mi, attende ad sapientiam meam,et prudentiae meae inclina aurem tuam,
PROV|5|2|ut custodias cogitationes,et disciplinam labia tua conservent.
PROV|5|3|Favum enim stillant labia meretricis,et nitidius oleo guttur eius;
PROV|5|4|novissima autem illius amara quasi absinthiumet acuta quasi gladius biceps.
PROV|5|5|Pedes eius descendunt in mortem,et ad inferos gressus illius tendunt;
PROV|5|6|cum non observet semitam vitae,vagi sunt gressus eius, et ipsa nescit.
PROV|5|7|Nunc ergo, fili mi, audi meet ne recedas a verbis oris mei.
PROV|5|8|Longe fac ab ea viam tuamet ne appropinques foribus domus eius.
PROV|5|9|Ne des alienis honorem tuumet annos tuos crudeli,
PROV|5|10|ne forte impleantur extranei viribus tuis,et labores tui sint in domo aliena,
PROV|5|11|et gemas in novissimis,quando consumpseris carnes tuas et corpus tuum
PROV|5|12|et dicas: " Cur detestatus sum disciplinam,et increpationes renuit cor meum,
PROV|5|13|nec audivi vocem docentium meet magistris non inclinavi aurem meam?
PROV|5|14|Paene fui in omni malo,in medio ecclesiae et synagogae ".
PROV|5|15|Bibe aquam de cisterna tuaet fluenta putei tui,
PROV|5|16|ne deriventur fontes tui foras,et in plateis rivi aquarum;
PROV|5|17|habeto eas solus,nec sint alieni participes tui.
PROV|5|18|Sit vena tua benedicta,et laetare cum muliere adulescentiae tuae;
PROV|5|19|cerva carissima et gratissimus hinnulus,blanditiae eius inebrient te in omni tempore,in amore eius delectare iugiter.
PROV|5|20|Quare seduceris, fili mi, ab alienaet foveris in sinu extraneae?
PROV|5|21|Quoniam ante Dominum viae hominis,et omnes gressus eius considerat.
PROV|5|22|Iniquitates suae capient impium,et funibus peccatorum suorum constringetur.
PROV|5|23|Ipse morietur, quia non habuit disciplinam,et in multitudine stultitiae suae decipietur.
PROV|6|1|Fili mi, si spoponderis pro amico tuo,defixisti apud extraneum manum tuam;
PROV|6|2|illaqueatus es verbis oris tuiet captus propriis sermonibus.
PROV|6|3|Fac ergo, quod dico, fili mi, et temetipsum libera,quia incidisti in manum proximi tui;discurre, prosternere, insta amico tuo.
PROV|6|4|Ne dederis somnum oculis tuisnec palpebris tuis dormitationem.
PROV|6|5|Eruere quasi dammula de rete,et quasi avis de manu aucupis.
PROV|6|6|Vade ad formicam, o piger,et considera vias eius et disce sapientiam.
PROV|6|7|Quae, cum non habeat ducemnec praeceptorem nec principem,
PROV|6|8|parat in aestate cibum sibiet congregat in messe, quod comedat.
PROV|6|9|Usquequo, piger, dormies?Quando consurges e somno tuo?
PROV|6|10|Paululum dormis, paululum dormitas,paululum conseres manus, ut dormias;
PROV|6|11|et veniet tibi quasi viator egestas,et pauperies quasi vir armatus.
PROV|6|12|Homo iniquus, vir inutilis,graditur ore perverso;
PROV|6|13|annuit oculis, terit pede,digito loquitur.
PROV|6|14|Prava in corde suo machinatur,malum in omni tempore, iurgia seminat.
PROV|6|15|Ideo extemplo veniet perditio sua,et subito conteretur nec habebit medicinam.
PROV|6|16|Sex sunt, quae odit Dominus,et septem detestatur anima eius:
PROV|6|17|oculos sublimes, linguam mendacem,manus effundentes innoxium sanguinem,
PROV|6|18|cor machinans cogitationes pravas,pedes veloces ad currendum in malum,
PROV|6|19|proferentem mendacia, testem fallacemet eum, qui seminat inter fratres discordias.
PROV|6|20|Conserva, fili mi, praecepta patris tuiet ne reicias legem matris tuae;
PROV|6|21|liga ea in corde tuo iugiteret circumda gutturi tuo.
PROV|6|22|Cum ambulaveris, dirigent te,cum dormieris, custodient teet, cum evigilaveris, colloquentur tecum.
PROV|6|23|Quia mandatum lucerna est, et lex lux,et via vitae increpatio disciplinae,
PROV|6|24|ut custodiant te a muliere malaet a blanda lingua extraneae;
PROV|6|25|non concupiscat pulchritudinem eius cor tuum,nec capiaris nutibus illius:
PROV|6|26|pretium enim scorti vix est torta panis,mulier autem viri pretiosam animam capit.
PROV|6|27|Numquid potest homo abscondere ignem in sinu suo,et vestimenta illius non ardebunt?
PROV|6|28|Aut ambulare super prunas,et non comburentur plantae eius?
PROV|6|29|Sic qui ingreditur ad mulierem proximi sui;non erit mundus, quicumque tetigerit eam.
PROV|6|30|Non contemptui erit fur, cum furatus fuerit,ut esurientem impleat animam.
PROV|6|31|Deprehensus quoque reddet septuplumet omnem substantiam domus suae tradet.
PROV|6|32|Qui autem adulter est cum muliere, vecors est;perdet animam suam, qui hoc fecerit.
PROV|6|33|Plagam et ignominiam congregat sibi,et opprobrium illius non delebitur.
PROV|6|34|Quia zelus est furor viri,et non parcet in die vindictae
PROV|6|35|nec accipiet personam tuam in piaculumnec suscipiet dona plurima.
PROV|7|1|Fili mi, custodi sermones meoset praecepta mea reconde tibi.
PROV|7|2|Serva mandata mea et vives,et legem meam quasi pupillam oculi tui.
PROV|7|3|Liga ea in digitis tuis,scribe illa in tabulis cordis tui.
PROV|7|4|Dic sapientiae: " Soror mea es "et prudentiam voca Amicam,
PROV|7|5|ut custodiat te a muliere extraneaet ab aliena, quae verba sua dulcia facit.
PROV|7|6|De fenestra enim domus meaeper cancellos prospexi
PROV|7|7|et video inter parvulos;considero inter filios vecordem iuvenem,
PROV|7|8|qui transit per plateam iuxta angulumet prope viam domus illius graditur
PROV|7|9|in obscuro advesperascente die,in mediis tenebris et caligine.
PROV|7|10|Et ecce, occurrit illi mulier ornatu meretricio,cauta corde, garrula et rebellans,
PROV|7|11|quietis impatiensnec valens in domo consistere pedibus suis:
PROV|7|12|nunc foris, nunc in plateiset iuxta angulos insidians.
PROV|7|13|Apprehensumque deosculatur iuvenemet procaci vultu blanditur dicens:
PROV|7|14|" Victimas pro salute vovi,hodie reddidi vota mea;
PROV|7|15|idcirco egressa sum in occursum tuumdesiderans te videre et repperi.
PROV|7|16|Stragulatis vestibus lectulum meum stravi,linteis pictis ex Aegypto;
PROV|7|17|aspersi cubile meum myrrhaet aloe et cinnamomo.
PROV|7|18|Veni, inebriemur voluptatibus,usque mane fruamur amoribus.
PROV|7|19|Non est enim vir in domo sua;abiit via longissima,
PROV|7|20|sacculum pecuniae secum tulit,in die plenae lunae reversurus est in domum suam ".
PROV|7|21|Irretivit eum multis sermonibuset blanditiis labiorum protraxit illum.
PROV|7|22|Stultus eam sequitur quasi bos ductus ad victimam,sicut irretitur vinculo cervus,
PROV|7|23|donec transfigat sagitta iecur eius;velut si avis festinet ad laqueumet nescit quod de periculo animae illius agitur.
PROV|7|24|Nunc ergo, fili mi, audi meet attende verbis oris mei.
PROV|7|25|Ne abstrahatur in viis illius mens tua,neque decipiaris semitis eius.
PROV|7|26|Multos enim vulneratos deiecit,et fortissimi quique interfecti sunt ab ea:
PROV|7|27|viae inferi domus eiuspenetrantes in interiora mortis.
PROV|8|1|Numquid non sapientia clamitat,et prudentia dat vocem suam?
PROV|8|2|In summis verticibussupra viam in mediis semitis stans,
PROV|8|3|iuxta portas ad introitum civitatis,in ipsis foribus conclamat:
PROV|8|4|" O viri, ad vos clamito,et vox mea ad filios hominum.
PROV|8|5|Intellegite, parvuli, astutiam;et insipientes, animadvertite.
PROV|8|6|Audite, quoniam de rebus magnis locutura sum,et aperientur labia mea, ut recta praedicent.
PROV|8|7|Veritatem meditabitur guttur meum,et labia mea detestabuntur impium.
PROV|8|8|Iusti sunt omnes sermones oris mei,non est in eis pravum quid neque perversum;
PROV|8|9|omnes recti sunt intellegentibuset aequi invenientibus scientiam.
PROV|8|10|Accipitc disciplinam meam et non pecuniam,doctrinam magis quam aurum electum.
PROV|8|11|Melior est enim sapientia gemmis,et omne desiderabile ei non potest comparari ".
PROV|8|12|Ego sapientia habito cum prudentiaet artem excogitandi invenio.
PROV|8|13|Timor Domini odisse malum;arrogantiam et superbiam et viam pravamet os bilingue detestor.
PROV|8|14|Meum est consilium et prudentia,mea est intellegentia, mea est fortitudo.
PROV|8|15|Per me reges regnant,et principes iusta decernunt;
PROV|8|16|per me duces imperant,et potentes decernunt iustitiam.
PROV|8|17|Ego diligentes me diligo;et, qui mane vigilant ad me, invenient me.
PROV|8|18|Mecum sunt divitiae et gloria,opes superbae et iustitia.
PROV|8|19|Melior est enim fructus meus auro et obryzo,et genimina mea argento electo.
PROV|8|20|In viis iustitiae ambulo,in medio semitarum iudicii,
PROV|8|21|ut ditem diligentes meet thesauros eorum repleam.
PROV|8|22|Dominus possedit me in initio viarum suarum,antequam quidquam faceret a principio;
PROV|8|23|ab aeterno ordinata sumet ex antiquis, antequam terra fieret.
PROV|8|24|Nondum erant abyssi, et ego iam concepta eram,necdum fontes graves aquis,
PROV|8|25|priusquam montes demergerentur,ante colles ego parturiebar.
PROV|8|26|Adhuc terram non fecerat et camposet initium glebae orbis terrae.
PROV|8|27|Quando praeparabat caelos, aderam,quando certa lege et gyro vallabat abyssos,
PROV|8|28|quando nubes firmabat sursum,et praevaluerunt fontes abyssi,
PROV|8|29|quando circumdabat mari terminum suumet aquis, ne transirent fines suos,quando iecit fundamenta terrae,
PROV|8|30|cum eo eram ut artifex:delectatio eius per singulos dies,ludens coram eo omni tempore,
PROV|8|31|ludens in orbe terrarum,et deliciae meae esse cum filiis hominum.
PROV|8|32|Nunc ergo, filii, audite me:beati, qui custodiunt vias meas;
PROV|8|33|audite disciplinam et estote sapienteset nolite abicere eam.
PROV|8|34|Beatus homo, qui audit meet qui vigilat ad fores meas cotidieet observat ad postes ostii mei.
PROV|8|35|Qui me invenerit, inveniet vitamet hauriet delicias a Domino.
PROV|8|36|Qui autem in me peccaverit, laedet animam suam:omnes, qui me oderunt, diligunt mortem.
PROV|9|1|Sapientia aedificavit sibi domum,excidit columnas septem;
PROV|9|2|immolavit victimas suas, miscuit vinumet proposuit mensam suam.
PROV|9|3|Misit ancillas suas, ut vocarentad arcem et ad excelsa civitatis:
PROV|9|4|" Si quis est parvulus, veniat ad me ".Et vecordi locuta est:
PROV|9|5|" Venite, comedite panem meumet bibite vinum, quod miscui vobis;
PROV|9|6|relinquite infantiam et viviteet ambulate per vias prudentiae ".
PROV|9|7|Qui erudit derisorem, ipse iniuriam sibi facit;et, qui arguit impium, sibi maculam generat.
PROV|9|8|Noli arguere derisorem, ne oderit te;argue sapientem, et diliget te.
PROV|9|9|Da sapienti, et sapientior fiet;doce iustum, et addet doctrinam.
PROV|9|10|Principium sapientiae timor Domini,et scientia Sancti est prudentia.
PROV|9|11|Per me enim multiplicabuntur dies tui,et addentur tibi anni vitae.
PROV|9|12|Si sapiens fueris, tibimetipsi eris;si autem illusor, solus portabis malum.
PROV|9|13|Mulier stulta est clamosa,fatua et nihil sciens;
PROV|9|14|sedit in foribus domus suaesuper sellam in excelsis urbis,
PROV|9|15|ut vocaret transeuntes per viamet pergentes itinere suo:
PROV|9|16|" Qui est parvulus, declinet ad me ".Et vecordi locuta est:
PROV|9|17|" Aquae furtivae dulciores sunt,et panis in abscondito suavior ".
PROV|9|18|Et ignoravit quod ibi sint umbrae,et in profundis inferni convivae eius.
PROV|10|1|Parabolae Salomonis.Filius sapiens laetificat pa trem,filius vero stultus maestitia est matris suae.
PROV|10|2|Nil proderunt thesauri impietatis,iustitia vero liberabit a morte.
PROV|10|3|Non affliget Dominus fame animam iustiet cupiditatem impiorum subvertet.
PROV|10|4|Egestatem operata est manus remissa,manus autem fortium divitias parat.
PROV|10|5|Qui congregat in messe, filius sapiens est;qui autem stertit aestate, filius confusionis.
PROV|10|6|Benedictiones Domini super caput iusti,os autem impiorum operit violentiam.
PROV|10|7|Memoria iusti in benedictione erit,et nomen impiorum putrescet.
PROV|10|8|Sapiens corde praecepta suscipit,et stultus labiis corruet.
PROV|10|9|Qui ambulat simpliciter, ambulat confidenter;qui autem depravat vias suas, manifestus erit.
PROV|10|10|Qui annuit oculo, dabit dolorem,et stultus labiis corruet.
PROV|10|11|Vena vitae os iusti,et os impiorum operit violentiam.
PROV|10|12|Odium suscitat rixas,et universa delicta operit caritas.
PROV|10|13|In labiis sapientis invenitur sapientia,et virga in dorso eius, qui indiget corde.
PROV|10|14|Sapientes recondunt scientiam,os autem stulti ruinae proximum est.
PROV|10|15|Substantia divitis urbs fortitudinis eius,ruina pauperum egestas eorum.
PROV|10|16|Opus iusti ad vitam,fructus autem impii ad peccatum.
PROV|10|17|Graditur ad vitam, qui custodit disciplinam;qui autem increpationes relinquit, errat.
PROV|10|18|Abscondunt odium labia mendacia;qui profert contumeliam, insipiens est.
PROV|10|19|In multiloquio non deerit peccatum;qui autem moderatur labia sua, prudentissimus est.
PROV|10|20|Argentum electum lingua iusti,cor autem impiorum pro nihilo.
PROV|10|21|Labia iusti erudiunt plurimos;qui autem indocti sunt, in cordis egestate morientur.
PROV|10|22|Benedictio Domini divites facit,nec addet ei labor quidquam.
PROV|10|23|Quasi per risum stultus operatur scelus,sapientia autem est viro prudentiae.
PROV|10|24|Quod timet impius, veniet super eum;desiderium suum iustis dabitur.
PROV|10|25|Quasi tempestas transiens non erit impius,iustus autem quasi fundamentum sempiternum.
PROV|10|26|Sicut acetum dentibus et fumus oculis,sic piger his, qui miserunt eum.
PROV|10|27|Timor Domini apponet dies,et anni impiorum breviabuntur.
PROV|10|28|Exspectatio iustorum laetitia,spes autem impiorum peribit.
PROV|10|29|Fortitudo simplici via Dominiet ruina his, qui operantur malum.
PROV|10|30|Iustus in aeternum non commovebitur,impii autem non habitabunt super terram.
PROV|10|31|Os iusti germinabit sapientiam,lingua prava abscindetur.
PROV|10|32|Labia iusti considerant placita,et os impiorum perversa.
PROV|11|1|Statera dolosa abominatio est apud Dominum,et pondus aequum voluntas eius.
PROV|11|2|Venit superbia, veniet et contumelia;apud humiles autem sapientia.
PROV|11|3|Simplicitas iustorum diriget eos,et supplantatio perversorum vastabit illos.
PROV|11|4|Non proderunt divitiae in die ultionis,iustitia autem liberabit a morte.
PROV|11|5|Iustitia simplicis diriget viam eius,et in impietate sua corruet impius.
PROV|11|6|Iustitia rectorum liberabit eos,et in insidiis suis capientur iniqui.
PROV|11|7|Mortuo homine impio, nulla erit ultra spes;et exspectatio divitiarum peribit.
PROV|11|8|Iustus de angustia liberatus est,et tradetur impius pro eo.
PROV|11|9|Simulator ore decipit amicum suum,iusti autem liberabuntur scientia.
PROV|11|10|In bonis iustorum exsultabit civitas,et in perditione impiorum erit laudatio.
PROV|11|11|Benedictione iustorum exaltabitur civitaset ore impiorum subvertetur.
PROV|11|12|Qui despicit amicum suum, indigens corde est,vir autem prudens tacebit.
PROV|11|13|Qui ambulat susurrans, revelat arcana;qui autem fidelis est animi, celat commissum.
PROV|11|14|Ubi non adsunt dispositiones, populus corruet;salus autem, ubi multa consilia.
PROV|11|15|Affligetur malo, qui fidem facit pro extraneo;qui autem odit sponsores, securus erit.
PROV|11|16|Mulier gratiosa inveniet gloriam,et robusti habebunt divitias.
PROV|11|17|Benefacit animae suae vir misericors;qui autem crudelis est, carnem suam affligit.
PROV|11|18|Impius facit opus fallax,seminanti autem iustitiam merces fidelis.
PROV|11|19|Firmus in iustitia praeparat vitam,et sectator malorum mortem.
PROV|11|20|Abominabile Domino cor pravum,et voluntas eius in iis, qui simpliciter ambulant.
PROV|11|21|Manus in manu, non erit impunitus malus,semen autem iustorum salvabitur.
PROV|11|22|Circulus aureus in naribus suismulier pulchra et fatua.
PROV|11|23|Desiderium iustorum omne bonum est,praestolatio impiorum furor.
PROV|11|24|Alii dividunt propria et ditiores fiunt,alii parciores iusto semper in egestate sunt.
PROV|11|25|Anima, quae benedicit, impinguabitur;et, qui inebriat, ipse quoque inebriatur.
PROV|11|26|Qui abscondit frumenta, maledicetur in populis,benedictio autem super caput vendentium.
PROV|11|27|Qui instanter quaerit bonum, quaerit beneplacitum;qui autem investigator malorum est, haec advenient ei.
PROV|11|28|Qui confidit in divitiis suis, corruet,iusti autem quasi virens folium germinabunt.
PROV|11|29|Qui conturbat domum suam, possidebit ventos;et, qui stultus est, serviet sapienti.
PROV|11|30|Fructus iusti lignum vitae;et suscipit animas, qui sapiens est.
PROV|11|31|Si iustus in terra rependitur,quanto magis impius et peccator.
PROV|12|1|Qui diligit disciplinam, diligit scientiam;qui autem odit increpationes, insipiens est.
PROV|12|2|Qui bonus est, hauriet gratiam a Domino,virum autem versutum ipse condemnabit.
PROV|12|3|Non roborabitur homo ex impietate,et radix iustorum non commovebitur.
PROV|12|4|Mulier diligens corona est viro suo,et quasi putredo in ossibus eius, quae est inhonesta.
PROV|12|5|Cogitationes iustorum iudicia,et consilia impiorum fraudulentia.
PROV|12|6|Verba impiorum insidiantur sanguini,os iustorum liberabit eos.
PROV|12|7|Subvertuntur impii et iam non sunt,domus autem iustorum permanebit.
PROV|12|8|Ad doctrinam suam laudabitur vir;qui autem perversus corde est, patebit contemptui.
PROV|12|9|Melior est pauper, qui ministrat sibi,quam gloriosus et indigens pane.
PROV|12|10|Curat iustus iumentorum suorum animas,viscera autem impiorum crudelia.
PROV|12|11|Qui operatur terram suam, satiabitur panibus;qui autem sectatur vana, vecors est.
PROV|12|12|Desiderat impius laqueum pessimorum,radix autem iustorum proficiet.
PROV|12|13|Propter peccata labiorum irretitur malus,effugiet autem iustus de angustia.
PROV|12|14|De fructu oris sui unusquisque replebitur bonis,et iuxta opera manuum suarum retribuetur ei.
PROV|12|15|Via stulti recta in oculis eius;qui autem sapiens est, audit consilia.
PROV|12|16|Fatuus statim indicat iram suam,dissimulat autem iniuriam callidus.
PROV|12|17|Qui spirat veritatem, index iustitiae est,testis autem mendax, fraudulentiae.
PROV|12|18|Est qui temere loquitur et quasi gladio pungit,lingua autem sapientium sanitas est.
PROV|12|19|Labium veritatis firmum erit in perpetuum,ad momentum autem lingua mendacii.
PROV|12|20|Dolus in corde cogitantium mala;qui autem pacis ineunt consilia, sequitur eos gaudium.
PROV|12|21|Nulla calamitas obveniet iusto,impii autem replebuntur malo.
PROV|12|22|Abominatio est Domino labia mendacia,qui autem fideliter agunt, placent ei.
PROV|12|23|Homo versutus celat scientiam,et cor insipientium provocat stultitiam.
PROV|12|24|Manus fortium dominabitur,quae autem remissa est, tributis serviet.
PROV|12|25|Maeror in corde viri humiliabit illum,et sermo bonus laetificabit eum.
PROV|12|26|In rectum ducit amicum iustus,iter autem impiorum decipiet eos.
PROV|12|27|Non assabit ignavia praedam suam,sed substantia pretiosa erit viro industrio.
PROV|12|28|In semita iustitiae vita,est autem etiam iter apertum ad mortem.
PROV|13|1|Filius sapiens disciplina patris;qui autem illusor est, non audit, cum arguitur.
PROV|13|2|De fructu oris sui homo satiabitur bonis,anima autem praevaricatorum violentia.
PROV|13|3|Qui custodit os suum, custodit animam suam;qui autem incautus est eloquio, ruina est ei.
PROV|13|4|Vult et non habet piger,anima autem operantium impinguabitur.
PROV|13|5|Verbum mendax iustus detestabitur,impius autem confundit et dehonestat.
PROV|13|6|Iustitia custodit innocentem in via,impietas autem peccatorem supplantat.
PROV|13|7|Est qui quasi dives habetur, cum nihil habeat;et est qui quasi pauper, cum in multis divitiis sit.
PROV|13|8|Redemptio animae viri divitiae suae;qui autem pauper est, increpationem non sustinet.
PROV|13|9|Lux iustorum laetificat,lucerna autem impiorum exstinguetur.
PROV|13|10|Inter superbos tantum iurgia sunt,et apud humiles sapientia.
PROV|13|11|Substantia festinata minuetur;qui autem colligit manu, multiplicat.
PROV|13|12|Spes, quae differtur, affligit animam,lignum vitae desiderium veniens.
PROV|13|13|Qui contemnit verbum, ipse se obligat;qui autem timet praeceptum, retribuetur ei.
PROV|13|14|Lex sapientis fons vitae,ut declinet a laqueis mortis.
PROV|13|15|Intellegentia bona dabit gratiam,in itinere infidelium vorago.
PROV|13|16|Omnis astutus agit cum consilio;qui autem fatuus est, aperit stultitiam.
PROV|13|17|Nuntius impius cadet in malum,legatus autem fidelis sanitas.
PROV|13|18|Egestas et ignominia ei, qui deserit disciplinam;qui autem acquiescit arguenti, glorificabitur.
PROV|13|19|Desiderium, si compleatur, delectat animam;detestantur stulti fugere mala.
PROV|13|20|Qui cum sapientibus graditur, sapiens erit;amicus stultorum malus efficietur.
PROV|13|21|Peccatores persequitur malum,et iustis retribuentur bona.
PROV|13|22|Bonus relinquit heredes filios et nepotes;et custoditur iusto substantia peccatoris.
PROV|13|23|Multi cibi in novalibus pauperum,et est qui perit, deficiente iudicio.
PROV|13|24|Qui parcit virgae, odit filium suum;qui autem diligit illum, instanter erudit.
PROV|13|25|Iustus comedit et replet animam suam,venter autem impiorum insaturabilis.
PROV|14|1|Sapientia mulierum aedificat domum suam,insipientia eam manibus destruet.
PROV|14|2|Ambulans recto itinere timet Deum;despicit illum, qui infami graditur via.
PROV|14|3|In ore stulti virga superbiae,labia autem sapientium custodiunt eos.
PROV|14|4|Ubi non sunt boves, praesepe vacuum est;plurimae autem segetes in fortitudine bovis.
PROV|14|5|Testis fidelis non mentitur,profert autem mendacium dolosus testis.
PROV|14|6|Quaerit derisor sapientiam et non invenit;doctrina prudentibus facilis.
PROV|14|7|Cede coram viro stulto,quia nescies labia prudentiae.
PROV|14|8|Sapientia callidi est intellegere viam suam,et imprudentia stultorum errans.
PROV|14|9|Stulti parvipendent peccatum,et inter iustos morabitur gratia.
PROV|14|10|Cor novit amaritudinem animae suae,in gaudio eius non miscebitur extraneus.
PROV|14|11|Domus impiorum delebitur,tabernacula vero iustorum germinabunt.
PROV|14|12|Est via, quae videtur homini recta,novissima autem eius deducunt ad mortem.
PROV|14|13|Etiam in risu cor dolore miscebitur,et extrema gaudii luctus occupat.
PROV|14|14|Viis suis replebitur stultus,et super eum erit vir bonus.
PROV|14|15|Simplex credit omni verbo,astutus considerat gressus suos.
PROV|14|16|Sapiens timet et declinat a malo,stultus transilit et confidit.
PROV|14|17|Impatiens operabitur stultitiam,et vir versutus odiosus est.
PROV|14|18|Possidebunt simplices stultitiam,et astuti coronabuntur scientia.
PROV|14|19|Procumbunt mali ante bonos,et impii ante portas iustorum.
PROV|14|20|Etiam proximo suo pauper odiosus erit,amici vero divitum multi.
PROV|14|21|Qui despicit proximum suum, peccat;qui autem miseretur pauperis, beatus erit.
PROV|14|22|Nonne errant, qui operantur malum?Misericordia et veritas iis, qui praeparant bona.
PROV|14|23|In omni labore erit abundantia;verbum autem labiorum tendit tantummodo ad egestatem.
PROV|14|24|Corona sapientium divitiae eorum,fatuitas stultorum fatuitas est.
PROV|14|25|Liberat animas testis fidelis,et profert mendacia versipellis.
PROV|14|26|In timore Domini fiducia fortis,et filiis eius erit spes.
PROV|14|27|Timor Domini fons vitae,declinans a laqueis mortis.
PROV|14|28|In multitudine populi dignitas regis,et in paucitate plebis ruina principis.
PROV|14|29|Qui patiens est, multa gubernatur prudentia;qui autem impatiens est, exaltat stultitiam.
PROV|14|30|Vita carnium sanitas cordis,putredo ossium invidia.
PROV|14|31|Qui calumniatur egentem, exprobrat Factori eius;honorat autem eum, qui miseretur pauperis.
PROV|14|32|In malitia sua impelletur impius,sperat autem iustus in integritate sua.
PROV|14|33|In corde prudentis requiescit sapientia,at in medio stultorum agnoscetur?
PROV|14|34|Iustitia elevat gentem,vituperium autem populorum est peccatum.
PROV|14|35|Acceptus est regi minister intellegens,et iracundia ei, qui turpiter agit.
PROV|15|1|Responsio mollis frangit iram,sermo durus suscitat furorem.
PROV|15|2|Lingua sapientium stillat scientiam,os fatuorum ebullit stultitiam.
PROV|15|3|In omni loco oculi Dominicontemplantur malos et bonos.
PROV|15|4|Lingua placabilis lignum vitae,sed obliquitas in ea conteret spiritum.
PROV|15|5|Stultus irridet disciplinam patris sui;qui autem custodit increpationes, astutior fiet.
PROV|15|6|In domo iusti divitiae plurimae,et in fructibus impii conturbatio.
PROV|15|7|Labia sapientium disseminabunt scientiam;cor stultorum non rectum erit.
PROV|15|8|Victimae impiorum abominabiles Domino;vota iustorum grata sunt ei.
PROV|15|9|Abominatio est Domino via impii;qui sequitur iustitiam, diligetur.
PROV|15|10|Admonitio mala deserenti viam;qui increpationes odit, morietur.
PROV|15|11|Infernus et Perditio coram Domino,quanto magis corda filiorum hominum!
PROV|15|12|Non amat derisor eum, qui se corripit,nec ad sapientes graditur.
PROV|15|13|Cor gaudens exhilarat faciem,in maerore animi deicitur spiritus.
PROV|15|14|Cor sapientis quaerit doctrinam,et os stultorum pascitur stultitia.
PROV|15|15|Omnes dies pauperis mali;hilaris autem corde quasi iuge convivium.
PROV|15|16|Melius est parum cum timore Dominiquam thesauri magni cum sollicitudine.
PROV|15|17|Melius est demensum holerum cum caritatequam vitulus saginatus cum odio.
PROV|15|18|Vir iracundus provocat rixas;qui patiens est, mitigat lites.
PROV|15|19|Iter pigrorum quasi saepes spinarum,via sollertium complanata.
PROV|15|20|Filius sapiens laetificat patrem,et stultus homo despicit matrem suam.
PROV|15|21|Stultitia gaudium sensu carenti;et vir prudens dirigit gressus suos.
PROV|15|22|Dissipantur cogitationes, ubi non est consilium;ubi vero sunt plures consiliarii, confirmantur.
PROV|15|23|Laetatur homo in responsione oris sui,et sermo opportunus est optimus.
PROV|15|24|Semita vitae sursum est viro erudito,ut declinet de inferno deorsum.
PROV|15|25|Domum superborum demolietur Dominuset firmos faciet terminos viduae.
PROV|15|26|Abominatio Domini cogitationes malae,et purus sermo pulcherrimus.
PROV|15|27|Conturbat domum suam, qui sectatur avaritiam;qui autem odit munera, vivet.
PROV|15|28|Mens iusti meditatur, ut respondeat;os impiorum redundat malis.
PROV|15|29|Longe est Dominus ab impiiset orationes iustorum exaudiet.
PROV|15|30|Lux oculorum laetificat animam,fama bona impinguat ossa.
PROV|15|31|Auris, quae audit increpationes vitae,in medio sapientium commorabitur.
PROV|15|32|Qui abicit disciplinam, despicit animam suam;qui autem acquiescit increpationibus, possessor est cordis.
PROV|15|33|Timor Domini disciplina sapientiae,et gloriam praecedit humilitas.
PROV|16|1|Hominis est animum praeparare,et Domini est responsio linguae.
PROV|16|2|Omnes viae hominis purae sunt oculis eius,spirituum ponderator est Dominus.
PROV|16|3|Revela Domino opera tua,et dirigentur cogitationes tuae.
PROV|16|4|Universa secundum proprium finem operatus est Dominus;impium quoque ad diem malum.
PROV|16|5|Abominatio Domini est omnis arrogans;manus in manu, non erit innocens.
PROV|16|6|Misericordia et veritate redimitur iniquitas,et in timore Domini declinatur a malo.
PROV|16|7|Cum placuerint Domino viae hominis,inimicos quoque eius convertet ad pacem.
PROV|16|8|Melius est parum cum iustitiaquam multi fructus sine aequitate.
PROV|16|9|Cor hominis disponit viam suam,sed Domini est dirigere gressus eius.
PROV|16|10|Divinatio in labiis regis,in iudicio non errabit os eius.
PROV|16|11|Pondus et statera iusta Domini sunt,et opera eius omnes lapides sacculi.
PROV|16|12|Abominantur reges agere impie,quoniam iustitia firmatur solium.
PROV|16|13|Voluntas regum labia iusta;qui recta loquitur, diligetur.
PROV|16|14|Indignatio regis nuntii mortis,et vir sapiens placabit eam.
PROV|16|15|In lumine vultus regis vita,et voluntas eius quasi imber serotinus.
PROV|16|16|Possidere sapientiam quanto melius est auro;et acquirere prudentiam pretiosius est argento.
PROV|16|17|Semita iustorum declinare a malo;custos animae suae, qui servat viam suam.
PROV|16|18|Contritionem praecedit superbia,et ante ruinam exaltatio spiritus.
PROV|16|19|Melius est humiliari cum mitibusquam dividere spolia cum superbis.
PROV|16|20|Eruditus in verbo reperiet bona;et, qui sperat in Domino, beatus est.
PROV|16|21|Qui sapiens est corde, appellabitur prudens;et dulcedo labiorum addet doctrinam.
PROV|16|22|Fons vitae eruditio possidentis;poena stultorum stultitia.
PROV|16|23|Cor sapientis erudiet os eiuset labiis eius addet doctrinam.
PROV|16|24|Favus mellis composita verba,dulcedo animae et sanitas ossium.
PROV|16|25|Est via, quae videtur homini recta,et novissima eius ducunt ad mortem.
PROV|16|26|Anima laborantis laborat sibi,quia compulit eum os suum.
PROV|16|27|Vir impius fodit malum,et in labiis eius quasi ignis ardens.
PROV|16|28|Homo perversus suscitat lites,et mussitator separat familiares.
PROV|16|29|Vir iniquus lactat amicum suumet ducit eum per viam non bonam.
PROV|16|30|Qui attonitis oculis cogitat prava,comprimens labia sua perficit malum.
PROV|16|31|Corona dignitatis canities,quae in viis iustitiae reperietur.
PROV|16|32|Melior est patiens viro forti,et, qui dominatur animo suo, expugnatore urbium.
PROV|16|33|Sortes mittuntur in sinum,sed a Domino temperantur.
PROV|17|1|Melior est buccella sicca cum pacequam domus plena victimis cum iurgio.
PROV|17|2|Servus sapiens dominabitur filiis inhonestiset inter fratres hereditatem dividet.
PROV|17|3|Sicut igne probatur argentum et aurum camino,ita corda probat Dominus.
PROV|17|4|Malus oboedit labio iniquo,et fallax obtemperat linguae mendaci.
PROV|17|5|Qui despicit pauperem, exprobrat Factori eius;et, qui in ruina laetatur alterius, non erit impunitus.
PROV|17|6|Corona senum filii filiorum,et gloria filiorum patres eorum.
PROV|17|7|Non decent stultum verba composita,nec principem labium mentiens.
PROV|17|8|Gemma gratissima munus in oculis domini eius;quocumque se verterit, prospere aget.
PROV|17|9|Qui celat delictum, quaerit amicitias;qui sermone repetit, separat foederatos.
PROV|17|10|Plus proficit correptio apud prudentemquam centum plagae apud stultum.
PROV|17|11|Semper iurgia quaerit malus;angelus autem crudelis mittetur contra eum.
PROV|17|12|Expedit magis ursae occurrere, raptis fetibus,quam fatuo confidenti in stultitia sua.
PROV|17|13|Qui reddit mala pro bonis,non recedet malum de domo eius.
PROV|17|14|Aquarum proruptio initium est iurgiorum;et, antequam exacerbetur contentio, desere.
PROV|17|15|Qui iustificat impium et qui condemnat iustum,abominabilis est uterque apud Dominum.
PROV|17|16|Ad quid pretium in manu stulti?Ad emendam sapientiam, cum careat corde?
PROV|17|17|Omni tempore diligit, qui amicus est,et frater ad angustiam natus est.
PROV|17|18|Stultus homo iungit manus,cum spoponderit pro amico suo.
PROV|17|19|Qui diligit delictum, diligit rixas;et, qui exaltat ostium, quaerit effracturam.
PROV|17|20|Qui perversi cordis est, non inveniet bonum;et, qui vertit linguam, incidet in malum.
PROV|17|21|Qui generat stultum, maerorem generat sibi,sed nec pater in fatuo laetabitur.
PROV|17|22|Animus gaudens aetatem floridam facit,spiritus tristis exsiccat ossa.
PROV|17|23|Munera de sinu impius accipit,ut pervertat semitas iudicii.
PROV|17|24|In facie prudentis lucet sapientia,oculi stultorum in finibus terrae.
PROV|17|25|Ira patris filius stultuset dolor matris, quae genuit eum.
PROV|17|26|Non est bonum multam inferre iustonec percutere principem contra rectitudinem.
PROV|17|27|Qui moderatur sermones suos, novit scientiam,et lenis spiritu est vir prudens.
PROV|17|28|Stultus quoque, si tacuerit, sapiens reputabituret, si compresserit labia sua, intellegens.
PROV|18|1|Occasiones quaerit, qui vult recedere ab amico;omni consilio exacerbatur.
PROV|18|2|Non delectatur stultus prudentiased in revelatione cordis sui.
PROV|18|3|Cum venerit impius, veniet et contemptio,et cum ignominia opprobrium.
PROV|18|4|Aqua profunda verba ex ore viri,et torrens redundans fons sapientiae.
PROV|18|5|Accipere personam impii non est bonum,ut declines iustum in iudicio.
PROV|18|6|Labia stulti miscent se rixis,et os eius plagas provocat.
PROV|18|7|Os stulti ruina eius,et labia ipsius laqueus animae eius.
PROV|18|8|Verba susurronis quasi dulcia,et ipsa perveniunt usque ad interiora ventris.
PROV|18|9|Qui mollis et dissolutus est in opere suo,frater est viri dissipantis.
PROV|18|10|Turris fortissima nomen Domini;ad ipsum currit iustus et exaltabitur.
PROV|18|11|Substantia divitis urbs roboris eiuset quasi murus excelsus in cogitatione eius.
PROV|18|12|Antequam conteratur, exaltatur cor hominis;et, antequam glorificetur, humiliatur.
PROV|18|13|Qui prius respondet quam audiat,stultitia est ei et contumelia.
PROV|18|14|Spiritus viri sustentat imbecillitatem suam;spiritum vero confractum, quis poterit sustinere?
PROV|18|15|Cor prudens possidebit scientiam,et auris sapientium quaerit doctrinam.
PROV|18|16|Donum hominis dilatat viam eiuset ante principes deducit eum.
PROV|18|17|Qui prior in contentione loquitur, putatur iustus;venit amicus eius et arguet eum.
PROV|18|18|Lites comprimit sorset inter potentes quoque diiudicat.
PROV|18|19|Frater, qui offenditur, durior est civitate firma,et lites quasi vectes urbium.
PROV|18|20|De fructu oris viri replebitur venter eius,et genimina labiorum ipsius saturabunt eum.
PROV|18|21|Mors et vita in manu linguae;qui diligunt eam, comedent fructus eius.
PROV|18|22|Qui invenit mulierem bonam, invenit bonumet hausit gratiam a Domino.
PROV|18|23|Cum obsecrationibus loquetur pauper,et dives effabitur rigide.
PROV|18|24|Vir cum amicis concuti potest,sed est amicus, qui adhaereat magis quam frater.
PROV|19|1|Melior est pauper, qui ambulat in simplicitate sua,quam qui torquet labia et est insipiens.
PROV|19|2|Ubi non est scientia animae, non est bonum;et, qui festinus est pedibus, offendit.
PROV|19|3|Stultitia hominis supplantat gressus eius,et contra Deum fervet animo suo.
PROV|19|4|Divitiae addunt amicos plurimos;pauper autem ab amico suo separatur.
PROV|19|5|Testis falsus non erit impunitus;et, qui mendacia loquitur, non effugiet.
PROV|19|6|Multi blandiuntur faciei potentis,et omnes amici sunt dona tribuenti.
PROV|19|7|Omnes fratres hominis pauperis oderunt eum,insu7per et amici procul recesserunt ab eo;qui tantum verba sectatur, nihil habebit.
PROV|19|8|Qui autem possessor est mentis, diligit animam suam,et custos prudentiae inveniet bona.
PROV|19|9|Falsus testis non erit impunitus;et, qui loquitur mendacia, peribit.
PROV|19|10|Non decent stultum deliciae,nec servum dominari principibus.
PROV|19|11|Doctrina viri mitigat iram eius,et gloria eius est iniqua praetergredi.
PROV|19|12|Sicut fremitus leonis ita et regis ira,et sicut ros super herbam ita et gratia eius.
PROV|19|13|Calamitas patris filius stultus;et tecta iugiter perstillantia litigiosa mulier.
PROV|19|14|Domus et divitiae hereditas patrum,a Domino autem uxor prudens.
PROV|19|15|Pigredo immittit soporem,et anima dissoluta esuriet.
PROV|19|16|Qui custodit mandatum, custodit animam suam;qui autem neglegit viam suam, mortificabitur.
PROV|19|17|Feneratur Domino, qui miseretur pauperis,et vicissitudinem suam reddet ei.
PROV|19|18|Erudi filium tuum, dum spes est;ad interfectionem autem eius ne ponas animam tuam.
PROV|19|19|Qui impatiens est, sustinebit multam;et, si eum abripere vis, aliud appones.
PROV|19|20|Audi consilium et suscipe disciplinam,ut sis sapiens in novissimis tuis.
PROV|19|21|Multae cogitationes in corde viri,voluntas autem Domini permanebit.
PROV|19|22|Desiderabile in homine est misericordia eius;et melior est pauper quam vir mendax.
PROV|19|23|Timor Domini ad vitam,et in plenitudine commorabitur absque visitatione mali.
PROV|19|24|Abscondit piger manum suam in catinonec ad os suum applicat eam.
PROV|19|25|Derisore flagellato vel parvulus sapientior erit;si autem corripueris sapientem, intelleget disciplinam.
PROV|19|26|Qui affligit patrem et fugat matrem,filius inhonestus et ignominiosus.
PROV|19|27|Acquiesce, fili, ut audias doctrinamnec erres a sermonibus scientiae.
PROV|19|28|Testis iniquus deridet iudicium,et os impiorum devorat iniquitatem.
PROV|19|29|Paratae sunt derisoribus virgae,et plagae stultorum corporibus.
PROV|20|1|Luxuriosa res vinum, et tumultuosa sicera;quicumque his delectatur, non erit sapiens.
PROV|20|2|Sicut rugitus leonis ita et terror regis:qui provocat eum, peccat in animam suam.
PROV|20|3|Honor est homini separari a contentionibus;omnes autem stulti miscentur contumeliis.
PROV|20|4|Propter frigus piger arare noluit;mendicabit ergo aestate, et non dabitur illi.
PROV|20|5|Sicut aqua profunda consilium in corde viri,sed homo sapiens exhauriet illud.
PROV|20|6|Multi homines misericordes vocantur;virum autem fidelem quis inveniet?
PROV|20|7|Iustus, qui ambulat in simplicitate sua,beatos post se filios derelinquet.
PROV|20|8|Rex, qui sedet in solio iudicii,dissipat omne malum intuitu suo.
PROV|20|9|Quis potest dicere: " Mundavi cor meum,purus sum a peccato "?
PROV|20|10|Pondus et pondus, mensura et mensura,utrumque abominabile est apud Dominum.
PROV|20|11|Ex studiis suis intellegitur puer,si munda et recta sint opera eius.
PROV|20|12|Aurem audientem et oculum videntem,Dominus fecit utrumque.
PROV|20|13|Noli diligere somnum, ne te egestas opprimat;aperi oculos tuos et saturare panibus.
PROV|20|14|" Malum est, malum est! " dicit omnis emptoret, cum recesserit, tunc gloriabitur.
PROV|20|15|Est aurum et multitudo gemmarumet vas pretiosum labia scientiae.
PROV|20|16|Tolle vestimentum eius, quia fideiussor exstitit alieni,et pro extraneis aufer pignus ab eo.
PROV|20|17|Suavis est homini panis mendacii,et postea implebitur os eius calculo.
PROV|20|18|Cogitationes consiliis firmantur,et dispensationibus tractanda sunt bella.
PROV|20|19|Ei, qui revelat mysteria et calumniaturet dilatat labia sua, ne commiscearis.
PROV|20|20|Qui maledicit patri suo et matri,exstinguetur lucerna eius in mediis tenebris.
PROV|20|21|Hereditas, ad quam festinatur in principio,in novissimo benedictione carebit.
PROV|20|22|Ne dicas: " Reddam malum ";exspecta Dominum, et liberabit te.
PROV|20|23|Abominatio est apud Dominum pondus et pondus;statera dolosa non est bona in oculis eius.
PROV|20|24|A Domino diriguntur gressus viri;quis autem hominum intellegere potest viam suam?
PROV|20|25|Laqueus est homini inconsulte dicere: " Sanctum! "et post vota retractare.
PROV|20|26|Ventilat impios rex sapienset incurvat super eos rotam.
PROV|20|27|Lucerna Domini spiraculum hominis,quae investigat omnia secreta ventris.
PROV|20|28|Misericordia et veritas custodiunt regem,et roboratur clementia thronus eius.
PROV|20|29|Ornamentum iuvenum fortitudo eorum,et honor senum canities.
PROV|20|30|Livor vulneris absterget mala,et plagae in secretioribus ventris.
PROV|21|1|Sicut rivi aquarum cor regis in manu Domini:quocumque voluerit, inclinabit illud.
PROV|21|2|Omnis via viri recta sibi videtur;appendit autem corda Dominus.
PROV|21|3|Facere misericordiam et iudiciummagis placet Domino quam victimae.
PROV|21|4|Exaltatio oculorum et dilatatio cordis,lucerna impiorum: peccatum.
PROV|21|5|Cogitationes sollertis semper in abundantiam;omnis autem festinus semper in egestate est.
PROV|21|6|Qui congregat thesauros lingua mendacii,vento impingetur ad laqueos mortis.
PROV|21|7|Violentia impiorum detrahet eos,quia noluerunt facere iudicium.
PROV|21|8|Perversa via viri aliena est;qui autem mundus est, rectum opus eius.
PROV|21|9|Melius est sedere in angulo domatisquam cum muliere litigiosa et in domo communi.
PROV|21|10|Anima impii desiderat malum;non miserebitur proximo suo.
PROV|21|11|Multato derisore sapientior erit parvulus;et, si instruatur sapiens, sumet scientiam.
PROV|21|12|Excogitat Iustus de domo impii,ut praecipitet impios in malum.
PROV|21|13|Qui obturat aurem suam ad clamorem pauperis,et ipse clamabit, et non exaudietur.
PROV|21|14|Munus absconditum exstinguit iras,et donum in sinu indignationem maximam.
PROV|21|15|Gaudium iusto est facere iudicium,et ruina operantibus iniquitatem.
PROV|21|16|Vir, qui erraverit a via prudentiae,in coetu umbrarum commorabitur.
PROV|21|17|Qui diligit convivia, in egestate erit;qui amat vinum et pinguia, non ditabitur.
PROV|21|18|Redemptio pro iusto impius,et pro rectis iniquus.
PROV|21|19|Melius est habitare in terra desertaquam cum muliere rixosa et iracunda.
PROV|21|20|Thesaurus desiderabilis et pinguis in habitaculo sapientis,et imprudens homo dissipabit illum.
PROV|21|21|Qui sequitur iustitiam et misericordiam,inveniet vitam et iustitiam et gloriam.
PROV|21|22|Civitatem fortium ascendit sapienset destruit robur fiduciae eius.
PROV|21|23|Qui custodit os suum et linguam suam,custodit ab angustiis animam suam.
PROV|21|24|Superbus et arrogans vocatur derisor,qui operatur in ira superbiae.
PROV|21|25|Desideria occidunt pigrum;noluerunt enim quidquam manus eius operari:
PROV|21|26|tota die concupiscit et desiderat;qui autem iustus est, tribuet et non parcit.
PROV|21|27|Hostiae impiorum abominabiles,eo magis quia offeruntur ex scelere.
PROV|21|28|Testis mendax peribit;vir oboediens loquetur in victoriam.
PROV|21|29|Vir impius obfirmat vultum suum;qui autem rectus est, corrigit viam suam.
PROV|21|30|Non est sapientia, non est prudentia,non est consilium contra Dominum.
PROV|21|31|Equus paratur ad diem belli,Dominus autem salutem tribuit.
PROV|22|1|Melius est nomen bonum quam divitiae multae,super argentum et aurum gratia bona.
PROV|22|2|Dives et pauper obviaverunt sibi:utriusque operator est Dominus.
PROV|22|3|Callidus vidit malum et abscondit se;simplices pertransierunt et afflicti sunt damno.
PROV|22|4|Praemium modestiae timor Domini,divitiae et gloria et vita.
PROV|22|5|Spinae et laquei in via perversi,custos autem animae suae longe recedit ab eis.
PROV|22|6|Institue adulescentem iuxta viam suam;etiam cum senuerit, non recedet ab ea.
PROV|22|7|Dives pauperibus imperat;et, qui accipit mutuum, servus est fenerantis.
PROV|22|8|Qui seminat iniquitatem, metet malaet virga irae suae consummabitur.
PROV|22|9|Qui bono oculo est, benedicetur,de panibus enim suis dedit pauperi.
PROV|22|10|Eice derisorem, et exibit cum eo iurgium;cessabuntque causae et contumeliae.
PROV|22|11|Qui diligit cordis munditiam,propter gratiam labiorum suorum habebit amicum regem.
PROV|22|12|Oculi Domini custodiunt scientiam,et supplantantur verba iniqui.
PROV|22|13|Dicit piger: " Leo est foris,in medio platearum occidendus sum ".
PROV|22|14|Fovea profunda os alienae;cui iratus est Dominus, incidet in eam.
PROV|22|15|Stultitia colligata est in corde pueri,et virga disciplinae fugabit eam.
PROV|22|16|Opprimis pauperem? Ipse augebit divitias suas.Donas ditiori? Ipse egebis.
PROV|22|17|Inclina aurem tuam et audi verba sapientium,appone autem cor ad doctrinam meam,
PROV|22|18|quia pulchra erunt, cum servaveris ea in ventre tuo,et redundabunt in labiis tuis.
PROV|22|19|Ut sit in Domino fiducia tua,ostendi ea tibi hodie.
PROV|22|20|Nonne descripsi ea tibi nudiustertiusin cogitationibus et scientia,
PROV|22|21|ut ostenderem tibi firmitatem verborum veritatis,ut respondeas illi, qui misit te?
PROV|22|22|Non facias violentiam pauperi, quia pauper est,neque conteras egenum in porta,
PROV|22|23|quia iudicabit Dominus causam eorum,et anima spoliabit spoliatores.
PROV|22|24|Noli esse amicus homini iracundoneque ambules cum viro furioso,
PROV|22|25|ne forte discas semitas eiuset sumas scandalum animae tuae.
PROV|22|26|Noli esse cum his, qui iungunt manus suaset qui vades se offerunt pro debitis:
PROV|22|27|si enim non habes unde restituas,quid causae est ut tollat lectum tuum subter te?
PROV|22|28|Ne transferas terminos antiquos,quos posuerunt patres tui.
PROV|22|29|Vidisti virum velocem in opere suo:coram regibus stabit nec erit ante ignobiles.
PROV|23|1|Quando sederis, ut comedas cum principe,diligenter attende, quae apposita sunt ante faciem tuam,
PROV|23|2|et statue cultrum in gutture tuo,si avidus es.
PROV|23|3|Ne desideres de cibis eius,quia est panis mendacii.
PROV|23|4|Noli laborare, ut diteris,sed in prudentia tua acquiesce.
PROV|23|5|Si erigas oculos tuos ad opes, iam non sunt;quia facient sibi pennas quasi aquilae et volabunt in caelum.
PROV|23|6|Ne comedas cum homine invidoet ne desideres cibos eius;
PROV|23|7|quoniam sicut aestimavit in animo suo,ita ipse est. Comede et bibe " dicet tibi,et mens eius non est tecum.
PROV|23|8|Buccellam, quam comederas, evomeset perdes pulchros sermones tuos.
PROV|23|9|In auribus insipientium ne loquaris,quia despicient doctrinam eloquii tui.
PROV|23|10|Ne attingas terminos viduaeet agrum pupillorum ne introeas:
PROV|23|11|redemptor enim illorum fortis est,et ipse iudicabit contra te causam illorum.
PROV|23|12|Introduc ad doctrinam cor tuumet aures tuas ad verba scientiae.
PROV|23|13|Noli subtrahere a puero disciplinam;si enim percusseris eum virga, non morietur:
PROV|23|14|tu virga percuties eumet animam eius de inferno liberabis.
PROV|23|15|Fili mi, si sapiens fuerit cor tuum,gaudebit tecum et cor meum,
PROV|23|16|et exsultabunt renes mei,cum locuta fuerint rectum labia tua.
PROV|23|17|Non aemuletur cor tuum peccatores,sed in timore Domini esto tota die,
PROV|23|18|quia est tibi posteritas,et praestolatio tua non auferetur.
PROV|23|19|Audi, fili mi, et esto sapienset dirige in via animum tuum.
PROV|23|20|Noli esse in conviviis potatorumnec in comissationibus carnis,
PROV|23|21|quia vacantes potibus et comissatores consumentur,et vestietur pannis dormitatio.
PROV|23|22|Audi patrem tuum, qui genuit te,et ne contemnas, cum senuerit mater tua.
PROV|23|23|Veritatem eme et noli vendere;sapientiam eme et doctrinam et intellegentiam.
PROV|23|24|Exsultat gaudio pater iusti;qui sapientem genuit, laetabitur in eo;
PROV|23|25|gaudeat pater tuus et mater tua,et exsultet, quae genuit te.
PROV|23|26|Praebe, fili mi, cor tuum mihi,et oculi tui vias meas custodiant.
PROV|23|27|Fovea enim profunda est meretrix,et puteus angustus aliena,
PROV|23|28|nam insidiatur ipsa in via quasi latroet iniquos in hominibus addet.
PROV|23|29|Cui " Vae "? Cui " Eheu "?Cui rixae? Cui querela?Cui sine causa vulnera? Cui suffusio oculorum?
PROV|23|30|His, qui commorantur in vinoet eunt, ut scrutentur mixtum.
PROV|23|31|Ne intuearis vinum, quando flavescit,cum splenduerit in calice color eius:ingreditur blande,
PROV|23|32|sed in novissimo mordebit ut coluberet sicut regulus vulnerat.
PROV|23|33|Oculi tui videbunt extranea,et cor tuum loquetur perversa;
PROV|23|34|et eris sicut dormiens in medio mariet quasi sopitus ad malum navis:
PROV|23|35|" Verberaverunt me, sed non dolui,percusserunt me, et ego non sensi;quando evigilabo et rursus illud requiram? ".
PROV|24|1|Ne aemuleris viros malosnec desideres esse cum eis,
PROV|24|2|quia rapinas meditatur mens eorum,et perniciem labia eorum loquuntur.
PROV|24|3|Sapientia aedificabitur domus,et prudentia roborabitur.
PROV|24|4|In doctrina replebuntur cellaria,universa substantia pretiosa et pulcherrima.
PROV|24|5|Vir sapiens fortis est,et vir doctus firmat robur.
PROV|24|6|Quia cum dispositione parabis tibi bellum,et erit salus, ubi multa consilia sunt.
PROV|24|7|Excelsa stulto sapientia,in porta non aperiet os suum.
PROV|24|8|Qui cogitat mala facere,vir perniciosus vocabitur.
PROV|24|9|Cogitatio stulti peccatum est,et abominatio hominum detractor.
PROV|24|10|Si fueris lassus in die angustiae,coartabitur fortitudo tua.
PROV|24|11|Erue eos, qui ducuntur ad mortem;et, qui trahuntur ad interitum, retine.
PROV|24|12|Si dixeris: " Nesciebamus hoc ";nonne qui ponderator est cordis, ipse intellegit,et servatorem animae tuae nihil fallitreddetque homini iuxta opera sua?
PROV|24|13|Comede, fili mi, mel, quia bonum estet favum dulcissimum gutturi tuo.
PROV|24|14|Sic, scito, est sapientia animae tuae;quam cum inveneris, erit tibi posteritas,et spes tua non peribit.
PROV|24|15|Ne insidieris, o nequam, domui iustineque vastes requiem eius.
PROV|24|16|Septies enim cadet iustus et resurget;impii autem corruent in malum.
PROV|24|17|Cum ceciderit inimicus tuus, ne gaudeas,et in ruina eius ne exsultet cor tuum,
PROV|24|18|ne forte videat Dominus, et displiceat eiet auferat ab eo iram suam.
PROV|24|19|Ne succendas ira in pessimosnec aemuleris impios,
PROV|24|20|quoniam non erit posteritas maligno,et lucerna impiorum exstinguetur.
PROV|24|21|Time Dominum, fili mi, et regemet cum nova sectantibus non commiscearis,
PROV|24|22|quoniam repente consurget perditio eorum,et ruinam utriusque quis novit?
PROV|24|23|Haec quoque sapientibus:Dignoscere personam in iudicio non est bonum.
PROV|24|24|Qui dicit impio: " Iustus es ",maledicent ei populi, et detestabuntur eum tribus.
PROV|24|25|Qui vero arguunt eum, laudabuntur,et super ipsos veniet benedictio boni.
PROV|24|26|Labia deosculatur,qui recta verba respondet.
PROV|24|27|Praepara foris opus tuumet diligenter exerce illud in agro tuo,ut postea aedifices domum tuam.
PROV|24|28|Ne sis testis frustra contra proximum tuumnec decipias quemquam labiis tuis.
PROV|24|29|Ne dicas: " Quomodo fecit mihi, sic faciam ei,reddam viro secundum opus suum ".
PROV|24|30|Per agrum hominis pigri transiviet per vineam viri sensu carentis:
PROV|24|31|et ecce totum repleverant urticae,et operuerant superficiem eius spinae,et maceria lapidum destructa erat;
PROV|24|32|quod cum vidissem, posui in corde meo,vidi, didici disciplinam:
PROV|24|33|" Parum dormies, modicum dormitabis,pauxillum manus conseres, ut quiescas,
PROV|24|34|et veniet tibi quasi cursor egestas,et mendicitas quasi vir armatus ".
PROV|25|1|Hae quoque parabolae Salomonis, quas transcripse runt viri Ezechiae regis Iudae.
PROV|25|2|Gloria Dei est celare verbum,et gloria regum investigare sermonem.
PROV|25|3|Caelum prae altitudine et terra prae profunditate,et cor regum inscrutabile.
PROV|25|4|Aufer scorias de argento,et egredietur vas pro argentario.
PROV|25|5|Aufer impium de conspectu regis,et firmabitur iustitia thronus eius.
PROV|25|6|Ne gloriosus appareas coram regeet in loco magnorum ne steteris.
PROV|25|7|Melius est enim ut dicatur tibi: " Ascende huc ",quam ut humilieris coram principe.
PROV|25|8|Quae viderunt oculi tui,ne proferas in iurgio cito,quoniam quid facies postea,cum dehonestaverit te amicus tuus?
PROV|25|9|Causam tuam tracta cum amico tuoet secretum extranei ne reveles,
PROV|25|10|ne forte insultet tibi, cum audierit,et contumelia tua revocari non poterit.
PROV|25|11|Mala aurea in ornatibus argenteis,verbum prolatum in tempore suo.
PROV|25|12|Inauris aurea et margaritum fulgenssapiens, qui arguit super aurem audientem.
PROV|25|13|Sicut frigus nivis in die messis,ita legatus fidelis ei, qui misit eum:animam ipsius recreat.
PROV|25|14|Nubes et ventus et pluviae non sequentesvir gloriosus et promissa non complens.
PROV|25|15|Patientia lenietur princeps,et lingua mollis confringet ossa.
PROV|25|16|Mel invenisti? Comede, quod sufficit tibi,ne forte satiatus evomas illud.
PROV|25|17|Subtrahe pedem tuum de domo proximi tui,ne quando satiatus oderit te.
PROV|25|18|Malleus et gladius et sagitta acutahomo, qui loquitur contra proximum suum falsum testimonium.
PROV|25|19|Dens putridus et pes vacillans,qui sperat super infideli in die angustiae.
PROV|25|20|Sicut exuens pallium in die frigoris,sicut acetum in nitro,qui cantat carmina cordi tristi.
PROV|25|21|Si esurierit inimicus tuus, ciba illum;si sitierit, pota illum:
PROV|25|22|prunas enim congregabis super caput eius,et Dominus reddet tibi.
PROV|25|23|Ventus aquilo parturit pluvias,et faciem tristem lingua detrahens.
PROV|25|24|Melius est sedere in angulo domatisquam cum muliere litigiosa et in domo communi.
PROV|25|25|Aqua frigida animae sitientiet nuntius bonus de terra longinqua.
PROV|25|26|Fons turbatus pede et vena corruptaiustus cadens coram impio.
PROV|25|27|Mel nimium comedere non est bonum,nec quaestus gloriae est gloria.
PROV|25|28|Urbs diruta et absque murovir, qui non potest cohibere spiritum suum.
PROV|26|1|Quomodo nix in aestate et pluvia in messe,sic indecens est stulto gloria.
PROV|26|2|Sicut avis ad alia transvolans et hirundo volitans,sic maledictum frustra prolatum non superveniet.
PROV|26|3|Flagellum equo et camus asinoet virga dorso stultorum.
PROV|26|4|Ne respondeas stulto iuxta stultitiam suam,ne tu quoque efficiaris ei similis;
PROV|26|5|responde stulto iuxta stultitiam suam,ne sibi sapiens esse videatur.
PROV|26|6|Amputat sibi pedes et iniuriam bibit,qui mittit verba per manum stulti.
PROV|26|7|Quomodo molles claudo tibiae,sic in ore stultorum parabola.
PROV|26|8|Sicut qui celat lapidem in acervo,ita qui tribuit insipienti honorem.
PROV|26|9|Spina crescens in manu temulenti,sic parabola in ore stultorum.
PROV|26|10|Sagittarius, qui conicit ad omnia,ita qui stultum conducit et qui vagos conducit.
PROV|26|11|Sicut canis, qui revertitur ad vomitum suum,sic stultus, qui iterat stultitiam suam.
PROV|26|12|Vidisti hominem sapientem sibi videri?Magis illo spem habebit stultus.
PROV|26|13|Dicit piger: " Leaena est in via,et leo in plateis ".
PROV|26|14|Ostium vertitur in cardine suo,et piger in lectulo suo.
PROV|26|15|Abscondit piger manum in catinoet laborat, si ad os suum eam converterit.
PROV|26|16|Sapientior sibi piger videturseptem viris respondentibus sententias.
PROV|26|17|Apprehendit auribus canem,qui transiens commiscetur rixae alterius.
PROV|26|18|Sicut insanit, qui mittit sagittaset lanceas in mortem,
PROV|26|19|ita vir, qui decipit amicum suumet dicit: " Nonne ludens feci? ".
PROV|26|20|Cum defecerint ligna, exstinguetur ignis,et, susurrone subtracto, iurgia conquiescent.
PROV|26|21|Sicut carbones ad prunas et ligna ad ignem,sic homo litigiosus ad inflammandas rixas.
PROV|26|22|Verba susurronis quasi dulciaet ipsa perveniunt ad intima ventris.
PROV|26|23|Sicut argentum sordidum ornans vas fictile,sic labia levia et cor malum.
PROV|26|24|Labiis suis se dissimulabit inimicus,cum in corde tractaverit dolos:
PROV|26|25|quando mollierit vocem suam, ne credideris ei,quoniam septem abominationes sunt in corde illius;
PROV|26|26|operiet odium fraudulenter,revelabitur autem malitia eius in concilio.
PROV|26|27|Qui fodit foveam, incidet in eam;et, qui volvit lapidem, revertetur ad eum.
PROV|26|28|Lingua fallax non amat veritatem,et os lubricum operatur ruinas.
PROV|27|1|Ne glorieris in crastinumignorans, quid superventura pariat dies.
PROV|27|2|Laudet te alienus et non os tuum,extraneus et non labia tua.
PROV|27|3|Grave est saxum et onerosa arena,sed ira stulti utroque gravior.
PROV|27|4|Saevitas et erumpens furor,et coram zelo consistere quis poterit?
PROV|27|5|Melior est manifesta correptioquam amor absconditus.
PROV|27|6|Veriora sunt vulnera diligentisquam fraudulenta oscula odientis.
PROV|27|7|Anima saturata calcabit favum,et anima esuriens etiam amarum pro dulci sumet.
PROV|27|8|Sicut avis transmigrans de nido suo,sic vir errans longe a loco suo.
PROV|27|9|Unguento et ture delectatur coret dulcedine amici in consilio ex animo.
PROV|27|10|Amicum tuum et amicum patris tui ne dimiseriset domum fratris tui ne ingrediaris in die afflictionis tuae.Melior est vicinus iuxta quam frater procul.
PROV|27|11|Stude sapientiae, fili mi, et laetifica cor meum,ut possim exprobranti mihi respondere sermonem.
PROV|27|12|Astutus videns malum absconditus est;simplices transeuntes multati sunt.
PROV|27|13|Tolle vestimentum eius, qui spopondit pro extraneo,et pro alienis aufer ei pignus.
PROV|27|14|Qui benedicit proximo suo voce grandi mane consurgens,maledictio reputabitur ei.
PROV|27|15|Tecta perstillantia in die frigoriset litigiosa mulier comparantur;
PROV|27|16|qui retinet eam, quasi qui ventum teneat,et oleum dextera sua tenere reperietur.
PROV|27|17|Ferrum ferro exacuitur,et homo exacuit faciem amici sui.
PROV|27|18|Qui servat ficum, comedet fructus eius;et, qui custos est domini sui, glorificabitur.
PROV|27|19|Quomodo in aqua facies prospicit ad faciem,sic cor hominis ad hominem.
PROV|27|20|Infernus et Perditio numquam implentur,similiter et oculi hominum insatiabiles.
PROV|27|21|Quomodo probatur in conflatorio argentum et in fornace aurum,sic probatur homo ore laudantis.
PROV|27|22|Si pilo contuderis stultum in pila quasi ptisanas,non auferetur ab eo stultitia eius.
PROV|27|23|Diligenter agnosce vultum pecoris tui;appone cor tuum ad greges,
PROV|27|24|non enim habebis iugiter divitias.Num corona tribuetur in generationem et generationem?
PROV|27|25|Nudata sunt prata, et apparuerunt herbae virentes,et collecta sunt fena de montibus;
PROV|27|26|agni ad vestimentum tuum,et haedi ad agri pretium;
PROV|27|27|sufficiat tibi lac caprarum in cibum tuumet in cibum domus tuae et ad victum ancillis tuis.
PROV|28|1|Fugit impius, nemine persequente;iustus autem quasi leo confidens.
PROV|28|2|Propter peccata terrae multi principes eius;et propter hominem intellegentem et sapientemrectus ordo longior erit.
PROV|28|3|Vir pauper et calumnians pauperessimilis est imbri vehementi, in quo paratur fames.
PROV|28|4|Qui derelinquunt legem, laudant impium;qui custodiunt, succenduntur contra eum.
PROV|28|5|Viri mali non intellegunt iudicium;qui autem requirunt Dominum, animadvertunt omnia.
PROV|28|6|Melior est pauper ambulans in simplicitate suaquam perversus in viis suis, quamquam dives.
PROV|28|7|Qui custodit legem, filius sapiens est;qui autem comissatores pascit, confundit patrem suum.
PROV|28|8|Qui coacervat divitias suas usuris et fenore,liberali in pauperes congregat eas.
PROV|28|9|Qui declinat aures suas, ne audiat legem,oratio quoque eius erit exsecrabilis.
PROV|28|10|Qui decipit iustos in via mala, in interitu suo corruet,et simplices possidebunt bona eius.
PROV|28|11|Sapiens sibi videtur vir dives,pauper autem prudens scrutabitur eum.
PROV|28|12|In exsultatione iustorum multa gloria est,et, cum exaltantur impii, abscondit se homo.
PROV|28|13|Qui abscondit scelera sua, non prosperabit;qui autem confessus fuerit et reliquerit ea,misericordiam consequetur.
PROV|28|14|Beatus homo, qui semper est pavidus;qui vero indurat cor suum, corruet in malum.
PROV|28|15|Leo rugiens et ursus esuriensprinceps impius super populum pauperem.
PROV|28|16|Dux indigens prudentia multos opprimet;qui autem odit avaritiam, longi fient dies eius.
PROV|28|17|Hominem, animae cuiusdam sanguine gravatum,si usque ad lacum fugerit, nemo sustineat.
PROV|28|18|Qui ambulat simpliciter, salvus erit;qui perversis graditur viis, subito concidet.
PROV|28|19|Qui operatur terram suam, satiabitur panibus;qui autem sectatur otium, replebitur egestate.
PROV|28|20|Vir fidelis multum laudabitur;qui autem festinat ditari, non erit innocens.
PROV|28|21|Qui dignoscit in iudicio faciem, non benefacit;et pro buccella panis praevaricatur homo.
PROV|28|22|Festinat ditari vir invidus,ignorat quod egestas superveniet ei.
PROV|28|23|Qui corripit hominem, gratiam postea invenietmagis quam ille, qui lingua blanditur.
PROV|28|24|Qui abripit aliquid a patre suo et a matreet dicit: " Hoc non est peccatum ",particeps homicidae est.
PROV|28|25|Qui desiderium dilatat, iurgia concitat;qui vero sperat in Domino, impinguabitur.
PROV|28|26|Qui confidit in corde suo, stultus est;qui autem graditur sapienter, ipse salvabitur.
PROV|28|27|Qui dat pauperi, non indigebit;qui autem occultat oculos, abundabit maledictis.
PROV|28|28|Cum surrexerint impii, abscondentur homines;cum illi perierint, multiplicabuntur iusti.
PROV|29|1|Vir, qui correptiones dura cervice contemnit,subito conteretur absque sanatione.
PROV|29|2|In multiplicatione iustorum laetabitur vulgus;et in dominatione impii gemet populus.
PROV|29|3|Vir, qui amat sapientiam, laetificat patrem suum;qui autem nutrit scorta, perdet substantiam.
PROV|29|4|Rex in iustitia erigit terram;vir acceptor donorum destruet eam.
PROV|29|5|Homo, qui blanditur amico suo,rete expandit gressibus eius.
PROV|29|6|In peccato vir iniquus irretitur laqueo,et iustus exsultabit atque gaudebit.
PROV|29|7|Novit iustus causam pauperum,impius ignorat scientiam.
PROV|29|8|Homines pestilentes dissipant civitatem;sapientes vero avertunt furorem.
PROV|29|9|Vir sapiens, si cum stulto iudicio contenderit,sive irascatur sive rideat, non inveniet requiem.
PROV|29|10|Viri sanguinum oderunt simplicem;iusti autem quaerunt animam eius.
PROV|29|11|Totum spiritum suum profert stultus;sapiens mitigat eum in posterum.
PROV|29|12|Princeps, qui libenter audit verba mendacii,omnes ministros habet impios.
PROV|29|13|Pauper et oppressor obviaverunt sibi,utriusque oculorum illuminator est Dominus.
PROV|29|14|Rex, qui iudicat in veritate pauperes,thronus eius in aeternum firmabitur.
PROV|29|15|Virga atque correptio tribuit sapientiam;puer autem, qui dimittitur voluntati suae, confundit matrem suam.
PROV|29|16|In multiplicatione impiorum multiplicabuntur scelera,et iusti ruinas eorum videbunt.
PROV|29|17|Erudi filium tuum, et refrigerabit teet dabit delicias animae tuae.
PROV|29|18|Cum visio defecerit, dissipabitur populus;qui vero custodit legem, beatus est.
PROV|29|19|Servus verbis non potest erudiri,quia intellegit et respondere contemnit.
PROV|29|20|Vidisti hominem velocem ad loquendum?Magis illo spem habebit insipiens.
PROV|29|21|Qui delicate a pueritia nutrit servum suum,postea sentiet eum contumacem.
PROV|29|22|Vir iracundus provocat rixas;et, qui ad indignandum facilis est, erit ad peccandum proclivior.
PROV|29|23|Superbia hominis humiliabit eum,et humilis spiritu suscipiet gloriam.
PROV|29|24|Qui cum fure participat, odit animam suam;adiuramentum audit et non indicat.
PROV|29|25|Timor hominis inducit laqueum;qui sperat in Domino, sublevabitur.
PROV|29|26|Multi requirunt faciem principis;et iudicium a Domino egreditur singulorum.
PROV|29|27|Abominantur iusti virum impium;et abominantur impii eos, qui recta sunt via.
PROV|30|1|Verba Agur filii Iaces ex Massa.Oraculum hominis ad Itiel,ad Itiel et Ucal.
PROV|30|2|Quoniam stultissimus sum virorum,et sapientia hominum non est mecum;
PROV|30|3|et non didici sapientiamet scientiam sanctorum non novi.
PROV|30|4|Quis ascendit in caelum atque descendit?Quis continuit spiritum in manibus suis?Quis colligavit aquas quasi in vestimento?Quis statuit omnes terminos terrae?Quod nomen est eius, et quod nomen filii eius, si nosti?
PROV|30|5|Omnis sermo Dei probatusclipeus est sperantibus in eum.
PROV|30|6|Ne addas quidquam verbis illius:et arguaris inveniarisque mendax.
PROV|30|7|Duo rogavi te,ne deneges mihi, antequam moriar:
PROV|30|8|vanitatem et verba mendacia longe fac a me,mendicitatem et divitias ne dederis mihi,tribue tantum victum demensum mihi,
PROV|30|9|ne forte satiatus illiciar ad negandumet dicam: " Quis est Dominus? "aut egestate compulsus fureret periurem nomen Dei mei.
PROV|30|10|Ne calumnieris servum ad dominum suum,ne forte maledicat tibi, et puniaris.
PROV|30|11|Generatio, quae patri suo maledicitet quae matri suae non benedicit.
PROV|30|12|Generatio, quae sibi munda videturet non est lota a sordibus suis.
PROV|30|13|Generatio, cuius oculi quam excelsi sunt,et palpebrae eius in alta surrectae!
PROV|30|14|Generatio, quae pro dentibus gladios habet,et cultri molares eius,ut comedat inopes de terraet pauperes ex hominibus.
PROV|30|15|Sanguisugae duae sunt filiae: Affer, affer! ".Tria sunt insaturabilia,et quattuor, quae numquam dicunt: " Sufficit! ":
PROV|30|16|infernus et venter sterilis,terra, quae non satiatur aqua,ignis, qui numquam dicit: " Sufficit! ".
PROV|30|17|Oculum, qui subsannat patremet qui despicit obsequium matris suae,effodiant eum corvi de torrente,et comedant eum filii aquilae.
PROV|30|18|Tria sunt nimis difficilia mihi,et quattuor penitus ignoro:
PROV|30|19|viam aquilae in caelo,viam colubri super petram,viam navis in medio mariet viam viri in adulescentula.
PROV|30|20|Talis est et via mulieris adulterae,quae comedit et tergens os suum dicit: Non sum operata malum ".
PROV|30|21|Per tria movetur terra,et quattuor non potest sustinere:
PROV|30|22|per servum, cum regnaverit,per stultum, cum saturatus fuerit cibo,
PROV|30|23|per odiosam mulierem, cum in matrimonio fuerit assumpta,et per ancillam, cum fuerit heres dominae suae.
PROV|30|24|Quattuor sunt minima terrae,et ipsa sunt sapientiora sapientibus:
PROV|30|25|formicae populus infirmus,quae praeparant in messe cibum sibi;
PROV|30|26|hyraces plebs invalida,qui collocant in petra cubile suum;
PROV|30|27|regem locusta non habetet egreditur universa per turmas suas;
PROV|30|28|stellio manibus nitituret moratur in aedibus regis.
PROV|30|29|Tria sunt, quae bene gradiuntur,et quattuor, quae incedunt feliciter:
PROV|30|30|leo fortissimus bestiarumad nullius pavebit occursum,
PROV|30|31|gallus succinctus lumbos et arieset rex, qui secum habet exercitum.
PROV|30|32|Si stultum te praebuisti, postquam elevatus es in sublime,et si considerasti, ori impone manum.
PROV|30|33|Qui enim fortiter premit lac, exprimit butyrum,et, qui vehementer emungit nares, elicit sanguinem,et, qui provocat iras, producit discordias.
PROV|31|1|Verba Lamuelis regis Massa, quae erudivit eum mater eius.
PROV|31|2|Quid, fili mi? Quid, fili uteri mei?Quid, fili votorum meorum?
PROV|31|3|Ne dederis mulieribus substantiam tuamet vias tuas illis, quae delent reges.
PROV|31|4|Non decet reges, o Lamuel, non decet reges bibere vinum,nec magistratus desiderare siceram,
PROV|31|5|ne forte bibant et obliviscantur iudiciorumet mutent causam omnium filiorum pauperis.
PROV|31|6|Date siceram pereuntiet vinum his, qui amaro sunt animo:
PROV|31|7|bibat et obliviscatur egestatis suaeet doloris sui non recordetur amplius.
PROV|31|8|Aperi os tuum pro mutoet causis omnium filiorum, qui pereunt;
PROV|31|9|aperi os tuum, decerne, quod iustum est,et iudica inopem et pauperem.
PROV|31|10|ALEPH. Mulierem fortem quis inveniet?Longe super gemmas pretium eius.
PROV|31|11|BETH. Confidit in ea cor viri sui et spoliis non indigebit.
PROV|31|12|GHIMEL. Reddet ei bonum et non malum omnibus diebus vitae suae.
PROV|31|13|DALETH. Quaesivit lanam et linumet operata est delectatione manuum suarum.
PROV|31|14|HE. Facta est quasi navis institorisde longe portans panem suum.
PROV|31|15|VAU. Et de nocte surrexitdeditque praedam domesticis suiset cibaria ancillis suis.
PROV|31|16|ZAIN. Consideravit agrum et emit eum;de fructu manuum suarum plantavit vineam.
PROV|31|17|HETH. Accinxit fortitudine lumbos suoset roboravit brachium suum.
PROV|31|18|TETH. Gustavit et vidit quia bona est negotiatio eius;non exstinguetur in nocte lucerna eius.
PROV|31|19|IOD. Manum suam misit ad colos,et digiti eius apprehenderunt fusum.
PROV|31|20|CAPH. Palmas suas aperuit inopiet manum suam extendit ad pauperem.
PROV|31|21|LAMED. Non timebit domui suae a frigoribus nivis:omnes enim domestici eius vestiti sunt duplicibus.
PROV|31|22|MEM. Stragulatam vestem fecit sibi;byssus et purpura indumentum eius.
PROV|31|23|NUN. Nobilis in portis vir eius,quando sederit cum senatoribus terrae.
PROV|31|24|SAMECH. Sindonem fecit et vendiditet cingulum tradidit Chananaeo.
PROV|31|25|Ain. Fortitudo et decor indumentum eius,et ridebit in die novissimo.
PROV|31|26|PHE. Os suum aperuit sapientiae,et lex clementiae in lingua eius.
PROV|31|27|SADE. Consideravit semitas domus suaeet panem otiosa non comedit.
PROV|31|28|COPH. Surrexerunt filii eius et beatissimam praedicaverunt,vir eius et laudavit eam:
PROV|31|29|RES. " Multae filiae fortiter operatae sunt,tu supergressa es universas ".
PROV|31|30|SIN. Fallax gratia et vana est pulchritudo;mulier timens Dominum ipsa laudabitur.
PROV|31|31|TAU. Date ei de fructu manuum suarum,et laudent eam in portis opera eius.
