COL|1|1|Paulus, apostolus Christi Iesu per voluntatem Dei, et Timo theus frater
COL|1|2|his, qui sunt Colossis, sanctis et fidelibus fratribus in Christo: gratia vobis et pax a Deo Patre nostro.
COL|1|3|Gratias agimus Deo Patri Domini nostri Iesu Christi semper pro vobis orantes,
COL|1|4|audientes fidem vestram in Christo Iesu et dilectionem, quam habetis in sanctos omnes,
COL|1|5|propter spem, quae reposita est vobis in caelis, quam ante audistis in verbo veritatis evangelii,
COL|1|6|quod pervenit ad vos, sicut et in universo mundo est fructificans et crescens, sicut et in vobis, ex ea die, qua audistis et cognovistis gratiam Dei in veritate;
COL|1|7|sicut didicistis ab Epaphra carissimo conservo nostro, qui est fidelis pro nobis minister Christi,
COL|1|8|qui etiam manifestavit nobis dilectionem vestram in Spiritu.
COL|1|9|Ideo et nos, ex qua die audivimus, non cessamus pro vobis orantes et postulantes, ut impleamini agnitione voluntatis eius in omni sapientia et intellectu spiritali,
COL|1|10|ut ambuletis digne Domino per omnia placentes, in omni opere bono fructificantes et crescentes in scientia Dei,
COL|1|11|in omni virtute confortati secundum potentiam claritatis eius in omnem patientiam et longanimitatem, cum gaudio
COL|1|12|gratias agentes Patri,qui idoneos vos fecit in partem sortis sanctorum in lumine;
COL|1|13|qui eripuit nos de potestate tenebrarumet transtulit in regnum Filii dilectionis suae,
COL|1|14|in quo habemus redemptionem,remissionem peccatorum;
COL|1|15|qui est imago Dei invisibilis,primogenitus omnis creaturae,
COL|1|16|quia in ipso condita sunt universa in caelis et in terra,visibilia et invisibilia,sive throni sive dominationessive principatus sive potestates.Omnia per ipsum et in ipsum creata sunt,
COL|1|17|et ipse est ante omnia,et omnia in ipso constant.
COL|1|18|Et ipse est caput corporis ecclesiae;qui est principium, primogenitus ex mortuis,ut sit in omnibus ipse primatum tenens,
COL|1|19|quia in ipso complacuit omnem plenitudinem habitare
COL|1|20|et per eum reconciliare omnia in ipsum,pacificans per sanguinem crucis eius,sive quae in terris sive quae in caelis sunt.
COL|1|21|Et vos, cum essetis aliquando alienati et inimici sensu in operibus malis,
COL|1|22|nunc autem reconciliavit in corpore carnis eius per mortem exhibere vos sanctos et immaculatos et irreprehensibiles coram ipso;
COL|1|23|si tamen permanetis in fide fundati et stabiles et immobiles a spe evangelii, quod audistis, quod praedicatum est in universa creatura, quae sub caelo est, cuius factus sum ego Paulus minister.
COL|1|24|Nunc gaudeo in passionibus pro vobis et adimpleo, ea quae desunt passionum Christi in carne mea pro corpore eius, quod est ecclesia,
COL|1|25|cuius factus sum ego minister secundum dispensationem Dei, quae data est mihi in vos, ut impleam verbum Dei;
COL|1|26|mysterium, quod absconditum fuit a saeculis et generationibus, nunc autem manifestatum est sanctis eius,
COL|1|27|quibus voluit Deus notas facere divitias gloriae mysterii huius in gentibus, quod est Christus in vobis, spes gloriae;
COL|1|28|quem nos annuntiamus, commonentes omnem hominem et docentes omnem hominem in omni sapientia, ut exhibeamus omnem hominem perfectum in Christo;
COL|1|29|ad quod et laboro certando secundum operationem eius, quae operatur in me in virtute.
COL|2|1|Volo enim vos scire qualem sollicitudinem habeam pro vo bis et pro his, qui sunt Laodiciae, et quicumque non viderunt faciem meam in carne,
COL|2|2|ut consolentur corda ipsorum instructi in caritate et in omnes divitias plenitudinis intellectus, in agnitionem mysterii Dei, Christi,
COL|2|3|in quo sunt omnes thesauri sapientiae et scientiae absconditi.
COL|2|4|Hoc dico, ut nemo vos decipiat in subtilitate sermonum.
COL|2|5|Nam etsi corpore absens sum, sed spiritu vobiscum sum, gaudens et videns ordinem vestrum et firmamentum eius, quae in Christum est, fidei vestrae.
COL|2|6|Sicut ergo accepistis Christum Iesum Dominum, in ipso ambulate,
COL|2|7|radicati et superaedificati in ipso et confirmati fide, sicut didicistis, abundantes in gratiarum actione.
COL|2|8|Videte, ne quis vos depraedetur per philosophiam et inanem fallaciam secundum traditionem hominum, secundum elementa mundi et non secundum Christum;
COL|2|9|quia in ipso inhabitat omnis plenitudo divinitatis corporaliter,
COL|2|10|et estis in illo repleti, qui est caput omnis principatus et potestatis;
COL|2|11|in quo et circumcisi estis circumcisione non manufacta in exspoliatione corporis carnis, in circumcisione Christi;
COL|2|12|consepulti ei in baptismo, in quo et conresuscitati estis per fidem operationis Dei, qui suscitavit illum a mortuis;
COL|2|13|et vos, cum mortui essetis in delictis et praeputio carnis vestrae, convivificavit cum illo, donans nobis omnia delicta,
COL|2|14|delens, quod adversum nos erat, chirographum decretis, quod erat contrarium nobis, et ipsum tulit de medio affigens illud cruci;
COL|2|15|exspolians principatus et potestates traduxit confidenter, triumphans illos in semetipso.
COL|2|16|Nemo ergo vos iudicet in cibo aut in potu aut ex parte diei festi aut neomeniae aut sabbatorum,
COL|2|17|quae sunt umbra futurorum, corpus autem Christi.
COL|2|18|Nemo vos bravio defraudet complacens sibi in humilitate et religione angelorum propter ea, quae vidit, ingrediens, frustra inflatus sensu carnis suae
COL|2|19|et non tenens caput, ex quo totum corpus per nexus et coniunctiones subministratum et compaginatum crescit in augmentum Dei.
COL|2|20|Si mortui estis cum Christo ab elementis mundi, quid tamquam viventes in mundo decretis subicimini:
COL|2|21|" Ne tetigeris neque gustaveris neque contrectaveris ",
COL|2|22|quae sunt omnia in corruptionem ipso usu secundum praecepta et doctrinas hominum?
COL|2|23|Quae sunt rationem quidem habentia sapientiae in superstitione et humilitate, et non parcendo corpori, non in honore aliquo ad saturitatem carnis.
COL|3|1|Igitur, si conresurrexistis Chri sto, quae sursum sunt quaerite, ubi Christus est in dextera Dei sedens;
COL|3|2|quae sursum sunt sapite, non quae supra terram.
COL|3|3|Mortui enim estis, et vita vestra abscondita est cum Christo in Deo!
COL|3|4|Cum Christus apparuerit, vita vestra, tunc et vos apparebitis cum ipso in gloria.
COL|3|5|Mortificate ergo membra, quae sunt super terram: fornicationem, immunditiam, libidinem, concupiscentiam malam et avaritiam, quae est simulacrorum servitus,
COL|3|6|propter quae venit ira Dei super filios incredulitatis;
COL|3|7|in quibus et vos ambulastis aliquando, cum viveretis in illis.
COL|3|8|Nunc autem deponite et vos omnia: iram, indignationem, malitiam, blasphemiam, turpem sermonem de ore vestro;
COL|3|9|nolite mentiri invicem, qui exuistis vos veterem hominem cum actibus eius
COL|3|10|et induistis novum, eum, qui renovatur in agnitionem secundum imaginem eius, qui creavit eum,
COL|3|11|ubi non est Graecus et Iudaeus, circumcisio et praeputium, barbarus, Scytha, servus, liber, sed omnia et in omnibus Christus.
COL|3|12|Induite vos ergo, sicut electi Dei, sancti et dilecti, viscera misericordiae, benignitatem, humilitatem, mansuetudinem, longanimitatem,
COL|3|13|supportantes invicem et donantes vobis ipsis, si quis adversus aliquem habet querelam; sicut et Dominus donavit vobis, ita et vos;
COL|3|14|super omnia autem haec: caritatem, quod est vinculum perfectionis.
COL|3|15|Et pax Christi dominetur in cordibus vestris, ad quam et vocati estis in uno corpore. Et grati estote.
COL|3|16|Verbum Christi habitet in vobis abundanter, in omni sapientia docentes et commonentes vosmetipsos psalmis, hymnis, canticis spiritalibus, in gratia cantantes in cordibus vestris Deo;
COL|3|17|et omne, quodcumque facitis in verbo aut in opere, omnia in nomine Domini Iesu gratias agentes Deo Patri per ipsum.
COL|3|18|Mulieres, subditae estote viris, sicut oportet in Domino.
COL|3|19|Viri, diligite uxores et nolite amari esse ad illas.
COL|3|20|Filii, oboedite parentibus per omnia; hoc enim placitum est in Domino.
COL|3|21|Patres, nolite ad indignationem provocare filios vestros, ut non pusillo animo fiant.
COL|3|22|Servi, oboedite per omnia dominis carnalibus, non ad oculum servientes, quasi hominibus placentes, sed in simplicitate cordis, timentes Dominum.
COL|3|23|Quodcumque facitis, ex animo operamini sicut Domino et non hominibus,
COL|3|24|scientes quod a Domino accipietis retributionem hereditatis. Domino Christo servite;
COL|3|25|qui enim iniuriam facit, recipiet id quod inique gessit, et non est personarum acceptio.
COL|4|1|Domini, quod iustum est et aequum, servis praestate, scien tes quoniam et vos Dominum habetis in caelo.
COL|4|2|Orationi instate, vigilantes in ea in gratiarum actione,
COL|4|3|orantes simul et pro nobis, ut Deus aperiat nobis ostium sermonis ad loquendum mysterium Christi, propter quod etiam vinctus sum,
COL|4|4|ut manifestem illud, ita ut oportet me loqui.
COL|4|5|In sapientia ambulate ad eos, qui foris sunt, tempus redimentes.
COL|4|6|Sermo vester semper sit in gratia, sale conditus, ut sciatis quomodo oporteat vos unicuique respondere.
COL|4|7|Quae circa me sunt, omnia vobis nota faciet Tychicus, carissimus frater et fidelis minister et conservus in Domino,
COL|4|8|quem misi ad vos ad hoc ipsum, ut cognoscatis, quae circa nos sunt, et consoletur corda vestra,
COL|4|9|cum Onesimo fideli et carissimo fratre, qui est ex vobis; omnia, quae hic aguntur, nota facient vobis.
COL|4|10|Salutat vos Aristarchus concaptivus meus et Marcus consobrinus Barnabae, de quo accepistis mandata - si venerit ad vos, excipite illum -
COL|4|11|et Iesus, qui dicitur Iustus, qui sunt ex circumcisione; hi soli adiutores in regno Dei, qui mihi fuerunt solacio.
COL|4|12|Salutat vos Epaphras, qui ex vobis est, servus Christi Iesu, semper certans pro vobis in orationibus, ut stetis perfecti et impleti in omni voluntate Dei.
COL|4|13|Testimonium enim illi perhibeo, quod habet multum laborem pro vobis et pro his, qui sunt Laodiciae et qui Hierapoli.
COL|4|14|Salutat vos Lucas, medicus carissimus, et Demas.
COL|4|15|Salutate fratres, qui sunt Laodiciae, et Nympham et, quae in domo eius est, ecclesiam.
COL|4|16|Et cum lecta fuerit apud vos epistula, facite ut et in Laodicensium ecclesia legatur, et eam, quae ex Laodicia est, vos quoque legatis.
COL|4|17|Et dicite Archippo: " Vide ministerium, quod accepisti in Domino, ut illud impleas ".
COL|4|18|Salutatio mea manu Pauli. Memores estote vinculorum meorum.Gratia vobiscum.
