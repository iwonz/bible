DAN|1|1|犹大 王 约雅敬 在位第三年， 巴比伦 王 尼布甲尼撒 来到 耶路撒冷 ，将城围困。
DAN|1|2|主将 犹大 王 约雅敬 和上帝殿中的一些器皿交在他的手中。他就把他们带到 示拿 地他神明的庙里，将器皿收入他神明的库房中。
DAN|1|3|王吩咐太监长 亚施毗拿 ，从 以色列 人的王室后裔和贵族中带进几个人来，
DAN|1|4|就是没有残疾、相貌俊美、通达各样学问 、知识聪明俱备、足能在王宫侍立的少年，要教他们 迦勒底 的文字和语言。
DAN|1|5|王从自己所用的膳和所饮的酒中，派给他们每日的分量，养育他们三年，好叫他们期满以后侍立在王面前。
DAN|1|6|他们中间有 犹大 人 但以理 、 哈拿尼雅 、 米沙利 和 亚撒利雅 。
DAN|1|7|太监长给他们另外起名，称 但以理 为 伯提沙撒 ，称 哈拿尼雅 为 沙得拉 ，称 米沙利 为 米煞 ，称 亚撒利雅 为 亚伯尼歌 。
DAN|1|8|但以理 却立志，不以王的膳和王所饮的酒玷污自己，于是恳求太监长容他不使自己玷污。
DAN|1|9|上帝使 但以理 在太监长眼前蒙恩，得怜悯。
DAN|1|10|太监长对 但以理 说：“我惧怕我主我王，他已经派给你们饮食，何必让他见你们的面貌比你们同年龄的少年憔悴呢？这样，你们就使我的头在王那里不保了。”
DAN|1|11|但以理 对太监长所派监管 但以理 、 哈拿尼雅 、 米沙利 、 亚撒利雅 的管理者说：
DAN|1|12|“请你考验仆人们十天，给我们素菜吃，清水喝，
DAN|1|13|然后你亲自观察我们的面貌和那用王膳的少年的面貌；就照你所观察的待你的仆人吧！”
DAN|1|14|管理者准许他们这件事，考验他们十天。
DAN|1|15|过了十天，他们的身材看来比所有享用王膳的少年更加俊美健壮，
DAN|1|16|于是管理者撤去王派给他们用的膳和所饮的酒，只给他们素菜。
DAN|1|17|这四个少年，上帝在各样文字学问上赐给他们知识和聪明； 但以理 又明白各样异象和梦兆。
DAN|1|18|王吩咐带他们进宫的日子到了，太监长就把他们带到 尼布甲尼撒 面前。
DAN|1|19|王与他们谈论，在所有少年中找不到人能与 但以理 、 哈拿尼雅 、 米沙利 、 亚撒利雅 相比，于是他们就在王面前侍立。
DAN|1|20|王考问他们一切智慧和聪明的事，发现他们比全国所有的术士和巫师胜过十倍。
DAN|1|21|到 居鲁士 王元年， 但以理 还健在。
DAN|2|1|尼布甲尼撒 在位第二年，他做了很多梦，心里烦乱，不能睡觉。
DAN|2|2|王吩咐人将术士、巫师、行邪术的和 迦勒底 人召来，要他们把王的梦告诉王；他们就来，站在王面前。
DAN|2|3|王对他们说：“我做了一个梦，心里烦乱，想要知道这是什么梦。”
DAN|2|4|迦勒底 人用 亚兰 话对王说：“愿王万岁！请将梦告诉仆人，我们就可以讲解。”
DAN|2|5|王回答 迦勒底 人说：“这事我已决定，你们若不把梦和梦的解释告诉我，就必被凌迟，你们的房屋必成粪堆；
DAN|2|6|但你们若能说出这个梦和梦的解释，就必从我得到礼物、赏赐和殊荣。现在，你们要把梦和梦的解释告诉我。”
DAN|2|7|他们再一次回答说：“请王将梦告诉仆人，我们就可以讲解。”
DAN|2|8|王回答说：“我确实知道你们是故意拖延，因为你们知道这事我已决定。
DAN|2|9|你们若不将梦告诉我，只有一个办法对待你们；因为你们彼此串通，向我胡言乱语，要等候情势改变。现在，你们要将梦告诉我，让我知道你们真能为我解梦。”
DAN|2|10|迦勒底 人回答王说：“世上没有人能解释王的事情；从来没有君王、大臣、掌权者向术士、巫师，或 迦勒底 人问过这样的事。
DAN|2|11|王所问的事很难，除了不与血肉之躯同住的上帝，没有人能在王面前解释。”
DAN|2|12|王因这事生气，大大震怒，吩咐灭绝 巴比伦 所有的智慧人。
DAN|2|13|命令发出，智慧人将要被杀，人就寻找 但以理 和他的同伴，要杀他们。
DAN|2|14|王的护卫长 亚略 奉命去杀 巴比伦 的智慧人， 但以理 用婉言和智慧回应，
DAN|2|15|向王的大臣 亚略 说：“王的命令为何这样紧急呢？” 亚略 就把事情告诉 但以理 。
DAN|2|16|于是 但以理 进去求王宽限，好为王解梦。
DAN|2|17|但以理 回到他的居所，把这事告诉他的同伴 哈拿尼雅 、 米沙利 、 亚撒利雅 ，
DAN|2|18|要他们祈求天上的上帝施怜悯，将这奥秘指明，免得 但以理 和他的同伴与 巴比伦 其余的智慧人一同灭亡。
DAN|2|19|这奥秘就在夜间异象中显明给 但以理 ， 但以理 就称颂天上的上帝。
DAN|2|20|但以理 说： “上帝的名是应当称颂的，从亘古直到永远！ 因为智慧和能力都属乎他。
DAN|2|21|他改变时间、季节， 他废王，立王； 将智慧赐给智慧人， 将知识赐给聪明人。
DAN|2|22|他显明深奥隐秘的事， 洞悉幽暗中的一切， 光明也与他同住。
DAN|2|23|我列祖的上帝啊，我感谢你，赞美你， 因你将智慧才能赐给我， 我们所求问的现在你已指明给我， 把王的事给我们指明。”
DAN|2|24|于是， 但以理 进到王所派灭绝 巴比伦 智慧人的 亚略 那里去，对他这样说：“不要灭绝 巴比伦 的智慧人，求你领我到王面前，我可以为王解梦。”
DAN|2|25|亚略 就急忙领 但以理 到王面前，对王这样说：“我在被掳的 犹大 人中找到一人，能将梦的解释告诉王。”
DAN|2|26|王对那称为 伯提沙撒 的 但以理 说：“你能将我所做的梦和梦的解释告诉我吗？”
DAN|2|27|但以理 回答王说：“王所问的那奥秘，智慧人、巫师、术士、观兆的都不能告诉王，
DAN|2|28|只有那在天上的上帝能显明奥秘。他已把日后将要发生的事指示 尼布甲尼撒 王。你在床上做的梦和你脑中的异象是这样：
DAN|2|29|你，王啊，你在床上所思想的是关乎日后的事，那显明奥秘的主已把将来要发生的事指示你。
DAN|2|30|至于我，那奥秘显明给我，并非因我智慧胜过一切活着的人，而是为了让王知道梦的解释，知道你心里的意念。
DAN|2|31|“你，王啊，你正观看，看哪，有一个很大的像，这像甚高，极其光耀，立在你面前，形状非常可怕。
DAN|2|32|这像的头是纯金的，胸膛和膀臂是银的，腹部和腰是铜的，
DAN|2|33|腿是铁的，脚是半铁半泥的。
DAN|2|34|你正观看，见有一块非人手凿出来的石头打在它半铁半泥的脚上，把脚砸碎；
DAN|2|35|于是铁、泥、铜、银、金都一同砸得粉碎，如夏天禾场上的糠秕，被风吹散，无处可寻。打碎这像的石头成了一座大山，覆盖全地。
DAN|2|36|“这就是那梦；我们要在王面前讲解那梦。
DAN|2|37|你，王啊，你是诸王之王。天上的上帝已将国度、权势、能力、尊荣都赐给你。
DAN|2|38|世人和走兽，并天空的飞鸟，不论居住何处，他都交在你的手中，令你掌管这一切。你就是那金的头。
DAN|2|39|在你以后必兴起另一国，不及于你；又有第三国如铜，必掌管全地。
DAN|2|40|第四国必坚壮如铁，就像铁能打碎砸碎一切；铁怎样压碎一切，那国也必照样打碎压碎。
DAN|2|41|你既看见像的脚和脚趾头，一半是陶匠的泥，一半是铁，那国将来也必分裂。你既看见铁和泥搀杂，那国也必有铁的力量。
DAN|2|42|那脚趾头既是半铁半泥，那国也必半强半弱。
DAN|2|43|你既看见铁和泥搀杂，他们必有混杂的后裔，却不能彼此相合，正如铁和泥不能相合。
DAN|2|44|当诸王在位的时候，天上的上帝必另立一个永不败坏的国度，这国度必不归给其他百姓，却要打碎灭绝所有的国度，存立到永远。
DAN|2|45|你既看见非人手凿出来的一块石头从山而出，打碎铁、铜、泥、银、金，那就是至大的上帝把将来要发生的事给王指明。这梦是确实的，这解释也是准确的。”
DAN|2|46|当时， 尼布甲尼撒 王脸伏于地，向 但以理 下拜，并且吩咐人给他奉上供物和香。
DAN|2|47|王对 但以理 说：“你既能讲明这奥秘，你们的上帝诚然是万神之神、万王之主，是奥秘的启示者。”
DAN|2|48|于是王使 但以理 高升，赏赐他极多的礼物，派他管理 巴比伦 全省，又立他为总理，掌管 巴比伦 所有的智慧人。
DAN|2|49|但以理 求王，王就派 沙得拉 、 米煞 、 亚伯尼歌 管理 巴比伦 省的事务，只是 但以理 仍在朝中侍立。
DAN|3|1|尼布甲尼撒 王造了一个金像，高六十肘，宽六肘，立在 巴比伦 省的 杜拉 平原。
DAN|3|2|尼布甲尼撒 王差人将总督、钦差、省长、参谋、财务、法官、地方官和各省的官员都召了来，为 尼布甲尼撒 王所立的像行开光礼。
DAN|3|3|于是总督、钦差、省长、参谋、财务、法官、地方官和各省的官员都聚集，站在 尼布甲尼撒 所立的像前，要为 尼布甲尼撒 王所立的像行开光礼。
DAN|3|4|那时传令的大声呼叫说：“各方、各国、各族 的人哪，有命令传给你们：
DAN|3|5|你们一听见角、号、琴、瑟、三角琴、鼓和各样乐器的声音，就当俯伏，拜 尼布甲尼撒 王所立的金像。
DAN|3|6|凡不俯伏下拜的，必立刻扔在烈火的窑中。”
DAN|3|7|因此百姓一听见角、号、琴、瑟、三角琴 和各样乐器的声音，各方、各国、各族的人就都俯伏，拜 尼布甲尼撒 王所立的金像。
DAN|3|8|在那时，有几个 迦勒底 人进前来控告 犹大 人。
DAN|3|9|他们对 尼布甲尼撒 王说：“愿王万岁！
DAN|3|10|你，王啊，你曾降旨，凡听见角、号、琴、瑟、三角琴、鼓和各样乐器声音的，都当俯伏拜这金像。
DAN|3|11|凡不俯伏下拜的，必扔在烈火的窑中。
DAN|3|12|现在有几个 犹大 人，就是王所派管理 巴比伦 省事务的 沙得拉 、 米煞 、 亚伯尼歌 ；王啊，这些人不理你的谕旨，不事奉你的神明，也不拜你所立的金像。”
DAN|3|13|当时， 尼布甲尼撒 大发烈怒，命令把 沙得拉 、 米煞 、 亚伯尼歌 带过来；他们就把这几个人带到王面前。
DAN|3|14|尼布甲尼撒 对他们说：“ 沙得拉 、 米煞 、 亚伯尼歌 ，你们不事奉我的神明，不拜我所立的金像，是真的吗？
DAN|3|15|现在，你们若准备好，一听见角、号、琴、瑟、三角琴、鼓和各样乐器的声音，就俯伏拜我所造的像；若不下拜，必立刻扔在烈火的窑中，有哪一个神明能救你们脱离我的手呢？”
DAN|3|16|沙得拉 、 米煞 、 亚伯尼歌 对王说：“ 尼布甲尼撒 啊，这件事我们不必回答你，
DAN|3|17|即便如此，我们所事奉的上帝能将我们从烈火的窑中救出来。王啊，他必救我们脱离你的手；
DAN|3|18|即或不然，王啊，你当知道，我们绝不事奉你的神明，也不拜你所立的金像。”
DAN|3|19|当时， 尼布甲尼撒 怒气填胸，向 沙得拉 、 米煞 、 亚伯尼歌 变了脸色，命令把窑烧热，比平常热七倍；
DAN|3|20|又命令他军中的几个壮士，把 沙得拉 、 米煞 、 亚伯尼歌 捆起来，扔在烈火的窑中。
DAN|3|21|这三人穿着内袍、外衣、头巾和其他的衣服，被捆起来扔在烈火的窑中。
DAN|3|22|因为王的命令紧急，窑又非常热，那抬 沙得拉 、 米煞 、 亚伯尼歌 的人都被火焰烧死。
DAN|3|23|但是这三个人， 沙得拉 、 米煞 、 亚伯尼歌 被捆绑着，掉进烈火的窑中。
DAN|3|24|那时， 尼布甲尼撒 王惊奇，急忙站起来，对谋士说：“我们捆起来扔在火里的不是三个人吗？”他们回答王说：“王啊，是的。”
DAN|3|25|王说：“看哪，我看见有四个人，并没有捆绑，在火中行走，也没有受伤；那第四个的相貌好像神明的儿子。”
DAN|3|26|于是 尼布甲尼撒 靠近烈火窑门，说：“至高上帝的仆人 沙得拉 、 米煞 、 亚伯尼歌 ，出来，来吧！” 沙得拉 、 米煞 、 亚伯尼歌 就从火中出来。
DAN|3|27|那些总督、钦差、省长和王的谋士一同聚集来看这三个人，见火不能伤他们的身体，头发没有烧焦，衣裳也没有变色，都没有火烧过的气味。
DAN|3|28|尼布甲尼撒 说：“ 沙得拉 、 米煞 、 亚伯尼歌 的上帝是应当称颂的！他差遣使者救护倚靠他的仆人，他们不遵王的命令，甚至舍身，在他们上帝以外不肯事奉敬拜别神。
DAN|3|29|现在我降旨，无论何方、何国、何族，凡有人毁谤 沙得拉 、 米煞 、 亚伯尼歌 的上帝，他必被凌迟，他的房屋必成粪堆，因为没有别神能像这样施行拯救。”
DAN|3|30|那时王在 巴比伦 省使 沙得拉 、 米煞 、 亚伯尼歌 高升。
DAN|4|1|尼布甲尼撒 王对住在全地各方、各国、各族的人说：“愿你们大享平安！
DAN|4|2|我乐意宣扬至高上帝向我所行的神迹奇事。
DAN|4|3|他的神迹何其大！ 他的奇事何其盛！ 他的国度存到永远； 他的权柄存到万代！
DAN|4|4|“我－ 尼布甲尼撒 安居在家中，在宫里享受荣华。
DAN|4|5|我做了一个梦，使我惧怕。我在床上的意念和脑中的异象，使我惊惶。
DAN|4|6|因此我降旨召 巴比伦 的智慧人全都到我面前，要他们将梦的解释告诉我。
DAN|4|7|于是那些术士、巫师、 迦勒底 人、观兆的都进来，我将那梦告诉他们，他们却不能把梦的解释告诉我。
DAN|4|8|最后， 但以理 ，就是按照我神明的名字称为 伯提沙撒 的，来到我面前，他里头有神圣神明的灵，我将梦告诉他：
DAN|4|9|‘术士的领袖 伯提沙撒 啊，我知道你里头有神圣神明的灵，什么奥秘都不能为难你。现在你要把我梦中所见的异象和梦的解释告诉我 。’
DAN|4|10|“我在床上脑中的异象是这样：我观看，看哪，大地中间有一棵树，极其高大。
DAN|4|11|那树渐长，而且茁壮，高得顶天，从地极都能看见，
DAN|4|12|叶子华美，果子甚多，可作所有动物的食物；野地的走兽卧在荫下，天空的飞鸟宿在枝上，凡有血肉的都从这树得食物。
DAN|4|13|“我观看，我在床上脑中的异象是这样，看哪，有守望者，就是神圣的一位，从天而降，
DAN|4|14|大声呼叫说：‘砍倒这树！砍下枝子！拔掉叶子！抛散果子！使走兽逃离树下，飞鸟躲开树枝。
DAN|4|15|树的残干却要留在地里，在田野的青草中用铁圈和铜圈套住。任他让天上的露水滴湿，和地上的走兽一同吃草，
DAN|4|16|使他的心改变，不再是人的心，而给他一个兽心，使他经过七个时期 。
DAN|4|17|这是众守望者所发的命令，是众圣者所作的决定，好叫世人知道至高者在人的国中掌权，要将国赐给谁就赐给谁，并且立极卑微的人执掌国权。’
DAN|4|18|“这是我－ 尼布甲尼撒 王所做的梦。 伯提沙撒 啊，你要说明这梦的解释；我国中所有的智慧人都不能把梦的解释告诉我，惟独你能，因你里头有神圣神明的灵。”
DAN|4|19|于是称为 伯提沙撒 的 但以理 惊骇片时，心意惊惶。王说：“ 伯提沙撒 啊，不要因梦和梦的解释惊惶。” 伯提沙撒 回答说：“我主啊，愿这梦归给恨恶你的人，这梦的解释归给你的敌人。
DAN|4|20|你所见的树渐长，而且茁壮，高得顶天，全地都能看见，
DAN|4|21|叶子华美，果子甚多，可作所有动物的食物；野地的走兽住在其下，天空的飞鸟宿在枝上。
DAN|4|22|“王啊，这成长又茁壮的树就是你。你的威势成长及于天，你的权柄达到地极。
DAN|4|23|王既看见一位神圣的守望者从天而降，说：‘将这树砍倒毁坏，树的残干却要留在地里，在田野的青草中用铁圈和铜圈套住。任他让天上的露水滴湿，与野地的走兽一同吃草，直到经过七个时期。’
DAN|4|24|“王啊，梦的解释就是这样：临到我主我王的事是出于至高者的命令。
DAN|4|25|你必被赶出离开世人，与野地的走兽同住，吃草如牛，让天上的露水滴湿，且要经过七个时期，直等到你知道至高者在人的国中掌权，要将国赐给谁就赐给谁。
DAN|4|26|这使树的残干存留的命令，是要等你知道天在掌权，你的国必定归你。
DAN|4|27|王啊，求你悦纳我的谏言，以施行公义除去罪过，以怜悯穷人除掉罪恶，或者你的平安可以延长。”
DAN|4|28|这些事都临到 尼布甲尼撒 王。
DAN|4|29|过了十二个月，他在 巴比伦 王宫顶上散步。
DAN|4|30|王说：“这大 巴比伦 岂不是我用大能大力建为首都，要显示我威严的荣耀吗？”
DAN|4|31|这话还在王口中的时候，有声音从天降下，说：“ 尼布甲尼撒 王啊，有话对你说，你的国离开你了。
DAN|4|32|你必被赶出离开世人，与野地的走兽同住，吃草如牛，且要经过七个时期；等你知道至高者在人的国中掌权，要将国赐给谁就赐给谁。”
DAN|4|33|当时这话就应验在 尼布甲尼撒 身上，他被赶出离开世人，吃草如牛，身体被天上的露水滴湿，头发长得像鹰的羽毛，指甲长得像鸟爪。
DAN|4|34|“时候到了，我－ 尼布甲尼撒 举目望天，我的知识复归于我，我就称颂至高者，赞美尊敬活到永远的上帝。 他的权柄存到永远， 他的国度存到万代。
DAN|4|35|地上所有的居民都算为虚无； 在天上万军和地上居民中， 他都凭自己的旨意行事。 无人能拦住他的手， 或问他说，你在做什么呢？
DAN|4|36|“那时，我的知识复归于我，威严和光荣也复归于我，使我的国度得荣耀，我的谋士和大臣也来朝见我。我又重建我的国度，更大的权势加添在我身上。
DAN|4|37|现在我－ 尼布甲尼撒 赞美、尊崇、恭敬天上的王，因为他所行的全都信实，他所做的尽都公平。那行事骄傲的，他能降为卑。”
DAN|5|1|伯沙撒 王为他的一千大臣摆设盛筵，与这一千人饮酒。
DAN|5|2|伯沙撒 在欢饮之间，吩咐人将他父 尼布甲尼撒 从 耶路撒冷 圣殿所掳掠的金银器皿拿来，好使王与大臣、王后、妃嫔用这器皿饮酒。
DAN|5|3|于是他们把圣殿，就是 耶路撒冷 上帝殿中所掳掠的金器皿拿来，王和大臣、王后、妃嫔就用这器皿饮酒。
DAN|5|4|他们饮酒，赞美金、银、铜、铁、木、石造的神明。
DAN|5|5|当时，忽然有人的指头出现，在灯台对面王宫粉刷的墙上写字。王看见写字的指头，
DAN|5|6|就变了脸色，心意惊惶，腰骨好像脱节，双膝彼此相碰，
DAN|5|7|大声吩咐将巫师、 迦勒底 人和观兆的领进来。王对 巴比伦 的智慧人说：“谁能读这文字，并且向我讲解它的意思，他必身穿紫袍，项带金链，在我国中位列第三。”
DAN|5|8|于是王所有的智慧人都进前来，他们却不能读那文字，也不能为王讲解它的意思。
DAN|5|9|伯沙撒 王就甚惊惶，脸色改变，他的大臣也都困惑。
DAN|5|10|太后 因王和他大臣所说的话，就进入宴会厅，说：“愿王万岁！你的心不要惊惶，脸不要变色。
DAN|5|11|在你国中有一人，他里头有神圣神明的灵，你父在世的日子，这人心中光明，又有聪明智慧，好像神明的智慧。你父 尼布甲尼撒 王，就是王的父，曾立他为术士、巫师、 迦勒底 人和观兆者的领袖，
DAN|5|12|都因他有美好的灵性，又有知识聪明，能解梦，释谜语，解疑惑。这人名叫 但以理 ， 尼布甲尼撒 王又称他为 伯提沙撒 ，现在可以召他来，他必解明这意思。”
DAN|5|13|于是 但以理 被领到王面前。王问 但以理 说：“你就是我父王从 犹大 带来、被掳的 犹大 人 但以理 吗？
DAN|5|14|我听说你里头有神明的灵，心中有光，又有聪明和高超的智慧。
DAN|5|15|现在智慧人和巫师都被带到我面前，要叫他们读这文字，为我讲解它的意思；无奈他们都不能讲解它的意思。
DAN|5|16|我听说你能讲解，能解疑惑；现在你若能读这文字，为我讲解它的意思，就必身穿紫袍，项戴金链，在我国中位列第三。”
DAN|5|17|但以理 回答王说：“你的礼物可以归你自己，你的赏赐可以归给别人；我却要为王读这文字，讲解它的意思。
DAN|5|18|你，王啊，至高的上帝曾将国度、大权、荣耀、威严赐给你父 尼布甲尼撒 ；
DAN|5|19|因上帝所赐给他的大权，各方、各国、各族的人都在他面前恐惧战兢，因他要杀就杀，要人活就活，要升就升，要降就降。
DAN|5|20|但他的心高傲，灵也刚愎，以致行事狂傲，就被革去国度的王位，夺走荣耀。
DAN|5|21|他被赶出离开世人，他的心变为兽心，与野驴同住，吃草如牛，身体被天上的露水滴湿，直到他知道，至高的上帝在人的国中掌权，凭自己的旨意立人治国。
DAN|5|22|伯沙撒 啊，你是他的儿子 ，你虽知道这一切，却不谦卑自己，
DAN|5|23|竟向天上的主自高，差人将他殿中的器皿拿到你面前，你和大臣、王后、妃嫔用这器皿饮酒。你又赞美那不能看、不能听、无知无识，用金、银、铜、铁、木、石造的神明，没有将荣耀归与那手中掌管你气息，管理你一切行动的上帝。
DAN|5|24|于是从他那里显出指头写这文字。
DAN|5|25|“所写的文字是：‘弥尼，弥尼，提客勒，乌法珥新 。’
DAN|5|26|解释是这样：弥尼就是上帝数算你国的年日到此完毕。
DAN|5|27|提客勒就是你被秤在天平上，秤出你的亏欠来。
DAN|5|28|毗勒斯 就是你的国要分裂，归给 玛代 人和 波斯 人。”
DAN|5|29|于是 伯沙撒 下令，人就把紫袍给 但以理 穿上，把金链给他戴在颈项上，又传令使他在国中位列第三。
DAN|5|30|当夜， 迦勒底 王 伯沙撒 被杀。
DAN|5|31|玛代 人 大流士 年六十二岁，取了 迦勒底 国。
DAN|6|1|大流士 随心所愿，立了一百二十个总督，治理全国，
DAN|6|2|又在他们以上立总长三人， 但以理 也在其中；使总督在他们三人面前呈报，免得王受亏损。
DAN|6|3|这 但以理 因有卓越的灵性，超乎其余的总长和总督，王想立他治理全国。
DAN|6|4|那时，总长和总督在治国的事务上寻找 但以理 的把柄，为要控告他；只是找不到任何的把柄和过失，因他忠心办事，毫无错误过失。
DAN|6|5|那些人就说：“我们要找 但以理 的把柄，若不从他上帝的律法中下手，就寻不着。”
DAN|6|6|于是，总长和总督纷纷聚集来见王，说：“ 大流士 王万岁！
DAN|6|7|国中的总长、钦差、总督、谋士和省长彼此商议，求王下旨，立一条禁令，三十天之内，不拘何人，若在王以外，或向神明或向人求什么，就必扔在狮子坑中。
DAN|6|8|王啊，现在求你立这禁令，在这文件上签署，使它不能更改；照 玛代 人和 波斯 人的例，绝不更动。”
DAN|6|9|于是 大流士 王在这禁令的文件上签署。
DAN|6|10|但以理 知道这文件已经签署，就进自己的家，他家楼上的窗户开向 耶路撒冷 。他一天三次，双膝跪着，在他的上帝面前祷告感谢，像平常一样。
DAN|6|11|于是，那些人纷纷聚集，发现 但以理 在他上帝面前祈祷恳求。
DAN|6|12|他们就进到王面前，向王提及禁令，说：“三十天之内不拘何人，若在王以外，或向神明或向人求什么，必被扔在狮子坑中，王不是在这禁令上签署了吗？”王回答说：“确有这事，照 玛代 人和 波斯 人的例是不可更改的。”
DAN|6|13|他们对王说：“王啊，那被掳的 犹大 人 但以理 不理会你，也不遵守你签署的禁令，竟一天三次祈祷。”
DAN|6|14|王听见这话，就甚愁烦，一心要救 但以理 ，直到日落的时候，他还在筹划解救他。
DAN|6|15|那些人就纷纷聚集到王那里，对王说：“王啊，当知道 玛代 人和 波斯 人有例，凡王所立的禁令和律例都不可更改。”
DAN|6|16|于是王下令，人就把 但以理 带来，扔在狮子坑中。王对 但以理 说：“你经常事奉的上帝，他必拯救你。”
DAN|6|17|有人搬来一块石头放在坑口，王用自己的玺和大臣的印，封闭那坑，使惩办 但以理 的事绝不更改。
DAN|6|18|王回到宫里，终夜禁食，不让人带乐器 到他面前，他也失眠了。
DAN|6|19|次日黎明，王起来，急忙往狮子坑那里去，
DAN|6|20|临近坑边，哀声呼叫 但以理 。王对 但以理 说：“永生上帝的仆人 但以理 啊，你经常事奉的上帝能救你脱离狮子吗？”
DAN|6|21|但以理 对王说：“愿王万岁！
DAN|6|22|我的上帝差遣使者封住狮子的口，叫狮子不伤我，因我在上帝面前无辜。王啊，在你面前我也没有做过任何亏损的事。”
DAN|6|23|王因此就甚喜乐，吩咐把 但以理 从坑里拉上来。于是 但以理 从坑里被拉上来，身上毫无损伤，因为他信靠他的上帝。
DAN|6|24|王下令，把那些控告 但以理 的人和他们的妻子儿女都带来，扔在狮子坑中。他们还没有到坑底，狮子就制伏他们，咬碎他们的骨头。
DAN|6|25|于是， 大流士 王传旨给住在全地各方、各国、各族的人说：“愿你们大享平安！
DAN|6|26|现在我降旨，我所统辖全国的人民，都要在 但以理 的上帝面前战兢畏惧。 因为他是活的上帝， 永远长存， 他的国度永不败坏， 他的权柄永存无极！
DAN|6|27|他庇护，搭救， 在天上地下施行神迹奇事， 救了 但以理 脱离狮子的口。”
DAN|6|28|如此，这 但以理 ，当 大流士 在位的时候和 波斯 的 居鲁士 在位的时候，大享亨通。
DAN|7|1|巴比伦 王 伯沙撒 元年， 但以理 在床上做梦，脑中看见异象，就记录这梦，述说其中的大意。
DAN|7|2|但以理 说： 我在夜间的异象中观看，看哪，天上四风，突然刮在大海之上。
DAN|7|3|有四只巨兽从海里上来，它们各不相同：
DAN|7|4|头一个像狮子，有鹰的翅膀；我正观看的时候，它的翅膀被拔去，它从地上被扶起来，用两脚站立，像人一样，还给了它人的心。
DAN|7|5|看哪，另有一兽如熊，就是第二兽，半身侧立，口里的牙齿中有三根獠牙 。有人吩咐这兽说：“起来，吞吃许多的肉。”
DAN|7|6|其后，我观看，看哪，另有一兽如豹，背上有四个鸟的翅膀；这兽有四个头，还给了它权柄。
DAN|7|7|其后，我在夜间的异象中观看，看哪，第四兽可怕可惧，极其强壮，有大铁牙，吞吃嚼碎，剩下的用脚践踏。这兽与前面所有的兽不同，它有十只角。
DAN|7|8|我正思考这些角的时候，看哪，其中又长出另一只小角；先前的角中有三只角在它面前连根被拔出。看哪，这角有眼，像人的眼，有口说夸大的话。
DAN|7|9|我正观看的时候， 有宝座设立， 上面坐着亘古常在者。 他的衣服洁白如雪， 头发如纯净的羊毛。 宝座是火焰， 其轮为烈火。
DAN|7|10|有火如河涌出， 从他面前流出来； 事奉他的有千千， 在他面前侍立的有万万； 他坐着要行审判 ， 案卷都展开了。
DAN|7|11|于是我观看，因这角说夸大的话，我正观看的时候，那兽被杀，身体被毁，扔在火中焚烧。
DAN|7|12|其余的兽，权柄都被夺去，生命却得以延续，直到所定的时候和日期。
DAN|7|13|我在夜间的异象中观看， 看哪，有一位像人子的， 驾着天上的云而来， 被领到亘古常在者面前。
DAN|7|14|他得了权柄、荣耀、国度， 使各方、各国、各族的人都事奉他。 他的权柄是永远的，不能废去， 他的国度必不败坏。
DAN|7|15|至于我－ 但以理 ，我的灵在我里面忧伤，我脑中的异象使我惊惶。
DAN|7|16|我走近其中一位侍立者，问他这一切的实情。他就告诉我，使我知道这事的解释：
DAN|7|17|这四只巨兽就是将要在世上兴起的四个王 。
DAN|7|18|然而，至高者的众圣者必要得到这国度，并且拥有它，直到永远，永永远远。
DAN|7|19|于是我想要更清楚知道第四兽的实情，它与一切的兽不同，甚是可怕，有铁牙铜爪，吞吃嚼碎，剩下的用脚践踏；
DAN|7|20|头上有十只角和那另长出的一角，三只角在这角面前掉落；这角有眼，有口说夸大的话，形状比它的同类更强。
DAN|7|21|我观看，这角与众圣者争战，胜了他们，
DAN|7|22|直到亘古常在者来到，为至高者的众圣者伸冤，众圣者得到国度的时候就到了。
DAN|7|23|那侍立者这样说： 第四兽就是世上要兴起的第四国， 与其他各国不同， 它要并吞全地， 并且践踏嚼碎。
DAN|7|24|至于那十只角，就是从这国中兴起的十个王； 后来又兴起另一王， 与先前的不相同， 他要制伏三个王。
DAN|7|25|他说话抵挡至高者， 折磨至高者的众圣者， 又改变节期和律法。 众圣者要交在他手中一年 、两年、又半年。
DAN|7|26|然而，他坐着要行审判； 他的权柄要被夺去， 毁坏，灭绝，一直到底。
DAN|7|27|国度、权柄和天下诸国的大权 必赐给至高者的众圣民。 他的国是永远的国， 所有掌权的都必事奉他，顺从他。
DAN|7|28|这事到此结束。我－ 但以理 因这些念头甚是惊惶，脸色也变了，却将这事记在心里。
DAN|8|1|伯沙撒 王在位第三年，有异象向我－ 但以理 显现，是在先前所见的异象之后。
DAN|8|2|我在异象中观看，见自己在 以拦 省 书珊 的城堡中；我在异象中又见自己在 乌莱河 边。
DAN|8|3|我举目观看，看哪，有一只公绵羊站在河边，它有两只角，这两角都高，一角高过另一角，后长出来的比较高。
DAN|8|4|我见那公绵羊向西、向北、向南抵撞，没有任何兽在它面前站立得住，没有能逃脱它手的；它任意而行，自高自大。
DAN|8|5|我正思想的时候，看哪，有一只公山羊从西而来，遍行全地，脚不着地。这山羊两眼当中有一只显眼的角。
DAN|8|6|它往我先前所见、站在河边、有双角的公绵羊那里，以猛烈的怒气向它直闯。
DAN|8|7|我见公山羊靠近公绵羊，向它发怒，攻击它，折断它的两角。公绵羊在公山羊面前站立不住；它把公绵羊撞倒在地，用脚践踏，没有能救公绵羊脱离它手的。
DAN|8|8|这公山羊长得极其高大，正强壮的时候，那大角折断了，从角的下面向天的四方 长出四只显眼的角来。
DAN|8|9|从四角中的一角又长出另一只小角，向南、向东、向佳美之地，日渐壮大。
DAN|8|10|它渐壮大，高及诸天万象，把一些天象和星辰摔落在地，用脚践踏。
DAN|8|11|它自高自大 ，自以为高及万象之君，它除掉经常献给君的祭，毁坏君的圣所。
DAN|8|12|因罪过的缘故，有军队和经常献的祭交给它。它把真理抛在地上，任意而行 ，无往不利。
DAN|8|13|我听见有一位圣者说话，又有一位圣者向那说话的圣者说：“这经常献的祭、带来荒凉的罪过、圣所与军队被践踏的异象，要持续到几时呢？”
DAN|8|14|他对我 说：“要到二千三百日，圣所就必洁净 。”
DAN|8|15|我－ 但以理 见了这异象，想要明白其中的意思。看哪，有一位形状像人的站在我面前。
DAN|8|16|我听见 乌莱河 中有人声呼叫说：“ 加百列 啊，要使这人明白这异象。”
DAN|8|17|他就来到我所站的地方。他一来，我就惊慌，脸伏于地。他对我说：“人子啊，你要明白，因为这是关乎末后时期的异象。”
DAN|8|18|他对我说话的时候，我正沉睡，脸伏于地。他就摸我，扶我站起来。
DAN|8|19|他说：“看哪，我要指示你恼怒结束的时候必成的事，因为这是关乎末后指定的时期。
DAN|8|20|你所看见那有双角的公绵羊就是 玛代 王和 波斯 王。
DAN|8|21|那公山羊就是 希腊 王；两眼当中的大角就是第一个王。
DAN|8|22|至于角折断了，又从角的下面长出四只角，意思就是有四个国要从这国兴起，只是权势都不及它。
DAN|8|23|这四国末期，恶贯满盈的时候，必有一王兴起，面貌凶恶，诡计多端。
DAN|8|24|他的权柄极大，却不是因自己的能力；他要施行惊人的毁灭，无往不利，任意而行，又要毁灭强有力的人和众圣民。
DAN|8|25|他用权术使手中的诡计成功；他的心自高自大，趁人无备的时候毁灭多人。他又起来攻击万君之君，至终却非因人的手而遭毁灭。
DAN|8|26|所说二千三百日 的异象是真的，但你要将这异象封住，因为它关乎未来许多的日子。”
DAN|8|27|于是我－ 但以理 昏倒，病了数日，然后起来办理王的事务。我因这异象惊骇不已，但还是不能了解。
DAN|9|1|玛代 族 亚哈随鲁 的儿子 大流士 被立为王，统治 迦勒底 国元年，
DAN|9|2|就是他在位第一年，我－ 但以理 从书上得知，耶和华的话临到 耶利米 先知，论 耶路撒冷 荒凉期满的年数为七十年。
DAN|9|3|我面向主上帝，禁食，披麻蒙灰，恳切祷告祈求。
DAN|9|4|我向耶和华－我的上帝祈祷、认罪，说：“主啊，你是大而可畏的上帝，向爱主、守主诫命的人守约施慈爱。
DAN|9|5|我们犯罪作恶，行恶叛逆，偏离你的诫命典章，
DAN|9|6|没有听从你仆人众先知奉你的名向我们君王、官长、祖先和这地所有百姓所说的话。
DAN|9|7|主啊，你是公义的，但我们 犹大 人和 耶路撒冷 的居民，并你所赶到各国的 以色列 众人，不论远近，因为背叛了你，脸上蒙羞，正如今日一样。
DAN|9|8|耶和华啊，我们和我们的君王、官长、祖先因得罪了你，脸上就都蒙羞。
DAN|9|9|主－我们的上帝是怜悯饶恕人的，我们却违背了他，
DAN|9|10|没有听从耶和华－我们上帝的话，没有遵行他藉仆人众先知向我们颁布的律法。
DAN|9|11|以色列 众人都犯了你的律法，偏离、不听从你的话；因此，你仆人 摩西 律法上所写的诅咒和誓言倾倒在我们身上，因我们得罪了上帝。
DAN|9|12|上帝使大灾祸临到我们，实现了警戒我们和审判我们官长的话；原来 耶路撒冷 所遭遇的灾祸是普天之下未曾有过的。
DAN|9|13|这一切灾祸临到我们，是照 摩西 律法上所写的，我们却没有求耶和华－我们上帝的恩惠，使我们回转离开罪孽，明白你的真理。
DAN|9|14|所以耶和华特意使这灾祸临到我们，耶和华－我们的上帝在他所行的事上都是公义的；我们并没有听从他的话。
DAN|9|15|主－我们的上帝啊，你曾用大能的手领你的子民出 埃及 地，使自己得了名声，正如今日一样，现在，我们犯了罪，作了恶。
DAN|9|16|主啊，求你按你丰盛的公义，使你的怒气和愤怒转离你的城 耶路撒冷 ，就是你的圣山。因我们的罪恶和我们祖先的罪孽， 耶路撒冷 和你的子民被四围的人羞辱。
DAN|9|17|我们的上帝啊，现在求你垂听你仆人的祈祷恳求，为你自己的缘故使你的脸向荒凉的圣所发光。
DAN|9|18|我的上帝啊，求你侧耳而听，睁眼而看，眷顾我们那荒凉之地和称为你名下的城。我们在你面前恳求，不是因自己的义，而是因你丰富的怜悯。
DAN|9|19|主啊，求你垂听！主啊，求你赦免！主啊，求你侧耳，求你实行！为你自己的缘故不要迟延。我的上帝啊，因这城和这民都是称为你名下的。”
DAN|9|20|我正说话、祷告，承认我的罪和我百姓 以色列 的罪，为我上帝的圣山，在耶和华－我的上帝面前恳求；
DAN|9|21|我正在祷告中说话，先前在异象中所见的那位 加百列 ，约在献晚祭的时候迅速飞到我这里来。
DAN|9|22|他指教我说 ：“ 但以理 啊，现在我来要使你有智慧，有聪明。
DAN|9|23|你刚开始恳求的时候，就有命令发出。现在我来告诉你，因你是蒙爱的；所以你要思想这事，明白这异象。
DAN|9|24|“为你百姓和你圣城，已经定了七十个七，要止住罪过，除净罪恶，赎尽罪孽，引进永恒的公义，封住异象和预言，并膏至圣所 。
DAN|9|25|你当知道，当明白，从发出命令恢复并重建 耶路撒冷 ，直到受膏的君出现，必有七个七和六十二个七。 耶路撒冷城 连街带濠都必在艰难中恢复并重建。
DAN|9|26|过了六十二个七，那受膏者 被剪除，一无所有；必有一王的百姓来毁灭这城和圣所，它的结局 必如洪水冲没。必有战争，一直到末了，荒凉的事已经定了。
DAN|9|27|在一七之期，他必与许多人坚立盟约；一七之半，他必使献祭与供献止息。那施行毁灭的可憎之物必立在圣殿里 ，直到所定的结局倾倒在那行毁灭者的身上。”
DAN|10|1|波斯 王 居鲁士 第三年，有话指示那称为 伯提沙撒 的 但以理 。这话是确实的，指着大战争； 但以理 明白这话，明白这异象。
DAN|10|2|那时，我－ 但以理 悲伤了三个七日；
DAN|10|3|美味我没有吃，酒和肉没有入我的口，也没有用油抹我的身，直到满了三个七日。
DAN|10|4|正月二十四日，我在 大河 ，就是 底格里斯河 边，
DAN|10|5|举目观看，看哪，有一人身穿细麻衣，腰束 乌法 的纯金腰带。
DAN|10|6|他的身体如水苍玉，面貌如闪电，眼目如火把，手臂和脚如明亮的铜，说话的声音像众人的声音。
DAN|10|7|我－ 但以理 一人看见这异象，跟我一起的人没有看见，却有极大的战兢落在他们身上，他们就逃跑躲避，
DAN|10|8|只剩下我一人。我看见这大异象就浑身无力，面容变色，毫无气力。
DAN|10|9|我听见他说话的声音；一听见他说话的声音，我就沉睡，脸伏于地。
DAN|10|10|看哪，有一只手摸我，使我膝盖和手掌战抖。
DAN|10|11|他对我说：“蒙爱的 但以理 啊，要思想我对你所说的话，只管站起来，因为我现在奉差遣来到你这里。”他对我说这话，我就战战兢兢地站起来。
DAN|10|12|他说：“ 但以理 啊，不要惧怕！因为自从第一日你立志要明白，又在你上帝面前刻苦自己，你的话已蒙应允；我就是因你的话而来。
DAN|10|13|但 波斯 国的领袖拦阻了我二十一天。看哪，天使长 中的一位 米迦勒 来帮助我，因为我被留在 波斯 诸王那里。
DAN|10|14|现在我来，要使你明白你百姓日后必遭遇的事，因为这异象关乎未来的日子。”
DAN|10|15|他向我这样说，我就脸面朝地，哑口无声。
DAN|10|16|看哪，有一位形状像人的，摸我的嘴唇，我就开口说话，向那站在我面前的说：“我主啊，因这异象使我感到剧痛，毫无气力。
DAN|10|17|我主的仆人怎能跟我主说话呢？我现在浑身无力，毫无气息。”
DAN|10|18|有一位形状像人的再一次摸我，使我有力量。
DAN|10|19|他说：“蒙爱的人哪，不要惧怕，愿你平安！你要刚强！要刚强！ ”他一对我说话，我就觉得有力量，说：“我主请说，因你使我有力量。”
DAN|10|20|他说：“你知道我为什么到你这里来吗？现在我要回去与 波斯 的领袖争战，我去了之后，看哪， 希腊 的领袖必来。
DAN|10|21|但我要将那记录在真理之书上的话告诉你。除了你们的天使 米迦勒 之外，没有人帮助我抵挡他们。”
DAN|11|1|“至于我，当 玛代 的 大流士 元年，我曾起来扶助 米迦勒 ，使他坚强。
DAN|11|2|现在我要指示你确实的事。” “看哪， 波斯 还有三个王要兴起，第四王必富足远胜诸王。他因富足成为强盛，就煽动各国攻击 希腊 国。
DAN|11|3|必有一个勇敢的王兴起，执掌大权，随意而行。
DAN|11|4|他正兴起的时候，他的国必瓦解，向天的四方 裂开，却不归他的后裔，也不如他当年统治的权威；他的国必被拔出，归给他后裔之外的人。
DAN|11|5|“南方的王必强盛，他的将帅中必有一个比他更强，执掌权柄，权柄甚大。
DAN|11|6|过了几年，他们必结盟，南方王的女儿必来到北方王那里，使约生效；但这女子不能保留实力，王的力量 也未能存留。这女子、带她来的、生她的 和当时扶助她的必被杀害 。
DAN|11|7|但从这女子的本家必另有一子 接续王位，他要率领军队进入北方王的堡垒，攻击他们，而且得胜，
DAN|11|8|把他们的神像和铸成的偶像，与金银宝器都掳掠到 埃及 去。数年之内，他不去攻击北方的王。
DAN|11|9|北方的王必侵入南方王的国土，但却要撤回本地。
DAN|11|10|“北方王的儿子们必动干戈，招聚许多军兵。他要前进，如洪水泛滥；要再度争战，直捣南方王的堡垒。
DAN|11|11|南方王必发烈怒，出来与北方王争战，摆列大军；北方王的军兵必败在南方王的手下。
DAN|11|12|这大军既被扫荡，南方王的心就自高；他虽使万人仆倒，却不能保持胜利。
DAN|11|13|“北方王要再度摆列大军，比先前更多。过了几年，他必率领大军，带极多的装备而来。
DAN|11|14|那时，必有许多人起来攻击南方王，并且你百姓中的残暴人要兴起，应验异象，他们却要败亡。
DAN|11|15|北方王必来建土堆攻取坚固城，南方的军兵抵挡不住，就是精选的部队也无力抵挡；
DAN|11|16|前来攻击南方王的必任意而行，无人在北方王面前站立得住。他要站在那佳美之地，用手施行毁灭。
DAN|11|17|“他必定意倾全国之力而来，与南方王订约，把自己的女儿 给南方王为妻，企图败坏他的国度。这计谋却未得逞，自己也得不到好处。
DAN|11|18|其后北方王必转头，夺取许多海岛。但有一将帅除掉北方王对人的羞辱，并且使羞辱归到他自己身上。
DAN|11|19|他必转头回到本地的堡垒，却要绊跌仆倒，归于无有。
DAN|11|20|“那时，有一人兴起接续他的王位，他为了王国的荣华，差官员横征暴敛。这王过不多时就死了，不是因怒气 ，也不是因战役。”
DAN|11|21|“后来，有一个卑鄙的人兴起接续他的王位，人未曾将国的尊荣给他，他却趁人无备的时候前来，用诡诈夺取政权。
DAN|11|22|势如洪水般的军兵在他面前被冲没，遭击溃；立约的领袖也是如此。
DAN|11|23|他与人结盟之后，却行诡诈。跟随他的人虽不多，他却日渐强盛。
DAN|11|24|他趁人无备的时候，来到国中极肥沃之地，做他祖宗和祖宗的祖宗未曾做过的事，瓜分掳物、掠物和财宝，又策划进攻堡垒；然而这都是暂时的。
DAN|11|25|“他必奋勇向前，率领大军攻击南方王；南方王以极强的大军迎战，却抵挡不住，因为有人设计谋害南方王。
DAN|11|26|吃王饷的使王败坏，王的军队必被冲没，仆倒被杀的甚多。
DAN|11|27|至于这二王，他们心怀恶计，同席吃饭却彼此说谎，但计谋不成，因为结局要在指定的时期来到。
DAN|11|28|北方王必带许多财宝回本地，但他的心反对圣约；他恣意横行，回到本地。
DAN|11|29|“到了指定的时期，他必返回，侵入南方。这一次却不像前一次，
DAN|11|30|因为 基提 的战船要来攻击他，他就丧胆而退。他恼恨圣约，恣意横行，要回来善待那些背弃圣约的人。
DAN|11|31|他要兴兵，这兵必亵渎圣所，就是堡垒，除掉经常献的祭，设立那施行毁灭的可憎之物。
DAN|11|32|他必用巧言奉承违背圣约的恶人；惟独认识上帝的子民必刚强行事。
DAN|11|33|民间的智慧人必训诲许多人，然而在一段日子里，他们必因刀剑、火烧、掳掠、抢夺而仆倒。
DAN|11|34|他们仆倒的时候，会得到少许援助，却有许多人用诡诈加入他们。
DAN|11|35|智慧人中有些人仆倒，为要使他们受熬炼，成为洁净、洁白，直到末了；因为还有一段日子才到所定的时期。
DAN|11|36|“王必任意而行，自高自大，超过所有的神明，又用荒谬的话攻击万神之神。他必行事亨通，直到主的愤怒结束，因为所定的事必然实现。
DAN|11|37|他不顾他祖宗的神明，也不顾妇女所仰慕的神明，任何神明他都不顾；因为他自大，高过一切，
DAN|11|38|以敬奉堡垒的神明取而代之，用金、银、宝石和珍宝敬奉他祖宗所不认识的神明。
DAN|11|39|他靠外邦神明的帮助，攻破最坚固的堡垒。凡承认他的，他要给他们许多尊荣，使他们管辖许多人，又分封土地作为报偿。
DAN|11|40|“到末了，南方王要与北方王交战。北方王要用战车、骑兵和许多战船，势如暴风来攻击他，又要侵入列国，如洪水泛滥。
DAN|11|41|他要侵入那佳美之地，许多国就被倾覆 ，但 以东 人、 摩押 人和大半的 亚扪 人必逃离他的手。
DAN|11|42|他要伸手攻击列国，连 埃及 地也不得逃脱。
DAN|11|43|他要掌管 埃及 的金银财宝和各样珍宝， 路比 人和 古实 人都跟从他的脚步。
DAN|11|44|但从东方和北方必有消息传来扰乱他，他就大发烈怒出去，要将许多人杀灭净尽。
DAN|11|45|他要在海和荣美的圣山之间搭起王宫的帐幕；然而他的结局到了，无人能帮助他。”
DAN|12|1|“那时，保佑你百姓的天使长 米迦勒 必站起来，并且有大艰难，自从有国以来直到此时，未曾有过这样的事。那时，你的百姓凡记录在册上的，必得拯救。
DAN|12|2|睡在地里尘埃中的必有多人醒过来；其中有得永生的，有受羞辱永远被憎恶的。
DAN|12|3|智慧人要发光，如同天上的光；那领许多人归于义的必发光如星，直到永永远远。
DAN|12|4|但以理 啊，你要隐藏这话，封闭这书，直到末时。必有许多人往来奔跑 ，知识 就必增长。”
DAN|12|5|我－ 但以理 观看，看哪，另有两个人站立：一个在河这边，一个在河那边。
DAN|12|6|其中一个对那在河水之上、穿细麻衣的说：“这奇异的事要到几时才应验呢？”
DAN|12|7|我听见那在河水之上、穿细麻衣的，向天举起左右手，指着那活到永远的起誓说：“要到一年 、两年，又半年，粉碎圣民力量结束的时候，这一切的事就要应验。”
DAN|12|8|我听了却不明白，就说：“我主啊，这些事的结局是怎样呢？”
DAN|12|9|他说：“ 但以理 ，去吧！因为这话已经隐藏封闭，直到末时。
DAN|12|10|必有许多人使自己洁净、洁白，且受熬炼；但恶人仍必行恶，没有一个恶人明白，惟独智慧人能明白。
DAN|12|11|从除掉经常献的祭，设立那施行毁灭的可憎之物的时候起，必有一千二百九十日。
DAN|12|12|那等候，直到一千三百三十五日的有福了。
DAN|12|13|“至于你，你要去等候结局。你必安息，到了末期，你必起来，享受你的福分。”
