1THESS|1|1|Paulus et Silvanus et Timotheus ecclesiae Thessalonicensium in Deo Patre et Domino Iesu Christo gratia vobis et pax
1THESS|1|2|gratias agimus Deo semper pro omnibus vobis memoriam facientes in orationibus nostris sine intermissione
1THESS|1|3|memores operis fidei vestrae et laboris et caritatis et sustinentiae spei Domini nostri Iesu Christi ante Deum et Patrem nostrum
1THESS|1|4|scientes fratres dilecti a Deo electionem vestram
1THESS|1|5|quia evangelium nostrum non fuit ad vos in sermone tantum sed et in virtute et in Spiritu Sancto et in plenitudine multa sicut scitis quales fuerimus vobis propter vos
1THESS|1|6|et vos imitatores nostri facti estis et Domini excipientes verbum in tribulatione multa cum gaudio Spiritus Sancti
1THESS|1|7|ita ut facti sitis forma omnibus credentibus in Macedonia et in Achaia
1THESS|1|8|a vobis enim diffamatus est sermo Domini non solum in Macedonia et in Achaia sed in omni loco fides vestra quae est ad Deum profecta est ita ut non sit nobis necesse quicquam loqui
1THESS|1|9|ipsi enim de nobis adnuntiant qualem introitum habuerimus ad vos et quomodo conversi estis ad Deum a simulacris servire Deo vivo et vero
1THESS|1|10|et expectare Filium eius de caelis quem suscitavit ex mortuis Iesum qui eripuit nos ab ira ventura
1THESS|2|1|nam ipsi scitis fratres introitum nostrum ad vos quia non inanis fuit
1THESS|2|2|sed ante passi et contumeliis affecti sicut scitis in Philippis fiduciam habuimus in Deo nostro loqui ad vos evangelium Dei in multa sollicitudine
1THESS|2|3|exhortatio enim nostra non de errore neque de inmunditia neque in dolo
1THESS|2|4|sed sicut probati sumus a Deo ut crederetur nobis evangelium ita loquimur non quasi hominibus placentes sed Deo qui probat corda nostra
1THESS|2|5|neque enim aliquando fuimus in sermone adulationis sicut scitis neque in occasione avaritiae Deus testis est
1THESS|2|6|nec quaerentes ab hominibus gloriam neque a vobis neque ab aliis
1THESS|2|7|cum possimus oneri esse ut Christi apostoli sed facti sumus lenes in medio vestrum tamquam si nutrix foveat filios suos
1THESS|2|8|ita desiderantes vos cupide volebamus tradere vobis non solum evangelium Dei sed etiam animas nostras quoniam carissimi nobis facti estis
1THESS|2|9|memores enim estis fratres laborem nostrum et fatigationem nocte et die operantes ne quem vestrum gravaremus praedicavimus in vobis evangelium Dei
1THESS|2|10|vos testes estis et Deus quam sancte et iuste et sine querella vobis qui credidistis fuimus
1THESS|2|11|sicut scitis qualiter unumquemque vestrum tamquam pater filios suos
1THESS|2|12|deprecantes vos et consolantes testificati sumus ut ambularetis digne Deo qui vocavit vos in suum regnum et gloriam
1THESS|2|13|ideo et nos gratias agimus Deo sine intermissione quoniam cum accepissetis a nobis verbum auditus Dei accepistis non ut verbum hominum sed sicut est vere verbum Dei qui operatur in vobis qui credidistis
1THESS|2|14|vos enim imitatores facti estis fratres ecclesiarum Dei quae sunt in Iudaea in Christo Iesu quia eadem passi estis et vos a contribulibus vestris sicut et ipsi a Iudaeis
1THESS|2|15|qui et Dominum occiderunt Iesum et prophetas et nos persecuti sunt et Deo non placent et omnibus hominibus adversantur
1THESS|2|16|prohibentes nos gentibus loqui ut salvae fiant ut impleant peccata sua semper praevenit autem ira Dei super illos usque in finem
1THESS|2|17|nos autem fratres desolati a vobis ad tempus horae aspectu non corde abundantius festinavimus faciem vestram videre cum multo desiderio
1THESS|2|18|quoniam voluimus venire ad vos ego quidem Paulus et semel et iterum et inpedivit nos Satanas
1THESS|2|19|quae est enim nostra spes aut gaudium aut corona gloriae nonne vos ante Dominum nostrum Iesum estis in adventu eius
1THESS|2|20|vos enim estis gloria nostra et gaudium
1THESS|3|1|propter quod non sustinentes amplius placuit nobis remanere Athenis solis
1THESS|3|2|et misimus Timotheum fratrem nostrum et ministrum Dei in evangelio Christi ad confirmandos vos et exhortandos pro fide vestra
1THESS|3|3|ut nemo moveatur in tribulationibus istis ipsi enim scitis quod in hoc positi sumus
1THESS|3|4|nam et cum apud vos essemus praedicebamus vobis passuros nos tribulationes sicut et factum est et scitis
1THESS|3|5|propterea et ego amplius non sustinens misi ad cognoscendam fidem vestram ne forte temptaverit vos is qui temptat et inanis fiat labor noster
1THESS|3|6|nunc autem veniente Timotheo ad nos a vobis et adnuntiante nobis fidem et caritatem vestram et quia memoriam nostri habetis bonam semper desiderantes nos videre sicut nos quoque vos
1THESS|3|7|ideo consolati sumus fratres in vobis in omni necessitate et tribulatione nostra per vestram fidem
1THESS|3|8|quoniam nunc vivimus si vos statis in Domino
1THESS|3|9|quam enim gratiarum actionem possumus Deo retribuere pro vobis in omni gaudio quo gaudemus propter vos ante Deum nostrum
1THESS|3|10|nocte et die abundantius orantes ut videamus faciem vestram et conpleamus ea quae desunt fidei vestrae
1THESS|3|11|ipse autem Deus et Pater noster et Dominus Iesus dirigat viam nostram ad vos
1THESS|3|12|vos autem Dominus multiplicet et abundare faciat caritatem in invicem et in omnes quemadmodum et nos in vobis
1THESS|3|13|ad confirmanda corda vestra sine querella in sanctitate ante Deum et Patrem nostrum in adventu Domini nostri Iesu cum omnibus sanctis eius amen
1THESS|4|1|de cetero ergo fratres rogamus vos et obsecramus in Domino Iesu ut quemadmodum accepistis a nobis quomodo vos oporteat ambulare et placere Deo sicut et ambulatis ut abundetis magis
1THESS|4|2|scitis enim quae praecepta dederimus vobis per Dominum Iesum
1THESS|4|3|haec est enim voluntas Dei sanctificatio vestra
1THESS|4|4|ut abstineatis vos a fornicatione ut sciat unusquisque vestrum suum vas possidere in sanctificatione et honore
1THESS|4|5|non in passione desiderii sicut et gentes quae ignorant Deum
1THESS|4|6|ut ne quis supergrediatur neque circumveniat in negotio fratrem suum quoniam vindex est Dominus de his omnibus sicut et praediximus vobis et testificati sumus
1THESS|4|7|non enim vocavit nos Deus in inmunditia sed in sanctificatione
1THESS|4|8|itaque qui spernit non hominem spernit sed Deum qui etiam dedit Spiritum suum Sanctum in vobis
1THESS|4|9|de caritate autem fraternitatis non necesse habemus scribere vobis ipsi enim vos a Deo didicistis ut diligatis invicem
1THESS|4|10|etenim facitis illud in omnes fratres in universa Macedonia rogamus autem vos fratres ut abundetis magis
1THESS|4|11|et operam detis ut quieti sitis et ut vestrum negotium agatis et operemini manibus vestris sicut praecepimus vobis
1THESS|4|12|et ut honeste ambuletis ad eos qui foris sunt et nullius aliquid desideretis
1THESS|4|13|nolumus autem vos ignorare fratres de dormientibus ut non contristemini sicut et ceteri qui spem non habent
1THESS|4|14|si enim credimus quod Iesus mortuus est et resurrexit ita et Deus eos qui dormierunt per Iesum adducet cum eo
1THESS|4|15|hoc enim vobis dicimus in verbo Domini quia nos qui vivimus qui residui sumus in adventum Domini non praeveniemus eos qui dormierunt
1THESS|4|16|quoniam ipse Dominus in iussu et in voce archangeli et in tuba Dei descendet de caelo et mortui qui in Christo sunt resurgent primi
1THESS|4|17|deinde nos qui vivimus qui relinquimur simul rapiemur cum illis in nubibus obviam Domino in aera et sic semper cum Domino erimus
1THESS|4|18|itaque consolamini invicem in verbis istis
1THESS|5|1|de temporibus autem et momentis fratres non indigetis ut scribamus vobis
1THESS|5|2|ipsi enim diligenter scitis quia dies Domini sicut fur in nocte ita veniet
1THESS|5|3|cum enim dixerint pax et securitas tunc repentinus eis superveniet interitus sicut dolor in utero habenti et non effugient
1THESS|5|4|vos autem fratres non estis in tenebris ut vos dies ille tamquam fur conprehendat
1THESS|5|5|omnes enim vos filii lucis estis et filii diei non sumus noctis neque tenebrarum
1THESS|5|6|igitur non dormiamus sicut ceteri sed vigilemus et sobrii simus
1THESS|5|7|qui enim dormiunt nocte dormiunt et qui ebrii sunt nocte ebrii sunt
1THESS|5|8|nos autem qui diei sumus sobrii simus induti loricam fidei et caritatis et galeam spem salutis
1THESS|5|9|quoniam non posuit nos Deus in iram sed in adquisitionem salutis per Dominum nostrum Iesum Christum
1THESS|5|10|qui mortuus est pro nobis ut sive vigilemus sive dormiamus simul cum illo vivamus
1THESS|5|11|propter quod consolamini invicem et aedificate alterutrum sicut et facitis
1THESS|5|12|rogamus autem vos fratres ut noveritis eos qui laborant inter vos et praesunt vobis in Domino et monent vos
1THESS|5|13|ut habeatis illos abundantius in caritate propter opus illorum pacem habete cum eis
1THESS|5|14|rogamus autem vos fratres corripite inquietos consolamini pusillianimes suscipite infirmos patientes estote ad omnes
1THESS|5|15|videte ne quis malum pro malo alicui reddat sed semper quod bonum est sectamini et in invicem et in omnes
1THESS|5|16|semper gaudete
1THESS|5|17|sine intermissione orate
1THESS|5|18|in omnibus gratias agite haec enim voluntas Dei est in Christo Iesu in omnibus vobis
1THESS|5|19|Spiritum nolite extinguere
1THESS|5|20|prophetias nolite spernere
1THESS|5|21|omnia autem probate quod bonum est tenete
1THESS|5|22|ab omni specie mala abstinete vos
1THESS|5|23|ipse autem Deus pacis sanctificet vos per omnia et integer spiritus vester et anima et corpus sine querella in adventu Domini nostri Iesu Christi servetur
1THESS|5|24|fidelis est qui vocavit vos qui etiam faciet
1THESS|5|25|fratres orate pro nobis
1THESS|5|26|salutate fratres omnes in osculo sancto
1THESS|5|27|adiuro vos per Dominum ut legatur epistula omnibus sanctis fratribus
1THESS|5|28|gratia Domini nostri Iesu Christi vobiscum amen
