ISA|1|1|Видение Исаии, сына Амосова, которое он видел о Иудее и Иерусалиме, во дни Озии, Иоафама, Ахаза, Езекии – царей Иудейских.
ISA|1|2|Слушайте, небеса, и внимай, земля, потому что Господь говорит: Я воспитал и возвысил сыновей, а они возмутились против Меня.
ISA|1|3|Вол знает владетеля своего, и осел – ясли господина своего; а Израиль не знает [Меня], народ Мой не разумеет.
ISA|1|4|Увы, народ грешный, народ обремененный беззакониями, племя злодеев, сыны погибельные! Оставили Господа, презрели Святаго Израилева, – повернулись назад.
ISA|1|5|Во что вас бить еще, продолжающие свое упорство? Вся голова в язвах, и все сердце исчахло.
ISA|1|6|От подошвы ноги до темени головы нет у него здорового места: язвы, пятна, гноящиеся раны, неочищенные и необвязанные и не смягченные елеем.
ISA|1|7|Земля ваша опустошена; города ваши сожжены огнем; поля ваши в ваших глазах съедают чужие; все опустело, как после разорения чужими.
ISA|1|8|И осталась дщерь Сиона, как шатер в винограднике, как шалаш в огороде, как осажденный город.
ISA|1|9|Если бы Господь Саваоф не оставил нам небольшого остатка, то мы были бы то же, что Содом, уподобились бы Гоморре.
ISA|1|10|Слушайте слово Господне, князья Содомские; внимай закону Бога нашего, народ Гоморрский!
ISA|1|11|К чему Мне множество жертв ваших? говорит Господь. Я пресыщен всесожжениями овнов и туком откормленного скота, и крови тельцов и агнцев и козлов не хочу.
ISA|1|12|Когда вы приходите являться пред лице Мое, кто требует от вас, чтобы вы топтали дворы Мои?
ISA|1|13|Не носите больше даров тщетных: курение отвратительно для Меня; новомесячий и суббот, праздничных собраний не могу терпеть: беззаконие – и празднование!
ISA|1|14|Новомесячия ваши и праздники ваши ненавидит душа Моя: они бремя для Меня; Мне тяжело нести их.
ISA|1|15|И когда вы простираете руки ваши, Я закрываю от вас очи Мои; и когда вы умножаете моления ваши, Я не слышу: ваши руки полны крови.
ISA|1|16|Омойтесь, очиститесь; удалите злые деяния ваши от очей Моих; перестаньте делать зло;
ISA|1|17|научитесь делать добро, ищите правды, спасайте угнетенного, защищайте сироту, вступайтесь за вдову.
ISA|1|18|Тогда придите – и рассудим, говорит Господь. Если будут грехи ваши, как багряное, – как снег убелю; если будут красны, как пурпур, – как волну убелю.
ISA|1|19|Если захотите и послушаетесь, то будете вкушать блага земли;
ISA|1|20|если же отречетесь и будете упорствовать, то меч пожрет вас: ибо уста Господни говорят.
ISA|1|21|Как сделалась блудницею верная столица, исполненная правосудия! Правда обитала в ней, а теперь – убийцы.
ISA|1|22|Серебро твое стало изгарью, вино твое испорчено водою;
ISA|1|23|князья твои – законопреступники и сообщники воров; все они любят подарки и гоняются за мздою; не защищают сироты, и дело вдовы не доходит до них.
ISA|1|24|Посему говорит Господь, Господь Саваоф, Сильный Израилев: о, удовлетворю Я Себя над противниками Моими и отмщу врагам Моим!
ISA|1|25|И обращу на тебя руку Мою и, как в щелочи, очищу с тебя примесь, и отделю от тебя все свинцовое;
ISA|1|26|и опять буду поставлять тебе судей, как прежде, и советников, как вначале; тогда будут говорить о тебе: "город правды, столица верная".
ISA|1|27|Сион спасется правосудием, и обратившиеся [сыны] его – правдою;
ISA|1|28|всем же отступникам и грешникам – погибель, и оставившие Господа истребятся.
ISA|1|29|Они будут постыжены за дубравы, которые столь вожделенны для вас, и посрамлены за сады, которые вы избрали себе;
ISA|1|30|ибо вы будете, как дуб, [которого] лист опал, и как сад, в котором нет воды.
ISA|1|31|И сильный будет отрепьем, и дело его – искрою; и будут гореть вместе, – и никто не потушит.
ISA|2|1|Слово, которое было в видении к Исаии, сыну Амосову, о Иудее и Иерусалиме.
ISA|2|2|И будет в последние дни, гора дома Господня будет поставлена во главу гор и возвысится над холмами, и потекут к ней все народы.
ISA|2|3|И пойдут многие народы и скажут: придите, и взойдем на гору Господню, в дом Бога Иаковлева, и научит Он нас Своим путям и будем ходить по стезям Его; ибо от Сиона выйдет закон, и слово Господне – из Иерусалима.
ISA|2|4|И будет Он судить народы, и обличит многие племена; и перекуют мечи свои на орала, и копья свои – на серпы: не поднимет народ на народ меча, и не будут более учиться воевать.
ISA|2|5|О, дом Иакова! Придите, и будем ходить во свете Господнем.
ISA|2|6|Но Ты отринул народ Твой, дом Иакова, потому что они многое переняли от востока: и чародеи [у них], как у Филистимлян, и с сынами чужих они в общении.
ISA|2|7|И наполнилась земля его серебром и золотом, и нет числа сокровищам его; и наполнилась земля его конями, и нет числа колесницам его;
ISA|2|8|и наполнилась земля его идолами: они поклоняются делу рук своих, тому, что сделали персты их.
ISA|2|9|И преклонился человек, и унизился муж, – и Ты не простишь их.
ISA|2|10|Иди в скалу и сокройся в землю от страха Господа и от славы величия Его.
ISA|2|11|Поникнут гордые взгляды человека, и высокое людское унизится; и один Господь будет высок в тот день.
ISA|2|12|Ибо [грядет] день Господа Саваофа на все гордое и высокомерное и на все превознесенное, – и оно будет унижено, –
ISA|2|13|и на все кедры Ливанские, высокие и превозносящиеся, и на все дубы Васанские,
ISA|2|14|и на все высокие горы, и на все возвышающиеся холмы,
ISA|2|15|и на всякую высокую башню, и на всякую крепкую стену,
ISA|2|16|и на все корабли Фарсисские, и на все вожделенные украшения их.
ISA|2|17|И падет величие человеческое, и высокое людское унизится; и один Господь будет высок в тот день,
ISA|2|18|и идолы совсем исчезнут.
ISA|2|19|И войдут [люди] в расселины скал и в пропасти земли от страха Господа и от славы величия Его, когда Он восстанет сокрушить землю.
ISA|2|20|В тот день человек бросит кротам и летучим мышам серебряных своих идолов и золотых своих идолов, которых сделал себе для поклонения им,
ISA|2|21|чтобы войти в ущелья скал и в расселины гор от страха Господа и от славы величия Его, когда Он восстанет сокрушить землю.
ISA|2|22|Перестаньте вы надеяться на человека, которого дыхание в ноздрях его, ибо что он значит?
ISA|3|1|Вот, Господь, Господь Саваоф, отнимет у Иерусалима и у Иуды посох и трость, всякое подкрепление хлебом и всякое подкрепление водою,
ISA|3|2|храброго вождя и воина, судью и пророка, и прозорливца и старца,
ISA|3|3|пятидесятника и вельможу и советника, и мудрого художника и искусного в слове.
ISA|3|4|И дам им отроков в начальники, и дети будут господствовать над ними.
ISA|3|5|И в народе один будет угнетаем другим, и каждый – ближним своим; юноша будет нагло превозноситься над старцем, и простолюдин над вельможею.
ISA|3|6|Тогда ухватится человек за брата своего, в семействе отца своего, [и скажет]: у тебя [есть] одежда, будь нашим вождем, и да будут эти развалины под рукою твоею.
ISA|3|7|А [он] с клятвою скажет: не могу исцелить [ран общества]; и в моем доме нет ни хлеба, ни одежды; не делайте меня вождем народа.
ISA|3|8|Так рушился Иерусалим, и пал Иуда, потому что язык их и дела их – против Господа, оскорбительны для очей славы Его.
ISA|3|9|Выражение лиц их свидетельствует против них, и о грехе своем они рассказывают открыто, как Содомляне, не скрывают: горе душе их! ибо сами на себя навлекают зло.
ISA|3|10|Скажите праведнику, что благо [ему], ибо он будет вкушать плоды дел своих;
ISA|3|11|а беззаконнику – горе, ибо будет ему возмездие за [дела] рук его.
ISA|3|12|Притеснители народа Моего – дети, и женщины господствуют над ним. Народ Мой! вожди твои вводят тебя в заблуждение и путь стезей твоих испортили.
ISA|3|13|Восстал Господь на суд – и стоит, чтобы судить народы.
ISA|3|14|Господь вступает в суд со старейшинами народа Своего и с князьями его: вы опустошили виноградник; награбленное у бедного – в ваших домах;
ISA|3|15|что вы тесните народ Мой и угнетаете бедных? говорит Господь, Господь Саваоф.
ISA|3|16|И сказал Господь: за то, что дочери Сиона надменны и ходят, подняв шею и обольщая взорами, и выступают величавою поступью и гремят цепочками на ногах, –
ISA|3|17|оголит Господь темя дочерей Сиона и обнажит Господь срамоту их;
ISA|3|18|в тот день отнимет Господь красивые цепочки на ногах и звездочки, и луночки,
ISA|3|19|серьги, и ожерелья, и опахала, увясла и запястья, и пояса, и сосудцы с духами, и привески волшебные,
ISA|3|20|перстни и кольца в носу,
ISA|3|21|верхнюю одежду и нижнюю, и платки, и кошельки,
ISA|3|22|светлые тонкие епанчи и повязки, и покрывала.
ISA|3|23|И будет вместо благовония зловоние, и вместо пояса будет веревка, и вместо завитых волос – плешь, и вместо широкой епанчи – узкое вретище, вместо красоты – клеймо.
ISA|3|24|Мужи твои падут от меча, и храбрые твои – на войне.
ISA|3|25|И будут воздыхать и плакать ворота [столицы],
ISA|3|26|и будет она сидеть на земле опустошенная.
ISA|4|1|И ухватятся семь женщин за одного мужчину в тот день, и скажут: "свой хлеб будем есть и свою одежду будем носить, только пусть будем называться твоим именем, – сними с нас позор".
ISA|4|2|В тот день отрасль Господа явится в красоте и чести, и плод земли – в величии и славе, для уцелевших [сынов] Израиля.
ISA|4|3|Тогда оставшиеся на Сионе и уцелевшие в Иерусалиме будут именоваться святыми, все вписанные в книгу для житья в Иерусалиме,
ISA|4|4|когда Господь омоет скверну дочерей Сиона и очистит кровь Иерусалима из среды его духом суда и духом огня.
ISA|4|5|И сотворит Господь над всяким местом горы Сиона и над собраниями ее облако и дым во время дня и блистание пылающего огня во время ночи; ибо над всем чтимым будет покров.
ISA|4|6|И будет шатер для осенения днем от зноя и для убежища и защиты от непогод и дождя.
ISA|5|1|Воспою Возлюбленному моему песнь Возлюбленного моего о винограднике Его. У Возлюбленного моего был виноградник на вершине утучненной горы,
ISA|5|2|и Он обнес его оградою, и очистил его от камней, и насадил в нем отборные виноградные лозы, и построил башню посреди его, и выкопал в нем точило, и ожидал, что он принесет добрые грозды, а он принес дикие ягоды.
ISA|5|3|И ныне, жители Иерусалима и мужи Иуды, рассудите Меня с виноградником Моим.
ISA|5|4|Что еще надлежало бы сделать для виноградника Моего, чего Я не сделал ему? Почему, когда Я ожидал, что он принесет добрые грозды, он принес дикие ягоды?
ISA|5|5|Итак Я скажу вам, что сделаю с виноградником Моим: отниму у него ограду, и будет он опустошаем; разрушу стены его, и будет попираем,
ISA|5|6|и оставлю его в запустении: не будут ни обрезывать, ни вскапывать его, – и зарастет он тернами и волчцами, и повелю облакам не проливать на него дождя.
ISA|5|7|Виноградник Господа Саваофа есть дом Израилев, и мужи Иуды – любимое насаждение Его. И ждал Он правосудия, но вот – кровопролитие; [ждал] правды, и вот – вопль.
ISA|5|8|Горе вам, прибавляющие дом к дому, присоединяющие поле к полю, так что [другим] не остается места, как будто вы одни поселены на земле.
ISA|5|9|В уши мои [сказал] Господь Саваоф: многочисленные домы эти будут пусты, большие и красивые – без жителей;
ISA|5|10|десять участков в винограднике дадут один бат, и хомер посеянного зерна едва принесет ефу.
ISA|5|11|Горе тем, которые с раннего утра ищут сикеры и до позднего вечера разгорячают себя вином;
ISA|5|12|и цитра и гусли, тимпан и свирель и вино на пиршествах их; а на дела Господа они не взирают и о деяниях рук Его не помышляют.
ISA|5|13|За то народ мой пойдет в плен непредвиденно, и вельможи его будут голодать, и богачи его будут томиться жаждою.
ISA|5|14|За то преисподняя расширилась и без меры раскрыла пасть свою: и сойдет [туда] слава их и богатство их, и шум их и [все], что веселит их.
ISA|5|15|И преклонится человек, и смирится муж, и глаза гордых поникнут;
ISA|5|16|а Господь Саваоф превознесется в суде, и Бог Святый явит святость Свою в правде.
ISA|5|17|И будут пастись овцы по своей воле, и чужие будут питаться оставленными жирными пажитями богатых.
ISA|5|18|Горе тем, которые влекут на себя беззаконие вервями суетности, и грех – как бы ремнями колесничными;
ISA|5|19|которые говорят: "пусть Он поспешит и ускорит дело Свое, чтобы мы видели, и пусть приблизится и придет в исполнение совет Святаго Израилева, чтобы мы узнали!"
ISA|5|20|Горе тем, которые зло называют добром, и добро – злом, тьму почитают светом, и свет – тьмою, горькое почитают сладким, и сладкое – горьким!
ISA|5|21|Горе тем, которые мудры в своих глазах и разумны пред самими собою!
ISA|5|22|Горе тем, которые храбры пить вино и сильны приготовлять крепкий напиток,
ISA|5|23|которые за подарки оправдывают виновного и правых лишают законного!
ISA|5|24|За то, как огонь съедает солому, и пламя истребляет сено, так истлеет корень их, и цвет их разнесется, как прах; потому что они отвергли закон Господа Саваофа и презрели слово Святаго Израилева.
ISA|5|25|За то возгорится гнев Господа на народ Его, и прострет Он руку Свою на него и поразит его, так что содрогнутся горы, и трупы их будут как помет на улицах. И при всем этом гнев Его не отвратится, и рука Его еще будет простерта.
ISA|5|26|И поднимет знамя народам дальним, и даст знак живущему на краю земли, – и вот, он легко и скоро придет;
ISA|5|27|не будет у него ни усталого, ни изнемогающего; ни один не задремлет и не заснет, и не снимется пояс с чресл его, и не разорвется ремень у обуви его;
ISA|5|28|стрелы его заострены, и все луки его натянуты; копыта коней его подобны кремню, и колеса его – как вихрь;
ISA|5|29|рев его – как рев львицы; он рыкает подобно скимнам, и заревет, и схватит добычу и унесет, и никто не отнимет.
ISA|5|30|И заревет на него в тот день как бы рев [разъяренного] моря; и взглянет он на землю, и вот – тьма, горе, и свет померк в облаках.
ISA|6|1|В год смерти царя Озии видел я Господа, сидящего на престоле высоком и превознесенном, и края риз Его наполняли весь храм.
ISA|6|2|Вокруг Него стояли Серафимы; у каждого из них по шести крыл: двумя закрывал каждый лице свое, и двумя закрывал ноги свои, и двумя летал.
ISA|6|3|И взывали они друг ко другу и говорили: Свят, Свят, Свят Господь Саваоф! вся земля полна славы Его!
ISA|6|4|И поколебались верхи врат от гласа восклицающих, и дом наполнился курениями.
ISA|6|5|И сказал я: горе мне! погиб я! ибо я человек с нечистыми устами, и живу среди народа также с нечистыми устами, – и глаза мои видели Царя, Господа Саваофа.
ISA|6|6|Тогда прилетел ко мне один из Серафимов, и в руке у него горящий уголь, который он взял клещами с жертвенника,
ISA|6|7|и коснулся уст моих и сказал: вот, это коснулось уст твоих, и беззаконие твое удалено от тебя, и грех твой очищен.
ISA|6|8|И услышал я голос Господа, говорящего: кого Мне послать? и кто пойдет для Нас? И я сказал: вот я, пошли меня.
ISA|6|9|И сказал Он: пойди и скажи этому народу: слухом услышите – и не уразумеете, и очами смотреть будете – и не увидите.
ISA|6|10|Ибо огрубело сердце народа сего, и ушами с трудом слышат, и очи свои сомкнули, да не узрят очами, и не услышат ушами, и не уразумеют сердцем, и не обратятся, чтобы Я исцелил их.
ISA|6|11|И сказал я: надолго ли, Господи? Он сказал: доколе не опустеют города, и останутся без жителей, и домы без людей, и доколе земля эта совсем не опустеет.
ISA|6|12|И удалит Господь людей, и великое запустение будет на этой земле.
ISA|6|13|И если еще останется десятая часть на ней и возвратится, и она опять будет разорена; [но] как от теревинфа и как от дуба, когда они и срублены, [остается] корень их, так святое семя [будет] корнем ее.
ISA|7|1|И было во дни Ахаза, сына Иоафамова, сына Озии, царя Иудейского, Рецин, царь Сирийский, и Факей, сын Ремалиин, царь Израильский, пошли против Иерусалима, чтобы завоевать его, но не могли завоевать.
ISA|7|2|И было возвещено дому Давидову и сказано: Сирияне расположились в земле Ефремовой; и всколебалось сердце его и сердце народа его, как колеблются от ветра дерева в лесу.
ISA|7|3|И сказал Господь Исаии: выйди ты и сын твой Шеар–ясув навстречу Ахазу, к концу водопровода верхнего пруда, на дорогу к полю белильничьему,
ISA|7|4|и скажи ему: наблюдай и будь спокоен; не страшись и да не унывает сердце твое от двух концов этих дымящихся головней, от разгоревшегося гнева Рецина и Сириян и сына Ремалиина.
ISA|7|5|Сирия, Ефрем и сын Ремалиин умышляют против тебя зло, говоря:
ISA|7|6|пойдем на Иудею и возмутим ее, и овладеем ею и поставим в ней царем сына Тавеилова.
ISA|7|7|Но Господь Бог так говорит: это не состоится и не сбудется;
ISA|7|8|ибо глава Сирии – Дамаск, и глава Дамаска – Рецин; а чрез шестьдесят пять лет Ефрем перестанет быть народом;
ISA|7|9|и глава Ефрема – Самария, и глава Самарии – сын Ремалиин. Если вы не верите, то потому, что вы не удостоверены.
ISA|7|10|И продолжал Господь говорить к Ахазу, и сказал:
ISA|7|11|проси себе знамения у Господа Бога твоего: проси или в глубине, или на высоте.
ISA|7|12|И сказал Ахаз: не буду просить и не буду искушать Господа.
ISA|7|13|Тогда сказал [Исаия]: слушайте же, дом Давидов! разве мало для вас затруднять людей, что вы хотите затруднять и Бога моего?
ISA|7|14|Итак Сам Господь даст вам знамение: се, Дева во чреве приимет и родит Сына, и нарекут имя Ему: Еммануил.
ISA|7|15|Он будет питаться молоком и медом, доколе не будет разуметь отвергать худое и избирать доброе;
ISA|7|16|ибо прежде нежели этот младенец будет разуметь отвергать худое и избирать доброе, земля та, которой ты страшишься, будет оставлена обоими царями ее.
ISA|7|17|Но наведет Господь на тебя и на народ твой и на дом отца твоего дни, какие не приходили со времени отпадения Ефрема от Иуды, наведет царя Ассирийского.
ISA|7|18|И будет в тот день: даст знак Господь мухе, которая при устье реки Египетской, и пчеле, которая в земле Ассирийской, –
ISA|7|19|и прилетят и усядутся все они по долинам опустелым и по расселинам скал, и по всем колючим кустарникам, и по всем деревам.
ISA|7|20|В тот день обреет Господь бритвою, нанятою по ту сторону реки, царем Ассирийским, голову и волоса на ногах, и даже отнимет бороду.
ISA|7|21|И будет в тот день: кто будет содержать корову и двух овец,
ISA|7|22|по изобилию молока, которое они дадут, будет есть масло; маслом и медом будут питаться все, оставшиеся в этой земле.
ISA|7|23|И будет в тот день: на всяком месте, где росла тысяча виноградных лоз на тысячу сребренников, будет терновник и колючий кустарник.
ISA|7|24|Со стрелами и луками будут ходить туда, ибо вся земля будет терновником и колючим кустарником.
ISA|7|25|И ни на одну из гор, которые расчищались бороздниками, не пойдешь, боясь терновника и колючего кустарника: туда будут выгонять волов, и мелкий скот будет топтать их.
ISA|8|1|И сказал мне Господь: возьми себе большой свиток и начертай на нем человеческим письмом: Магер–шелал–хаш–баз.
ISA|8|2|И я взял себе верных свидетелей: Урию священника и Захарию, сына Варахиина, –
ISA|8|3|и приступил я к пророчице, и она зачала и родила сына. И сказал мне Господь: нареки ему имя: Магер–шелал–хаш–баз,
ISA|8|4|ибо прежде нежели дитя будет уметь выговорить: отец мой, мать моя, – богатства Дамаска и добычи Самарийские понесут перед царем Ассирийским.
ISA|8|5|И продолжал Господь говорить ко мне и сказал еще:
ISA|8|6|за то, что этот народ пренебрегает водами Силоама, текущими тихо, и восхищается Рецином и сыном Ремалииным,
ISA|8|7|наведет на него Господь воды реки бурные и большие – царя Ассирийского со всею славою его; и поднимется она во всех протоках своих и выступит из всех берегов своих;
ISA|8|8|и пойдет по Иудее, наводнит ее и высоко поднимется – дойдет до шеи; и распростертие крыльев ее будет во всю широту земли Твоей, Еммануил!
ISA|8|9|Враждуйте, народы, но трепещите, и внимайте, все отдаленные земли! Вооружайтесь, но трепещите; вооружайтесь, но трепещите!
ISA|8|10|Замышляйте замыслы, но они рушатся; говорите слово, но оно не состоится: ибо с нами Бог!
ISA|8|11|Ибо так говорил мне Господь, [держа на мне] крепкую руку и внушая мне не ходить путем сего народа, и сказал:
ISA|8|12|"Не называйте заговором всего того, что народ сей называет заговором; и не бойтесь того, чего он боится, и не страшитесь.
ISA|8|13|Господа Саваофа – Его чтите свято, и Он – страх ваш, и Он – трепет ваш!
ISA|8|14|И будет Он освящением и камнем преткновения, и скалою соблазна для обоих домов Израиля, петлею и сетью для жителей Иерусалима.
ISA|8|15|И многие из них преткнутся и упадут, и разобьются, и запутаются в сети, и будут уловлены.
ISA|8|16|Завяжи свидетельство, и запечатай откровение при учениках Моих".
ISA|8|17|Итак я надеюсь на Господа, сокрывшего лице Свое от дома Иаковлева, и уповаю на Него.
ISA|8|18|Вот я и дети, которых дал мне Господь, как указания и предзнаменования в Израиле от Господа Саваофа, живущего на горе Сионе.
ISA|8|19|И когда скажут вам: обратитесь к вызывателям умерших и к чародеям, к шептунам и чревовещателям, – тогда отвечайте: не должен ли народ обращаться к своему Богу? спрашивают ли мертвых о живых?
ISA|8|20|[Обращайтесь] к закону и откровению. Если они не говорят, как это слово, то нет в них света.
ISA|8|21|И будут они бродить по земле, жестоко угнетенные и голодные; и во время голода будут злиться, хулить царя своего и Бога своего.
ISA|8|22|И взглянут вверх, и посмотрят на землю; и вот – горе и мрак, густая тьма, и будут повержены во тьму. Но не всегда будет мрак там, где теперь он сгустел.
ISA|8|23|Прежнее время умалило землю Завулонову и землю Неффалимову; но последующее возвеличит приморский путь, Заиорданскую страну, Галилею языческую.
ISA|9|1|Народ, ходящий во тьме, увидит свет великий; на живущих в стране тени смертной свет воссияет.
ISA|9|2|Ты умножишь народ, увеличишь радость его. Он будет веселиться пред Тобою, как веселятся во время жатвы, как радуются при разделе добычи.
ISA|9|3|Ибо ярмо, тяготившее его, и жезл, поражавший его, и трость притеснителя его Ты сокрушишь, как в день Мадиама.
ISA|9|4|Ибо всякая обувь воина во время брани и одежда, обагренная кровью, будут отданы на сожжение, в пищу огню.
ISA|9|5|Ибо младенец родился нам – Сын дан нам; владычество на раменах Его, и нарекут имя Ему: Чудный, Советник, Бог крепкий, Отец вечности, Князь мира.
ISA|9|6|Умножению владычества Его и мира нет предела на престоле Давида и в царстве его, чтобы Ему утвердить его и укрепить его судом и правдою отныне и до века. Ревность Господа Саваофа соделает это.
ISA|9|7|Слово посылает Господь на Иакова, и оно нисходит на Израиля,
ISA|9|8|чтобы знал весь народ, Ефрем и жители Самарии, которые с гордостью и надменным сердцем говорят:
ISA|9|9|кирпичи пали – построим из тесаного камня; сикоморы вырублены – заменим их кедрами.
ISA|9|10|И воздвигнет Господь против него врагов Рецина, и неприятелей его вооружит:
ISA|9|11|Сириян с востока, а Филистимлян с запада; и будут они пожирать Израиля полным ртом. При всем этом не отвратится гнев Его, и рука Его еще простерта.
ISA|9|12|Но народ не обращается к Биющему его, и к Господу Саваофу не прибегает.
ISA|9|13|И отсечет Господь у Израиля голову и хвост, пальму и трость, в один день:
ISA|9|14|старец и знатный, – это голова; а пророк–лжеучитель есть хвост.
ISA|9|15|И вожди сего народа введут его в заблуждение, и водимые ими погибнут.
ISA|9|16|Поэтому о юношах его не порадуется Господь, и сирот его и вдов его не помилует: ибо все они – лицемеры и злодеи, и уста всех говорят нечестиво. При всем этом не отвратится гнев Его, и рука Его еще простерта.
ISA|9|17|Ибо беззаконие, как огонь, разгорелось, пожирает терновник и колючий кустарник и пылает в чащах леса, и поднимаются столбы дыма.
ISA|9|18|Ярость Господа Саваофа опалит землю, и народ сделается как бы пищею огня; не пощадит человек брата своего.
ISA|9|19|И будут резать по правую сторону, и останутся голодны; и будут есть по левую, и не будут сыты; каждый будет пожирать плоть мышцы своей:
ISA|9|20|Манассия – Ефрема, и Ефрем – Манассию, оба вместе – Иуду. При всем этом не отвратится гнев Его, и рука Его еще простерта.
ISA|10|1|Горе тем, которые постановляют несправедливые законы и пишут жестокие решения,
ISA|10|2|чтобы устранить бедных от правосудия и похитить права у малосильных из народа Моего, чтобы вдов сделать добычею своею и ограбить сирот.
ISA|10|3|И что вы будете делать в день посещения, когда придет гибель издалека? К кому прибегнете за помощью? И где оставите богатство ваше?
ISA|10|4|Без Меня согнутся между узниками и падут между убитыми. При всем этом не отвратится гнев Его, и рука Его еще простерта.
ISA|10|5|О, Ассур, жезл гнева Моего! и бич в руке его – Мое негодование!
ISA|10|6|Я пошлю его против народа нечестивого и против народа гнева Моего, дам ему повеление ограбить грабежом и добыть добычу и попирать его, как грязь на улицах.
ISA|10|7|Но он не так подумает и не так помыслит сердце его; у него будет на сердце – разорить и истребить немало народов.
ISA|10|8|Ибо он скажет: "не все ли цари князья мои?
ISA|10|9|Халне не то же ли, что Кархемис? Емаф не то же ли, что Арпад? Самария не то же ли, что Дамаск?
ISA|10|10|Так как рука моя овладела царствами идольскими, в которых кумиров более, нежели в Иерусалиме и Самарии, –
ISA|10|11|то не сделаю ли того же с Иерусалимом и изваяниями его, что сделал с Самариею и идолами ее?"
ISA|10|12|И будет, когда Господь совершит все Свое дело на горе Сионе и в Иерусалиме, скажет: посмотрю на успех надменного сердца царя Ассирийского и на тщеславие высоко поднятых глаз его.
ISA|10|13|Он говорит: "силою руки моей и моею мудростью я сделал это, потому что я умен: и переставляю пределы народов, и расхищаю сокровища их, и низвергаю с престолов, как исполин;
ISA|10|14|и рука моя захватила богатство народов, как гнезда; и как забирают оставленные в них яйца, так забрал я всю землю, и никто не пошевелил крылом, и не открыл рта, и не пискнул".
ISA|10|15|Величается ли секира пред тем, кто рубит ею? Пила гордится ли пред тем, кто двигает ее? Как будто жезл восстает против того, кто поднимает его; как будто палка поднимается на того, кто не дерево!
ISA|10|16|За то Господь, Господь Саваоф, пошлет чахлость на тучных его, и между знаменитыми его возжет пламя, как пламя огня.
ISA|10|17|Свет Израиля будет огнем, и Святый его – пламенем, которое сожжет и пожрет терны его и волчцы его в один день;
ISA|10|18|и славный лес его и сад его, от души до тела, истребит; и он будет, как чахлый умирающий.
ISA|10|19|И остаток дерев леса его так будет малочислен, что дитя в состоянии будет сделать опись.
ISA|10|20|И будет в тот день: остаток Израиля и спасшиеся из дома Иакова не будут более полагаться на того, кто поразил их, но возложат упование на Господа, Святаго Израилева, чистосердечно.
ISA|10|21|Остаток обратится, остаток Иакова – к Богу сильному.
ISA|10|22|Ибо, хотя бы народа у тебя, Израиль, [было] столько, сколько песку морского, только остаток его обратится; истребление определено изобилующею правдою;
ISA|10|23|ибо определенное истребление совершит Господь, Господь Саваоф, во всей земле.
ISA|10|24|Посему так говорит Господь, Господь Саваоф: народ Мой, живущий на Сионе! не бойся Ассура. Он поразит тебя жезлом и трость свою поднимет на тебя, как Египет.
ISA|10|25|Еще немного, очень немного, и пройдет Мое негодование, и ярость Моя [обратится] на истребление их.
ISA|10|26|И поднимет Господь Саваоф бич на него, как во время поражения Мадиама у скалы Орива, или как [простер] на море жезл, и поднимет его, как на Египет.
ISA|10|27|И будет в тот день: снимется с рамен твоих бремя его, и ярмо его – с шеи твоей; и распадется ярмо от тука.
ISA|10|28|Он идет на Аиаф, проходит Мигрон, в Михмасе складывает свои запасы.
ISA|10|29|Проходят теснины; в Геве ночлег их; Рама трясется; Гива Саулова разбежалась.
ISA|10|30|Вой голосом твоим, дочь Галима; пусть услышит тебя Лаис, бедный Анафоф!
ISA|10|31|Мадмена разбежалась, жители Гевима спешат уходить.
ISA|10|32|Еще день простоит он в Нове; грозит рукою своею горе Сиону, холму Иерусалимскому.
ISA|10|33|Вот, Господь, Господь Саваоф, страшною силою сорвет ветви дерев, и величающиеся ростом будут срублены, высокие – повержены на землю.
ISA|10|34|И посечет чащу леса железом, и Ливан падет от Всемогущего.
ISA|11|1|И произойдет отрасль от корня Иессеева, и ветвь произрастет от корня его;
ISA|11|2|и почиет на нем Дух Господень, дух премудрости и разума, дух совета и крепости, дух ведения и благочестия;
ISA|11|3|и страхом Господним исполнится, и будет судить не по взгляду очей Своих и не по слуху ушей Своих решать дела.
ISA|11|4|Он будет судить бедных по правде, и дела страдальцев земли решать по истине; и жезлом уст Своих поразит землю, и духом уст Своих убьет нечестивого.
ISA|11|5|И будет препоясанием чресл Его правда, и препоясанием бедр Его – истина.
ISA|11|6|Тогда волк будет жить вместе с ягненком, и барс будет лежать вместе с козленком; и теленок, и молодой лев, и вол будут вместе, и малое дитя будет водить их.
ISA|11|7|И корова будет пастись с медведицею, и детеныши их будут лежать вместе, и лев, как вол, будет есть солому.
ISA|11|8|И младенец будет играть над норою аспида, и дитя протянет руку свою на гнездо змеи.
ISA|11|9|Не будут делать зла и вреда на всей святой горе Моей, ибо земля будет наполнена ведением Господа, как воды наполняют море.
ISA|11|10|И будет в тот день: к корню Иессееву, который станет, как знамя для народов, обратятся язычники, – и покой его будет слава.
ISA|11|11|И будет в тот день: Господь снова прострет руку Свою, чтобы возвратить Себе остаток народа Своего, какой останется у Ассура, и в Египте, и в Патросе, и у Хуса, и у Елама, и в Сеннааре, и в Емафе, и на островах моря.
ISA|11|12|И поднимет знамя язычникам, и соберет изгнанников Израиля, и рассеянных Иудеев созовет от четырех концов земли.
ISA|11|13|И прекратится зависть Ефрема, и враждующие против Иуды будут истреблены. Ефрем не будет завидовать Иуде, и Иуда не будет притеснять Ефрема.
ISA|11|14|И полетят на плеча Филистимлян к западу, ограбят всех детей Востока; на Едома и Моава наложат руку свою, и дети Аммона будут подданными им.
ISA|11|15|И иссушит Господь залив моря Египетского, и прострет руку Свою на реку в сильном ветре Своем, и разобьет ее на семь ручьев, так что в сандалиях могут переходить ее.
ISA|11|16|Тогда для остатка народа Его, который останется у Ассура, будет большая дорога, как это было для Израиля, когда он выходил из земли Египетской.
ISA|12|1|И скажешь в тот день: славлю Тебя, Господи; Ты гневался на меня, но отвратил гнев Твой и утешил меня.
ISA|12|2|Вот, Бог – спасение мое: уповаю на Него и не боюсь; ибо Господь – сила моя, и пение мое – Господь; и Он был мне во спасение.
ISA|12|3|И в радости будете почерпать воду из источников спасения,
ISA|12|4|и скажете в тот день: славьте Господа, призывайте имя Его; возвещайте в народах дела Его; напоминайте, что велико имя Его;
ISA|12|5|пойте Господу, ибо Он соделал великое, – да знают это по всей земле.
ISA|12|6|Веселись и радуйся, жительница Сиона, ибо велик посреди тебя Святый Израилев.
ISA|13|1|Пророчество о Вавилоне, которое изрек Исаия, сын Амосов.
ISA|13|2|Поднимите знамя на открытой горе, возвысьте голос; махните им рукою, чтобы шли в ворота властелинов.
ISA|13|3|Я дал повеление избранным Моим и призвал для [совершения] гнева Моего сильных Моих, торжествующих в величии Моем.
ISA|13|4|Большой шум на горах, как бы от многолюдного народа, мятежный шум царств и народов, собравшихся вместе: Господь Саваоф обозревает боевое войско.
ISA|13|5|Идут из отдаленной страны, от края неба, Господь и орудия гнева Его, чтобы сокрушить всю землю.
ISA|13|6|Рыдайте, ибо день Господа близок, идет как разрушительная сила от Всемогущего.
ISA|13|7|От того руки у всех опустились, и сердце у каждого человека растаяло.
ISA|13|8|Ужаснулись, судороги и боли схватили их; мучатся, как рождающая, с изумлением смотрят друг на друга, лица у них разгорелись.
ISA|13|9|Вот, приходит день Господа лютый, с гневом и пылающею яростью, чтобы сделать землю пустынею и истребить с нее грешников ее.
ISA|13|10|Звезды небесные и светила не дают от себя света; солнце меркнет при восходе своем, и луна не сияет светом своим.
ISA|13|11|Я накажу мир за зло, и нечестивых – за беззакония их, и положу конец высокоумию гордых, и уничижу надменность притеснителей;
ISA|13|12|сделаю то, что люди будут дороже чистого золота, и мужи – дороже золота Офирского.
ISA|13|13|Для сего потрясу небо, и земля сдвинется с места своего от ярости Господа Саваофа, в день пылающего гнева Его.
ISA|13|14|Тогда каждый, как преследуемая серна и как покинутые овцы, обратится к народу своему, и каждый побежит в свою землю.
ISA|13|15|Но кто попадется, будет пронзен, и кого схватят, тот падет от меча.
ISA|13|16|И младенцы их будут разбиты пред глазами их; домы их будут разграблены и жены их обесчещены.
ISA|13|17|Вот, Я подниму против них Мидян, которые не ценят серебра и не пристрастны к золоту.
ISA|13|18|Луки их сразят юношей и не пощадят плода чрева: глаз их не сжалится над детьми.
ISA|13|19|И Вавилон, краса царств, гордость Халдеев, будет ниспровержен Богом, как Содом и Гоморра,
ISA|13|20|не заселится никогда, и в роды родов не будет жителей в нем; не раскинет Аравитянин шатра своего, и пастухи со стадами не будут отдыхать там.
ISA|13|21|Но будут обитать в нем звери пустыни, и домы наполнятся филинами; и страусы поселятся, и косматые будут скакать там.
ISA|13|22|Шакалы будут выть в чертогах их, и гиены – в увеселительных домах.
ISA|14|1|Близко время его, и не замедлят дни его, ибо помилует Господь Иакова и снова возлюбит Израиля; и поселит их на земле их, и присоединятся к ним иноземцы и прилепятся к дому Иакова.
ISA|14|2|И возьмут их народы, и приведут на место их, и дом Израиля усвоит их себе на земле Господней рабами и рабынями, и возьмет в плен пленивших его, и будет господствовать над угнетателями своими.
ISA|14|3|И будет в тот день: когда Господь устроит тебя от скорби твоей и от страха и от тяжкого рабства, которому ты порабощен был,
ISA|14|4|ты произнесешь победную песнь на царя Вавилонского и скажешь: как не стало мучителя, пресеклось грабительство!
ISA|14|5|Сокрушил Господь жезл нечестивых, скипетр владык,
ISA|14|6|поражавший народы в ярости ударами неотвратимыми, во гневе господствовавший над племенами с неудержимым преследованием.
ISA|14|7|Вся земля отдыхает, покоится, восклицает от радости;
ISA|14|8|и кипарисы радуются о тебе, и кедры ливанские, [говоря]: "с тех пор, как ты заснул, никто не приходит рубить нас".
ISA|14|9|Ад преисподний пришел в движение ради тебя, чтобы встретить тебя при входе твоем; пробудил для тебя Рефаимов, всех вождей земли; поднял всех царей языческих с престолов их.
ISA|14|10|Все они будут говорить тебе: и ты сделался бессильным, как мы! и ты стал подобен нам!
ISA|14|11|В преисподнюю низвержена гордыня твоя со всем шумом твоим; под тобою подстилается червь, и черви – покров твой.
ISA|14|12|Как упал ты с неба, денница, сын зари! разбился о землю, попиравший народы.
ISA|14|13|А говорил в сердце своем: "взойду на небо, выше звезд Божиих вознесу престол мой и сяду на горе в сонме богов, на краю севера;
ISA|14|14|взойду на высоты облачные, буду подобен Всевышнему".
ISA|14|15|Но ты низвержен в ад, в глубины преисподней.
ISA|14|16|Видящие тебя всматриваются в тебя, размышляют о тебе: "тот ли это человек, который колебал землю, потрясал царства,
ISA|14|17|вселенную сделал пустынею и разрушал города ее, пленников своих не отпускал домой?"
ISA|14|18|Все цари народов, все лежат с честью, каждый в своей усыпальнице;
ISA|14|19|а ты повержен вне гробницы своей, как презренная ветвь, как одежда убитых, сраженных мечом, которых опускают в каменные рвы, – ты, как попираемый труп,
ISA|14|20|не соединишься с ними в могиле; ибо ты разорил землю твою, убил народ твой: во веки не помянется племя злодеев.
ISA|14|21|Готовьте заклание сыновьям его за беззаконие отца их, чтобы не восстали и не завладели землею и не наполнили вселенной неприятелями.
ISA|14|22|И восстану на них, говорит Господь Саваоф, и истреблю имя Вавилона и весь остаток, и сына и внука, говорит Господь.
ISA|14|23|И сделаю его владением ежей и болотом, и вымету его метлою истребительною, говорит Господь Саваоф.
ISA|14|24|С клятвою говорит Господь Саваоф: как Я помыслил, так и будет; как Я определил, так и состоится,
ISA|14|25|чтобы сокрушить Ассура в земле Моей и растоптать его на горах Моих; и спадет с них ярмо его, и снимется бремя его с рамен их.
ISA|14|26|Таково определение, постановленное о всей земле, и вот рука, простертая на все народы,
ISA|14|27|ибо Господь Саваоф определил, и кто может отменить это? рука Его простерта, – и кто отвратит ее?
ISA|14|28|В год смерти царя Ахаза было такое пророческое слово:
ISA|14|29|не радуйся, земля Филистимская, что сокрушен жезл, который поражал тебя, ибо из корня змеиного выйдет аспид, и плодом его будет летучий дракон.
ISA|14|30|Тогда беднейшие будут накормлены, и нищие будут покоиться в безопасности; а твой корень уморю голодом, и он убьет остаток твой.
ISA|14|31|Рыдайте, ворота! вой голосом, город! Распадешься ты, вся земля Филистимская, ибо от севера дым идет, и нет отсталого в полчищах их.
ISA|14|32|Что же скажут вестники народа? – То, что Господь утвердил Сион, и в нем найдут убежище бедные из народа Его.
ISA|15|1|Пророчество о Моаве. – Так! ночью будет разорен Ар–Моав и уничтожен; так! ночью будет разорен Кир–Моав и уничтожен!
ISA|15|2|Он восходит к Баиту и Дивону, восходит на высоты, чтобы плакать; Моав рыдает над Нево и Медевою; у всех их острижены головы, у всех обриты бороды.
ISA|15|3|На улицах его препоясываются вретищем; на кровлях его и площадях его все рыдает, утопает в слезах.
ISA|15|4|И вопит Есевон и Елеала; голос их слышится до самой Иаацы; за ними и воины Моава рыдают; душа его возмущена в нем.
ISA|15|5|Рыдает сердце мое о Моаве; бегут из него к Сигору, до третьей Эглы; восходят на Лухит с плачем; по дороге Хоронаимской поднимают страшный крик;
ISA|15|6|потому что воды Нимрима иссякли, луга засохли, трава выгорела, не стало зелени.
ISA|15|7|Поэтому они остатки стяжания и, что сбережено ими, переносят за реку Аравийскую.
ISA|15|8|Ибо вопль по всем пределам Моава, до Эглаима плач его и до Беэр–Елима плач его;
ISA|15|9|потому что воды Димона наполнились кровью, и Я наведу на Димон еще новое – львов на убежавших из Моава и на оставшихся в стране.
ISA|16|1|Посылайте агнцев владетелю земли из Селы в пустыне на гору дочери Сиона;
ISA|16|2|ибо блуждающей птице, выброшенной из гнезда, будут подобны дочери Моава у бродов Арнонских.
ISA|16|3|"Составь совет, постанови решение; осени нас среди полудня, как ночью, тенью твоею, укрой изгнанных, не выдай скитающихся.
ISA|16|4|Пусть поживут у тебя мои изгнанные Моавитяне; будь им покровом от грабителя: ибо притеснителя не станет, грабеж прекратится, попирающие исчезнут с земли.
ISA|16|5|И утвердится престол милостью, и воссядет на нем в истине, в шатре Давидовом, судия, ищущий правды и стремящийся к правосудию".
ISA|16|6|"Слыхали мы о гордости Моава, гордости чрезмерной, о надменности его и высокомерии и неистовстве его: неискренна речь его".
ISA|16|7|Поэтому возрыдает Моав о Моаве, – все будут рыдать; стенайте о твердынях Кирхарешета: они совершенно разрушены.
ISA|16|8|Поля Есевонские оскудели, также и виноградник Севамский; властители народов истребили лучшие лозы его, которые достигали до Иазера, расстилались по пустыне; побеги их расширялись, переходили за море.
ISA|16|9|Посему [и] я буду плакать о лозе Севамской плачем Иазера, буду обливать тебя слезами моими, Есевон и Елеала; ибо во время собирания винограда твоего и во время жатвы твоей нет более шумной радости.
ISA|16|10|Исчезло с плодоносной земли веселье и ликование, и в виноградниках не поют, не ликуют; виноградарь не топчет винограда в точилах: Я прекратил ликование.
ISA|16|11|От того внутренность моя стонет о Моаве, как гусли, и сердце мое – о Кирхарешете.
ISA|16|12|Хотя и явится Моав, и будет до утомления [подвизаться] на высотах, и придет к святилищу своему помолиться, но ничто не поможет.
ISA|16|13|Вот слово, которое изрек Господь о Моаве издавна.
ISA|16|14|Ныне же так говорит Господь: чрез три года, считая годами наемничьими, величие Моава будет унижено со всем великим многолюдством, и остаток [будет] очень малый и незначительный.
ISA|17|1|Пророчество о Дамаске. – Вот, Дамаск исключается из [числа] городов и будет грудою развалин.
ISA|17|2|Города Ароерские будут покинуты, – останутся для стад, которые будут отдыхать там, и некому будет пугать их.
ISA|17|3|Не станет твердыни Ефремовой и царства Дамасского с остальною Сириею; с ними будет то же, что со славою сынов Израиля, говорит Господь Саваоф.
ISA|17|4|И будет в тот день: умалится слава Иакова, и тучное тело его сделается тощим.
ISA|17|5|То же будет, что по собрании хлеба жнецом, когда рука его пожнет колосья, и когда соберут колосья в долине Рефаимской.
ISA|17|6|И останутся у него, как бывает при обивании маслин, две–три ягоды на самой вершине, или четыре–пять на плодоносных ветвях, говорит Господь, Бог Израилев.
ISA|17|7|В тот день обратит человек взор свой к Творцу своему, и глаза его будут устремлены к Святому Израилеву;
ISA|17|8|и не взглянет на жертвенники, на дело рук своих, и не посмотрит на то, что сделали персты его, на кумиры Астарты и Ваала.
ISA|17|9|В тот день укрепленные города его будут, как развалины в лесах и на вершинах гор, оставленные пред сынами Израиля, – и будет пусто.
ISA|17|10|Ибо ты забыл Бога спасения твоего, и не воспоминал о скале прибежища твоего; от того развел увеселительные сады и насадил черенки от чужой лозы.
ISA|17|11|В день насаждения твоего ты заботился, чтобы оно росло и чтобы посеянное тобою рано расцвело; но в день собирания не куча жатвы будет, но скорбь жестокая.
ISA|17|12|Увы! шум народов многих! шумят они, как шумит море. Рев племен! они ревут, как ревут сильные воды.
ISA|17|13|Ревут народы, как ревут сильные воды; но Он погрозил им и они далеко побежали, и были гонимы, как прах по горам от ветра и как пыль от вихря.
ISA|17|14|Вечер – и вот ужас! и прежде утра уже нет его. Такова участь грабителей наших, жребий разорителей наших.
ISA|18|1|Горе земле, осеняющей крыльями по ту сторону рек Ефиопских,
ISA|18|2|посылающей послов по морю, и в папировых суднах по водам! Идите, быстрые послы, к народу крепкому и бодрому, к народу страшному от начала и доныне, к народу рослому и [все] попирающему, которого землю разрезывают реки.
ISA|18|3|Все вы, населяющие вселенную и живущие на земле! смотрите, когда знамя поднимется на горах, и, когда загремит труба, слушайте!
ISA|18|4|Ибо так Господь сказал мне: Я спокойно смотрю из жилища Моего, как светлая теплота после дождя, как облако росы во время жатвенного зноя.
ISA|18|5|Ибо прежде собирания винограда, когда он отцветет, и грозд начнет созревать, Он отрежет ножом ветви и отнимет, и отрубит отрасли.
ISA|18|6|И оставят все хищным птицам на горах и зверям полевым; и птицы будут проводить там лето, а все звери полевые будут зимовать там.
ISA|18|7|В то время будет принесен дар Господу Саваофу от народа крепкого и бодрого, от народа страшного от начала и доныне, от народа рослого и [все] попирающего, которого землю разрезывают реки, – к месту имени Господа Саваофа, на гору Сион.
ISA|19|1|Пророчество о Египте. – Вот, Господь восседит на облаке легком и грядет в Египет. И потрясутся от лица Его идолы Египетские, и сердце Египта растает в нем.
ISA|19|2|Я вооружу Египтян против Египтян; и будут сражаться брат против брата и друг против друга, город с городом, царство с царством.
ISA|19|3|И дух Египта изнеможет в нем, и разрушу совет его, и прибегнут они к идолам и к чародеям, и к вызывающим мертвых и к гадателям.
ISA|19|4|И предам Египтян в руки властителя жестокого, и свирепый царь будет господствовать над ними, говорит Господь, Господь Саваоф.
ISA|19|5|И истощатся воды в море и река иссякнет и высохнет;
ISA|19|6|и оскудеют реки, и каналы Египетские обмелеют и высохнут; камыш и тростник завянут.
ISA|19|7|Поля при реке, по берегам реки, и все, посеянное при реке, засохнет, развеется и исчезнет.
ISA|19|8|И восплачут рыбаки, и возрыдают все, бросающие уду в реку, и ставящие сети в воде впадут в уныние;
ISA|19|9|и будут в смущении обрабатывающие лен и ткачи белых полотен;
ISA|19|10|и будут сокрушены сети, и все, которые содержат садки для живой рыбы, упадут в духе.
ISA|19|11|Так! обезумели князья Цоанские; совет мудрых советников фараоновых стал бессмысленным. Как скажете вы фараону: "я сын мудрецов, сын царей древних?"
ISA|19|12|Где они? где твои мудрецы? пусть они теперь скажут тебе; пусть узнают, что Господь Саваоф определил о Египте.
ISA|19|13|Обезумели князья Цоанские; обманулись князья Мемфисские, и совратил Египет с пути главы племен его.
ISA|19|14|Господь послал в него дух опьянения; и они ввели Египет в заблуждение во всех делах его, подобно тому, как пьяный бродит по блевотине своей.
ISA|19|15|И не будет в Египте такого дела, которое совершить умели бы голова и хвост, пальма и трость.
ISA|19|16|В тот день Египтяне будут подобны женщинам, и вострепещут и убоятся движения руки Господа Саваофа, которую Он поднимет на них.
ISA|19|17|Земля Иудина сделается ужасом для Египта; кто вспомнит о ней, тот затрепещет от определения Господа Саваофа, которое Он постановил о нем.
ISA|19|18|В тот день пять городов в земле Египетской будут говорить языком Ханаанским и клясться Господом Саваофом; один назовется городом солнца.
ISA|19|19|В тот день жертвенник Господу будет посреди земли Египетской, и памятник Господу – у пределов ее.
ISA|19|20|И будет он знамением и свидетельством о Господе Саваофе в земле Египетской, потому что они воззовут к Господу по причине притеснителей, и Он пошлет им спасителя и заступника, и избавит их.
ISA|19|21|И Господь явит Себя в Египте; и Египтяне в тот день познают Господа и принесут жертвы и дары, и дадут обеты Господу, и исполнят.
ISA|19|22|И поразит Господь Египет; поразит и исцелит; они обратятся к Господу, и Он услышит их, и исцелит их.
ISA|19|23|В тот день из Египта в Ассирию будет большая дорога, и будет приходить Ассур в Египет, и Египтяне – в Ассирию; и Египтяне вместе с Ассириянами будут служить Господу.
ISA|19|24|В тот день Израиль будет третьим с Египтом и Ассириею; благословение будет посреди земли,
ISA|19|25|которую благословит Господь Саваоф, говоря: благословен народ Мой – Египтяне, и дело рук Моих – Ассирияне, и наследие Мое – Израиль.
ISA|20|1|В год, когда Тартан пришел к Азоту, быв послан от Саргона, царя Ассирийского, и воевал против Азота, и взял его,
ISA|20|2|в то самое время Господь сказал Исаии, сыну Амосову, так: пойди и сними вретище с чресл твоих и сбрось сандалии твои с ног твоих. Он так и сделал: ходил нагой и босой.
ISA|20|3|И сказал Господь: как раб Мой Исаия ходил нагой и босой три года, в указание и предзнаменование о Египте и Ефиопии,
ISA|20|4|так поведет царь Ассирийский пленников из Египта и переселенцев из Ефиопии, молодых и старых, нагими и босыми и с обнаженными чреслами, в посрамление Египту.
ISA|20|5|Тогда ужаснутся и устыдятся из–за Ефиопии, надежды своей, и из–за Египта, которым хвалились.
ISA|20|6|И скажут в тот день жители этой страны: вот каковы те, на которых мы надеялись и к которым прибегали за помощью, чтобы спастись от царя Ассирийского! и как спаслись бы мы?
ISA|21|1|Пророчество о пустыне приморской. – Как бури на юге носятся, идет он от пустыни, из земли страшной.
ISA|21|2|Грозное видение показано мне: грабитель грабит, опустошитель опустошает; восходи, Елам, осаждай, Мид! всем стенаниям я положу конец.
ISA|21|3|От этого чресла мои трясутся; муки схватили меня, как муки рождающей. Я взволнован от того, что слышу; я смущен от того, что вижу.
ISA|21|4|Сердце мое трепещет; дрожь бьет меня; отрадная ночь моя превратилась в ужас для меня.
ISA|21|5|Приготовляют стол, расстилают покрывала, – едят, пьют. "Вставайте, князья, мажьте щиты!"
ISA|21|6|Ибо так сказал мне Господь: пойди, поставь сторожа; пусть он сказывает, что увидит.
ISA|21|7|И увидел он едущих попарно всадников на конях, всадников на ослах, всадников на верблюдах; и вслушивался он прилежно, с большим вниманием, –
ISA|21|8|и закричал, [как] лев: господин мой! на страже стоял я весь день, и на месте моем оставался целые ночи:
ISA|21|9|и вот, едут люди, всадники на конях попарно. Потом он возгласил и сказал: пал, пал Вавилон, и все идолы богов его лежат на земле разбитые.
ISA|21|10|О, измолоченный мой и сын гумна моего! Что слышал я от Господа Саваофа, Бога Израилева, то и возвестил вам.
ISA|21|11|Пророчество о Думе. – Кричат мне с Сеира: сторож! сколько ночи? сторож! сколько ночи?
ISA|21|12|Сторож отвечает: приближается утро, но еще ночь. Если вы настоятельно спрашиваете, то обратитесь и приходите.
ISA|21|13|Пророчество об Аравии. – В лесу Аравийском ночуйте, караваны Деданские!
ISA|21|14|Живущие в земле Фемайской! несите воды навстречу жаждущим; с хлебом встречайте бегущих,
ISA|21|15|ибо они от мечей бегут, от меча обнаженного и от лука натянутого, и от лютости войны.
ISA|21|16|Ибо так сказал мне Господь: еще год, равный году наемничьему, и вся слава Кидарова исчезнет,
ISA|21|17|и луков у храбрых сынов Кидара останется немного: так сказал Господь, Бог Израилев.
ISA|22|1|Пророчество о долине видения. – Что с тобою, что ты весь взошел на кровли?
ISA|22|2|Город шумный, волнующийся, город ликующий! Пораженные твои не мечом убиты и не в битве умерли;
ISA|22|3|все вожди твои бежали вместе, но были связаны стрелками; все найденные у тебя связаны вместе, как ни далеко бежали.
ISA|22|4|Потому говорю: оставьте меня, я буду плакать горько; не усиливайтесь утешать меня в разорении дочери народа моего.
ISA|22|5|Ибо день смятения и попрания и замешательства в долине видения от Господа, Бога Саваофа. Ломают стену, и крик восходит на горы.
ISA|22|6|И Елам несет колчан; люди на колесницах [и] всадники, и Кир обнажает щит.
ISA|22|7|И вот, лучшие долины твои полны колесницами, и всадники выстроились против ворот,
ISA|22|8|и снимают покров с Иудеи; и ты в тот день обращаешь взор на запас оружия в доме кедровом.
ISA|22|9|Но вы видите, что много проломов в стене города Давидова, и собираете воды в нижнем пруде;
ISA|22|10|и отмечаете домы в Иерусалиме, и разрушаете домы, чтобы укрепить стену;
ISA|22|11|и устрояете между двумя стенами хранилище для вод старого пруда. А на Того, Кто это делает, не взираете, и не смотрите на Того, Кто издавна определил это.
ISA|22|12|И Господь, Господь Саваоф, призывает вас в этот день плакать и сетовать, и остричь волоса и препоясаться вретищем.
ISA|22|13|Но вот, веселье и радость! Убивают волов, и режут овец; едят мясо, и пьют вино: "будем есть и пить, ибо завтра умрем!"
ISA|22|14|И открыл мне в уши Господь Саваоф: не будет прощено вам это нечестие, доколе не умрете, сказал Господь, Господь Саваоф.
ISA|22|15|Так сказал Господь, Господь Саваоф: ступай, пойди к этому царедворцу, к Севне, начальнику дворца [и скажи ему]:
ISA|22|16|что у тебя здесь, и кто здесь у тебя, что ты здесь высекаешь себе гробницу? – Он высекает себе гробницу на возвышенности, вырубает в скале жилище себе.
ISA|22|17|Вот, Господь перебросит тебя, как бросает сильный человек, и сожмет тебя в ком;
ISA|22|18|свернув тебя в сверток, бросит тебя, как меч, в землю обширную; там ты умрешь, и там великолепные колесницы твои будут поношением для дома господина твоего.
ISA|22|19|И столкну тебя с места твоего, и свергну тебя со степени твоей.
ISA|22|20|И будет в тот день, призову раба Моего Елиакима, сына Хелкиина,
ISA|22|21|и одену его в одежду твою, и поясом твоим опояшу его, и власть твою передам в руки его; и будет он отцом для жителей Иерусалима и для дома Иудина.
ISA|22|22|И ключ дома Давидова возложу на рамена его; отворит он, и никто не запрет; запрет он, и никто не отворит.
ISA|22|23|И укреплю его как гвоздь в твердом месте; и будет он как седалище славы для дома отца своего.
ISA|22|24|И будет висеть на нем вся слава дома отца его, детей и внуков, всей домашней утвари до последних музыкальных орудий.
ISA|22|25|В тот день, говорит Господь Саваоф, пошатнется гвоздь, укрепленный в твердом месте, и будет выбит, и упадет, и распадется вся тяжесть, которая на нем: ибо Господь говорит.
ISA|23|1|Пророчество о Тире. – Рыдайте, корабли Фарсиса, ибо он разрушен; нет домов, и некому входить в домы. Так им возвещено из земли Киттийской.
ISA|23|2|Умолкните, обитатели острова, который наполняли купцы Сидонские, плавающие по морю.
ISA|23|3|По великим водам привозились в него семена Сихора, жатва [большой] реки, и был он торжищем народов.
ISA|23|4|Устыдись, Сидон; ибо [вот что] говорит море, крепость морская: "как бы ни мучилась я родами и ни рождала, и ни воспитывала юношей, ни возращала девиц".
ISA|23|5|Когда весть дойдет до Египтян, содрогнутся они, услышав о Тире.
ISA|23|6|Переселяйтесь в Фарсис, рыдайте, обитатели острова!
ISA|23|7|Это ли ваш ликующий город, которого начало от дней древних? Ноги его несут его скитаться в стране далекой.
ISA|23|8|Кто определил это Тиру, который раздавал венцы, которого купцы [были] князья, торговцы – знаменитости земли?
ISA|23|9|Господь Саваоф определил это, чтобы посрамить надменность всякой славы, чтобы унизить все знаменитости земли.
ISA|23|10|Ходи по земле твоей, дочь Фарсиса, как река: нет более препоны.
ISA|23|11|Он простер руку Свою на море, потряс царства; Господь дал повеление о Ханаане разрушить крепости его
ISA|23|12|и сказал: ты не будешь более ликовать, посрамленная девица, дочь Сидона! Вставай, иди в Киттим, [но] и там не будет тебе покоя.
ISA|23|13|Вот земля Халдеев. Этого народа прежде не было; Ассур положил ему начало из обитателей пустынь. Они ставят башни свои, разрушают чертоги его, превращают его в развалины.
ISA|23|14|Рыдайте, корабли Фарсисские! Ибо твердыня ваша разорена.
ISA|23|15|И будет в тот день, забудут Тир на семьдесят лет, в мере дней одного царя. По окончании же семидесяти лет с Тиром будет то же, что поют о блуднице:
ISA|23|16|"возьми цитру, ходи по городу, забытая блудница! Играй складно, пой много песен, чтобы вспомнили о тебе".
ISA|23|17|И будет, по истечении семидесяти лет, Господь посетит Тир; и он снова начнет получать прибыль свою и будет блудодействовать со всеми царствами земными по всей вселенной.
ISA|23|18|Но торговля его и прибыль его будут посвящаемы Господу; не будут заперты и уложены в кладовые, ибо к живущим пред лицем Господа будет переходить прибыль от торговли его, чтобы они ели до сытости и имели одежду прочную.
ISA|24|1|Вот, Господь опустошает землю и делает ее бесплодною; изменяет вид ее и рассевает живущих на ней.
ISA|24|2|И что будет с народом, то и со священником; что со слугою, то и с господином его; что со служанкою, то и с госпожею ее; что с покупающим, то и с продающим; что с заемщиком, то и с заимодавцем; что с ростовщиком, то и с дающим в рост.
ISA|24|3|Земля опустошена вконец и совершенно разграблена, ибо Господь изрек слово сие.
ISA|24|4|Сетует, уныла земля; поникла, уныла вселенная; поникли возвышавшиеся над народом земли.
ISA|24|5|И земля осквернена под живущими на ней, ибо они преступили законы, изменили устав, нарушили вечный завет.
ISA|24|6|За то проклятие поедает землю, и несут наказание живущие на ней; за то сожжены обитатели земли, и немного осталось людей.
ISA|24|7|Плачет сок грозда; болит виноградная лоза; воздыхают все веселившиеся сердцем.
ISA|24|8|Прекратилось веселье с тимпанами; умолк шум веселящихся; затихли звуки гуслей;
ISA|24|9|уже не пьют вина с песнями; горька сикера для пьющих ее.
ISA|24|10|Разрушен опустевший город, все домы заперты, нельзя войти.
ISA|24|11|Плачут о вине на улицах; помрачилась всякая радость; изгнано всякое веселие земли.
ISA|24|12|В городе осталось запустение, и ворота развалились.
ISA|24|13|А посреди земли, между народами, будет то же, что бывает при обивании маслин, при обирании [винограда], когда кончена уборка.
ISA|24|14|Они возвысят голос свой, восторжествуют в величии Господа, громко будут восклицать с моря.
ISA|24|15|Итак славьте Господа на востоке, на островах морских – имя Господа, Бога Израилева.
ISA|24|16|От края земли мы слышим песнь: "Слава Праведному!" И сказал я: беда мне, беда мне! увы мне! злодеи злодействуют, и злодействуют злодеи злодейски.
ISA|24|17|Ужас и яма и петля для тебя, житель земли!
ISA|24|18|Тогда побежавший от крика ужаса упадет в яму; и кто выйдет из ямы, попадет в петлю; ибо окна с [небесной] высоты растворятся, и основания земли потрясутся.
ISA|24|19|Земля сокрушается, земля распадается, земля сильно потрясена;
ISA|24|20|шатается земля, как пьяный, и качается, как колыбель, и беззаконие ее тяготеет на ней; она упадет, и уже не встанет.
ISA|24|21|И будет в тот день: посетит Господь воинство выспреннее на высоте и царей земных на земле.
ISA|24|22|И будут собраны вместе, как узники, в ров, и будут заключены в темницу, и после многих дней будут наказаны.
ISA|24|23|И покраснеет луна, и устыдится солнце, когда Господь Саваоф воцарится на горе Сионе и в Иерусалиме, и пред старейшинами его [будет] слава.
ISA|25|1|Господи! Ты Бог мой; превознесу Тебя, восхвалю имя Твое, ибо Ты совершил дивное; предопределения древние истинны, аминь.
ISA|25|2|Ты превратил город в груду камней, твердую крепость в развалины; чертогов иноплеменников уже не стало в городе; вовек не будет он восстановлен.
ISA|25|3|Посему будут прославлять Тебя народы сильные; города страшных племен будут бояться Тебя,
ISA|25|4|ибо Ты был убежищем бедного, убежищем нищего в тесное для него время, защитою от бури, тенью от зноя; ибо гневное дыхание тиранов было подобно буре против стены.
ISA|25|5|Как зной в месте безводном, Ты укротил буйство врагов; [как] зной тенью облака, подавлено ликование притеснителей.
ISA|25|6|И сделает Господь Саваоф на горе сей для всех народов трапезу из тучных яств, трапезу из чистых вин, из тука костей и самых чистых вин;
ISA|25|7|и уничтожит на горе сей покрывало, покрывающее все народы, покрывало, лежащее на всех племенах.
ISA|25|8|Поглощена будет смерть навеки, и отрет Господь Бог слезы со всех лиц, и снимет поношение с народа Своего по всей земле; ибо так говорит Господь.
ISA|25|9|И скажут в тот день: вот Он, Бог наш! на Него мы уповали, и Он спас нас! Сей есть Господь; на Него уповали мы; возрадуемся и возвеселимся во спасении Его!
ISA|25|10|Ибо рука Господа почиет на горе сей, и Моав будет попран на месте своем, как попирается солома в навозе.
ISA|25|11|И хотя он распрострет посреди его руки свои, как плавающий распростирает их для плавания; [но Бог] унизит гордость его вместе с лукавством рук его.
ISA|25|12|И твердыню высоких стен твоих обрушит, низвергнет, повергнет на землю, в прах.
ISA|26|1|В тот день будет воспета песнь сия в земле Иудиной: город крепкий у нас; спасение дал Он вместо стены и вала.
ISA|26|2|Отворите ворота; да войдет народ праведный, хранящий истину.
ISA|26|3|Твердого духом Ты хранишь в совершенном мире, ибо на Тебя уповает он.
ISA|26|4|Уповайте на Господа вовеки, ибо Господь Бог есть твердыня вечная:
ISA|26|5|Он ниспроверг живших на высоте, высоко стоявший город; поверг его, поверг на землю, бросил его в прах.
ISA|26|6|Нога попирает его, ноги бедного, стопы нищих.
ISA|26|7|Путь праведника прям; Ты уравниваешь стезю праведника.
ISA|26|8|И на пути судов Твоих, Господи, мы уповали на Тебя; к имени Твоему и к воспоминанию о Тебе стремилась душа наша.
ISA|26|9|Душею моею я стремился к Тебе ночью, и духом моим я буду искать Тебя во внутренности моей с раннего утра: ибо когда суды Твои [совершаются] на земле, тогда живущие в мире научаются правде.
ISA|26|10|Если нечестивый будет помилован, то не научится он правде, – будет злодействовать в земле правых и не будет взирать на величие Господа.
ISA|26|11|Господи! рука Твоя была высоко поднята, но они не видали ее; увидят и устыдятся ненавидящие народ Твой; огонь пожрет врагов Твоих.
ISA|26|12|Господи! Ты даруешь нам мир; ибо и все дела наши Ты устрояешь для нас.
ISA|26|13|Господи Боже наш! другие владыки кроме Тебя господствовали над нами; но чрез Тебя только мы славим имя Твое.
ISA|26|14|Мертвые не оживут; рефаимы не встанут, потому что Ты посетил и истребил их, и уничтожил всякую память о них.
ISA|26|15|Ты умножил народ, Господи, умножил народ, – прославил Себя, распространил все пределы земли.
ISA|26|16|Господи! в бедствии он искал Тебя; изливал тихие моления, когда наказание Твое постигало его.
ISA|26|17|Как беременная женщина, при наступлении родов, мучится, вопит от болей своих, так были мы пред Тобою, Господи.
ISA|26|18|Были беременны, мучились, – и рождали как бы ветер; спасения не доставили земле, и прочие жители вселенной не пали.
ISA|26|19|Оживут мертвецы Твои, восстанут мертвые тела! Воспряните и торжествуйте, поверженные в прахе: ибо роса Твоя – роса растений, и земля извергнет мертвецов.
ISA|26|20|Пойди, народ мой, войди в покои твои и запри за собой двери твои, укройся на мгновение, доколе не пройдет гнев;
ISA|26|21|ибо вот, Господь выходит из жилища Своего наказать обитателей земли за их беззаконие, и земля откроет поглощенную ею кровь и уже не скроет убитых своих.
ISA|27|1|В тот день поразит Господь мечом Своим тяжелым, и большим и крепким, левиафана, змея прямо бегущего, и левиафана, змея изгибающегося, и убьет чудовище морское.
ISA|27|2|В тот день воспойте о нем – о возлюбленном винограднике:
ISA|27|3|Я, Господь, хранитель его, в каждое мгновение напояю его; ночью и днем стерегу его, чтобы кто не ворвался в него.
ISA|27|4|Гнева нет во Мне. Но если бы кто противопоставил Мне [в нем] волчцы и терны, Я войною пойду против него, выжгу его совсем.
ISA|27|5|Разве прибегнет к защите Моей и заключит мир со Мною? тогда пусть заключит мир со Мною.
ISA|27|6|В грядущие [дни] укоренится Иаков, даст отпрыск и расцветет Израиль; и наполнится плодами вселенная.
ISA|27|7|Так ли Он поражал его, как поражал поражавших его? Так ли убивал его, как убиты убивавшие его?
ISA|27|8|Мерою Ты наказывал его, когда отвергал его; выбросил его сильным дуновением Своим как бы в день восточного ветра.
ISA|27|9|И чрез это загладится беззаконие Иакова; и плодом сего будет снятие греха с него, когда все камни жертвенников он обратит в куски извести, и не будут уже стоять дубравы и истуканы солнца.
ISA|27|10|Ибо укрепленный город опустеет, жилища [будут] покинуты и заброшены, как пустыня. Там будет пастись теленок, и там он будет покоиться и объедать ветви его.
ISA|27|11|Когда ветви его засохнут, их обломают; женщины придут и сожгут их. Так как это народ безрассудный, то не сжалится над ним Творец его, и не помилует его Создатель его.
ISA|27|12|Но будет в тот день: Господь потрясет все от великой реки до потока Египетского, и вы, сыны Израиля, будете собраны один к другому;
ISA|27|13|и будет в тот день: вострубит великая труба, и придут затерявшиеся в Ассирийской земле и изгнанные в землю Египетскую и поклонятся Господу на горе святой в Иерусалиме.
ISA|28|1|Горе венку гордости пьяных Ефремлян, увядшему цветку красивого убранства его, который на вершине тучной долины сраженных вином!
ISA|28|2|Вот, крепкий и сильный у Господа, как ливень с градом и губительный вихрь, как разлившееся наводнение бурных вод, с силою повергает его на землю.
ISA|28|3|Ногами попирается венок гордости пьяных Ефремлян.
ISA|28|4|И с увядшим цветком красивого убранства его, который на вершине тучной долины, делается то же, что бывает с созревшею прежде времени смоквою, которую, как скоро кто увидит, тотчас берет в руку и проглатывает ее.
ISA|28|5|В тот день Господь Саваоф будет великолепным венцом и славною диадемою для остатка народа Своего,
ISA|28|6|и духом правосудия для сидящего в судилище и мужеством для отражающих неприятеля до ворот.
ISA|28|7|Но и эти шатаются от вина и сбиваются с пути от сикеры; священник и пророк спотыкаются от крепких напитков; побеждены вином, обезумели от сикеры, в видении ошибаются, в суждении спотыкаются.
ISA|28|8|Ибо все столы наполнены отвратительною блевотиною, нет [чистого] места.
ISA|28|9|А [говорят]: "кого хочет он учить ведению? и кого вразумлять проповедью? отнятых от грудного молока, отлученных от сосцов [матери]?
ISA|28|10|Ибо все заповедь на заповедь, заповедь на заповедь, правило на правило, правило на правило, тут немного и там немного".
ISA|28|11|За то лепечущими устами и на чужом языке будут говорить к этому народу.
ISA|28|12|Им говорили: "вот – покой, дайте покой утружденному, и вот успокоение". Но они не хотели слушать.
ISA|28|13|И стало у них словом Господа: заповедь на заповедь, заповедь на заповедь, правило на правило, правило на правило, тут немного, там немного, – так что они пойдут, и упадут навзничь, и разобьются, и попадут в сеть и будут уловлены.
ISA|28|14|Итак слушайте слово Господне, хульники, правители народа сего, который в Иерусалиме.
ISA|28|15|Так как вы говорите: "мы заключили союз со смертью и с преисподнею сделали договор: когда всепоражающий бич будет проходить, он не дойдет до нас, – потому что ложь сделали мы убежищем для себя, и обманом прикроем себя".
ISA|28|16|Посему так говорит Господь Бог: вот, Я полагаю в основание на Сионе камень, камень испытанный, краеугольный, драгоценный, крепко утвержденный: верующий в него не постыдится.
ISA|28|17|И поставлю суд мерилом и правду весами; и градом истребится убежище лжи, и воды потопят место укрывательства.
ISA|28|18|И союз ваш со смертью рушится, и договор ваш с преисподнею не устоит. Когда пойдет всепоражающий бич, вы будете попраны.
ISA|28|19|Как скоро он пойдет, схватит вас; ходить же будет каждое утро, день и ночь, и один слух о нем будет внушать ужас.
ISA|28|20|Слишком коротка будет постель, чтобы протянуться; слишком узко и одеяло, чтобы завернуться в него.
ISA|28|21|Ибо восстанет Господь, как на горе Перациме; разгневается, как на долине Гаваонской, чтобы сделать дело Свое, необычайное дело, и совершить действие Свое, чудное Свое действие.
ISA|28|22|Итак не кощунствуйте, чтобы узы ваши не стали крепче; ибо я слышал от Господа, Бога Саваофа, что истребление определено для всей земли.
ISA|28|23|Приклоните ухо, и послушайте моего голоса; будьте внимательны, и выслушайте речь мою.
ISA|28|24|Всегда ли земледелец пашет для посева, бороздит и боронит землю свою?
ISA|28|25|Нет; когда уровняет поверхность ее, он сеет чернуху, или рассыпает тмин, или разбрасывает пшеницу рядами, и ячмень в определенном месте, и полбу рядом с ним.
ISA|28|26|И такому порядку учит его Бог его; Он наставляет его.
ISA|28|27|Ибо не молотят чернухи катком зубчатым, и колес молотильных не катают по тмину; но палкою выколачивают чернуху, и тмин – палкою.
ISA|28|28|Зерновой хлеб вымолачивают, но не разбивают его; и водят по нему молотильные колеса с конями их, но не растирают его.
ISA|28|29|И это происходит от Господа Саваофа: дивны судьбы Его, велика премудрость Его!
ISA|29|1|Горе Ариилу, Ариилу, городу, в котором жил Давид! приложите год к году; пусть заколают жертвы.
ISA|29|2|Но Я стесню Ариил, и будет плач и сетование; и он останется у Меня, как Ариил.
ISA|29|3|Я расположусь станом вокруг тебя и стесню тебя стражею наблюдательною, и воздвигну против тебя укрепления.
ISA|29|4|И будешь унижен, с земли будешь говорить, и глуха будет речь твоя из–под праха, и голос твой будет, как голос чревовещателя, и из–под праха шептать будет речь твоя.
ISA|29|5|Множество врагов твоих будет, как мелкая пыль, и полчище лютых, как разлетающаяся плева; и это совершится внезапно, в одно мгновение.
ISA|29|6|Господь Саваоф посетит тебя громом и землетрясением, и сильным гласом, бурею и вихрем, и пламенем всепожирающего огня.
ISA|29|7|И как сон, как ночное сновидение, будет множество всех народов, воюющих против Ариила, и всех выступивших против него и укреплений его и стеснивших его.
ISA|29|8|И как голодному снится, будто он ест, но пробуждается, и душа его тоща; и как жаждущему снится, будто он пьет, но пробуждается, и вот он томится, и душа его жаждет: то же будет и множеству всех народов, воюющих против горы Сиона.
ISA|29|9|Изумляйтесь и дивитесь: они ослепили других, и сами ослепли; они пьяны, но не от вина, – шатаются, но не от сикеры;
ISA|29|10|ибо навел на вас Господь дух усыпления и сомкнул глаза ваши, пророки, и закрыл ваши головы, прозорливцы.
ISA|29|11|И всякое пророчество для вас то же, что слова в запечатанной книге, которую подают умеющему читать книгу и говорят: "прочитай ее"; и тот отвечает: "не могу, потому что она запечатана".
ISA|29|12|И передают книгу тому, кто читать не умеет, и говорят: "прочитай ее"; и тот отвечает: "я не умею читать".
ISA|29|13|И сказал Господь: так как этот народ приближается ко Мне устами своими, и языком своим чтит Меня, сердце же его далеко отстоит от Меня, и благоговение их предо Мною есть изучение заповедей человеческих;
ISA|29|14|то вот, Я еще необычайно поступлю с этим народом, чудно и дивно, так что мудрость мудрецов его погибнет, и разума у разумных его не станет.
ISA|29|15|Горе тем, которые думают скрыться в глубину, чтобы замысл свой утаить от Господа, которые делают дела свои во мраке и говорят: "кто увидит нас? и кто узнает нас?"
ISA|29|16|Какое безрассудство! Разве можно считать горшечника, как глину? Скажет ли изделие о сделавшем его: "не он сделал меня"? и скажет ли произведение о художнике своем: "он не разумеет"?
ISA|29|17|Еще немного, очень немного, и Ливан не превратится ли в сад, а сад не будут ли почитать, как лес?
ISA|29|18|И в тот день глухие услышат слова книги, и прозрят из тьмы и мрака глаза слепых.
ISA|29|19|И страждущие более и более будут радоваться о Господе, и бедные люди будут торжествовать о Святом Израиля,
ISA|29|20|потому что не будет более обидчика, и хульник исчезнет, и будут истреблены все поборники неправды,
ISA|29|21|которые запутывают человека в словах, и требующему суда у ворот расставляют сети, и отталкивают правого.
ISA|29|22|Посему так говорит о доме Иакова Господь, Который искупил Авраама: тогда Иаков не будет в стыде, и лице его более не побледнеет.
ISA|29|23|Ибо когда увидит у себя детей своих, дело рук Моих, то они свято будут чтить имя Мое и свято чтить Святаго Иаковлева, и благоговеть пред Богом Израилевым.
ISA|29|24|Тогда блуждающие духом познают мудрость, и непокорные научатся послушанию.
ISA|30|1|Горе непокорным сынам, говорит Господь, которые делают совещания, но без Меня, и заключают союзы, но не по духу Моему, чтобы прилагать грех ко греху:
ISA|30|2|не вопросив уст Моих, идут в Египет, чтобы подкрепить себя силою фараона и укрыться под тенью Египта.
ISA|30|3|Но сила фараона будет для вас стыдом, и убежище под тенью Египта – бесчестием;
ISA|30|4|потому что князья его уже в Цоане, и послы его дошли до Ханеса.
ISA|30|5|Все они будут постыжены из–за народа, [который] бесполезен для них; не будет от него ни помощи, ни пользы, но – стыд и срам.
ISA|30|6|Тяжести на животных, [идущих] на юг, по земле угнетения и тесноты, откуда [выходят] львицы и львы, аспиды и летучие змеи; они несут на хребтах ослов богатства свои и на горбах верблюдов сокровища свои к народу, который не принесет им пользы.
ISA|30|7|Ибо помощь Египта будет тщетна и напрасна; потому Я сказал им: сила их – сидеть спокойно.
ISA|30|8|Теперь пойди, начертай это на доске у них, и впиши это в книгу, чтобы осталось на будущее время, навсегда, навеки.
ISA|30|9|Ибо это народ мятежный, дети лживые, дети, которые не хотят слушать закона Господня,
ISA|30|10|которые провидящим говорят: "перестаньте провидеть", и пророкам: "не пророчествуйте нам правды, говорите нам лестное, предсказывайте приятное;
ISA|30|11|сойдите с дороги, уклонитесь от пути; устраните от глаз наших Святаго Израилева."
ISA|30|12|Посему так говорит Святый Израилев: так как вы отвергаете слово сие, а надеетесь на обман и неправду, и опираетесь на то:
ISA|30|13|то беззаконие это будет для вас, как угрожающая падением трещина, обнаружившаяся в высокой стене, которой разрушение настанет внезапно, в одно мгновение.
ISA|30|14|И Он разрушит ее, как сокрушают глиняный сосуд, разбивая его без пощады, так что в обломках его не найдется и черепка, чтобы взять огня с очага или зачерпнуть воды из водоема;
ISA|30|15|ибо так говорит Господь Бог, Святый Израилев: оставаясь на месте и в покое, вы спаслись бы; в тишине и уповании крепость ваша; но вы не хотели
ISA|30|16|и говорили: "нет, мы на конях убежим", – за то и побежите; "мы на быстрых ускачем", – за то и преследующие вас будут быстры.
ISA|30|17|От угрозы одного [побежит] тысяча, от угрозы пятерых побежите так, что остаток ваш будет как веха на вершине горы и как знамя на холме.
ISA|30|18|И потому Господь медлит, чтобы помиловать вас, и потому еще удерживается, чтобы сжалиться над вами; ибо Господь есть Бог правды: блаженны все уповающие на Него!
ISA|30|19|Народ будет жить на Сионе в Иерусалиме; ты не будешь много плакать, – Он помилует тебя, по голосу вопля твоего, и как только услышит его, ответит тебе.
ISA|30|20|И даст вам Господь хлеб в горести и воду в нужде; и учители твои уже не будут скрываться, и глаза твои будут видеть учителей твоих;
ISA|30|21|и уши твои будут слышать слово, говорящее позади тебя: "вот путь, идите по нему", если бы вы уклонились направо и если бы вы уклонились налево.
ISA|30|22|Тогда вы будете считать скверною оклад идолов из серебра твоего и оклад истуканов из золота твоего; ты бросишь их, как нечистоту; ты скажешь им: прочь отсюда.
ISA|30|23|И Он даст дождь на семя твое, которым засеешь поле, и хлеб, плод земли, и он будет обилен и сочен; стада твои в тот день будут пастись на обширных пастбищах.
ISA|30|24|И волы и ослы, возделывающие поле, будут есть корм соленый, очищенный лопатою и веялом.
ISA|30|25|И на всякой горе высокой и на всяком холме возвышенном потекут ручьи, потоки вод, в день великого поражения, когда упадут башни.
ISA|30|26|И свет луны будет, как свет солнца, а свет солнца будет светлее всемеро, как свет семи дней, в тот день, когда Господь обвяжет рану народа Своего и исцелит нанесенные ему язвы.
ISA|30|27|Вот, имя Господа идет издали, горит гнев Его, и пламя его сильно, уста Его исполнены негодования, и язык Его, как огонь поедающий,
ISA|30|28|и дыхание Его, как разлившийся поток, который поднимается даже до шеи, чтобы развеять народы до истощания; и будет в челюстях народов узда, направляющая к заблуждению.
ISA|30|29|А у вас будут песни, как в ночь священного праздника, и веселие сердца, как у идущего со свирелью на гору Господню, к твердыне Израилевой.
ISA|30|30|И возгремит Господь величественным гласом Своим и явит тяготеющую мышцу Свою в сильном гневе и в пламени поедающего огня, в буре и в наводнении и в каменном граде.
ISA|30|31|Ибо от гласа Господа содрогнется Ассур, жезлом поражаемый.
ISA|30|32|И всякое движение определенного ему жезла, который Господь направит на него, будет с тимпанами и цитрами, и Он пойдет против него войною опустошительною.
ISA|30|33|Ибо Тофет давно уже устроен; он приготовлен и для царя, глубок и широк; в костре его много огня и дров; дуновение Господа, как поток серы, зажжет его.
ISA|31|1|Горе тем, которые идут в Египет за помощью, надеются на коней и полагаются на колесницы, потому что их много, и на всадников, потому что они весьма сильны, а на Святаго Израилева не взирают и к Господу не прибегают!
ISA|31|2|Но премудр Он; и наведет бедствие, и не отменит слов Своих; восстанет против дома нечестивых и против помощи делающих беззаконие.
ISA|31|3|И Египтяне – люди, а не Бог; и кони их – плоть, а не дух. И прострет руку Свою Господь, и споткнется защитник, и упадет защищаемый, и все вместе погибнут.
ISA|31|4|Ибо так сказал мне Господь: как лев, как скимен, ревущий над своею добычею, хотя бы множество пастухов кричало на него, от крика их не содрогнется и множеству их не уступит, – так Господь Саваоф сойдет сразиться за гору Сион и за холм его.
ISA|31|5|Как птицы – птенцов, так Господь Саваоф покроет Иерусалим, защитит и избавит, пощадит и спасет.
ISA|31|6|Обратитесь к Тому, от Которого вы столько отпали, сыны Израиля!
ISA|31|7|В тот день отбросит каждый человек своих серебряных идолов и золотых своих идолов, которых руки ваши сделали вам на грех.
ISA|31|8|И Ассур падет не от человеческого меча, и не человеческий меч потребит его, – он избежит от меча, и юноши его будут податью.
ISA|31|9|И от страха пробежит мимо крепости своей; и князья его будут пугаться знамени, говорит Господь, Которого огонь на Сионе и горнило в Иерусалиме.
ISA|32|1|Вот, Царь будет царствовать по правде, и князья будут править по закону;
ISA|32|2|и каждый из них будет как защита от ветра и покров от непогоды, как источники вод в степи, как тень от высокой скалы в земле жаждущей.
ISA|32|3|И очи видящих не будут закрываемы, и уши слышащих будут внимать.
ISA|32|4|И сердце легкомысленных будет уметь рассуждать; и косноязычные будут говорить ясно.
ISA|32|5|Невежду уже не будут называть почтенным, и о коварном не скажут, что он честный.
ISA|32|6|Ибо невежда говорит глупое, и сердце его помышляет о беззаконном, чтобы действовать лицемерно и произносить хулу на Господа, душу голодного лишать хлеба и отнимать питье у жаждущего.
ISA|32|7|У коварного и действования гибельные: он замышляет ковы, чтобы погубить бедного словами лжи, хотя бы бедный был и прав.
ISA|32|8|А честный и мыслит о честном и твердо стоит во всем, что честно.
ISA|32|9|Женщины беспечные! встаньте, послушайте голоса моего; дочери беззаботные! приклоните слух к моим словам.
ISA|32|10|Еще несколько дней сверх года, и ужаснетесь, беспечные! ибо не будет обирания винограда, и время жатвы не настанет.
ISA|32|11|Содрогнитесь, беззаботные! ужаснитесь, беспечные! сбросьте одежды, обнажитесь и препояшьте чресла.
ISA|32|12|Будут бить себя в грудь о прекрасных полях, о виноградной лозе плодовитой.
ISA|32|13|На земле народа моего будут расти терны и волчцы, равно и на всех домах веселья в ликующем городе;
ISA|32|14|ибо чертоги будут оставлены; шумный город будет покинут; Офел и башня навсегда будут служить, вместо пещер, убежищем диких ослов и пасущихся стад,
ISA|32|15|доколе не излиется на нас Дух свыше, и пустыня не сделается садом, а сад не будут считать лесом.
ISA|32|16|Тогда суд водворится в этой пустыне, и правосудие будет пребывать на плодоносном поле.
ISA|32|17|И делом правды будет мир, и плодом правосудия – спокойствие и безопасность вовеки.
ISA|32|18|Тогда народ мой будет жить в обители мира и в селениях безопасных, и в покоищах блаженных.
ISA|32|19|И град будет падать на лес, и город спустится в долину.
ISA|32|20|Блаженны вы, сеющие при всех водах и посылающие туда вола и осла.
ISA|33|1|Горе тебе, опустошитель, который не был опустошаем, и грабитель, которого не грабили! Когда кончишь опустошение, будешь опустошен и ты; когда прекратишь грабительства, разграбят и тебя.
ISA|33|2|Господи! помилуй нас; на Тебя уповаем мы; будь нашею мышцею с раннего утра и спасением нашим во время тесное.
ISA|33|3|От грозного гласа [Твоего] побегут народы; когда восстанешь, рассеются племена,
ISA|33|4|и будут собирать добычу вашу, как собирает гусеница; бросятся на нее, как бросается саранча.
ISA|33|5|Высок Господь, живущий в вышних; Он наполнит Сион судом и правдою.
ISA|33|6|И настанут безопасные времена твои, изобилие спасения, мудрости и ведения; страх Господень будет сокровищем твоим.
ISA|33|7|Вот, сильные их кричат на улицах; послы для мира горько плачут.
ISA|33|8|Опустели дороги; не стало путешествующих; он нарушил договор, разрушил города, – ни во что ставит людей.
ISA|33|9|Земля сетует, сохнет; Ливан постыжен, увял; Сарон похож стал на пустыню, и обнажены от листьев своих Васан и Кармил.
ISA|33|10|Ныне Я восстану, говорит Господь, ныне поднимусь, ныне вознесусь.
ISA|33|11|Вы беременны сеном, разродитесь соломою; дыхание ваше – огонь, который пожрет вас.
ISA|33|12|И будут народы, [как] горящая известь, [как] срубленный терновник, будут сожжены в огне.
ISA|33|13|Слушайте, дальние, что сделаю Я; и вы, ближние, познайте могущество Мое.
ISA|33|14|Устрашились грешники на Сионе; трепет овладел нечестивыми: "кто из нас может жить при огне пожирающем? кто из нас может жить при вечном пламени?" –
ISA|33|15|Тот, кто ходит в правде и говорит истину; кто презирает корысть от притеснения, удерживает руки свои от взяток, затыкает уши свои, чтобы не слышать о кровопролитии, и закрывает глаза свои, чтобы не видеть зла;
ISA|33|16|тот будет обитать на высотах; убежище его – неприступные скалы; хлеб будет дан ему; вода у него не иссякнет.
ISA|33|17|Глаза твои увидят Царя в красоте Его, узрят землю отдаленную;
ISA|33|18|сердце твое будет [только] вспоминать об ужасах: "где делавший перепись? где весивший [дань]? где осматривающий башни?"
ISA|33|19|Не увидишь более народа свирепого, народа с глухою, невнятною речью, с языком странным, непонятным.
ISA|33|20|Взгляни на Сион, город праздничных собраний наших; глаза твои увидят Иерусалим, жилище мирное, непоколебимую скинию; столпы ее никогда не исторгнутся, и ни одна вервь ее не порвется.
ISA|33|21|Там у нас великий Господь будет вместо рек, вместо широких каналов; туда не войдет ни одно весельное судно, и не пройдет большой корабль.
ISA|33|22|Ибо Господь – судия наш, Господь – законодатель наш, Господь – царь наш; Он спасет нас.
ISA|33|23|Ослабли веревки твои, не могут удержать мачты и натянуть паруса. Тогда будет большой раздел добычи, так что и хромые пойдут на грабеж.
ISA|33|24|И ни один из жителей не скажет: "я болен"; народу, живущему там, будут отпущены согрешения.
ISA|34|1|Приступите, народы, слушайте и внимайте, племена! да слышит земля и все, что наполняет ее, вселенная и все рождающееся в ней!
ISA|34|2|Ибо гнев Господа на все народы, и ярость Его на все воинство их. Он предал их заклятию, отдал их на заклание.
ISA|34|3|И убитые их будут разбросаны, и от трупов их поднимется смрад, и горы размокнут от крови их.
ISA|34|4|И истлеет все небесное воинство; и небеса свернутся, как свиток книжный; и все воинство их падет, как спадает лист с виноградной лозы, и как увядший лист – со смоковницы.
ISA|34|5|Ибо упился меч Мой на небесах: вот, для суда нисходит он на Едом и на народ, преданный Мною заклятию.
ISA|34|6|Меч Господа наполнится кровью, утучнеет от тука, от крови агнцев и козлов, от тука с почек овнов: ибо жертва у Господа в Восоре и большое заклание в земле Едома.
ISA|34|7|И буйволы падут с ними и тельцы вместе с волами, и упьется земля их кровью, и прах их утучнеет от тука.
ISA|34|8|Ибо день мщения у Господа, год возмездия за Сион.
ISA|34|9|И превратятся реки его в смолу, и прах его – в серу, и будет земля его горящею смолою:
ISA|34|10|не будет гаснуть ни днем, ни ночью; вечно будет восходить дым ее; будет от рода в род оставаться опустелою; во веки веков никто не пройдет по ней;
ISA|34|11|и завладеют ею пеликан и еж; и филин и ворон поселятся в ней; и протянут по ней вервь разорения и отвес уничтожения.
ISA|34|12|Никого не останется там из знатных ее, кого можно было бы призвать на царство, и все князья ее будут ничто.
ISA|34|13|И зарастут дворцы ее колючими растениями, крапивою и репейником – твердыни ее; и будет она жилищем шакалов, пристанищем страусов.
ISA|34|14|И звери пустыни будут встречаться с дикими кошками, и лешие будут перекликаться один с другим; там будет отдыхать ночное привидение и находить себе покой.
ISA|34|15|Там угнездится летучий змей, будет класть яйца и выводить детей и собирать их под тень свою; там и коршуны будут собираться один к другому.
ISA|34|16|Отыщите в книге Господней и прочитайте; ни одно из сих не преминет придти, и одно другим не заменится. Ибо сами уста Его повелели, и сам дух Его соберет их.
ISA|34|17|И Сам Он бросил им жребий, и Его рука разделила им ее мерою; во веки будут они владеть ею, из рода в род будут жить на ней.
ISA|35|1|Возвеселится пустыня и сухая земля, и возрадуется страна необитаемая и расцветет как нарцисс;
ISA|35|2|великолепно будет цвести и радоваться, будет торжествовать и ликовать; слава Ливана дастся ей, великолепие Кармила и Сарона; они увидят славу Господа, величие Бога нашего.
ISA|35|3|Укрепите ослабевшие руки и утвердите колени дрожащие;
ISA|35|4|скажите робким душею: будьте тверды, не бойтесь; вот Бог ваш, придет отмщение, воздаяние Божие; Он придет и спасет вас.
ISA|35|5|Тогда откроются глаза слепых, и уши глухих отверзутся.
ISA|35|6|Тогда хромой вскочит, как олень, и язык немого будет петь; ибо пробьются воды в пустыне, и в степи – потоки.
ISA|35|7|И превратится призрак вод в озеро, и жаждущая земля – в источники вод; в жилище шакалов, где они покоятся, будет место для тростника и камыша.
ISA|35|8|И будет там большая дорога, и путь по ней назовется путем святым: нечистый не будет ходить по нему; но он будет для них [одних]; идущие этим путем, даже и неопытные, не заблудятся.
ISA|35|9|Льва не будет там, и хищный зверь не взойдет на него; его не найдется там, а будут ходить искупленные.
ISA|35|10|И возвратятся избавленные Господом, придут на Сион с радостным восклицанием; и радость вечная будет над головою их; они найдут радость и веселье, а печаль и воздыхание удалятся.
ISA|36|1|И было в четырнадцатый год царя Езекии, пошел Сеннахирим, царь Ассирийский, против всех укрепленных городов Иудеи и взял их.
ISA|36|2|И послал царь Ассирийский из Лахиса в Иерусалим к царю Езекии Рабсака с большим войском; и он остановился у водопровода верхнего пруда на дороге поля белильничьего.
ISA|36|3|И вышел к нему Елиаким, сын Хелкиин, начальник дворца, и Севна писец, и Иоах, сын Асафов, дееписатель.
ISA|36|4|И сказал им Рабсак: скажите Езекии: так говорит царь великий, царь Ассирийский: что это за упование, на которое ты уповаешь?
ISA|36|5|Я думаю, [что] это одни пустые слова, [а] для войны нужны совет и сила: итак на кого ты уповаешь, что отложился от меня?
ISA|36|6|Вот, ты думаешь опереться на Египет, на эту трость надломленную, которая, если кто опрется на нее, войдет тому в руку и проколет ее! Таков фараон, царь Египетский, для всех уповающих на него.
ISA|36|7|А если скажешь мне: "на Господа, Бога нашего мы уповаем", то на того ли, которого высоты и жертвенники отменил Езекия и сказал Иуде и Иерусалиму: "пред сим только жертвенником поклоняйтесь"?
ISA|36|8|Итак вступи в союз с господином моим, царем Ассирийским; я дам тебе две тысячи коней; можешь ли достать себе всадников на них?
ISA|36|9|И как ты хочешь заставить отступить вождя, одного из малейших рабов господина моего, надеясь на Египет, ради колесниц и коней?
ISA|36|10|Да разве я без воли Господней пошел на землю сию, чтобы разорить ее? Господь сказал мне: пойди на землю сию и разори ее.
ISA|36|11|И сказал Елиаким и Севна и Иоах Рабсаку: говори рабам твоим по–арамейски, потому что мы понимаем, а не говори с нами по–иудейски, вслух народа, который на стене.
ISA|36|12|И сказал Рабсак: разве [только] к господину твоему и к тебе послал меня господин мой сказать слова сии? Нет, [также] и к людям, которые сидят на стене, чтобы есть помет свой и пить мочу свою с вами.
ISA|36|13|И встал Рабсак, и возгласил громким голосом по–иудейски, и сказал: слушайте слово царя великого, царя Ассирийского!
ISA|36|14|Так говорит царь: пусть не обольщает вас Езекия, ибо он не может спасти вас;
ISA|36|15|и пусть не обнадеживает вас Езекия Господом, говоря: "спасет нас Господь; не будет город сей отдан в руки царя Ассирийского".
ISA|36|16|Не слушайте Езекии, ибо так говорит царь Ассирийский: примиритесь со мною и выйдите ко мне, и пусть каждый ест плоды виноградной лозы своей и смоковницы своей, и пусть каждый пьет воду из своего колодезя,
ISA|36|17|доколе я не приду и не возьму вас в землю такую же, как и ваша земля, в землю хлеба и вина, в землю плодов и виноградников.
ISA|36|18|[Итак] да не обольщает вас Езекия, говоря: "Господь спасет нас". Спасли ли боги народов, каждый свою землю, от руки царя Ассирийского?
ISA|36|19|Где боги Емафа и Арпада? Где боги Сепарваима? Спасли ли они Самарию от руки моей?
ISA|36|20|Который из всех богов земель сих спас землю свою от руки моей? Так неужели спасет Господь Иерусалим от руки моей?
ISA|36|21|Но они молчали и не отвечали ему ни слова, потому что от царя дано было приказание: не отвечайте ему.
ISA|36|22|И пришел Елиаким, сын Хелкиин, начальник дворца, и Севна писец, и Иоах, сын Асафов, дееписатель, к Езекии в разодранных одеждах и пересказали ему слова Рабсака.
ISA|37|1|Когда услышал это царь Езекия, то разодрал одежды свои и покрылся вретищем, и пошел в дом Господень;
ISA|37|2|и послал Елиакима, начальника дворца, и Севну писца, и старших священников, покрытых вретищами, к пророку Исаии, сыну Амосову.
ISA|37|3|И они сказали ему: так говорит Езекия: день скорби и наказания и посрамления день сей, ибо младенцы дошли до отверстия утробы матерней, а силы нет родить.
ISA|37|4|Может быть, услышит Господь Бог твой слова Рабсака, которого послал царь Ассирийский, господин его, хулить Бога живаго и поносить словами, какие слышал Господь, Бог твой; вознеси же молитву об оставшихся, которые находятся еще в живых.
ISA|37|5|И пришли слуги царя Езекии к Исаии.
ISA|37|6|И сказал им Исаия: так скажите господину вашему: так говорит Господь: не бойся слов, которые слышал ты, которыми поносили Меня слуги царя Ассирийского.
ISA|37|7|Вот, Я пошлю в него дух, и он услышит весть, и возвратится в землю свою, и Я поражу его мечом в земле его.
ISA|37|8|И возвратился Рабсак и нашел царя Ассирийского воюющим против Ливны; ибо он слышал, что тот отошел от Лахиса.
ISA|37|9|И услышал он о Тиргаке, царе Ефиопском; [ему] сказали: вот, он вышел сразиться с тобою. Услышав это, он послал послов к Езекии, сказав:
ISA|37|10|так скажите Езекии, царю Иудейскому: пусть не обманывает тебя Бог твой, на Которого ты уповаешь, думая: "не будет отдан Иерусалим в руки царя Ассирийского".
ISA|37|11|Вот, ты слышал, что сделали цари Ассирийские со всеми землями, положив на них заклятие; ты ли уцелеешь?
ISA|37|12|Боги народов, которых разорили отцы мои, спасли ли их, [спасли] [ли] Гозан и Харан, и Рецеф, и сынов Едена, что в Фалассаре?
ISA|37|13|Где царь Емафа и царь Арпада, и царь города Сепарваима, Ены и Иввы?
ISA|37|14|И взял Езекия письмо из руки послов и прочитал его, и пошел в дом Господень, и развернул его Езекия пред лицем Господним;
ISA|37|15|и молился Езекия пред лицем Господним и говорил:
ISA|37|16|Господи Саваоф, Боже Израилев, седящий на Херувимах! Ты один Бог всех царств земли; Ты сотворил небо и землю.
ISA|37|17|Приклони, Господи, ухо Твое и услышь; открой, Господи, очи Твои и воззри, и услышь слова Сеннахирима, который послал поносить Тебя, Бога живаго.
ISA|37|18|Правда, о, Господи! цари Ассирийские опустошили все страны и земли их
ISA|37|19|и побросали богов их в огонь; но это были не боги, а изделие рук человеческих, дерево и камень, потому и истребили их.
ISA|37|20|И ныне, Господи Боже наш, спаси нас от руки его; и узнают все царства земли, что Ты, Господи, Бог один.
ISA|37|21|И послал Исаия, сын Амосов, к Езекии сказать: так говорит Господь, Бог Израилев: о чем ты молился Мне против Сеннахирима, царя Ассирийского, –
ISA|37|22|вот слово, которое Господь изрек о нем: презрит тебя, посмеется над тобою девствующая дочь Сиона, покачает вслед тебя головою дочь Иерусалима.
ISA|37|23|Кого ты порицал и поносил? и на кого возвысил голос и поднял так высоко глаза твои? на Святаго Израилева.
ISA|37|24|Чрез рабов твоих ты порицал Господа и сказал: "со множеством колесниц моих я взошел на высоту гор, на ребра Ливана, и срубил рослые кедры его, отличные кипарисы его, и пришел на самую вершину его, в рощу сада его;
ISA|37|25|и откапывал я, и пил воду; и осушу ступнями ног моих все реки Египетские".
ISA|37|26|Разве не слышал ты, что Я издавна сделал это, в древние дни предначертал это, а ныне выполнил тем, что ты опустошаешь крепкие города, [превращая] их в груды развалин?
ISA|37|27|И жители их сделались маломощны, трепещут и остаются в стыде; они стали как трава на поле и нежная зелень, как порост на кровлях и опаленный хлеб, прежде нежели выколосился.
ISA|37|28|Сядешь ли ты, выйдешь ли, войдешь ли, Я знаю [все, знаю] и дерзость твою против Меня.
ISA|37|29|За твою дерзость против Меня и за то, что надмение твое дошло до ушей Моих, Я вложу кольцо Мое в ноздри твои и удила Мои в рот твой, и возвращу тебя назад тою же дорогою, которою ты пришел.
ISA|37|30|И вот, тебе, Езекия, знамение: ешьте в этот год выросшее от упавшего зерна, и на другой год – самородное; а на третий год сейте и жните, и садите виноградные сады, и ешьте плоды их.
ISA|37|31|И уцелевший в доме Иудином остаток пустит опять корень внизу и принесет плод вверху,
ISA|37|32|ибо из Иерусалима произойдет остаток, и спасенное – от горы Сиона. Ревность Господа Саваофа соделает это.
ISA|37|33|Посему так говорит Господь о царе Ассирийском: "не войдет он в этот город и не бросит туда стрелы, и не приступит к нему со щитом, и не насыплет против него вала.
ISA|37|34|По той же дороге, по которой пришел, возвратится, а в город сей не войдет, говорит Господь.
ISA|37|35|Я буду охранять город сей, чтобы спасти его ради Себя и ради Давида, раба Моего".
ISA|37|36|И вышел Ангел Господень и поразил в стане Ассирийском сто восемьдесят пять тысяч [человек]. И встали поутру, и вот, все тела мертвые.
ISA|37|37|И отступил, и пошел, и возвратился Сеннахирим, царь Ассирийский, и жил в Ниневии.
ISA|37|38|И когда он поклонялся в доме Нисроха, бога своего, Адрамелех и Шарецер, сыновья его, убили его мечом, а сами убежали в землю Араратскую. И воцарился Асардан, сын его, вместо него.
ISA|38|1|В те дни Езекия заболел смертельно. И пришел к нему пророк Исаия, сын Амосов, и сказал ему: так говорит Господь: сделай завещание для дома твоего, ибо ты умрешь, не выздоровеешь.
ISA|38|2|Тогда Езекия отворотился лицем к стене и молился Господу, говоря:
ISA|38|3|"о, Господи! вспомни, что я ходил пред лицем Твоим верно и с преданным [Тебе] сердцем и делал угодное в очах Твоих". И заплакал Езекия сильно.
ISA|38|4|И было слово Господне к Исаии, и сказано:
ISA|38|5|пойди и скажи Езекии: так говорит Господь, Бог Давида, отца твоего: Я услышал молитву твою, увидел слезы твои, и вот, Я прибавлю к дням твоим пятнадцать лет,
ISA|38|6|и от руки царя Ассирийского спасу тебя и город сей и защищу город сей.
ISA|38|7|И вот тебе знамение от Господа, что Господь исполнит слово, которое Он изрек.
ISA|38|8|Вот, я возвращу назад на десять ступеней солнечную тень, которая прошла по ступеням Ахазовым. И возвратилось солнце на десять ступеней по ступеням, по которым оно сходило.
ISA|38|9|Молитва Езекии, царя Иудейского, когда он болен был и выздоровел от болезни:
ISA|38|10|"Я сказал в себе: в преполовение дней моих должен я идти во врата преисподней; я лишен остатка лет моих.
ISA|38|11|Я говорил: не увижу я Господа, Господа на земле живых; не увижу больше человека между живущими в мире;
ISA|38|12|жилище мое снимается с места и уносится от меня, как шалаш пастушеский; я должен отрезать подобно ткачу жизнь мою; Он отрежет меня от основы; день и ночь я ждал, что Ты пошлешь мне кончину.
ISA|38|13|Я ждал до утра; подобно льву, Он сокрушал все кости мои; день и ночь я ждал, что Ты пошлешь мне кончину.
ISA|38|14|Как журавль, как ласточка издавал я звуки, тосковал как голубь; уныло смотрели глаза мои к небу: Господи! тесно мне; спаси меня.
ISA|38|15|Что скажу я? Он сказал мне, Он и сделал. Тихо буду проводить все годы жизни моей, помня горесть души моей.
ISA|38|16|Господи! так живут, и во всем этом жизнь моего духа; Ты исцелишь меня, даруешь мне жизнь.
ISA|38|17|Вот, во благо мне была сильная горесть, и Ты избавил душу мою от рва погибели, бросил все грехи мои за хребет Свой.
ISA|38|18|Ибо не преисподняя славит Тебя, не смерть восхваляет Тебя, не нисшедшие в могилу уповают на истину Твою.
ISA|38|19|Живой, только живой прославит Тебя, как я ныне: отец возвестит детям истину Твою.
ISA|38|20|Господь спасет меня; и мы во все дни жизни нашей [со звуками] струн моих будем воспевать песни в доме Господнем".
ISA|38|21|И сказал Исаия: пусть принесут пласт смокв и обложат им нарыв; и он выздоровеет.
ISA|38|22|А Езекия сказал: какое знамение, что я буду ходить в дом Господень?
ISA|39|1|В то время Меродах Валадан, сын Валадана, царь Вавилонский, прислал к Езекии письмо и дары, ибо слышал, что он был болен и выздоровел.
ISA|39|2|И обрадовался посланным Езекия, и показал им дом сокровищ своих, серебро и золото, и ароматы, и драгоценные масти, весь оружейный свой дом и все, что находилось в сокровищницах его; ничего не осталось, чего не показал бы им Езекия в доме своем и во всем владении своем.
ISA|39|3|И пришел пророк Исаия к царю Езекии и сказал ему: что говорили эти люди? и откуда они приходили к тебе? Езекия сказал: из далекой земли приходили они ко мне, из Вавилона.
ISA|39|4|И сказал [Исаия]: что видели они в доме твоем? Езекия сказал: видели все, что есть в доме моем; ничего не осталось в сокровищницах моих, чего я не показал бы им.
ISA|39|5|И сказал Исаия Езекии: выслушай слово Господа Саваофа:
ISA|39|6|вот, придут дни, и все, что есть в доме твоем и что собрали отцы твои до сего дня, будет унесено в Вавилон; ничего не останется, говорит Господь.
ISA|39|7|И возьмут из сыновей твоих, которые произойдут от тебя, которых ты родишь, – и они будут евнухами во дворце царя Вавилонского.
ISA|39|8|И сказал Езекия Исаии: благо слово Господне, которое ты изрек; потому что, присовокупил он, мир и благосостояние пребудут во дни мои.
ISA|40|1|Утешайте, утешайте народ Мой, говорит Бог ваш;
ISA|40|2|говорите к сердцу Иерусалима и возвещайте ему, что исполнилось время борьбы его, что за неправды его сделано удовлетворение, ибо он от руки Господней принял вдвое за все грехи свои.
ISA|40|3|Глас вопиющего в пустыне: приготовьте путь Господу, прямыми сделайте в степи стези Богу нашему;
ISA|40|4|всякий дол да наполнится, и всякая гора и холм да понизятся, кривизны выпрямятся и неровные пути сделаются гладкими;
ISA|40|5|и явится слава Господня, и узрит всякая плоть [спасение Божие]; ибо уста Господни изрекли это.
ISA|40|6|Голос говорит: возвещай! И сказал: что мне возвещать? Всякая плоть – трава, и вся красота ее – как цвет полевой.
ISA|40|7|Засыхает трава, увядает цвет, когда дунет на него дуновение Господа: так и народ – трава.
ISA|40|8|Трава засыхает, цвет увядает, а слово Бога нашего пребудет вечно.
ISA|40|9|Взойди на высокую гору, благовествующий Сион! возвысь с силою голос твой, благовествующий Иерусалим! возвысь, не бойся; скажи городам Иудиным: вот Бог ваш!
ISA|40|10|Вот, Господь Бог грядет с силою, и мышца Его со властью. Вот, награда Его с Ним и воздаяние Его пред лицем Его.
ISA|40|11|Как пастырь Он будет пасти стадо Свое; агнцев будет брать на руки и носить на груди Своей, и водить дойных.
ISA|40|12|Кто исчерпал воды горстью своею и пядью измерил небеса, и вместил в меру прах земли, и взвесил на весах горы и на чашах весовых холмы?
ISA|40|13|Кто уразумел дух Господа, и был советником у Него и учил Его?
ISA|40|14|С кем советуется Он, и кто вразумляет Его и наставляет Его на путь правды, и учит Его знанию, и указывает Ему путь мудрости?
ISA|40|15|Вот народы – как капля из ведра, и считаются как пылинка на весах. Вот, острова как порошинку поднимает Он.
ISA|40|16|И Ливана недостаточно для жертвенного огня, и животных на нем – для всесожжения.
ISA|40|17|Все народы пред Ним как ничто, – менее ничтожества и пустоты считаются у Него.
ISA|40|18|Итак кому уподобите вы Бога? И какое подобие найдете Ему?
ISA|40|19|Идола выливает художник, и золотильщик покрывает его золотом и приделывает серебряные цепочки.
ISA|40|20|А кто беден для такого приношения, выбирает негниющее дерево, приискивает себе искусного художника, чтобы сделать идола, который стоял бы твердо.
ISA|40|21|Разве не знаете? разве вы не слышали? разве вам не говорено было от начала? разве вы не уразумели из оснований земли?
ISA|40|22|Он есть Тот, Который восседает над кругом земли, и живущие на ней – как саранча [пред Ним]; Он распростер небеса, как тонкую ткань, и раскинул их, как шатер для жилья.
ISA|40|23|Он обращает князей в ничто, делает чем–то пустым судей земли.
ISA|40|24|Едва они посажены, едва посеяны, едва укоренился в земле ствол их, и как только Он дохнул на них, они высохли, и вихрь унес их, как солому.
ISA|40|25|Кому же вы уподобите Меня и с кем сравните? говорит Святый.
ISA|40|26|Поднимите глаза ваши на высоту [небес] и посмотрите, кто сотворил их? Кто выводит воинство их счетом? Он всех их называет по имени: по множеству могущества и великой силе у Него ничто не выбывает.
ISA|40|27|Как же говоришь ты, Иаков, и высказываешь, Израиль: "путь мой сокрыт от Господа, и дело мое забыто у Бога моего"?
ISA|40|28|Разве ты не знаешь? разве ты не слышал, что вечный Господь Бог, сотворивший концы земли, не утомляется и не изнемогает? разум Его неисследим.
ISA|40|29|Он дает утомленному силу, и изнемогшему дарует крепость.
ISA|40|30|Утомляются и юноши и ослабевают, и молодые люди падают,
ISA|40|31|а надеющиеся на Господа обновятся в силе: поднимут крылья, как орлы, потекут – и не устанут, пойдут – и не утомятся.
ISA|41|1|Умолкните предо Мною, острова, и народы да обновят свои силы; пусть они приблизятся и скажут: "станем вместе на суд".
ISA|41|2|Кто воздвиг от востока мужа правды, призвал его следовать за собою, предал ему народы и покорил царей? Он обратил их мечом его в прах, луком его в солому, разносимую ветром.
ISA|41|3|Он гонит их, идет спокойно дорогою, по которой никогда не ходил ногами своими.
ISA|41|4|Кто сделал и совершил это? Тот, Кто от начала вызывает роды; Я – Господь первый, и в последних – Я тот же.
ISA|41|5|Увидели острова и ужаснулись, концы земли затрепетали. Они сблизились и сошлись;
ISA|41|6|каждый помогает своему товарищу и говорит своему брату: "крепись!"
ISA|41|7|Кузнец ободряет плавильщика, разглаживающий листы молотом – кующего на наковальне, говоря о спайке: "хороша"; и укрепляет гвоздями, чтобы было твердо.
ISA|41|8|А ты, Израиль, раб Мой, Иаков, которого Я избрал, семя Авраама, друга Моего, –
ISA|41|9|ты, которого Я взял от концов земли и призвал от краев ее, и сказал тебе: "ты Мой раб, Я избрал тебя и не отвергну тебя":
ISA|41|10|не бойся, ибо Я с тобою; не смущайся, ибо Я Бог твой; Я укреплю тебя, и помогу тебе, и поддержу тебя десницею правды Моей.
ISA|41|11|Вот, в стыде и посрамлении останутся все, раздраженные против тебя; будут как ничто и погибнут препирающиеся с тобою.
ISA|41|12|Будешь искать их, и не найдешь их, враждующих против тебя; борющиеся с тобою будут как ничто, совершенно ничто;
ISA|41|13|ибо Я Господь, Бог твой; держу тебя за правую руку твою, говорю тебе: "не бойся, Я помогаю тебе".
ISA|41|14|Не бойся, червь Иаков, малолюдный Израиль, – Я помогаю тебе, говорит Господь и Искупитель твой, Святый Израилев.
ISA|41|15|Вот, Я сделал тебя острым молотилом, новым, зубчатым; ты будешь молотить и растирать горы, и холмы сделаешь, как мякину.
ISA|41|16|Ты будешь веять их, и ветер разнесет их, и вихрь развеет их; а ты возрадуешься о Господе, будешь хвалиться Святым Израилевым.
ISA|41|17|Бедные и нищие ищут воды, и нет [ее]; язык их сохнет от жажды: Я, Господь, услышу их, Я, Бог Израилев, не оставлю их.
ISA|41|18|Открою на горах реки и среди долин источники; пустыню сделаю озером и сухую землю – источниками воды;
ISA|41|19|посажу в пустыне кедр, ситтим и мирту и маслину; насажу в степи кипарис, явор и бук вместе,
ISA|41|20|чтобы увидели и познали, и рассмотрели и уразумели, что рука Господня соделала это, и Святый Израилев сотворил сие.
ISA|41|21|Представьте дело ваше, говорит Господь; приведите ваши доказательства, говорит Царь Иакова.
ISA|41|22|Пусть они представят и скажут нам, что произойдет; пусть возвестят что–либо прежде, нежели оно произошло, и мы вникнем умом своим и узнаем, как оно кончилось, или пусть предвозвестят нам о будущем.
ISA|41|23|Скажите, что произойдет в будущем, и мы будем знать, что вы боги, или сделайте что–нибудь, доброе ли, худое ли, чтобы мы изумились и вместе с вами увидели.
ISA|41|24|Но вы ничто, и дело ваше ничтожно; мерзость тот, кто избирает вас.
ISA|41|25|Я воздвиг его от севера, и он придет; от восхода солнца будет призывать имя Мое и попирать владык, как грязь, и топтать, как горшечник глину.
ISA|41|26|Кто возвестил об этом изначала, чтобы нам знать, и задолго пред тем, чтобы нам можно было сказать: "правда"? Но никто не сказал, никто не возвестил, никто не слыхал слов ваших.
ISA|41|27|Я первый [сказал] Сиону: "вот оно!" и дал Иерусалиму благовестника.
ISA|41|28|Итак Я смотрел, и не было никого, и между ними не нашлось советника, чтоб Я мог спросить их, и они дали ответ.
ISA|41|29|Вот, все они ничто, ничтожны и дела их; ветер и пустота истуканы их.
ISA|42|1|Вот, Отрок Мой, Которого Я держу за руку, избранный Мой, к которому благоволит душа Моя. Положу дух Мой на Него, и возвестит народам суд;
ISA|42|2|не возопиет и не возвысит голоса Своего, и не даст услышать его на улицах;
ISA|42|3|трости надломленной не переломит, и льна курящегося не угасит; будет производить суд по истине;
ISA|42|4|не ослабеет и не изнеможет, доколе на земле не утвердит суда, и на закон Его будут уповать острова.
ISA|42|5|Так говорит Господь Бог, сотворивший небеса и пространство их, распростерший землю с произведениями ее, дающий дыхание народу на ней и дух ходящим по ней.
ISA|42|6|Я, Господь, призвал Тебя в правду, и буду держать Тебя за руку и хранить Тебя, и поставлю Тебя в завет для народа, во свет для язычников,
ISA|42|7|чтобы открыть глаза слепых, чтобы узников вывести из заключения и сидящих во тьме – из темницы.
ISA|42|8|Я Господь, это – Мое имя, и не дам славы Моей иному и хвалы Моей истуканам.
ISA|42|9|Вот, [предсказанное] прежде сбылось, и новое Я возвещу; прежде нежели оно произойдет, Я возвещу вам.
ISA|42|10|Пойте Господу новую песнь, хвалу Ему от концов земли, вы, плавающие по морю, и все, наполняющее его, острова и живущие на них.
ISA|42|11|Да возвысит голос пустыня и города ее, селения, где обитает Кидар; да торжествуют живущие на скалах, да возглашают с вершин гор.
ISA|42|12|Да воздадут Господу славу, и хвалу Его да возвестят на островах.
ISA|42|13|Господь выйдет, как исполин, как муж браней возбудит ревность; воззовет и поднимет воинский крик, и покажет Себя сильным против врагов Своих.
ISA|42|14|Долго молчал Я, терпел, удерживался; теперь буду кричать, как рождающая, буду разрушать и поглощать все;
ISA|42|15|опустошу горы и холмы, и всю траву их иссушу; и реки сделаю островами, и осушу озера;
ISA|42|16|и поведу слепых дорогою, которой они не знают, неизвестными путями буду вести их; мрак сделаю светом пред ними, и кривые пути – прямыми: вот что Я сделаю для них и не оставлю их.
ISA|42|17|Тогда обратятся вспять и великим стыдом покроются надеющиеся на идолов, говорящие истуканам: "вы наши боги".
ISA|42|18|Слушайте, глухие, и смотрите, слепые, чтобы видеть.
ISA|42|19|Кто так слеп, как раб Мой, и глух, как вестник Мой, Мною посланный? Кто так слеп, как возлюбленный, так слеп, как раб Господа?
ISA|42|20|Ты видел многое, но не замечал; уши были открыты, но не слышал.
ISA|42|21|Господу угодно было, ради правды Своей, возвеличить и прославить закон.
ISA|42|22|Но это народ разоренный и разграбленный; все они связаны в подземельях и сокрыты в темницах; сделались добычею, и нет избавителя; ограблены, и никто не говорит: "отдай назад!"
ISA|42|23|Кто из вас приклонил к этому ухо, вникнул и выслушал это для будущего?
ISA|42|24|Кто предал Иакова на разорение и Израиля грабителям? не Господь ли, против Которого мы грешили? Не хотели они ходить путями Его и не слушали закона Его.
ISA|42|25|И Он излил на них ярость гнева Своего и лютость войны: она окружила их пламенем со всех сторон, но они не примечали; и горела у них, но они не уразумели этого сердцем.
ISA|43|1|Ныне же так говорит Господь, сотворивший тебя, Иаков, и устроивший тебя, Израиль: не бойся, ибо Я искупил тебя, назвал тебя по имени твоему; ты Мой.
ISA|43|2|Будешь ли переходить через воды, Я с тобою, – через реки ли, они не потопят тебя; пойдешь ли через огонь, не обожжешься, и пламя не опалит тебя.
ISA|43|3|Ибо Я Господь, Бог твой, Святый Израилев, Спаситель твой; в выкуп за тебя отдал Египет, Ефиопию и Савею за тебя.
ISA|43|4|Так как ты дорог в очах Моих, многоценен, и Я возлюбил тебя, то отдам [других] людей за тебя, и народы за душу твою.
ISA|43|5|Не бойся, ибо Я с тобою; от востока приведу племя твое и от запада соберу тебя.
ISA|43|6|Северу скажу: "отдай"; и югу: "не удерживай; веди сыновей Моих издалека и дочерей Моих от концов земли,
ISA|43|7|каждого кто называется Моим именем, кого Я сотворил для славы Моей, образовал и устроил.
ISA|43|8|Выведи народ слепой, хотя у него есть глаза, и глухой, хотя у него есть уши".
ISA|43|9|Пусть все народы соберутся вместе, и совокупятся племена. Кто между ними предсказал это? пусть возвестят, что было от начала; пусть представят свидетелей от себя и оправдаются, чтобы можно было услышать и сказать: "правда!"
ISA|43|10|А Мои свидетели, говорит Господь, вы и раб Мой, которого Я избрал, чтобы вы знали и верили Мне, и разумели, что это Я: прежде Меня не было Бога и после Меня не будет.
ISA|43|11|Я, Я Господь, и нет Спасителя кроме Меня.
ISA|43|12|Я предрек и спас, и возвестил; а иного нет у вас, и вы – свидетели Мои, говорит Господь, что Я Бог;
ISA|43|13|от [начала] дней Я Тот же, и никто не спасет от руки Моей; Я сделаю, и кто отменит это?
ISA|43|14|Так говорит Господь, Искупитель ваш, Святый Израилев: ради вас Я послал в Вавилон и сокрушил все запоры и Халдеев, величавшихся кораблями.
ISA|43|15|Я Господь, Святый ваш, Творец Израиля, Царь ваш.
ISA|43|16|Так говорит Господь, открывший в море дорогу, в сильных водах стезю,
ISA|43|17|выведший колесницы и коней, войско и силу; все легли вместе, не встали; потухли как светильня, погасли.
ISA|43|18|Но вы не вспоминаете прежнего и о древнем не помышляете.
ISA|43|19|Вот, Я делаю новое; ныне же оно явится; неужели вы и этого не хотите знать? Я проложу дорогу в степи, реки в пустыне.
ISA|43|20|Полевые звери прославят Меня, шакалы и страусы, потому что Я в пустынях дам воду, реки в сухой степи, чтобы поить избранный народ Мой.
ISA|43|21|Этот народ Я образовал для Себя; он будет возвещать славу Мою.
ISA|43|22|А ты, Иаков, не взывал ко Мне; ты, Израиль, не трудился для Меня.
ISA|43|23|Ты не приносил Мне агнцев твоих во всесожжение и жертвами твоими не чтил Меня. Я не заставлял тебя служить Мне хлебным приношением и не отягощал тебя фимиамом.
ISA|43|24|Ты не покупал Мне благовонной трости за серебро и туком жертв твоих не насыщал Меня; но ты грехами твоими затруднял Меня, беззакониями твоими отягощал Меня.
ISA|43|25|Я, Я Сам изглаживаю преступления твои ради Себя Самого и грехов твоих не помяну:
ISA|43|26|припомни Мне; станем судиться; говори ты, чтоб оправдаться.
ISA|43|27|Праотец твой согрешил, и ходатаи твои отступили от Меня.
ISA|43|28|За то Я предстоятелей святилища лишил священства и Иакова предал на заклятие и Израиля на поругание.
ISA|44|1|А ныне слушай, Иаков, раб Мой, и Израиль, которого Я избрал.
ISA|44|2|Так говорит Господь, создавший тебя и образовавший тебя, помогающий тебе от утробы матерней: не бойся, раб Мой, Иаков, и возлюбленный [Израиль], которого Я избрал;
ISA|44|3|ибо Я изолью воды на жаждущее и потоки на иссохшее; излию дух Мой на племя твое и благословение Мое на потомков твоих.
ISA|44|4|И будут расти между травою, как ивы при потоках вод.
ISA|44|5|Один скажет: "я Господень", другой назовется именем Иакова; а иной напишет рукою своею: "я Господень", и прозовется именем Израиля.
ISA|44|6|Так говорит Господь, Царь Израиля, и Искупитель его, Господь Саваоф: Я первый и Я последний, и кроме Меня нет Бога,
ISA|44|7|ибо кто как Я? Пусть он расскажет, возвестит и в порядке представит Мне [все] с того времени, как Я устроил народ древний, или пусть возвестят наступающее и будущее.
ISA|44|8|Не бойтесь и не страшитесь: не издавна ли Я возвестил тебе и предсказал? И вы Мои свидетели. Есть ли Бог кроме Меня? нет другой твердыни, никакой не знаю.
ISA|44|9|Делающие идолов все ничтожны, и вожделеннейшие их не приносят никакой пользы, и они сами себе свидетели в том. Они не видят и не разумеют, и потому будут посрамлены.
ISA|44|10|Кто сделал бога и вылил идола, не приносящего никакой пользы?
ISA|44|11|Все участвующие в этом будут постыжены, ибо и художники сами из людей же; пусть все они соберутся и станут; они устрашатся, и все будут постыжены.
ISA|44|12|Кузнец делает из железа топор и работает на угольях, молотами обделывает его и трудится над ним сильною рукою своею до того, что становится голоден и бессилен, не пьет воды и изнемогает.
ISA|44|13|Плотник [выбрав дерево], протягивает по нему линию, остроконечным орудием делает на нем очертание, потом обделывает его резцом и округляет его, и выделывает из него образ человека красивого вида, чтобы поставить его в доме.
ISA|44|14|Он рубит себе кедры, берет сосну и дуб, которые выберет между деревьями в лесу, садит ясень, а дождь возращает его.
ISA|44|15|И это служит человеку топливом, и [часть] из этого употребляет он на то, чтобы ему было тепло, и разводит огонь, и печет хлеб. И из того же делает бога, и поклоняется ему, делает идола, и повергается перед ним.
ISA|44|16|Часть дерева сожигает в огне, другою частью варит мясо в пищу, жарит жаркое и ест досыта, а также греется и говорит: "хорошо, я согрелся; почувствовал огонь".
ISA|44|17|А из остатков от того делает бога, идола своего, поклоняется ему, повергается перед ним и молится ему, и говорит: "спаси меня, ибо ты бог мой".
ISA|44|18|Не знают и не разумеют они: Он закрыл глаза их, чтобы не видели, [и] сердца их, чтобы не разумели.
ISA|44|19|И не возьмет он этого к своему сердцу, и нет у него столько знания и смысла, чтобы сказать: "половину его я сжег в огне и на угольях его испек хлеб, изжарил мясо и съел; а из остатка его сделаю ли я мерзость? буду ли поклоняться куску дерева?"
ISA|44|20|Он гоняется за пылью; обманутое сердце ввело его в заблуждение, и он не может освободить души своей и сказать: "не обман ли в правой руке моей?"
ISA|44|21|Помни это, Иаков и Израиль, ибо ты раб Мой; Я образовал тебя: раб Мой ты, Израиль, не забывай Меня.
ISA|44|22|Изглажу беззакония твои, как туман, и грехи твои, как облако; обратись ко Мне, ибо Я искупил тебя.
ISA|44|23|Торжествуйте, небеса, ибо Господь соделал это. Восклицайте, глубины земли; шумите от радости, горы, лес и все деревья в нем; ибо искупил Господь Иакова и прославится в Израиле.
ISA|44|24|Так говорит Господь, искупивший тебя и образовавший тебя от утробы матерней: Я Господь, Который сотворил все, один распростер небеса и Своею силою разостлал землю,
ISA|44|25|Который делает ничтожными знамения лжепророков и обнаруживает безумие волшебников, мудрецов прогоняет назад и знание их делает глупостью,
ISA|44|26|Который утверждает слово раба Своего и приводит в исполнение изречение Своих посланников, Который говорит Иерусалиму: "ты будешь населен", и городам Иудиным: "вы будете построены, и развалины его Я восстановлю",
ISA|44|27|Который бездне говорит: "иссохни!" и реки твои Я иссушу,
ISA|44|28|Который говорит о Кире: пастырь Мой, и он исполнит всю волю Мою и скажет Иерусалиму: "ты будешь построен!" и храму: "ты будешь основан!"
ISA|45|1|Так говорит Господь помазаннику Своему Киру: Я держу тебя за правую руку, чтобы покорить тебе народы, и сниму поясы с чресл царей, чтоб отворялись для тебя двери, и ворота не затворялись;
ISA|45|2|Я пойду пред тобою и горы уровняю, медные двери сокрушу и запоры железные сломаю;
ISA|45|3|и отдам тебе хранимые во тьме сокровища и сокрытые богатства, дабы ты познал, что Я Господь, называющий тебя по имени, Бог Израилев.
ISA|45|4|Ради Иакова, раба Моего, и Израиля, избранного Моего, Я назвал тебя по имени, почтил тебя, хотя ты не знал Меня.
ISA|45|5|Я Господь, и нет иного; нет Бога кроме Меня; Я препоясал тебя, хотя ты не знал Меня,
ISA|45|6|дабы узнали от восхода солнца и от запада, что нет кроме Меня; Я Господь, и нет иного.
ISA|45|7|Я образую свет и творю тьму, делаю мир и произвожу бедствия; Я, Господь, делаю все это.
ISA|45|8|Кропите, небеса, свыше, и облака да проливают правду; да раскроется земля и приносит спасение, и да произрастает вместе правда. Я, Господь, творю это.
ISA|45|9|Горе тому, кто препирается с Создателем своим, черепок из черепков земных! Скажет ли глина горшечнику: "что ты делаешь?" и твое дело [скажет ли о тебе]: "у него нет рук?"
ISA|45|10|Горе тому, кто говорит отцу: "зачем ты произвел [меня] на свет?", а матери: "зачем ты родила [меня]?"
ISA|45|11|Так говорит Господь, Святый Израиля и Создатель его: вы спрашиваете Меня о будущем сыновей Моих и хотите Мне указывать в деле рук Моих?
ISA|45|12|Я создал землю и сотворил на ней человека; Я – Мои руки распростерли небеса, и всему воинству их дал закон Я.
ISA|45|13|Я воздвиг его в правде и уровняю все пути его. Он построит город Мой и отпустит пленных Моих, не за выкуп и не за дары, говорит Господь Саваоф.
ISA|45|14|Так говорит Господь: труды Египтян и торговля Ефиоплян, и Савейцы, люди рослые, к тебе перейдут и будут твоими; они последуют за тобою, в цепях придут и повергнутся пред тобою, и будут умолять тебя, [говоря]: у тебя только Бог, и нет иного Бога.
ISA|45|15|Истинно Ты Бог сокровенный, Бог Израилев, Спаситель.
ISA|45|16|Все они будут постыжены и посрамлены; вместе с ними со стыдом пойдут и все, делающие идолов.
ISA|45|17|Израиль же будет спасен спасением вечным в Господе; вы не будете постыжены и посрамлены во веки веков.
ISA|45|18|Ибо так говорит Господь, сотворивший небеса, Он, Бог, образовавший землю и создавший ее; Он утвердил ее, не напрасно сотворил ее; Он образовал ее для жительства: Я Господь, и нет иного.
ISA|45|19|Не тайно Я говорил, не в темном месте земли; не говорил Я племени Иакова: "напрасно ищете Меня". Я Господь, изрекающий правду, открывающий истину.
ISA|45|20|Соберитесь и придите, приблизьтесь все, уцелевшие из народов. Невежды те, которые носят деревянного своего идола и молятся богу, который не спасает.
ISA|45|21|Объявите и скажите, посоветовавшись между собою: кто возвестил это из древних времен, наперед сказал это? Не Я ли, Господь? и нет иного Бога кроме Меня, Бога праведного и спасающего нет кроме Меня.
ISA|45|22|Ко Мне обратитесь, и будете спасены, все концы земли, ибо я Бог, и нет иного.
ISA|45|23|Мною клянусь: из уст Моих исходит правда, слово неизменное, что предо Мною преклонится всякое колено, Мною будет клясться всякий язык.
ISA|45|24|Только у Господа, будут говорить о Мне, правда и сила; к Нему придут и устыдятся все, враждовавшие против Него.
ISA|45|25|Господом будет оправдано и прославлено все племя Израилево.
ISA|46|1|Пал Вил, низвергся Нево; истуканы их – на скоте и вьючных животных; ваша ноша сделалась бременем для усталых животных.
ISA|46|2|Низверглись, пали вместе; не могли защитить носивших, и сами пошли в плен.
ISA|46|3|Послушайте меня, дом Иаковлев и весь остаток дома Израилева, принятые [Мною] от чрева, носимые Мною от утробы [матерней]:
ISA|46|4|и до старости вашей Я тот же буду, и до седины вашей Я же буду носить [вас]; Я создал и буду носить, поддерживать и охранять вас.
ISA|46|5|Кому уподобите Меня, и [с кем] сравните, и с кем сличите, чтобы мы были сходны?
ISA|46|6|Высыпают золото из кошелька и весят серебро на весах, и нанимают серебряника, чтобы он сделал из него бога; кланяются ему и повергаются перед ним;
ISA|46|7|поднимают его на плечи, несут его и ставят его на свое место; он стоит, с места своего не двигается; кричат к нему, – он не отвечает, не спасает от беды.
ISA|46|8|Вспомните это и покажите себя мужами; примите это, отступники, к сердцу;
ISA|46|9|вспомните прежде бывшее, от [начала] века, ибо Я Бог, и нет иного Бога, и нет подобного Мне.
ISA|46|10|Я возвещаю от начала, что будет в конце, и от древних времен то, что еще не сделалось, говорю: Мой совет состоится, и все, что Мне угодно, Я сделаю.
ISA|46|11|Я воззвал орла от востока, из дальней страны, исполнителя определения Моего. Я сказал, и приведу это в исполнение; предначертал, и сделаю.
ISA|46|12|Послушайте Меня, жестокие сердцем, далекие от правды:
ISA|46|13|Я приблизил правду Мою, она не далеко, и спасение Мое не замедлит; и дам Сиону спасение, Израилю славу Мою.
ISA|47|1|Сойди и сядь на прах, девица, дочь Вавилона; сиди на земле: престола нет, дочь Халдеев, и вперед не будут называть тебя нежною и роскошною.
ISA|47|2|Возьми жернова и мели муку; сними покрывало твое, подбери подол, открой голени, переходи через реки:
ISA|47|3|откроется нагота твоя, и даже виден будет стыд твой. Совершу мщение и не пощажу никого.
ISA|47|4|Искупитель наш – Господь Саваоф имя Ему, Святый Израилев.
ISA|47|5|Сиди молча и уйди в темноту, дочь Халдеев: ибо вперед не будут называть тебя госпожею царств.
ISA|47|6|Я прогневался на народ Мой, уничижил наследие Мое и предал их в руки твои; [а] ты не оказала им милосердия, на старца налагала крайне тяжкое иго твое.
ISA|47|7|И ты говорила: "вечно буду госпожею", а не представляла того в уме твоем, не помышляла, что будет после.
ISA|47|8|Но ныне выслушай это, изнеженная, живущая беспечно, говорящая в сердце своем: "я, – и другой подобной мне нет; не буду сидеть вдовою и не буду знать потери детей".
ISA|47|9|Но внезапно, в один день, придет к тебе то и другое, потеря детей и вдовство; в полной мере придут они на тебя, несмотря на множество чародейств твоих и на великую силу волшебств твоих.
ISA|47|10|Ибо ты надеялась на злодейство твое, говорила: "никто не видит меня". Мудрость твоя и знание твое – они сбили тебя с пути; и ты говорила в сердце твоем: "я, и никто кроме меня".
ISA|47|11|И придет на тебя бедствие: ты не узнаешь, откуда оно поднимется; и нападет на тебя беда, которой ты не в силах будешь отвратить, и внезапно придет на тебя пагуба, о которой ты и не думаешь.
ISA|47|12|Оставайся же с твоими волшебствами и со множеством чародейств твоих, которыми ты занималась от юности твоей: может быть, пособишь себе, может быть, устоишь.
ISA|47|13|Ты утомлена множеством советов твоих; пусть же выступят наблюдатели небес и звездочеты и предвещатели по новолуниям, и спасут тебя от того, что должно приключиться тебе.
ISA|47|14|Вот они, как солома: огонь сожег их, – не избавили души своей от пламени; не осталось угля, чтобы погреться, ни огня, чтобы посидеть перед ним.
ISA|47|15|Такими стали для тебя те, с которыми ты трудилась, с которыми вела торговлю от юности твоей. Каждый побрел в свою сторону; никто не спасает тебя.
ISA|48|1|Слушайте это, дом Иакова, называющиеся именем Израиля и происшедшие от источника Иудина, клянущиеся именем Господа и исповедающие Бога Израилева, хотя не по истине и не по правде.
ISA|48|2|Ибо они называют себя [происходящими] от святого города и опираются на Бога Израилева; Господь Саваоф – имя Ему.
ISA|48|3|Прежнее Я задолго объявлял; из Моих уст выходило оно, и Я возвещал это и внезапно делал, и все сбывалось.
ISA|48|4|Я знал, что ты упорен, и что в шее твоей жилы железные, и лоб твой – медный;
ISA|48|5|поэтому и объявлял тебе задолго, прежде нежели это приходило, и предъявлял тебе, чтобы ты не сказал: "идол мой сделал это, и истукан мой и изваянный мой повелел этому быть".
ISA|48|6|Ты слышал, – посмотри на все это! и неужели вы не признаете этого? А ныне Я возвещаю тебе новое и сокровенное, и ты не знал этого.
ISA|48|7|Оно произошло ныне, а не задолго и не за день, и ты не слыхал о том, чтобы ты не сказал: "вот! я знал это".
ISA|48|8|Ты и не слыхал и не знал об этом, и ухо твое не было прежде открыто; ибо Я знал, что ты поступишь вероломно, и от самого чрева [матернего] ты прозван отступником.
ISA|48|9|Ради имени Моего отлагал гнев Мой, и ради славы Моей удерживал Себя от истребления тебя.
ISA|48|10|Вот, Я расплавил тебя, но не как серебро; испытал тебя в горниле страдания.
ISA|48|11|Ради Себя, ради Себя Самого делаю это, – ибо какое было бы нарекание [на имя Мое]! славы Моей не дам иному.
ISA|48|12|Послушай Меня, Иаков и Израиль, призванный Мой: Я тот же, Я первый и Я последний.
ISA|48|13|Моя рука основала землю, и Моя десница распростерла небеса; призову их, и они предстанут вместе.
ISA|48|14|Соберитесь все и слушайте: кто между ними предсказал это? Господь возлюбил его, и он исполнит волю Его над Вавилоном и явит мышцу Его над Халдеями.
ISA|48|15|Я, Я сказал, и призвал его; Я привел его, и путь его будет благоуспешен.
ISA|48|16|Приступите ко Мне, слушайте это: Я и сначала говорил не тайно; с того времени, как это происходит, Я был там; и ныне послал Меня Господь Бог и Дух Его.
ISA|48|17|Так говорит Господь, Искупитель твой, Святый Израилев: Я Господь, Бог твой, научающий тебя полезному, ведущий тебя по тому пути, по которому должно тебе идти.
ISA|48|18|О, если бы ты внимал заповедям Моим! тогда мир твой был бы как река, и правда твоя – как волны морские.
ISA|48|19|И семя твое было бы как песок, и происходящие из чресл твоих – как песчинки: не изгладилось бы, не истребилось бы имя его предо Мною.
ISA|48|20|Выходите из Вавилона, бегите от Халдеев, со гласом радости возвещайте и проповедуйте это, распространяйте эту весть до пределов земли; говорите: "Господь искупил раба Своего Иакова".
ISA|48|21|И не жаждут они в пустынях, чрез которые Он ведет их: Он источает им воду из камня; рассекает скалу, и льются воды.
ISA|48|22|Нечестивым же нет мира, говорит Господь.
ISA|49|1|Слушайте Меня, острова, и внимайте, народы дальние: Господь призвал Меня от чрева, от утробы матери Моей называл имя Мое;
ISA|49|2|и соделал уста Мои как острый меч; тенью руки Своей покрывал Меня, и соделал Меня стрелою изостренною; в колчане Своем хранил Меня;
ISA|49|3|и сказал Мне: Ты раб Мой, Израиль, в Тебе Я прославлюсь.
ISA|49|4|А Я сказал: напрасно Я трудился, ни на что и вотще истощал силу Свою. Но Мое право у Господа, и награда Моя у Бога Моего.
ISA|49|5|И ныне говорит Господь, образовавший Меня от чрева в раба Себе, чтобы обратить к Нему Иакова и чтобы Израиль собрался к Нему; Я почтен в очах Господа, и Бог Мой – сила Моя.
ISA|49|6|И Он сказал: мало того, что Ты будешь рабом Моим для восстановления колен Иаковлевых и для возвращения остатков Израиля, но Я сделаю Тебя светом народов, чтобы спасение Мое простерлось до концов земли.
ISA|49|7|Так говорит Господь, Искупитель Израиля, Святый Его, презираемому всеми, поносимому народом, рабу властелинов: цари увидят, и встанут; князья поклонятся ради Господа, Который верен, ради Святаго Израилева, Который избрал Тебя.
ISA|49|8|Так говорит Господь: во время благоприятное Я услышал Тебя, и в день спасения помог Тебе; и Я буду охранять Тебя, и сделаю Тебя заветом народа, чтобы восстановить землю, чтобы возвратить наследникам наследия опустошенные,
ISA|49|9|сказать узникам: "выходите", и тем, которые во тьме: "покажитесь". Они при дорогах будут пасти, и по всем холмам будут пажити их;
ISA|49|10|не будут терпеть голода и жажды, и не поразит их зной и солнце; ибо Милующий их будет вести их и приведет их к источникам вод.
ISA|49|11|И все горы Мои сделаю путем, и дороги Мои будут подняты.
ISA|49|12|Вот, одни придут издалека; и вот, одни от севера и моря, а другие из земли Синим.
ISA|49|13|Радуйтесь, небеса, и веселись, земля, и восклицайте, горы, от радости; ибо утешил Господь народ Свой и помиловал страдальцев Своих.
ISA|49|14|А Сион говорил: "оставил меня Господь, и Бог мой забыл меня!"
ISA|49|15|Забудет ли женщина грудное дитя свое, чтобы не пожалеть сына чрева своего? но если бы и она забыла, то Я не забуду тебя.
ISA|49|16|Вот, Я начертал тебя на дланях [Моих]; стены твои всегда предо Мною.
ISA|49|17|Сыновья твои поспешат [к тебе], а разорители и опустошители твои уйдут от тебя.
ISA|49|18|Возведи очи твои и посмотри вокруг, – все они собираются, идут к тебе. Живу Я! говорит Господь, – всеми ими ты облечешься, как убранством, и нарядишься ими, как невеста.
ISA|49|19|Ибо развалины твои и пустыни твои, и разоренная земля твоя будут теперь слишком тесны для жителей, и поглощавшие тебя удалятся от тебя.
ISA|49|20|Дети, которые будут у тебя после потери прежних, будут говорить вслух тебе: "тесно для меня место; уступи мне, чтобы я мог жить".
ISA|49|21|И ты скажешь в сердце твоем: кто мне родил их? я была бездетна и бесплодна, отведена в плен и удалена; кто же возрастил их? вот, я оставалась одинокою; где же они были?
ISA|49|22|Так говорит Господь Бог: вот, Я подниму руку Мою к народам, и выставлю знамя Мое племенам, и принесут сыновей твоих на руках и дочерей твоих на плечах.
ISA|49|23|И будут цари питателями твоими, и царицы их кормилицами твоими; лицом до земли будут кланяться тебе и лизать прах ног твоих, и узнаешь, что Я Господь, что надеющиеся на Меня не постыдятся.
ISA|49|24|Может ли быть отнята у сильного добыча, и могут ли быть отняты у победителя взятые в плен?
ISA|49|25|Да! так говорит Господь: и плененные сильным будут отняты, и добыча тирана будет избавлена; потому что Я буду состязаться с противниками твоими и сыновей твоих Я спасу;
ISA|49|26|и притеснителей твоих накормлю собственною их плотью, и они будут упоены кровью своею, как молодым вином; и всякая плоть узнает, что Я Господь, Спаситель твой и Искупитель твой, Сильный Иаковлев.
ISA|50|1|Так говорит Господь: где разводное письмо вашей матери, с которым Я отпустил ее? или которому из Моих заимодавцев Я продал вас? Вот, вы проданы за грехи ваши, и за преступления ваши отпущена мать ваша.
ISA|50|2|Почему, когда Я приходил, никого не было, и когда Я звал, никто не отвечал? Разве рука Моя коротка стала для того, чтобы избавлять, или нет силы во Мне, чтобы спасать? Вот, прещением Моим Я иссушаю море, превращаю реки в пустыню; рыбы в них гниют от недостатка воды и умирают от жажды.
ISA|50|3|Я облекаю небеса мраком, и вретище делаю покровом их.
ISA|50|4|Господь Бог дал Мне язык мудрых, чтобы Я мог словом подкреплять изнемогающего; каждое утро Он пробуждает, пробуждает ухо Мое, чтобы Я слушал, подобно учащимся.
ISA|50|5|Господь Бог открыл Мне ухо, и Я не воспротивился, не отступил назад.
ISA|50|6|Я предал хребет Мой биющим и ланиты Мои поражающим; лица Моего не закрывал от поруганий и оплевания.
ISA|50|7|И Господь Бог помогает Мне: поэтому Я не стыжусь, поэтому Я держу лице Мое, как кремень, и знаю, что не останусь в стыде.
ISA|50|8|Близок оправдывающий Меня: кто хочет состязаться со Мною? станем вместе. Кто хочет судиться со Мною? пусть подойдет ко Мне.
ISA|50|9|Вот, Господь Бог помогает Мне: кто осудит Меня? Вот, все они, как одежда, обветшают; моль съест их.
ISA|50|10|Кто из вас боится Господа, слушается гласа Раба Его? Кто ходит во мраке, без света, да уповает на имя Господа и да утверждается в Боге своем.
ISA|50|11|Вот, все вы, которые возжигаете огонь, вооруженные зажигательными стрелами, – идите в пламень огня вашего и стрел, раскаленных вами! Это будет вам от руки Моей; в мучении умрете.
ISA|51|1|Послушайте Меня, стремящиеся к правде, ищущие Господа! Взгляните на скалу, из которой вы иссечены, в глубину рва, из которого вы извлечены.
ISA|51|2|Посмотрите на Авраама, отца вашего, и на Сарру, родившую вас: ибо Я призвал его одного и благословил его, и размножил его.
ISA|51|3|Так, Господь утешит Сион, утешит все развалины его и сделает пустыни его, как рай, и степь его, как сад Господа; радость и веселие будет в нем, славословие и песнопение.
ISA|51|4|Послушайте Меня, народ Мой, и племя Мое, приклоните ухо ко Мне! ибо от Меня произойдет закон, и суд Мой поставлю во свет для народов.
ISA|51|5|Правда Моя близка; спасение Мое восходит, и мышца Моя будет судить народы; острова будут уповать на Меня и надеяться на мышцу Мою.
ISA|51|6|Поднимите глаза ваши к небесам, и посмотрите на землю вниз: ибо небеса исчезнут, как дым, и земля обветшает, как одежда, и жители ее также вымрут; а Мое спасение пребудет вечным, и правда Моя не престанет.
ISA|51|7|Послушайте Меня, знающие правду, народ, у которого в сердце закон Мой! Не бойтесь поношения от людей, и злословия их не страшитесь.
ISA|51|8|Ибо, как одежду, съест их моль и, как волну, съест их червь; а правда Моя пребудет вовек, и спасение Мое – в роды родов.
ISA|51|9|Восстань, восстань, облекись крепостью, мышца Господня! Восстань, как в дни древние, в роды давние! Не ты ли сразила Раава, поразила крокодила?
ISA|51|10|Не ты ли иссушила море, воды великой бездны, превратила глубины моря в дорогу, чтобы прошли искупленные?
ISA|51|11|И возвратятся избавленные Господом и придут на Сион с пением, и радость вечная над головою их; они найдут радость и веселье: печаль и вздохи удалятся.
ISA|51|12|Я, Я Сам – Утешитель ваш. Кто ты, что боишься человека, который умирает, и сына человеческого, который то же, что трава,
ISA|51|13|и забываешь Господа, Творца своего, распростершего небеса и основавшего землю; и непрестанно, всякий день страшишься ярости притеснителя, как бы он готов был истребить? Но где ярость притеснителя?
ISA|51|14|Скоро освобожден будет пленный, и не умрет в яме и не будет нуждаться в хлебе.
ISA|51|15|Я Господь, Бог твой, возмущающий море, так что волны его ревут: Господь Саваоф – имя Его.
ISA|51|16|И Я вложу слова Мои в уста твои, и тенью руки Моей покрою тебя, чтобы устроить небеса и утвердить землю и сказать Сиону: "ты Мой народ".
ISA|51|17|Воспряни, воспряни, восстань, Иерусалим, ты, который из руки Господа выпил чашу ярости Его, выпил до дна чашу опьянения, осушил.
ISA|51|18|Некому было вести его из всех сыновей, рожденных им, и некому было поддержать его за руку из всех сыновей, [которых] он возрастил.
ISA|51|19|Тебя постигли два [бедствия], кто пожалеет о тебе? – опустошение и истребление, голод и меч: кем я утешу тебя?
ISA|51|20|Сыновья твои изнемогли, лежат по углам всех улиц, как серна в тенетах, исполненные гнева Господа, прещения Бога твоего.
ISA|51|21|Итак выслушай это, страдалец и опьяневший, но не от вина.
ISA|51|22|Так говорит Господь твой, Господь и Бог твой, отмщающий за Свой народ: вот, Я беру из руки твоей чашу опьянения, дрожжи из чаши ярости Моей: ты не будешь уже пить их,
ISA|51|23|и подам ее в руки мучителям твоим, которые говорили тебе: "пади ниц, чтобы нам пройти по тебе"; и ты хребет твой делал как бы землею и улицею для проходящих.
ISA|52|1|Восстань, восстань, облекись в силу твою, Сион! Облекись в одежды величия твоего, Иерусалим, город святый! ибо уже не будет более входить в тебя необрезанный и нечистый.
ISA|52|2|Отряси с себя прах; встань, пленный Иерусалим! сними цепи с шеи твоей, пленная дочь Сиона!
ISA|52|3|ибо так говорит Господь: за ничто были вы проданы, и без серебра будете выкуплены;
ISA|52|4|ибо так говорит Господь Бог: народ Мой ходил прежде в Египет, чтобы там пожить, и Ассур теснил его ни за что.
ISA|52|5|И теперь что у Меня здесь? говорит Господь; народ Мой взят даром, властители их неистовствуют, говорит Господь, и постоянно, всякий день имя Мое бесславится.
ISA|52|6|Поэтому народ Мой узнает имя Мое; поэтому [узнает] в тот день, что Я тот же, Который сказал: "вот Я!"
ISA|52|7|Как прекрасны на горах ноги благовестника, возвещающего мир, благовествующего радость, проповедующего спасение, говорящего Сиону: "воцарился Бог твой!"
ISA|52|8|Голос сторожей твоих – они возвысили голос, и все вместе ликуют, ибо своими глазами видят, что Господь возвращается в Сион.
ISA|52|9|Торжествуйте, пойте вместе, развалины Иерусалима, ибо утешил Господь народ Свой, искупил Иерусалим.
ISA|52|10|Обнажил Господь святую мышцу Свою пред глазами всех народов; и все концы земли увидят спасение Бога нашего.
ISA|52|11|Идите, идите, выходите оттуда; не касайтесь нечистого; выходите из среды его, очистите себя, носящие сосуды Господни!
ISA|52|12|ибо вы выйдете неторопливо, и не побежите; потому что впереди вас пойдет Господь, и Бог Израилев будет стражем позади вас.
ISA|52|13|Вот, раб Мой будет благоуспешен, возвысится и вознесется, и возвеличится.
ISA|52|14|Как многие изумлялись, [смотря] на Тебя, – столько был обезображен паче всякого человека лик Его, и вид Его – паче сынов человеческих!
ISA|52|15|Так многие народы приведет Он в изумление; цари закроют пред Ним уста свои, ибо они увидят то, о чем не было говорено им, и узнают то, чего не слыхали.
ISA|53|1|Кто поверил слышанному от нас, и кому открылась мышца Господня?
ISA|53|2|Ибо Он взошел пред Ним, как отпрыск и как росток из сухой земли; нет в Нем ни вида, ни величия; и мы видели Его, и не было в Нем вида, который привлекал бы нас к Нему.
ISA|53|3|Он был презрен и умален пред людьми, муж скорбей и изведавший болезни, и мы отвращали от Него лице свое; Он был презираем, и мы ни во что ставили Его.
ISA|53|4|Но Он взял на Себя наши немощи и понес наши болезни; а мы думали, [что] Он был поражаем, наказуем и уничижен Богом.
ISA|53|5|Но Он изъязвлен был за грехи наши и мучим за беззакония наши; наказание мира нашего [было] на Нем, и ранами Его мы исцелились.
ISA|53|6|Все мы блуждали, как овцы, совратились каждый на свою дорогу: и Господь возложил на Него грехи всех нас.
ISA|53|7|Он истязуем был, но страдал добровольно и не открывал уст Своих; как овца, веден был Он на заклание, и как агнец пред стригущим его безгласен, так Он не отверзал уст Своих.
ISA|53|8|От уз и суда Он был взят; но род Его кто изъяснит? ибо Он отторгнут от земли живых; за преступления народа Моего претерпел казнь.
ISA|53|9|Ему назначали гроб со злодеями, но Он погребен у богатого, потому что не сделал греха, и не было лжи в устах Его.
ISA|53|10|Но Господу угодно было поразить Его, и Он предал Его мучению; когда же душа Его принесет жертву умилостивления, Он узрит потомство долговечное, и воля Господня благоуспешно будет исполняться рукою Его.
ISA|53|11|На подвиг души Своей Он будет смотреть с довольством; чрез познание Его Он, Праведник, Раб Мой, оправдает многих и грехи их на Себе понесет.
ISA|53|12|Посему Я дам Ему часть между великими, и с сильными будет делить добычу, за то, что предал душу Свою на смерть, и к злодеям причтен был, тогда как Он понес на Себе грех многих и за преступников сделался ходатаем.
ISA|54|1|Возвеселись, неплодная, нерождающая; воскликни и возгласи, немучившаяся родами; потому что у оставленной гораздо более детей, нежели у имеющей мужа, говорит Господь.
ISA|54|2|Распространи место шатра твоего, расширь покровы жилищ твоих; не стесняйся, пусти длиннее верви твои и утверди колья твои;
ISA|54|3|ибо ты распространишься направо и налево, и потомство твое завладеет народами и населит опустошенные города.
ISA|54|4|Не бойся, ибо не будешь постыжена; не смущайся, ибо не будешь в поругании: ты забудешь посрамление юности твоей и не будешь более вспоминать о бесславии вдовства твоего.
ISA|54|5|Ибо твой Творец есть супруг твой; Господь Саваоф – имя Его; и Искупитель твой – Святый Израилев: Богом всей земли назовется Он.
ISA|54|6|Ибо как жену, оставленную и скорбящую духом, призывает тебя Господь, и [как] жену юности, которая была отвержена, говорит Бог твой.
ISA|54|7|На малое время Я оставил тебя, но с великою милостью восприму тебя.
ISA|54|8|В жару гнева Я сокрыл от тебя лице Мое на время, но вечною милостью помилую тебя, говорит Искупитель твой, Господь.
ISA|54|9|Ибо это для Меня, как воды Ноя: как Я поклялся, что воды Ноя не придут более на землю, так поклялся не гневаться на тебя и не укорять тебя.
ISA|54|10|Горы сдвинутся и холмы поколеблются, – а милость Моя не отступит от тебя, и завет мира Моего не поколеблется, говорит милующий тебя Господь.
ISA|54|11|Бедная, бросаемая бурею, безутешная! Вот, Я положу камни твои на рубине и сделаю основание твое из сапфиров;
ISA|54|12|и сделаю окна твои из рубинов и ворота твои – из жемчужин, и всю ограду твою – из драгоценных камней.
ISA|54|13|И все сыновья твои будут научены Господом, и великий мир будет у сыновей твоих.
ISA|54|14|Ты утвердишься правдою, будешь далека от угнетения, ибо тебе бояться нечего, и от ужаса, ибо он не приблизится к тебе.
ISA|54|15|Вот, будут вооружаться [против тебя], но не от Меня; кто бы ни вооружился против тебя, падет.
ISA|54|16|Вот, Я сотворил кузнеца, который раздувает угли в огне и производит орудие для своего дела, – и Я творю губителя для истребления.
ISA|54|17|Ни одно орудие, сделанное против тебя, не будет успешно; и всякий язык, который будет состязаться с тобою на суде, – ты обвинишь. Это есть наследие рабов Господа, оправдание их от Меня, говорит Господь.
ISA|55|1|Жаждущие! идите все к водам; даже и вы, у которых нет серебра, идите, покупайте и ешьте; идите, покупайте без серебра и без платы вино и молоко.
ISA|55|2|Для чего вам отвешивать серебро за то, что не хлеб, и трудовое свое за то, что не насыщает? Послушайте Меня внимательно и вкушайте благо, и душа ваша да насладится туком.
ISA|55|3|Приклоните ухо ваше и придите ко Мне: послушайте, и жива будет душа ваша, – и дам вам завет вечный, неизменные милости, [обещанные] Давиду.
ISA|55|4|Вот, Я дал Его свидетелем для народов, вождем и наставником народам.
ISA|55|5|Вот, ты призовешь народ, которого ты не знал, и народы, которые тебя не знали, поспешат к тебе ради Господа Бога твоего и ради Святаго Израилева, ибо Он прославил тебя.
ISA|55|6|Ищите Господа, когда можно найти Его; призывайте Его, когда Он близко.
ISA|55|7|Да оставит нечестивый путь свой и беззаконник – помыслы свои, и да обратится к Господу, и Он помилует его, и к Богу нашему, ибо Он многомилостив.
ISA|55|8|Мои мысли – не ваши мысли, ни ваши пути – пути Мои, говорит Господь.
ISA|55|9|Но как небо выше земли, так пути Мои выше путей ваших, и мысли Мои выше мыслей ваших.
ISA|55|10|Как дождь и снег нисходит с неба и туда не возвращается, но напояет землю и делает ее способною рождать и произращать, чтобы она давала семя тому, кто сеет, и хлеб тому, кто ест, –
ISA|55|11|так и слово Мое, которое исходит из уст Моих, – оно не возвращается ко Мне тщетным, но исполняет то, что Мне угодно, и совершает то, для чего Я послал его.
ISA|55|12|Итак вы выйдете с веселием и будете провожаемы с миром; горы и холмы будут петь пред вами песнь, и все дерева в поле рукоплескать вам.
ISA|55|13|Вместо терновника вырастет кипарис; вместо крапивы возрастет мирт; и это будет во славу Господа, в знамение вечное, несокрушимое.
ISA|56|1|Так говорит Господь: сохраняйте суд и делайте правду; ибо близко спасение Мое и откровение правды Моей.
ISA|56|2|Блажен муж, который делает это, и сын человеческий, который крепко держится этого, который хранит субботу от осквернения и оберегает руку свою, чтобы не сделать никакого зла.
ISA|56|3|Да не говорит сын иноплеменника, присоединившийся к Господу: "Господь совсем отделил меня от Своего народа", и да не говорит евнух: "вот я сухое дерево".
ISA|56|4|Ибо Господь так говорит об евнухах: которые хранят Мои субботы и избирают угодное Мне, и крепко держатся завета Моего, –
ISA|56|5|тем дам Я в доме Моем и в стенах Моих место и имя лучшее, нежели сыновьям и дочерям; дам им вечное имя, которое не истребится.
ISA|56|6|И сыновей иноплеменников, присоединившихся к Господу, чтобы служить Ему и любить имя Господа, быть рабами Его, всех, хранящих субботу от осквернения ее и твердо держащихся завета Моего,
ISA|56|7|Я приведу на святую гору Мою и обрадую их в Моем доме молитвы; всесожжения их и жертвы их [будут] благоприятны на жертвеннике Моем, ибо дом Мой назовется домом молитвы для всех народов.
ISA|56|8|Господь Бог, собирающий рассеянных Израильтян, говорит: к собранным у него Я буду еще собирать других.
ISA|56|9|Все звери полевые, все звери лесные! идите есть.
ISA|56|10|Стражи их слепы все и невежды: все они немые псы, не могущие лаять, бредящие лежа, любящие спать.
ISA|56|11|И это псы, жадные душею, не знающие сытости; и это пастыри бессмысленные: все смотрят на свою дорогу, каждый до последнего, на свою корысть;
ISA|56|12|приходите, [говорят], я достану вина, и мы напьемся сикеры; и завтра то же будет, что сегодня, да еще и больше.
ISA|57|1|Праведник умирает, и никто не принимает этого к сердцу; и мужи благочестивые восхищаются [от земли], и никто не помыслит, что праведник восхищается от зла.
ISA|57|2|Он отходит к миру; ходящие прямым путем будут покоиться на ложах своих.
ISA|57|3|Но приблизьтесь сюда вы, сыновья чародейки, семя прелюбодея и блудницы!
ISA|57|4|Над кем вы глумитесь? против кого расширяете рот, высовываете язык? не дети ли вы преступления, семя лжи,
ISA|57|5|разжигаемые похотью к идолам под каждым ветвистым деревом, заколающие детей при ручьях, между расселинами скал?
ISA|57|6|В гладких камнях ручьев доля твоя; они, они жребий твой; им ты делаешь возлияние и приносишь жертвы: могу ли Я быть доволен этим?
ISA|57|7|На высокой и выдающейся горе ты ставишь ложе твое и туда восходишь приносить жертву.
ISA|57|8|За дверью также и за косяками ставишь памяти твои; ибо, отвратившись от Меня, ты обнажаешься и восходишь; распространяешь ложе твое и договариваешься с теми из них, с которыми любишь лежать, высматриваешь место.
ISA|57|9|Ты ходила также к царю с благовонною мастью и умножила масти твои, и далеко посылала послов твоих, и унижалась до преисподней.
ISA|57|10|От долгого пути твоего утомлялась, но не говорила: "надежда потеряна!"; все еще находила живость в руке твоей, и потому не чувствовала ослабления.
ISA|57|11|Кого же ты испугалась и устрашилась, что сделалась неверною и Меня перестала помнить и хранить в твоем сердце? не от того ли, что Я молчал, и притом долго, ты перестала бояться Меня?
ISA|57|12|Я покажу правду твою и дела твои, – и они будут не в пользу тебе.
ISA|57|13|Когда ты будешь вопить, спасет ли тебя сборище твое? – всех их унесет ветер, развеет дуновение; а надеющийся на Меня наследует землю и будет владеть святою горою Моею.
ISA|57|14|И сказал: поднимайте, поднимайте, ровняйте путь, убирайте преграду с пути народа Моего.
ISA|57|15|Ибо так говорит Высокий и Превознесенный, вечно Живущий, – Святый имя Его: Я живу на высоте [небес] и во святилище, и также с сокрушенными и смиренными духом, чтобы оживлять дух смиренных и оживлять сердца сокрушенных.
ISA|57|16|Ибо не вечно буду Я вести тяжбу и не до конца гневаться; иначе изнеможет предо Мною дух и всякое дыхание, Мною сотворенное.
ISA|57|17|За грех корыстолюбия его Я гневался и поражал его, скрывал лице и негодовал; но он, отвратившись, пошел по пути своего сердца.
ISA|57|18|Я видел пути его, и исцелю его, и буду водить его и утешать его и сетующих его.
ISA|57|19|Я исполню слово: мир, мир дальнему и ближнему, говорит Господь, и исцелю его.
ISA|57|20|А нечестивые – как море взволнованное, которое не может успокоиться и которого воды выбрасывают ил и грязь.
ISA|57|21|Нет мира нечестивым, говорит Бог мой.
ISA|58|1|Взывай громко, не удерживайся; возвысь голос твой, подобно трубе, и укажи народу Моему на беззакония его, и дому Иаковлеву – на грехи его.
ISA|58|2|Они каждый день ищут Меня и хотят знать пути Мои, как бы народ, поступающий праведно и не оставляющий законов Бога своего; они вопрошают Меня о судах правды, желают приближения к Богу:
ISA|58|3|"Почему мы постимся, а Ты не видишь? смиряем души свои, а Ты не знаешь?" – Вот, в день поста вашего вы исполняете волю вашу и требуете тяжких трудов от других.
ISA|58|4|Вот, вы поститесь для ссор и распрей и для того, чтобы дерзкою рукою бить других; вы не поститесь в это время так, чтобы голос ваш был услышан на высоте.
ISA|58|5|Таков ли тот пост, который Я избрал, день, в который томит человек душу свою, когда гнет голову свою, как тростник, и подстилает под себя рубище и пепел? Это ли назовешь постом и днем, угодным Господу?
ISA|58|6|Вот пост, который Я избрал: разреши оковы неправды, развяжи узы ярма, и угнетенных отпусти на свободу, и расторгни всякое ярмо;
ISA|58|7|раздели с голодным хлеб твой, и скитающихся бедных введи в дом; когда увидишь нагого, одень его, и от единокровного твоего не укрывайся.
ISA|58|8|Тогда откроется, как заря, свет твой, и исцеление твое скоро возрастет, и правда твоя пойдет пред тобою, и слава Господня будет сопровождать тебя.
ISA|58|9|Тогда ты воззовешь, и Господь услышит; возопиешь, и Он скажет: "вот Я!" Когда ты удалишь из среды твоей ярмо, перестанешь поднимать перст и говорить оскорбительное,
ISA|58|10|и отдашь голодному душу твою и напитаешь душу страдальца: тогда свет твой взойдет во тьме, и мрак твой [будет] как полдень;
ISA|58|11|и будет Господь вождем твоим всегда, и во время засухи будет насыщать душу твою и утучнять кости твои, и ты будешь, как напоенный водою сад и как источник, которого воды никогда не иссякают.
ISA|58|12|И застроятся [потомками] твоими пустыни вековые: ты восстановишь основания многих поколений, и будут называть тебя восстановителем развалин, возобновителем путей для населения.
ISA|58|13|Если ты удержишь ногу твою ради субботы от исполнения прихотей твоих во святый день Мой, и будешь называть субботу отрадою, святым днем Господним, чествуемым, и почтишь ее тем, что не будешь заниматься обычными твоими делами, угождать твоей прихоти и пустословить, –
ISA|58|14|то будешь иметь радость в Господе, и Я возведу тебя на высоты земли и дам вкусить тебе наследие Иакова, отца твоего: уста Господни изрекли это.
ISA|59|1|Вот, рука Господа не сократилась на то, чтобы спасать, и ухо Его не отяжелело для того, чтобы слышать.
ISA|59|2|Но беззакония ваши произвели разделение между вами и Богом вашим, и грехи ваши отвращают лице [Его] от вас, чтобы не слышать.
ISA|59|3|Ибо руки ваши осквернены кровью и персты ваши – беззаконием; уста ваши говорят ложь, язык ваш произносит неправду.
ISA|59|4|Никто не возвышает голоса за правду, и никто не вступается за истину; надеются на пустое и говорят ложь, зачинают зло и рождают злодейство;
ISA|59|5|высиживают змеиные яйца и ткут паутину; кто поест яиц их, – умрет, а если раздавит, – выползет ехидна.
ISA|59|6|Паутины их для одежды негодны, и они не покроются своим произведением; дела их – дела неправедные, и насилие в руках их.
ISA|59|7|Ноги их бегут ко злу, и они спешат на пролитие невинной крови; мысли их – мысли нечестивые; опустошение и гибель на стезях их.
ISA|59|8|Пути мира они не знают, и нет суда на стезях их; пути их искривлены, и никто, идущий по ним, не знает мира.
ISA|59|9|Потому–то и далек от нас суд, и правосудие не достигает до нас; ждем света, и вот тьма, – озарения, и ходим во мраке.
ISA|59|10|Осязаем, как слепые стену, и, как без глаз, ходим ощупью; спотыкаемся в полдень, как в сумерки, между живыми – как мертвые.
ISA|59|11|Все мы ревем, как медведи, и стонем, как голуби; ожидаем суда, и нет [его], – спасения, но оно далеко от нас.
ISA|59|12|Ибо преступления наши многочисленны пред Тобою, и грехи наши свидетельствуют против нас; ибо преступления наши с нами, и беззакония наши мы знаем.
ISA|59|13|Мы изменили и солгали пред Господом, и отступили от Бога нашего; говорили клевету и измену, зачинали и рождали из сердца лживые слова.
ISA|59|14|И суд отступил назад, и правда стала вдали, ибо истина преткнулась на площади, и честность не может войти.
ISA|59|15|И не стало истины, и удаляющийся от зла подвергается оскорблению. И Господь увидел это, и противно было очам Его, что нет суда.
ISA|59|16|И видел, что нет человека, и дивился, что нет заступника; и помогла Ему мышца Его, и правда Его поддержала Его.
ISA|59|17|И Он возложил на Себя правду, как броню, и шлем спасения на главу Свою; и облекся в ризу мщения, как в одежду, и покрыл Себя ревностью, как плащом.
ISA|59|18|По мере возмездия, по этой мере Он воздаст противникам Своим – яростью, врагам Своим – местью, островам воздаст должное.
ISA|59|19|И убоятся имени Господа на западе и славы Его – на восходе солнца. Если враг придет как река, дуновение Господа прогонит его.
ISA|59|20|И придет Искупитель Сиона и [сынов] Иакова, обратившихся от нечестия, говорит Господь.
ISA|59|21|И вот завет Мой с ними, говорит Господь: Дух Мой, Который на тебе, и слова Мои, которые вложил Я в уста твои, не отступят от уст твоих и от уст потомства твоего, и от уст потомков потомства твоего, говорит Господь, отныне и до века.
ISA|60|1|Восстань, светись, [Иерусалим], ибо пришел свет твой, и слава Господня взошла над тобою.
ISA|60|2|Ибо вот, тьма покроет землю, и мрак – народы; а над тобою воссияет Господь, и слава Его явится над тобою.
ISA|60|3|И придут народы к свету твоему, и цари – к восходящему над тобою сиянию.
ISA|60|4|Возведи очи твои и посмотри вокруг: все они собираются, идут к тебе; сыновья твои издалека идут и дочерей твоих на руках несут.
ISA|60|5|Тогда увидишь, и возрадуешься, и затрепещет и расширится сердце твое, потому что богатство моря обратится к тебе, достояние народов придет к тебе.
ISA|60|6|Множество верблюдов покроет тебя – дромадеры из Мадиама и Ефы; все они из Савы придут, принесут золото и ладан и возвестят славу Господа.
ISA|60|7|Все овцы Кидарские будут собраны к тебе; овны Неваиофские послужат тебе: взойдут на алтарь Мой жертвою благоугодною, и Я прославлю дом славы Моей.
ISA|60|8|Кто это летят, как облака, и как голуби – к голубятням своим?
ISA|60|9|Так, Меня ждут острова и впереди их – корабли Фарсисские, чтобы перевезти сынов твоих издалека и с ними серебро их и золото их, во имя Господа Бога твоего и Святаго Израилева, потому что Он прославил тебя.
ISA|60|10|Тогда сыновья иноземцев будут строить стены твои, и цари их – служить тебе; ибо во гневе Моем Я поражал тебя, но в благоволении Моем буду милостив к тебе.
ISA|60|11|И будут всегда отверсты врата твои, не будут затворяться ни днем ни ночью, чтобы приносимо было к тебе достояние народов и приводимы были цари их.
ISA|60|12|Ибо народ и царства, которые не захотят служить тебе, – погибнут, и такие народы совершенно истребятся.
ISA|60|13|Слава Ливана придет к тебе, кипарис и певг и вместе кедр, чтобы украсить место святилища Моего, и Я прославлю подножие ног Моих.
ISA|60|14|И придут к тебе с покорностью сыновья угнетавших тебя, и падут к стопам ног твоих все, презиравшие тебя, и назовут тебя городом Господа, Сионом Святаго Израилева.
ISA|60|15|Вместо того, что ты был оставлен и ненавидим, так что никто не проходил чрез [тебя], Я соделаю тебя величием навеки, радостью в роды родов.
ISA|60|16|Ты будешь насыщаться молоком народов, и груди царские сосать будешь, и узнаешь, что Я Господь – Спаситель твой и Искупитель твой, Сильный Иаковлев.
ISA|60|17|Вместо меди буду доставлять тебе золото, и вместо железа серебро, и вместо дерева медь, и вместо камней железо; и поставлю правителем твоим мир и надзирателями твоими – правду.
ISA|60|18|Не слышно будет более насилия в земле твоей, опустошения и разорения – в пределах твоих; и будешь называть стены твои спасением и ворота твои – славою.
ISA|60|19|Не будет уже солнце служить тебе светом дневным, и сияние луны – светить тебе; но Господь будет тебе вечным светом, и Бог твой – славою твоею.
ISA|60|20|Не зайдет уже солнце твое, и луна твоя не сокроется, ибо Господь будет для тебя вечным светом, и окончатся дни сетования твоего.
ISA|60|21|И народ твой весь будет праведный, на веки наследует землю, – отрасль насаждения Моего, дело рук Моих, к прославлению Моему.
ISA|60|22|От малого произойдет тысяча, и от самого слабого – сильный народ. Я, Господь, ускорю совершить это в свое время.
ISA|61|1|Дух Господа Бога на Мне, ибо Господь помазал Меня благовествовать нищим, послал Меня исцелять сокрушенных сердцем, проповедывать пленным освобождение и узникам открытие темницы,
ISA|61|2|проповедывать лето Господне благоприятное и день мщения Бога нашего, утешить всех сетующих,
ISA|61|3|возвестить сетующим на Сионе, что им вместо пепла дастся украшение, вместо плача – елей радости, вместо унылого духа – славная одежда, и назовут их сильными правдою, насаждением Господа во славу Его.
ISA|61|4|И застроят пустыни вековые, восстановят древние развалины и возобновят города разоренные, остававшиеся в запустении с давних родов.
ISA|61|5|И придут иноземцы и будут пасти стада ваши; и сыновья чужестранцев [будут] вашими земледельцами и вашими виноградарями.
ISA|61|6|А вы будете называться священниками Господа, служителями Бога нашего будут именовать вас; будете пользоваться достоянием народов и славиться славою их.
ISA|61|7|За посрамление вам будет вдвое; за поношение они будут радоваться своей доле, потому что в земле своей вдвое получат; веселие вечное будет у них.
ISA|61|8|Ибо Я, Господь, люблю правосудие, ненавижу грабительство с насилием, и воздам награду им по истине, и завет вечный поставлю с ними;
ISA|61|9|и будет известно между народами семя их, и потомство их – среди племен; все видящие их познают, что они семя, благословенное Господом.
ISA|61|10|Радостью буду радоваться о Господе, возвеселится душа моя о Боге моем; ибо Он облек меня в ризы спасения, одеждою правды одел меня, как на жениха возложил венец и, как невесту, украсил убранством.
ISA|61|11|Ибо, как земля производит растения свои, и как сад произращает посеянное в нем, так Господь Бог проявит правду и славу пред всеми народами.
ISA|62|1|Не умолкну ради Сиона, и ради Иерусалима не успокоюсь, доколе не взойдет, как свет, правда его и спасение его – как горящий светильник.
ISA|62|2|И увидят народы правду твою и все цари – славу твою, и назовут тебя новым именем, которое нарекут уста Господа.
ISA|62|3|И будешь венцом славы в руке Господа и царскою диадемою на длани Бога твоего.
ISA|62|4|Не будут уже называть тебя "оставленным", и землю твою не будут более называть "пустынею", но будут называть тебя: "Мое благоволение к нему", а землю твою – "замужнею", ибо Господь благоволит к тебе, и земля твоя сочетается.
ISA|62|5|Как юноша сочетается с девою, так сочетаются с тобою сыновья твои; и [как] жених радуется о невесте, так будет радоваться о тебе Бог твой.
ISA|62|6|На стенах твоих, Иерусалим, Я поставил сторожей, [которые] не будут умолкать ни днем, ни ночью. О, вы, напоминающие о Господе! не умолкайте, –
ISA|62|7|не умолкайте пред Ним, доколе Он не восстановит и доколе не сделает Иерусалима славою на земле.
ISA|62|8|Господь поклялся десницею Своею и крепкою мышцею Своею: не дам зерна твоего более в пищу врагам твоим, и сыновья чужих не будут пить вина твоего, над которым ты трудился;
ISA|62|9|но собирающие его будут есть его и славить Господа, и обирающие виноград будут пить [вино] его во дворах святилища Моего.
ISA|62|10|Проходите, проходите в ворота, приготовляйте путь народу! Ровняйте, ровняйте дорогу, убирайте камни, поднимите знамя для народов!
ISA|62|11|Вот, Господь объявляет до конца земли: скажите дщери Сиона: грядет Спаситель твой; награда Его с Ним и воздаяние Его пред Ним.
ISA|62|12|И назовут их народом святым, искупленным от Господа, а тебя назовут взысканным городом, неоставленным.
ISA|63|1|Кто это идет от Едома, в червленых ризах от Восора, столь величественный в Своей одежде, выступающий в полноте силы Своей? "Я – изрекающий правду, сильный, чтобы спасать".
ISA|63|2|Отчего же одеяние Твое красно, и ризы у Тебя, как у топтавшего в точиле?
ISA|63|3|"Я топтал точило один, и из народов никого не было со Мною; и Я топтал их во гневе Моем и попирал их в ярости Моей; кровь их брызгала на ризы Мои, и Я запятнал все одеяние Свое;
ISA|63|4|ибо день мщения – в сердце Моем, и год Моих искупленных настал.
ISA|63|5|Я смотрел, и не было помощника; дивился, что не было поддерживающего; но помогла Мне мышца Моя, и ярость Моя – она поддержала Меня:
ISA|63|6|и попрал Я народы во гневе Моем, и сокрушил их в ярости Моей, и вылил на землю кровь их".
ISA|63|7|Воспомяну милости Господни и славу Господню за все, что Господь даровал нам, и великую благость [Его] к дому Израилеву, какую оказал Он ему по милосердию Своему и по множеству щедрот Своих.
ISA|63|8|Он сказал: "подлинно они народ Мой, дети, которые не солгут", и Он был для них Спасителем.
ISA|63|9|Во всякой скорби их Он не оставлял их, и Ангел лица Его спасал их; по любви Своей и благосердию Своему Он искупил их, взял и носил их во все дни древние.
ISA|63|10|Но они возмутились и огорчили Святаго Духа Его; поэтому Он обратился в неприятеля их: Сам воевал против них.
ISA|63|11|Тогда народ Его вспомнил древние дни, Моисеевы: где Тот, Который вывел их из моря с пастырем овец Своих? где Тот, Который вложил в сердце его Святаго Духа Своего,
ISA|63|12|Который вел Моисея за правую руку величественною мышцею Своею, разделил пред ними воды, чтобы сделать Себе вечное имя,
ISA|63|13|Который вел их чрез бездны, как коня по степи, [и] они не спотыкались?
ISA|63|14|Как стадо сходит в долину, Дух Господень вел их к покою. Так вел Ты народ Твой, чтобы сделать Себе славное имя.
ISA|63|15|Призри с небес и посмотри из жилища святыни Твоей и славы Твоей: где ревность Твоя и могущество Твое? – благоутробие Твое и милости Твои ко мне удержаны.
ISA|63|16|Только Ты – Отец наш; ибо Авраам не узнает нас, и Израиль не признает нас своими; Ты, Господи, Отец наш, от века имя Твое: "Искупитель наш".
ISA|63|17|Для чего, Господи, Ты попустил нам совратиться с путей Твоих, ожесточиться сердцу нашему, чтобы не бояться Тебя? обратись ради рабов Твоих, ради колен наследия Твоего.
ISA|63|18|Короткое время владел им народ святыни Твоей: враги наши попрали святилище Твое.
ISA|63|19|Мы сделались такими, над которыми Ты как бы никогда не владычествовал и над которыми не именовалось имя Твое.
ISA|64|1|О, если бы Ты расторг небеса [и] сошел! горы растаяли бы от лица Твоего,
ISA|64|2|как от плавящего огня, как от кипятящего воду, чтобы имя Твое сделать известным врагам Твоим; от лица Твоего содрогнулись бы народы.
ISA|64|3|Когда Ты совершал страшные дела, нами неожиданные, и нисходил, – горы таяли от лица Твоего.
ISA|64|4|Ибо от века не слыхали, не внимали ухом, и никакой глаз не видал другого бога, кроме Тебя, который столько сделал бы для надеющихся на него.
ISA|64|5|Ты милостиво встречал радующегося и делающего правду, поминающего Тебя на путях Твоих. Но вот, Ты прогневался, потому что мы издавна грешили; и как же мы будем спасены?
ISA|64|6|Все мы сделались – как нечистый, и вся праведность наша – как запачканная одежда; и все мы поблекли, как лист, и беззакония наши, как ветер, уносят нас.
ISA|64|7|И нет призывающего имя Твое, который положил бы крепко держаться за Тебя; поэтому Ты сокрыл от нас лице Твое и оставил нас погибать от беззаконий наших.
ISA|64|8|Но ныне, Господи, Ты – Отец наш; мы – глина, а Ты – образователь наш, и все мы – дело руки Твоей.
ISA|64|9|Не гневайся, Господи, без меры, и не вечно помни беззаконие. Воззри же: мы все народ Твой.
ISA|64|10|Города святыни Твоей сделались пустынею; пустынею стал Сион; Иерусалим опустошен.
ISA|64|11|Дом освящения нашего и славы нашей, где отцы наши прославляли Тебя, сожжен огнем, и все драгоценности наши разграблены.
ISA|64|12|После этого будешь ли еще удерживаться, Господи, будешь ли молчать и карать нас без меры?
ISA|65|1|Я открылся не вопрошавшим обо Мне; Меня нашли не искавшие Меня. "Вот Я! вот Я!" говорил Я народу, не именовавшемуся именем Моим.
ISA|65|2|Всякий день простирал Я руки Мои к народу непокорному, ходившему путем недобрым, по своим помышлениям, –
ISA|65|3|к народу, который постоянно оскорбляет Меня в лице, приносит жертвы в рощах и сожигает фимиам на черепках,
ISA|65|4|сидит в гробах и ночует в пещерах; ест свиное мясо, и мерзкое варево в сосудах у него;
ISA|65|5|который говорит: "остановись, не подходи ко мне, потому что я свят для тебя". Они – дым для обоняния Моего, огонь, горящий всякий день.
ISA|65|6|Вот что написано пред лицем Моим: не умолчу, но воздам, воздам в недро их
ISA|65|7|беззакония ваши, говорит Господь, и вместе беззакония отцов ваших, которые воскуряли фимиам на горах, и на холмах поносили Меня; и отмерю в недра их прежние деяния их.
ISA|65|8|Так говорит Господь: когда в виноградной кисти находится сок, тогда говорят: "не повреди ее, ибо в ней благословение"; то же сделаю Я и ради рабов Моих, чтобы не всех погубить.
ISA|65|9|И произведу от Иакова семя, и от Иуды наследника гор Моих, и наследуют это избранные Мои, и рабы Мои будут жить там.
ISA|65|10|И будет Сарон пастбищем для овец и долина Ахор – местом отдыха для волов народа Моего, который взыскал Меня.
ISA|65|11|А вас, которые оставили Господа, забыли святую гору Мою, приготовляете трапезу для Гада и растворяете полную чашу для Мени, –
ISA|65|12|вас обрекаю Я мечу, и все вы преклонитесь на заклание: потому что Я звал, и вы не отвечали; говорил, и вы не слушали, но делали злое в очах Моих и избирали то, что было неугодно Мне.
ISA|65|13|Посему так говорит Господь Бог: вот, рабы Мои будут есть, а вы будете голодать; рабы Мои будут пить, а вы будете томиться жаждою;
ISA|65|14|рабы Мои будут веселиться, а вы будете в стыде; рабы Мои будут петь от сердечной радости, а вы будете кричать от сердечной скорби и рыдать от сокрушения духа.
ISA|65|15|И оставите имя ваше избранным Моим для проклятия; и убьет тебя Господь Бог, а рабов Своих назовет иным именем,
ISA|65|16|которым кто будет благословлять себя на земле, будет благословляться Богом истины; и кто будет клясться на земле, будет клясться Богом истины, – потому что прежние скорби будут забыты и сокрыты от очей Моих.
ISA|65|17|Ибо вот, Я творю новое небо и новую землю, и прежние уже не будут воспоминаемы и не придут на сердце.
ISA|65|18|А вы будете веселиться и радоваться вовеки о том, что Я творю: ибо вот, Я творю Иерусалим веселием и народ его радостью.
ISA|65|19|И буду радоваться о Иерусалиме и веселиться о народе Моем; и не услышится в нем более голос плача и голос вопля.
ISA|65|20|Там не будет более малолетнего и старца, который не достигал бы полноты дней своих; ибо столетний будет умирать юношею, но столетний грешник будет проклинаем.
ISA|65|21|И буду строить домы и жить в них, и насаждать виноградники и есть плоды их.
ISA|65|22|Не будут строить, чтобы другой жил, не будут насаждать, чтобы другой ел; ибо дни народа Моего будут, как дни дерева, и избранные Мои долго будут пользоваться изделием рук своих.
ISA|65|23|Не будут трудиться напрасно и рождать детей на горе; ибо будут семенем, благословенным от Господа, и потомки их с ними.
ISA|65|24|И будет, прежде нежели они воззовут, Я отвечу; они еще будут говорить, и Я уже услышу.
ISA|65|25|Волк и ягненок будут пастись вместе, и лев, как вол, будет есть солому, а для змея прах будет пищею: они не будут причинять зла и вреда на всей святой горе Моей, говорит Господь.
ISA|66|1|Так говорит Господь: небо – престол Мой, а земля – подножие ног Моих; где же построите вы дом для Меня, и где место покоя Моего?
ISA|66|2|Ибо все это соделала рука Моя, и все сие было, говорит Господь. А вот на кого Я призрю: на смиренного и сокрушенного духом и на трепещущего пред словом Моим.
ISA|66|3|Заколающий вола – то же, что убивающий человека; приносящий агнца в жертву – то же, что задушающий пса; приносящий семидал – то же, что приносящий свиную кровь; воскуряющий фимиам – то же, что молящийся идолу; и как они избрали собственные свои пути, и душа их находит удовольствие в мерзостях их, –
ISA|66|4|так и Я употреблю их обольщение и наведу на них ужасное для них: потому что Я звал, и не было отвечающего, говорил, и они не слушали, а делали злое в очах Моих и избирали то, что неугодно Мне.
ISA|66|5|Выслушайте слово Господа, трепещущие пред словом Его: ваши братья, ненавидящие вас и изгоняющие вас за имя Мое, говорят: "пусть явит Себя в славе Господь, и мы посмотрим на веселие ваше". Но они будут постыжены.
ISA|66|6|Вот, шум из города, голос из храма, голос Господа, воздающего возмездие врагам Своим.
ISA|66|7|Еще не мучилась родами, а родила; прежде нежели наступили боли ее, разрешилась сыном.
ISA|66|8|Кто слыхал таковое? кто видал подобное этому? возникала ли страна в один день? рождался ли народ в один раз, как Сион, едва начал родами мучиться, родил сынов своих?
ISA|66|9|Доведу ли Я до родов, и не дам родить? говорит Господь. Или, давая силу родить, заключу ли [утробу]? говорит Бог твой.
ISA|66|10|Возвеселитесь с Иерусалимом и радуйтесь о нем, все любящие его! возрадуйтесь с ним радостью, все сетовавшие о нем,
ISA|66|11|чтобы вам питаться и насыщаться от сосцов утешений его, упиваться и наслаждаться преизбытком славы его.
ISA|66|12|Ибо так говорит Господь: вот, Я направляю к нему мир как реку, и богатство народов – как разливающийся поток для наслаждения вашего; на руках будут носить вас и на коленях ласкать.
ISA|66|13|Как утешает кого–либо мать его, так утешу Я вас, и вы будете утешены в Иерусалиме.
ISA|66|14|И увидите это, и возрадуется сердце ваше, и кости ваши расцветут, как молодая зелень, и откроется рука Господа рабам Его, а на врагов Своих Он разгневается.
ISA|66|15|Ибо вот, придет Господь в огне, и колесницы Его – как вихрь, чтобы излить гнев Свой с яростью и прещение Свое с пылающим огнем.
ISA|66|16|Ибо Господь с огнем и мечом Своим произведет суд над всякою плотью, и много будет пораженных Господом.
ISA|66|17|Те, которые освящают и очищают себя в рощах, один за другим, едят свиное мясо и мерзость и мышей, – все погибнут, говорит Господь.
ISA|66|18|Ибо Я [знаю] деяния их и мысли их; и вот, приду собрать все народы и языки, и они придут и увидят славу Мою.
ISA|66|19|И положу на них знамение, и пошлю из спасенных от них к народам: в Фарсис, к Пулу и Луду, к натягивающим лук, к Тубалу и Явану, на дальние острова, которые не слышали обо Мне и не видели славы Моей: и они возвестят народам славу Мою
ISA|66|20|и представят всех братьев ваших от всех народов в дар Господу на конях и колесницах, и на носилках, и на мулах, и на быстрых верблюдах, на святую гору Мою, в Иерусалим, говорит Господь, – подобно тому, как сыны Израилевы приносят дар в дом Господа в чистом сосуде.
ISA|66|21|Из них буду брать также в священники и левиты, говорит Господь.
ISA|66|22|Ибо, как новое небо и новая земля, которые Я сотворю, всегда будут пред лицем Моим, говорит Господь, так будет и семя ваше и имя ваше.
ISA|66|23|Тогда из месяца в месяц и из субботы в субботу будет приходить всякая плоть пред лице Мое на поклонение, говорит Господь.
ISA|66|24|И будут выходить и увидят трупы людей, отступивших от Меня: ибо червь их не умрет, и огонь их не угаснет; и будут они мерзостью для всякой плоти.
