JER|1|1|The words of Jeremiah son of Hilkiah, one of the priests at Anathoth in the territory of Benjamin.
JER|1|2|The word of the LORD came to him in the thirteenth year of the reign of Josiah son of Amon king of Judah,
JER|1|3|and through the reign of Jehoiakim son of Josiah king of Judah, down to the fifth month of the eleventh year of Zedekiah son of Josiah king of Judah, when the people of Jerusalem went into exile.
JER|1|4|The word of the LORD came to me, saying,
JER|1|5|"Before I formed you in the womb I knew you, before you were born I set you apart; I appointed you as a prophet to the nations."
JER|1|6|"Ah, Sovereign LORD," I said, "I do not know how to speak; I am only a child."
JER|1|7|But the LORD said to me, "Do not say, 'I am only a child.' You must go to everyone I send you to and say whatever I command you.
JER|1|8|Do not be afraid of them, for I am with you and will rescue you," declares the LORD.
JER|1|9|Then the LORD reached out his hand and touched my mouth and said to me, "Now, I have put my words in your mouth.
JER|1|10|See, today I appoint you over nations and kingdoms to uproot and tear down, to destroy and overthrow, to build and to plant."
JER|1|11|The word of the LORD came to me: "What do you see, Jeremiah?I see the branch of an almond tree," I replied.
JER|1|12|The LORD said to me, "You have seen correctly, for I am watching to see that my word is fulfilled."
JER|1|13|The word of the LORD came to me again: "What do you see?I see a boiling pot, tilting away from the north," I answered.
JER|1|14|The LORD said to me, "From the north disaster will be poured out on all who live in the land.
JER|1|15|I am about to summon all the peoples of the northern kingdoms," declares the LORD. "Their kings will come and set up their thrones in the entrance of the gates of Jerusalem; they will come against all her surrounding walls and against all the towns of Judah.
JER|1|16|I will pronounce my judgments on my people because of their wickedness in forsaking me, in burning incense to other gods and in worshiping what their hands have made.
JER|1|17|"Get yourself ready! Stand up and say to them whatever I command you. Do not be terrified by them, or I will terrify you before them.
JER|1|18|Today I have made you a fortified city, an iron pillar and a bronze wall to stand against the whole land-against the kings of Judah, its officials, its priests and the people of the land.
JER|1|19|They will fight against you but will not overcome you, for I am with you and will rescue you," declares the LORD.
JER|2|1|The word of the LORD came to me:
JER|2|2|"Go and proclaim in the hearing of Jerusalem: "'I remember the devotion of your youth, how as a bride you loved me and followed me through the desert, through a land not sown.
JER|2|3|Israel was holy to the LORD, the firstfruits of his harvest; all who devoured her were held guilty, and disaster overtook them,'" declares the LORD.
JER|2|4|Hear the word of the LORD, O house of Jacob, all you clans of the house of Israel.
JER|2|5|This is what the LORD says: "What fault did your fathers find in me, that they strayed so far from me? They followed worthless idols and became worthless themselves.
JER|2|6|They did not ask, 'Where is the LORD, who brought us up out of Egypt and led us through the barren wilderness, through a land of deserts and rifts, a land of drought and darkness, a land where no one travels and no one lives?'
JER|2|7|I brought you into a fertile land to eat its fruit and rich produce. But you came and defiled my land and made my inheritance detestable.
JER|2|8|The priests did not ask, 'Where is the LORD?' Those who deal with the law did not know me; the leaders rebelled against me. The prophets prophesied by Baal, following worthless idols.
JER|2|9|"Therefore I bring charges against you again," declares the LORD. "And I will bring charges against your children's children.
JER|2|10|Cross over to the coasts of Kittim and look, send to Kedar and observe closely; see if there has ever been anything like this:
JER|2|11|Has a nation ever changed its gods? (Yet they are not gods at all.) But my people have exchanged their Glory for worthless idols.
JER|2|12|Be appalled at this, O heavens, and shudder with great horror," declares the LORD.
JER|2|13|"My people have committed two sins: They have forsaken me, the spring of living water, and have dug their own cisterns, broken cisterns that cannot hold water.
JER|2|14|Is Israel a servant, a slave by birth? Why then has he become plunder?
JER|2|15|Lions have roared; they have growled at him. They have laid waste his land; his towns are burned and deserted.
JER|2|16|Also, the men of Memphis and Tahpanhes have shaved the crown of your head.
JER|2|17|Have you not brought this on yourselves by forsaking the LORD your God when he led you in the way?
JER|2|18|Now why go to Egypt to drink water from the Shihor? And why go to Assyria to drink water from the River?
JER|2|19|Your wickedness will punish you; your backsliding will rebuke you. Consider then and realize how evil and bitter it is for you when you forsake the LORD your God and have no awe of me," declares the Lord, the LORD Almighty.
JER|2|20|"Long ago you broke off your yoke and tore off your bonds; you said, 'I will not serve you!' Indeed, on every high hill and under every spreading tree you lay down as a prostitute.
JER|2|21|I had planted you like a choice vine of sound and reliable stock. How then did you turn against me into a corrupt, wild vine?
JER|2|22|Although you wash yourself with soda and use an abundance of soap, the stain of your guilt is still before me," declares the Sovereign LORD.
JER|2|23|"How can you say, 'I am not defiled; I have not run after the Baals'? See how you behaved in the valley; consider what you have done. You are a swift she-camel running here and there,
JER|2|24|a wild donkey accustomed to the desert, sniffing the wind in her craving- in her heat who can restrain her? Any males that pursue her need not tire themselves; at mating time they will find her.
JER|2|25|Do not run until your feet are bare and your throat is dry. But you said, 'It's no use! I love foreign gods, and I must go after them.'
JER|2|26|"As a thief is disgraced when he is caught, so the house of Israel is disgraced- they, their kings and their officials, their priests and their prophets.
JER|2|27|They say to wood, 'You are my father,' and to stone, 'You gave me birth.' They have turned their backs to me and not their faces; yet when they are in trouble, they say, 'Come and save us!'
JER|2|28|Where then are the gods you made for yourselves? Let them come if they can save you when you are in trouble! For you have as many gods as you have towns, O Judah.
JER|2|29|"Why do you bring charges against me? You have all rebelled against me," declares the LORD.
JER|2|30|"In vain I punished your people; they did not respond to correction. Your sword has devoured your prophets like a ravening lion.
JER|2|31|"You of this generation, consider the word of the LORD: "Have I been a desert to Israel or a land of great darkness? Why do my people say, 'We are free to roam; we will come to you no more'?
JER|2|32|Does a maiden forget her jewelry, a bride her wedding ornaments? Yet my people have forgotten me, days without number.
JER|2|33|How skilled you are at pursuing love! Even the worst of women can learn from your ways.
JER|2|34|On your clothes men find the lifeblood of the innocent poor, though you did not catch them breaking in. Yet in spite of all this
JER|2|35|you say, 'I am innocent; he is not angry with me.' But I will pass judgment on you because you say, 'I have not sinned.'
JER|2|36|Why do you go about so much, changing your ways? You will be disappointed by Egypt as you were by Assyria.
JER|2|37|You will also leave that place with your hands on your head, for the LORD has rejected those you trust; you will not be helped by them.
JER|3|1|"If a man divorces his wife and she leaves him and marries another man, should he return to her again? Would not the land be completely defiled? But you have lived as a prostitute with many lovers- would you now return to me?" declares the LORD.
JER|3|2|"Look up to the barren heights and see. Is there any place where you have not been ravished? By the roadside you sat waiting for lovers, sat like a nomad in the desert. You have defiled the land with your prostitution and wickedness.
JER|3|3|Therefore the showers have been withheld, and no spring rains have fallen. Yet you have the brazen look of a prostitute; you refuse to blush with shame.
JER|3|4|Have you not just called to me: 'My Father, my friend from my youth,
JER|3|5|will you always be angry? Will your wrath continue forever?' This is how you talk, but you do all the evil you can."
JER|3|6|During the reign of King Josiah, the LORD said to me, "Have you seen what faithless Israel has done? She has gone up on every high hill and under every spreading tree and has committed adultery there.
JER|3|7|I thought that after she had done all this she would return to me but she did not, and her unfaithful sister Judah saw it.
JER|3|8|I gave faithless Israel her certificate of divorce and sent her away because of all her adulteries. Yet I saw that her unfaithful sister Judah had no fear; she also went out and committed adultery.
JER|3|9|Because Israel's immorality mattered so little to her, she defiled the land and committed adultery with stone and wood.
JER|3|10|In spite of all this, her unfaithful sister Judah did not return to me with all her heart, but only in pretense," declares the LORD.
JER|3|11|The LORD said to me, "Faithless Israel is more righteous than unfaithful Judah.
JER|3|12|Go, proclaim this message toward the north: "'Return, faithless Israel,' declares the LORD, 'I will frown on you no longer, for I am merciful,' declares the LORD, 'I will not be angry forever.
JER|3|13|Only acknowledge your guilt- you have rebelled against the LORD your God, you have scattered your favors to foreign gods under every spreading tree, and have not obeyed me,'" declares the LORD.
JER|3|14|"Return, faithless people," declares the LORD, "for I am your husband. I will choose you-one from a town and two from a clan-and bring you to Zion.
JER|3|15|Then I will give you shepherds after my own heart, who will lead you with knowledge and understanding.
JER|3|16|In those days, when your numbers have increased greatly in the land," declares the LORD, "men will no longer say, 'The ark of the covenant of the LORD.' It will never enter their minds or be remembered; it will not be missed, nor will another one be made.
JER|3|17|At that time they will call Jerusalem The Throne of the LORD, and all nations will gather in Jerusalem to honor the name of the LORD. No longer will they follow the stubbornness of their evil hearts.
JER|3|18|In those days the house of Judah will join the house of Israel, and together they will come from a northern land to the land I gave your forefathers as an inheritance.
JER|3|19|"I myself said, "'How gladly would I treat you like sons and give you a desirable land, the most beautiful inheritance of any nation.' I thought you would call me 'Father' and not turn away from following me.
JER|3|20|But like a woman unfaithful to her husband, so you have been unfaithful to me, O house of Israel," declares the LORD.
JER|3|21|A cry is heard on the barren heights, the weeping and pleading of the people of Israel, because they have perverted their ways and have forgotten the LORD their God.
JER|3|22|"Return, faithless people; I will cure you of backsliding.Yes, we will come to you, for you are the LORD our God.
JER|3|23|Surely the idolatrous commotion on the hills and mountains is a deception; surely in the LORD our God is the salvation of Israel.
JER|3|24|From our youth shameful gods have consumed the fruits of our fathers' labor- their flocks and herds, their sons and daughters.
JER|3|25|Let us lie down in our shame, and let our disgrace cover us. We have sinned against the LORD our God, both we and our fathers; from our youth till this day we have not obeyed the LORD our God."
JER|4|1|"If you will return, O Israel, return to me," declares the LORD. "If you put your detestable idols out of my sight and no longer go astray,
JER|4|2|and if in a truthful, just and righteous way you swear, 'As surely as the LORD lives,' then the nations will be blessed by him and in him they will glory."
JER|4|3|This is what the LORD says to the men of Judah and to Jerusalem: "Break up your unplowed ground and do not sow among thorns.
JER|4|4|Circumcise yourselves to the LORD, circumcise your hearts, you men of Judah and people of Jerusalem, or my wrath will break out and burn like fire because of the evil you have done- burn with no one to quench it.
JER|4|5|"Announce in Judah and proclaim in Jerusalem and say: 'Sound the trumpet throughout the land!' Cry aloud and say: 'Gather together! Let us flee to the fortified cities!'
JER|4|6|Raise the signal to go to Zion! Flee for safety without delay! For I am bringing disaster from the north, even terrible destruction."
JER|4|7|A lion has come out of his lair; a destroyer of nations has set out. He has left his place to lay waste your land. Your towns will lie in ruins without inhabitant.
JER|4|8|So put on sackcloth, lament and wail, for the fierce anger of the LORD has not turned away from us.
JER|4|9|"In that day," declares the LORD, "the king and the officials will lose heart, the priests will be horrified, and the prophets will be appalled."
JER|4|10|Then I said, "Ah, Sovereign LORD, how completely you have deceived this people and Jerusalem by saying, 'You will have peace,' when the sword is at our throats."
JER|4|11|At that time this people and Jerusalem will be told, "A scorching wind from the barren heights in the desert blows toward my people, but not to winnow or cleanse;
JER|4|12|a wind too strong for that comes from me. Now I pronounce my judgments against them."
JER|4|13|Look! He advances like the clouds, his chariots come like a whirlwind, his horses are swifter than eagles. Woe to us! We are ruined!
JER|4|14|O Jerusalem, wash the evil from your heart and be saved. How long will you harbor wicked thoughts?
JER|4|15|A voice is announcing from Dan, proclaiming disaster from the hills of Ephraim.
JER|4|16|"Tell this to the nations, proclaim it to Jerusalem: 'A besieging army is coming from a distant land, raising a war cry against the cities of Judah.
JER|4|17|They surround her like men guarding a field, because she has rebelled against me,'" declares the LORD.
JER|4|18|"Your own conduct and actions have brought this upon you. This is your punishment. How bitter it is! How it pierces to the heart!"
JER|4|19|Oh, my anguish, my anguish! I writhe in pain. Oh, the agony of my heart! My heart pounds within me, I cannot keep silent. For I have heard the sound of the trumpet; I have heard the battle cry.
JER|4|20|Disaster follows disaster; the whole land lies in ruins. In an instant my tents are destroyed, my shelter in a moment.
JER|4|21|How long must I see the battle standard and hear the sound of the trumpet?
JER|4|22|"My people are fools; they do not know me. They are senseless children; they have no understanding. They are skilled in doing evil; they know not how to do good."
JER|4|23|I looked at the earth, and it was formless and empty; and at the heavens, and their light was gone.
JER|4|24|I looked at the mountains, and they were quaking; all the hills were swaying.
JER|4|25|I looked, and there were no people; every bird in the sky had flown away.
JER|4|26|I looked, and the fruitful land was a desert; all its towns lay in ruins before the LORD, before his fierce anger.
JER|4|27|This is what the LORD says: "The whole land will be ruined, though I will not destroy it completely.
JER|4|28|Therefore the earth will mourn and the heavens above grow dark, because I have spoken and will not relent, I have decided and will not turn back."
JER|4|29|At the sound of horsemen and archers every town takes to flight. Some go into the thickets; some climb up among the rocks. All the towns are deserted; no one lives in them.
JER|4|30|What are you doing, O devastated one? Why dress yourself in scarlet and put on jewels of gold? Why shade your eyes with paint? You adorn yourself in vain. Your lovers despise you; they seek your life.
JER|4|31|I hear a cry as of a woman in labor, a groan as of one bearing her first child- the cry of the Daughter of Zion gasping for breath, stretching out her hands and saying, "Alas! I am fainting; my life is given over to murderers."
JER|5|1|"Go up and down the streets of Jerusalem, look around and consider, search through her squares. If you can find but one person who deals honestly and seeks the truth, I will forgive this city.
JER|5|2|Although they say, 'As surely as the LORD lives,' still they are swearing falsely."
JER|5|3|O LORD, do not your eyes look for truth? You struck them, but they felt no pain; you crushed them, but they refused correction. They made their faces harder than stone and refused to repent.
JER|5|4|I thought, "These are only the poor; they are foolish, for they do not know the way of the LORD, the requirements of their God.
JER|5|5|So I will go to the leaders and speak to them; surely they know the way of the LORD, the requirements of their God." But with one accord they too had broken off the yoke and torn off the bonds.
JER|5|6|Therefore a lion from the forest will attack them, a wolf from the desert will ravage them, a leopard will lie in wait near their towns to tear to pieces any who venture out, for their rebellion is great and their backslidings many.
JER|5|7|"Why should I forgive you? Your children have forsaken me and sworn by gods that are not gods. I supplied all their needs, yet they committed adultery and thronged to the houses of prostitutes.
JER|5|8|They are well-fed, lusty stallions, each neighing for another man's wife.
JER|5|9|Should I not punish them for this?" declares the LORD. "Should I not avenge myself on such a nation as this?
JER|5|10|"Go through her vineyards and ravage them, but do not destroy them completely. Strip off her branches, for these people do not belong to the LORD.
JER|5|11|The house of Israel and the house of Judah have been utterly unfaithful to me," declares the LORD.
JER|5|12|They have lied about the LORD; they said, "He will do nothing! No harm will come to us; we will never see sword or famine.
JER|5|13|The prophets are but wind and the word is not in them; so let what they say be done to them."
JER|5|14|Therefore this is what the LORD God Almighty says: "Because the people have spoken these words, I will make my words in your mouth a fire and these people the wood it consumes.
JER|5|15|O house of Israel," declares the LORD, "I am bringing a distant nation against you- an ancient and enduring nation, a people whose language you do not know, whose speech you do not understand.
JER|5|16|Their quivers are like an open grave; all of them are mighty warriors.
JER|5|17|They will devour your harvests and food, devour your sons and daughters; they will devour your flocks and herds, devour your vines and fig trees. With the sword they will destroy the fortified cities in which you trust.
JER|5|18|"Yet even in those days," declares the LORD, "I will not destroy you completely.
JER|5|19|And when the people ask, 'Why has the LORD our God done all this to us?' you will tell them, 'As you have forsaken me and served foreign gods in your own land, so now you will serve foreigners in a land not your own.'
JER|5|20|"Announce this to the house of Jacob and proclaim it in Judah:
JER|5|21|Hear this, you foolish and senseless people, who have eyes but do not see, who have ears but do not hear:
JER|5|22|Should you not fear me?" declares the LORD. "Should you not tremble in my presence? I made the sand a boundary for the sea, an everlasting barrier it cannot cross. The waves may roll, but they cannot prevail; they may roar, but they cannot cross it.
JER|5|23|But these people have stubborn and rebellious hearts; they have turned aside and gone away.
JER|5|24|They do not say to themselves, 'Let us fear the LORD our God, who gives autumn and spring rains in season, who assures us of the regular weeks of harvest.'
JER|5|25|Your wrongdoings have kept these away; your sins have deprived you of good.
JER|5|26|"Among my people are wicked men who lie in wait like men who snare birds and like those who set traps to catch men.
JER|5|27|Like cages full of birds, their houses are full of deceit; they have become rich and powerful
JER|5|28|and have grown fat and sleek. Their evil deeds have no limit; they do not plead the case of the fatherless to win it, they do not defend the rights of the poor.
JER|5|29|Should I not punish them for this?" declares the LORD. "Should I not avenge myself on such a nation as this?
JER|5|30|"A horrible and shocking thing has happened in the land:
JER|5|31|The prophets prophesy lies, the priests rule by their own authority, and my people love it this way. But what will you do in the end?
JER|6|1|"Flee for safety, people of Benjamin! Flee from Jerusalem! Sound the trumpet in Tekoa! Raise the signal over Beth Hakkerem! For disaster looms out of the north, even terrible destruction.
JER|6|2|I will destroy the Daughter of Zion, so beautiful and delicate.
JER|6|3|Shepherds with their flocks will come against her; they will pitch their tents around her, each tending his own portion."
JER|6|4|"Prepare for battle against her! Arise, let us attack at noon! But, alas, the daylight is fading, and the shadows of evening grow long.
JER|6|5|So arise, let us attack at night and destroy her fortresses!"
JER|6|6|This is what the LORD Almighty says: "Cut down the trees and build siege ramps against Jerusalem. This city must be punished; it is filled with oppression.
JER|6|7|As a well pours out its water, so she pours out her wickedness. Violence and destruction resound in her; her sickness and wounds are ever before me.
JER|6|8|Take warning, O Jerusalem, or I will turn away from you and make your land desolate so no one can live in it."
JER|6|9|This is what the LORD Almighty says: "Let them glean the remnant of Israel as thoroughly as a vine; pass your hand over the branches again, like one gathering grapes."
JER|6|10|To whom can I speak and give warning? Who will listen to me? Their ears are closed so they cannot hear. The word of the LORD is offensive to them; they find no pleasure in it.
JER|6|11|But I am full of the wrath of the LORD, and I cannot hold it in. "Pour it out on the children in the street and on the young men gathered together; both husband and wife will be caught in it, and the old, those weighed down with years.
JER|6|12|Their houses will be turned over to others, together with their fields and their wives, when I stretch out my hand against those who live in the land," declares the LORD.
JER|6|13|"From the least to the greatest, all are greedy for gain; prophets and priests alike, all practice deceit.
JER|6|14|They dress the wound of my people as though it were not serious. 'Peace, peace,' they say, when there is no peace.
JER|6|15|Are they ashamed of their loathsome conduct? No, they have no shame at all; they do not even know how to blush. So they will fall among the fallen; they will be brought down when I punish them," says the LORD.
JER|6|16|This is what the LORD says: "Stand at the crossroads and look; ask for the ancient paths, ask where the good way is, and walk in it, and you will find rest for your souls. But you said, 'We will not walk in it.'
JER|6|17|I appointed watchmen over you and said, 'Listen to the sound of the trumpet!' But you said, 'We will not listen.'
JER|6|18|Therefore hear, O nations; observe, O witnesses, what will happen to them.
JER|6|19|Hear, O earth: I am bringing disaster on this people, the fruit of their schemes, because they have not listened to my words and have rejected my law.
JER|6|20|What do I care about incense from Sheba or sweet calamus from a distant land? Your burnt offerings are not acceptable; your sacrifices do not please me."
JER|6|21|Therefore this is what the LORD says: "I will put obstacles before this people. Fathers and sons alike will stumble over them; neighbors and friends will perish."
JER|6|22|This is what the LORD says: "Look, an army is coming from the land of the north; a great nation is being stirred up from the ends of the earth.
JER|6|23|They are armed with bow and spear; they are cruel and show no mercy. They sound like the roaring sea as they ride on their horses; they come like men in battle formation to attack you, O Daughter of Zion."
JER|6|24|We have heard reports about them, and our hands hang limp. Anguish has gripped us, pain like that of a woman in labor.
JER|6|25|Do not go out to the fields or walk on the roads, for the enemy has a sword, and there is terror on every side.
JER|6|26|O my people, put on sackcloth and roll in ashes; mourn with bitter wailing as for an only son, for suddenly the destroyer will come upon us.
JER|6|27|"I have made you a tester of metals and my people the ore, that you may observe and test their ways.
JER|6|28|They are all hardened rebels, going about to slander. They are bronze and iron; they all act corruptly.
JER|6|29|The bellows blow fiercely to burn away the lead with fire, but the refining goes on in vain; the wicked are not purged out.
JER|6|30|They are called rejected silver, because the LORD has rejected them."
JER|7|1|This is the word that came to Jeremiah from the LORD:
JER|7|2|"Stand at the gate of the LORD's house and there proclaim this message: "'Hear the word of the LORD, all you people of Judah who come through these gates to worship the LORD.
JER|7|3|This is what the LORD Almighty, the God of Israel, says: Reform your ways and your actions, and I will let you live in this place.
JER|7|4|Do not trust in deceptive words and say, "This is the temple of the LORD, the temple of the LORD, the temple of the LORD!"
JER|7|5|If you really change your ways and your actions and deal with each other justly,
JER|7|6|if you do not oppress the alien, the fatherless or the widow and do not shed innocent blood in this place, and if you do not follow other gods to your own harm,
JER|7|7|then I will let you live in this place, in the land I gave your forefathers for ever and ever.
JER|7|8|But look, you are trusting in deceptive words that are worthless.
JER|7|9|"'Will you steal and murder, commit adultery and perjury, burn incense to Baal and follow other gods you have not known,
JER|7|10|and then come and stand before me in this house, which bears my Name, and say, "We are safe"-safe to do all these detestable things?
JER|7|11|Has this house, which bears my Name, become a den of robbers to you? But I have been watching! declares the LORD.
JER|7|12|"'Go now to the place in Shiloh where I first made a dwelling for my Name, and see what I did to it because of the wickedness of my people Israel.
JER|7|13|While you were doing all these things, declares the LORD, I spoke to you again and again, but you did not listen; I called you, but you did not answer.
JER|7|14|Therefore, what I did to Shiloh I will now do to the house that bears my Name, the temple you trust in, the place I gave to you and your fathers.
JER|7|15|I will thrust you from my presence, just as I did all your brothers, the people of Ephraim.'
JER|7|16|"So do not pray for this people nor offer any plea or petition for them; do not plead with me, for I will not listen to you.
JER|7|17|Do you not see what they are doing in the towns of Judah and in the streets of Jerusalem?
JER|7|18|The children gather wood, the fathers light the fire, and the women knead the dough and make cakes of bread for the Queen of Heaven. They pour out drink offerings to other gods to provoke me to anger.
JER|7|19|But am I the one they are provoking? declares the LORD. Are they not rather harming themselves, to their own shame?
JER|7|20|"'Therefore this is what the Sovereign LORD says: My anger and my wrath will be poured out on this place, on man and beast, on the trees of the field and on the fruit of the ground, and it will burn and not be quenched.
JER|7|21|"'This is what the LORD Almighty, the God of Israel, says: Go ahead, add your burnt offerings to your other sacrifices and eat the meat yourselves!
JER|7|22|For when I brought your forefathers out of Egypt and spoke to them, I did not just give them commands about burnt offerings and sacrifices,
JER|7|23|but I gave them this command: Obey me, and I will be your God and you will be my people. Walk in all the ways I command you, that it may go well with you.
JER|7|24|But they did not listen or pay attention; instead, they followed the stubborn inclinations of their evil hearts. They went backward and not forward.
JER|7|25|From the time your forefathers left Egypt until now, day after day, again and again I sent you my servants the prophets.
JER|7|26|But they did not listen to me or pay attention. They were stiff-necked and did more evil than their forefathers.'
JER|7|27|"When you tell them all this, they will not listen to you; when you call to them, they will not answer.
JER|7|28|Therefore say to them, 'This is the nation that has not obeyed the LORD its God or responded to correction. Truth has perished; it has vanished from their lips.
JER|7|29|Cut off your hair and throw it away; take up a lament on the barren heights, for the LORD has rejected and abandoned this generation that is under his wrath.
JER|7|30|"'The people of Judah have done evil in my eyes, declares the LORD. They have set up their detestable idols in the house that bears my Name and have defiled it.
JER|7|31|They have built the high places of Topheth in the Valley of Ben Hinnom to burn their sons and daughters in the fire-something I did not command, nor did it enter my mind.
JER|7|32|So beware, the days are coming, declares the LORD, when people will no longer call it Topheth or the Valley of Ben Hinnom, but the Valley of Slaughter, for they will bury the dead in Topheth until there is no more room.
JER|7|33|Then the carcasses of this people will become food for the birds of the air and the beasts of the earth, and there will be no one to frighten them away.
JER|7|34|I will bring an end to the sounds of joy and gladness and to the voices of bride and bridegroom in the towns of Judah and the streets of Jerusalem, for the land will become desolate.
JER|8|1|"'At that time, declares the LORD, the bones of the kings and officials of Judah, the bones of the priests and prophets, and the bones of the people of Jerusalem will be removed from their graves.
JER|8|2|They will be exposed to the sun and the moon and all the stars of the heavens, which they have loved and served and which they have followed and consulted and worshiped. They will not be gathered up or buried, but will be like refuse lying on the ground.
JER|8|3|Wherever I banish them, all the survivors of this evil nation will prefer death to life, declares the LORD Almighty.'
JER|8|4|"Say to them, 'This is what the LORD says: "'When men fall down, do they not get up? When a man turns away, does he not return?
JER|8|5|Why then have these people turned away? Why does Jerusalem always turn away? They cling to deceit; they refuse to return.
JER|8|6|I have listened attentively, but they do not say what is right. No one repents of his wickedness, saying, "What have I done?" Each pursues his own course like a horse charging into battle.
JER|8|7|Even the stork in the sky knows her appointed seasons, and the dove, the swift and the thrush observe the time of their migration. But my people do not know the requirements of the LORD.
JER|8|8|"'How can you say, "We are wise, for we have the law of the LORD," when actually the lying pen of the scribes has handled it falsely?
JER|8|9|The wise will be put to shame; they will be dismayed and trapped. Since they have rejected the word of the LORD, what kind of wisdom do they have?
JER|8|10|Therefore I will give their wives to other men and their fields to new owners. From the least to the greatest, all are greedy for gain; prophets and priests alike, all practice deceit.
JER|8|11|They dress the wound of my people as though it were not serious. "Peace, peace," they say, when there is no peace.
JER|8|12|Are they ashamed of their loathsome conduct? No, they have no shame at all; they do not even know how to blush. So they will fall among the fallen; they will be brought down when they are punished, says the LORD.
JER|8|13|"'I will take away their harvest, declares the LORD. There will be no grapes on the vine. There will be no figs on the tree, and their leaves will wither. What I have given them will be taken from them. '"
JER|8|14|"Why are we sitting here? Gather together! Let us flee to the fortified cities and perish there! For the LORD our God has doomed us to perish and given us poisoned water to drink, because we have sinned against him.
JER|8|15|We hoped for peace but no good has come, for a time of healing but there was only terror.
JER|8|16|The snorting of the enemy's horses is heard from Dan; at the neighing of their stallions the whole land trembles. They have come to devour the land and everything in it, the city and all who live there."
JER|8|17|"See, I will send venomous snakes among you, vipers that cannot be charmed, and they will bite you," declares the LORD.
JER|8|18|O my Comforter in sorrow, my heart is faint within me.
JER|8|19|Listen to the cry of my people from a land far away: "Is the LORD not in Zion? Is her King no longer there?Why have they provoked me to anger with their images, with their worthless foreign idols?"
JER|8|20|"The harvest is past, the summer has ended, and we are not saved."
JER|8|21|Since my people are crushed, I am crushed; I mourn, and horror grips me.
JER|8|22|Is there no balm in Gilead? Is there no physician there? Why then is there no healing for the wound of my people?
JER|9|1|Oh, that my head were a spring of water and my eyes a fountain of tears! I would weep day and night for the slain of my people.
JER|9|2|Oh, that I had in the desert a lodging place for travelers, so that I might leave my people and go away from them; for they are all adulterers, a crowd of unfaithful people.
JER|9|3|"They make ready their tongue like a bow, to shoot lies; it is not by truth that they triumph in the land. They go from one sin to another; they do not acknowledge me," declares the LORD.
JER|9|4|"Beware of your friends; do not trust your brothers. For every brother is a deceiver, and every friend a slanderer.
JER|9|5|Friend deceives friend, and no one speaks the truth. They have taught their tongues to lie; they weary themselves with sinning.
JER|9|6|You live in the midst of deception; in their deceit they refuse to acknowledge me," declares the LORD.
JER|9|7|Therefore this is what the LORD Almighty says: "See, I will refine and test them, for what else can I do because of the sin of my people?
JER|9|8|Their tongue is a deadly arrow; it speaks with deceit. With his mouth each speaks cordially to his neighbor, but in his heart he sets a trap for him.
JER|9|9|Should I not punish them for this?" declares the LORD. "Should I not avenge myself on such a nation as this?"
JER|9|10|I will weep and wail for the mountains and take up a lament concerning the desert pastures. They are desolate and untraveled, and the lowing of cattle is not heard. The birds of the air have fled and the animals are gone.
JER|9|11|"I will make Jerusalem a heap of ruins, a haunt of jackals; and I will lay waste the towns of Judah so no one can live there."
JER|9|12|What man is wise enough to understand this? Who has been instructed by the LORD and can explain it? Why has the land been ruined and laid waste like a desert that no one can cross?
JER|9|13|The LORD said, "It is because they have forsaken my law, which I set before them; they have not obeyed me or followed my law.
JER|9|14|Instead, they have followed the stubbornness of their hearts; they have followed the Baals, as their fathers taught them."
JER|9|15|Therefore, this is what the LORD Almighty, the God of Israel, says: "See, I will make this people eat bitter food and drink poisoned water.
JER|9|16|I will scatter them among nations that neither they nor their fathers have known, and I will pursue them with the sword until I have destroyed them."
JER|9|17|This is what the LORD Almighty says: "Consider now! Call for the wailing women to come; send for the most skillful of them.
JER|9|18|Let them come quickly and wail over us till our eyes overflow with tears and water streams from our eyelids.
JER|9|19|The sound of wailing is heard from Zion: 'How ruined we are! How great is our shame! We must leave our land because our houses are in ruins.'"
JER|9|20|Now, O women, hear the word of the LORD; open your ears to the words of his mouth. Teach your daughters how to wail; teach one another a lament.
JER|9|21|Death has climbed in through our windows and has entered our fortresses; it has cut off the children from the streets and the young men from the public squares.
JER|9|22|Say, "This is what the LORD declares: "'The dead bodies of men will lie like refuse on the open field, like cut grain behind the reaper, with no one to gather them.'"
JER|9|23|This is what the LORD says: "Let not the wise man boast of his wisdom or the strong man boast of his strength or the rich man boast of his riches,
JER|9|24|but let him who boasts boast about this: that he understands and knows me, that I am the LORD, who exercises kindness, justice and righteousness on earth, for in these I delight," declares the LORD.
JER|9|25|"The days are coming," declares the LORD, "when I will punish all who are circumcised only in the flesh-
JER|9|26|Egypt, Judah, Edom, Ammon, Moab and all who live in the desert in distant places. For all these nations are really uncircumcised, and even the whole house of Israel is uncircumcised in heart."
JER|10|1|Hear what the LORD says to you, O house of Israel.
JER|10|2|This is what the LORD says: "Do not learn the ways of the nations or be terrified by signs in the sky, though the nations are terrified by them.
JER|10|3|For the customs of the peoples are worthless; they cut a tree out of the forest, and a craftsman shapes it with his chisel.
JER|10|4|They adorn it with silver and gold; they fasten it with hammer and nails so it will not totter.
JER|10|5|Like a scarecrow in a melon patch, their idols cannot speak; they must be carried because they cannot walk. Do not fear them; they can do no harm nor can they do any good."
JER|10|6|No one is like you, O LORD; you are great, and your name is mighty in power.
JER|10|7|Who should not revere you, O King of the nations? This is your due. Among all the wise men of the nations and in all their kingdoms, there is no one like you.
JER|10|8|They are all senseless and foolish; they are taught by worthless wooden idols.
JER|10|9|Hammered silver is brought from Tarshish and gold from Uphaz. What the craftsman and goldsmith have made is then dressed in blue and purple- all made by skilled workers.
JER|10|10|But the LORD is the true God; he is the living God, the eternal King. When he is angry, the earth trembles; the nations cannot endure his wrath.
JER|10|11|"Tell them this: 'These gods, who did not make the heavens and the earth, will perish from the earth and from under the heavens.'"
JER|10|12|But God made the earth by his power; he founded the world by his wisdom and stretched out the heavens by his understanding.
JER|10|13|When he thunders, the waters in the heavens roar; he makes clouds rise from the ends of the earth. He sends lightning with the rain and brings out the wind from his storehouses.
JER|10|14|Everyone is senseless and without knowledge; every goldsmith is shamed by his idols. His images are a fraud; they have no breath in them.
JER|10|15|They are worthless, the objects of mockery; when their judgment comes, they will perish.
JER|10|16|He who is the Portion of Jacob is not like these, for he is the Maker of all things, including Israel, the tribe of his inheritance- the LORD Almighty is his name.
JER|10|17|Gather up your belongings to leave the land, you who live under siege.
JER|10|18|For this is what the LORD says: "At this time I will hurl out those who live in this land; I will bring distress on them so that they may be captured."
JER|10|19|Woe to me because of my injury! My wound is incurable! Yet I said to myself, "This is my sickness, and I must endure it."
JER|10|20|My tent is destroyed; all its ropes are snapped. My sons are gone from me and are no more; no one is left now to pitch my tent or to set up my shelter.
JER|10|21|The shepherds are senseless and do not inquire of the LORD; so they do not prosper and all their flock is scattered.
JER|10|22|Listen! The report is coming- a great commotion from the land of the north! It will make the towns of Judah desolate, a haunt of jackals.
JER|10|23|I know, O LORD, that a man's life is not his own; it is not for man to direct his steps.
JER|10|24|Correct me, LORD, but only with justice- not in your anger, lest you reduce me to nothing.
JER|10|25|Pour out your wrath on the nations that do not acknowledge you, on the peoples who do not call on your name. For they have devoured Jacob; they have devoured him completely and destroyed his homeland.
JER|11|1|This is the word that came to Jeremiah from the LORD:
JER|11|2|"Listen to the terms of this covenant and tell them to the people of Judah and to those who live in Jerusalem.
JER|11|3|Tell them that this is what the LORD, the God of Israel, says: 'Cursed is the man who does not obey the terms of this covenant-
JER|11|4|the terms I commanded your forefathers when I brought them out of Egypt, out of the iron-smelting furnace.' I said, 'Obey me and do everything I command you, and you will be my people, and I will be your God.
JER|11|5|Then I will fulfill the oath I swore to your forefathers, to give them a land flowing with milk and honey'-the land you possess today." I answered, "Amen, LORD."
JER|11|6|The LORD said to me, "Proclaim all these words in the towns of Judah and in the streets of Jerusalem: 'Listen to the terms of this covenant and follow them.
JER|11|7|From the time I brought your forefathers up from Egypt until today, I warned them again and again, saying, "Obey me."
JER|11|8|But they did not listen or pay attention; instead, they followed the stubbornness of their evil hearts. So I brought on them all the curses of the covenant I had commanded them to follow but that they did not keep.'"
JER|11|9|Then the LORD said to me, "There is a conspiracy among the people of Judah and those who live in Jerusalem.
JER|11|10|They have returned to the sins of their forefathers, who refused to listen to my words. They have followed other gods to serve them. Both the house of Israel and the house of Judah have broken the covenant I made with their forefathers.
JER|11|11|Therefore this is what the LORD says: 'I will bring on them a disaster they cannot escape. Although they cry out to me, I will not listen to them.
JER|11|12|The towns of Judah and the people of Jerusalem will go and cry out to the gods to whom they burn incense, but they will not help them at all when disaster strikes.
JER|11|13|You have as many gods as you have towns, O Judah; and the altars you have set up to burn incense to that shameful god Baal are as many as the streets of Jerusalem.'
JER|11|14|"Do not pray for this people nor offer any plea or petition for them, because I will not listen when they call to me in the time of their distress.
JER|11|15|"What is my beloved doing in my temple as she works out her evil schemes with many? Can consecrated meat avert your punishment? When you engage in your wickedness, then you rejoice. "
JER|11|16|The LORD called you a thriving olive tree with fruit beautiful in form. But with the roar of a mighty storm he will set it on fire, and its branches will be broken.
JER|11|17|The LORD Almighty, who planted you, has decreed disaster for you, because the house of Israel and the house of Judah have done evil and provoked me to anger by burning incense to Baal.
JER|11|18|Because the LORD revealed their plot to me, I knew it, for at that time he showed me what they were doing.
JER|11|19|I had been like a gentle lamb led to the slaughter; I did not realize that they had plotted against me, saying, "Let us destroy the tree and its fruit; let us cut him off from the land of the living, that his name be remembered no more."
JER|11|20|But, O LORD Almighty, you who judge righteously and test the heart and mind, let me see your vengeance upon them, for to you I have committed my cause.
JER|11|21|"Therefore this is what the LORD says about the men of Anathoth who are seeking your life and saying, 'Do not prophesy in the name of the LORD or you will die by our hands'-
JER|11|22|therefore this is what the LORD Almighty says: 'I will punish them. Their young men will die by the sword, their sons and daughters by famine.
JER|11|23|Not even a remnant will be left to them, because I will bring disaster on the men of Anathoth in the year of their punishment.'"
JER|12|1|You are always righteous, O LORD, when I bring a case before you. Yet I would speak with you about your justice: Why does the way of the wicked prosper? Why do all the faithless live at ease?
JER|12|2|You have planted them, and they have taken root; they grow and bear fruit. You are always on their lips but far from their hearts.
JER|12|3|Yet you know me, O LORD; you see me and test my thoughts about you. Drag them off like sheep to be butchered! Set them apart for the day of slaughter!
JER|12|4|How long will the land lie parched and the grass in every field be withered? Because those who live in it are wicked, the animals and birds have perished. Moreover, the people are saying, "He will not see what happens to us."
JER|12|5|"If you have raced with men on foot and they have worn you out, how can you compete with horses? If you stumble in safe country, how will you manage in the thickets by the Jordan?
JER|12|6|Your brothers, your own family- even they have betrayed you; they have raised a loud cry against you. Do not trust them, though they speak well of you.
JER|12|7|"I will forsake my house, abandon my inheritance; I will give the one I love into the hands of her enemies.
JER|12|8|My inheritance has become to me like a lion in the forest. She roars at me; therefore I hate her.
JER|12|9|Has not my inheritance become to me like a speckled bird of prey that other birds of prey surround and attack? Go and gather all the wild beasts; bring them to devour.
JER|12|10|Many shepherds will ruin my vineyard and trample down my field; they will turn my pleasant field into a desolate wasteland.
JER|12|11|It will be made a wasteland, parched and desolate before me; the whole land will be laid waste because there is no one who cares.
JER|12|12|Over all the barren heights in the desert destroyers will swarm, for the sword of the LORD will devour from one end of the land to the other; no one will be safe.
JER|12|13|They will sow wheat but reap thorns; they will wear themselves out but gain nothing. So bear the shame of your harvest because of the LORD's fierce anger."
JER|12|14|This is what the LORD says: "As for all my wicked neighbors who seize the inheritance I gave my people Israel, I will uproot them from their lands and I will uproot the house of Judah from among them.
JER|12|15|But after I uproot them, I will again have compassion and will bring each of them back to his own inheritance and his own country.
JER|12|16|And if they learn well the ways of my people and swear by my name, saying, 'As surely as the LORD lives'-even as they once taught my people to swear by Baal-then they will be established among my people.
JER|12|17|But if any nation does not listen, I will completely uproot and destroy it," declares the LORD.
JER|13|1|This is what the LORD said to me: "Go and buy a linen belt and put it around your waist, but do not let it touch water."
JER|13|2|So I bought a belt, as the LORD directed, and put it around my waist.
JER|13|3|Then the word of the LORD came to me a second time:
JER|13|4|"Take the belt you bought and are wearing around your waist, and go now to Perath and hide it there in a crevice in the rocks."
JER|13|5|So I went and hid it at Perath, as the LORD told me.
JER|13|6|Many days later the LORD said to me, "Go now to Perath and get the belt I told you to hide there."
JER|13|7|So I went to Perath and dug up the belt and took it from the place where I had hidden it, but now it was ruined and completely useless.
JER|13|8|Then the word of the LORD came to me:
JER|13|9|"This is what the LORD says: 'In the same way I will ruin the pride of Judah and the great pride of Jerusalem.
JER|13|10|These wicked people, who refuse to listen to my words, who follow the stubbornness of their hearts and go after other gods to serve and worship them, will be like this belt-completely useless!
JER|13|11|For as a belt is bound around a man's waist, so I bound the whole house of Israel and the whole house of Judah to me,' declares the LORD, 'to be my people for my renown and praise and honor. But they have not listened.'
JER|13|12|"Say to them: 'This is what the LORD, the God of Israel, says: Every wineskin should be filled with wine.' And if they say to you, 'Don't we know that every wineskin should be filled with wine?'
JER|13|13|then tell them, 'This is what the LORD says: I am going to fill with drunkenness all who live in this land, including the kings who sit on David's throne, the priests, the prophets and all those living in Jerusalem.
JER|13|14|I will smash them one against the other, fathers and sons alike, declares the LORD. I will allow no pity or mercy or compassion to keep me from destroying them.'"
JER|13|15|Hear and pay attention, do not be arrogant, for the LORD has spoken.
JER|13|16|Give glory to the LORD your God before he brings the darkness, before your feet stumble on the darkening hills. You hope for light, but he will turn it to thick darkness and change it to deep gloom.
JER|13|17|But if you do not listen, I will weep in secret because of your pride; my eyes will weep bitterly, overflowing with tears, because the LORD's flock will be taken captive.
JER|13|18|Say to the king and to the queen mother, "Come down from your thrones, for your glorious crowns will fall from your heads."
JER|13|19|The cities in the Negev will be shut up, and there will be no one to open them. All Judah will be carried into exile, carried completely away.
JER|13|20|Lift up your eyes and see those who are coming from the north. Where is the flock that was entrusted to you, the sheep of which you boasted?
JER|13|21|What will you say when the LORD sets over you those you cultivated as your special allies? Will not pain grip you like that of a woman in labor?
JER|13|22|And if you ask yourself, "Why has this happened to me?"- it is because of your many sins that your skirts have been torn off and your body mistreated.
JER|13|23|Can the Ethiopian change his skin or the leopard its spots? Neither can you do good who are accustomed to doing evil.
JER|13|24|"I will scatter you like chaff driven by the desert wind.
JER|13|25|This is your lot, the portion I have decreed for you," declares the LORD, "because you have forgotten me and trusted in false gods.
JER|13|26|I will pull up your skirts over your face that your shame may be seen-
JER|13|27|your adulteries and lustful neighings, your shameless prostitution! I have seen your detestable acts on the hills and in the fields. Woe to you, O Jerusalem! How long will you be unclean?"
JER|14|1|This is the word of the LORD to Jeremiah concerning the drought:
JER|14|2|"Judah mourns, her cities languish; they wail for the land, and a cry goes up from Jerusalem.
JER|14|3|The nobles send their servants for water; they go to the cisterns but find no water. They return with their jars unfilled; dismayed and despairing, they cover their heads.
JER|14|4|The ground is cracked because there is no rain in the land; the farmers are dismayed and cover their heads.
JER|14|5|Even the doe in the field deserts her newborn fawn because there is no grass.
JER|14|6|Wild donkeys stand on the barren heights and pant like jackals; their eyesight fails for lack of pasture."
JER|14|7|Although our sins testify against us, O LORD, do something for the sake of your name. For our backsliding is great; we have sinned against you.
JER|14|8|O Hope of Israel, its Savior in times of distress, why are you like a stranger in the land, like a traveler who stays only a night?
JER|14|9|Why are you like a man taken by surprise, like a warrior powerless to save? You are among us, O LORD, and we bear your name; do not forsake us!
JER|14|10|This is what the LORD says about this people: "They greatly love to wander; they do not restrain their feet. So the LORD does not accept them; he will now remember their wickedness and punish them for their sins."
JER|14|11|Then the LORD said to me, "Do not pray for the well-being of this people.
JER|14|12|Although they fast, I will not listen to their cry; though they offer burnt offerings and grain offerings, I will not accept them. Instead, I will destroy them with the sword, famine and plague."
JER|14|13|But I said, "Ah, Sovereign LORD, the prophets keep telling them, 'You will not see the sword or suffer famine. Indeed, I will give you lasting peace in this place.'"
JER|14|14|Then the LORD said to me, "The prophets are prophesying lies in my name. I have not sent them or appointed them or spoken to them. They are prophesying to you false visions, divinations, idolatries and the delusions of their own minds.
JER|14|15|Therefore, this is what the LORD says about the prophets who are prophesying in my name: I did not send them, yet they are saying, 'No sword or famine will touch this land.' Those same prophets will perish by sword and famine.
JER|14|16|And the people they are prophesying to will be thrown out into the streets of Jerusalem because of the famine and sword. There will be no one to bury them or their wives, their sons or their daughters. I will pour out on them the calamity they deserve.
JER|14|17|"Speak this word to them: "'Let my eyes overflow with tears night and day without ceasing; for my virgin daughter-my people- has suffered a grievous wound, a crushing blow.
JER|14|18|If I go into the country, I see those slain by the sword; if I go into the city, I see the ravages of famine. Both prophet and priest have gone to a land they know not.'"
JER|14|19|Have you rejected Judah completely? Do you despise Zion? Why have you afflicted us so that we cannot be healed? We hoped for peace but no good has come, for a time of healing but there is only terror.
JER|14|20|O LORD, we acknowledge our wickedness and the guilt of our fathers; we have indeed sinned against you.
JER|14|21|For the sake of your name do not despise us; do not dishonor your glorious throne. Remember your covenant with us and do not break it.
JER|14|22|Do any of the worthless idols of the nations bring rain? Do the skies themselves send down showers? No, it is you, O LORD our God. Therefore our hope is in you, for you are the one who does all this.
JER|15|1|Then the LORD said to me: "Even if Moses and Samuel were to stand before me, my heart would not go out to this people. Send them away from my presence! Let them go!
JER|15|2|And if they ask you, 'Where shall we go?' tell them, 'This is what the LORD says: "'Those destined for death, to death; those for the sword, to the sword; those for starvation, to starvation; those for captivity, to captivity.'
JER|15|3|"I will send four kinds of destroyers against them," declares the LORD, "the sword to kill and the dogs to drag away and the birds of the air and the beasts of the earth to devour and destroy.
JER|15|4|I will make them abhorrent to all the kingdoms of the earth because of what Manasseh son of Hezekiah king of Judah did in Jerusalem.
JER|15|5|"Who will have pity on you, O Jerusalem? Who will mourn for you? Who will stop to ask how you are?
JER|15|6|You have rejected me," declares the LORD. "You keep on backsliding. So I will lay hands on you and destroy you; I can no longer show compassion.
JER|15|7|I will winnow them with a winnowing fork at the city gates of the land. I will bring bereavement and destruction on my people, for they have not changed their ways.
JER|15|8|I will make their widows more numerous than the sand of the sea. At midday I will bring a destroyer against the mothers of their young men; suddenly I will bring down on them anguish and terror.
JER|15|9|The mother of seven will grow faint and breathe her last. Her sun will set while it is still day; she will be disgraced and humiliated. I will put the survivors to the sword before their enemies," declares the LORD.
JER|15|10|Alas, my mother, that you gave me birth, a man with whom the whole land strives and contends! I have neither lent nor borrowed, yet everyone curses me.
JER|15|11|The LORD said, "Surely I will deliver you for a good purpose; surely I will make your enemies plead with you in times of disaster and times of distress.
JER|15|12|"Can a man break iron- iron from the north-or bronze?
JER|15|13|Your wealth and your treasures I will give as plunder, without charge, because of all your sins throughout your country.
JER|15|14|I will enslave you to your enemies in a land you do not know, for my anger will kindle a fire that will burn against you."
JER|15|15|You understand, O LORD; remember me and care for me. Avenge me on my persecutors. You are long-suffering-do not take me away; think of how I suffer reproach for your sake.
JER|15|16|When your words came, I ate them; they were my joy and my heart's delight, for I bear your name, O LORD God Almighty.
JER|15|17|I never sat in the company of revelers, never made merry with them; I sat alone because your hand was on me and you had filled me with indignation.
JER|15|18|Why is my pain unending and my wound grievous and incurable? Will you be to me like a deceptive brook, like a spring that fails?
JER|15|19|Therefore this is what the LORD says: "If you repent, I will restore you that you may serve me; if you utter worthy, not worthless, words, you will be my spokesman. Let this people turn to you, but you must not turn to them.
JER|15|20|I will make you a wall to this people, a fortified wall of bronze; they will fight against you but will not overcome you, for I am with you to rescue and save you," declares the LORD.
JER|15|21|"I will save you from the hands of the wicked and redeem you from the grasp of the cruel."
JER|16|1|Then the word of the LORD came to me:
JER|16|2|"You must not marry and have sons or daughters in this place."
JER|16|3|For this is what the LORD says about the sons and daughters born in this land and about the women who are their mothers and the men who are their fathers:
JER|16|4|"They will die of deadly diseases. They will not be mourned or buried but will be like refuse lying on the ground. They will perish by sword and famine, and their dead bodies will become food for the birds of the air and the beasts of the earth."
JER|16|5|For this is what the LORD says: "Do not enter a house where there is a funeral meal; do not go to mourn or show sympathy, because I have withdrawn my blessing, my love and my pity from this people," declares the LORD.
JER|16|6|"Both high and low will die in this land. They will not be buried or mourned, and no one will cut himself or shave his head for them.
JER|16|7|No one will offer food to comfort those who mourn for the dead-not even for a father or a mother-nor will anyone give them a drink to console them.
JER|16|8|"And do not enter a house where there is feasting and sit down to eat and drink.
JER|16|9|For this is what the LORD Almighty, the God of Israel, says: Before your eyes and in your days I will bring an end to the sounds of joy and gladness and to the voices of bride and bridegroom in this place.
JER|16|10|"When you tell these people all this and they ask you, 'Why has the LORD decreed such a great disaster against us? What wrong have we done? What sin have we committed against the LORD our God?'
JER|16|11|then say to them, 'It is because your fathers forsook me,' declares the LORD, 'and followed other gods and served and worshiped them. They forsook me and did not keep my law.
JER|16|12|But you have behaved more wickedly than your fathers. See how each of you is following the stubbornness of his evil heart instead of obeying me.
JER|16|13|So I will throw you out of this land into a land neither you nor your fathers have known, and there you will serve other gods day and night, for I will show you no favor.'
JER|16|14|"However, the days are coming," declares the LORD, "when men will no longer say, 'As surely as the LORD lives, who brought the Israelites up out of Egypt,'
JER|16|15|but they will say, 'As surely as the LORD lives, who brought the Israelites up out of the land of the north and out of all the countries where he had banished them.' For I will restore them to the land I gave their forefathers.
JER|16|16|"But now I will send for many fishermen," declares the LORD, "and they will catch them. After that I will send for many hunters, and they will hunt them down on every mountain and hill and from the crevices of the rocks.
JER|16|17|My eyes are on all their ways; they are not hidden from me, nor is their sin concealed from my eyes.
JER|16|18|I will repay them double for their wickedness and their sin, because they have defiled my land with the lifeless forms of their vile images and have filled my inheritance with their detestable idols."
JER|16|19|O LORD, my strength and my fortress, my refuge in time of distress, to you the nations will come from the ends of the earth and say, "Our fathers possessed nothing but false gods, worthless idols that did them no good.
JER|16|20|Do men make their own gods? Yes, but they are not gods!"
JER|16|21|"Therefore I will teach them- this time I will teach them my power and might. Then they will know that my name is the LORD.
JER|17|1|"Judah's sin is engraved with an iron tool, inscribed with a flint point, on the tablets of their hearts and on the horns of their altars.
JER|17|2|Even their children remember their altars and Asherah poles beside the spreading trees and on the high hills.
JER|17|3|My mountain in the land and your wealth and all your treasures I will give away as plunder, together with your high places, because of sin throughout your country.
JER|17|4|Through your own fault you will lose the inheritance I gave you. I will enslave you to your enemies in a land you do not know, for you have kindled my anger, and it will burn forever."
JER|17|5|This is what the LORD says: "Cursed is the one who trusts in man, who depends on flesh for his strength and whose heart turns away from the LORD.
JER|17|6|He will be like a bush in the wastelands; he will not see prosperity when it comes. He will dwell in the parched places of the desert, in a salt land where no one lives.
JER|17|7|"But blessed is the man who trusts in the LORD, whose confidence is in him.
JER|17|8|He will be like a tree planted by the water that sends out its roots by the stream. It does not fear when heat comes; its leaves are always green. It has no worries in a year of drought and never fails to bear fruit."
JER|17|9|The heart is deceitful above all things and beyond cure. Who can understand it?
JER|17|10|"I the LORD search the heart and examine the mind, to reward a man according to his conduct, according to what his deeds deserve."
JER|17|11|Like a partridge that hatches eggs it did not lay is the man who gains riches by unjust means. When his life is half gone, they will desert him, and in the end he will prove to be a fool.
JER|17|12|A glorious throne, exalted from the beginning, is the place of our sanctuary.
JER|17|13|O LORD, the hope of Israel, all who forsake you will be put to shame. Those who turn away from you will be written in the dust because they have forsaken the LORD, the spring of living water.
JER|17|14|Heal me, O LORD, and I will be healed; save me and I will be saved, for you are the one I praise.
JER|17|15|They keep saying to me, "Where is the word of the LORD? Let it now be fulfilled!"
JER|17|16|I have not run away from being your shepherd; you know I have not desired the day of despair. What passes my lips is open before you.
JER|17|17|Do not be a terror to me; you are my refuge in the day of disaster.
JER|17|18|Let my persecutors be put to shame, but keep me from shame; let them be terrified, but keep me from terror. Bring on them the day of disaster; destroy them with double destruction.
JER|17|19|This is what the LORD said to me: "Go and stand at the gate of the people, through which the kings of Judah go in and out; stand also at all the other gates of Jerusalem.
JER|17|20|Say to them, 'Hear the word of the LORD, O kings of Judah and all people of Judah and everyone living in Jerusalem who come through these gates.
JER|17|21|This is what the LORD says: Be careful not to carry a load on the Sabbath day or bring it through the gates of Jerusalem.
JER|17|22|Do not bring a load out of your houses or do any work on the Sabbath, but keep the Sabbath day holy, as I commanded your forefathers.
JER|17|23|Yet they did not listen or pay attention; they were stiff-necked and would not listen or respond to discipline.
JER|17|24|But if you are careful to obey me, declares the LORD, and bring no load through the gates of this city on the Sabbath, but keep the Sabbath day holy by not doing any work on it,
JER|17|25|then kings who sit on David's throne will come through the gates of this city with their officials. They and their officials will come riding in chariots and on horses, accompanied by the men of Judah and those living in Jerusalem, and this city will be inhabited forever.
JER|17|26|People will come from the towns of Judah and the villages around Jerusalem, from the territory of Benjamin and the western foothills, from the hill country and the Negev, bringing burnt offerings and sacrifices, grain offerings, incense and thank offerings to the house of the LORD.
JER|17|27|But if you do not obey me to keep the Sabbath day holy by not carrying any load as you come through the gates of Jerusalem on the Sabbath day, then I will kindle an unquenchable fire in the gates of Jerusalem that will consume her fortresses.'"
JER|18|1|This is the word that came to Jeremiah from the LORD:
JER|18|2|"Go down to the potter's house, and there I will give you my message."
JER|18|3|So I went down to the potter's house, and I saw him working at the wheel.
JER|18|4|But the pot he was shaping from the clay was marred in his hands; so the potter formed it into another pot, shaping it as seemed best to him.
JER|18|5|Then the word of the LORD came to me:
JER|18|6|"O house of Israel, can I not do with you as this potter does?" declares the LORD. "Like clay in the hand of the potter, so are you in my hand, O house of Israel.
JER|18|7|If at any time I announce that a nation or kingdom is to be uprooted, torn down and destroyed,
JER|18|8|and if that nation I warned repents of its evil, then I will relent and not inflict on it the disaster I had planned.
JER|18|9|And if at another time I announce that a nation or kingdom is to be built up and planted,
JER|18|10|and if it does evil in my sight and does not obey me, then I will reconsider the good I had intended to do for it.
JER|18|11|"Now therefore say to the people of Judah and those living in Jerusalem, 'This is what the LORD says: Look! I am preparing a disaster for you and devising a plan against you. So turn from your evil ways, each one of you, and reform your ways and your actions.'
JER|18|12|But they will reply, 'It's no use. We will continue with our own plans; each of us will follow the stubbornness of his evil heart.'"
JER|18|13|Therefore this is what the LORD says: "Inquire among the nations: Who has ever heard anything like this? A most horrible thing has been done by Virgin Israel.
JER|18|14|Does the snow of Lebanon ever vanish from its rocky slopes? Do its cool waters from distant sources ever cease to flow?
JER|18|15|Yet my people have forgotten me; they burn incense to worthless idols, which made them stumble in their ways and in the ancient paths. They made them walk in bypaths and on roads not built up.
JER|18|16|Their land will be laid waste, an object of lasting scorn; all who pass by will be appalled and will shake their heads.
JER|18|17|Like a wind from the east, I will scatter them before their enemies; I will show them my back and not my face in the day of their disaster."
JER|18|18|They said, "Come, let's make plans against Jeremiah; for the teaching of the law by the priest will not be lost, nor will counsel from the wise, nor the word from the prophets. So come, let's attack him with our tongues and pay no attention to anything he says."
JER|18|19|Listen to me, O LORD; hear what my accusers are saying!
JER|18|20|Should good be repaid with evil? Yet they have dug a pit for me. Remember that I stood before you and spoke in their behalf to turn your wrath away from them.
JER|18|21|So give their children over to famine; hand them over to the power of the sword. Let their wives be made childless and widows; let their men be put to death, their young men slain by the sword in battle.
JER|18|22|Let a cry be heard from their houses when you suddenly bring invaders against them, for they have dug a pit to capture me and have hidden snares for my feet.
JER|18|23|But you know, O LORD, all their plots to kill me. Do not forgive their crimes or blot out their sins from your sight. Let them be overthrown before you; deal with them in the time of your anger.
JER|19|1|This is what the LORD says: "Go and buy a clay jar from a potter. Take along some of the elders of the people and of the priests
JER|19|2|and go out to the Valley of Ben Hinnom, near the entrance of the Potsherd Gate. There proclaim the words I tell you,
JER|19|3|and say, 'Hear the word of the LORD, O kings of Judah and people of Jerusalem. This is what the LORD Almighty, the God of Israel, says: Listen! I am going to bring a disaster on this place that will make the ears of everyone who hears of it tingle.
JER|19|4|For they have forsaken me and made this a place of foreign gods; they have burned sacrifices in it to gods that neither they nor their fathers nor the kings of Judah ever knew, and they have filled this place with the blood of the innocent.
JER|19|5|They have built the high places of Baal to burn their sons in the fire as offerings to Baal-something I did not command or mention, nor did it enter my mind.
JER|19|6|So beware, the days are coming, declares the LORD, when people will no longer call this place Topheth or the Valley of Ben Hinnom, but the Valley of Slaughter.
JER|19|7|"'In this place I will ruin the plans of Judah and Jerusalem. I will make them fall by the sword before their enemies, at the hands of those who seek their lives, and I will give their carcasses as food to the birds of the air and the beasts of the earth.
JER|19|8|I will devastate this city and make it an object of scorn; all who pass by will be appalled and will scoff because of all its wounds.
JER|19|9|I will make them eat the flesh of their sons and daughters, and they will eat one another's flesh during the stress of the siege imposed on them by the enemies who seek their lives.'
JER|19|10|"Then break the jar while those who go with you are watching,
JER|19|11|and say to them, 'This is what the LORD Almighty says: I will smash this nation and this city just as this potter's jar is smashed and cannot be repaired. They will bury the dead in Topheth until there is no more room.
JER|19|12|This is what I will do to this place and to those who live here, declares the LORD. I will make this city like Topheth.
JER|19|13|The houses in Jerusalem and those of the kings of Judah will be defiled like this place, Topheth-all the houses where they burned incense on the roofs to all the starry hosts and poured out drink offerings to other gods.'"
JER|19|14|Jeremiah then returned from Topheth, where the LORD had sent him to prophesy, and stood in the court of the LORD's temple and said to all the people,
JER|19|15|"This is what the LORD Almighty, the God of Israel, says: 'Listen! I am going to bring on this city and the villages around it every disaster I pronounced against them, because they were stiff-necked and would not listen to my words.'"
JER|20|1|When the priest Pashhur son of Immer, the chief officer in the temple of the LORD, heard Jeremiah prophesying these things,
JER|20|2|he had Jeremiah the prophet beaten and put in the stocks at the Upper Gate of Benjamin at the LORD's temple.
JER|20|3|The next day, when Pashhur released him from the stocks, Jeremiah said to him, "The LORD's name for you is not Pashhur, but Magor-Missabib.
JER|20|4|For this is what the LORD says: 'I will make you a terror to yourself and to all your friends; with your own eyes you will see them fall by the sword of their enemies. I will hand all Judah over to the king of Babylon, who will carry them away to Babylon or put them to the sword.
JER|20|5|I will hand over to their enemies all the wealth of this city-all its products, all its valuables and all the treasures of the kings of Judah. They will take it away as plunder and carry it off to Babylon.
JER|20|6|And you, Pashhur, and all who live in your house will go into exile to Babylon. There you will die and be buried, you and all your friends to whom you have prophesied lies.'"
JER|20|7|O LORD, you deceived me, and I was deceived; you overpowered me and prevailed. I am ridiculed all day long; everyone mocks me.
JER|20|8|Whenever I speak, I cry out proclaiming violence and destruction. So the word of the LORD has brought me insult and reproach all day long.
JER|20|9|But if I say, "I will not mention him or speak any more in his name," his word is in my heart like a fire, a fire shut up in my bones. I am weary of holding it in; indeed, I cannot.
JER|20|10|I hear many whispering, "Terror on every side! Report him! Let's report him!" All my friends are waiting for me to slip, saying, "Perhaps he will be deceived; then we will prevail over him and take our revenge on him."
JER|20|11|But the LORD is with me like a mighty warrior; so my persecutors will stumble and not prevail. They will fail and be thoroughly disgraced; their dishonor will never be forgotten.
JER|20|12|O LORD Almighty, you who examine the righteous and probe the heart and mind, let me see your vengeance upon them, for to you I have committed my cause.
JER|20|13|Sing to the LORD! Give praise to the LORD! He rescues the life of the needy from the hands of the wicked.
JER|20|14|Cursed be the day I was born! May the day my mother bore me not be blessed!
JER|20|15|Cursed be the man who brought my father the news, who made him very glad, saying, "A child is born to you-a son!"
JER|20|16|May that man be like the towns the LORD overthrew without pity. May he hear wailing in the morning, a battle cry at noon.
JER|20|17|For he did not kill me in the womb, with my mother as my grave, her womb enlarged forever.
JER|20|18|Why did I ever come out of the womb to see trouble and sorrow and to end my days in shame?
JER|21|1|The word came to Jeremiah from the LORD when King Zedekiah sent to him Pashhur son of Malkijah and the priest Zephaniah son of Maaseiah. They said:
JER|21|2|"Inquire now of the LORD for us because Nebuchadnezzar king of Babylon is attacking us. Perhaps the LORD will perform wonders for us as in times past so that he will withdraw from us."
JER|21|3|But Jeremiah answered them, "Tell Zedekiah,
JER|21|4|'This is what the LORD, the God of Israel, says: I am about to turn against you the weapons of war that are in your hands, which you are using to fight the king of Babylon and the Babylonians who are outside the wall besieging you. And I will gather them inside this city.
JER|21|5|I myself will fight against you with an outstretched hand and a mighty arm in anger and fury and great wrath.
JER|21|6|I will strike down those who live in this city-both men and animals-and they will die of a terrible plague.
JER|21|7|After that, declares the LORD, I will hand over Zedekiah king of Judah, his officials and the people in this city who survive the plague, sword and famine, to Nebuchadnezzar king of Babylon and to their enemies who seek their lives. He will put them to the sword; he will show them no mercy or pity or compassion.'
JER|21|8|"Furthermore, tell the people, 'This is what the LORD says: See, I am setting before you the way of life and the way of death.
JER|21|9|Whoever stays in this city will die by the sword, famine or plague. But whoever goes out and surrenders to the Babylonians who are besieging you will live; he will escape with his life.
JER|21|10|I have determined to do this city harm and not good, declares the LORD. It will be given into the hands of the king of Babylon, and he will destroy it with fire.'
JER|21|11|"Moreover, say to the royal house of Judah, 'Hear the word of the LORD;
JER|21|12|O house of David, this is what the LORD says: "'Administer justice every morning; rescue from the hand of his oppressor the one who has been robbed, or my wrath will break out and burn like fire because of the evil you have done- burn with no one to quench it.
JER|21|13|I am against you, Jerusalem, you who live above this valley on the rocky plateau, declares the LORD - you who say, "Who can come against us? Who can enter our refuge?"
JER|21|14|I will punish you as your deeds deserve, declares the LORD. I will kindle a fire in your forests that will consume everything around you.'"
JER|22|1|This is what the LORD says: "Go down to the palace of the king of Judah and proclaim this message there:
JER|22|2|'Hear the word of the LORD, O king of Judah, you who sit on David's throne-you, your officials and your people who come through these gates.
JER|22|3|This is what the LORD says: Do what is just and right. Rescue from the hand of his oppressor the one who has been robbed. Do no wrong or violence to the alien, the fatherless or the widow, and do not shed innocent blood in this place.
JER|22|4|For if you are careful to carry out these commands, then kings who sit on David's throne will come through the gates of this palace, riding in chariots and on horses, accompanied by their officials and their people.
JER|22|5|But if you do not obey these commands, declares the LORD, I swear by myself that this palace will become a ruin.'"
JER|22|6|For this is what the LORD says about the palace of the king of Judah: "Though you are like Gilead to me, like the summit of Lebanon, I will surely make you like a desert, like towns not inhabited.
JER|22|7|I will send destroyers against you, each man with his weapons, and they will cut up your fine cedar beams and throw them into the fire.
JER|22|8|"People from many nations will pass by this city and will ask one another, 'Why has the LORD done such a thing to this great city?'
JER|22|9|And the answer will be: 'Because they have forsaken the covenant of the LORD their God and have worshiped and served other gods.'"
JER|22|10|Do not weep for the dead king or mourn his loss; rather, weep bitterly for him who is exiled, because he will never return nor see his native land again.
JER|22|11|For this is what the LORD says about Shallum son of Josiah, who succeeded his father as king of Judah but has gone from this place: "He will never return.
JER|22|12|He will die in the place where they have led him captive; he will not see this land again."
JER|22|13|"Woe to him who builds his palace by unrighteousness, his upper rooms by injustice, making his countrymen work for nothing, not paying them for their labor.
JER|22|14|He says, 'I will build myself a great palace with spacious upper rooms.' So he makes large windows in it, panels it with cedar and decorates it in red.
JER|22|15|"Does it make you a king to have more and more cedar? Did not your father have food and drink? He did what was right and just, so all went well with him.
JER|22|16|He defended the cause of the poor and needy, and so all went well. Is that not what it means to know me?" declares the LORD.
JER|22|17|"But your eyes and your heart are set only on dishonest gain, on shedding innocent blood and on oppression and extortion."
JER|22|18|Therefore this is what the LORD says about Jehoiakim son of Josiah king of Judah: "They will not mourn for him: 'Alas, my brother! Alas, my sister!' They will not mourn for him: 'Alas, my master! Alas, his splendor!'
JER|22|19|He will have the burial of a donkey- dragged away and thrown outside the gates of Jerusalem."
JER|22|20|"Go up to Lebanon and cry out, let your voice be heard in Bashan, cry out from Abarim, for all your allies are crushed.
JER|22|21|I warned you when you felt secure, but you said, 'I will not listen!' This has been your way from your youth; you have not obeyed me.
JER|22|22|The wind will drive all your shepherds away, and your allies will go into exile. Then you will be ashamed and disgraced because of all your wickedness.
JER|22|23|You who live in 'Lebanon, 'who are nestled in cedar buildings, how you will groan when pangs come upon you, pain like that of a woman in labor!
JER|22|24|"As surely as I live," declares the LORD, "even if you, Jehoiachin son of Jehoiakim king of Judah, were a signet ring on my right hand, I would still pull you off.
JER|22|25|I will hand you over to those who seek your life, those you fear-to Nebuchadnezzar king of Babylon and to the Babylonians.
JER|22|26|I will hurl you and the mother who gave you birth into another country, where neither of you was born, and there you both will die.
JER|22|27|You will never come back to the land you long to return to."
JER|22|28|Is this man Jehoiachin a despised, broken pot, an object no one wants? Why will he and his children be hurled out, cast into a land they do not know?
JER|22|29|O land, land, land, hear the word of the LORD!
JER|22|30|This is what the LORD says: "Record this man as if childless, a man who will not prosper in his lifetime, for none of his offspring will prosper, none will sit on the throne of David or rule anymore in Judah."
JER|23|1|"Woe to the shepherds who are destroying and scattering the sheep of my pasture!" declares the LORD.
JER|23|2|Therefore this is what the LORD, the God of Israel, says to the shepherds who tend my people: "Because you have scattered my flock and driven them away and have not bestowed care on them, I will bestow punishment on you for the evil you have done," declares the LORD.
JER|23|3|"I myself will gather the remnant of my flock out of all the countries where I have driven them and will bring them back to their pasture, where they will be fruitful and increase in number.
JER|23|4|I will place shepherds over them who will tend them, and they will no longer be afraid or terrified, nor will any be missing," declares the LORD.
JER|23|5|"The days are coming," declares the LORD, "when I will raise up to David a righteous Branch, a King who will reign wisely and do what is just and right in the land.
JER|23|6|In his days Judah will be saved and Israel will live in safety. This is the name by which he will be called: The LORD Our Righteousness.
JER|23|7|"So then, the days are coming," declares the LORD, "when people will no longer say, 'As surely as the LORD lives, who brought the Israelites up out of Egypt,'
JER|23|8|but they will say, 'As surely as the LORD lives, who brought the descendants of Israel up out of the land of the north and out of all the countries where he had banished them.' Then they will live in their own land."
JER|23|9|Concerning the prophets: My heart is broken within me; all my bones tremble. I am like a drunken man, like a man overcome by wine, because of the LORD and his holy words.
JER|23|10|The land is full of adulterers; because of the curse the land lies parched and the pastures in the desert are withered. The prophets follow an evil course and use their power unjustly.
JER|23|11|"Both prophet and priest are godless; even in my temple I find their wickedness," declares the LORD.
JER|23|12|"Therefore their path will become slippery; they will be banished to darkness and there they will fall. I will bring disaster on them in the year they are punished," declares the LORD.
JER|23|13|"Among the prophets of Samaria I saw this repulsive thing: They prophesied by Baal and led my people Israel astray.
JER|23|14|And among the prophets of Jerusalem I have seen something horrible: They commit adultery and live a lie. They strengthen the hands of evildoers, so that no one turns from his wickedness. They are all like Sodom to me; the people of Jerusalem are like Gomorrah."
JER|23|15|Therefore, this is what the LORD Almighty says concerning the prophets: "I will make them eat bitter food and drink poisoned water, because from the prophets of Jerusalem ungodliness has spread throughout the land."
JER|23|16|This is what the LORD Almighty says: "Do not listen to what the prophets are prophesying to you; they fill you with false hopes. They speak visions from their own minds, not from the mouth of the LORD.
JER|23|17|They keep saying to those who despise me, 'The LORD says: You will have peace.' And to all who follow the stubbornness of their hearts they say, 'No harm will come to you.'
JER|23|18|But which of them has stood in the council of the LORD to see or to hear his word? Who has listened and heard his word?
JER|23|19|See, the storm of the LORD will burst out in wrath, a whirlwind swirling down on the heads of the wicked.
JER|23|20|The anger of the LORD will not turn back until he fully accomplishes the purposes of his heart. In days to come you will understand it clearly.
JER|23|21|I did not send these prophets, yet they have run with their message; I did not speak to them, yet they have prophesied.
JER|23|22|But if they had stood in my council, they would have proclaimed my words to my people and would have turned them from their evil ways and from their evil deeds.
JER|23|23|"Am I only a God nearby," declares the LORD, "and not a God far away?
JER|23|24|Can anyone hide in secret places so that I cannot see him?" declares the LORD. "Do not I fill heaven and earth?" declares the LORD.
JER|23|25|"I have heard what the prophets say who prophesy lies in my name. They say, 'I had a dream! I had a dream!'
JER|23|26|How long will this continue in the hearts of these lying prophets, who prophesy the delusions of their own minds?
JER|23|27|They think the dreams they tell one another will make my people forget my name, just as their fathers forgot my name through Baal worship.
JER|23|28|Let the prophet who has a dream tell his dream, but let the one who has my word speak it faithfully. For what has straw to do with grain?" declares the LORD.
JER|23|29|"Is not my word like fire," declares the LORD, "and like a hammer that breaks a rock in pieces?
JER|23|30|"Therefore," declares the LORD, "I am against the prophets who steal from one another words supposedly from me.
JER|23|31|Yes," declares the LORD, "I am against the prophets who wag their own tongues and yet declare, 'The LORD declares.'
JER|23|32|Indeed, I am against those who prophesy false dreams," declares the LORD. "They tell them and lead my people astray with their reckless lies, yet I did not send or appoint them. They do not benefit these people in the least," declares the LORD.
JER|23|33|"When these people, or a prophet or a priest, ask you, 'What is the oracle of the LORD?' say to them, 'What oracle? I will forsake you, declares the LORD.'
JER|23|34|If a prophet or a priest or anyone else claims, 'This is the oracle of the LORD,' I will punish that man and his household.
JER|23|35|This is what each of you keeps on saying to his friend or relative: 'What is the LORD's answer?' or 'What has the LORD spoken?'
JER|23|36|But you must not mention 'the oracle of the LORD 'again, because every man's own word becomes his oracle and so you distort the words of the living God, the LORD Almighty, our God.
JER|23|37|This is what you keep saying to a prophet: 'What is the LORD's answer to you?' or 'What has the LORD spoken?'
JER|23|38|Although you claim, 'This is the oracle of the LORD,' this is what the LORD says: You used the words, 'This is the oracle of the LORD,' even though I told you that you must not claim, 'This is the oracle of the LORD.'
JER|23|39|Therefore, I will surely forget you and cast you out of my presence along with the city I gave to you and your fathers.
JER|23|40|I will bring upon you everlasting disgrace-everlasting shame that will not be forgotten."
JER|24|1|After Jehoiachin son of Jehoiakim king of Judah and the officials, the craftsmen and the artisans of Judah were carried into exile from Jerusalem to Babylon by Nebuchadnezzar king of Babylon, the LORD showed me two baskets of figs placed in front of the temple of the LORD.
JER|24|2|One basket had very good figs, like those that ripen early; the other basket had very poor figs, so bad they could not be eaten.
JER|24|3|Then the LORD asked me, "What do you see, Jeremiah?Figs," I answered. "The good ones are very good, but the poor ones are so bad they cannot be eaten."
JER|24|4|Then the word of the LORD came to me:
JER|24|5|"This is what the LORD, the God of Israel, says: 'Like these good figs, I regard as good the exiles from Judah, whom I sent away from this place to the land of the Babylonians.
JER|24|6|My eyes will watch over them for their good, and I will bring them back to this land. I will build them up and not tear them down; I will plant them and not uproot them.
JER|24|7|I will give them a heart to know me, that I am the LORD. They will be my people, and I will be their God, for they will return to me with all their heart.
JER|24|8|"'But like the poor figs, which are so bad they cannot be eaten,' says the LORD, 'so will I deal with Zedekiah king of Judah, his officials and the survivors from Jerusalem, whether they remain in this land or live in Egypt.
JER|24|9|I will make them abhorrent and an offense to all the kingdoms of the earth, a reproach and a byword, an object of ridicule and cursing, wherever I banish them.
JER|24|10|I will send the sword, famine and plague against them until they are destroyed from the land I gave to them and their fathers.'"
JER|25|1|The word came to Jeremiah concerning all the people of Judah in the fourth year of Jehoiakim son of Josiah king of Judah, which was the first year of Nebuchadnezzar king of Babylon.
JER|25|2|So Jeremiah the prophet said to all the people of Judah and to all those living in Jerusalem:
JER|25|3|For twenty-three years-from the thirteenth year of Josiah son of Amon king of Judah until this very day-the word of the LORD has come to me and I have spoken to you again and again, but you have not listened.
JER|25|4|And though the LORD has sent all his servants the prophets to you again and again, you have not listened or paid any attention.
JER|25|5|They said, "Turn now, each of you, from your evil ways and your evil practices, and you can stay in the land the LORD gave to you and your fathers for ever and ever.
JER|25|6|Do not follow other gods to serve and worship them; do not provoke me to anger with what your hands have made. Then I will not harm you."
JER|25|7|"But you did not listen to me," declares the LORD, "and you have provoked me with what your hands have made, and you have brought harm to yourselves."
JER|25|8|Therefore the LORD Almighty says this: "Because you have not listened to my words,
JER|25|9|I will summon all the peoples of the north and my servant Nebuchadnezzar king of Babylon," declares the LORD, "and I will bring them against this land and its inhabitants and against all the surrounding nations. I will completely destroy them and make them an object of horror and scorn, and an everlasting ruin.
JER|25|10|I will banish from them the sounds of joy and gladness, the voices of bride and bridegroom, the sound of millstones and the light of the lamp.
JER|25|11|This whole country will become a desolate wasteland, and these nations will serve the king of Babylon seventy years.
JER|25|12|"But when the seventy years are fulfilled, I will punish the king of Babylon and his nation, the land of the Babylonians, for their guilt," declares the LORD, "and will make it desolate forever.
JER|25|13|I will bring upon that land all the things I have spoken against it, all that are written in this book and prophesied by Jeremiah against all the nations.
JER|25|14|They themselves will be enslaved by many nations and great kings; I will repay them according to their deeds and the work of their hands."
JER|25|15|This is what the LORD, the God of Israel, said to me: "Take from my hand this cup filled with the wine of my wrath and make all the nations to whom I send you drink it.
JER|25|16|When they drink it, they will stagger and go mad because of the sword I will send among them."
JER|25|17|So I took the cup from the LORD's hand and made all the nations to whom he sent me drink it:
JER|25|18|Jerusalem and the towns of Judah, its kings and officials, to make them a ruin and an object of horror and scorn and cursing, as they are today;
JER|25|19|Pharaoh king of Egypt, his attendants, his officials and all his people,
JER|25|20|and all the foreign people there; all the kings of Uz; all the kings of the Philistines (those of Ashkelon, Gaza, Ekron, and the people left at Ashdod);
JER|25|21|Edom, Moab and Ammon;
JER|25|22|all the kings of Tyre and Sidon; the kings of the coastlands across the sea;
JER|25|23|Dedan, Tema, Buz and all who are in distant places;
JER|25|24|all the kings of Arabia and all the kings of the foreign people who live in the desert;
JER|25|25|all the kings of Zimri, Elam and Media;
JER|25|26|and all the kings of the north, near and far, one after the other-all the kingdoms on the face of the earth. And after all of them, the king of Sheshach will drink it too.
JER|25|27|"Then tell them, 'This is what the LORD Almighty, the God of Israel, says: Drink, get drunk and vomit, and fall to rise no more because of the sword I will send among you.'
JER|25|28|But if they refuse to take the cup from your hand and drink, tell them, 'This is what the LORD Almighty says: You must drink it!
JER|25|29|See, I am beginning to bring disaster on the city that bears my Name, and will you indeed go unpunished? You will not go unpunished, for I am calling down a sword upon all who live on the earth, declares the LORD Almighty.'
JER|25|30|"Now prophesy all these words against them and say to them: "'The LORD will roar from on high; he will thunder from his holy dwelling and roar mightily against his land. He will shout like those who tread the grapes, shout against all who live on the earth.
JER|25|31|The tumult will resound to the ends of the earth, for the LORD will bring charges against the nations; he will bring judgment on all mankind and put the wicked to the sword,'" declares the LORD.
JER|25|32|This is what the LORD Almighty says: "Look! Disaster is spreading from nation to nation; a mighty storm is rising from the ends of the earth."
JER|25|33|At that time those slain by the LORD will be everywhere-from one end of the earth to the other. They will not be mourned or gathered up or buried, but will be like refuse lying on the ground.
JER|25|34|Weep and wail, you shepherds; roll in the dust, you leaders of the flock. For your time to be slaughtered has come; you will fall and be shattered like fine pottery.
JER|25|35|The shepherds will have nowhere to flee, the leaders of the flock no place to escape.
JER|25|36|Hear the cry of the shepherds, the wailing of the leaders of the flock, for the LORD is destroying their pasture.
JER|25|37|The peaceful meadows will be laid waste because of the fierce anger of the LORD.
JER|25|38|Like a lion he will leave his lair, and their land will become desolate because of the sword of the oppressor and because of the LORD's fierce anger.
JER|26|1|Early in the reign of Jehoiakim son of Josiah king of Judah, this word came from the LORD:
JER|26|2|"This is what the LORD says: Stand in the courtyard of the LORD's house and speak to all the people of the towns of Judah who come to worship in the house of the LORD. Tell them everything I command you; do not omit a word.
JER|26|3|Perhaps they will listen and each will turn from his evil way. Then I will relent and not bring on them the disaster I was planning because of the evil they have done.
JER|26|4|Say to them, 'This is what the LORD says: If you do not listen to me and follow my law, which I have set before you,
JER|26|5|and if you do not listen to the words of my servants the prophets, whom I have sent to you again and again (though you have not listened),
JER|26|6|then I will make this house like Shiloh and this city an object of cursing among all the nations of the earth.'"
JER|26|7|The priests, the prophets and all the people heard Jeremiah speak these words in the house of the LORD.
JER|26|8|But as soon as Jeremiah finished telling all the people everything the LORD had commanded him to say, the priests, the prophets and all the people seized him and said, "You must die!
JER|26|9|Why do you prophesy in the LORD's name that this house will be like Shiloh and this city will be desolate and deserted?" And all the people crowded around Jeremiah in the house of the LORD.
JER|26|10|When the officials of Judah heard about these things, they went up from the royal palace to the house of the LORD and took their places at the entrance of the New Gate of the LORD's house.
JER|26|11|Then the priests and the prophets said to the officials and all the people, "This man should be sentenced to death because he has prophesied against this city. You have heard it with your own ears!"
JER|26|12|Then Jeremiah said to all the officials and all the people: "The LORD sent me to prophesy against this house and this city all the things you have heard.
JER|26|13|Now reform your ways and your actions and obey the LORD your God. Then the LORD will relent and not bring the disaster he has pronounced against you.
JER|26|14|As for me, I am in your hands; do with me whatever you think is good and right.
JER|26|15|Be assured, however, that if you put me to death, you will bring the guilt of innocent blood on yourselves and on this city and on those who live in it, for in truth the LORD has sent me to you to speak all these words in your hearing."
JER|26|16|Then the officials and all the people said to the priests and the prophets, "This man should not be sentenced to death! He has spoken to us in the name of the LORD our God."
JER|26|17|Some of the elders of the land stepped forward and said to the entire assembly of people,
JER|26|18|"Micah of Moresheth prophesied in the days of Hezekiah king of Judah. He told all the people of Judah, 'This is what the LORD Almighty says: "'Zion will be plowed like a field, Jerusalem will become a heap of rubble, the temple hill a mound overgrown with thickets.'
JER|26|19|"Did Hezekiah king of Judah or anyone else in Judah put him to death? Did not Hezekiah fear the LORD and seek his favor? And did not the LORD relent, so that he did not bring the disaster he pronounced against them? We are about to bring a terrible disaster on ourselves!"
JER|26|20|(Now Uriah son of Shemaiah from Kiriath Jearim was another man who prophesied in the name of the LORD; he prophesied the same things against this city and this land as Jeremiah did.
JER|26|21|When King Jehoiakim and all his officers and officials heard his words, the king sought to put him to death. But Uriah heard of it and fled in fear to Egypt.
JER|26|22|King Jehoiakim, however, sent Elnathan son of Acbor to Egypt, along with some other men.
JER|26|23|They brought Uriah out of Egypt and took him to King Jehoiakim, who had him struck down with a sword and his body thrown into the burial place of the common people.)
JER|26|24|Furthermore, Ahikam son of Shaphan supported Jeremiah, and so he was not handed over to the people to be put to death.
JER|27|1|Early in the reign of Zedekiah son of Josiah king of Judah, this word came to Jeremiah from the LORD:
JER|27|2|This is what the LORD said to me: "Make a yoke out of straps and crossbars and put it on your neck.
JER|27|3|Then send word to the kings of Edom, Moab, Ammon, Tyre and Sidon through the envoys who have come to Jerusalem to Zedekiah king of Judah.
JER|27|4|Give them a message for their masters and say, 'This is what the LORD Almighty, the God of Israel, says: "Tell this to your masters:
JER|27|5|With my great power and outstretched arm I made the earth and its people and the animals that are on it, and I give it to anyone I please.
JER|27|6|Now I will hand all your countries over to my servant Nebuchadnezzar king of Babylon; I will make even the wild animals subject to him.
JER|27|7|All nations will serve him and his son and his grandson until the time for his land comes; then many nations and great kings will subjugate him.
JER|27|8|"'"If, however, any nation or kingdom will not serve Nebuchadnezzar king of Babylon or bow its neck under his yoke, I will punish that nation with the sword, famine and plague, declares the LORD, until I destroy it by his hand.
JER|27|9|So do not listen to your prophets, your diviners, your interpreters of dreams, your mediums or your sorcerers who tell you, 'You will not serve the king of Babylon.'
JER|27|10|They prophesy lies to you that will only serve to remove you far from your lands; I will banish you and you will perish.
JER|27|11|But if any nation will bow its neck under the yoke of the king of Babylon and serve him, I will let that nation remain in its own land to till it and to live there, declares the LORD."'"
JER|27|12|I gave the same message to Zedekiah king of Judah. I said, "Bow your neck under the yoke of the king of Babylon; serve him and his people, and you will live.
JER|27|13|Why will you and your people die by the sword, famine and plague with which the LORD has threatened any nation that will not serve the king of Babylon?
JER|27|14|Do not listen to the words of the prophets who say to you, 'You will not serve the king of Babylon,' for they are prophesying lies to you.
JER|27|15|'I have not sent them,' declares the LORD. 'They are prophesying lies in my name. Therefore, I will banish you and you will perish, both you and the prophets who prophesy to you.'"
JER|27|16|Then I said to the priests and all these people, "This is what the LORD says: Do not listen to the prophets who say, 'Very soon now the articles from the LORD's house will be brought back from Babylon.' They are prophesying lies to you.
JER|27|17|Do not listen to them. Serve the king of Babylon, and you will live. Why should this city become a ruin?
JER|27|18|If they are prophets and have the word of the LORD, let them plead with the LORD Almighty that the furnishings remaining in the house of the LORD and in the palace of the king of Judah and in Jerusalem not be taken to Babylon.
JER|27|19|For this is what the LORD Almighty says about the pillars, the Sea, the movable stands and the other furnishings that are left in this city,
JER|27|20|which Nebuchadnezzar king of Babylon did not take away when he carried Jehoiachin son of Jehoiakim king of Judah into exile from Jerusalem to Babylon, along with all the nobles of Judah and Jerusalem-
JER|27|21|yes, this is what the LORD Almighty, the God of Israel, says about the things that are left in the house of the LORD and in the palace of the king of Judah and in Jerusalem:
JER|27|22|'They will be taken to Babylon and there they will remain until the day I come for them,' declares the LORD. 'Then I will bring them back and restore them to this place.'"
JER|28|1|In the fifth month of that same year, the fourth year, early in the reign of Zedekiah king of Judah, the prophet Hananiah son of Azzur, who was from Gibeon, said to me in the house of the LORD in the presence of the priests and all the people:
JER|28|2|"This is what the LORD Almighty, the God of Israel, says: 'I will break the yoke of the king of Babylon.
JER|28|3|Within two years I will bring back to this place all the articles of the LORD's house that Nebuchadnezzar king of Babylon removed from here and took to Babylon.
JER|28|4|I will also bring back to this place Jehoiachin son of Jehoiakim king of Judah and all the other exiles from Judah who went to Babylon,' declares the LORD, 'for I will break the yoke of the king of Babylon.'"
JER|28|5|Then the prophet Jeremiah replied to the prophet Hananiah before the priests and all the people who were standing in the house of the LORD.
JER|28|6|He said, "Amen! May the LORD do so! May the LORD fulfill the words you have prophesied by bringing the articles of the LORD's house and all the exiles back to this place from Babylon.
JER|28|7|Nevertheless, listen to what I have to say in your hearing and in the hearing of all the people:
JER|28|8|From early times the prophets who preceded you and me have prophesied war, disaster and plague against many countries and great kingdoms.
JER|28|9|But the prophet who prophesies peace will be recognized as one truly sent by the LORD only if his prediction comes true."
JER|28|10|Then the prophet Hananiah took the yoke off the neck of the prophet Jeremiah and broke it,
JER|28|11|and he said before all the people, "This is what the LORD says: 'In the same way will I break the yoke of Nebuchadnezzar king of Babylon off the neck of all the nations within two years.'" At this, the prophet Jeremiah went on his way.
JER|28|12|Shortly after the prophet Hananiah had broken the yoke off the neck of the prophet Jeremiah, the word of the LORD came to Jeremiah:
JER|28|13|"Go and tell Hananiah, 'This is what the LORD says: You have broken a wooden yoke, but in its place you will get a yoke of iron.
JER|28|14|This is what the LORD Almighty, the God of Israel, says: I will put an iron yoke on the necks of all these nations to make them serve Nebuchadnezzar king of Babylon, and they will serve him. I will even give him control over the wild animals.'"
JER|28|15|Then the prophet Jeremiah said to Hananiah the prophet, "Listen, Hananiah! The LORD has not sent you, yet you have persuaded this nation to trust in lies.
JER|28|16|Therefore, this is what the LORD says: 'I am about to remove you from the face of the earth. This very year you are going to die, because you have preached rebellion against the LORD.'"
JER|28|17|In the seventh month of that same year, Hananiah the prophet died.
JER|29|1|This is the text of the letter that the prophet Jeremiah sent from Jerusalem to the surviving elders among the exiles and to the priests, the prophets and all the other people Nebuchadnezzar had carried into exile from Jerusalem to Babylon.
JER|29|2|(This was after King Jehoiachin and the queen mother, the court officials and the leaders of Judah and Jerusalem, the craftsmen and the artisans had gone into exile from Jerusalem.)
JER|29|3|He entrusted the letter to Elasah son of Shaphan and to Gemariah son of Hilkiah, whom Zedekiah king of Judah sent to King Nebuchadnezzar in Babylon. It said:
JER|29|4|This is what the LORD Almighty, the God of Israel, says to all those I carried into exile from Jerusalem to Babylon:
JER|29|5|"Build houses and settle down; plant gardens and eat what they produce.
JER|29|6|Marry and have sons and daughters; find wives for your sons and give your daughters in marriage, so that they too may have sons and daughters. Increase in number there; do not decrease.
JER|29|7|Also, seek the peace and prosperity of the city to which I have carried you into exile. Pray to the LORD for it, because if it prospers, you too will prosper."
JER|29|8|Yes, this is what the LORD Almighty, the God of Israel, says: "Do not let the prophets and diviners among you deceive you. Do not listen to the dreams you encourage them to have.
JER|29|9|They are prophesying lies to you in my name. I have not sent them," declares the LORD.
JER|29|10|This is what the LORD says: "When seventy years are completed for Babylon, I will come to you and fulfill my gracious promise to bring you back to this place.
JER|29|11|For I know the plans I have for you," declares the LORD, "plans to prosper you and not to harm you, plans to give you hope and a future.
JER|29|12|Then you will call upon me and come and pray to me, and I will listen to you.
JER|29|13|You will seek me and find me when you seek me with all your heart.
JER|29|14|I will be found by you," declares the LORD, "and will bring you back from captivity. I will gather you from all the nations and places where I have banished you," declares the LORD, "and will bring you back to the place from which I carried you into exile."
JER|29|15|You may say, "The LORD has raised up prophets for us in Babylon,"
JER|29|16|but this is what the LORD says about the king who sits on David's throne and all the people who remain in this city, your countrymen who did not go with you into exile-
JER|29|17|yes, this is what the LORD Almighty says: "I will send the sword, famine and plague against them and I will make them like poor figs that are so bad they cannot be eaten.
JER|29|18|I will pursue them with the sword, famine and plague and will make them abhorrent to all the kingdoms of the earth and an object of cursing and horror, of scorn and reproach, among all the nations where I drive them.
JER|29|19|For they have not listened to my words," declares the LORD, "words that I sent to them again and again by my servants the prophets. And you exiles have not listened either," declares the LORD.
JER|29|20|Therefore, hear the word of the LORD, all you exiles whom I have sent away from Jerusalem to Babylon.
JER|29|21|This is what the LORD Almighty, the God of Israel, says about Ahab son of Kolaiah and Zedekiah son of Maaseiah, who are prophesying lies to you in my name: "I will hand them over to Nebuchadnezzar king of Babylon, and he will put them to death before your very eyes.
JER|29|22|Because of them, all the exiles from Judah who are in Babylon will use this curse: 'The LORD treat you like Zedekiah and Ahab, whom the king of Babylon burned in the fire.'
JER|29|23|For they have done outrageous things in Israel; they have committed adultery with their neighbors' wives and in my name have spoken lies, which I did not tell them to do. I know it and am a witness to it," declares the LORD.
JER|29|24|Tell Shemaiah the Nehelamite,
JER|29|25|"This is what the LORD Almighty, the God of Israel, says: You sent letters in your own name to all the people in Jerusalem, to Zephaniah son of Maaseiah the priest, and to all the other priests. You said to Zephaniah,
JER|29|26|'The LORD has appointed you priest in place of Jehoiada to be in charge of the house of the LORD; you should put any madman who acts like a prophet into the stocks and neck-irons.
JER|29|27|So why have you not reprimanded Jeremiah from Anathoth, who poses as a prophet among you?
JER|29|28|He has sent this message to us in Babylon: It will be a long time. Therefore build houses and settle down; plant gardens and eat what they produce.'"
JER|29|29|Zephaniah the priest, however, read the letter to Jeremiah the prophet.
JER|29|30|Then the word of the LORD came to Jeremiah:
JER|29|31|"Send this message to all the exiles: 'This is what the LORD says about Shemaiah the Nehelamite: Because Shemaiah has prophesied to you, even though I did not send him, and has led you to believe a lie,
JER|29|32|this is what the LORD says: I will surely punish Shemaiah the Nehelamite and his descendants. He will have no one left among this people, nor will he see the good things I will do for my people, declares the LORD, because he has preached rebellion against me.'"
JER|30|1|This is the word that came to Jeremiah from the LORD:
JER|30|2|"This is what the LORD, the God of Israel, says: 'Write in a book all the words I have spoken to you.
JER|30|3|The days are coming,' declares the LORD, 'when I will bring my people Israel and Judah back from captivity and restore them to the land I gave their forefathers to possess,' says the LORD."
JER|30|4|These are the words the LORD spoke concerning Israel and Judah:
JER|30|5|"This is what the LORD says: "'Cries of fear are heard- terror, not peace.
JER|30|6|Ask and see: Can a man bear children? Then why do I see every strong man with his hands on his stomach like a woman in labor, every face turned deathly pale?
JER|30|7|How awful that day will be! None will be like it. It will be a time of trouble for Jacob, but he will be saved out of it.
JER|30|8|"'In that day,' declares the LORD Almighty, 'I will break the yoke off their necks and will tear off their bonds; no longer will foreigners enslave them.
JER|30|9|Instead, they will serve the LORD their God and David their king, whom I will raise up for them.
JER|30|10|"'So do not fear, O Jacob my servant; do not be dismayed, O Israel,' declares the LORD. 'I will surely save you out of a distant place, your descendants from the land of their exile. Jacob will again have peace and security, and no one will make him afraid.
JER|30|11|I am with you and will save you,' declares the LORD. 'Though I completely destroy all the nations among which I scatter you, I will not completely destroy you. I will discipline you but only with justice; I will not let you go entirely unpunished.'
JER|30|12|"This is what the LORD says: "'Your wound is incurable, your injury beyond healing.
JER|30|13|There is no one to plead your cause, no remedy for your sore, no healing for you.
JER|30|14|All your allies have forgotten you; they care nothing for you. I have struck you as an enemy would and punished you as would the cruel, because your guilt is so great and your sins so many.
JER|30|15|Why do you cry out over your wound, your pain that has no cure? Because of your great guilt and many sins I have done these things to you.
JER|30|16|"'But all who devour you will be devoured; all your enemies will go into exile. Those who plunder you will be plundered; all who make spoil of you I will despoil.
JER|30|17|But I will restore you to health and heal your wounds,' declares the LORD, 'because you are called an outcast, Zion for whom no one cares.'
JER|30|18|"This is what the LORD says: "'I will restore the fortunes of Jacob's tents and have compassion on his dwellings; the city will be rebuilt on her ruins, and the palace will stand in its proper place.
JER|30|19|From them will come songs of thanksgiving and the sound of rejoicing. I will add to their numbers, and they will not be decreased; I will bring them honor, and they will not be disdained.
JER|30|20|Their children will be as in days of old, and their community will be established before me; I will punish all who oppress them.
JER|30|21|Their leader will be one of their own; their ruler will arise from among them. I will bring him near and he will come close to me, for who is he who will devote himself to be close to me?' declares the LORD.
JER|30|22|"'So you will be my people, and I will be your God.'"
JER|30|23|See, the storm of the LORD will burst out in wrath, a driving wind swirling down on the heads of the wicked.
JER|30|24|The fierce anger of the LORD will not turn back until he fully accomplishes the purposes of his heart. In days to come you will understand this.
JER|31|1|"At that time," declares the LORD, "I will be the God of all the clans of Israel, and they will be my people."
JER|31|2|This is what the LORD says: "The people who survive the sword will find favor in the desert; I will come to give rest to Israel."
JER|31|3|The LORD appeared to us in the past, saying: "I have loved you with an everlasting love; I have drawn you with loving-kindness.
JER|31|4|I will build you up again and you will be rebuilt, O Virgin Israel. Again you will take up your tambourines and go out to dance with the joyful.
JER|31|5|Again you will plant vineyards on the hills of Samaria; the farmers will plant them and enjoy their fruit.
JER|31|6|There will be a day when watchmen cry out on the hills of Ephraim, 'Come, let us go up to Zion, to the LORD our God.'"
JER|31|7|This is what the LORD says: "Sing with joy for Jacob; shout for the foremost of the nations. Make your praises heard, and say, 'O LORD, save your people, the remnant of Israel.'
JER|31|8|See, I will bring them from the land of the north and gather them from the ends of the earth. Among them will be the blind and the lame, expectant mothers and women in labor; a great throng will return.
JER|31|9|They will come with weeping; they will pray as I bring them back. I will lead them beside streams of water on a level path where they will not stumble, because I am Israel's father, and Ephraim is my firstborn son.
JER|31|10|"Hear the word of the LORD, O nations; proclaim it in distant coastlands: 'He who scattered Israel will gather them and will watch over his flock like a shepherd.'
JER|31|11|For the LORD will ransom Jacob and redeem them from the hand of those stronger than they.
JER|31|12|They will come and shout for joy on the heights of Zion; they will rejoice in the bounty of the LORD - the grain, the new wine and the oil, the young of the flocks and herds. They will be like a well-watered garden, and they will sorrow no more.
JER|31|13|Then maidens will dance and be glad, young men and old as well. I will turn their mourning into gladness; I will give them comfort and joy instead of sorrow.
JER|31|14|I will satisfy the priests with abundance, and my people will be filled with my bounty," declares the LORD.
JER|31|15|This is what the LORD says: "A voice is heard in Ramah, mourning and great weeping, Rachel weeping for her children and refusing to be comforted, because her children are no more."
JER|31|16|This is what the LORD says: "Restrain your voice from weeping and your eyes from tears, for your work will be rewarded," declares the LORD. "They will return from the land of the enemy.
JER|31|17|So there is hope for your future," declares the LORD. "Your children will return to their own land.
JER|31|18|"I have surely heard Ephraim's moaning: 'You disciplined me like an unruly calf, and I have been disciplined. Restore me, and I will return, because you are the LORD my God.
JER|31|19|After I strayed, I repented; after I came to understand, I beat my breast. I was ashamed and humiliated because I bore the disgrace of my youth.'
JER|31|20|Is not Ephraim my dear son, the child in whom I delight? Though I often speak against him, I still remember him. Therefore my heart yearns for him; I have great compassion for him," declares the LORD.
JER|31|21|"Set up road signs; put up guideposts. Take note of the highway, the road that you take. Return, O Virgin Israel, return to your towns.
JER|31|22|How long will you wander, O unfaithful daughter? The LORD will create a new thing on earth- a woman will surround a man."
JER|31|23|This is what the LORD Almighty, the God of Israel, says: "When I bring them back from captivity, the people in the land of Judah and in its towns will once again use these words: 'The LORD bless you, O righteous dwelling, O sacred mountain.'
JER|31|24|People will live together in Judah and all its towns-farmers and those who move about with their flocks.
JER|31|25|I will refresh the weary and satisfy the faint."
JER|31|26|At this I awoke and looked around. My sleep had been pleasant to me.
JER|31|27|"The days are coming," declares the LORD, "when I will plant the house of Israel and the house of Judah with the offspring of men and of animals.
JER|31|28|Just as I watched over them to uproot and tear down, and to overthrow, destroy and bring disaster, so I will watch over them to build and to plant," declares the LORD.
JER|31|29|"In those days people will no longer say, 'The fathers have eaten sour grapes, and the children's teeth are set on edge.'
JER|31|30|Instead, everyone will die for his own sin; whoever eats sour grapes-his own teeth will be set on edge.
JER|31|31|"The time is coming," declares the LORD, "when I will make a new covenant with the house of Israel and with the house of Judah.
JER|31|32|It will not be like the covenant I made with their forefathers when I took them by the hand to lead them out of Egypt, because they broke my covenant, though I was a husband to them, "declares the LORD.
JER|31|33|"This is the covenant I will make with the house of Israel after that time," declares the LORD. "I will put my law in their minds and write it on their hearts. I will be their God, and they will be my people.
JER|31|34|No longer will a man teach his neighbor, or a man his brother, saying, 'Know the LORD,' because they will all know me, from the least of them to the greatest," declares the LORD. "For I will forgive their wickedness and will remember their sins no more."
JER|31|35|This is what the LORD says, he who appoints the sun to shine by day, who decrees the moon and stars to shine by night, who stirs up the sea so that its waves roar- the LORD Almighty is his name:
JER|31|36|"Only if these decrees vanish from my sight," declares the LORD, "will the descendants of Israel ever cease to be a nation before me."
JER|31|37|This is what the LORD says: "Only if the heavens above can be measured and the foundations of the earth below be searched out will I reject all the descendants of Israel because of all they have done," declares the LORD.
JER|31|38|"The days are coming," declares the LORD, "when this city will be rebuilt for me from the Tower of Hananel to the Corner Gate.
JER|31|39|The measuring line will stretch from there straight to the hill of Gareb and then turn to Goah.
JER|31|40|The whole valley where dead bodies and ashes are thrown, and all the terraces out to the Kidron Valley on the east as far as the corner of the Horse Gate, will be holy to the LORD. The city will never again be uprooted or demolished."
JER|32|1|This is the word that came to Jeremiah from the LORD in the tenth year of Zedekiah king of Judah, which was the eighteenth year of Nebuchadnezzar.
JER|32|2|The army of the king of Babylon was then besieging Jerusalem, and Jeremiah the prophet was confined in the courtyard of the guard in the royal palace of Judah.
JER|32|3|Now Zedekiah king of Judah had imprisoned him there, saying, "Why do you prophesy as you do? You say, 'This is what the LORD says: I am about to hand this city over to the king of Babylon, and he will capture it.
JER|32|4|Zedekiah king of Judah will not escape out of the hands of the Babylonians but will certainly be handed over to the king of Babylon, and will speak with him face to face and see him with his own eyes.
JER|32|5|He will take Zedekiah to Babylon, where he will remain until I deal with him, declares the LORD. If you fight against the Babylonians, you will not succeed.'"
JER|32|6|Jeremiah said, "The word of the LORD came to me:
JER|32|7|Hanamel son of Shallum your uncle is going to come to you and say, 'Buy my field at Anathoth, because as nearest relative it is your right and duty to buy it.'
JER|32|8|"Then, just as the LORD had said, my cousin Hanamel came to me in the courtyard of the guard and said, 'Buy my field at Anathoth in the territory of Benjamin. Since it is your right to redeem it and possess it, buy it for yourself.'"I knew that this was the word of the LORD;
JER|32|9|so I bought the field at Anathoth from my cousin Hanamel and weighed out for him seventeen shekels of silver.
JER|32|10|I signed and sealed the deed, had it witnessed, and weighed out the silver on the scales.
JER|32|11|I took the deed of purchase-the sealed copy containing the terms and conditions, as well as the unsealed copy-
JER|32|12|and I gave this deed to Baruch son of Neriah, the son of Mahseiah, in the presence of my cousin Hanamel and of the witnesses who had signed the deed and of all the Jews sitting in the courtyard of the guard.
JER|32|13|"In their presence I gave Baruch these instructions:
JER|32|14|'This is what the LORD Almighty, the God of Israel, says: Take these documents, both the sealed and unsealed copies of the deed of purchase, and put them in a clay jar so they will last a long time.
JER|32|15|For this is what the LORD Almighty, the God of Israel, says: Houses, fields and vineyards will again be bought in this land.'
JER|32|16|"After I had given the deed of purchase to Baruch son of Neriah, I prayed to the LORD:
JER|32|17|"Ah, Sovereign LORD, you have made the heavens and the earth by your great power and outstretched arm. Nothing is too hard for you.
JER|32|18|You show love to thousands but bring the punishment for the fathers' sins into the laps of their children after them. O great and powerful God, whose name is the LORD Almighty,
JER|32|19|great are your purposes and mighty are your deeds. Your eyes are open to all the ways of men; you reward everyone according to his conduct and as his deeds deserve.
JER|32|20|You performed miraculous signs and wonders in Egypt and have continued them to this day, both in Israel and among all mankind, and have gained the renown that is still yours.
JER|32|21|You brought your people Israel out of Egypt with signs and wonders, by a mighty hand and an outstretched arm and with great terror.
JER|32|22|You gave them this land you had sworn to give their forefathers, a land flowing with milk and honey.
JER|32|23|They came in and took possession of it, but they did not obey you or follow your law; they did not do what you commanded them to do. So you brought all this disaster upon them.
JER|32|24|"See how the siege ramps are built up to take the city. Because of the sword, famine and plague, the city will be handed over to the Babylonians who are attacking it. What you said has happened, as you now see.
JER|32|25|And though the city will be handed over to the Babylonians, you, O Sovereign LORD, say to me, 'Buy the field with silver and have the transaction witnessed.'"
JER|32|26|Then the word of the LORD came to Jeremiah:
JER|32|27|"I am the LORD, the God of all mankind. Is anything too hard for me?
JER|32|28|Therefore, this is what the LORD says: I am about to hand this city over to the Babylonians and to Nebuchadnezzar king of Babylon, who will capture it.
JER|32|29|The Babylonians who are attacking this city will come in and set it on fire; they will burn it down, along with the houses where the people provoked me to anger by burning incense on the roofs to Baal and by pouring out drink offerings to other gods.
JER|32|30|"The people of Israel and Judah have done nothing but evil in my sight from their youth; indeed, the people of Israel have done nothing but provoke me with what their hands have made, declares the LORD.
JER|32|31|From the day it was built until now, this city has so aroused my anger and wrath that I must remove it from my sight.
JER|32|32|The people of Israel and Judah have provoked me by all the evil they have done-they, their kings and officials, their priests and prophets, the men of Judah and the people of Jerusalem.
JER|32|33|They turned their backs to me and not their faces; though I taught them again and again, they would not listen or respond to discipline.
JER|32|34|They set up their abominable idols in the house that bears my Name and defiled it.
JER|32|35|They built high places for Baal in the Valley of Ben Hinnom to sacrifice their sons and daughters to Molech, though I never commanded, nor did it enter my mind, that they should do such a detestable thing and so make Judah sin.
JER|32|36|"You are saying about this city, 'By the sword, famine and plague it will be handed over to the king of Babylon'; but this is what the LORD, the God of Israel, says:
JER|32|37|I will surely gather them from all the lands where I banish them in my furious anger and great wrath; I will bring them back to this place and let them live in safety.
JER|32|38|They will be my people, and I will be their God.
JER|32|39|I will give them singleness of heart and action, so that they will always fear me for their own good and the good of their children after them.
JER|32|40|I will make an everlasting covenant with them: I will never stop doing good to them, and I will inspire them to fear me, so that they will never turn away from me.
JER|32|41|I will rejoice in doing them good and will assuredly plant them in this land with all my heart and soul.
JER|32|42|"This is what the LORD says: As I have brought all this great calamity on this people, so I will give them all the prosperity I have promised them.
JER|32|43|Once more fields will be bought in this land of which you say, 'It is a desolate waste, without men or animals, for it has been handed over to the Babylonians.'
JER|32|44|Fields will be bought for silver, and deeds will be signed, sealed and witnessed in the territory of Benjamin, in the villages around Jerusalem, in the towns of Judah and in the towns of the hill country, of the western foothills and of the Negev, because I will restore their fortunes, declares the LORD."
JER|33|1|While Jeremiah was still confined in the courtyard of the guard, the word of the LORD came to him a second time:
JER|33|2|"This is what the LORD says, he who made the earth, the LORD who formed it and established it-the LORD is his name:
JER|33|3|'Call to me and I will answer you and tell you great and unsearchable things you do not know.'
JER|33|4|For this is what the LORD, the God of Israel, says about the houses in this city and the royal palaces of Judah that have been torn down to be used against the siege ramps and the sword
JER|33|5|in the fight with the Babylonians: 'They will be filled with the dead bodies of the men I will slay in my anger and wrath. I will hide my face from this city because of all its wickedness.
JER|33|6|"'Nevertheless, I will bring health and healing to it; I will heal my people and will let them enjoy abundant peace and security.
JER|33|7|I will bring Judah and Israel back from captivity and will rebuild them as they were before.
JER|33|8|I will cleanse them from all the sin they have committed against me and will forgive all their sins of rebellion against me.
JER|33|9|Then this city will bring me renown, joy, praise and honor before all nations on earth that hear of all the good things I do for it; and they will be in awe and will tremble at the abundant prosperity and peace I provide for it.'
JER|33|10|"This is what the LORD says: 'You say about this place, "It is a desolate waste, without men or animals." Yet in the towns of Judah and the streets of Jerusalem that are deserted, inhabited by neither men nor animals, there will be heard once more
JER|33|11|the sounds of joy and gladness, the voices of bride and bridegroom, and the voices of those who bring thank offerings to the house of the LORD, saying, "Give thanks to the LORD Almighty, for the LORD is good; his love endures forever." For I will restore the fortunes of the land as they were before,' says the LORD.
JER|33|12|"This is what the LORD Almighty says: 'In this place, desolate and without men or animals-in all its towns there will again be pastures for shepherds to rest their flocks.
JER|33|13|In the towns of the hill country, of the western foothills and of the Negev, in the territory of Benjamin, in the villages around Jerusalem and in the towns of Judah, flocks will again pass under the hand of the one who counts them,' says the LORD.
JER|33|14|"'The days are coming,' declares the LORD, 'when I will fulfill the gracious promise I made to the house of Israel and to the house of Judah.
JER|33|15|"'In those days and at that time I will make a righteous Branch sprout from David's line; he will do what is just and right in the land.
JER|33|16|In those days Judah will be saved and Jerusalem will live in safety. This is the name by which it will be called: The LORD Our Righteousness.'
JER|33|17|For this is what the LORD says: 'David will never fail to have a man to sit on the throne of the house of Israel,
JER|33|18|nor will the priests, who are Levites, ever fail to have a man to stand before me continually to offer burnt offerings, to burn grain offerings and to present sacrifices.'"
JER|33|19|The word of the LORD came to Jeremiah:
JER|33|20|"This is what the LORD says: 'If you can break my covenant with the day and my covenant with the night, so that day and night no longer come at their appointed time,
JER|33|21|then my covenant with David my servant-and my covenant with the Levites who are priests ministering before me-can be broken and David will no longer have a descendant to reign on his throne.
JER|33|22|I will make the descendants of David my servant and the Levites who minister before me as countless as the stars of the sky and as measureless as the sand on the seashore.'"
JER|33|23|The word of the LORD came to Jeremiah:
JER|33|24|"Have you not noticed that these people are saying, 'The LORD has rejected the two kingdoms he chose'? So they despise my people and no longer regard them as a nation.
JER|33|25|This is what the LORD says: 'If I have not established my covenant with day and night and the fixed laws of heaven and earth,
JER|33|26|then I will reject the descendants of Jacob and David my servant and will not choose one of his sons to rule over the descendants of Abraham, Isaac and Jacob. For I will restore their fortunes and have compassion on them.'"
JER|34|1|While Nebuchadnezzar king of Babylon and all his army and all the kingdoms and peoples in the empire he ruled were fighting against Jerusalem and all its surrounding towns, this word came to Jeremiah from the LORD:
JER|34|2|"This is what the LORD, the God of Israel, says: Go to Zedekiah king of Judah and tell him, 'This is what the LORD says: I am about to hand this city over to the king of Babylon, and he will burn it down.
JER|34|3|You will not escape from his grasp but will surely be captured and handed over to him. You will see the king of Babylon with your own eyes, and he will speak with you face to face. And you will go to Babylon.
JER|34|4|"'Yet hear the promise of the LORD, O Zedekiah king of Judah. This is what the LORD says concerning you: You will not die by the sword;
JER|34|5|you will die peacefully. As people made a funeral fire in honor of your fathers, the former kings who preceded you, so they will make a fire in your honor and lament, "Alas, O master!" I myself make this promise, declares the LORD.'"
JER|34|6|Then Jeremiah the prophet told all this to Zedekiah king of Judah, in Jerusalem,
JER|34|7|while the army of the king of Babylon was fighting against Jerusalem and the other cities of Judah that were still holding out-Lachish and Azekah. These were the only fortified cities left in Judah.
JER|34|8|The word came to Jeremiah from the LORD after King Zedekiah had made a covenant with all the people in Jerusalem to proclaim freedom for the slaves.
JER|34|9|Everyone was to free his Hebrew slaves, both male and female; no one was to hold a fellow Jew in bondage.
JER|34|10|So all the officials and people who entered into this covenant agreed that they would free their male and female slaves and no longer hold them in bondage. They agreed, and set them free.
JER|34|11|But afterward they changed their minds and took back the slaves they had freed and enslaved them again.
JER|34|12|Then the word of the LORD came to Jeremiah:
JER|34|13|"This is what the LORD, the God of Israel, says: I made a covenant with your forefathers when I brought them out of Egypt, out of the land of slavery. I said,
JER|34|14|'Every seventh year each of you must free any fellow Hebrew who has sold himself to you. After he has served you six years, you must let him go free.' Your fathers, however, did not listen to me or pay attention to me.
JER|34|15|Recently you repented and did what is right in my sight: Each of you proclaimed freedom to his countrymen. You even made a covenant before me in the house that bears my Name.
JER|34|16|But now you have turned around and profaned my name; each of you has taken back the male and female slaves you had set free to go where they wished. You have forced them to become your slaves again.
JER|34|17|"Therefore, this is what the LORD says: You have not obeyed me; you have not proclaimed freedom for your fellow countrymen. So I now proclaim 'freedom' for you, declares the LORD -'freedom' to fall by the sword, plague and famine. I will make you abhorrent to all the kingdoms of the earth.
JER|34|18|The men who have violated my covenant and have not fulfilled the terms of the covenant they made before me, I will treat like the calf they cut in two and then walked between its pieces.
JER|34|19|The leaders of Judah and Jerusalem, the court officials, the priests and all the people of the land who walked between the pieces of the calf,
JER|34|20|I will hand over to their enemies who seek their lives. Their dead bodies will become food for the birds of the air and the beasts of the earth.
JER|34|21|"I will hand Zedekiah king of Judah and his officials over to their enemies who seek their lives, to the army of the king of Babylon, which has withdrawn from you.
JER|34|22|I am going to give the order, declares the LORD, and I will bring them back to this city. They will fight against it, take it and burn it down. And I will lay waste the towns of Judah so no one can live there."
JER|35|1|This is the word that came to Jeremiah from the LORD during the reign of Jehoiakim son of Josiah king of Judah:
JER|35|2|"Go to the Recabite family and invite them to come to one of the side rooms of the house of the LORD and give them wine to drink."
JER|35|3|So I went to get Jaazaniah son of Jeremiah, the son of Habazziniah, and his brothers and all his sons-the whole family of the Recabites.
JER|35|4|I brought them into the house of the LORD, into the room of the sons of Hanan son of Igdaliah the man of God. It was next to the room of the officials, which was over that of Maaseiah son of Shallum the doorkeeper.
JER|35|5|Then I set bowls full of wine and some cups before the men of the Recabite family and said to them, "Drink some wine."
JER|35|6|But they replied, "We do not drink wine, because our forefather Jonadab son of Recab gave us this command: 'Neither you nor your descendants must ever drink wine.
JER|35|7|Also you must never build houses, sow seed or plant vineyards; you must never have any of these things, but must always live in tents. Then you will live a long time in the land where you are nomads.'
JER|35|8|We have obeyed everything our forefather Jonadab son of Recab commanded us. Neither we nor our wives nor our sons and daughters have ever drunk wine
JER|35|9|or built houses to live in or had vineyards, fields or crops.
JER|35|10|We have lived in tents and have fully obeyed everything our forefather Jonadab commanded us.
JER|35|11|But when Nebuchadnezzar king of Babylon invaded this land, we said, 'Come, we must go to Jerusalem to escape the Babylonian and Aramean armies.' So we have remained in Jerusalem."
JER|35|12|Then the word of the LORD came to Jeremiah, saying:
JER|35|13|"This is what the LORD Almighty, the God of Israel, says: Go and tell the men of Judah and the people of Jerusalem, 'Will you not learn a lesson and obey my words?' declares the LORD.
JER|35|14|'Jonadab son of Recab ordered his sons not to drink wine and this command has been kept. To this day they do not drink wine, because they obey their forefather's command. But I have spoken to you again and again, yet you have not obeyed me.
JER|35|15|Again and again I sent all my servants the prophets to you. They said, "Each of you must turn from your wicked ways and reform your actions; do not follow other gods to serve them. Then you will live in the land I have given to you and your fathers." But you have not paid attention or listened to me.
JER|35|16|The descendants of Jonadab son of Recab have carried out the command their forefather gave them, but these people have not obeyed me.'
JER|35|17|"Therefore, this is what the LORD God Almighty, the God of Israel, says: 'Listen! I am going to bring on Judah and on everyone living in Jerusalem every disaster I pronounced against them. I spoke to them, but they did not listen; I called to them, but they did not answer.'"
JER|35|18|Then Jeremiah said to the family of the Recabites, "This is what the LORD Almighty, the God of Israel, says: 'You have obeyed the command of your forefather Jonadab and have followed all his instructions and have done everything he ordered.'
JER|35|19|Therefore, this is what the LORD Almighty, the God of Israel, says: 'Jonadab son of Recab will never fail to have a man to serve me.'"
JER|36|1|In the fourth year of Jehoiakim son of Josiah king of Judah, this word came to Jeremiah from the LORD:
JER|36|2|"Take a scroll and write on it all the words I have spoken to you concerning Israel, Judah and all the other nations from the time I began speaking to you in the reign of Josiah till now.
JER|36|3|Perhaps when the people of Judah hear about every disaster I plan to inflict on them, each of them will turn from his wicked way; then I will forgive their wickedness and their sin."
JER|36|4|So Jeremiah called Baruch son of Neriah, and while Jeremiah dictated all the words the LORD had spoken to him, Baruch wrote them on the scroll.
JER|36|5|Then Jeremiah told Baruch, "I am restricted; I cannot go to the LORD's temple.
JER|36|6|So you go to the house of the LORD on a day of fasting and read to the people from the scroll the words of the LORD that you wrote as I dictated. Read them to all the people of Judah who come in from their towns.
JER|36|7|Perhaps they will bring their petition before the LORD, and each will turn from his wicked ways, for the anger and wrath pronounced against this people by the LORD are great."
JER|36|8|Baruch son of Neriah did everything Jeremiah the prophet told him to do; at the LORD's temple he read the words of the LORD from the scroll.
JER|36|9|In the ninth month of the fifth year of Jehoiakim son of Josiah king of Judah, a time of fasting before the LORD was proclaimed for all the people in Jerusalem and those who had come from the towns of Judah.
JER|36|10|From the room of Gemariah son of Shaphan the secretary, which was in the upper courtyard at the entrance of the New Gate of the temple, Baruch read to all the people at the LORD's temple the words of Jeremiah from the scroll.
JER|36|11|When Micaiah son of Gemariah, the son of Shaphan, heard all the words of the LORD from the scroll,
JER|36|12|he went down to the secretary's room in the royal palace, where all the officials were sitting: Elishama the secretary, Delaiah son of Shemaiah, Elnathan son of Acbor, Gemariah son of Shaphan, Zedekiah son of Hananiah, and all the other officials.
JER|36|13|After Micaiah told them everything he had heard Baruch read to the people from the scroll,
JER|36|14|all the officials sent Jehudi son of Nethaniah, the son of Shelemiah, the son of Cushi, to say to Baruch, "Bring the scroll from which you have read to the people and come." So Baruch son of Neriah went to them with the scroll in his hand.
JER|36|15|They said to him, "Sit down, please, and read it to us." So Baruch read it to them.
JER|36|16|When they heard all these words, they looked at each other in fear and said to Baruch, "We must report all these words to the king."
JER|36|17|Then they asked Baruch, "Tell us, how did you come to write all this? Did Jeremiah dictate it?"
JER|36|18|"Yes," Baruch replied, "he dictated all these words to me, and I wrote them in ink on the scroll."
JER|36|19|Then the officials said to Baruch, "You and Jeremiah, go and hide. Don't let anyone know where you are."
JER|36|20|After they put the scroll in the room of Elishama the secretary, they went to the king in the courtyard and reported everything to him.
JER|36|21|The king sent Jehudi to get the scroll, and Jehudi brought it from the room of Elishama the secretary and read it to the king and all the officials standing beside him.
JER|36|22|It was the ninth month and the king was sitting in the winter apartment, with a fire burning in the firepot in front of him.
JER|36|23|Whenever Jehudi had read three or four columns of the scroll, the king cut them off with a scribe's knife and threw them into the firepot, until the entire scroll was burned in the fire.
JER|36|24|The king and all his attendants who heard all these words showed no fear, nor did they tear their clothes.
JER|36|25|Even though Elnathan, Delaiah and Gemariah urged the king not to burn the scroll, he would not listen to them.
JER|36|26|Instead, the king commanded Jerahmeel, a son of the king, Seraiah son of Azriel and Shelemiah son of Abdeel to arrest Baruch the scribe and Jeremiah the prophet. But the LORD had hidden them.
JER|36|27|After the king burned the scroll containing the words that Baruch had written at Jeremiah's dictation, the word of the LORD came to Jeremiah:
JER|36|28|"Take another scroll and write on it all the words that were on the first scroll, which Jehoiakim king of Judah burned up.
JER|36|29|Also tell Jehoiakim king of Judah, 'This is what the LORD says: You burned that scroll and said, "Why did you write on it that the king of Babylon would certainly come and destroy this land and cut off both men and animals from it?"
JER|36|30|Therefore, this is what the LORD says about Jehoiakim king of Judah: He will have no one to sit on the throne of David; his body will be thrown out and exposed to the heat by day and the frost by night.
JER|36|31|I will punish him and his children and his attendants for their wickedness; I will bring on them and those living in Jerusalem and the people of Judah every disaster I pronounced against them, because they have not listened.'"
JER|36|32|So Jeremiah took another scroll and gave it to the scribe Baruch son of Neriah, and as Jeremiah dictated, Baruch wrote on it all the words of the scroll that Jehoiakim king of Judah had burned in the fire. And many similar words were added to them.
JER|37|1|Zedekiah son of Josiah was made king of Judah by Nebuchadnezzar king of Babylon; he reigned in place of Jehoiachin son of Jehoiakim.
JER|37|2|Neither he nor his attendants nor the people of the land paid any attention to the words the LORD had spoken through Jeremiah the prophet.
JER|37|3|King Zedekiah, however, sent Jehucal son of Shelemiah with the priest Zephaniah son of Maaseiah to Jeremiah the prophet with this message: "Please pray to the LORD our God for us."
JER|37|4|Now Jeremiah was free to come and go among the people, for he had not yet been put in prison.
JER|37|5|Pharaoh's army had marched out of Egypt, and when the Babylonians who were besieging Jerusalem heard the report about them, they withdrew from Jerusalem.
JER|37|6|Then the word of the LORD came to Jeremiah the prophet:
JER|37|7|"This is what the LORD, the God of Israel, says: Tell the king of Judah, who sent you to inquire of me, 'Pharaoh's army, which has marched out to support you, will go back to its own land, to Egypt.
JER|37|8|Then the Babylonians will return and attack this city; they will capture it and burn it down.'
JER|37|9|"This is what the LORD says: Do not deceive yourselves, thinking, 'The Babylonians will surely leave us.' They will not!
JER|37|10|Even if you were to defeat the entire Babylonian army that is attacking you and only wounded men were left in their tents, they would come out and burn this city down."
JER|37|11|After the Babylonian army had withdrawn from Jerusalem because of Pharaoh's army,
JER|37|12|Jeremiah started to leave the city to go to the territory of Benjamin to get his share of the property among the people there.
JER|37|13|But when he reached the Benjamin Gate, the captain of the guard, whose name was Irijah son of Shelemiah, the son of Hananiah, arrested him and said, "You are deserting to the Babylonians!"
JER|37|14|"That's not true!" Jeremiah said. "I am not deserting to the Babylonians." But Irijah would not listen to him; instead, he arrested Jeremiah and brought him to the officials.
JER|37|15|They were angry with Jeremiah and had him beaten and imprisoned in the house of Jonathan the secretary, which they had made into a prison.
JER|37|16|Jeremiah was put into a vaulted cell in a dungeon, where he remained a long time.
JER|37|17|Then King Zedekiah sent for him and had him brought to the palace, where he asked him privately, "Is there any word from the LORD?Yes," Jeremiah replied, "you will be handed over to the king of Babylon."
JER|37|18|Then Jeremiah said to King Zedekiah, "What crime have I committed against you or your officials or this people, that you have put me in prison?
JER|37|19|Where are your prophets who prophesied to you, 'The king of Babylon will not attack you or this land'?
JER|37|20|But now, my lord the king, please listen. Let me bring my petition before you: Do not send me back to the house of Jonathan the secretary, or I will die there."
JER|37|21|King Zedekiah then gave orders for Jeremiah to be placed in the courtyard of the guard and given bread from the street of the bakers each day until all the bread in the city was gone. So Jeremiah remained in the courtyard of the guard.
JER|38|1|Shephatiah son of Mattan, Gedaliah son of Pashhur, Jehucal son of Shelemiah, and Pashhur son of Malkijah heard what Jeremiah was telling all the people when he said,
JER|38|2|"This is what the LORD says: 'Whoever stays in this city will die by the sword, famine or plague, but whoever goes over to the Babylonians will live. He will escape with his life; he will live.'
JER|38|3|And this is what the LORD says: 'This city will certainly be handed over to the army of the king of Babylon, who will capture it.'"
JER|38|4|Then the officials said to the king, "This man should be put to death. He is discouraging the soldiers who are left in this city, as well as all the people, by the things he is saying to them. This man is not seeking the good of these people but their ruin."
JER|38|5|"He is in your hands," King Zedekiah answered. "The king can do nothing to oppose you."
JER|38|6|So they took Jeremiah and put him into the cistern of Malkijah, the king's son, which was in the courtyard of the guard. They lowered Jeremiah by ropes into the cistern; it had no water in it, only mud, and Jeremiah sank down into the mud.
JER|38|7|But Ebed-Melech, a Cushite, an official in the royal palace, heard that they had put Jeremiah into the cistern. While the king was sitting in the Benjamin Gate,
JER|38|8|Ebed-Melech went out of the palace and said to him,
JER|38|9|"My lord the king, these men have acted wickedly in all they have done to Jeremiah the prophet. They have thrown him into a cistern, where he will starve to death when there is no longer any bread in the city."
JER|38|10|Then the king commanded Ebed-Melech the Cushite, "Take thirty men from here with you and lift Jeremiah the prophet out of the cistern before he dies."
JER|38|11|So Ebed-Melech took the men with him and went to a room under the treasury in the palace. He took some old rags and worn-out clothes from there and let them down with ropes to Jeremiah in the cistern.
JER|38|12|Ebed-Melech the Cushite said to Jeremiah, "Put these old rags and worn-out clothes under your arms to pad the ropes." Jeremiah did so,
JER|38|13|and they pulled him up with the ropes and lifted him out of the cistern. And Jeremiah remained in the courtyard of the guard.
JER|38|14|Then King Zedekiah sent for Jeremiah the prophet and had him brought to the third entrance to the temple of the LORD. "I am going to ask you something," the king said to Jeremiah. "Do not hide anything from me."
JER|38|15|Jeremiah said to Zedekiah, "If I give you an answer, will you not kill me? Even if I did give you counsel, you would not listen to me."
JER|38|16|But King Zedekiah swore this oath secretly to Jeremiah: "As surely as the LORD lives, who has given us breath, I will neither kill you nor hand you over to those who are seeking your life."
JER|38|17|Then Jeremiah said to Zedekiah, "This is what the LORD God Almighty, the God of Israel, says: 'If you surrender to the officers of the king of Babylon, your life will be spared and this city will not be burned down; you and your family will live.
JER|38|18|But if you will not surrender to the officers of the king of Babylon, this city will be handed over to the Babylonians and they will burn it down; you yourself will not escape from their hands.'"
JER|38|19|King Zedekiah said to Jeremiah, "I am afraid of the Jews who have gone over to the Babylonians, for the Babylonians may hand me over to them and they will mistreat me."
JER|38|20|"They will not hand you over," Jeremiah replied. "Obey the LORD by doing what I tell you. Then it will go well with you, and your life will be spared.
JER|38|21|But if you refuse to surrender, this is what the LORD has revealed to me:
JER|38|22|All the women left in the palace of the king of Judah will be brought out to the officials of the king of Babylon. Those women will say to you: "'They misled you and overcame you- those trusted friends of yours. Your feet are sunk in the mud; your friends have deserted you.'
JER|38|23|"All your wives and children will be brought out to the Babylonians. You yourself will not escape from their hands but will be captured by the king of Babylon; and this city will be burned down."
JER|38|24|Then Zedekiah said to Jeremiah, "Do not let anyone know about this conversation, or you may die.
JER|38|25|If the officials hear that I talked with you, and they come to you and say, 'Tell us what you said to the king and what the king said to you; do not hide it from us or we will kill you,'
JER|38|26|then tell them, 'I was pleading with the king not to send me back to Jonathan's house to die there.'"
JER|38|27|All the officials did come to Jeremiah and question him, and he told them everything the king had ordered him to say. So they said no more to him, for no one had heard his conversation with the king.
JER|38|28|And Jeremiah remained in the courtyard of the guard until the day Jerusalem was captured.
JER|39|1|This is how Jerusalem was taken: In the ninth year of Zedekiah king of Judah, in the tenth month, Nebuchadnezzar king of Babylon marched against Jerusalem with his whole army and laid siege to it.
JER|39|2|And on the ninth day of the fourth month of Zedekiah's eleventh year, the city wall was broken through.
JER|39|3|Then all the officials of the king of Babylon came and took seats in the Middle Gate: Nergal-Sharezer of Samgar, Nebo-Sarsekim a chief officer, Nergal-Sharezer a high official and all the other officials of the king of Babylon.
JER|39|4|When Zedekiah king of Judah and all the soldiers saw them, they fled; they left the city at night by way of the king's garden, through the gate between the two walls, and headed toward the Arabah.
JER|39|5|But the Babylonian army pursued them and overtook Zedekiah in the plains of Jericho. They captured him and took him to Nebuchadnezzar king of Babylon at Riblah in the land of Hamath, where he pronounced sentence on him.
JER|39|6|There at Riblah the king of Babylon slaughtered the sons of Zedekiah before his eyes and also killed all the nobles of Judah.
JER|39|7|Then he put out Zedekiah's eyes and bound him with bronze shackles to take him to Babylon.
JER|39|8|The Babylonians set fire to the royal palace and the houses of the people and broke down the walls of Jerusalem.
JER|39|9|Nebuzaradan commander of the imperial guard carried into exile to Babylon the people who remained in the city, along with those who had gone over to him, and the rest of the people.
JER|39|10|But Nebuzaradan the commander of the guard left behind in the land of Judah some of the poor people, who owned nothing; and at that time he gave them vineyards and fields.
JER|39|11|Now Nebuchadnezzar king of Babylon had given these orders about Jeremiah through Nebuzaradan commander of the imperial guard:
JER|39|12|"Take him and look after him; don't harm him but do for him whatever he asks."
JER|39|13|So Nebuzaradan the commander of the guard, Nebushazban a chief officer, Nergal-Sharezer a high official and all the other officers of the king of Babylon
JER|39|14|sent and had Jeremiah taken out of the courtyard of the guard. They turned him over to Gedaliah son of Ahikam, the son of Shaphan, to take him back to his home. So he remained among his own people.
JER|39|15|While Jeremiah had been confined in the courtyard of the guard, the word of the LORD came to him:
JER|39|16|"Go and tell Ebed-Melech the Cushite, 'This is what the LORD Almighty, the God of Israel, says: I am about to fulfill my words against this city through disaster, not prosperity. At that time they will be fulfilled before your eyes.
JER|39|17|But I will rescue you on that day, declares the LORD; you will not be handed over to those you fear.
JER|39|18|I will save you; you will not fall by the sword but will escape with your life, because you trust in me, declares the LORD.'"
JER|40|1|The word came to Jeremiah from the LORD after Nebuzaradan commander of the imperial guard had released him at Ramah. He had found Jeremiah bound in chains among all the captives from Jerusalem and Judah who were being carried into exile to Babylon.
JER|40|2|When the commander of the guard found Jeremiah, he said to him, "The LORD your God decreed this disaster for this place.
JER|40|3|And now the LORD has brought it about; he has done just as he said he would. All this happened because you people sinned against the LORD and did not obey him.
JER|40|4|But today I am freeing you from the chains on your wrists. Come with me to Babylon, if you like, and I will look after you; but if you do not want to, then don't come. Look, the whole country lies before you; go wherever you please."
JER|40|5|However, before Jeremiah turned to go, Nebuzaradan added, "Go back to Gedaliah son of Ahikam, the son of Shaphan, whom the king of Babylon has appointed over the towns of Judah, and live with him among the people, or go anywhere else you please." Then the commander gave him provisions and a present and let him go.
JER|40|6|So Jeremiah went to Gedaliah son of Ahikam at Mizpah and stayed with him among the people who were left behind in the land.
JER|40|7|When all the army officers and their men who were still in the open country heard that the king of Babylon had appointed Gedaliah son of Ahikam as governor over the land and had put him in charge of the men, women and children who were the poorest in the land and who had not been carried into exile to Babylon,
JER|40|8|they came to Gedaliah at Mizpah-Ishmael son of Nethaniah, Johanan and Jonathan the sons of Kareah, Seraiah son of Tanhumeth, the sons of Ephai the Netophathite, and Jaazaniah the son of the Maacathite, and their men.
JER|40|9|Gedaliah son of Ahikam, the son of Shaphan, took an oath to reassure them and their men. "Do not be afraid to serve the Babylonians, "he said. "Settle down in the land and serve the king of Babylon, and it will go well with you.
JER|40|10|I myself will stay at Mizpah to represent you before the Babylonians who come to us, but you are to harvest the wine, summer fruit and oil, and put them in your storage jars, and live in the towns you have taken over."
JER|40|11|When all the Jews in Moab, Ammon, Edom and all the other countries heard that the king of Babylon had left a remnant in Judah and had appointed Gedaliah son of Ahikam, the son of Shaphan, as governor over them,
JER|40|12|they all came back to the land of Judah, to Gedaliah at Mizpah, from all the countries where they had been scattered. And they harvested an abundance of wine and summer fruit.
JER|40|13|Johanan son of Kareah and all the army officers still in the open country came to Gedaliah at Mizpah
JER|40|14|and said to him, "Don't you know that Baalis king of the Ammonites has sent Ishmael son of Nethaniah to take your life?" But Gedaliah son of Ahikam did not believe them.
JER|40|15|Then Johanan son of Kareah said privately to Gedaliah in Mizpah, "Let me go and kill Ishmael son of Nethaniah, and no one will know it. Why should he take your life and cause all the Jews who are gathered around you to be scattered and the remnant of Judah to perish?"
JER|40|16|But Gedaliah son of Ahikam said to Johanan son of Kareah, "Don't do such a thing! What you are saying about Ishmael is not true."
JER|41|1|In the seventh month Ishmael son of Nethaniah, the son of Elishama, who was of royal blood and had been one of the king's officers, came with ten men to Gedaliah son of Ahikam at Mizpah. While they were eating together there,
JER|41|2|Ishmael son of Nethaniah and the ten men who were with him got up and struck down Gedaliah son of Ahikam, the son of Shaphan, with the sword, killing the one whom the king of Babylon had appointed as governor over the land.
JER|41|3|Ishmael also killed all the Jews who were with Gedaliah at Mizpah, as well as the Babylonian soldiers who were there.
JER|41|4|The day after Gedaliah's assassination, before anyone knew about it,
JER|41|5|eighty men who had shaved off their beards, torn their clothes and cut themselves came from Shechem, Shiloh and Samaria, bringing grain offerings and incense with them to the house of the LORD.
JER|41|6|Ishmael son of Nethaniah went out from Mizpah to meet them, weeping as he went. When he met them, he said, "Come to Gedaliah son of Ahikam."
JER|41|7|When they went into the city, Ishmael son of Nethaniah and the men who were with him slaughtered them and threw them into a cistern.
JER|41|8|But ten of them said to Ishmael, "Don't kill us! We have wheat and barley, oil and honey, hidden in a field." So he let them alone and did not kill them with the others.
JER|41|9|Now the cistern where he threw all the bodies of the men he had killed along with Gedaliah was the one King Asa had made as part of his defense against Baasha king of Israel. Ishmael son of Nethaniah filled it with the dead.
JER|41|10|Ishmael made captives of all the rest of the people who were in Mizpah-the king's daughters along with all the others who were left there, over whom Nebuzaradan commander of the imperial guard had appointed Gedaliah son of Ahikam. Ishmael son of Nethaniah took them captive and set out to cross over to the Ammonites.
JER|41|11|When Johanan son of Kareah and all the army officers who were with him heard about all the crimes Ishmael son of Nethaniah had committed,
JER|41|12|they took all their men and went to fight Ishmael son of Nethaniah. They caught up with him near the great pool in Gibeon.
JER|41|13|When all the people Ishmael had with him saw Johanan son of Kareah and the army officers who were with him, they were glad.
JER|41|14|All the people Ishmael had taken captive at Mizpah turned and went over to Johanan son of Kareah.
JER|41|15|But Ishmael son of Nethaniah and eight of his men escaped from Johanan and fled to the Ammonites.
JER|41|16|Then Johanan son of Kareah and all the army officers who were with him led away all the survivors from Mizpah whom he had recovered from Ishmael son of Nethaniah after he had assassinated Gedaliah son of Ahikam: the soldiers, women, children and court officials he had brought from Gibeon.
JER|41|17|And they went on, stopping at Geruth Kimham near Bethlehem on their way to Egypt
JER|41|18|to escape the Babylonians. They were afraid of them because Ishmael son of Nethaniah had killed Gedaliah son of Ahikam, whom the king of Babylon had appointed as governor over the land.
JER|42|1|Then all the army officers, including Johanan son of Kareah and Jezaniah son of Hoshaiah, and all the people from the least to the greatest approached
JER|42|2|Jeremiah the prophet and said to him, "Please hear our petition and pray to the LORD your God for this entire remnant. For as you now see, though we were once many, now only a few are left.
JER|42|3|Pray that the LORD your God will tell us where we should go and what we should do."
JER|42|4|"I have heard you," replied Jeremiah the prophet. "I will certainly pray to the LORD your God as you have requested; I will tell you everything the LORD says and will keep nothing back from you."
JER|42|5|Then they said to Jeremiah, "May the LORD be a true and faithful witness against us if we do not act in accordance with everything the LORD your God sends you to tell us.
JER|42|6|Whether it is favorable or unfavorable, we will obey the LORD our God, to whom we are sending you, so that it will go well with us, for we will obey the LORD our God."
JER|42|7|Ten days later the word of the LORD came to Jeremiah.
JER|42|8|So he called together Johanan son of Kareah and all the army officers who were with him and all the people from the least to the greatest.
JER|42|9|He said to them, "This is what the LORD, the God of Israel, to whom you sent me to present your petition, says:
JER|42|10|'If you stay in this land, I will build you up and not tear you down; I will plant you and not uproot you, for I am grieved over the disaster I have inflicted on you.
JER|42|11|Do not be afraid of the king of Babylon, whom you now fear. Do not be afraid of him, declares the LORD, for I am with you and will save you and deliver you from his hands.
JER|42|12|I will show you compassion so that he will have compassion on you and restore you to your land.'
JER|42|13|"However, if you say, 'We will not stay in this land,' and so disobey the LORD your God,
JER|42|14|and if you say, 'No, we will go and live in Egypt, where we will not see war or hear the trumpet or be hungry for bread,'
JER|42|15|then hear the word of the LORD, O remnant of Judah. This is what the LORD Almighty, the God of Israel, says: 'If you are determined to go to Egypt and you do go to settle there,
JER|42|16|then the sword you fear will overtake you there, and the famine you dread will follow you into Egypt, and there you will die.
JER|42|17|Indeed, all who are determined to go to Egypt to settle there will die by the sword, famine and plague; not one of them will survive or escape the disaster I will bring on them.'
JER|42|18|This is what the LORD Almighty, the God of Israel, says: 'As my anger and wrath have been poured out on those who lived in Jerusalem, so will my wrath be poured out on you when you go to Egypt. You will be an object of cursing and horror, of condemnation and reproach; you will never see this place again.'
JER|42|19|"O remnant of Judah, the LORD has told you, 'Do not go to Egypt.' Be sure of this: I warn you today
JER|42|20|that you made a fatal mistake when you sent me to the LORD your God and said, 'Pray to the LORD our God for us; tell us everything he says and we will do it.'
JER|42|21|I have told you today, but you still have not obeyed the LORD your God in all he sent me to tell you.
JER|42|22|So now, be sure of this: You will die by the sword, famine and plague in the place where you want to go to settle."
JER|43|1|When Jeremiah finished telling the people all the words of the LORD their God-everything the LORD had sent him to tell them-
JER|43|2|Azariah son of Hoshaiah and Johanan son of Kareah and all the arrogant men said to Jeremiah, "You are lying! The LORD our God has not sent you to say, 'You must not go to Egypt to settle there.'
JER|43|3|But Baruch son of Neriah is inciting you against us to hand us over to the Babylonians, so they may kill us or carry us into exile to Babylon."
JER|43|4|So Johanan son of Kareah and all the army officers and all the people disobeyed the LORD's command to stay in the land of Judah.
JER|43|5|Instead, Johanan son of Kareah and all the army officers led away all the remnant of Judah who had come back to live in the land of Judah from all the nations where they had been scattered.
JER|43|6|They also led away all the men, women and children and the king's daughters whom Nebuzaradan commander of the imperial guard had left with Gedaliah son of Ahikam, the son of Shaphan, and Jeremiah the prophet and Baruch son of Neriah.
JER|43|7|So they entered Egypt in disobedience to the LORD and went as far as Tahpanhes.
JER|43|8|In Tahpanhes the word of the LORD came to Jeremiah:
JER|43|9|"While the Jews are watching, take some large stones with you and bury them in clay in the brick pavement at the entrance to Pharaoh's palace in Tahpanhes.
JER|43|10|Then say to them, 'This is what the LORD Almighty, the God of Israel, says: I will send for my servant Nebuchadnezzar king of Babylon, and I will set his throne over these stones I have buried here; he will spread his royal canopy above them.
JER|43|11|He will come and attack Egypt, bringing death to those destined for death, captivity to those destined for captivity, and the sword to those destined for the sword.
JER|43|12|He will set fire to the temples of the gods of Egypt; he will burn their temples and take their gods captive. As a shepherd wraps his garment around him, so will he wrap Egypt around himself and depart from there unscathed.
JER|43|13|There in the temple of the sun in Egypt he will demolish the sacred pillars and will burn down the temples of the gods of Egypt.'"
JER|44|1|This word came to Jeremiah concerning all the Jews living in Lower Egypt-in Migdol, Tahpanhes and Memphis -and in Upper Egypt:
JER|44|2|"This is what the LORD Almighty, the God of Israel, says: You saw the great disaster I brought on Jerusalem and on all the towns of Judah. Today they lie deserted and in ruins
JER|44|3|because of the evil they have done. They provoked me to anger by burning incense and by worshiping other gods that neither they nor you nor your fathers ever knew.
JER|44|4|Again and again I sent my servants the prophets, who said, 'Do not do this detestable thing that I hate!'
JER|44|5|But they did not listen or pay attention; they did not turn from their wickedness or stop burning incense to other gods.
JER|44|6|Therefore, my fierce anger was poured out; it raged against the towns of Judah and the streets of Jerusalem and made them the desolate ruins they are today.
JER|44|7|"Now this is what the LORD God Almighty, the God of Israel, says: Why bring such great disaster on yourselves by cutting off from Judah the men and women, the children and infants, and so leave yourselves without a remnant?
JER|44|8|Why provoke me to anger with what your hands have made, burning incense to other gods in Egypt, where you have come to live? You will destroy yourselves and make yourselves an object of cursing and reproach among all the nations on earth.
JER|44|9|Have you forgotten the wickedness committed by your fathers and by the kings and queens of Judah and the wickedness committed by you and your wives in the land of Judah and the streets of Jerusalem?
JER|44|10|To this day they have not humbled themselves or shown reverence, nor have they followed my law and the decrees I set before you and your fathers.
JER|44|11|"Therefore, this is what the LORD Almighty, the God of Israel, says: I am determined to bring disaster on you and to destroy all Judah.
JER|44|12|I will take away the remnant of Judah who were determined to go to Egypt to settle there. They will all perish in Egypt; they will fall by the sword or die from famine. From the least to the greatest, they will die by sword or famine. They will become an object of cursing and horror, of condemnation and reproach.
JER|44|13|I will punish those who live in Egypt with the sword, famine and plague, as I punished Jerusalem.
JER|44|14|None of the remnant of Judah who have gone to live in Egypt will escape or survive to return to the land of Judah, to which they long to return and live; none will return except a few fugitives."
JER|44|15|Then all the men who knew that their wives were burning incense to other gods, along with all the women who were present-a large assembly-and all the people living in Lower and Upper Egypt, said to Jeremiah,
JER|44|16|"We will not listen to the message you have spoken to us in the name of the LORD!
JER|44|17|We will certainly do everything we said we would: We will burn incense to the Queen of Heaven and will pour out drink offerings to her just as we and our fathers, our kings and our officials did in the towns of Judah and in the streets of Jerusalem. At that time we had plenty of food and were well off and suffered no harm.
JER|44|18|But ever since we stopped burning incense to the Queen of Heaven and pouring out drink offerings to her, we have had nothing and have been perishing by sword and famine."
JER|44|19|The women added, "When we burned incense to the Queen of Heaven and poured out drink offerings to her, did not our husbands know that we were making cakes like her image and pouring out drink offerings to her?"
JER|44|20|Then Jeremiah said to all the people, both men and women, who were answering him,
JER|44|21|"Did not the LORD remember and think about the incense burned in the towns of Judah and the streets of Jerusalem by you and your fathers, your kings and your officials and the people of the land?
JER|44|22|When the LORD could no longer endure your wicked actions and the detestable things you did, your land became an object of cursing and a desolate waste without inhabitants, as it is today.
JER|44|23|Because you have burned incense and have sinned against the LORD and have not obeyed him or followed his law or his decrees or his stipulations, this disaster has come upon you, as you now see."
JER|44|24|Then Jeremiah said to all the people, including the women, "Hear the word of the LORD, all you people of Judah in Egypt.
JER|44|25|This is what the LORD Almighty, the God of Israel, says: You and your wives have shown by your actions what you promised when you said, 'We will certainly carry out the vows we made to burn incense and pour out drink offerings to the Queen of Heaven.'"Go ahead then, do what you promised! Keep your vows!
JER|44|26|But hear the word of the LORD, all Jews living in Egypt: 'I swear by my great name,' says the LORD, 'that no one from Judah living anywhere in Egypt will ever again invoke my name or swear, "As surely as the Sovereign LORD lives."
JER|44|27|For I am watching over them for harm, not for good; the Jews in Egypt will perish by sword and famine until they are all destroyed.
JER|44|28|Those who escape the sword and return to the land of Judah from Egypt will be very few. Then the whole remnant of Judah who came to live in Egypt will know whose word will stand-mine or theirs.
JER|44|29|"'This will be the sign to you that I will punish you in this place,' declares the LORD, 'so that you will know that my threats of harm against you will surely stand.'
JER|44|30|This is what the LORD says: 'I am going to hand Pharaoh Hophra king of Egypt over to his enemies who seek his life, just as I handed Zedekiah king of Judah over to Nebuchadnezzar king of Babylon, the enemy who was seeking his life.'"
JER|45|1|This is what Jeremiah the prophet told Baruch son of Neriah in the fourth year of Jehoiakim son of Josiah king of Judah, after Baruch had written on a scroll the words Jeremiah was then dictating:
JER|45|2|"This is what the LORD, the God of Israel, says to you, Baruch:
JER|45|3|You said, 'Woe to me! The LORD has added sorrow to my pain; I am worn out with groaning and find no rest.'"
JER|45|4|The LORD said, "Say this to him: 'This is what the LORD says: I will overthrow what I have built and uproot what I have planted, throughout the land.
JER|45|5|Should you then seek great things for yourself? Seek them not. For I will bring disaster on all people, declares the LORD, but wherever you go I will let you escape with your life.'"
JER|46|1|This is the word of the LORD that came to Jeremiah the prophet concerning the nations:
JER|46|2|Concerning Egypt: This is the message against the army of Pharaoh Neco king of Egypt, which was defeated at Carchemish on the Euphrates River by Nebuchadnezzar king of Babylon in the fourth year of Jehoiakim son of Josiah king of Judah:
JER|46|3|"Prepare your shields, both large and small, and march out for battle!
JER|46|4|Harness the horses, mount the steeds! Take your positions with helmets on! Polish your spears, put on your armor!
JER|46|5|What do I see? They are terrified, they are retreating, their warriors are defeated. They flee in haste without looking back, and there is terror on every side," declares the LORD.
JER|46|6|"The swift cannot flee nor the strong escape. In the north by the River Euphrates they stumble and fall.
JER|46|7|"Who is this that rises like the Nile, like rivers of surging waters?
JER|46|8|Egypt rises like the Nile, like rivers of surging waters. She says, 'I will rise and cover the earth; I will destroy cities and their people.'
JER|46|9|Charge, O horses! Drive furiously, O charioteers! March on, O warriors- men of Cush and Put who carry shields, men of Lydia who draw the bow.
JER|46|10|But that day belongs to the LORD, the Lord Almighty- a day of vengeance, for vengeance on his foes. The sword will devour till it is satisfied, till it has quenched its thirst with blood. For the Lord, the LORD Almighty, will offer sacrifice in the land of the north by the River Euphrates.
JER|46|11|"Go up to Gilead and get balm, O Virgin Daughter of Egypt. But you multiply remedies in vain; there is no healing for you.
JER|46|12|The nations will hear of your shame; your cries will fill the earth. One warrior will stumble over another; both will fall down together."
JER|46|13|This is the message the LORD spoke to Jeremiah the prophet about the coming of Nebuchadnezzar king of Babylon to attack Egypt:
JER|46|14|"Announce this in Egypt, and proclaim it in Migdol; proclaim it also in Memphis and Tahpanhes: 'Take your positions and get ready, for the sword devours those around you.'
JER|46|15|Why will your warriors be laid low? They cannot stand, for the LORD will push them down.
JER|46|16|They will stumble repeatedly; they will fall over each other. They will say, 'Get up, let us go back to our own people and our native lands, away from the sword of the oppressor.'
JER|46|17|There they will exclaim, 'Pharaoh king of Egypt is only a loud noise; he has missed his opportunity.'
JER|46|18|"As surely as I live," declares the King, whose name is the LORD Almighty, "one will come who is like Tabor among the mountains, like Carmel by the sea.
JER|46|19|Pack your belongings for exile, you who live in Egypt, for Memphis will be laid waste and lie in ruins without inhabitant.
JER|46|20|"Egypt is a beautiful heifer, but a gadfly is coming against her from the north.
JER|46|21|The mercenaries in her ranks are like fattened calves. They too will turn and flee together, they will not stand their ground, for the day of disaster is coming upon them, the time for them to be punished.
JER|46|22|Egypt will hiss like a fleeing serpent as the enemy advances in force; they will come against her with axes, like men who cut down trees.
JER|46|23|They will chop down her forest," declares the LORD, "dense though it be. They are more numerous than locusts, they cannot be counted.
JER|46|24|The Daughter of Egypt will be put to shame, handed over to the people of the north."
JER|46|25|The LORD Almighty, the God of Israel, says: "I am about to bring punishment on Amon god of Thebes, on Pharaoh, on Egypt and her gods and her kings, and on those who rely on Pharaoh.
JER|46|26|I will hand them over to those who seek their lives, to Nebuchadnezzar king of Babylon and his officers. Later, however, Egypt will be inhabited as in times past," declares the LORD.
JER|46|27|"Do not fear, O Jacob my servant; do not be dismayed, O Israel. I will surely save you out of a distant place, your descendants from the land of their exile. Jacob will again have peace and security, and no one will make him afraid.
JER|46|28|Do not fear, O Jacob my servant, for I am with you," declares the LORD. "Though I completely destroy all the nations among which I scatter you, I will not completely destroy you. I will discipline you but only with justice; I will not let you go entirely unpunished."
JER|47|1|This is the word of the LORD that came to Jeremiah the prophet concerning the Philistines before Pharaoh attacked Gaza:
JER|47|2|This is what the LORD says: "See how the waters are rising in the north; they will become an overflowing torrent. They will overflow the land and everything in it, the towns and those who live in them. The people will cry out; all who dwell in the land will wail
JER|47|3|at the sound of the hoofs of galloping steeds, at the noise of enemy chariots and the rumble of their wheels. Fathers will not turn to help their children; their hands will hang limp.
JER|47|4|For the day has come to destroy all the Philistines and to cut off all survivors who could help Tyre and Sidon. The LORD is about to destroy the Philistines, the remnant from the coasts of Caphtor.
JER|47|5|Gaza will shave her head in mourning; Ashkelon will be silenced. O remnant on the plain, how long will you cut yourselves?
JER|47|6|"'Ah, sword of the LORD,' you cry, 'how long till you rest? Return to your scabbard; cease and be still.'
JER|47|7|But how can it rest when the LORD has commanded it, when he has ordered it to attack Ashkelon and the coast?"
JER|48|1|Concerning Moab: This is what the LORD Almighty, the God of Israel, says: "Woe to Nebo, for it will be ruined. Kiriathaim will be disgraced and captured; the stronghold will be disgraced and shattered.
JER|48|2|Moab will be praised no more; in Heshbon men will plot her downfall: 'Come, let us put an end to that nation.' You too, O Madmen, will be silenced; the sword will pursue you.
JER|48|3|Listen to the cries from Horonaim, cries of great havoc and destruction.
JER|48|4|Moab will be broken; her little ones will cry out.
JER|48|5|They go up the way to Luhith, weeping bitterly as they go; on the road down to Horonaim anguished cries over the destruction are heard.
JER|48|6|Flee! Run for your lives; become like a bush in the desert.
JER|48|7|Since you trust in your deeds and riches, you too will be taken captive, and Chemosh will go into exile, together with his priests and officials.
JER|48|8|The destroyer will come against every town, and not a town will escape. The valley will be ruined and the plateau destroyed, because the LORD has spoken.
JER|48|9|Put salt on Moab, for she will be laid waste; her towns will become desolate, with no one to live in them.
JER|48|10|"A curse on him who is lax in doing the LORD's work! A curse on him who keeps his sword from bloodshed!
JER|48|11|"Moab has been at rest from youth, like wine left on its dregs, not poured from one jar to another- she has not gone into exile. So she tastes as she did, and her aroma is unchanged.
JER|48|12|But days are coming," declares the LORD, "when I will send men who pour from jars, and they will pour her out; they will empty her jars and smash her jugs.
JER|48|13|Then Moab will be ashamed of Chemosh, as the house of Israel was ashamed when they trusted in Bethel.
JER|48|14|"How can you say, 'We are warriors, men valiant in battle'?
JER|48|15|Moab will be destroyed and her towns invaded; her finest young men will go down in the slaughter," declares the King, whose name is the LORD Almighty.
JER|48|16|"The fall of Moab is at hand; her calamity will come quickly.
JER|48|17|Mourn for her, all who live around her, all who know her fame; say, 'How broken is the mighty scepter, how broken the glorious staff!'
JER|48|18|"Come down from your glory and sit on the parched ground, O inhabitants of the Daughter of Dibon, for he who destroys Moab will come up against you and ruin your fortified cities.
JER|48|19|Stand by the road and watch, you who live in Aroer. Ask the man fleeing and the woman escaping, ask them, 'What has happened?'
JER|48|20|Moab is disgraced, for she is shattered. Wail and cry out! Announce by the Arnon that Moab is destroyed.
JER|48|21|Judgment has come to the plateau- to Holon, Jahzah and Mephaath,
JER|48|22|to Dibon, Nebo and Beth Diblathaim,
JER|48|23|to Kiriathaim, Beth Gamul and Beth Meon,
JER|48|24|to Kerioth and Bozrah- to all the towns of Moab, far and near.
JER|48|25|Moab's horn is cut off; her arm is broken," declares the LORD.
JER|48|26|"Make her drunk, for she has defied the LORD. Let Moab wallow in her vomit; let her be an object of ridicule.
JER|48|27|Was not Israel the object of your ridicule? Was she caught among thieves, that you shake your head in scorn whenever you speak of her?
JER|48|28|Abandon your towns and dwell among the rocks, you who live in Moab. Be like a dove that makes its nest at the mouth of a cave.
JER|48|29|"We have heard of Moab's pride- her overweening pride and conceit, her pride and arrogance and the haughtiness of her heart.
JER|48|30|I know her insolence but it is futile," declares the LORD, "and her boasts accomplish nothing.
JER|48|31|Therefore I wail over Moab, for all Moab I cry out, I moan for the men of Kir Hareseth.
JER|48|32|I weep for you, as Jazer weeps, O vines of Sibmah. Your branches spread as far as the sea; they reached as far as the sea of Jazer. The destroyer has fallen on your ripened fruit and grapes.
JER|48|33|Joy and gladness are gone from the orchards and fields of Moab. I have stopped the flow of wine from the presses; no one treads them with shouts of joy. Although there are shouts, they are not shouts of joy.
JER|48|34|"The sound of their cry rises from Heshbon to Elealeh and Jahaz, from Zoar as far as Horonaim and Eglath Shelishiyah, for even the waters of Nimrim are dried up.
JER|48|35|In Moab I will put an end to those who make offerings on the high places and burn incense to their gods," declares the LORD.
JER|48|36|"So my heart laments for Moab like a flute; it laments like a flute for the men of Kir Hareseth. The wealth they acquired is gone.
JER|48|37|Every head is shaved and every beard cut off; every hand is slashed and every waist is covered with sackcloth.
JER|48|38|On all the roofs in Moab and in the public squares there is nothing but mourning, for I have broken Moab like a jar that no one wants," declares the LORD.
JER|48|39|"How shattered she is! How they wail! How Moab turns her back in shame! Moab has become an object of ridicule, an object of horror to all those around her."
JER|48|40|This is what the LORD says: "Look! An eagle is swooping down, spreading its wings over Moab.
JER|48|41|Kerioth will be captured and the strongholds taken. In that day the hearts of Moab's warriors will be like the heart of a woman in labor.
JER|48|42|Moab will be destroyed as a nation because she defied the LORD.
JER|48|43|Terror and pit and snare await you, O people of Moab," declares the LORD.
JER|48|44|"Whoever flees from the terror will fall into a pit, whoever climbs out of the pit will be caught in a snare; for I will bring upon Moab the year of her punishment," declares the LORD.
JER|48|45|"In the shadow of Heshbon the fugitives stand helpless, for a fire has gone out from Heshbon, a blaze from the midst of Sihon; it burns the foreheads of Moab, the skulls of the noisy boasters.
JER|48|46|Woe to you, O Moab! The people of Chemosh are destroyed; your sons are taken into exile and your daughters into captivity.
JER|48|47|"Yet I will restore the fortunes of Moab in days to come," declares the LORD. Here ends the judgment on Moab.
JER|49|1|Concerning the Ammonites: This is what the LORD says: "Has Israel no sons? Has she no heirs? Why then has Molech taken possession of Gad? Why do his people live in its towns?
JER|49|2|But the days are coming," declares the LORD, "when I will sound the battle cry against Rabbah of the Ammonites; it will become a mound of ruins, and its surrounding villages will be set on fire. Then Israel will drive out those who drove her out," says the LORD.
JER|49|3|"Wail, O Heshbon, for Ai is destroyed! Cry out, O inhabitants of Rabbah! Put on sackcloth and mourn; rush here and there inside the walls, for Molech will go into exile, together with his priests and officials.
JER|49|4|Why do you boast of your valleys, boast of your valleys so fruitful? O unfaithful daughter, you trust in your riches and say, 'Who will attack me?'
JER|49|5|I will bring terror on you from all those around you," declares the Lord, the LORD Almighty. "Every one of you will be driven away, and no one will gather the fugitives.
JER|49|6|"Yet afterward, I will restore the fortunes of the Ammonites," declares the LORD.
JER|49|7|Concerning Edom: This is what the LORD Almighty says: "Is there no longer wisdom in Teman? Has counsel perished from the prudent? Has their wisdom decayed?
JER|49|8|Turn and flee, hide in deep caves, you who live in Dedan, for I will bring disaster on Esau at the time I punish him.
JER|49|9|If grape pickers came to you, would they not leave a few grapes? If thieves came during the night, would they not steal only as much as they wanted?
JER|49|10|But I will strip Esau bare; I will uncover his hiding places, so that he cannot conceal himself. His children, relatives and neighbors will perish, and he will be no more.
JER|49|11|Leave your orphans; I will protect their lives. Your widows too can trust in me."
JER|49|12|This is what the LORD says: "If those who do not deserve to drink the cup must drink it, why should you go unpunished? You will not go unpunished, but must drink it.
JER|49|13|I swear by myself," declares the LORD, "that Bozrah will become a ruin and an object of horror, of reproach and of cursing; and all its towns will be in ruins forever."
JER|49|14|I have heard a message from the LORD: An envoy was sent to the nations to say, "Assemble yourselves to attack it! Rise up for battle!"
JER|49|15|"Now I will make you small among the nations, despised among men.
JER|49|16|The terror you inspire and the pride of your heart have deceived you, you who live in the clefts of the rocks, who occupy the heights of the hill. Though you build your nest as high as the eagle's, from there I will bring you down," declares the LORD.
JER|49|17|"Edom will become an object of horror; all who pass by will be appalled and will scoff because of all its wounds.
JER|49|18|As Sodom and Gomorrah were overthrown, along with their neighboring towns," says the LORD, "so no one will live there; no man will dwell in it.
JER|49|19|"Like a lion coming up from Jordan's thickets to a rich pastureland, I will chase Edom from its land in an instant. Who is the chosen one I will appoint for this? Who is like me and who can challenge me? And what shepherd can stand against me?"
JER|49|20|Therefore, hear what the LORD has planned against Edom, what he has purposed against those who live in Teman: The young of the flock will be dragged away; he will completely destroy their pasture because of them.
JER|49|21|At the sound of their fall the earth will tremble; their cry will resound to the Red Sea.
JER|49|22|Look! An eagle will soar and swoop down, spreading its wings over Bozrah. In that day the hearts of Edom's warriors will be like the heart of a woman in labor.
JER|49|23|Concerning Damascus: "Hamath and Arpad are dismayed, for they have heard bad news. They are disheartened, troubled like the restless sea.
JER|49|24|Damascus has become feeble, she has turned to flee and panic has gripped her; anguish and pain have seized her, pain like that of a woman in labor.
JER|49|25|Why has the city of renown not been abandoned, the town in which I delight?
JER|49|26|Surely, her young men will fall in the streets; all her soldiers will be silenced in that day," declares the LORD Almighty.
JER|49|27|"I will set fire to the walls of Damascus; it will consume the fortresses of Ben-Hadad."
JER|49|28|Concerning Kedar and the kingdoms of Hazor, which Nebuchadnezzar king of Babylon attacked: This is what the LORD says: "Arise, and attack Kedar and destroy the people of the East.
JER|49|29|Their tents and their flocks will be taken; their shelters will be carried off with all their goods and camels. Men will shout to them, 'Terror on every side!'
JER|49|30|"Flee quickly away! Stay in deep caves, you who live in Hazor," declares the LORD. "Nebuchadnezzar king of Babylon has plotted against you; he has devised a plan against you.
JER|49|31|"Arise and attack a nation at ease, which lives in confidence," declares the LORD, "a nation that has neither gates nor bars; its people live alone.
JER|49|32|Their camels will become plunder, and their large herds will be booty. I will scatter to the winds those who are in distant places and will bring disaster on them from every side," declares the LORD.
JER|49|33|"Hazor will become a haunt of jackals, a desolate place forever. No one will live there; no man will dwell in it."
JER|49|34|This is the word of the LORD that came to Jeremiah the prophet concerning Elam, early in the reign of Zedekiah king of Judah:
JER|49|35|This is what the LORD Almighty says: "See, I will break the bow of Elam, the mainstay of their might.
JER|49|36|I will bring against Elam the four winds from the four quarters of the heavens; I will scatter them to the four winds, and there will not be a nation where Elam's exiles do not go.
JER|49|37|I will shatter Elam before their foes, before those who seek their lives; I will bring disaster upon them, even my fierce anger," declares the LORD. "I will pursue them with the sword until I have made an end of them.
JER|49|38|I will set my throne in Elam and destroy her king and officials," declares the LORD.
JER|49|39|"Yet I will restore the fortunes of Elam in days to come," declares the LORD.
JER|50|1|This is the word the LORD spoke through Jeremiah the prophet concerning Babylon and the land of the Babylonians:
JER|50|2|"Announce and proclaim among the nations, lift up a banner and proclaim it; keep nothing back, but say, 'Babylon will be captured; Bel will be put to shame, Marduk filled with terror. Her images will be put to shame and her idols filled with terror.'
JER|50|3|A nation from the north will attack her and lay waste her land. No one will live in it; both men and animals will flee away.
JER|50|4|"In those days, at that time," declares the LORD, "the people of Israel and the people of Judah together will go in tears to seek the LORD their God.
JER|50|5|They will ask the way to Zion and turn their faces toward it. They will come and bind themselves to the LORD in an everlasting covenant that will not be forgotten.
JER|50|6|"My people have been lost sheep; their shepherds have led them astray and caused them to roam on the mountains. They wandered over mountain and hill and forgot their own resting place.
JER|50|7|Whoever found them devoured them; their enemies said, 'We are not guilty, for they sinned against the LORD, their true pasture, the LORD, the hope of their fathers.'
JER|50|8|"Flee out of Babylon; leave the land of the Babylonians, and be like the goats that lead the flock.
JER|50|9|For I will stir up and bring against Babylon an alliance of great nations from the land of the north. They will take up their positions against her, and from the north she will be captured. Their arrows will be like skilled warriors who do not return empty-handed.
JER|50|10|So Babylonia will be plundered; all who plunder her will have their fill," declares the LORD.
JER|50|11|"Because you rejoice and are glad, you who pillage my inheritance, because you frolic like a heifer threshing grain and neigh like stallions,
JER|50|12|your mother will be greatly ashamed; she who gave you birth will be disgraced. She will be the least of the nations- a wilderness, a dry land, a desert.
JER|50|13|Because of the LORD's anger she will not be inhabited but will be completely desolate. All who pass Babylon will be horrified and scoff because of all her wounds.
JER|50|14|"Take up your positions around Babylon, all you who draw the bow. Shoot at her! Spare no arrows, for she has sinned against the LORD.
JER|50|15|Shout against her on every side! She surrenders, her towers fall, her walls are torn down. Since this is the vengeance of the LORD, take vengeance on her; do to her as she has done to others.
JER|50|16|Cut off from Babylon the sower, and the reaper with his sickle at harvest. Because of the sword of the oppressor let everyone return to his own people, let everyone flee to his own land.
JER|50|17|"Israel is a scattered flock that lions have chased away. The first to devour him was the king of Assyria; the last to crush his bones was Nebuchadnezzar king of Babylon."
JER|50|18|Therefore this is what the LORD Almighty, the God of Israel, says: "I will punish the king of Babylon and his land as I punished the king of Assyria.
JER|50|19|But I will bring Israel back to his own pasture and he will graze on Carmel and Bashan; his appetite will be satisfied on the hills of Ephraim and Gilead.
JER|50|20|In those days, at that time," declares the LORD, "search will be made for Israel's guilt, but there will be none, and for the sins of Judah, but none will be found, for I will forgive the remnant I spare.
JER|50|21|"Attack the land of Merathaim and those who live in Pekod. Pursue, kill and completely destroy them," declares the LORD. "Do everything I have commanded you.
JER|50|22|The noise of battle is in the land, the noise of great destruction!
JER|50|23|How broken and shattered is the hammer of the whole earth! How desolate is Babylon among the nations!
JER|50|24|I set a trap for you, O Babylon, and you were caught before you knew it; you were found and captured because you opposed the LORD.
JER|50|25|The LORD has opened his arsenal and brought out the weapons of his wrath, for the Sovereign LORD Almighty has work to do in the land of the Babylonians.
JER|50|26|Come against her from afar. Break open her granaries; pile her up like heaps of grain. Completely destroy her and leave her no remnant.
JER|50|27|Kill all her young bulls; let them go down to the slaughter! Woe to them! For their day has come, the time for them to be punished.
JER|50|28|Listen to the fugitives and refugees from Babylon declaring in Zion how the LORD our God has taken vengeance, vengeance for his temple.
JER|50|29|"Summon archers against Babylon, all those who draw the bow. Encamp all around her; let no one escape. Repay her for her deeds; do to her as she has done. For she has defied the LORD, the Holy One of Israel.
JER|50|30|Therefore, her young men will fall in the streets; all her soldiers will be silenced in that day," declares the LORD.
JER|50|31|"See, I am against you, O arrogant one," declares the Lord, the LORD Almighty, "for your day has come, the time for you to be punished.
JER|50|32|The arrogant one will stumble and fall and no one will help her up; I will kindle a fire in her towns that will consume all who are around her."
JER|50|33|This is what the LORD Almighty says: "The people of Israel are oppressed, and the people of Judah as well. All their captors hold them fast, refusing to let them go.
JER|50|34|Yet their Redeemer is strong; the LORD Almighty is his name. He will vigorously defend their cause so that he may bring rest to their land, but unrest to those who live in Babylon.
JER|50|35|"A sword against the Babylonians!" declares the LORD - "against those who live in Babylon and against her officials and wise men!
JER|50|36|A sword against her false prophets! They will become fools. A sword against her warriors! They will be filled with terror.
JER|50|37|A sword against her horses and chariots and all the foreigners in her ranks! They will become women. A sword against her treasures! They will be plundered.
JER|50|38|A drought on her waters! They will dry up. For it is a land of idols, idols that will go mad with terror.
JER|50|39|"So desert creatures and hyenas will live there, and there the owl will dwell. It will never again be inhabited or lived in from generation to generation.
JER|50|40|As God overthrew Sodom and Gomorrah along with their neighboring towns," declares the LORD, "so no one will live there; no man will dwell in it.
JER|50|41|"Look! An army is coming from the north; a great nation and many kings are being stirred up from the ends of the earth.
JER|50|42|They are armed with bows and spears; they are cruel and without mercy. They sound like the roaring sea as they ride on their horses; they come like men in battle formation to attack you, O Daughter of Babylon.
JER|50|43|The king of Babylon has heard reports about them, and his hands hang limp. Anguish has gripped him, pain like that of a woman in labor.
JER|50|44|Like a lion coming up from Jordan's thickets to a rich pastureland, I will chase Babylon from its land in an instant. Who is the chosen one I will appoint for this? Who is like me and who can challenge me? And what shepherd can stand against me?"
JER|50|45|Therefore, hear what the LORD has planned against Babylon, what he has purposed against the land of the Babylonians: The young of the flock will be dragged away; he will completely destroy their pasture because of them.
JER|50|46|At the sound of Babylon's capture the earth will tremble; its cry will resound among the nations.
JER|51|1|This is what the LORD says: "See, I will stir up the spirit of a destroyer against Babylon and the people of Leb Kamai.
JER|51|2|I will send foreigners to Babylon to winnow her and to devastate her land; they will oppose her on every side in the day of her disaster.
JER|51|3|Let not the archer string his bow, nor let him put on his armor. Do not spare her young men; completely destroy her army.
JER|51|4|They will fall down slain in Babylon, fatally wounded in her streets.
JER|51|5|For Israel and Judah have not been forsaken by their God, the LORD Almighty, though their land is full of guilt before the Holy One of Israel.
JER|51|6|"Flee from Babylon! Run for your lives! Do not be destroyed because of her sins. It is time for the LORD's vengeance; he will pay her what she deserves.
JER|51|7|Babylon was a gold cup in the LORD's hand; she made the whole earth drunk. The nations drank her wine; therefore they have now gone mad.
JER|51|8|Babylon will suddenly fall and be broken. Wail over her! Get balm for her pain; perhaps she can be healed.
JER|51|9|"'We would have healed Babylon, but she cannot be healed; let us leave her and each go to his own land, for her judgment reaches to the skies, it rises as high as the clouds.'
JER|51|10|"'The LORD has vindicated us; come, let us tell in Zion what the LORD our God has done.'
JER|51|11|"Sharpen the arrows, take up the shields! The LORD has stirred up the kings of the Medes, because his purpose is to destroy Babylon. The LORD will take vengeance, vengeance for his temple.
JER|51|12|Lift up a banner against the walls of Babylon! Reinforce the guard, station the watchmen, prepare an ambush! The LORD will carry out his purpose, his decree against the people of Babylon.
JER|51|13|You who live by many waters and are rich in treasures, your end has come, the time for you to be cut off.
JER|51|14|The LORD Almighty has sworn by himself: I will surely fill you with men, as with a swarm of locusts, and they will shout in triumph over you.
JER|51|15|"He made the earth by his power; he founded the world by his wisdom and stretched out the heavens by his understanding.
JER|51|16|When he thunders, the waters in the heavens roar; he makes clouds rise from the ends of the earth. He sends lightning with the rain and brings out the wind from his storehouses.
JER|51|17|"Every man is senseless and without knowledge; every goldsmith is shamed by his idols. His images are a fraud; they have no breath in them.
JER|51|18|They are worthless, the objects of mockery; when their judgment comes, they will perish.
JER|51|19|He who is the Portion of Jacob is not like these, for he is the Maker of all things, including the tribe of his inheritance- the LORD Almighty is his name.
JER|51|20|"You are my war club, my weapon for battle- with you I shatter nations, with you I destroy kingdoms,
JER|51|21|with you I shatter horse and rider, with you I shatter chariot and driver,
JER|51|22|with you I shatter man and woman, with you I shatter old man and youth, with you I shatter young man and maiden,
JER|51|23|with you I shatter shepherd and flock, with you I shatter farmer and oxen, with you I shatter governors and officials.
JER|51|24|"Before your eyes I will repay Babylon and all who live in Babylonia for all the wrong they have done in Zion," declares the LORD.
JER|51|25|"I am against you, O destroying mountain, you who destroy the whole earth," declares the LORD. "I will stretch out my hand against you, roll you off the cliffs, and make you a burned-out mountain.
JER|51|26|No rock will be taken from you for a cornerstone, nor any stone for a foundation, for you will be desolate forever," declares the LORD.
JER|51|27|"Lift up a banner in the land! Blow the trumpet among the nations! Prepare the nations for battle against her; summon against her these kingdoms: Ararat, Minni and Ashkenaz. Appoint a commander against her; send up horses like a swarm of locusts.
JER|51|28|Prepare the nations for battle against her- the kings of the Medes, their governors and all their officials, and all the countries they rule.
JER|51|29|The land trembles and writhes, for the LORD's purposes against Babylon stand- to lay waste the land of Babylon so that no one will live there.
JER|51|30|Babylon's warriors have stopped fighting; they remain in their strongholds. Their strength is exhausted; they have become like women. Her dwellings are set on fire; the bars of her gates are broken.
JER|51|31|One courier follows another and messenger follows messenger to announce to the king of Babylon that his entire city is captured,
JER|51|32|the river crossings seized, the marshes set on fire, and the soldiers terrified."
JER|51|33|This is what the LORD Almighty, the God of Israel, says: "The Daughter of Babylon is like a threshing floor at the time it is trampled; the time to harvest her will soon come."
JER|51|34|"Nebuchadnezzar king of Babylon has devoured us, he has thrown us into confusion, he has made us an empty jar. Like a serpent he has swallowed us and filled his stomach with our delicacies, and then has spewed us out.
JER|51|35|May the violence done to our flesh be upon Babylon," say the inhabitants of Zion. "May our blood be on those who live in Babylonia," says Jerusalem.
JER|51|36|Therefore, this is what the LORD says: "See, I will defend your cause and avenge you; I will dry up her sea and make her springs dry.
JER|51|37|Babylon will be a heap of ruins, a haunt of jackals, an object of horror and scorn, a place where no one lives.
JER|51|38|Her people all roar like young lions, they growl like lion cubs.
JER|51|39|But while they are aroused, I will set out a feast for them and make them drunk, so that they shout with laughter- then sleep forever and not awake," declares the LORD.
JER|51|40|"I will bring them down like lambs to the slaughter, like rams and goats.
JER|51|41|"How Sheshach will be captured, the boast of the whole earth seized! What a horror Babylon will be among the nations!
JER|51|42|The sea will rise over Babylon; its roaring waves will cover her.
JER|51|43|Her towns will be desolate, a dry and desert land, a land where no one lives, through which no man travels.
JER|51|44|I will punish Bel in Babylon and make him spew out what he has swallowed. The nations will no longer stream to him. And the wall of Babylon will fall.
JER|51|45|"Come out of her, my people! Run for your lives! Run from the fierce anger of the LORD.
JER|51|46|Do not lose heart or be afraid when rumors are heard in the land; one rumor comes this year, another the next, rumors of violence in the land and of ruler against ruler.
JER|51|47|For the time will surely come when I will punish the idols of Babylon; her whole land will be disgraced and her slain will all lie fallen within her.
JER|51|48|Then heaven and earth and all that is in them will shout for joy over Babylon, for out of the north destroyers will attack her," declares the LORD.
JER|51|49|"Babylon must fall because of Israel's slain, just as the slain in all the earth have fallen because of Babylon.
JER|51|50|You who have escaped the sword, leave and do not linger! Remember the LORD in a distant land, and think on Jerusalem."
JER|51|51|"We are disgraced, for we have been insulted and shame covers our faces, because foreigners have entered the holy places of the LORD's house."
JER|51|52|"But days are coming," declares the LORD, "when I will punish her idols, and throughout her land the wounded will groan.
JER|51|53|Even if Babylon reaches the sky and fortifies her lofty stronghold, I will send destroyers against her," declares the LORD.
JER|51|54|"The sound of a cry comes from Babylon, the sound of great destruction from the land of the Babylonians.
JER|51|55|The LORD will destroy Babylon; he will silence her noisy din. Waves of enemies will rage like great waters; the roar of their voices will resound.
JER|51|56|A destroyer will come against Babylon; her warriors will be captured, and their bows will be broken. For the LORD is a God of retribution; he will repay in full.
JER|51|57|I will make her officials and wise men drunk, her governors, officers and warriors as well; they will sleep forever and not awake," declares the King, whose name is the LORD Almighty.
JER|51|58|This is what the LORD Almighty says: "Babylon's thick wall will be leveled and her high gates set on fire; the peoples exhaust themselves for nothing, the nations' labor is only fuel for the flames."
JER|51|59|This is the message Jeremiah gave to the staff officer Seraiah son of Neriah, the son of Mahseiah, when he went to Babylon with Zedekiah king of Judah in the fourth year of his reign.
JER|51|60|Jeremiah had written on a scroll about all the disasters that would come upon Babylon-all that had been recorded concerning Babylon.
JER|51|61|He said to Seraiah, "When you get to Babylon, see that you read all these words aloud.
JER|51|62|Then say, 'O LORD, you have said you will destroy this place, so that neither man nor animal will live in it; it will be desolate forever.'
JER|51|63|When you finish reading this scroll, tie a stone to it and throw it into the Euphrates.
JER|51|64|Then say, 'So will Babylon sink to rise no more because of the disaster I will bring upon her. And her people will fall.'" The words of Jeremiah end here.
JER|52|1|Zedekiah was twenty-one years old when he became king, and he reigned in Jerusalem eleven years. His mother's name was Hamutal daughter of Jeremiah; she was from Libnah.
JER|52|2|He did evil in the eyes of the LORD, just as Jehoiakim had done.
JER|52|3|It was because of the LORD's anger that all this happened to Jerusalem and Judah, and in the end he thrust them from his presence. Now Zedekiah rebelled against the king of Babylon.
JER|52|4|So in the ninth year of Zedekiah's reign, on the tenth day of the tenth month, Nebuchadnezzar king of Babylon marched against Jerusalem with his whole army. They camped outside the city and built siege works all around it.
JER|52|5|The city was kept under siege until the eleventh year of King Zedekiah.
JER|52|6|By the ninth day of the fourth month the famine in the city had become so severe that there was no food for the people to eat.
JER|52|7|Then the city wall was broken through, and the whole army fled. They left the city at night through the gate between the two walls near the king's garden, though the Babylonians were surrounding the city. They fled toward the Arabah,
JER|52|8|but the Babylonian army pursued King Zedekiah and overtook him in the plains of Jericho. All his soldiers were separated from him and scattered,
JER|52|9|and he was captured. He was taken to the king of Babylon at Riblah in the land of Hamath, where he pronounced sentence on him.
JER|52|10|There at Riblah the king of Babylon slaughtered the sons of Zedekiah before his eyes; he also killed all the officials of Judah.
JER|52|11|Then he put out Zedekiah's eyes, bound him with bronze shackles and took him to Babylon, where he put him in prison till the day of his death.
JER|52|12|On the tenth day of the fifth month, in the nineteenth year of Nebuchadnezzar king of Babylon, Nebuzaradan commander of the imperial guard, who served the king of Babylon, came to Jerusalem.
JER|52|13|He set fire to the temple of the LORD, the royal palace and all the houses of Jerusalem. Every important building he burned down.
JER|52|14|The whole Babylonian army under the commander of the imperial guard broke down all the walls around Jerusalem.
JER|52|15|Nebuzaradan the commander of the guard carried into exile some of the poorest people and those who remained in the city, along with the rest of the craftsmen and those who had gone over to the king of Babylon.
JER|52|16|But Nebuzaradan left behind the rest of the poorest people of the land to work the vineyards and fields.
JER|52|17|The Babylonians broke up the bronze pillars, the movable stands and the bronze Sea that were at the temple of the LORD and they carried all the bronze to Babylon.
JER|52|18|They also took away the pots, shovels, wick trimmers, sprinkling bowls, dishes and all the bronze articles used in the temple service.
JER|52|19|The commander of the imperial guard took away the basins, censers, sprinkling bowls, pots, lampstands, dishes and bowls used for drink offerings-all that were made of pure gold or silver.
JER|52|20|The bronze from the two pillars, the Sea and the twelve bronze bulls under it, and the movable stands, which King Solomon had made for the temple of the LORD, was more than could be weighed.
JER|52|21|Each of the pillars was eighteen cubits high and twelve cubits in circumference; each was four fingers thick, and hollow.
JER|52|22|The bronze capital on top of the one pillar was five cubits high and was decorated with a network and pomegranates of bronze all around. The other pillar, with its pomegranates, was similar.
JER|52|23|There were ninety-six pomegranates on the sides; the total number of pomegranates above the surrounding network was a hundred.
JER|52|24|The commander of the guard took as prisoners Seraiah the chief priest, Zephaniah the priest next in rank and the three doorkeepers.
JER|52|25|Of those still in the city, he took the officer in charge of the fighting men, and seven royal advisers. He also took the secretary who was chief officer in charge of conscripting the people of the land and sixty of his men who were found in the city.
JER|52|26|Nebuzaradan the commander took them all and brought them to the king of Babylon at Riblah.
JER|52|27|There at Riblah, in the land of Hamath, the king had them executed. So Judah went into captivity, away from her land.
JER|52|28|This is the number of the people Nebuchadnezzar carried into exile: in the seventh year, 3,023 Jews;
JER|52|29|in Nebuchadnezzar's eighteenth year, 832 people from Jerusalem;
JER|52|30|in his twenty-third year, 745 Jews taken into exile by Nebuzaradan the commander of the imperial guard. There were 4,600 people in all.
JER|52|31|In the thirty-seventh year of the exile of Jehoiachin king of Judah, in the year Evil-Merodach became king of Babylon, he released Jehoiachin king of Judah and freed him from prison on the twenty-fifth day of the twelfth month.
JER|52|32|He spoke kindly to him and gave him a seat of honor higher than those of the other kings who were with him in Babylon.
JER|52|33|So Jehoiachin put aside his prison clothes and for the rest of his life ate regularly at the king's table.
JER|52|34|Day by day the king of Babylon gave Jehoiachin a regular allowance as long as he lived, till the day of his death.
