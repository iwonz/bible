AMOS|1|1|Слова Амоса, одного из пастухов Фекойских, которые он [слышал] в видении об Израиле во дни Озии, царя Иудейского, и во дни Иеровоама, сына Иоасова, царя Израильского, за два года перед землетрясением.
AMOS|1|2|И сказал он: Господь возгремит с Сиона и даст глас Свой из Иерусалима, и восплачут хижины пастухов, и иссохнет вершина Кармила.
AMOS|1|3|Так говорит Господь: за три преступления Дамаска и за четыре не пощажу его, потому что они молотили Галаад железными молотилами.
AMOS|1|4|И пошлю огонь на дом Азаила, и пожрет он чертоги Венадада.
AMOS|1|5|И сокрушу затворы Дамаска, и истреблю жителей долины Авен и держащего скипетр – из дома Еденова, и пойдет народ Арамейский в плен в Кир, говорит Господь.
AMOS|1|6|Так говорит Господь: за три преступления Газы и за четыре не пощажу ее, потому что они вывели всех в плен, чтобы предать их Едому.
AMOS|1|7|И пошлю огонь в стены Газы, – и пожрет чертоги ее.
AMOS|1|8|И истреблю жителей Азота и держащего скипетр в Аскалоне, и обращу руку Мою на Екрон, и погибнет остаток Филистимлян, говорит Господь Бог.
AMOS|1|9|Так говорит Господь: за три преступления Тира и за четыре не пощажу его, потому что они передали всех пленных Едому и не вспомнили братского союза.
AMOS|1|10|Пошлю огонь в стены Тира, и пожрет чертоги его.
AMOS|1|11|Так говорит Господь: за три преступления Едома и за четыре не пощажу его, потому что он преследовал брата своего мечом, подавил чувства родства, свирепствовал постоянно во гневе своем и всегда сохранял ярость свою.
AMOS|1|12|И пошлю огонь на Феман, и пожрет чертоги Восора.
AMOS|1|13|Так говорит Господь: за три преступления сынов Аммоновых и за четыре не пощажу их, потому что они рассекали беременных в Галааде, чтобы расширить пределы свои.
AMOS|1|14|И запалю огонь в стенах Раввы, и пожрет чертоги ее, среди крика в день брани, с вихрем в день бури.
AMOS|1|15|И пойдет царь их в плен, он и князья его вместе с ним, говорит Господь.
AMOS|2|1|Так говорит Господь: за три преступления Моава и за четыре не пощажу его, потому что он пережег кости царя Едомского в известь.
AMOS|2|2|И пошлю огонь на Моава, и пожрет чертоги Кериофа, и погибнет Моав среди разгрома с шумом, при звуке трубы.
AMOS|2|3|Истреблю судью из среды его и умерщвлю всех князей его вместе с ним, говорит Господь.
AMOS|2|4|Так говорит Господь: за три преступления Иуды и за четыре не пощажу его, потому что отвергли закон Господень и постановлений Его не сохранили, и идолы их, вслед которых ходили отцы их, совратили их с пути.
AMOS|2|5|И пошлю огонь на Иуду, и пожрет чертоги Иерусалима.
AMOS|2|6|Так говорит Господь: за три преступления Израиля и за четыре не пощажу его, потому что продают правого за серебро и бедного – за пару сандалий.
AMOS|2|7|Жаждут, чтобы прах земной был на голове бедных, и путь кротких извращают; даже отец и сын ходят к одной женщине, чтобы бесславить святое имя Мое.
AMOS|2|8|На одеждах, взятых в залог, возлежат при всяком жертвеннике, и вино, [взыскиваемое] с обвиненных, пьют в доме богов своих.
AMOS|2|9|А Я истребил перед лицем их Аморрея, которого высота была как высота кедра и который был крепок как дуб; Я истребил плод его вверху и корни его внизу.
AMOS|2|10|Вас же Я вывел из земли Египетской и водил вас в пустыне сорок лет, чтобы вам наследовать землю Аморрейскую.
AMOS|2|11|Из сыновей ваших Я избирал в пророки и из юношей ваших – в назореи; не так ли это, сыны Израиля? говорит Господь.
AMOS|2|12|А вы назореев поили вином и пророкам приказывали, говоря: "не пророчествуйте".
AMOS|2|13|Вот, Я придавлю вас, как давит колесница, нагруженная снопами, –
AMOS|2|14|и у проворного не станет силы бежать, и крепкий не удержит крепости своей, и храбрый не спасет своей жизни,
AMOS|2|15|ни стреляющий из лука не устоит, ни скороход не убежит, ни сидящий на коне не спасет своей жизни.
AMOS|2|16|И самый отважный из храбрых убежит нагой в тот день, говорит Господь.
AMOS|3|1|Слушайте слово сие, которое Господь изрек на вас, сыны Израилевы, на все племя, которое вывел Я из земли Египетской, говоря:
AMOS|3|2|только вас признал Я из всех племен земли, потому и взыщу с вас за все беззакония ваши.
AMOS|3|3|Пойдут ли двое вместе, не сговорившись между собою?
AMOS|3|4|Ревет ли лев в лесу, когда нет перед ним добычи? подает ли свой голос львенок из логовища своего, когда он ничего не поймал?
AMOS|3|5|Попадет ли птица в петлю на земле, когда силка нет для нее? Поднимется ли с земли петля, когда ничего не попало в нее?
AMOS|3|6|Трубит ли в городе труба, – и народ не испугался бы? Бывает ли в городе бедствие, которое не Господь попустил бы?
AMOS|3|7|Ибо Господь Бог ничего не делает, не открыв Своей тайны рабам Своим, пророкам.
AMOS|3|8|Лев начал рыкать, – кто не содрогнется? Господь Бог сказал, – кто не будет пророчествовать?
AMOS|3|9|Провозгласите на кровлях в Азоте и на кровлях в земле Египетской и скажите: соберитесь на горы Самарии и посмотрите на великое бесчинство в ней и на притеснения среди нее.
AMOS|3|10|Они не умеют поступать справедливо, говорит Господь: насилием и грабежом собирают сокровища в чертоги свои.
AMOS|3|11|Посему так говорит Господь Бог: вот неприятель, и притом вокруг всей земли! он низложит могущество твое, и ограблены будут чертоги твои.
AMOS|3|12|Так говорит Господь: как [иногда] пастух исторгает из пасти львиной две голени или часть уха, так спасены будут сыны Израилевы, сидящие в Самарии в углу постели и в Дамаске на ложе.
AMOS|3|13|Слушайте и засвидетельствуйте дому Иакова, говорит Господь Бог, Бог Саваоф.
AMOS|3|14|Ибо в тот день, когда Я взыщу с Израиля за преступления его, взыщу и за жертвенники в Вефиле, и отсечены будут роги алтаря, и падут на землю.
AMOS|3|15|И поражу дом зимний вместе с домом летним, и исчезнут домы с украшениями из слоновой кости, и не станет многих домов, говорит Господь.
AMOS|4|1|Слушайте слово сие, телицы Васанские, которые на горе Самарийской, вы, притесняющие бедных, угнетающие нищих, говорящие господам своим: "подавай, и мы будем пить!"
AMOS|4|2|Клялся Господь Бог святостью Своею, что вот, придут на вас дни, когда повлекут вас крюками и остальных ваших удами.
AMOS|4|3|И сквозь проломы стен выйдете, каждая, как случится, и бросите все убранство чертогов, говорит Господь.
AMOS|4|4|Идите в Вефиль – и грешите, в Галгал – и умножайте преступления; приносите жертвы ваши каждое утро, десятины ваши хотя через каждые три дня.
AMOS|4|5|Приносите в жертву благодарения квасное, провозглашайте о добровольных приношениях ваших и разглашайте о них, ибо это вы любите, сыны Израилевы, говорит Господь Бог.
AMOS|4|6|За то и дал Я вам голые зубы во всех городах ваших и недостаток хлеба во всех селениях ваших; но вы не обратились ко Мне, говорит Господь.
AMOS|4|7|И удерживал от вас дождь за три месяца до жатвы; проливал дождь на один город, а на другой город не проливал дождя; один участок напояем был дождем, а другой, не окропленный дождем, засыхал.
AMOS|4|8|И сходились два–три города в один город, чтобы напиться воды, и не могли досыта напиться; но и тогда вы не обратились ко Мне, говорит Господь.
AMOS|4|9|Я поражал вас ржою и блеклостью хлеба; множество садов ваших и виноградников ваших, и смоковниц ваших, и маслин ваших пожирала гусеница, – и при всем том вы не обратились ко Мне, говорит Господь.
AMOS|4|10|Посылал Я на вас моровую язву, подобную Египетской, убивал мечом юношей ваших, отводя коней в плен, так что смрад от станов ваших поднимался в ноздри ваши; и при всем том вы не обратились ко Мне, говорит Господь.
AMOS|4|11|Производил Я среди вас разрушения, как разрушил Бог Содом и Гоморру, и вы были выхвачены, как головня из огня, – и при всем том вы не обратились ко Мне, говорит Господь.
AMOS|4|12|Посему так поступлю Я с тобою, Израиль; и как Я так поступлю с тобою, то приготовься к сретению Бога твоего, Израиль,
AMOS|4|13|ибо вот Он, Который образует горы, и творит ветер, и объявляет человеку намерения его, утренний свет обращает в мрак, и шествует превыше земли; Господь Бог Саваоф – имя Ему.
AMOS|5|1|Слушайте это слово, в котором я подниму плач о вас, дом Израилев.
AMOS|5|2|Упала, не встает более дева Израилева! повержена на земле своей, и некому поднять ее.
AMOS|5|3|Ибо так говорит Господь Бог: город, выступавший тысячею, останется только с сотнею, и выступавший сотнею, останется с десятком у дома Израилева.
AMOS|5|4|Ибо так говорит Господь дому Израилеву: взыщите Меня, и будете живы.
AMOS|5|5|Не ищите Вефиля и не ходите в Галгал, и в Вирсавию не странствуйте, ибо Галгал весь пойдет в плен и Вефиль обратится в ничто.
AMOS|5|6|Взыщите Господа, и будете живы, чтобы Он не устремился на дом Иосифов как огонь, который пожрет его, и некому будет погасить его в Вефиле.
AMOS|5|7|О, вы, которые суд превращаете в отраву и правду повергаете на землю!
AMOS|5|8|Кто сотворил семизвездие и Орион, и претворяет смертную тень в ясное утро, а день делает темным как ночь, призывает воды морские и разливает их по лицу земли? – Господь имя Ему!
AMOS|5|9|Он укрепляет опустошителя против сильного, и опустошитель входит в крепость.
AMOS|5|10|А они ненавидят обличающего в воротах и гнушаются тем, кто говорит правду.
AMOS|5|11|Итак за то, что вы попираете бедного и берете от него подарки хлебом, вы построите домы из тесаных камней, но жить не будете в них; разведете прекрасные виноградники, а вино из них не будете пить.
AMOS|5|12|Ибо Я знаю, как многочисленны преступления ваши и как тяжки грехи ваши: вы враги правого, берете взятки и извращаете в суде дела бедных.
AMOS|5|13|Поэтому разумный безмолвствует в это время, ибо злое это время.
AMOS|5|14|Ищите добра, а не зла, чтобы вам остаться в живых, – и тогда Господь Бог Саваоф будет с вами, как вы говорите.
AMOS|5|15|Возненавидьте зло и возлюбите добро, и восстановите у ворот правосудие; может быть, Господь Бог Саваоф помилует остаток Иосифов.
AMOS|5|16|Посему так говорит Господь Бог Саваоф, Вседержитель: на всех улицах будет плач, и на всех дорогах будут восклицать: "увы, увы!", и призовут земледельца сетовать и искусных в плачевных песнях – плакать,
AMOS|5|17|и во всех виноградниках будет плач, ибо Я пройду среди тебя, говорит Господь.
AMOS|5|18|Горе желающим дня Господня! для чего вам этот день Господень? он тьма, а не свет,
AMOS|5|19|то же, как если бы кто убежал от льва, и попался бы ему навстречу медведь, или если бы пришел домой и оперся рукою о стену, и змея ужалила бы его.
AMOS|5|20|Разве день Господень не мрак, а свет? он тьма, и нет в нем сияния.
AMOS|5|21|Ненавижу, отвергаю праздники ваши и не обоняю жертв во время торжественных собраний ваших.
AMOS|5|22|Если вознесете Мне всесожжение и хлебное приношение, Я не приму их и не призрю на благодарственную жертву из тучных тельцов ваших.
AMOS|5|23|Удали от Меня шум песней твоих, ибо звуков гуслей твоих Я не буду слушать.
AMOS|5|24|Пусть, как вода, течет суд, и правда – как сильный поток!
AMOS|5|25|Приносили ли вы Мне жертвы и хлебные дары в пустыне в течение сорока лет, дом Израилев?
AMOS|5|26|Вы носили скинию Молохову и звезду бога вашего Ремфана, изображения, которые вы сделали для себя.
AMOS|5|27|За то Я переселю вас за Дамаск, говорит Господь; Бог Саваоф – имя Ему!
AMOS|6|1|Горе беспечным на Сионе и надеющимся на гору Самарийскую именитым первенствующего народа, к которым приходит дом Израиля!
AMOS|6|2|Пройдите в Калне и посмотрите, оттуда перейдите в Емаф великий и спуститесь в Геф Филистимский: не лучше ли они сих царств? не обширнее ли пределы их пределов ваших?
AMOS|6|3|Вы, которые день бедствия считаете далеким и приближаете торжество насилия, –
AMOS|6|4|вы, которые лежите на ложах из слоновой кости и нежитесь на постелях ваших, едите лучших овнов из стада и тельцов с тучного пастбища,
AMOS|6|5|поете под звуки гуслей, думая, что владеете музыкальным орудием, как Давид,
AMOS|6|6|пьете из чаш вино, мажетесь наилучшими мастями, и не болезнуете о бедствии Иосифа!
AMOS|6|7|За то ныне пойдут они в плен во главе пленных, и кончится ликование изнеженных.
AMOS|6|8|Клянется Господь Бог Самим Собою, и так говорит Господь Бог Саваоф: гнушаюсь высокомерием Иакова и ненавижу чертоги его, и предам город и все, что наполняет его.
AMOS|6|9|И будет: если в каком доме останется десять человек, то умрут и они,
AMOS|6|10|и возьмет их родственник их или сожигатель, чтобы вынести кости их из дома, и скажет находящемуся при доме: есть ли еще у тебя кто? Тот ответит: нет никого. И скажет сей: молчи! ибо нельзя упоминать имени Господня.
AMOS|6|11|Ибо вот, Господь даст повеление и поразит большие дома расселинами, а малые дома – трещинами.
AMOS|6|12|Бегают ли кони по скале? можно ли распахивать ее волами? Вы между тем суд превращаете в яд и плод правды в горечь;
AMOS|6|13|вы, которые восхищаетесь ничтожными вещами и говорите: "не своею ли силою мы приобрели себе могущество?"
AMOS|6|14|Вот Я, говорит Господь Бог Саваоф, воздвигну народ против вас, дом Израилев, и будут теснить вас от входа в Емаф до потока в пустыне.
AMOS|7|1|Такое видение открыл мне Господь Бог: вот, Он создал саранчу в начале произрастания поздней травы, и это была трава после царского покоса.
AMOS|7|2|И было, когда она окончила есть траву на земле, я сказал: Господи Боже! пощади; как устоит Иаков? он очень мал.
AMOS|7|3|И пожалел Господь о том; "не будет сего", сказал Господь.
AMOS|7|4|Такое видение открыл мне Господь Бог: вот, Господь Бог произвел для суда огонь, – и он пожрал великую пучину, пожрал и часть земли.
AMOS|7|5|И сказал я: Господи Боже! останови; как устоит Иаков? он очень мал.
AMOS|7|6|И пожалел Господь о том; "и этого не будет", сказал Господь Бог.
AMOS|7|7|Такое видение открыл Он мне: вот, Господь стоял на отвесной стене, и в руке у Него свинцовый отвес.
AMOS|7|8|И сказал мне Господь: что ты видишь, Амос? Я ответил: отвес. И Господь сказал: вот, положу отвес среди народа Моего, Израиля; не буду более прощать ему.
AMOS|7|9|И опустошены будут [жертвенные] высоты Исааковы, и разрушены будут святилища Израилевы, и восстану с мечом против дома Иеровоамова.
AMOS|7|10|И послал Амасия, священник Вефильский, к Иеровоаму, царю Израильскому, сказать: Амос производит возмущение против тебя среди дома Израилева; земля не может терпеть всех слов его.
AMOS|7|11|Ибо так говорит Амос: "от меча умрет Иеровоам, а Израиль непременно отведен будет пленным из земли своей".
AMOS|7|12|И сказал Амасия Амосу: провидец! пойди и удались в землю Иудину; там ешь хлеб, и там пророчествуй,
AMOS|7|13|а в Вефиле больше не пророчествуй, ибо он святыня царя и дом царский.
AMOS|7|14|И отвечал Амос и сказал Амасии: я не пророк и не сын пророка; я был пастух и собирал сикоморы.
AMOS|7|15|Но Господь взял меня от овец и сказал мне Господь: "иди, пророчествуй к народу Моему, Израилю".
AMOS|7|16|Теперь выслушай слово Господне. Ты говоришь: "не пророчествуй на Израиля и не произноси слов на дом Исааков".
AMOS|7|17|За это, вот что говорит Господь: жена твоя будет обесчещена в городе, сыновья и дочери твои падут от меча, земля твоя будет разделена межевою вервью, а ты умрешь в земле нечистой, и Израиль непременно выведен будет из земли своей.
AMOS|8|1|Такое видение открыл мне Господь Бог: вот корзина со спелыми плодами.
AMOS|8|2|И сказал Он: что ты видишь, Амос? Я ответил: корзину со спелыми плодами. Тогда Господь сказал мне: приспел конец народу Моему, Израилю: не буду более прощать ему.
AMOS|8|3|Песни чертога в тот день обратятся в рыдание, говорит Господь Бог; много будет трупов, на всяком месте будут бросать их молча.
AMOS|8|4|Выслушайте это, алчущие поглотить бедных и погубить нищих, –
AMOS|8|5|вы, которые говорите: "когда–то пройдет новолуние, чтобы нам продавать хлеб, и суббота, чтобы открыть житницы, уменьшить меру, увеличить цену сикля и обманывать неверными весами,
AMOS|8|6|чтобы покупать неимущих за серебро и бедных за пару обуви, а высевки из хлеба продавать".
AMOS|8|7|Клялся Господь славою Иакова: поистине во веки не забуду ни одного из дел их!
AMOS|8|8|Не поколеблется ли от этого земля, и не восплачет ли каждый, живущий на ней? Взволнуется вся она, как река, и будет подниматься и опускаться, как река Египетская.
AMOS|8|9|И будет в тот день, говорит Господь Бог: произведу закат солнца в полдень и омрачу землю среди светлого дня.
AMOS|8|10|И обращу праздники ваши в сетование и все песни ваши в плач, и возложу на все чресла вретище и плешь на всякую голову; и произведу [в] [стране] плач, как о единственном сыне, и конец ее будет – как горький день.
AMOS|8|11|Вот наступают дни, говорит Господь Бог, когда Я пошлю на землю голод, – не голод хлеба, не жажду воды, но жажду слышания слов Господних.
AMOS|8|12|И будут ходить от моря до моря и скитаться от севера к востоку, ища слова Господня, и не найдут его.
AMOS|8|13|В тот день истаявать будут от жажды красивые девы и юноши,
AMOS|8|14|которые клянутся грехом Самарийским и говорят: "жив бог твой, Дан! и жив путь в Вирсавию!" – Они падут и уже не встанут.
AMOS|9|1|Видел я Господа стоящим над жертвенником, и Он сказал: ударь в притолоку над воротами, чтобы потряслись косяки, и обрушь их на головы всех их, остальных же из них Я поражу мечом: не убежит у них никто бегущий и не спасется из них никто, желающий спастись.
AMOS|9|2|Хотя бы они зарылись в преисподнюю, и оттуда рука Моя возьмет их; хотя бы взошли на небо, и оттуда свергну их.
AMOS|9|3|И хотя бы они скрылись на вершине Кармила, и там отыщу и возьму их; хотя бы сокрылись от очей Моих на дне моря, и там повелю морскому змею уязвить их.
AMOS|9|4|И если пойдут в плен впереди врагов своих, то повелю мечу и там убить их. Обращу на них очи Мои на беду им, а не во благо.
AMOS|9|5|Ибо Господь Бог Саваоф коснется земли, – и она растает, и восплачут все живущие на ней; и поднимется вся она как река, и опустится как река Египетская.
AMOS|9|6|Он устроил горние чертоги Свои на небесах и свод Свой утвердил на земле, призывает воды морские, и изливает их по лицу земли; Господь имя Ему.
AMOS|9|7|Не таковы ли, как сыны Ефиоплян, и вы для Меня, сыны Израилевы? говорит Господь. Не Я ли вывел Израиля из земли Египетской и Филистимлян – из Кафтора, и Арамлян – из Кира?
AMOS|9|8|Вот, очи Господа Бога – на грешное царство, и Я истреблю его с лица земли; но дом Иакова не совсем истреблю, говорит Господь.
AMOS|9|9|Ибо вот, Я повелю и рассыплю дом Израилев по всем народам, как рассыпают зерна в решете, и ни одно не падает на землю.
AMOS|9|10|От меча умрут все грешники из народа Моего, которые говорят: "не постигнет нас и не придет к нам это бедствие!"
AMOS|9|11|В тот день Я восстановлю скинию Давидову падшую, заделаю трещины в ней и разрушенное восстановлю, и устрою ее, как в дни древние,
AMOS|9|12|чтобы они овладели остатком Едома и всеми народами, между которыми возвестится имя Мое, говорит Господь, творящий все сие.
AMOS|9|13|Вот, наступят дни, говорит Господь, когда пахарь застанет еще жнеца, а топчущий виноград – сеятеля; и горы источать будут виноградный сок, и все холмы потекут.
AMOS|9|14|И возвращу из плена народ Мой, Израиля, и застроят опустевшие города и поселятся в них, насадят виноградники и будут пить вино из них, разведут сады и станут есть плоды из них.
AMOS|9|15|И водворю их на земле их, и они не будут более исторгаемы из земли своей, которую Я дал им, говорит Господь Бог твой.
