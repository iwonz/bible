TITUS|1|1|上帝的僕人、耶穌基督的使徒 保羅 ，為了使上帝的選民信從與認識合乎敬虔的真理—
TITUS|1|2|這真理是在盼望那無謊言的上帝在萬古之先所應許的永生，
TITUS|1|3|到了適當的時機，藉著傳揚福音，把他的道顯明了；這傳揚的責任是按著我們的救主上帝的命令交託給我的—
TITUS|1|4|我寫信給在共同的信仰上作我真兒子的 提多 。願恩惠、平安 從父上帝和我們的救主基督耶穌歸給你！
TITUS|1|5|我從前把你留在 克里特 ，是要你將那沒有辦完的事都辦妥，又照我所吩咐你的，在各城設立長老。
TITUS|1|6|若有無可指責的人，只作一個婦人的丈夫，兒女也是信主的，沒有人告他們放蕩，不受約束，就可以設立。
TITUS|1|7|監督既然是上帝的管家，必須無可指責、不自負、不暴躁、不酗酒、不好鬥、不貪財；
TITUS|1|8|卻要樂意接待外人、好善、克己、正直、聖潔、節制，
TITUS|1|9|堅守合乎教義的可靠之道，就能將健全的教導勸勉人，又能駁倒爭辯的人。
TITUS|1|10|因為也有許多人不受約束，說空話欺哄人，尤其是那些奉割禮的人。
TITUS|1|11|這些人的口必須堵住，因為他們貪不義之財，將不該教導的事教導人，敗壞人的全家。
TITUS|1|12|克里特 人中有一個本地的先知說：「 克里特 人常說謊話，是惡獸，貪吃懶做。」
TITUS|1|13|這個見證是真的。為這緣故，你要嚴厲地責備他們，使他們在信仰上健全。
TITUS|1|14|不要聽 猶太 人無稽的傳說和背棄真理之人的命令。
TITUS|1|15|在潔淨的人，凡物都潔淨；在污穢不信的人，甚麼都不潔淨，連心地和天良也都污穢了。
TITUS|1|16|他們宣稱認識上帝，卻在行為上否認他；他們是可憎惡的，是悖逆的，不配做任何好事。
TITUS|2|1|至於你，你所講的總要合乎那健全的教導。
TITUS|2|2|勸老年人要有節制、端正、克己，在信心、愛心、耐心上都要健全。
TITUS|2|3|又要勸年長的婦女在操守上恭正，不說讒言，不作酒的奴隸，用善道教導人，
TITUS|2|4|好指教年輕的婦女愛丈夫，愛兒女，
TITUS|2|5|克己，貞潔，理家，善良，順服自己的丈夫，免得上帝的道被毀謗。
TITUS|2|6|同樣，要勸年輕人凡事克己。
TITUS|2|7|你要顯出自己是好行為的榜樣，在教導上要正直、莊重，
TITUS|2|8|言語健全，無可指責，使那反對的人，因說不出我們有甚麼不好而自覺羞愧。
TITUS|2|9|要勸僕人順服自己的主人，凡事討他的喜悅，不可頂撞他，
TITUS|2|10|不可私竊財物；要凡事顯出完美的忠誠，好事事都能榮耀我們救主上帝的教導。
TITUS|2|11|因為，上帝救眾人的恩典已經顯明出來，
TITUS|2|12|訓練我們除去不敬虔的心和世俗的情慾，在今世過克己、正直、敬虔的生活，
TITUS|2|13|等候福樂的盼望，並等候至大的上帝和我們的救主 耶穌基督的榮耀顯現。
TITUS|2|14|他為我們的緣故捨己，為了要贖我們脫離一切罪惡，又潔淨我們作他自己的子民，熱心為善。
TITUS|2|15|這些事你要講明，要充分運用你的職權勸勉人，責備人。不要讓任何人輕看你。
TITUS|3|1|你要提醒眾人，叫他們順服執政的、掌權的，要服從，預備行各樣善事。
TITUS|3|2|不要毀謗，不要爭吵，要和氣，對眾人總要顯出溫柔。
TITUS|3|3|我們從前也是無知、悖逆、受迷惑，作各樣私慾和宴樂的奴隸，在惡毒、嫉妒中度日，是可恨的，而且彼此相恨。
TITUS|3|4|但到了我們救主上帝的恩慈和慈愛顯明的時候，
TITUS|3|5|他救了我們，並不是因我們自己所行的義，而是照他的憐憫，藉著重生的洗和聖靈的更新。
TITUS|3|6|聖靈就是上帝藉著我們的救主耶穌基督厚厚地澆灌在我們身上的，
TITUS|3|7|好讓我們因他的恩得稱為義，可以憑著永生的盼望成為後嗣 。
TITUS|3|8|這話是可信的。 我願你堅持這些事，使那些已信上帝的人留心行善 。這都是美好且對人有益的。
TITUS|3|9|要遠避愚拙的辯論、家譜、紛爭和因律法而起的爭辯，因為這都是虛妄無益的。
TITUS|3|10|分門結黨的人，警戒過一兩次後就要拒絕跟他來往；
TITUS|3|11|因為你知道這樣的人已經背道，常常犯罪，自己定自己的罪了。
TITUS|3|12|我打發 亞提馬 或 推基古 到你那裏去的時候，你要趕緊往 尼哥坡里 來見我，因為我已經決定在那裏過冬。
TITUS|3|13|你要趕緊給 西納 律師和 亞波羅 送行，讓他們沒有缺乏。
TITUS|3|14|我們的人也該學習行善，幫助有迫切需要的人，這樣才不會不結果子。
TITUS|3|15|跟我同在一起的人都向你問安。請代向在信仰上愛我們的人問安。願恩惠與你們眾人同在！
